VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tt_tinyQV
  CLASS BLOCK ;
  FOREIGN tt_um_tt_tinyQV ;
  ORIGIN 0.000 0.000 ;
  SIZE 1071.840 BY 710.640 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 21.580 3.560 23.780 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 60.450 3.560 62.650 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 99.320 3.560 101.520 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 138.190 3.560 140.390 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 177.060 3.560 179.260 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 215.930 3.560 218.130 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 254.800 3.560 257.000 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 293.670 3.560 295.870 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 332.540 3.560 334.740 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 371.410 3.560 373.610 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 410.280 3.560 412.480 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 449.150 3.560 451.350 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 488.020 3.560 490.220 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 526.890 3.560 529.090 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 565.760 3.560 567.960 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 604.630 3.560 606.830 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 643.500 3.560 645.700 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 682.370 3.560 684.570 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 721.240 3.560 723.440 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 760.110 3.560 762.310 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 798.980 3.560 801.180 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 837.850 3.560 840.050 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 876.720 3.560 878.920 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 915.590 3.560 917.790 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 954.460 3.560 956.660 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 993.330 3.560 995.530 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1032.200 3.560 1034.400 707.080 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 15.380 3.560 17.580 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 54.250 3.560 56.450 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 93.120 3.560 95.320 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 131.990 3.560 134.190 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 170.860 3.560 173.060 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 209.730 3.560 211.930 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 248.600 3.560 250.800 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 287.470 3.560 289.670 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 326.340 3.560 328.540 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 365.210 3.560 367.410 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 404.080 3.560 406.280 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 442.950 3.560 445.150 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 481.820 3.560 484.020 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 520.690 3.560 522.890 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 559.560 3.560 561.760 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 598.430 3.560 600.630 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 637.300 3.560 639.500 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 676.170 3.560 678.370 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 715.040 3.560 717.240 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 753.910 3.560 756.110 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 792.780 3.560 794.980 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 831.650 3.560 833.850 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 870.520 3.560 872.720 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 909.390 3.560 911.590 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 948.260 3.560 950.460 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 987.130 3.560 989.330 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1026.000 3.560 1028.200 707.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1064.870 3.560 1067.070 707.080 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.076800 ;
    ANTENNADIFFAREA 12.092400 ;
    PORT
      LAYER Metal5 ;
        RECT 187.050 709.640 187.350 710.640 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 190.890 709.640 191.190 710.640 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal5 ;
        RECT 183.210 709.640 183.510 710.640 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal5 ;
        RECT 179.370 709.640 179.670 710.640 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal5 ;
        RECT 175.530 709.640 175.830 710.640 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal5 ;
        RECT 171.690 709.640 171.990 710.640 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.038400 ;
    ANTENNADIFFAREA 6.046200 ;
    PORT
      LAYER Metal5 ;
        RECT 167.850 709.640 168.150 710.640 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal5 ;
        RECT 164.010 709.640 164.310 710.640 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal5 ;
        RECT 160.170 709.640 160.470 710.640 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal5 ;
        RECT 156.330 709.640 156.630 710.640 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal5 ;
        RECT 152.490 709.640 152.790 710.640 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 148.650 709.640 148.950 710.640 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal5 ;
        RECT 144.810 709.640 145.110 710.640 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal5 ;
        RECT 140.970 709.640 141.270 710.640 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 137.130 709.640 137.430 710.640 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal5 ;
        RECT 133.290 709.640 133.590 710.640 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal5 ;
        RECT 129.450 709.640 129.750 710.640 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 125.610 709.640 125.910 710.640 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 121.770 709.640 122.070 710.640 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.413600 ;
    PORT
      LAYER Metal5 ;
        RECT 56.490 709.640 56.790 710.640 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.413600 ;
    PORT
      LAYER Metal5 ;
        RECT 52.650 709.640 52.950 710.640 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.413600 ;
    PORT
      LAYER Metal5 ;
        RECT 48.810 709.640 49.110 710.640 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.413600 ;
    PORT
      LAYER Metal5 ;
        RECT 44.970 709.640 45.270 710.640 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.413600 ;
    PORT
      LAYER Metal5 ;
        RECT 41.130 709.640 41.430 710.640 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.943800 ;
    ANTENNADIFFAREA 0.706800 ;
    PORT
      LAYER Metal5 ;
        RECT 37.290 709.640 37.590 710.640 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.413600 ;
    PORT
      LAYER Metal5 ;
        RECT 33.450 709.640 33.750 710.640 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.413600 ;
    PORT
      LAYER Metal5 ;
        RECT 29.610 709.640 29.910 710.640 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.413600 ;
    PORT
      LAYER Metal5 ;
        RECT 87.210 709.640 87.510 710.640 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal5 ;
        RECT 83.370 709.640 83.670 710.640 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.135700 ;
    PORT
      LAYER Metal5 ;
        RECT 79.530 709.640 79.830 710.640 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.413600 ;
    PORT
      LAYER Metal5 ;
        RECT 75.690 709.640 75.990 710.640 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.124800 ;
    PORT
      LAYER Metal5 ;
        RECT 71.850 709.640 72.150 710.640 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.135700 ;
    PORT
      LAYER Metal5 ;
        RECT 68.010 709.640 68.310 710.640 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.413600 ;
    PORT
      LAYER Metal5 ;
        RECT 64.170 709.640 64.470 710.640 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.413600 ;
    PORT
      LAYER Metal5 ;
        RECT 60.330 709.640 60.630 710.640 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal5 ;
        RECT 117.930 709.640 118.230 710.640 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal5 ;
        RECT 114.090 709.640 114.390 710.640 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.023000 ;
    PORT
      LAYER Metal5 ;
        RECT 110.250 709.640 110.550 710.640 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal5 ;
        RECT 106.410 709.640 106.710 710.640 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.023000 ;
    PORT
      LAYER Metal5 ;
        RECT 102.570 709.640 102.870 710.640 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.023000 ;
    PORT
      LAYER Metal5 ;
        RECT 98.730 709.640 99.030 710.640 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.845800 ;
    PORT
      LAYER Metal5 ;
        RECT 94.890 709.640 95.190 710.640 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.988000 ;
    PORT
      LAYER Metal5 ;
        RECT 91.050 709.640 91.350 710.640 ;
    END
  END uo_out[7]
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 1068.960 707.010 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 1068.960 707.080 ;
      LAYER Metal2 ;
        RECT 2.605 3.680 1070.065 708.640 ;
      LAYER Metal3 ;
        RECT 3.260 3.635 1070.020 710.365 ;
      LAYER Metal4 ;
        RECT 3.695 3.680 1068.625 710.320 ;
      LAYER Metal5 ;
        RECT 24.380 709.430 29.400 709.640 ;
        RECT 30.120 709.430 33.240 709.640 ;
        RECT 33.960 709.430 37.080 709.640 ;
        RECT 37.800 709.430 40.920 709.640 ;
        RECT 41.640 709.430 44.760 709.640 ;
        RECT 45.480 709.430 48.600 709.640 ;
        RECT 49.320 709.430 52.440 709.640 ;
        RECT 53.160 709.430 56.280 709.640 ;
        RECT 57.000 709.430 60.120 709.640 ;
        RECT 60.840 709.430 63.960 709.640 ;
        RECT 64.680 709.430 67.800 709.640 ;
        RECT 68.520 709.430 71.640 709.640 ;
        RECT 72.360 709.430 75.480 709.640 ;
        RECT 76.200 709.430 79.320 709.640 ;
        RECT 80.040 709.430 83.160 709.640 ;
        RECT 83.880 709.430 87.000 709.640 ;
        RECT 87.720 709.430 90.840 709.640 ;
        RECT 91.560 709.430 94.680 709.640 ;
        RECT 95.400 709.430 98.520 709.640 ;
        RECT 99.240 709.430 102.360 709.640 ;
        RECT 103.080 709.430 106.200 709.640 ;
        RECT 106.920 709.430 110.040 709.640 ;
        RECT 110.760 709.430 113.880 709.640 ;
        RECT 114.600 709.430 117.720 709.640 ;
        RECT 118.440 709.430 121.560 709.640 ;
        RECT 122.280 709.430 125.400 709.640 ;
        RECT 126.120 709.430 129.240 709.640 ;
        RECT 129.960 709.430 133.080 709.640 ;
        RECT 133.800 709.430 136.920 709.640 ;
        RECT 137.640 709.430 140.760 709.640 ;
        RECT 141.480 709.430 144.600 709.640 ;
        RECT 145.320 709.430 148.440 709.640 ;
        RECT 149.160 709.430 152.280 709.640 ;
        RECT 153.000 709.430 156.120 709.640 ;
        RECT 156.840 709.430 159.960 709.640 ;
        RECT 160.680 709.430 163.800 709.640 ;
        RECT 164.520 709.430 167.640 709.640 ;
        RECT 168.360 709.430 171.480 709.640 ;
        RECT 172.200 709.430 175.320 709.640 ;
        RECT 176.040 709.430 179.160 709.640 ;
        RECT 179.880 709.430 183.000 709.640 ;
        RECT 183.720 709.430 186.840 709.640 ;
        RECT 187.560 709.430 190.680 709.640 ;
        RECT 191.400 709.430 1064.260 709.640 ;
        RECT 24.380 707.290 1064.260 709.430 ;
        RECT 24.380 12.875 54.040 707.290 ;
        RECT 56.660 12.875 60.240 707.290 ;
        RECT 62.860 12.875 92.910 707.290 ;
        RECT 95.530 12.875 99.110 707.290 ;
        RECT 101.730 12.875 131.780 707.290 ;
        RECT 134.400 12.875 137.980 707.290 ;
        RECT 140.600 12.875 170.650 707.290 ;
        RECT 173.270 12.875 176.850 707.290 ;
        RECT 179.470 12.875 209.520 707.290 ;
        RECT 212.140 12.875 215.720 707.290 ;
        RECT 218.340 12.875 248.390 707.290 ;
        RECT 251.010 12.875 254.590 707.290 ;
        RECT 257.210 12.875 287.260 707.290 ;
        RECT 289.880 12.875 293.460 707.290 ;
        RECT 296.080 12.875 326.130 707.290 ;
        RECT 328.750 12.875 332.330 707.290 ;
        RECT 334.950 12.875 365.000 707.290 ;
        RECT 367.620 12.875 371.200 707.290 ;
        RECT 373.820 12.875 403.870 707.290 ;
        RECT 406.490 12.875 410.070 707.290 ;
        RECT 412.690 12.875 442.740 707.290 ;
        RECT 445.360 12.875 448.940 707.290 ;
        RECT 451.560 12.875 481.610 707.290 ;
        RECT 484.230 12.875 487.810 707.290 ;
        RECT 490.430 12.875 520.480 707.290 ;
        RECT 523.100 12.875 526.680 707.290 ;
        RECT 529.300 12.875 559.350 707.290 ;
        RECT 561.970 12.875 565.550 707.290 ;
        RECT 568.170 12.875 598.220 707.290 ;
        RECT 600.840 12.875 604.420 707.290 ;
        RECT 607.040 12.875 637.090 707.290 ;
        RECT 639.710 12.875 643.290 707.290 ;
        RECT 645.910 12.875 675.960 707.290 ;
        RECT 678.580 12.875 682.160 707.290 ;
        RECT 684.780 12.875 714.830 707.290 ;
        RECT 717.450 12.875 721.030 707.290 ;
        RECT 723.650 12.875 753.700 707.290 ;
        RECT 756.320 12.875 759.900 707.290 ;
        RECT 762.520 12.875 792.570 707.290 ;
        RECT 795.190 12.875 798.770 707.290 ;
        RECT 801.390 12.875 831.440 707.290 ;
        RECT 834.060 12.875 837.640 707.290 ;
        RECT 840.260 12.875 870.310 707.290 ;
        RECT 872.930 12.875 876.510 707.290 ;
        RECT 879.130 12.875 909.180 707.290 ;
        RECT 911.800 12.875 915.380 707.290 ;
        RECT 918.000 12.875 948.050 707.290 ;
        RECT 950.670 12.875 954.250 707.290 ;
        RECT 956.870 12.875 986.920 707.290 ;
        RECT 989.540 12.875 993.120 707.290 ;
        RECT 995.740 12.875 1025.790 707.290 ;
        RECT 1028.410 12.875 1031.990 707.290 ;
        RECT 1034.610 12.875 1064.260 707.290 ;
  END
END tt_um_tt_tinyQV
END LIBRARY

