module tt_um_pqn (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire \pqn_inst.a[0] ;
 wire \pqn_inst.a[10] ;
 wire \pqn_inst.a[11] ;
 wire \pqn_inst.a[12] ;
 wire \pqn_inst.a[13] ;
 wire \pqn_inst.a[14] ;
 wire \pqn_inst.a[15] ;
 wire \pqn_inst.a[1] ;
 wire \pqn_inst.a[2] ;
 wire \pqn_inst.a[3] ;
 wire \pqn_inst.a[4] ;
 wire \pqn_inst.a[5] ;
 wire \pqn_inst.a[6] ;
 wire \pqn_inst.a[7] ;
 wire \pqn_inst.a[8] ;
 wire \pqn_inst.a[9] ;
 wire \pqn_inst.b[0] ;
 wire \pqn_inst.b[10] ;
 wire \pqn_inst.b[11] ;
 wire \pqn_inst.b[12] ;
 wire \pqn_inst.b[13] ;
 wire \pqn_inst.b[14] ;
 wire \pqn_inst.b[15] ;
 wire \pqn_inst.b[1] ;
 wire \pqn_inst.b[2] ;
 wire \pqn_inst.b[3] ;
 wire \pqn_inst.b[4] ;
 wire \pqn_inst.b[5] ;
 wire \pqn_inst.b[6] ;
 wire \pqn_inst.b[7] ;
 wire \pqn_inst.b[8] ;
 wire \pqn_inst.b[9] ;
 wire \pqn_inst.done ;
 wire \pqn_inst.multi.result[0] ;
 wire \pqn_inst.multi.result[10] ;
 wire \pqn_inst.multi.result[11] ;
 wire \pqn_inst.multi.result[12] ;
 wire \pqn_inst.multi.result[13] ;
 wire \pqn_inst.multi.result[14] ;
 wire \pqn_inst.multi.result[15] ;
 wire \pqn_inst.multi.result[1] ;
 wire \pqn_inst.multi.result[2] ;
 wire \pqn_inst.multi.result[3] ;
 wire \pqn_inst.multi.result[4] ;
 wire \pqn_inst.multi.result[5] ;
 wire \pqn_inst.multi.result[6] ;
 wire \pqn_inst.multi.result[7] ;
 wire \pqn_inst.multi.result[8] ;
 wire \pqn_inst.multi.result[9] ;
 wire \pqn_inst.multi.stage[0] ;
 wire \pqn_inst.multi.stage[1] ;
 wire \pqn_inst.multi.stage[2] ;
 wire \pqn_inst.multi.stage[3] ;
 wire \pqn_inst.multi.start ;
 wire \pqn_inst.multi.temp[0] ;
 wire \pqn_inst.multi.temp[1] ;
 wire \pqn_inst.multi.temp[2] ;
 wire \pqn_inst.multi.temp[3] ;
 wire \pqn_inst.multi.temp[4] ;
 wire \pqn_inst.multi.temp[5] ;
 wire \pqn_inst.multi.temp[6] ;
 wire \pqn_inst.multi.temp[7] ;
 wire \pqn_inst.multi.temp[8] ;
 wire \pqn_inst.multi.temp[9] ;
 wire \pqn_inst.n[0] ;
 wire \pqn_inst.n[10] ;
 wire \pqn_inst.n[11] ;
 wire \pqn_inst.n[12] ;
 wire \pqn_inst.n[13] ;
 wire \pqn_inst.n[14] ;
 wire \pqn_inst.n[15] ;
 wire \pqn_inst.n[1] ;
 wire \pqn_inst.n[2] ;
 wire \pqn_inst.n[3] ;
 wire \pqn_inst.n[4] ;
 wire \pqn_inst.n[5] ;
 wire \pqn_inst.n[6] ;
 wire \pqn_inst.n[7] ;
 wire \pqn_inst.n[8] ;
 wire \pqn_inst.n[9] ;
 wire \pqn_inst.stage[0] ;
 wire \pqn_inst.stage[1] ;
 wire \pqn_inst.stage[2] ;
 wire \pqn_inst.stage[3] ;
 wire \pqn_inst.v[0] ;
 wire \pqn_inst.v[10] ;
 wire \pqn_inst.v[11] ;
 wire \pqn_inst.v[12] ;
 wire \pqn_inst.v[13] ;
 wire \pqn_inst.v[14] ;
 wire \pqn_inst.v[15] ;
 wire \pqn_inst.v[1] ;
 wire \pqn_inst.v[2] ;
 wire \pqn_inst.v[3] ;
 wire \pqn_inst.v[4] ;
 wire \pqn_inst.v[5] ;
 wire \pqn_inst.v[6] ;
 wire \pqn_inst.v[7] ;
 wire \pqn_inst.v[8] ;
 wire \pqn_inst.v[9] ;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire clknet_0_clk;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;

 sg13g2_inv_1 _1543_ (.Y(_0715_),
    .A(\pqn_inst.stage[3] ));
 sg13g2_inv_1 _1544_ (.Y(_0716_),
    .A(net483));
 sg13g2_inv_1 _1545_ (.Y(_0717_),
    .A(\pqn_inst.n[10] ));
 sg13g2_inv_1 _1546_ (.Y(_0718_),
    .A(net268));
 sg13g2_inv_1 _1547_ (.Y(_0719_),
    .A(net289));
 sg13g2_inv_1 _1548_ (.Y(_0720_),
    .A(net239));
 sg13g2_inv_1 _1549_ (.Y(_0721_),
    .A(net218));
 sg13g2_inv_1 _1550_ (.Y(_0722_),
    .A(net231));
 sg13g2_inv_1 _1551_ (.Y(_0723_),
    .A(net201));
 sg13g2_inv_1 _1552_ (.Y(_0724_),
    .A(net211));
 sg13g2_inv_1 _1553_ (.Y(_0725_),
    .A(net205));
 sg13g2_inv_1 _1554_ (.Y(_0726_),
    .A(net260));
 sg13g2_inv_1 _1555_ (.Y(_0727_),
    .A(net236));
 sg13g2_inv_1 _1556_ (.Y(_0728_),
    .A(net238));
 sg13g2_inv_1 _1557_ (.Y(_0729_),
    .A(net273));
 sg13g2_inv_1 _1558_ (.Y(_0730_),
    .A(net229));
 sg13g2_inv_1 _1559_ (.Y(_0731_),
    .A(net267));
 sg13g2_inv_1 _1560_ (.Y(_0732_),
    .A(net291));
 sg13g2_inv_1 _1561_ (.Y(_0733_),
    .A(net290));
 sg13g2_inv_2 _1562_ (.Y(_0734_),
    .A(net251));
 sg13g2_inv_1 _1563_ (.Y(_0735_),
    .A(net270));
 sg13g2_inv_1 _1564_ (.Y(_0736_),
    .A(net275));
 sg13g2_inv_1 _1565_ (.Y(_0737_),
    .A(net271));
 sg13g2_inv_1 _1566_ (.Y(_0738_),
    .A(net200));
 sg13g2_inv_1 _1567_ (.Y(_0739_),
    .A(\pqn_inst.a[12] ));
 sg13g2_inv_1 _1568_ (.Y(_0740_),
    .A(\pqn_inst.a[11] ));
 sg13g2_inv_1 _1569_ (.Y(_0741_),
    .A(\pqn_inst.a[10] ));
 sg13g2_inv_1 _1570_ (.Y(_0742_),
    .A(\pqn_inst.a[9] ));
 sg13g2_inv_1 _1571_ (.Y(_0743_),
    .A(\pqn_inst.a[8] ));
 sg13g2_inv_1 _1572_ (.Y(_0744_),
    .A(\pqn_inst.a[7] ));
 sg13g2_inv_1 _1573_ (.Y(_0745_),
    .A(\pqn_inst.a[6] ));
 sg13g2_inv_1 _1574_ (.Y(_0746_),
    .A(\pqn_inst.a[5] ));
 sg13g2_inv_1 _1575_ (.Y(_0747_),
    .A(net170));
 sg13g2_inv_1 _1576_ (.Y(_0748_),
    .A(\pqn_inst.a[3] ));
 sg13g2_inv_1 _1577_ (.Y(_0749_),
    .A(\pqn_inst.a[2] ));
 sg13g2_inv_1 _1578_ (.Y(_0750_),
    .A(\pqn_inst.a[1] ));
 sg13g2_inv_1 _1579_ (.Y(_0751_),
    .A(net185));
 sg13g2_inv_1 _1580_ (.Y(_0752_),
    .A(\pqn_inst.b[15] ));
 sg13g2_inv_1 _1581_ (.Y(_0753_),
    .A(\pqn_inst.b[11] ));
 sg13g2_inv_1 _1582_ (.Y(_0754_),
    .A(\pqn_inst.b[10] ));
 sg13g2_inv_1 _1583_ (.Y(_0755_),
    .A(\pqn_inst.b[8] ));
 sg13g2_inv_1 _1584_ (.Y(_0756_),
    .A(\pqn_inst.b[3] ));
 sg13g2_inv_1 _1585_ (.Y(_0757_),
    .A(\pqn_inst.b[2] ));
 sg13g2_inv_1 _1586_ (.Y(_0758_),
    .A(\pqn_inst.b[0] ));
 sg13g2_inv_1 _1587_ (.Y(_0759_),
    .A(net495));
 sg13g2_inv_1 _1588_ (.Y(_0760_),
    .A(\pqn_inst.multi.stage[2] ));
 sg13g2_inv_1 _1589_ (.Y(_0761_),
    .A(net499));
 sg13g2_inv_1 _1590_ (.Y(_0762_),
    .A(net501));
 sg13g2_inv_1 _1591_ (.Y(_0763_),
    .A(net227));
 sg13g2_inv_4 _1592_ (.A(net486),
    .Y(_0764_));
 sg13g2_inv_2 _1593_ (.Y(_0765_),
    .A(\pqn_inst.multi.result[13] ));
 sg13g2_inv_4 _1594_ (.A(net279),
    .Y(_0766_));
 sg13g2_inv_1 _1595_ (.Y(_0767_),
    .A(\pqn_inst.multi.result[9] ));
 sg13g2_inv_2 _1596_ (.Y(_0768_),
    .A(\pqn_inst.multi.result[8] ));
 sg13g2_inv_1 _1597_ (.Y(_0769_),
    .A(\pqn_inst.multi.result[7] ));
 sg13g2_inv_2 _1598_ (.Y(_0770_),
    .A(\pqn_inst.multi.result[6] ));
 sg13g2_inv_4 _1599_ (.A(\pqn_inst.multi.result[5] ),
    .Y(_0771_));
 sg13g2_inv_2 _1600_ (.Y(_0772_),
    .A(net286));
 sg13g2_inv_2 _1601_ (.Y(_0773_),
    .A(net284));
 sg13g2_inv_1 _1602_ (.Y(_0774_),
    .A(net171));
 sg13g2_inv_1 _1603_ (.Y(_0775_),
    .A(net225));
 sg13g2_inv_1 _1604_ (.Y(_0776_),
    .A(net222));
 sg13g2_inv_1 _1605_ (.Y(_0777_),
    .A(\pqn_inst.multi.temp[2] ));
 sg13g2_inv_2 _1606_ (.Y(_0778_),
    .A(net521));
 sg13g2_inv_1 _1607_ (.Y(_0779_),
    .A(_0000_));
 sg13g2_inv_1 _1608_ (.Y(_0780_),
    .A(_0004_));
 sg13g2_inv_1 _1609_ (.Y(_0781_),
    .A(_0005_));
 sg13g2_inv_1 _1610_ (.Y(_0782_),
    .A(_0030_));
 sg13g2_inv_1 _1611_ (.Y(_0783_),
    .A(_0033_));
 sg13g2_inv_1 _1612_ (.Y(_0784_),
    .A(_0035_));
 sg13g2_inv_1 _1613_ (.Y(_0785_),
    .A(net494));
 sg13g2_inv_1 _1614_ (.Y(_0786_),
    .A(net529));
 sg13g2_and2_2 _1615_ (.A(net499),
    .B(net501),
    .X(_0787_));
 sg13g2_nor4_2 _1616_ (.A(net480),
    .B(net473),
    .C(net469),
    .Y(_0788_),
    .D(net466));
 sg13g2_nand3_1 _1617_ (.B(net497),
    .C(_0787_),
    .A(net496),
    .Y(_0789_));
 sg13g2_nand2b_1 _1618_ (.Y(_0790_),
    .B(\pqn_inst.b[12] ),
    .A_N(net501));
 sg13g2_a21oi_1 _1619_ (.A1(\pqn_inst.b[13] ),
    .A2(net501),
    .Y(_0791_),
    .B1(net499));
 sg13g2_nor2b_1 _1620_ (.A(net501),
    .B_N(net499),
    .Y(_0792_));
 sg13g2_nand2b_1 _1621_ (.Y(_0793_),
    .B(_0792_),
    .A_N(\pqn_inst.b[14] ));
 sg13g2_a221oi_1 _1622_ (.B2(_0791_),
    .C1(net473),
    .B1(_0790_),
    .A1(_0752_),
    .Y(_0794_),
    .A2(_0787_));
 sg13g2_a21oi_1 _1623_ (.A1(\pqn_inst.b[9] ),
    .A2(\pqn_inst.multi.stage[0] ),
    .Y(_0795_),
    .B1(net500));
 sg13g2_o21ai_1 _1624_ (.B1(_0795_),
    .Y(_0796_),
    .A1(_0755_),
    .A2(net502));
 sg13g2_a221oi_1 _1625_ (.B2(_0754_),
    .C1(net497),
    .B1(_0792_),
    .A1(_0753_),
    .Y(_0797_),
    .A2(_0787_));
 sg13g2_a221oi_1 _1626_ (.B2(_0797_),
    .C1(net480),
    .B1(_0796_),
    .A1(_0793_),
    .Y(_0798_),
    .A2(_0794_));
 sg13g2_mux4_1 _1627_ (.S0(net502),
    .A0(\pqn_inst.b[4] ),
    .A1(\pqn_inst.b[5] ),
    .A2(\pqn_inst.b[6] ),
    .A3(\pqn_inst.b[7] ),
    .S1(net500),
    .X(_0799_));
 sg13g2_a21oi_1 _1628_ (.A1(\pqn_inst.b[1] ),
    .A2(net502),
    .Y(_0800_),
    .B1(net500));
 sg13g2_o21ai_1 _1629_ (.B1(_0800_),
    .Y(_0801_),
    .A1(_0758_),
    .A2(net502));
 sg13g2_a221oi_1 _1630_ (.B2(_0757_),
    .C1(net497),
    .B1(_0792_),
    .A1(_0756_),
    .Y(_0802_),
    .A2(_0787_));
 sg13g2_a221oi_1 _1631_ (.B2(_0802_),
    .C1(net495),
    .B1(_0801_),
    .A1(net498),
    .Y(_0803_),
    .A2(_0799_));
 sg13g2_nor2_1 _1632_ (.A(net438),
    .B(net434),
    .Y(_0804_));
 sg13g2_or3_1 _1633_ (.A(_0751_),
    .B(net440),
    .C(net436),
    .X(_0805_));
 sg13g2_nor3_2 _1634_ (.A(net454),
    .B(net438),
    .C(net434),
    .Y(_0806_));
 sg13g2_nor4_2 _1635_ (.A(_0033_),
    .B(net459),
    .C(net440),
    .Y(_0807_),
    .D(net436));
 sg13g2_a21oi_2 _1636_ (.B1(_0807_),
    .Y(_0808_),
    .A2(_0805_),
    .A1(net459));
 sg13g2_a21o_1 _1637_ (.A2(_0805_),
    .A1(net459),
    .B1(_0807_),
    .X(_0809_));
 sg13g2_nor2_1 _1638_ (.A(net502),
    .B(_0808_),
    .Y(_0810_));
 sg13g2_and4_1 _1639_ (.A(net475),
    .B(net470),
    .C(net468),
    .D(_0807_),
    .X(_0811_));
 sg13g2_and2_1 _1640_ (.A(net478),
    .B(_0811_),
    .X(_0812_));
 sg13g2_a21oi_1 _1641_ (.A1(_0764_),
    .A2(_0812_),
    .Y(_0813_),
    .B1(net137));
 sg13g2_nand2_1 _1642_ (.Y(_0814_),
    .A(net137),
    .B(_0812_));
 sg13g2_nor2_1 _1643_ (.A(net486),
    .B(_0814_),
    .Y(_0815_));
 sg13g2_nor3_1 _1644_ (.A(net492),
    .B(_0813_),
    .C(_0815_),
    .Y(_0055_));
 sg13g2_nor2_2 _1645_ (.A(_0764_),
    .B(net492),
    .Y(_0816_));
 sg13g2_nand2b_1 _1646_ (.Y(_0817_),
    .B(net486),
    .A_N(net492));
 sg13g2_or3_1 _1647_ (.A(_0750_),
    .B(net440),
    .C(net436),
    .X(_0818_));
 sg13g2_nor4_1 _1648_ (.A(_0030_),
    .B(net459),
    .C(net440),
    .D(net436),
    .Y(_0819_));
 sg13g2_a21oi_1 _1649_ (.A1(net461),
    .A2(_0818_),
    .Y(_0820_),
    .B1(_0819_));
 sg13g2_a21o_1 _1650_ (.A2(_0818_),
    .A1(net461),
    .B1(_0819_),
    .X(_0821_));
 sg13g2_a221oi_1 _1651_ (.B2(net461),
    .C1(net502),
    .B1(_0818_),
    .A1(_0782_),
    .Y(_0822_),
    .A2(_0806_));
 sg13g2_a221oi_1 _1652_ (.B2(_0783_),
    .C1(net468),
    .B1(_0806_),
    .A1(net459),
    .Y(_0823_),
    .A2(_0805_));
 sg13g2_or3_1 _1653_ (.A(net500),
    .B(_0822_),
    .C(_0823_),
    .X(_0824_));
 sg13g2_nor4_2 _1654_ (.A(net498),
    .B(net499),
    .C(_0822_),
    .Y(_0825_),
    .D(_0823_));
 sg13g2_nand2_1 _1655_ (.Y(_0826_),
    .A(net478),
    .B(_0825_));
 sg13g2_nand3_1 _1656_ (.B(\pqn_inst.multi.temp[1] ),
    .C(_0825_),
    .A(net477),
    .Y(_0827_));
 sg13g2_a21oi_1 _1657_ (.A1(net477),
    .A2(_0825_),
    .Y(_0828_),
    .B1(\pqn_inst.multi.temp[1] ));
 sg13g2_xor2_1 _1658_ (.B(_0826_),
    .A(net174),
    .X(_0829_));
 sg13g2_nor2_2 _1659_ (.A(net486),
    .B(net492),
    .Y(_0830_));
 sg13g2_or2_1 _1660_ (.X(_0831_),
    .B(net492),
    .A(net486));
 sg13g2_xor2_1 _1661_ (.B(_0829_),
    .A(_0814_),
    .X(_0832_));
 sg13g2_a22oi_1 _1662_ (.Y(_0833_),
    .B1(_0830_),
    .B2(_0832_),
    .A2(net453),
    .A1(net174));
 sg13g2_inv_1 _1663_ (.Y(_0056_),
    .A(_0833_));
 sg13g2_nand2_1 _1664_ (.Y(_0834_),
    .A(net138),
    .B(net453));
 sg13g2_o21ai_1 _1665_ (.B1(_0827_),
    .Y(_0835_),
    .A1(_0814_),
    .A2(_0828_));
 sg13g2_or3_1 _1666_ (.A(_0749_),
    .B(net440),
    .C(_0803_),
    .X(_0836_));
 sg13g2_nor4_2 _1667_ (.A(_0035_),
    .B(net460),
    .C(net440),
    .Y(_0837_),
    .D(net436));
 sg13g2_a21oi_2 _1668_ (.B1(_0837_),
    .Y(_0838_),
    .A2(_0836_),
    .A1(net460));
 sg13g2_a21o_1 _1669_ (.A2(_0836_),
    .A1(net460),
    .B1(_0837_),
    .X(_0839_));
 sg13g2_a221oi_1 _1670_ (.B2(net460),
    .C1(net502),
    .B1(_0836_),
    .A1(_0784_),
    .Y(_0840_),
    .A2(_0806_));
 sg13g2_a221oi_1 _1671_ (.B2(net461),
    .C1(net468),
    .B1(_0818_),
    .A1(_0782_),
    .Y(_0841_),
    .A2(_0806_));
 sg13g2_nor2_1 _1672_ (.A(_0840_),
    .B(_0841_),
    .Y(_0842_));
 sg13g2_o21ai_1 _1673_ (.B1(net499),
    .Y(_0843_),
    .A1(net501),
    .A2(_0808_));
 sg13g2_o21ai_1 _1674_ (.B1(net470),
    .Y(_0844_),
    .A1(_0840_),
    .A2(_0841_));
 sg13g2_nand3_1 _1675_ (.B(_0843_),
    .C(_0844_),
    .A(net475),
    .Y(_0845_));
 sg13g2_nand4_1 _1676_ (.B(_0031_),
    .C(_0843_),
    .A(net475),
    .Y(_0846_),
    .D(_0844_));
 sg13g2_xor2_1 _1677_ (.B(_0846_),
    .A(_0034_),
    .X(_0847_));
 sg13g2_and2_1 _1678_ (.A(_0835_),
    .B(_0847_),
    .X(_0848_));
 sg13g2_o21ai_1 _1679_ (.B1(_0830_),
    .Y(_0849_),
    .A1(_0835_),
    .A2(_0847_));
 sg13g2_o21ai_1 _1680_ (.B1(_0834_),
    .Y(_0057_),
    .A1(_0848_),
    .A2(_0849_));
 sg13g2_nor2_1 _1681_ (.A(_0777_),
    .B(_0846_),
    .Y(_0850_));
 sg13g2_a21oi_1 _1682_ (.A1(_0835_),
    .A2(_0847_),
    .Y(_0851_),
    .B1(_0850_));
 sg13g2_a21o_1 _1683_ (.A2(_0847_),
    .A1(_0835_),
    .B1(_0850_),
    .X(_0852_));
 sg13g2_or3_1 _1684_ (.A(_0748_),
    .B(_0798_),
    .C(net436),
    .X(_0853_));
 sg13g2_nor4_2 _1685_ (.A(_0036_),
    .B(net459),
    .C(net440),
    .Y(_0854_),
    .D(net436));
 sg13g2_a21oi_2 _1686_ (.B1(_0854_),
    .Y(_0855_),
    .A2(_0853_),
    .A1(net459));
 sg13g2_a21o_1 _1687_ (.A2(_0853_),
    .A1(net459),
    .B1(_0854_),
    .X(_0856_));
 sg13g2_mux4_1 _1688_ (.S0(net468),
    .A0(_0808_),
    .A1(_0820_),
    .A2(_0838_),
    .A3(_0855_),
    .S1(net471),
    .X(_0857_));
 sg13g2_mux4_1 _1689_ (.S0(net468),
    .A0(_0809_),
    .A1(_0821_),
    .A2(_0839_),
    .A3(_0856_),
    .S1(net471),
    .X(_0858_));
 sg13g2_nor2_2 _1690_ (.A(net498),
    .B(_0857_),
    .Y(_0859_));
 sg13g2_nand2_2 _1691_ (.Y(_0860_),
    .A(_0031_),
    .B(_0859_));
 sg13g2_nor2_1 _1692_ (.A(_0776_),
    .B(_0860_),
    .Y(_0861_));
 sg13g2_xnor2_1 _1693_ (.Y(_0862_),
    .A(\pqn_inst.multi.temp[3] ),
    .B(_0860_));
 sg13g2_xnor2_1 _1694_ (.Y(_0863_),
    .A(_0776_),
    .B(_0860_));
 sg13g2_a21oi_1 _1695_ (.A1(_0851_),
    .A2(_0863_),
    .Y(_0864_),
    .B1(net462));
 sg13g2_o21ai_1 _1696_ (.B1(_0864_),
    .Y(_0865_),
    .A1(_0851_),
    .A2(_0863_));
 sg13g2_o21ai_1 _1697_ (.B1(_0865_),
    .Y(_0058_),
    .A1(_0776_),
    .A2(net463));
 sg13g2_nand2_1 _1698_ (.Y(_0866_),
    .A(net160),
    .B(net453));
 sg13g2_a21oi_1 _1699_ (.A1(_0852_),
    .A2(_0862_),
    .Y(_0867_),
    .B1(_0861_));
 sg13g2_a21o_1 _1700_ (.A2(_0862_),
    .A1(_0852_),
    .B1(_0861_),
    .X(_0868_));
 sg13g2_nand4_1 _1701_ (.B(net470),
    .C(net468),
    .A(net498),
    .Y(_0869_),
    .D(_0809_));
 sg13g2_or3_1 _1702_ (.A(_0747_),
    .B(net441),
    .C(net437),
    .X(_0870_));
 sg13g2_nor4_2 _1703_ (.A(_0038_),
    .B(net458),
    .C(net440),
    .Y(_0871_),
    .D(net436));
 sg13g2_a21oi_2 _1704_ (.B1(_0871_),
    .Y(_0872_),
    .A2(_0870_),
    .A1(net457));
 sg13g2_a21o_1 _1705_ (.A2(_0870_),
    .A1(net457),
    .B1(_0871_),
    .X(_0873_));
 sg13g2_mux2_1 _1706_ (.A0(_0856_),
    .A1(_0873_),
    .S(net467),
    .X(_0874_));
 sg13g2_mux4_1 _1707_ (.S0(net467),
    .A0(_0820_),
    .A1(_0838_),
    .A2(_0855_),
    .A3(_0872_),
    .S1(net471),
    .X(_0875_));
 sg13g2_o21ai_1 _1708_ (.B1(_0869_),
    .Y(_0876_),
    .A1(net498),
    .A2(_0875_));
 sg13g2_nand2_1 _1709_ (.Y(_0877_),
    .A(_0031_),
    .B(_0876_));
 sg13g2_xor2_1 _1710_ (.B(_0877_),
    .A(_0037_),
    .X(_0878_));
 sg13g2_and2_1 _1711_ (.A(_0868_),
    .B(_0878_),
    .X(_0879_));
 sg13g2_o21ai_1 _1712_ (.B1(_0830_),
    .Y(_0880_),
    .A1(_0868_),
    .A2(_0878_));
 sg13g2_o21ai_1 _1713_ (.B1(_0866_),
    .Y(_0059_),
    .A1(_0879_),
    .A2(_0880_));
 sg13g2_nand3_1 _1714_ (.B(net494),
    .C(_0876_),
    .A(\pqn_inst.multi.temp[4] ),
    .Y(_0881_));
 sg13g2_nor2b_1 _1715_ (.A(_0879_),
    .B_N(_0881_),
    .Y(_0882_));
 sg13g2_or4_1 _1716_ (.A(net475),
    .B(net499),
    .C(_0822_),
    .D(_0823_),
    .X(_0883_));
 sg13g2_or3_1 _1717_ (.A(_0746_),
    .B(net441),
    .C(net437),
    .X(_0884_));
 sg13g2_nor4_2 _1718_ (.A(_0039_),
    .B(net458),
    .C(net441),
    .Y(_0885_),
    .D(net437));
 sg13g2_a21oi_2 _1719_ (.B1(_0885_),
    .Y(_0886_),
    .A2(_0884_),
    .A1(net457));
 sg13g2_a21o_1 _1720_ (.A2(_0884_),
    .A1(net458),
    .B1(_0885_),
    .X(_0887_));
 sg13g2_mux4_1 _1721_ (.S0(net467),
    .A0(_0838_),
    .A1(_0855_),
    .A2(_0872_),
    .A3(_0886_),
    .S1(net471),
    .X(_0888_));
 sg13g2_o21ai_1 _1722_ (.B1(_0883_),
    .Y(_0889_),
    .A1(net498),
    .A2(_0888_));
 sg13g2_nand2_1 _1723_ (.Y(_0890_),
    .A(net494),
    .B(_0889_));
 sg13g2_nand3_1 _1724_ (.B(net494),
    .C(_0889_),
    .A(\pqn_inst.multi.temp[5] ),
    .Y(_0891_));
 sg13g2_a21oi_1 _1725_ (.A1(net494),
    .A2(_0889_),
    .Y(_0892_),
    .B1(\pqn_inst.multi.temp[5] ));
 sg13g2_xnor2_1 _1726_ (.Y(_0893_),
    .A(\pqn_inst.multi.temp[5] ),
    .B(_0890_));
 sg13g2_o21ai_1 _1727_ (.B1(_0764_),
    .Y(_0894_),
    .A1(_0882_),
    .A2(_0893_));
 sg13g2_a21oi_1 _1728_ (.A1(_0882_),
    .A2(_0893_),
    .Y(_0895_),
    .B1(_0894_));
 sg13g2_nand2b_1 _1729_ (.Y(_0896_),
    .B(net203),
    .A_N(net492));
 sg13g2_a21oi_1 _1730_ (.A1(net462),
    .A2(_0896_),
    .Y(_0060_),
    .B1(_0895_));
 sg13g2_a21oi_1 _1731_ (.A1(_0881_),
    .A2(_0891_),
    .Y(_0897_),
    .B1(_0892_));
 sg13g2_and2_1 _1732_ (.A(_0878_),
    .B(_0893_),
    .X(_0898_));
 sg13g2_a21oi_1 _1733_ (.A1(_0868_),
    .A2(_0898_),
    .Y(_0899_),
    .B1(_0897_));
 sg13g2_or3_1 _1734_ (.A(_0745_),
    .B(net441),
    .C(net437),
    .X(_0900_));
 sg13g2_nor4_2 _1735_ (.A(_0040_),
    .B(net457),
    .C(net441),
    .Y(_0901_),
    .D(net437));
 sg13g2_a21oi_2 _1736_ (.B1(_0901_),
    .Y(_0902_),
    .A2(_0900_),
    .A1(net458));
 sg13g2_a21o_1 _1737_ (.A2(_0900_),
    .A1(net457),
    .B1(_0901_),
    .X(_0903_));
 sg13g2_mux2_1 _1738_ (.A0(_0887_),
    .A1(_0903_),
    .S(net467),
    .X(_0904_));
 sg13g2_mux4_1 _1739_ (.S0(net467),
    .A0(_0855_),
    .A1(_0872_),
    .A2(_0886_),
    .A3(_0902_),
    .S1(net470),
    .X(_0905_));
 sg13g2_mux4_1 _1740_ (.S0(net470),
    .A0(_0810_),
    .A1(_0842_),
    .A2(_0874_),
    .A3(_0904_),
    .S1(net476),
    .X(_0906_));
 sg13g2_and3_1 _1741_ (.X(_0907_),
    .A(\pqn_inst.multi.temp[6] ),
    .B(net494),
    .C(_0906_));
 sg13g2_a21oi_1 _1742_ (.A1(net494),
    .A2(_0906_),
    .Y(_0908_),
    .B1(\pqn_inst.multi.temp[6] ));
 sg13g2_or2_1 _1743_ (.X(_0909_),
    .B(_0908_),
    .A(_0907_));
 sg13g2_or2_1 _1744_ (.X(_0910_),
    .B(_0909_),
    .A(_0899_));
 sg13g2_a21oi_1 _1745_ (.A1(_0899_),
    .A2(_0909_),
    .Y(_0911_),
    .B1(_0831_));
 sg13g2_a22oi_1 _1746_ (.Y(_0912_),
    .B1(_0910_),
    .B2(_0911_),
    .A2(net453),
    .A1(net165));
 sg13g2_inv_1 _1747_ (.Y(_0061_),
    .A(_0912_));
 sg13g2_nor2b_1 _1748_ (.A(_0907_),
    .B_N(_0910_),
    .Y(_0913_));
 sg13g2_or3_1 _1749_ (.A(_0744_),
    .B(net441),
    .C(net437),
    .X(_0914_));
 sg13g2_nor4_2 _1750_ (.A(_0041_),
    .B(net457),
    .C(net441),
    .Y(_0915_),
    .D(net437));
 sg13g2_a21oi_2 _1751_ (.B1(_0915_),
    .Y(_0916_),
    .A2(_0914_),
    .A1(net457));
 sg13g2_a21o_1 _1752_ (.A2(_0914_),
    .A1(net457),
    .B1(_0915_),
    .X(_0917_));
 sg13g2_mux4_1 _1753_ (.S0(net467),
    .A0(_0872_),
    .A1(_0886_),
    .A2(_0902_),
    .A3(_0916_),
    .S1(net470),
    .X(_0918_));
 sg13g2_mux4_1 _1754_ (.S0(net467),
    .A0(_0873_),
    .A1(_0887_),
    .A2(_0903_),
    .A3(_0917_),
    .S1(net470),
    .X(_0919_));
 sg13g2_mux2_1 _1755_ (.A0(_0857_),
    .A1(_0918_),
    .S(net475),
    .X(_0920_));
 sg13g2_mux2_1 _1756_ (.A0(_0858_),
    .A1(_0919_),
    .S(net476),
    .X(_0921_));
 sg13g2_a21oi_1 _1757_ (.A1(net494),
    .A2(_0921_),
    .Y(_0922_),
    .B1(\pqn_inst.multi.temp[7] ));
 sg13g2_o21ai_1 _1758_ (.B1(_0775_),
    .Y(_0923_),
    .A1(_0785_),
    .A2(_0920_));
 sg13g2_nor3_2 _1759_ (.A(_0775_),
    .B(_0785_),
    .C(_0920_),
    .Y(_0924_));
 sg13g2_nor2_1 _1760_ (.A(_0922_),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_or2_1 _1761_ (.X(_0926_),
    .B(_0925_),
    .A(_0913_));
 sg13g2_a21oi_1 _1762_ (.A1(_0913_),
    .A2(_0925_),
    .Y(_0927_),
    .B1(net488));
 sg13g2_a221oi_1 _1763_ (.B2(_0927_),
    .C1(net493),
    .B1(_0926_),
    .A1(net488),
    .Y(_0062_),
    .A2(_0775_));
 sg13g2_nor4_2 _1764_ (.A(_0907_),
    .B(_0908_),
    .C(_0922_),
    .Y(_0928_),
    .D(_0924_));
 sg13g2_nand3_1 _1765_ (.B(_0893_),
    .C(_0928_),
    .A(_0878_),
    .Y(_0929_));
 sg13g2_a221oi_1 _1766_ (.B2(_0897_),
    .C1(_0924_),
    .B1(_0928_),
    .A1(_0907_),
    .Y(_0930_),
    .A2(_0923_));
 sg13g2_o21ai_1 _1767_ (.B1(_0930_),
    .Y(_0931_),
    .A1(_0867_),
    .A2(_0929_));
 sg13g2_nor2_1 _1768_ (.A(net478),
    .B(_0811_),
    .Y(_0932_));
 sg13g2_or3_1 _1769_ (.A(_0743_),
    .B(net439),
    .C(net435),
    .X(_0933_));
 sg13g2_nor4_2 _1770_ (.A(_0042_),
    .B(net456),
    .C(net439),
    .Y(_0934_),
    .D(net435));
 sg13g2_a21oi_2 _1771_ (.B1(_0934_),
    .Y(_0935_),
    .A2(_0933_),
    .A1(net456));
 sg13g2_a21o_1 _1772_ (.A2(_0933_),
    .A1(net456),
    .B1(_0934_),
    .X(_0936_));
 sg13g2_mux4_1 _1773_ (.S0(net467),
    .A0(_0886_),
    .A1(_0902_),
    .A2(_0916_),
    .A3(_0935_),
    .S1(net470),
    .X(_0937_));
 sg13g2_mux4_1 _1774_ (.S0(net466),
    .A0(_0887_),
    .A1(_0903_),
    .A2(_0917_),
    .A3(_0936_),
    .S1(net472),
    .X(_0938_));
 sg13g2_mux2_1 _1775_ (.A0(_0875_),
    .A1(_0937_),
    .S(net475),
    .X(_0939_));
 sg13g2_a21oi_1 _1776_ (.A1(net478),
    .A2(_0939_),
    .Y(_0940_),
    .B1(_0932_));
 sg13g2_nand2_1 _1777_ (.Y(_0941_),
    .A(net171),
    .B(_0940_));
 sg13g2_xnor2_1 _1778_ (.Y(_0942_),
    .A(\pqn_inst.multi.temp[8] ),
    .B(_0940_));
 sg13g2_nand2b_1 _1779_ (.Y(_0943_),
    .B(_0942_),
    .A_N(_0931_));
 sg13g2_nand2b_1 _1780_ (.Y(_0944_),
    .B(_0931_),
    .A_N(_0942_));
 sg13g2_nand3_1 _1781_ (.B(_0943_),
    .C(_0944_),
    .A(_0830_),
    .Y(_0945_));
 sg13g2_o21ai_1 _1782_ (.B1(_0945_),
    .Y(_0063_),
    .A1(_0774_),
    .A2(net463));
 sg13g2_nor2_1 _1783_ (.A(net477),
    .B(_0825_),
    .Y(_0946_));
 sg13g2_or3_1 _1784_ (.A(_0742_),
    .B(net439),
    .C(net434),
    .X(_0947_));
 sg13g2_nor4_2 _1785_ (.A(_0043_),
    .B(net454),
    .C(net438),
    .Y(_0948_),
    .D(net434));
 sg13g2_a21oi_2 _1786_ (.B1(_0948_),
    .Y(_0949_),
    .A2(_0947_),
    .A1(net456));
 sg13g2_a21o_1 _1787_ (.A2(_0947_),
    .A1(net456),
    .B1(_0948_),
    .X(_0950_));
 sg13g2_mux4_1 _1788_ (.S0(net466),
    .A0(_0902_),
    .A1(_0916_),
    .A2(_0935_),
    .A3(_0949_),
    .S1(net472),
    .X(_0951_));
 sg13g2_mux2_1 _1789_ (.A0(_0888_),
    .A1(_0951_),
    .S(net475),
    .X(_0952_));
 sg13g2_a21oi_2 _1790_ (.B1(_0946_),
    .Y(_0953_),
    .A2(_0952_),
    .A1(net477));
 sg13g2_nand2_1 _1791_ (.Y(_0954_),
    .A(\pqn_inst.multi.temp[9] ),
    .B(_0953_));
 sg13g2_nor2_1 _1792_ (.A(\pqn_inst.multi.temp[9] ),
    .B(_0953_),
    .Y(_0955_));
 sg13g2_xor2_1 _1793_ (.B(_0953_),
    .A(net199),
    .X(_0956_));
 sg13g2_nand3_1 _1794_ (.B(_0944_),
    .C(_0956_),
    .A(_0941_),
    .Y(_0957_));
 sg13g2_a21oi_1 _1795_ (.A1(_0941_),
    .A2(_0944_),
    .Y(_0958_),
    .B1(_0956_));
 sg13g2_nor2_1 _1796_ (.A(net486),
    .B(_0958_),
    .Y(_0959_));
 sg13g2_nand2b_1 _1797_ (.Y(_0960_),
    .B(net199),
    .A_N(net493));
 sg13g2_a22oi_1 _1798_ (.Y(_0064_),
    .B1(_0960_),
    .B2(net462),
    .A2(_0959_),
    .A1(_0957_));
 sg13g2_o21ai_1 _1799_ (.B1(_0954_),
    .Y(_0961_),
    .A1(_0941_),
    .A2(_0955_));
 sg13g2_nor2b_1 _1800_ (.A(_0942_),
    .B_N(_0956_),
    .Y(_0962_));
 sg13g2_a21oi_1 _1801_ (.A1(_0931_),
    .A2(_0962_),
    .Y(_0963_),
    .B1(_0961_));
 sg13g2_or3_1 _1802_ (.A(_0741_),
    .B(net438),
    .C(net434),
    .X(_0964_));
 sg13g2_nor4_2 _1803_ (.A(_0044_),
    .B(net455),
    .C(net438),
    .Y(_0965_),
    .D(net434));
 sg13g2_a21oi_2 _1804_ (.B1(_0965_),
    .Y(_0966_),
    .A2(_0964_),
    .A1(net455));
 sg13g2_a21o_1 _1805_ (.A2(_0964_),
    .A1(net455),
    .B1(_0965_),
    .X(_0967_));
 sg13g2_mux4_1 _1806_ (.S0(net466),
    .A0(_0916_),
    .A1(_0935_),
    .A2(_0949_),
    .A3(_0966_),
    .S1(net472),
    .X(_0968_));
 sg13g2_mux2_1 _1807_ (.A0(_0905_),
    .A1(_0968_),
    .S(net474),
    .X(_0969_));
 sg13g2_mux2_1 _1808_ (.A0(_0845_),
    .A1(_0969_),
    .S(net477),
    .X(_0970_));
 sg13g2_xnor2_1 _1809_ (.Y(_0971_),
    .A(_0773_),
    .B(_0970_));
 sg13g2_nor2_1 _1810_ (.A(_0963_),
    .B(_0971_),
    .Y(_0972_));
 sg13g2_a21oi_1 _1811_ (.A1(_0963_),
    .A2(_0971_),
    .Y(_0973_),
    .B1(net462));
 sg13g2_nand2b_1 _1812_ (.Y(_0974_),
    .B(_0973_),
    .A_N(_0972_));
 sg13g2_o21ai_1 _1813_ (.B1(_0974_),
    .Y(_0065_),
    .A1(_0773_),
    .A2(_0817_));
 sg13g2_nor2_1 _1814_ (.A(_0017_),
    .B(_0970_),
    .Y(_0975_));
 sg13g2_or2_1 _1815_ (.X(_0976_),
    .B(_0975_),
    .A(_0972_));
 sg13g2_nor3_1 _1816_ (.A(_0740_),
    .B(net438),
    .C(net435),
    .Y(_0977_));
 sg13g2_nor2_1 _1817_ (.A(_0789_),
    .B(_0977_),
    .Y(_0978_));
 sg13g2_or4_1 _1818_ (.A(_0045_),
    .B(net454),
    .C(net438),
    .D(net434),
    .X(_0979_));
 sg13g2_nor2b_1 _1819_ (.A(_0978_),
    .B_N(_0979_),
    .Y(_0980_));
 sg13g2_o21ai_1 _1820_ (.B1(_0979_),
    .Y(_0981_),
    .A1(_0789_),
    .A2(_0977_));
 sg13g2_mux4_1 _1821_ (.S0(net465),
    .A0(_0936_),
    .A1(_0950_),
    .A2(_0967_),
    .A3(_0981_),
    .S1(net469),
    .X(_0982_));
 sg13g2_mux2_1 _1822_ (.A0(_0919_),
    .A1(_0982_),
    .S(net473),
    .X(_0983_));
 sg13g2_mux2_2 _1823_ (.A0(_0859_),
    .A1(_0983_),
    .S(net477),
    .X(_0984_));
 sg13g2_nand2_1 _1824_ (.Y(_0985_),
    .A(net507),
    .B(_0984_));
 sg13g2_xnor2_1 _1825_ (.Y(_0986_),
    .A(net507),
    .B(_0984_));
 sg13g2_o21ai_1 _1826_ (.B1(_0764_),
    .Y(_0987_),
    .A1(_0976_),
    .A2(_0986_));
 sg13g2_a21oi_1 _1827_ (.A1(_0976_),
    .A2(_0986_),
    .Y(_0988_),
    .B1(_0987_));
 sg13g2_nand2b_1 _1828_ (.Y(_0989_),
    .B(net507),
    .A_N(net493));
 sg13g2_a21oi_1 _1829_ (.A1(net462),
    .A2(_0989_),
    .Y(_0066_),
    .B1(_0988_));
 sg13g2_nand2_1 _1830_ (.Y(_0990_),
    .A(net255),
    .B(_0816_));
 sg13g2_nor2_1 _1831_ (.A(_0971_),
    .B(_0986_),
    .Y(_0991_));
 sg13g2_and2_1 _1832_ (.A(_0962_),
    .B(_0991_),
    .X(_0992_));
 sg13g2_nand2_1 _1833_ (.Y(_0993_),
    .A(_0931_),
    .B(_0992_));
 sg13g2_and2_1 _1834_ (.A(_0961_),
    .B(_0991_),
    .X(_0994_));
 sg13g2_o21ai_1 _1835_ (.B1(_0975_),
    .Y(_0995_),
    .A1(net507),
    .A2(_0984_));
 sg13g2_nand2_1 _1836_ (.Y(_0996_),
    .A(_0985_),
    .B(_0995_));
 sg13g2_a221oi_1 _1837_ (.B2(_0931_),
    .C1(_0996_),
    .B1(_0992_),
    .A1(_0961_),
    .Y(_0997_),
    .A2(_0991_));
 sg13g2_nor3_1 _1838_ (.A(_0739_),
    .B(net438),
    .C(net434),
    .Y(_0998_));
 sg13g2_nor2_1 _1839_ (.A(_0789_),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_or4_1 _1840_ (.A(_0046_),
    .B(net455),
    .C(net439),
    .D(net435),
    .X(_1000_));
 sg13g2_nor2b_1 _1841_ (.A(_0999_),
    .B_N(_1000_),
    .Y(_1001_));
 sg13g2_o21ai_1 _1842_ (.B1(_1000_),
    .Y(_1002_),
    .A1(_0789_),
    .A2(_0998_));
 sg13g2_mux4_1 _1843_ (.S0(net465),
    .A0(_0950_),
    .A1(_0967_),
    .A2(_0981_),
    .A3(_1002_),
    .S1(net469),
    .X(_1003_));
 sg13g2_mux2_2 _1844_ (.A0(_0938_),
    .A1(_1003_),
    .S(net474),
    .X(_1004_));
 sg13g2_mux2_1 _1845_ (.A0(_0876_),
    .A1(_1004_),
    .S(net477),
    .X(_1005_));
 sg13g2_xnor2_1 _1846_ (.Y(_1006_),
    .A(\pqn_inst.multi.result[2] ),
    .B(_1005_));
 sg13g2_nor2_1 _1847_ (.A(_0997_),
    .B(_1006_),
    .Y(_1007_));
 sg13g2_a21o_1 _1848_ (.A2(_1006_),
    .A1(_0997_),
    .B1(net462),
    .X(_1008_));
 sg13g2_o21ai_1 _1849_ (.B1(_0990_),
    .Y(_0067_),
    .A1(_1007_),
    .A2(_1008_));
 sg13g2_nor2b_1 _1850_ (.A(_0020_),
    .B_N(_1005_),
    .Y(_1009_));
 sg13g2_nor2_1 _1851_ (.A(_1007_),
    .B(_1009_),
    .Y(_1010_));
 sg13g2_a21oi_1 _1852_ (.A1(\pqn_inst.a[13] ),
    .A2(_0804_),
    .Y(_1011_),
    .B1(_0789_));
 sg13g2_nand2b_1 _1853_ (.Y(_1012_),
    .B(_0806_),
    .A_N(_0047_));
 sg13g2_nor2b_1 _1854_ (.A(_1011_),
    .B_N(_1012_),
    .Y(_1013_));
 sg13g2_nand2b_1 _1855_ (.Y(_1014_),
    .B(_1012_),
    .A_N(_1011_));
 sg13g2_mux4_1 _1856_ (.S0(net465),
    .A0(_0966_),
    .A1(_0980_),
    .A2(_1001_),
    .A3(_1013_),
    .S1(net469),
    .X(_1015_));
 sg13g2_and2_1 _1857_ (.A(net497),
    .B(_0951_),
    .X(_1016_));
 sg13g2_a21oi_1 _1858_ (.A1(net473),
    .A2(_1015_),
    .Y(_1017_),
    .B1(_1016_));
 sg13g2_mux4_1 _1859_ (.S0(net475),
    .A0(_0824_),
    .A1(_0888_),
    .A2(_0951_),
    .A3(_1015_),
    .S1(net477),
    .X(_1018_));
 sg13g2_nand2_1 _1860_ (.Y(_1019_),
    .A(_0772_),
    .B(_1018_));
 sg13g2_inv_1 _1861_ (.Y(_1020_),
    .A(_1019_));
 sg13g2_nor2_1 _1862_ (.A(_0772_),
    .B(_1018_),
    .Y(_1021_));
 sg13g2_nor2_1 _1863_ (.A(_1020_),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_or2_1 _1864_ (.X(_1023_),
    .B(_1022_),
    .A(_1010_));
 sg13g2_nor3_1 _1865_ (.A(_1007_),
    .B(_1009_),
    .C(_1021_),
    .Y(_1024_));
 sg13g2_a21oi_1 _1866_ (.A1(_1010_),
    .A2(_1022_),
    .Y(_1025_),
    .B1(net487));
 sg13g2_a221oi_1 _1867_ (.B2(_1025_),
    .C1(net493),
    .B1(_1023_),
    .A1(net487),
    .Y(_0068_),
    .A2(_0772_));
 sg13g2_nand2_1 _1868_ (.Y(_1026_),
    .A(net506),
    .B(_0816_));
 sg13g2_nand2_1 _1869_ (.Y(_1027_),
    .A(\pqn_inst.a[14] ),
    .B(_0804_));
 sg13g2_nor2b_1 _1870_ (.A(_0048_),
    .B_N(_0806_),
    .Y(_1028_));
 sg13g2_a21oi_1 _1871_ (.A1(net454),
    .A2(_1027_),
    .Y(_1029_),
    .B1(_1028_));
 sg13g2_a21o_1 _1872_ (.A2(_1027_),
    .A1(net454),
    .B1(_1028_),
    .X(_1030_));
 sg13g2_mux2_1 _1873_ (.A0(_1013_),
    .A1(_1029_),
    .S(net465),
    .X(_1031_));
 sg13g2_mux4_1 _1874_ (.S0(net465),
    .A0(_0981_),
    .A1(_1002_),
    .A2(_1014_),
    .A3(_1030_),
    .S1(net469),
    .X(_1032_));
 sg13g2_nor2_1 _1875_ (.A(net474),
    .B(_0968_),
    .Y(_1033_));
 sg13g2_a21o_1 _1876_ (.A2(_1032_),
    .A1(net473),
    .B1(_1033_),
    .X(_1034_));
 sg13g2_mux2_1 _1877_ (.A0(_0906_),
    .A1(_1034_),
    .S(net479),
    .X(_1035_));
 sg13g2_xnor2_1 _1878_ (.Y(_1036_),
    .A(net506),
    .B(_1035_));
 sg13g2_nor3_2 _1879_ (.A(_1020_),
    .B(_1024_),
    .C(_1036_),
    .Y(_1037_));
 sg13g2_o21ai_1 _1880_ (.B1(_1036_),
    .Y(_1038_),
    .A1(_1020_),
    .A2(_1024_));
 sg13g2_nand2_1 _1881_ (.Y(_1039_),
    .A(_0830_),
    .B(_1038_));
 sg13g2_o21ai_1 _1882_ (.B1(_1026_),
    .Y(_0069_),
    .A1(_1037_),
    .A2(_1039_));
 sg13g2_nor2b_1 _1883_ (.A(net272),
    .B_N(_1035_),
    .Y(_1040_));
 sg13g2_nand2b_1 _1884_ (.Y(_1041_),
    .B(_1035_),
    .A_N(_0023_));
 sg13g2_nand2_1 _1885_ (.Y(_1042_),
    .A(\pqn_inst.a[15] ),
    .B(_0804_));
 sg13g2_a22oi_1 _1886_ (.Y(_1043_),
    .B1(_1042_),
    .B2(net454),
    .A2(_0806_),
    .A1(\pqn_inst.a[15] ));
 sg13g2_nand3_1 _1887_ (.B(net465),
    .C(_0806_),
    .A(\pqn_inst.a[15] ),
    .Y(_1044_));
 sg13g2_o21ai_1 _1888_ (.B1(_1044_),
    .Y(_1045_),
    .A1(net465),
    .A2(_1030_));
 sg13g2_mux4_1 _1889_ (.S0(net465),
    .A0(_1002_),
    .A1(_1014_),
    .A2(_1030_),
    .A3(_1043_),
    .S1(net469),
    .X(_1046_));
 sg13g2_mux2_2 _1890_ (.A0(_0982_),
    .A1(_1046_),
    .S(net474),
    .X(_1047_));
 sg13g2_mux2_1 _1891_ (.A0(_0921_),
    .A1(_1047_),
    .S(net479),
    .X(_1048_));
 sg13g2_nor2_1 _1892_ (.A(\pqn_inst.multi.result[5] ),
    .B(_1048_),
    .Y(_1049_));
 sg13g2_nand2_1 _1893_ (.Y(_1050_),
    .A(\pqn_inst.multi.result[5] ),
    .B(_1048_));
 sg13g2_xnor2_1 _1894_ (.Y(_1051_),
    .A(\pqn_inst.multi.result[5] ),
    .B(_1048_));
 sg13g2_o21ai_1 _1895_ (.B1(_1051_),
    .Y(_1052_),
    .A1(_1037_),
    .A2(_1040_));
 sg13g2_nor3_1 _1896_ (.A(_1037_),
    .B(_1040_),
    .C(_1051_),
    .Y(_1053_));
 sg13g2_nor2_1 _1897_ (.A(net487),
    .B(_1053_),
    .Y(_1054_));
 sg13g2_a221oi_1 _1898_ (.B2(_1054_),
    .C1(net492),
    .B1(_1052_),
    .A1(net487),
    .Y(_0070_),
    .A2(_0771_));
 sg13g2_a21oi_1 _1899_ (.A1(_1009_),
    .A2(_1019_),
    .Y(_1055_),
    .B1(_1021_));
 sg13g2_nor3_1 _1900_ (.A(_1036_),
    .B(_1051_),
    .C(_1055_),
    .Y(_1056_));
 sg13g2_o21ai_1 _1901_ (.B1(_1050_),
    .Y(_1057_),
    .A1(_1041_),
    .A2(_1049_));
 sg13g2_nor2_1 _1902_ (.A(_1056_),
    .B(_1057_),
    .Y(_1058_));
 sg13g2_nor3_1 _1903_ (.A(_1006_),
    .B(_1036_),
    .C(_1051_),
    .Y(_1059_));
 sg13g2_nand2_1 _1904_ (.Y(_1060_),
    .A(_1022_),
    .B(_1059_));
 sg13g2_nor4_1 _1905_ (.A(_0994_),
    .B(_0996_),
    .C(_1056_),
    .D(_1057_),
    .Y(_1061_));
 sg13g2_a22oi_1 _1906_ (.Y(_1062_),
    .B1(_1061_),
    .B2(_0993_),
    .A2(_1060_),
    .A1(_1058_));
 sg13g2_nand2b_1 _1907_ (.Y(_1063_),
    .B(_1043_),
    .A_N(_0054_));
 sg13g2_mux2_1 _1908_ (.A0(_1031_),
    .A1(_1063_),
    .S(net469),
    .X(_1064_));
 sg13g2_nor2_1 _1909_ (.A(net497),
    .B(_1064_),
    .Y(_1065_));
 sg13g2_a21oi_2 _1910_ (.B1(_1065_),
    .Y(_1066_),
    .A2(_1003_),
    .A1(net497));
 sg13g2_mux2_1 _1911_ (.A0(_0939_),
    .A1(_1066_),
    .S(net479),
    .X(_1067_));
 sg13g2_nor2_1 _1912_ (.A(_0770_),
    .B(_1067_),
    .Y(_1068_));
 sg13g2_or2_1 _1913_ (.X(_1069_),
    .B(_1067_),
    .A(_0770_));
 sg13g2_xnor2_1 _1914_ (.Y(_1070_),
    .A(_0770_),
    .B(_1067_));
 sg13g2_nor2b_1 _1915_ (.A(_1062_),
    .B_N(_1070_),
    .Y(_1071_));
 sg13g2_a221oi_1 _1916_ (.B2(_0993_),
    .C1(_1070_),
    .B1(_1061_),
    .A1(_1058_),
    .Y(_1072_),
    .A2(_1060_));
 sg13g2_or2_1 _1917_ (.X(_1073_),
    .B(_1072_),
    .A(net486));
 sg13g2_a21oi_1 _1918_ (.A1(net486),
    .A2(net285),
    .Y(_1074_),
    .B1(net492));
 sg13g2_o21ai_1 _1919_ (.B1(_1074_),
    .Y(_0071_),
    .A1(_1071_),
    .A2(_1073_));
 sg13g2_nor2_1 _1920_ (.A(net473),
    .B(_1015_),
    .Y(_1075_));
 sg13g2_nor2_1 _1921_ (.A(_0032_),
    .B(_1045_),
    .Y(_1076_));
 sg13g2_a21o_1 _1922_ (.A2(_1076_),
    .A1(net473),
    .B1(_1075_),
    .X(_1077_));
 sg13g2_nor2_1 _1923_ (.A(net479),
    .B(_0952_),
    .Y(_1078_));
 sg13g2_and2_1 _1924_ (.A(net480),
    .B(_1077_),
    .X(_1079_));
 sg13g2_nor3_1 _1925_ (.A(\pqn_inst.multi.result[7] ),
    .B(_1078_),
    .C(_1079_),
    .Y(_1080_));
 sg13g2_inv_1 _1926_ (.Y(_1081_),
    .A(_1080_));
 sg13g2_o21ai_1 _1927_ (.B1(\pqn_inst.multi.result[7] ),
    .Y(_1082_),
    .A1(_1078_),
    .A2(_1079_));
 sg13g2_nand2b_1 _1928_ (.Y(_1083_),
    .B(_1082_),
    .A_N(_1080_));
 sg13g2_o21ai_1 _1929_ (.B1(_1083_),
    .Y(_1084_),
    .A1(_1068_),
    .A2(_1072_));
 sg13g2_nor3_1 _1930_ (.A(_1068_),
    .B(_1072_),
    .C(_1083_),
    .Y(_1085_));
 sg13g2_nor2_1 _1931_ (.A(net488),
    .B(_1085_),
    .Y(_1086_));
 sg13g2_a221oi_1 _1932_ (.B2(_1086_),
    .C1(net493),
    .B1(_1084_),
    .A1(net488),
    .Y(_0072_),
    .A2(_0769_));
 sg13g2_nand2_1 _1933_ (.Y(_1087_),
    .A(net265),
    .B(net453));
 sg13g2_nand2_1 _1934_ (.Y(_1088_),
    .A(net497),
    .B(_1032_));
 sg13g2_nor2_1 _1935_ (.A(_0032_),
    .B(_1063_),
    .Y(_1089_));
 sg13g2_a21oi_1 _1936_ (.A1(net473),
    .A2(_1089_),
    .Y(_1090_),
    .B1(net495));
 sg13g2_and2_1 _1937_ (.A(net495),
    .B(_0969_),
    .X(_1091_));
 sg13g2_a21o_1 _1938_ (.A2(_1090_),
    .A1(_1088_),
    .B1(_1091_),
    .X(_1092_));
 sg13g2_inv_1 _1939_ (.Y(_1093_),
    .A(_1092_));
 sg13g2_xnor2_1 _1940_ (.Y(_1094_),
    .A(_0768_),
    .B(_1092_));
 sg13g2_a21oi_1 _1941_ (.A1(_1069_),
    .A2(_1082_),
    .Y(_1095_),
    .B1(_1080_));
 sg13g2_a21oi_2 _1942_ (.B1(_1095_),
    .Y(_1096_),
    .A2(_1081_),
    .A1(_1072_));
 sg13g2_nor2_1 _1943_ (.A(_1094_),
    .B(_1096_),
    .Y(_1097_));
 sg13g2_a21o_1 _1944_ (.A2(_1096_),
    .A1(_1094_),
    .B1(net462),
    .X(_1098_));
 sg13g2_o21ai_1 _1945_ (.B1(_1087_),
    .Y(_0073_),
    .A1(_1097_),
    .A2(_1098_));
 sg13g2_nor2_2 _1946_ (.A(net496),
    .B(_0029_),
    .Y(_1099_));
 sg13g2_a22oi_1 _1947_ (.Y(_1100_),
    .B1(_1046_),
    .B2(_1099_),
    .A2(_0983_),
    .A1(net496));
 sg13g2_nor2_1 _1948_ (.A(net464),
    .B(_1100_),
    .Y(_1101_));
 sg13g2_xnor2_1 _1949_ (.Y(_1102_),
    .A(\pqn_inst.multi.result[9] ),
    .B(_1100_));
 sg13g2_inv_1 _1950_ (.Y(_1103_),
    .A(_1102_));
 sg13g2_a21o_1 _1951_ (.A2(_1093_),
    .A1(\pqn_inst.multi.result[8] ),
    .B1(_1097_),
    .X(_1104_));
 sg13g2_or2_1 _1952_ (.X(_1105_),
    .B(_1104_),
    .A(_1103_));
 sg13g2_a21oi_1 _1953_ (.A1(_1103_),
    .A2(_1104_),
    .Y(_1106_),
    .B1(net489));
 sg13g2_a221oi_1 _1954_ (.B2(_1106_),
    .C1(net158),
    .B1(_1105_),
    .A1(net489),
    .Y(_0074_),
    .A2(net464));
 sg13g2_nor2_1 _1955_ (.A(_1094_),
    .B(_1103_),
    .Y(_1107_));
 sg13g2_nor4_1 _1956_ (.A(_1070_),
    .B(_1083_),
    .C(_1094_),
    .D(_1103_),
    .Y(_1108_));
 sg13g2_a21oi_1 _1957_ (.A1(\pqn_inst.multi.result[8] ),
    .A2(_1093_),
    .Y(_1109_),
    .B1(_1101_));
 sg13g2_a21oi_1 _1958_ (.A1(net464),
    .A2(_1100_),
    .Y(_1110_),
    .B1(_1109_));
 sg13g2_a221oi_1 _1959_ (.B2(_1062_),
    .C1(_1110_),
    .B1(_1108_),
    .A1(_1095_),
    .Y(_1111_),
    .A2(_1107_));
 sg13g2_nor2b_1 _1960_ (.A(_1064_),
    .B_N(_1099_),
    .Y(_1112_));
 sg13g2_a21oi_2 _1961_ (.B1(_1112_),
    .Y(_1113_),
    .A2(_1004_),
    .A1(net495));
 sg13g2_nor2b_1 _1962_ (.A(_1113_),
    .B_N(net505),
    .Y(_1114_));
 sg13g2_xnor2_1 _1963_ (.Y(_1115_),
    .A(net505),
    .B(_1113_));
 sg13g2_nor2b_1 _1964_ (.A(_1115_),
    .B_N(_1111_),
    .Y(_1116_));
 sg13g2_nor2b_1 _1965_ (.A(_1111_),
    .B_N(_1115_),
    .Y(_1117_));
 sg13g2_nor3_1 _1966_ (.A(net462),
    .B(_1116_),
    .C(_1117_),
    .Y(_1118_));
 sg13g2_a21o_1 _1967_ (.A2(net453),
    .A1(net505),
    .B1(_1118_),
    .X(_0075_));
 sg13g2_a22oi_1 _1968_ (.Y(_1119_),
    .B1(_1076_),
    .B2(_1099_),
    .A2(_1017_),
    .A1(net495));
 sg13g2_and2_1 _1969_ (.A(_0766_),
    .B(_1119_),
    .X(_1120_));
 sg13g2_nand2b_1 _1970_ (.Y(_1121_),
    .B(\pqn_inst.multi.result[11] ),
    .A_N(_1119_));
 sg13g2_nor2b_1 _1971_ (.A(_1120_),
    .B_N(_1121_),
    .Y(_1122_));
 sg13g2_nor2_1 _1972_ (.A(_1114_),
    .B(_1117_),
    .Y(_1123_));
 sg13g2_or2_1 _1973_ (.X(_1124_),
    .B(_1123_),
    .A(_1122_));
 sg13g2_a21oi_1 _1974_ (.A1(_1122_),
    .A2(_1123_),
    .Y(_1125_),
    .B1(net485));
 sg13g2_a221oi_1 _1975_ (.B2(_1125_),
    .C1(net491),
    .B1(_1124_),
    .A1(net485),
    .Y(_0076_),
    .A2(_0766_));
 sg13g2_nand2_1 _1976_ (.Y(_1126_),
    .A(net504),
    .B(net453));
 sg13g2_nand2_1 _1977_ (.Y(_1127_),
    .A(_1115_),
    .B(_1122_));
 sg13g2_nand2b_1 _1978_ (.Y(_1128_),
    .B(_1121_),
    .A_N(_1114_));
 sg13g2_nor2b_1 _1979_ (.A(_1120_),
    .B_N(_1128_),
    .Y(_1129_));
 sg13g2_nand2b_1 _1980_ (.Y(_1130_),
    .B(_1128_),
    .A_N(_1120_));
 sg13g2_o21ai_1 _1981_ (.B1(_1130_),
    .Y(_1131_),
    .A1(_1111_),
    .A2(_1127_));
 sg13g2_a22oi_1 _1982_ (.Y(_1132_),
    .B1(_1089_),
    .B2(_1099_),
    .A2(_1034_),
    .A1(net495));
 sg13g2_xnor2_1 _1983_ (.Y(_1133_),
    .A(net504),
    .B(_1132_));
 sg13g2_and2_1 _1984_ (.A(_1131_),
    .B(_1133_),
    .X(_1134_));
 sg13g2_o21ai_1 _1985_ (.B1(_0830_),
    .Y(_1135_),
    .A1(_1131_),
    .A2(_1133_));
 sg13g2_o21ai_1 _1986_ (.B1(_1126_),
    .Y(_0077_),
    .A1(_1134_),
    .A2(_1135_));
 sg13g2_nor2_1 _1987_ (.A(net287),
    .B(_1132_),
    .Y(_1136_));
 sg13g2_a21oi_1 _1988_ (.A1(_1131_),
    .A2(_1133_),
    .Y(_1137_),
    .B1(_1136_));
 sg13g2_nand2_2 _1989_ (.Y(_1138_),
    .A(net496),
    .B(_1047_));
 sg13g2_xor2_1 _1990_ (.B(_1138_),
    .A(_0025_),
    .X(_1139_));
 sg13g2_or2_1 _1991_ (.X(_1140_),
    .B(_1139_),
    .A(_1137_));
 sg13g2_a21oi_1 _1992_ (.A1(_1137_),
    .A2(_1139_),
    .Y(_1141_),
    .B1(net485));
 sg13g2_a221oi_1 _1993_ (.B2(_1141_),
    .C1(net491),
    .B1(_1140_),
    .A1(net485),
    .Y(_0078_),
    .A2(_0765_));
 sg13g2_nand2_1 _1994_ (.Y(_1142_),
    .A(_1133_),
    .B(_1139_));
 sg13g2_inv_1 _1995_ (.Y(_1143_),
    .A(_1142_));
 sg13g2_nand3_1 _1996_ (.B(_1122_),
    .C(_1143_),
    .A(_1115_),
    .Y(_1144_));
 sg13g2_nor2_1 _1997_ (.A(_0765_),
    .B(_1138_),
    .Y(_1145_));
 sg13g2_a221oi_1 _1998_ (.B2(_1129_),
    .C1(_1145_),
    .B1(_1143_),
    .A1(_1136_),
    .Y(_1146_),
    .A2(_1139_));
 sg13g2_o21ai_1 _1999_ (.B1(_1146_),
    .Y(_1147_),
    .A1(_1111_),
    .A2(_1144_));
 sg13g2_nor2_2 _2000_ (.A(net480),
    .B(_1066_),
    .Y(_1148_));
 sg13g2_xnor2_1 _2001_ (.Y(_1149_),
    .A(_0026_),
    .B(_1148_));
 sg13g2_o21ai_1 _2002_ (.B1(_0830_),
    .Y(_1150_),
    .A1(_1147_),
    .A2(_1149_));
 sg13g2_a21oi_1 _2003_ (.A1(_1147_),
    .A2(_1149_),
    .Y(_1151_),
    .B1(_1150_));
 sg13g2_a21o_1 _2004_ (.A2(net453),
    .A1(net503),
    .B1(_1151_),
    .X(_0079_));
 sg13g2_a22oi_1 _2005_ (.Y(_1152_),
    .B1(_1149_),
    .B2(_1147_),
    .A2(_1148_),
    .A1(net503));
 sg13g2_nand2_1 _2006_ (.Y(_1153_),
    .A(net496),
    .B(_1077_));
 sg13g2_xnor2_1 _2007_ (.Y(_1154_),
    .A(_0028_),
    .B(_1153_));
 sg13g2_a221oi_1 _2008_ (.B2(_1147_),
    .C1(_1154_),
    .B1(_1149_),
    .A1(net503),
    .Y(_1155_),
    .A2(_1148_));
 sg13g2_nand2b_1 _2009_ (.Y(_1156_),
    .B(_1154_),
    .A_N(_1152_));
 sg13g2_nor2_1 _2010_ (.A(net485),
    .B(_1155_),
    .Y(_1157_));
 sg13g2_a221oi_1 _2011_ (.B2(_1157_),
    .C1(net491),
    .B1(_1156_),
    .A1(_0763_),
    .Y(_0080_),
    .A2(net485));
 sg13g2_nor3_1 _2012_ (.A(net177),
    .B(net489),
    .C(net454),
    .Y(_1158_));
 sg13g2_nor2_1 _2013_ (.A(net501),
    .B(_0764_),
    .Y(_1159_));
 sg13g2_nor3_1 _2014_ (.A(net491),
    .B(net178),
    .C(_1159_),
    .Y(_0081_));
 sg13g2_nor4_2 _2015_ (.A(net469),
    .B(net466),
    .C(net485),
    .Y(_1160_),
    .D(net456));
 sg13g2_a21oi_1 _2016_ (.A1(net501),
    .A2(_0764_),
    .Y(_1161_),
    .B1(net499));
 sg13g2_nor3_1 _2017_ (.A(net491),
    .B(_1160_),
    .C(_1161_),
    .Y(_0082_));
 sg13g2_xnor2_1 _2018_ (.Y(_1162_),
    .A(net259),
    .B(_0787_));
 sg13g2_nor3_1 _2019_ (.A(net485),
    .B(net454),
    .C(_1162_),
    .Y(_1163_));
 sg13g2_nor2_1 _2020_ (.A(net497),
    .B(_0764_),
    .Y(_1164_));
 sg13g2_nor3_1 _2021_ (.A(net491),
    .B(_1163_),
    .C(_1164_),
    .Y(_0083_));
 sg13g2_a21oi_1 _2022_ (.A1(net498),
    .A2(_1160_),
    .Y(_1165_),
    .B1(net495));
 sg13g2_nor2_1 _2023_ (.A(net491),
    .B(net254),
    .Y(_0084_));
 sg13g2_nand2_1 _2024_ (.Y(_0085_),
    .A(net529),
    .B(net463));
 sg13g2_nor2_1 _2025_ (.A(\pqn_inst.stage[3] ),
    .B(net463),
    .Y(_1166_));
 sg13g2_or2_2 _2026_ (.X(_1167_),
    .B(\pqn_inst.stage[1] ),
    .A(\pqn_inst.stage[2] ));
 sg13g2_a21oi_2 _2027_ (.B1(net463),
    .Y(_1168_),
    .A2(_1167_),
    .A1(\pqn_inst.stage[3] ));
 sg13g2_nor2b_2 _2028_ (.A(\pqn_inst.stage[3] ),
    .B_N(\pqn_inst.stage[2] ),
    .Y(_1169_));
 sg13g2_nor2_2 _2029_ (.A(net481),
    .B(net483),
    .Y(_1170_));
 sg13g2_and2_2 _2030_ (.A(_0716_),
    .B(_1169_),
    .X(_1171_));
 sg13g2_and2_2 _2031_ (.A(_1169_),
    .B(_1170_),
    .X(_1172_));
 sg13g2_nand2_2 _2032_ (.Y(_1173_),
    .A(_1169_),
    .B(_1170_));
 sg13g2_nor2_1 _2033_ (.A(_0715_),
    .B(_1167_),
    .Y(_1174_));
 sg13g2_and2_1 _2034_ (.A(\pqn_inst.stage[1] ),
    .B(net482),
    .X(_1175_));
 sg13g2_a22oi_1 _2035_ (.Y(_1176_),
    .B1(_1175_),
    .B2(_1169_),
    .A2(_1174_),
    .A1(_0716_));
 sg13g2_and2_2 _2036_ (.A(_1168_),
    .B(_1176_),
    .X(_1177_));
 sg13g2_nand2_1 _2037_ (.Y(_1178_),
    .A(_1168_),
    .B(_1176_));
 sg13g2_nand2_2 _2038_ (.Y(_1179_),
    .A(_1173_),
    .B(_1177_));
 sg13g2_nor2_2 _2039_ (.A(\pqn_inst.stage[3] ),
    .B(\pqn_inst.stage[2] ),
    .Y(_1180_));
 sg13g2_nor2_2 _2040_ (.A(\pqn_inst.stage[3] ),
    .B(_1167_),
    .Y(_1181_));
 sg13g2_and2_1 _2041_ (.A(_1170_),
    .B(_1180_),
    .X(_1182_));
 sg13g2_nand2_1 _2042_ (.Y(_1183_),
    .A(_1170_),
    .B(_1180_));
 sg13g2_nor2_1 _2043_ (.A(net410),
    .B(net450),
    .Y(_1184_));
 sg13g2_and2_2 _2044_ (.A(net481),
    .B(_1180_),
    .X(_1185_));
 sg13g2_nand2_1 _2045_ (.Y(_1186_),
    .A(net481),
    .B(_1180_));
 sg13g2_nor2_1 _2046_ (.A(net482),
    .B(_1186_),
    .Y(_1187_));
 sg13g2_nand2_1 _2047_ (.Y(_1188_),
    .A(_0716_),
    .B(net447));
 sg13g2_nand2_2 _2048_ (.Y(_1189_),
    .A(net481),
    .B(_1171_));
 sg13g2_and2_1 _2049_ (.A(net482),
    .B(_1169_),
    .X(_1190_));
 sg13g2_nand2_1 _2050_ (.Y(_1191_),
    .A(net482),
    .B(_1169_));
 sg13g2_nand2b_1 _2051_ (.Y(_1192_),
    .B(_1169_),
    .A_N(net481));
 sg13g2_nor2_1 _2052_ (.A(net481),
    .B(net443),
    .Y(_1193_));
 sg13g2_nand2b_2 _2053_ (.Y(_1194_),
    .B(net444),
    .A_N(net481));
 sg13g2_nand2_1 _2054_ (.Y(_1195_),
    .A(_1189_),
    .B(_1194_));
 sg13g2_nor2_2 _2055_ (.A(net431),
    .B(net417),
    .Y(_1196_));
 sg13g2_inv_1 _2056_ (.Y(_1197_),
    .A(net408));
 sg13g2_nor2_2 _2057_ (.A(_0716_),
    .B(net446),
    .Y(_1198_));
 sg13g2_nand2_2 _2058_ (.Y(_1199_),
    .A(_1175_),
    .B(_1180_));
 sg13g2_nand3_1 _2059_ (.B(_1194_),
    .C(_1199_),
    .A(_1189_),
    .Y(_1200_));
 sg13g2_inv_1 _2060_ (.Y(_1201_),
    .A(net416));
 sg13g2_nor2_1 _2061_ (.A(_0016_),
    .B(_1200_),
    .Y(_1202_));
 sg13g2_nor2_1 _2062_ (.A(_0017_),
    .B(net446),
    .Y(_1203_));
 sg13g2_o21ai_1 _2063_ (.B1(net425),
    .Y(_1204_),
    .A1(_1202_),
    .A2(_1203_));
 sg13g2_o21ai_1 _2064_ (.B1(_1204_),
    .Y(_1205_),
    .A1(_0003_),
    .A2(net408));
 sg13g2_a22oi_1 _2065_ (.Y(_1206_),
    .B1(net402),
    .B2(_1205_),
    .A2(net409),
    .A1(net148));
 sg13g2_nor2_1 _2066_ (.A(net516),
    .B(net149),
    .Y(_0086_));
 sg13g2_nand2_1 _2067_ (.Y(_1207_),
    .A(net135),
    .B(net409));
 sg13g2_nand2_1 _2068_ (.Y(_1208_),
    .A(net482),
    .B(_0019_));
 sg13g2_a22oi_1 _2069_ (.Y(_1209_),
    .B1(_1208_),
    .B2(net447),
    .A2(net417),
    .A1(_0780_));
 sg13g2_o21ai_1 _2070_ (.B1(_1209_),
    .Y(_1210_),
    .A1(_0018_),
    .A2(_1200_));
 sg13g2_nand2_1 _2071_ (.Y(_1211_),
    .A(_0004_),
    .B(net431));
 sg13g2_nand3_1 _2072_ (.B(_1210_),
    .C(_1211_),
    .A(net402),
    .Y(_1212_));
 sg13g2_a21oi_1 _2073_ (.A1(_1207_),
    .A2(_1212_),
    .Y(_0087_),
    .B1(net517));
 sg13g2_a22oi_1 _2074_ (.Y(_1213_),
    .B1(_1201_),
    .B2(_0049_),
    .A2(_1185_),
    .A1(_0020_));
 sg13g2_nor2_1 _2075_ (.A(net432),
    .B(_1213_),
    .Y(_1214_));
 sg13g2_a21oi_1 _2076_ (.A1(_0006_),
    .A2(_1197_),
    .Y(_1215_),
    .B1(_1214_));
 sg13g2_a22oi_1 _2077_ (.Y(_1216_),
    .B1(net402),
    .B2(_1215_),
    .A2(net409),
    .A1(net193));
 sg13g2_nor2_1 _2078_ (.A(net511),
    .B(net194),
    .Y(_0088_));
 sg13g2_nand3_1 _2079_ (.B(_1189_),
    .C(_1194_),
    .A(_0052_),
    .Y(_1217_));
 sg13g2_a21oi_1 _2080_ (.A1(_0007_),
    .A2(_1195_),
    .Y(_1218_),
    .B1(_1198_));
 sg13g2_a21oi_1 _2081_ (.A1(net482),
    .A2(_0021_),
    .Y(_1219_),
    .B1(net446));
 sg13g2_a21oi_1 _2082_ (.A1(_1217_),
    .A2(_1218_),
    .Y(_1220_),
    .B1(_1219_));
 sg13g2_a21oi_1 _2083_ (.A1(_0007_),
    .A2(net431),
    .Y(_1221_),
    .B1(_1220_));
 sg13g2_a22oi_1 _2084_ (.Y(_1222_),
    .B1(net401),
    .B2(_1221_),
    .A2(net410),
    .A1(net152));
 sg13g2_nor2_1 _2085_ (.A(net511),
    .B(net153),
    .Y(_0089_));
 sg13g2_nor2_1 _2086_ (.A(_0053_),
    .B(net416),
    .Y(_1223_));
 sg13g2_nor2_1 _2087_ (.A(_0023_),
    .B(_1199_),
    .Y(_1224_));
 sg13g2_o21ai_1 _2088_ (.B1(net425),
    .Y(_1225_),
    .A1(_1223_),
    .A2(_1224_));
 sg13g2_o21ai_1 _2089_ (.B1(_1225_),
    .Y(_1226_),
    .A1(_0022_),
    .A2(_1196_));
 sg13g2_a22oi_1 _2090_ (.Y(_1227_),
    .B1(net402),
    .B2(_1226_),
    .A2(_1179_),
    .A1(net146));
 sg13g2_nor2_1 _2091_ (.A(net516),
    .B(net147),
    .Y(_0090_));
 sg13g2_nand2_1 _2092_ (.Y(_1228_),
    .A(_0771_),
    .B(_1185_));
 sg13g2_o21ai_1 _2093_ (.B1(_1228_),
    .Y(_1229_),
    .A1(\pqn_inst.n[5] ),
    .A2(net416));
 sg13g2_o21ai_1 _2094_ (.B1(net402),
    .Y(_1230_),
    .A1(uo_out[5]),
    .A2(_1196_));
 sg13g2_a21oi_1 _2095_ (.A1(net426),
    .A2(_1229_),
    .Y(_1231_),
    .B1(_1230_));
 sg13g2_nor2_2 _2096_ (.A(_1179_),
    .B(_1183_),
    .Y(_1232_));
 sg13g2_a221oi_1 _2097_ (.B2(net2),
    .C1(_1231_),
    .B1(_1232_),
    .A1(net233),
    .Y(_1233_),
    .A2(net409));
 sg13g2_nor2_1 _2098_ (.A(net516),
    .B(_1233_),
    .Y(_0091_));
 sg13g2_nand2_1 _2099_ (.Y(_1234_),
    .A(_0770_),
    .B(net447));
 sg13g2_o21ai_1 _2100_ (.B1(_1234_),
    .Y(_1235_),
    .A1(\pqn_inst.n[6] ),
    .A2(net416));
 sg13g2_o21ai_1 _2101_ (.B1(net402),
    .Y(_1236_),
    .A1(uo_out[6]),
    .A2(_1196_));
 sg13g2_a21oi_1 _2102_ (.A1(net425),
    .A2(_1235_),
    .Y(_1237_),
    .B1(_1236_));
 sg13g2_a221oi_1 _2103_ (.B2(net3),
    .C1(_1237_),
    .B1(_1232_),
    .A1(net232),
    .Y(_1238_),
    .A2(net409));
 sg13g2_nor2_1 _2104_ (.A(net518),
    .B(_1238_),
    .Y(_0092_));
 sg13g2_nand2_1 _2105_ (.Y(_1239_),
    .A(_0769_),
    .B(net447));
 sg13g2_o21ai_1 _2106_ (.B1(_1239_),
    .Y(_1240_),
    .A1(\pqn_inst.n[7] ),
    .A2(net416));
 sg13g2_o21ai_1 _2107_ (.B1(net402),
    .Y(_1241_),
    .A1(uo_out[7]),
    .A2(net408));
 sg13g2_a21oi_1 _2108_ (.A1(net426),
    .A2(_1240_),
    .Y(_1242_),
    .B1(_1241_));
 sg13g2_a221oi_1 _2109_ (.B2(net4),
    .C1(_1242_),
    .B1(_1232_),
    .A1(net221),
    .Y(_1243_),
    .A2(net409));
 sg13g2_nor2_1 _2110_ (.A(net515),
    .B(_1243_),
    .Y(_0093_));
 sg13g2_nand2_1 _2111_ (.Y(_1244_),
    .A(_0768_),
    .B(net447));
 sg13g2_o21ai_1 _2112_ (.B1(_1244_),
    .Y(_1245_),
    .A1(\pqn_inst.n[8] ),
    .A2(net416));
 sg13g2_o21ai_1 _2113_ (.B1(net402),
    .Y(_1246_),
    .A1(uio_out[0]),
    .A2(net408));
 sg13g2_a21oi_1 _2114_ (.A1(net427),
    .A2(_1245_),
    .Y(_1247_),
    .B1(_1246_));
 sg13g2_a221oi_1 _2115_ (.B2(net5),
    .C1(_1247_),
    .B1(_1232_),
    .A1(net220),
    .Y(_1248_),
    .A2(net409));
 sg13g2_nor2_1 _2116_ (.A(net516),
    .B(_1248_),
    .Y(_0094_));
 sg13g2_nand2_1 _2117_ (.Y(_1249_),
    .A(_0767_),
    .B(net447));
 sg13g2_o21ai_1 _2118_ (.B1(_1249_),
    .Y(_1250_),
    .A1(\pqn_inst.n[9] ),
    .A2(net416));
 sg13g2_o21ai_1 _2119_ (.B1(net401),
    .Y(_1251_),
    .A1(uio_out[1]),
    .A2(net408));
 sg13g2_a21oi_1 _2120_ (.A1(net427),
    .A2(_1250_),
    .Y(_1252_),
    .B1(_1251_));
 sg13g2_a221oi_1 _2121_ (.B2(net6),
    .C1(_1252_),
    .B1(_1232_),
    .A1(net234),
    .Y(_1253_),
    .A2(net409));
 sg13g2_nor2_1 _2122_ (.A(net516),
    .B(_1253_),
    .Y(_0095_));
 sg13g2_nand2_1 _2123_ (.Y(_1254_),
    .A(_0717_),
    .B(_1201_));
 sg13g2_o21ai_1 _2124_ (.B1(_1254_),
    .Y(_1255_),
    .A1(net505),
    .A2(_1199_));
 sg13g2_o21ai_1 _2125_ (.B1(net401),
    .Y(_1256_),
    .A1(uio_out[2]),
    .A2(net408));
 sg13g2_a21o_1 _2126_ (.A2(_1255_),
    .A1(net427),
    .B1(_1256_),
    .X(_1257_));
 sg13g2_a22oi_1 _2127_ (.Y(_1258_),
    .B1(_1232_),
    .B2(net7),
    .A2(net410),
    .A1(net224));
 sg13g2_nand3_1 _2128_ (.B(_1257_),
    .C(_1258_),
    .A(net526),
    .Y(_0096_));
 sg13g2_nand2_1 _2129_ (.Y(_1259_),
    .A(_0766_),
    .B(net447));
 sg13g2_o21ai_1 _2130_ (.B1(_1259_),
    .Y(_1260_),
    .A1(net484),
    .A2(net416));
 sg13g2_o21ai_1 _2131_ (.B1(net401),
    .Y(_1261_),
    .A1(uio_out[3]),
    .A2(net408));
 sg13g2_a21o_1 _2132_ (.A2(_1260_),
    .A1(net427),
    .B1(_1261_),
    .X(_1262_));
 sg13g2_a22oi_1 _2133_ (.Y(_1263_),
    .B1(_1232_),
    .B2(net8),
    .A2(net410),
    .A1(net219));
 sg13g2_nand3_1 _2134_ (.B(_1262_),
    .C(_1263_),
    .A(net526),
    .Y(_0097_));
 sg13g2_o21ai_1 _2135_ (.B1(_1199_),
    .Y(_1264_),
    .A1(_0779_),
    .A2(net417));
 sg13g2_a21oi_1 _2136_ (.A1(_0014_),
    .A2(net417),
    .Y(_1265_),
    .B1(_1264_));
 sg13g2_a21oi_1 _2137_ (.A1(net483),
    .A2(_0024_),
    .Y(_1266_),
    .B1(net446));
 sg13g2_nand2_1 _2138_ (.Y(_1267_),
    .A(_0014_),
    .B(net428));
 sg13g2_o21ai_1 _2139_ (.B1(net401),
    .Y(_1268_),
    .A1(_1265_),
    .A2(_1266_));
 sg13g2_nor2b_1 _2140_ (.A(_1268_),
    .B_N(_1267_),
    .Y(_1269_));
 sg13g2_a21oi_1 _2141_ (.A1(net166),
    .A2(net410),
    .Y(_1270_),
    .B1(_1269_));
 sg13g2_nor2_1 _2142_ (.A(net510),
    .B(net167),
    .Y(_0098_));
 sg13g2_mux2_1 _2143_ (.A0(_0001_),
    .A1(_0015_),
    .S(net417),
    .X(_1271_));
 sg13g2_nand2_2 _2144_ (.Y(_1272_),
    .A(_0015_),
    .B(net429));
 sg13g2_a22oi_1 _2145_ (.Y(_1273_),
    .B1(_1271_),
    .B2(net446),
    .A2(_1198_),
    .A1(_0025_));
 sg13g2_nand3_1 _2146_ (.B(_1272_),
    .C(_1273_),
    .A(net401),
    .Y(_1274_));
 sg13g2_a21oi_1 _2147_ (.A1(net179),
    .A2(net410),
    .Y(_1275_),
    .B1(net510));
 sg13g2_nand2_1 _2148_ (.Y(_0099_),
    .A(_1274_),
    .B(_1275_));
 sg13g2_a21oi_1 _2149_ (.A1(_0781_),
    .A2(net417),
    .Y(_1276_),
    .B1(net447));
 sg13g2_o21ai_1 _2150_ (.B1(_1276_),
    .Y(_1277_),
    .A1(_0002_),
    .A2(net417));
 sg13g2_nand2_1 _2151_ (.Y(_1278_),
    .A(_0026_),
    .B(_1198_));
 sg13g2_nand2_2 _2152_ (.Y(_1279_),
    .A(_0005_),
    .B(net428));
 sg13g2_nand4_1 _2153_ (.B(_1277_),
    .C(_1278_),
    .A(net401),
    .Y(_1280_),
    .D(_1279_));
 sg13g2_a21oi_1 _2154_ (.A1(net181),
    .A2(net410),
    .Y(_1281_),
    .B1(net511));
 sg13g2_nand2_1 _2155_ (.Y(_0100_),
    .A(_1280_),
    .B(_1281_));
 sg13g2_mux2_1 _2156_ (.A0(_0027_),
    .A1(_0050_),
    .S(net417),
    .X(_1282_));
 sg13g2_nand2_2 _2157_ (.Y(_1283_),
    .A(_0050_),
    .B(net428));
 sg13g2_a22oi_1 _2158_ (.Y(_1284_),
    .B1(_1282_),
    .B2(net446),
    .A2(_1198_),
    .A1(_0028_));
 sg13g2_nand3_1 _2159_ (.B(_1283_),
    .C(_1284_),
    .A(net401),
    .Y(_1285_));
 sg13g2_a21oi_1 _2160_ (.A1(net195),
    .A2(net410),
    .Y(_1286_),
    .B1(net509));
 sg13g2_nand2_1 _2161_ (.Y(_0101_),
    .A(_1285_),
    .B(_1286_));
 sg13g2_or2_1 _2162_ (.X(_1287_),
    .B(_1181_),
    .A(_1171_));
 sg13g2_nor4_2 _2163_ (.A(\pqn_inst.stage[3] ),
    .B(net463),
    .C(_1185_),
    .Y(_1288_),
    .D(_1193_));
 sg13g2_nand3_1 _2164_ (.B(net446),
    .C(_1194_),
    .A(_1166_),
    .Y(_1289_));
 sg13g2_o21ai_1 _2165_ (.B1(_1288_),
    .Y(_1290_),
    .A1(net519),
    .A2(_1287_));
 sg13g2_a21oi_1 _2166_ (.A1(_0773_),
    .A2(_1287_),
    .Y(_1291_),
    .B1(_1290_));
 sg13g2_o21ai_1 _2167_ (.B1(net528),
    .Y(_1292_),
    .A1(net200),
    .A2(_1291_));
 sg13g2_a21oi_1 _2168_ (.A1(net200),
    .A2(_1291_),
    .Y(_0102_),
    .B1(_1292_));
 sg13g2_nand2_1 _2169_ (.Y(_1293_),
    .A(\pqn_inst.v[1] ),
    .B(net508));
 sg13g2_nor2_1 _2170_ (.A(\pqn_inst.v[1] ),
    .B(net508),
    .Y(_1294_));
 sg13g2_xor2_1 _2171_ (.B(net508),
    .A(\pqn_inst.v[1] ),
    .X(_1295_));
 sg13g2_nor2b_1 _2172_ (.A(\pqn_inst.v[0] ),
    .B_N(\pqn_inst.multi.result[0] ),
    .Y(_1296_));
 sg13g2_xnor2_1 _2173_ (.Y(_1297_),
    .A(_1295_),
    .B(_1296_));
 sg13g2_a21oi_2 _2174_ (.B1(_1171_),
    .Y(_1298_),
    .A2(_1181_),
    .A1(net482));
 sg13g2_a21o_1 _2175_ (.A2(_1181_),
    .A1(net482),
    .B1(_1171_),
    .X(_1299_));
 sg13g2_nand2_1 _2176_ (.Y(_1300_),
    .A(\pqn_inst.v[0] ),
    .B(\pqn_inst.multi.result[0] ));
 sg13g2_xnor2_1 _2177_ (.Y(_1301_),
    .A(_1295_),
    .B(_1300_));
 sg13g2_o21ai_1 _2178_ (.B1(\pqn_inst.v[1] ),
    .Y(_1302_),
    .A1(\pqn_inst.v[0] ),
    .A2(net524));
 sg13g2_nand3_1 _2179_ (.B(_0738_),
    .C(net519),
    .A(_0737_),
    .Y(_1303_));
 sg13g2_nand3_1 _2180_ (.B(_1302_),
    .C(_1303_),
    .A(_1298_),
    .Y(_1304_));
 sg13g2_a21oi_1 _2181_ (.A1(net422),
    .A2(_1301_),
    .Y(_1305_),
    .B1(net451));
 sg13g2_a22oi_1 _2182_ (.Y(_1306_),
    .B1(_1304_),
    .B2(_1305_),
    .A2(_1297_),
    .A1(net452));
 sg13g2_o21ai_1 _2183_ (.B1(net528),
    .Y(_1307_),
    .A1(net414),
    .A2(_1306_));
 sg13g2_a21oi_1 _2184_ (.A1(_0737_),
    .A2(net414),
    .Y(_0103_),
    .B1(_1307_));
 sg13g2_and2_1 _2185_ (.A(\pqn_inst.v[2] ),
    .B(\pqn_inst.multi.result[2] ),
    .X(_1308_));
 sg13g2_xnor2_1 _2186_ (.Y(_1309_),
    .A(\pqn_inst.v[2] ),
    .B(\pqn_inst.multi.result[2] ));
 sg13g2_inv_1 _2187_ (.Y(_1310_),
    .A(_1309_));
 sg13g2_nand2b_1 _2188_ (.Y(_1311_),
    .B(\pqn_inst.v[1] ),
    .A_N(net508));
 sg13g2_o21ai_1 _2189_ (.B1(_1311_),
    .Y(_1312_),
    .A1(_1295_),
    .A2(_1296_));
 sg13g2_xnor2_1 _2190_ (.Y(_1313_),
    .A(_1309_),
    .B(_1312_));
 sg13g2_o21ai_1 _2191_ (.B1(_1293_),
    .Y(_1314_),
    .A1(_1294_),
    .A2(_1300_));
 sg13g2_o21ai_1 _2192_ (.B1(net422),
    .Y(_1315_),
    .A1(_1310_),
    .A2(_1314_));
 sg13g2_a21o_1 _2193_ (.A2(_1314_),
    .A1(_1310_),
    .B1(_1315_),
    .X(_1316_));
 sg13g2_nand2b_1 _2194_ (.Y(_1317_),
    .B(\pqn_inst.v[2] ),
    .A_N(net524));
 sg13g2_xor2_1 _2195_ (.B(net524),
    .A(\pqn_inst.v[2] ),
    .X(_1318_));
 sg13g2_xor2_1 _2196_ (.B(_1318_),
    .A(_1302_),
    .X(_1319_));
 sg13g2_a21oi_1 _2197_ (.A1(_1298_),
    .A2(_1319_),
    .Y(_1320_),
    .B1(net451));
 sg13g2_a22oi_1 _2198_ (.Y(_1321_),
    .B1(_1316_),
    .B2(_1320_),
    .A2(_1313_),
    .A1(net451));
 sg13g2_o21ai_1 _2199_ (.B1(net1),
    .Y(_1322_),
    .A1(net415),
    .A2(_1321_));
 sg13g2_a21oi_1 _2200_ (.A1(_0736_),
    .A2(net414),
    .Y(_0104_),
    .B1(_1322_));
 sg13g2_nand2_1 _2201_ (.Y(_1323_),
    .A(\pqn_inst.v[3] ),
    .B(\pqn_inst.multi.result[3] ));
 sg13g2_xor2_1 _2202_ (.B(\pqn_inst.multi.result[3] ),
    .A(\pqn_inst.v[3] ),
    .X(_1324_));
 sg13g2_xnor2_1 _2203_ (.Y(_1325_),
    .A(\pqn_inst.v[3] ),
    .B(\pqn_inst.multi.result[3] ));
 sg13g2_a21oi_2 _2204_ (.B1(_1308_),
    .Y(_1326_),
    .A2(_1314_),
    .A1(_1310_));
 sg13g2_nand2b_1 _2205_ (.Y(_1327_),
    .B(_1324_),
    .A_N(_1326_));
 sg13g2_xnor2_1 _2206_ (.Y(_1328_),
    .A(_1325_),
    .B(_1326_));
 sg13g2_o21ai_1 _2207_ (.B1(_1317_),
    .Y(_1329_),
    .A1(_1302_),
    .A2(_1318_));
 sg13g2_and2_1 _2208_ (.A(\pqn_inst.v[3] ),
    .B(_1329_),
    .X(_1330_));
 sg13g2_nor2_2 _2209_ (.A(\pqn_inst.v[3] ),
    .B(_1329_),
    .Y(_1331_));
 sg13g2_o21ai_1 _2210_ (.B1(_1298_),
    .Y(_1332_),
    .A1(_1330_),
    .A2(_1331_));
 sg13g2_o21ai_1 _2211_ (.B1(_1332_),
    .Y(_1333_),
    .A1(net424),
    .A2(_1328_));
 sg13g2_nand2_1 _2212_ (.Y(_1334_),
    .A(net448),
    .B(_1333_));
 sg13g2_nor2_1 _2213_ (.A(_0736_),
    .B(\pqn_inst.multi.result[2] ),
    .Y(_1335_));
 sg13g2_a21oi_1 _2214_ (.A1(_1309_),
    .A2(_1312_),
    .Y(_1336_),
    .B1(_1335_));
 sg13g2_xnor2_1 _2215_ (.Y(_1337_),
    .A(_1325_),
    .B(_1336_));
 sg13g2_a21oi_1 _2216_ (.A1(net451),
    .A2(_1337_),
    .Y(_1338_),
    .B1(net415));
 sg13g2_a221oi_1 _2217_ (.B2(_1338_),
    .C1(net515),
    .B1(_1334_),
    .A1(_0735_),
    .Y(_0105_),
    .A2(net414));
 sg13g2_and2_1 _2218_ (.A(\pqn_inst.v[4] ),
    .B(\pqn_inst.multi.result[4] ),
    .X(_1339_));
 sg13g2_xnor2_1 _2219_ (.Y(_1340_),
    .A(\pqn_inst.v[4] ),
    .B(net506));
 sg13g2_inv_1 _2220_ (.Y(_1341_),
    .A(_1340_));
 sg13g2_and2_1 _2221_ (.A(_1323_),
    .B(_1327_),
    .X(_1342_));
 sg13g2_o21ai_1 _2222_ (.B1(_1323_),
    .Y(_1343_),
    .A1(_1325_),
    .A2(_1326_));
 sg13g2_nand2_1 _2223_ (.Y(_1344_),
    .A(_1341_),
    .B(_1343_));
 sg13g2_a21oi_1 _2224_ (.A1(_1340_),
    .A2(_1342_),
    .Y(_1345_),
    .B1(net424));
 sg13g2_xor2_1 _2225_ (.B(net524),
    .A(\pqn_inst.v[4] ),
    .X(_1346_));
 sg13g2_nand2_1 _2226_ (.Y(_1347_),
    .A(_1331_),
    .B(_1346_));
 sg13g2_nor2_1 _2227_ (.A(_1331_),
    .B(_1346_),
    .Y(_1348_));
 sg13g2_nor2_1 _2228_ (.A(net422),
    .B(_1348_),
    .Y(_1349_));
 sg13g2_a22oi_1 _2229_ (.Y(_1350_),
    .B1(_1347_),
    .B2(_1349_),
    .A2(_1345_),
    .A1(_1344_));
 sg13g2_or2_1 _2230_ (.X(_1351_),
    .B(_1350_),
    .A(net451));
 sg13g2_nand2_1 _2231_ (.Y(_1352_),
    .A(\pqn_inst.v[3] ),
    .B(_0772_));
 sg13g2_o21ai_1 _2232_ (.B1(_1352_),
    .Y(_1353_),
    .A1(_1324_),
    .A2(_1336_));
 sg13g2_and2_1 _2233_ (.A(_1340_),
    .B(_1353_),
    .X(_1354_));
 sg13g2_o21ai_1 _2234_ (.B1(net451),
    .Y(_1355_),
    .A1(_1340_),
    .A2(_1353_));
 sg13g2_nor2_1 _2235_ (.A(_1354_),
    .B(_1355_),
    .Y(_1356_));
 sg13g2_nor2_1 _2236_ (.A(net415),
    .B(_1356_),
    .Y(_1357_));
 sg13g2_a221oi_1 _2237_ (.B2(_1357_),
    .C1(net515),
    .B1(_1351_),
    .A1(_0734_),
    .Y(_0106_),
    .A2(net414));
 sg13g2_xnor2_1 _2238_ (.Y(_1358_),
    .A(\pqn_inst.v[5] ),
    .B(net524));
 sg13g2_inv_1 _2239_ (.Y(_1359_),
    .A(_1358_));
 sg13g2_a21oi_1 _2240_ (.A1(\pqn_inst.v[4] ),
    .A2(net519),
    .Y(_1360_),
    .B1(_1348_));
 sg13g2_nor2_1 _2241_ (.A(\pqn_inst.v[5] ),
    .B(\pqn_inst.multi.result[5] ),
    .Y(_1361_));
 sg13g2_xnor2_1 _2242_ (.Y(_1362_),
    .A(\pqn_inst.v[5] ),
    .B(\pqn_inst.multi.result[5] ));
 sg13g2_nand2b_1 _2243_ (.Y(_1363_),
    .B(_1344_),
    .A_N(_1339_));
 sg13g2_a21oi_1 _2244_ (.A1(_1362_),
    .A2(_1363_),
    .Y(_1364_),
    .B1(net424));
 sg13g2_o21ai_1 _2245_ (.B1(_1364_),
    .Y(_1365_),
    .A1(_1362_),
    .A2(_1363_));
 sg13g2_a21oi_1 _2246_ (.A1(_1358_),
    .A2(_1360_),
    .Y(_0171_),
    .B1(net422));
 sg13g2_o21ai_1 _2247_ (.B1(_0171_),
    .Y(_0172_),
    .A1(_1358_),
    .A2(_1360_));
 sg13g2_nand3_1 _2248_ (.B(_1365_),
    .C(_0172_),
    .A(net448),
    .Y(_0173_));
 sg13g2_nor2_1 _2249_ (.A(_0734_),
    .B(net506),
    .Y(_0174_));
 sg13g2_nor2_1 _2250_ (.A(_1354_),
    .B(_0174_),
    .Y(_0175_));
 sg13g2_xnor2_1 _2251_ (.Y(_0176_),
    .A(_1362_),
    .B(_0175_));
 sg13g2_a21oi_1 _2252_ (.A1(net451),
    .A2(_0176_),
    .Y(_0177_),
    .B1(net414));
 sg13g2_a221oi_1 _2253_ (.B2(_0177_),
    .C1(net515),
    .B1(_0173_),
    .A1(_0733_),
    .Y(_0107_),
    .A2(net414));
 sg13g2_nor2_1 _2254_ (.A(_0732_),
    .B(_0770_),
    .Y(_0178_));
 sg13g2_xnor2_1 _2255_ (.Y(_0179_),
    .A(\pqn_inst.v[6] ),
    .B(\pqn_inst.multi.result[6] ));
 sg13g2_inv_1 _2256_ (.Y(_0180_),
    .A(_0179_));
 sg13g2_a221oi_1 _2257_ (.B2(_1343_),
    .C1(_1339_),
    .B1(_1341_),
    .A1(\pqn_inst.v[5] ),
    .Y(_0181_),
    .A2(\pqn_inst.multi.result[5] ));
 sg13g2_nor3_1 _2258_ (.A(_1361_),
    .B(_0179_),
    .C(_0181_),
    .Y(_0182_));
 sg13g2_or3_1 _2259_ (.A(_1361_),
    .B(_0179_),
    .C(_0181_),
    .X(_0183_));
 sg13g2_o21ai_1 _2260_ (.B1(_0179_),
    .Y(_0184_),
    .A1(_1361_),
    .A2(_0181_));
 sg13g2_and2_1 _2261_ (.A(_0183_),
    .B(_0184_),
    .X(_0185_));
 sg13g2_xor2_1 _2262_ (.B(net525),
    .A(\pqn_inst.v[6] ),
    .X(_0186_));
 sg13g2_a21oi_1 _2263_ (.A1(_0733_),
    .A2(_0734_),
    .Y(_0187_),
    .B1(net525));
 sg13g2_a21oi_1 _2264_ (.A1(_1348_),
    .A2(_1358_),
    .Y(_0188_),
    .B1(_0187_));
 sg13g2_nor2_1 _2265_ (.A(_0186_),
    .B(_0188_),
    .Y(_0189_));
 sg13g2_a21oi_1 _2266_ (.A1(_0186_),
    .A2(_0188_),
    .Y(_0190_),
    .B1(net423));
 sg13g2_nor2b_1 _2267_ (.A(_0189_),
    .B_N(_0190_),
    .Y(_0191_));
 sg13g2_a21oi_1 _2268_ (.A1(net423),
    .A2(_0185_),
    .Y(_0192_),
    .B1(_0191_));
 sg13g2_or2_1 _2269_ (.X(_0193_),
    .B(_0192_),
    .A(net452));
 sg13g2_nor2_1 _2270_ (.A(\pqn_inst.v[5] ),
    .B(_0771_),
    .Y(_0194_));
 sg13g2_a221oi_1 _2271_ (.B2(_1353_),
    .C1(_0174_),
    .B1(_1340_),
    .A1(\pqn_inst.v[5] ),
    .Y(_0195_),
    .A2(_0771_));
 sg13g2_or3_1 _2272_ (.A(_0180_),
    .B(_0194_),
    .C(_0195_),
    .X(_0196_));
 sg13g2_o21ai_1 _2273_ (.B1(_0180_),
    .Y(_0197_),
    .A1(_0194_),
    .A2(_0195_));
 sg13g2_and2_1 _2274_ (.A(net451),
    .B(_0197_),
    .X(_0198_));
 sg13g2_a21oi_1 _2275_ (.A1(_0196_),
    .A2(_0198_),
    .Y(_0199_),
    .B1(net414));
 sg13g2_a221oi_1 _2276_ (.B2(_0199_),
    .C1(net515),
    .B1(_0193_),
    .A1(_0732_),
    .Y(_0108_),
    .A2(net415));
 sg13g2_xnor2_1 _2277_ (.Y(_0200_),
    .A(\pqn_inst.v[7] ),
    .B(net524));
 sg13g2_a21oi_1 _2278_ (.A1(\pqn_inst.v[6] ),
    .A2(net519),
    .Y(_0201_),
    .B1(_0189_));
 sg13g2_nand2_1 _2279_ (.Y(_0202_),
    .A(\pqn_inst.v[7] ),
    .B(\pqn_inst.multi.result[7] ));
 sg13g2_xnor2_1 _2280_ (.Y(_0203_),
    .A(\pqn_inst.v[7] ),
    .B(\pqn_inst.multi.result[7] ));
 sg13g2_inv_1 _2281_ (.Y(_0204_),
    .A(_0203_));
 sg13g2_o21ai_1 _2282_ (.B1(_0204_),
    .Y(_0205_),
    .A1(_0178_),
    .A2(_0182_));
 sg13g2_nand3b_1 _2283_ (.B(_0183_),
    .C(_0203_),
    .Y(_0206_),
    .A_N(_0178_));
 sg13g2_nand2_1 _2284_ (.Y(_0207_),
    .A(_0205_),
    .B(_0206_));
 sg13g2_or2_1 _2285_ (.X(_0208_),
    .B(_0201_),
    .A(_0200_));
 sg13g2_a21oi_1 _2286_ (.A1(_0200_),
    .A2(_0201_),
    .Y(_0209_),
    .B1(net423));
 sg13g2_a22oi_1 _2287_ (.Y(_0210_),
    .B1(_0208_),
    .B2(_0209_),
    .A2(_0207_),
    .A1(net423));
 sg13g2_nand2_1 _2288_ (.Y(_0211_),
    .A(net448),
    .B(_0210_));
 sg13g2_nand2_1 _2289_ (.Y(_0212_),
    .A(\pqn_inst.v[6] ),
    .B(_0770_));
 sg13g2_a21o_1 _2290_ (.A2(_0212_),
    .A1(_0196_),
    .B1(_0204_),
    .X(_0213_));
 sg13g2_nand3_1 _2291_ (.B(_0204_),
    .C(_0212_),
    .A(_0196_),
    .Y(_0214_));
 sg13g2_nand3_1 _2292_ (.B(_0213_),
    .C(_0214_),
    .A(net452),
    .Y(_0215_));
 sg13g2_and2_1 _2293_ (.A(_1288_),
    .B(_0215_),
    .X(_0216_));
 sg13g2_a221oi_1 _2294_ (.B2(_0216_),
    .C1(net516),
    .B1(_0211_),
    .A1(_0731_),
    .Y(_0109_),
    .A2(net415));
 sg13g2_nor2_1 _2295_ (.A(_0730_),
    .B(_0768_),
    .Y(_0217_));
 sg13g2_xnor2_1 _2296_ (.Y(_0218_),
    .A(\pqn_inst.v[8] ),
    .B(\pqn_inst.multi.result[8] ));
 sg13g2_a21oi_2 _2297_ (.B1(_0218_),
    .Y(_0219_),
    .A2(_0205_),
    .A1(_0202_));
 sg13g2_nand3_1 _2298_ (.B(_0205_),
    .C(_0218_),
    .A(_0202_),
    .Y(_0220_));
 sg13g2_nand2_1 _2299_ (.Y(_0221_),
    .A(net422),
    .B(_0220_));
 sg13g2_xor2_1 _2300_ (.B(net522),
    .A(\pqn_inst.v[8] ),
    .X(_0222_));
 sg13g2_nand2b_1 _2301_ (.Y(_0223_),
    .B(_0200_),
    .A_N(_0186_));
 sg13g2_nor4_1 _2302_ (.A(_1331_),
    .B(_1346_),
    .C(_1359_),
    .D(_0223_),
    .Y(_0224_));
 sg13g2_a21oi_1 _2303_ (.A1(_0731_),
    .A2(_0732_),
    .Y(_0225_),
    .B1(net523));
 sg13g2_nor3_1 _2304_ (.A(_0187_),
    .B(_0224_),
    .C(_0225_),
    .Y(_0226_));
 sg13g2_or2_1 _2305_ (.X(_0227_),
    .B(_0226_),
    .A(_0222_));
 sg13g2_a21oi_1 _2306_ (.A1(_0222_),
    .A2(_0226_),
    .Y(_0228_),
    .B1(net422));
 sg13g2_a21oi_1 _2307_ (.A1(_0227_),
    .A2(_0228_),
    .Y(_0229_),
    .B1(net450));
 sg13g2_o21ai_1 _2308_ (.B1(_0229_),
    .Y(_0230_),
    .A1(_0219_),
    .A2(_0221_));
 sg13g2_o21ai_1 _2309_ (.B1(_0213_),
    .Y(_0231_),
    .A1(_0731_),
    .A2(\pqn_inst.multi.result[7] ));
 sg13g2_xnor2_1 _2310_ (.Y(_0232_),
    .A(_0218_),
    .B(_0231_));
 sg13g2_a21oi_1 _2311_ (.A1(net450),
    .A2(_0232_),
    .Y(_0233_),
    .B1(net413));
 sg13g2_a22oi_1 _2312_ (.Y(_0234_),
    .B1(_0230_),
    .B2(_0233_),
    .A2(net413),
    .A1(net229));
 sg13g2_nor2_1 _2313_ (.A(net514),
    .B(_0234_),
    .Y(_0110_));
 sg13g2_nand2_1 _2314_ (.Y(_0235_),
    .A(_0729_),
    .B(_0767_));
 sg13g2_nand2_1 _2315_ (.Y(_0236_),
    .A(\pqn_inst.v[9] ),
    .B(\pqn_inst.multi.result[9] ));
 sg13g2_nand2_1 _2316_ (.Y(_0237_),
    .A(_0235_),
    .B(_0236_));
 sg13g2_nor2_1 _2317_ (.A(_0217_),
    .B(_0219_),
    .Y(_0238_));
 sg13g2_xnor2_1 _2318_ (.Y(_0239_),
    .A(\pqn_inst.v[9] ),
    .B(net522));
 sg13g2_o21ai_1 _2319_ (.B1(_0227_),
    .Y(_0240_),
    .A1(_0730_),
    .A2(net522));
 sg13g2_xnor2_1 _2320_ (.Y(_0241_),
    .A(_0237_),
    .B(_0238_));
 sg13g2_o21ai_1 _2321_ (.B1(net424),
    .Y(_0242_),
    .A1(_0239_),
    .A2(_0240_));
 sg13g2_a21o_1 _2322_ (.A2(_0240_),
    .A1(_0239_),
    .B1(_0242_),
    .X(_0243_));
 sg13g2_o21ai_1 _2323_ (.B1(_0243_),
    .Y(_0244_),
    .A1(net424),
    .A2(_0241_));
 sg13g2_nor2_1 _2324_ (.A(_0730_),
    .B(\pqn_inst.multi.result[8] ),
    .Y(_0245_));
 sg13g2_a21oi_1 _2325_ (.A1(_0218_),
    .A2(_0231_),
    .Y(_0246_),
    .B1(_0245_));
 sg13g2_xnor2_1 _2326_ (.Y(_0247_),
    .A(_0237_),
    .B(_0246_));
 sg13g2_nand2_1 _2327_ (.Y(_0248_),
    .A(net450),
    .B(_0247_));
 sg13g2_a21oi_1 _2328_ (.A1(net448),
    .A2(_0244_),
    .Y(_0249_),
    .B1(net413));
 sg13g2_a221oi_1 _2329_ (.B2(_0249_),
    .C1(net514),
    .B1(_0248_),
    .A1(_0729_),
    .Y(_0111_),
    .A2(net413));
 sg13g2_nand2_1 _2330_ (.Y(_0250_),
    .A(\pqn_inst.v[10] ),
    .B(net505));
 sg13g2_xnor2_1 _2331_ (.Y(_0251_),
    .A(\pqn_inst.v[10] ),
    .B(net505));
 sg13g2_o21ai_1 _2332_ (.B1(_0235_),
    .Y(_0252_),
    .A1(_0217_),
    .A2(_0219_));
 sg13g2_nand3_1 _2333_ (.B(_0251_),
    .C(_0252_),
    .A(_0236_),
    .Y(_0253_));
 sg13g2_a21o_1 _2334_ (.A2(_0252_),
    .A1(_0236_),
    .B1(_0251_),
    .X(_0254_));
 sg13g2_and2_1 _2335_ (.A(net422),
    .B(_0253_),
    .X(_0255_));
 sg13g2_xor2_1 _2336_ (.B(net521),
    .A(\pqn_inst.v[10] ),
    .X(_0256_));
 sg13g2_nand2b_1 _2337_ (.Y(_0257_),
    .B(_0239_),
    .A_N(_0227_));
 sg13g2_o21ai_1 _2338_ (.B1(net519),
    .Y(_0258_),
    .A1(\pqn_inst.v[9] ),
    .A2(\pqn_inst.v[8] ));
 sg13g2_a21o_1 _2339_ (.A2(_0258_),
    .A1(_0257_),
    .B1(_0256_),
    .X(_0259_));
 sg13g2_nand3_1 _2340_ (.B(_0257_),
    .C(_0258_),
    .A(_0256_),
    .Y(_0260_));
 sg13g2_nand3_1 _2341_ (.B(_0259_),
    .C(_0260_),
    .A(net424),
    .Y(_0261_));
 sg13g2_nand2_1 _2342_ (.Y(_0262_),
    .A(net448),
    .B(_0261_));
 sg13g2_a21o_1 _2343_ (.A2(_0255_),
    .A1(_0254_),
    .B1(_0262_),
    .X(_0263_));
 sg13g2_nor2_1 _2344_ (.A(\pqn_inst.v[9] ),
    .B(net464),
    .Y(_0264_));
 sg13g2_nand2_1 _2345_ (.Y(_0265_),
    .A(\pqn_inst.v[9] ),
    .B(net464));
 sg13g2_o21ai_1 _2346_ (.B1(_0265_),
    .Y(_0266_),
    .A1(_0246_),
    .A2(_0264_));
 sg13g2_xnor2_1 _2347_ (.Y(_0267_),
    .A(_0251_),
    .B(_0266_));
 sg13g2_a21oi_1 _2348_ (.A1(net449),
    .A2(_0267_),
    .Y(_0268_),
    .B1(net412));
 sg13g2_a22oi_1 _2349_ (.Y(_0269_),
    .B1(_0263_),
    .B2(_0268_),
    .A2(net413),
    .A1(net238));
 sg13g2_nor2_1 _2350_ (.A(net512),
    .B(_0269_),
    .Y(_0112_));
 sg13g2_nor2_1 _2351_ (.A(\pqn_inst.v[11] ),
    .B(\pqn_inst.multi.result[11] ),
    .Y(_0270_));
 sg13g2_nand2_1 _2352_ (.Y(_0271_),
    .A(\pqn_inst.v[11] ),
    .B(\pqn_inst.multi.result[11] ));
 sg13g2_nor2b_1 _2353_ (.A(_0270_),
    .B_N(_0271_),
    .Y(_0272_));
 sg13g2_inv_1 _2354_ (.Y(_0273_),
    .A(_0272_));
 sg13g2_nand2_1 _2355_ (.Y(_0274_),
    .A(_0250_),
    .B(_0254_));
 sg13g2_xnor2_1 _2356_ (.Y(_0275_),
    .A(_0273_),
    .B(_0274_));
 sg13g2_xor2_1 _2357_ (.B(net520),
    .A(\pqn_inst.v[11] ),
    .X(_0276_));
 sg13g2_o21ai_1 _2358_ (.B1(_0259_),
    .Y(_0277_),
    .A1(_0728_),
    .A2(net521));
 sg13g2_xor2_1 _2359_ (.B(_0277_),
    .A(_0276_),
    .X(_0278_));
 sg13g2_o21ai_1 _2360_ (.B1(net448),
    .Y(_0279_),
    .A1(net421),
    .A2(_0278_));
 sg13g2_a21oi_1 _2361_ (.A1(net421),
    .A2(_0275_),
    .Y(_0280_),
    .B1(_0279_));
 sg13g2_nor2_1 _2362_ (.A(_0728_),
    .B(net505),
    .Y(_0281_));
 sg13g2_a21oi_2 _2363_ (.B1(_0281_),
    .Y(_0282_),
    .A2(_0266_),
    .A1(_0251_));
 sg13g2_and2_1 _2364_ (.A(_0273_),
    .B(_0282_),
    .X(_0283_));
 sg13g2_o21ai_1 _2365_ (.B1(net449),
    .Y(_0284_),
    .A1(_0273_),
    .A2(_0282_));
 sg13g2_o21ai_1 _2366_ (.B1(_1288_),
    .Y(_0285_),
    .A1(_0283_),
    .A2(_0284_));
 sg13g2_a21oi_1 _2367_ (.A1(net263),
    .A2(net412),
    .Y(_0286_),
    .B1(net512));
 sg13g2_o21ai_1 _2368_ (.B1(_0286_),
    .Y(_0113_),
    .A1(_0280_),
    .A2(_0285_));
 sg13g2_nand2_1 _2369_ (.Y(_0287_),
    .A(\pqn_inst.v[12] ),
    .B(net504));
 sg13g2_xnor2_1 _2370_ (.Y(_0288_),
    .A(\pqn_inst.v[12] ),
    .B(net504));
 sg13g2_a21o_1 _2371_ (.A2(_0254_),
    .A1(_0250_),
    .B1(_0270_),
    .X(_0289_));
 sg13g2_a21o_1 _2372_ (.A2(_0289_),
    .A1(_0271_),
    .B1(_0288_),
    .X(_0290_));
 sg13g2_nand3_1 _2373_ (.B(_0288_),
    .C(_0289_),
    .A(_0271_),
    .Y(_0291_));
 sg13g2_nand3_1 _2374_ (.B(_0290_),
    .C(_0291_),
    .A(net421),
    .Y(_0292_));
 sg13g2_xor2_1 _2375_ (.B(net520),
    .A(\pqn_inst.v[12] ),
    .X(_0293_));
 sg13g2_nor3_1 _2376_ (.A(_0256_),
    .B(_0257_),
    .C(_0276_),
    .Y(_0294_));
 sg13g2_o21ai_1 _2377_ (.B1(net519),
    .Y(_0295_),
    .A1(\pqn_inst.v[11] ),
    .A2(\pqn_inst.v[10] ));
 sg13g2_nand2_1 _2378_ (.Y(_0296_),
    .A(_0258_),
    .B(_0295_));
 sg13g2_nor2_1 _2379_ (.A(_0294_),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_or2_1 _2380_ (.X(_0298_),
    .B(_0297_),
    .A(_0293_));
 sg13g2_a21oi_1 _2381_ (.A1(_0293_),
    .A2(_0297_),
    .Y(_0299_),
    .B1(net421));
 sg13g2_a21oi_1 _2382_ (.A1(_0298_),
    .A2(_0299_),
    .Y(_0300_),
    .B1(net449));
 sg13g2_nor2_1 _2383_ (.A(\pqn_inst.v[11] ),
    .B(_0766_),
    .Y(_0301_));
 sg13g2_nand2_1 _2384_ (.Y(_0302_),
    .A(\pqn_inst.v[11] ),
    .B(_0766_));
 sg13g2_o21ai_1 _2385_ (.B1(_0302_),
    .Y(_0303_),
    .A1(_0282_),
    .A2(_0301_));
 sg13g2_xnor2_1 _2386_ (.Y(_0304_),
    .A(_0288_),
    .B(_0303_));
 sg13g2_a221oi_1 _2387_ (.B2(net449),
    .C1(net412),
    .B1(_0304_),
    .A1(_0292_),
    .Y(_0305_),
    .A2(_0300_));
 sg13g2_nor2_1 _2388_ (.A(net512),
    .B(_0305_),
    .Y(_0306_));
 sg13g2_o21ai_1 _2389_ (.B1(_0306_),
    .Y(_0114_),
    .A1(_0726_),
    .A2(_1288_));
 sg13g2_nor2_1 _2390_ (.A(net490),
    .B(\pqn_inst.multi.result[13] ),
    .Y(_0307_));
 sg13g2_nand2_1 _2391_ (.Y(_0308_),
    .A(net490),
    .B(\pqn_inst.multi.result[13] ));
 sg13g2_nand2b_1 _2392_ (.Y(_0309_),
    .B(_0308_),
    .A_N(_0307_));
 sg13g2_nand2_1 _2393_ (.Y(_0310_),
    .A(_0287_),
    .B(_0290_));
 sg13g2_xor2_1 _2394_ (.B(_0310_),
    .A(_0309_),
    .X(_0311_));
 sg13g2_o21ai_1 _2395_ (.B1(_0298_),
    .Y(_0312_),
    .A1(_0726_),
    .A2(net520));
 sg13g2_nand2b_1 _2396_ (.Y(_0313_),
    .B(net520),
    .A_N(net490));
 sg13g2_nor2b_1 _2397_ (.A(net520),
    .B_N(\pqn_inst.v[13] ),
    .Y(_0314_));
 sg13g2_xor2_1 _2398_ (.B(net520),
    .A(net490),
    .X(_0315_));
 sg13g2_xnor2_1 _2399_ (.Y(_0316_),
    .A(_0312_),
    .B(_0315_));
 sg13g2_a21oi_1 _2400_ (.A1(net424),
    .A2(_0316_),
    .Y(_0317_),
    .B1(net449));
 sg13g2_o21ai_1 _2401_ (.B1(_0317_),
    .Y(_0318_),
    .A1(net424),
    .A2(_0311_));
 sg13g2_nor2_1 _2402_ (.A(_0726_),
    .B(net504),
    .Y(_0319_));
 sg13g2_a21oi_2 _2403_ (.B1(_0319_),
    .Y(_0320_),
    .A2(_0303_),
    .A1(_0288_));
 sg13g2_a21oi_1 _2404_ (.A1(_0309_),
    .A2(_0320_),
    .Y(_0321_),
    .B1(net448));
 sg13g2_o21ai_1 _2405_ (.B1(_0321_),
    .Y(_0322_),
    .A1(_0309_),
    .A2(_0320_));
 sg13g2_nand3_1 _2406_ (.B(_0318_),
    .C(_0322_),
    .A(_1288_),
    .Y(_0323_));
 sg13g2_a21oi_1 _2407_ (.A1(net490),
    .A2(net412),
    .Y(_0324_),
    .B1(net512));
 sg13g2_nand2_1 _2408_ (.Y(_0115_),
    .A(_0323_),
    .B(_0324_));
 sg13g2_nand2_1 _2409_ (.Y(_0325_),
    .A(\pqn_inst.v[14] ),
    .B(\pqn_inst.multi.result[14] ));
 sg13g2_xnor2_1 _2410_ (.Y(_0326_),
    .A(\pqn_inst.v[14] ),
    .B(net503));
 sg13g2_a21o_1 _2411_ (.A2(_0290_),
    .A1(_0287_),
    .B1(_0307_),
    .X(_0327_));
 sg13g2_a21o_1 _2412_ (.A2(_0327_),
    .A1(_0308_),
    .B1(_0326_),
    .X(_0328_));
 sg13g2_nand3_1 _2413_ (.B(_0326_),
    .C(_0327_),
    .A(_0308_),
    .Y(_0329_));
 sg13g2_nand3_1 _2414_ (.B(_0328_),
    .C(_0329_),
    .A(net421),
    .Y(_0330_));
 sg13g2_xor2_1 _2415_ (.B(net520),
    .A(\pqn_inst.v[14] ),
    .X(_0331_));
 sg13g2_a21oi_1 _2416_ (.A1(_0312_),
    .A2(_0313_),
    .Y(_0332_),
    .B1(_0314_));
 sg13g2_nor2_1 _2417_ (.A(_0331_),
    .B(_0332_),
    .Y(_0333_));
 sg13g2_nand2_1 _2418_ (.Y(_0334_),
    .A(_0331_),
    .B(_0332_));
 sg13g2_nor2_1 _2419_ (.A(net421),
    .B(_0333_),
    .Y(_0335_));
 sg13g2_a21oi_1 _2420_ (.A1(_0334_),
    .A2(_0335_),
    .Y(_0336_),
    .B1(net449));
 sg13g2_nor2_1 _2421_ (.A(net490),
    .B(_0765_),
    .Y(_0337_));
 sg13g2_nand2_1 _2422_ (.Y(_0338_),
    .A(net490),
    .B(_0765_));
 sg13g2_o21ai_1 _2423_ (.B1(_0338_),
    .Y(_0339_),
    .A1(_0320_),
    .A2(_0337_));
 sg13g2_xnor2_1 _2424_ (.Y(_0340_),
    .A(_0326_),
    .B(_0339_));
 sg13g2_a221oi_1 _2425_ (.B2(net449),
    .C1(net412),
    .B1(_0340_),
    .A1(_0330_),
    .Y(_0341_),
    .A2(_0336_));
 sg13g2_a21oi_1 _2426_ (.A1(net264),
    .A2(net412),
    .Y(_0342_),
    .B1(net512));
 sg13g2_nand2b_1 _2427_ (.Y(_0116_),
    .B(_0342_),
    .A_N(_0341_));
 sg13g2_xor2_1 _2428_ (.B(\pqn_inst.multi.result[15] ),
    .A(\pqn_inst.v[15] ),
    .X(_0343_));
 sg13g2_a21o_1 _2429_ (.A2(_0328_),
    .A1(_0325_),
    .B1(_0343_),
    .X(_0344_));
 sg13g2_nand3_1 _2430_ (.B(_0328_),
    .C(_0343_),
    .A(_0325_),
    .Y(_0345_));
 sg13g2_nand3_1 _2431_ (.B(_0344_),
    .C(_0345_),
    .A(net421),
    .Y(_0346_));
 sg13g2_a21oi_1 _2432_ (.A1(\pqn_inst.v[14] ),
    .A2(net519),
    .Y(_0347_),
    .B1(_0333_));
 sg13g2_xnor2_1 _2433_ (.Y(_0348_),
    .A(\pqn_inst.v[15] ),
    .B(net520));
 sg13g2_or2_1 _2434_ (.X(_0349_),
    .B(_0348_),
    .A(_0347_));
 sg13g2_a21oi_1 _2435_ (.A1(_0347_),
    .A2(_0348_),
    .Y(_0350_),
    .B1(net421));
 sg13g2_a21oi_1 _2436_ (.A1(_0349_),
    .A2(_0350_),
    .Y(_0351_),
    .B1(net449));
 sg13g2_nor2b_1 _2437_ (.A(net503),
    .B_N(\pqn_inst.v[14] ),
    .Y(_0352_));
 sg13g2_a21oi_1 _2438_ (.A1(_0326_),
    .A2(_0339_),
    .Y(_0353_),
    .B1(_0352_));
 sg13g2_or2_1 _2439_ (.X(_0354_),
    .B(_0353_),
    .A(_0343_));
 sg13g2_a21oi_1 _2440_ (.A1(_0343_),
    .A2(_0353_),
    .Y(_0355_),
    .B1(net448));
 sg13g2_a22oi_1 _2441_ (.Y(_0356_),
    .B1(_0354_),
    .B2(_0355_),
    .A2(_0351_),
    .A1(_0346_));
 sg13g2_a21oi_1 _2442_ (.A1(net230),
    .A2(net412),
    .Y(_0357_),
    .B1(net513));
 sg13g2_o21ai_1 _2443_ (.B1(_0357_),
    .Y(_0117_),
    .A1(net412),
    .A2(_0356_));
 sg13g2_nand2b_1 _2444_ (.Y(_0358_),
    .B(net432),
    .A_N(_0003_));
 sg13g2_a21oi_1 _2445_ (.A1(_0778_),
    .A2(_1198_),
    .Y(_0359_),
    .B1(net419));
 sg13g2_a221oi_1 _2446_ (.B2(_0359_),
    .C1(net517),
    .B1(_0358_),
    .A1(_0751_),
    .Y(_0118_),
    .A2(net418));
 sg13g2_a21oi_1 _2447_ (.A1(uio_out[7]),
    .A2(_0778_),
    .Y(_0360_),
    .B1(_1199_));
 sg13g2_nor2_1 _2448_ (.A(_1287_),
    .B(_0360_),
    .Y(_0361_));
 sg13g2_nand3_1 _2449_ (.B(_1211_),
    .C(_0361_),
    .A(_1192_),
    .Y(_0362_));
 sg13g2_a21oi_1 _2450_ (.A1(net175),
    .A2(net418),
    .Y(_0363_),
    .B1(net517));
 sg13g2_o21ai_1 _2451_ (.B1(_0363_),
    .Y(_0119_),
    .A1(net418),
    .A2(_0362_));
 sg13g2_o21ai_1 _2452_ (.B1(_1199_),
    .Y(_0364_),
    .A1(net523),
    .A2(_1194_));
 sg13g2_nor2_1 _2453_ (.A(net431),
    .B(_0360_),
    .Y(_0365_));
 sg13g2_o21ai_1 _2454_ (.B1(_1177_),
    .Y(_0366_),
    .A1(_0006_),
    .A2(net426));
 sg13g2_a21oi_1 _2455_ (.A1(_0364_),
    .A2(_0365_),
    .Y(_0367_),
    .B1(_0366_));
 sg13g2_o21ai_1 _2456_ (.B1(net529),
    .Y(_0368_),
    .A1(net191),
    .A2(_1177_));
 sg13g2_nor2_1 _2457_ (.A(_0367_),
    .B(_0368_),
    .Y(_0120_));
 sg13g2_o21ai_1 _2458_ (.B1(_0365_),
    .Y(_0369_),
    .A1(net523),
    .A2(_1192_));
 sg13g2_a21oi_1 _2459_ (.A1(_0007_),
    .A2(net431),
    .Y(_0370_),
    .B1(net419));
 sg13g2_a22oi_1 _2460_ (.Y(_0371_),
    .B1(_0369_),
    .B2(_0370_),
    .A2(net419),
    .A1(net168));
 sg13g2_nor2_1 _2461_ (.A(net517),
    .B(net169),
    .Y(_0121_));
 sg13g2_and4_1 _2462_ (.A(uio_out[7]),
    .B(uio_out[6]),
    .C(uio_out[5]),
    .D(uio_out[4]),
    .X(_0372_));
 sg13g2_nor2b_1 _2463_ (.A(_0051_),
    .B_N(uio_out[2]),
    .Y(_0373_));
 sg13g2_o21ai_1 _2464_ (.B1(_0372_),
    .Y(_0374_),
    .A1(uio_out[3]),
    .A2(_0373_));
 sg13g2_nor4_1 _2465_ (.A(uo_out[7]),
    .B(uo_out[6]),
    .C(uo_out[5]),
    .D(uo_out[4]),
    .Y(_0375_));
 sg13g2_nand3b_1 _2466_ (.B(uio_out[2]),
    .C(uio_out[1]),
    .Y(_0376_),
    .A_N(uio_out[3]));
 sg13g2_nor2_1 _2467_ (.A(uio_out[0]),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_nor4_1 _2468_ (.A(uo_out[3]),
    .B(uo_out[2]),
    .C(uo_out[1]),
    .D(uo_out[0]),
    .Y(_0378_));
 sg13g2_xor2_1 _2469_ (.B(_0374_),
    .A(_0050_),
    .X(_0379_));
 sg13g2_nand4_1 _2470_ (.B(_0375_),
    .C(_0377_),
    .A(_0372_),
    .Y(_0380_),
    .D(_0378_));
 sg13g2_and2_2 _2471_ (.A(_0379_),
    .B(_0380_),
    .X(_0381_));
 sg13g2_nand2_1 _2472_ (.Y(_0382_),
    .A(_0379_),
    .B(_0380_));
 sg13g2_a21oi_1 _2473_ (.A1(_0379_),
    .A2(_0380_),
    .Y(_0383_),
    .B1(net523));
 sg13g2_nor2_1 _2474_ (.A(net522),
    .B(_1189_),
    .Y(_0384_));
 sg13g2_nor2_1 _2475_ (.A(_1172_),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_nor2_1 _2476_ (.A(net411),
    .B(_0385_),
    .Y(_0386_));
 sg13g2_nand2_1 _2477_ (.Y(_0387_),
    .A(uio_out[7]),
    .B(_1198_));
 sg13g2_o21ai_1 _2478_ (.B1(_0387_),
    .Y(_0388_),
    .A1(_0364_),
    .A2(_0386_));
 sg13g2_and2_1 _2479_ (.A(uo_out[4]),
    .B(net431),
    .X(_0389_));
 sg13g2_nor3_1 _2480_ (.A(net418),
    .B(_1181_),
    .C(_0389_),
    .Y(_0390_));
 sg13g2_a221oi_1 _2481_ (.B2(_0390_),
    .C1(net517),
    .B1(_0388_),
    .A1(_0747_),
    .Y(_0122_),
    .A2(net419));
 sg13g2_nor2_1 _2482_ (.A(_1193_),
    .B(_0382_),
    .Y(_0391_));
 sg13g2_nand2_1 _2483_ (.Y(_0392_),
    .A(net523),
    .B(_1195_));
 sg13g2_and3_1 _2484_ (.X(_0393_),
    .A(net523),
    .B(_0379_),
    .C(_0380_));
 sg13g2_nand3_1 _2485_ (.B(_0379_),
    .C(_0380_),
    .A(net523),
    .Y(_0394_));
 sg13g2_a21oi_1 _2486_ (.A1(_1172_),
    .A2(_0394_),
    .Y(_0395_),
    .B1(_1198_));
 sg13g2_o21ai_1 _2487_ (.B1(_0395_),
    .Y(_0396_),
    .A1(_0391_),
    .A2(_0392_));
 sg13g2_o21ai_1 _2488_ (.B1(_1177_),
    .Y(_0397_),
    .A1(_0008_),
    .A2(net426));
 sg13g2_a21oi_1 _2489_ (.A1(_0387_),
    .A2(_0396_),
    .Y(_0398_),
    .B1(_0397_));
 sg13g2_o21ai_1 _2490_ (.B1(net529),
    .Y(_0399_),
    .A1(net189),
    .A2(_1177_));
 sg13g2_nor2_1 _2491_ (.A(_0398_),
    .B(_0399_),
    .Y(_0123_));
 sg13g2_nand2_1 _2492_ (.Y(_0400_),
    .A(_1171_),
    .B(_0381_));
 sg13g2_a22oi_1 _2493_ (.Y(_0401_),
    .B1(_0400_),
    .B2(net446),
    .A2(_1198_),
    .A1(uio_out[7]));
 sg13g2_nand2_1 _2494_ (.Y(_0402_),
    .A(net133),
    .B(net418));
 sg13g2_a21oi_1 _2495_ (.A1(_0009_),
    .A2(net431),
    .Y(_0403_),
    .B1(net418));
 sg13g2_o21ai_1 _2496_ (.B1(_0403_),
    .Y(_0404_),
    .A1(_0384_),
    .A2(_0401_));
 sg13g2_a21oi_1 _2497_ (.A1(_0402_),
    .A2(_0404_),
    .Y(_0124_),
    .B1(net517));
 sg13g2_a21oi_1 _2498_ (.A1(_1172_),
    .A2(_0381_),
    .Y(_0405_),
    .B1(_0384_));
 sg13g2_nand2_1 _2499_ (.Y(_0406_),
    .A(_1199_),
    .B(_0405_));
 sg13g2_o21ai_1 _2500_ (.B1(_1177_),
    .Y(_0407_),
    .A1(_0010_),
    .A2(net426));
 sg13g2_a21oi_1 _2501_ (.A1(_0387_),
    .A2(_0406_),
    .Y(_0408_),
    .B1(_0407_));
 sg13g2_o21ai_1 _2502_ (.B1(net527),
    .Y(_0409_),
    .A1(net197),
    .A2(_1177_));
 sg13g2_nor2_1 _2503_ (.A(_0408_),
    .B(_0409_),
    .Y(_0125_));
 sg13g2_nand3_1 _2504_ (.B(net522),
    .C(_1171_),
    .A(net481),
    .Y(_0410_));
 sg13g2_nand2b_1 _2505_ (.Y(_0411_),
    .B(_0410_),
    .A_N(_0401_));
 sg13g2_a21oi_1 _2506_ (.A1(_0011_),
    .A2(net430),
    .Y(_0412_),
    .B1(net418));
 sg13g2_a22oi_1 _2507_ (.Y(_0413_),
    .B1(_0411_),
    .B2(_0412_),
    .A2(net418),
    .A1(net183));
 sg13g2_nor2_1 _2508_ (.A(net511),
    .B(net184),
    .Y(_0126_));
 sg13g2_nand2_1 _2509_ (.Y(_0414_),
    .A(_0051_),
    .B(net430));
 sg13g2_and2_2 _2510_ (.A(_1177_),
    .B(_0401_),
    .X(_0415_));
 sg13g2_a22oi_1 _2511_ (.Y(_0416_),
    .B1(_0414_),
    .B2(_0415_),
    .A2(net420),
    .A1(net144));
 sg13g2_nor2_1 _2512_ (.A(net511),
    .B(net145),
    .Y(_0127_));
 sg13g2_nand2_1 _2513_ (.Y(_0417_),
    .A(_0012_),
    .B(net428));
 sg13g2_a22oi_1 _2514_ (.Y(_0418_),
    .B1(_0415_),
    .B2(_0417_),
    .A2(net420),
    .A1(net140));
 sg13g2_nor2_1 _2515_ (.A(net509),
    .B(net141),
    .Y(_0128_));
 sg13g2_nand2_1 _2516_ (.Y(_0419_),
    .A(_0013_),
    .B(net428));
 sg13g2_a22oi_1 _2517_ (.Y(_0420_),
    .B1(_0415_),
    .B2(_0419_),
    .A2(net420),
    .A1(net142));
 sg13g2_nor2_1 _2518_ (.A(net509),
    .B(net143),
    .Y(_0129_));
 sg13g2_a22oi_1 _2519_ (.Y(_0421_),
    .B1(_1267_),
    .B2(_0415_),
    .A2(net420),
    .A1(net150));
 sg13g2_nor2_1 _2520_ (.A(net509),
    .B(net151),
    .Y(_0130_));
 sg13g2_a22oi_1 _2521_ (.Y(_0422_),
    .B1(_1272_),
    .B2(_0415_),
    .A2(net420),
    .A1(net154));
 sg13g2_nor2_1 _2522_ (.A(net509),
    .B(net155),
    .Y(_0131_));
 sg13g2_a22oi_1 _2523_ (.Y(_0423_),
    .B1(_1279_),
    .B2(_0415_),
    .A2(net420),
    .A1(net156));
 sg13g2_nor2_1 _2524_ (.A(net509),
    .B(net157),
    .Y(_0132_));
 sg13g2_a22oi_1 _2525_ (.Y(_0424_),
    .B1(_1283_),
    .B2(_0415_),
    .A2(net420),
    .A1(net187));
 sg13g2_nor2_1 _2526_ (.A(net509),
    .B(net188),
    .Y(_0133_));
 sg13g2_a21oi_1 _2527_ (.A1(_0764_),
    .A2(_0789_),
    .Y(_0134_),
    .B1(net491));
 sg13g2_o21ai_1 _2528_ (.B1(\pqn_inst.stage[3] ),
    .Y(_0425_),
    .A1(net463),
    .A2(_1167_));
 sg13g2_o21ai_1 _2529_ (.B1(_0425_),
    .Y(_0426_),
    .A1(net463),
    .A2(_1176_));
 sg13g2_nor2_2 _2530_ (.A(_0715_),
    .B(_0426_),
    .Y(_0427_));
 sg13g2_o21ai_1 _2531_ (.B1(net528),
    .Y(_0428_),
    .A1(net210),
    .A2(net405));
 sg13g2_a21oi_1 _2532_ (.A1(_0738_),
    .A2(net407),
    .Y(_0135_),
    .B1(_0428_));
 sg13g2_o21ai_1 _2533_ (.B1(net528),
    .Y(_0429_),
    .A1(net216),
    .A2(net405));
 sg13g2_a21oi_1 _2534_ (.A1(_0737_),
    .A2(net405),
    .Y(_0136_),
    .B1(_0429_));
 sg13g2_o21ai_1 _2535_ (.B1(net528),
    .Y(_0430_),
    .A1(net214),
    .A2(net405));
 sg13g2_a21oi_1 _2536_ (.A1(_0736_),
    .A2(net406),
    .Y(_0137_),
    .B1(_0430_));
 sg13g2_o21ai_1 _2537_ (.B1(net526),
    .Y(_0431_),
    .A1(net208),
    .A2(net405));
 sg13g2_a21oi_1 _2538_ (.A1(_0735_),
    .A2(net405),
    .Y(_0138_),
    .B1(_0431_));
 sg13g2_o21ai_1 _2539_ (.B1(net528),
    .Y(_0432_),
    .A1(uo_out[4]),
    .A2(net406));
 sg13g2_a21oi_1 _2540_ (.A1(_0734_),
    .A2(net406),
    .Y(_0139_),
    .B1(_0432_));
 sg13g2_o21ai_1 _2541_ (.B1(net527),
    .Y(_0433_),
    .A1(net240),
    .A2(net405));
 sg13g2_a21oi_1 _2542_ (.A1(_0733_),
    .A2(net405),
    .Y(_0140_),
    .B1(_0433_));
 sg13g2_o21ai_1 _2543_ (.B1(net528),
    .Y(_0434_),
    .A1(net245),
    .A2(net406));
 sg13g2_a21oi_1 _2544_ (.A1(_0732_),
    .A2(net406),
    .Y(_0141_),
    .B1(_0434_));
 sg13g2_o21ai_1 _2545_ (.B1(net527),
    .Y(_0435_),
    .A1(net247),
    .A2(net406));
 sg13g2_a21oi_1 _2546_ (.A1(_0731_),
    .A2(net406),
    .Y(_0142_),
    .B1(_0435_));
 sg13g2_o21ai_1 _2547_ (.B1(net527),
    .Y(_0436_),
    .A1(net242),
    .A2(net407));
 sg13g2_a21oi_1 _2548_ (.A1(_0730_),
    .A2(net407),
    .Y(_0143_),
    .B1(_0436_));
 sg13g2_o21ai_1 _2549_ (.B1(net526),
    .Y(_0437_),
    .A1(net243),
    .A2(net404));
 sg13g2_a21oi_1 _2550_ (.A1(_0729_),
    .A2(net404),
    .Y(_0144_),
    .B1(_0437_));
 sg13g2_o21ai_1 _2551_ (.B1(net526),
    .Y(_0438_),
    .A1(net258),
    .A2(net404));
 sg13g2_a21oi_1 _2552_ (.A1(_0728_),
    .A2(net404),
    .Y(_0145_),
    .B1(_0438_));
 sg13g2_a21oi_1 _2553_ (.A1(\pqn_inst.v[11] ),
    .A2(net404),
    .Y(_0439_),
    .B1(net512));
 sg13g2_o21ai_1 _2554_ (.B1(_0439_),
    .Y(_0146_),
    .A1(_0727_),
    .A2(net404));
 sg13g2_a21oi_1 _2555_ (.A1(\pqn_inst.v[12] ),
    .A2(net403),
    .Y(_0440_),
    .B1(net513));
 sg13g2_o21ai_1 _2556_ (.B1(_0440_),
    .Y(_0147_),
    .A1(_0725_),
    .A2(net403));
 sg13g2_a21oi_1 _2557_ (.A1(net490),
    .A2(net403),
    .Y(_0441_),
    .B1(net512));
 sg13g2_o21ai_1 _2558_ (.B1(_0441_),
    .Y(_0148_),
    .A1(_0724_),
    .A2(net403));
 sg13g2_a21oi_1 _2559_ (.A1(\pqn_inst.v[14] ),
    .A2(net403),
    .Y(_0442_),
    .B1(net512));
 sg13g2_o21ai_1 _2560_ (.B1(_0442_),
    .Y(_0149_),
    .A1(_0723_),
    .A2(net403));
 sg13g2_a21oi_1 _2561_ (.A1(net230),
    .A2(net403),
    .Y(_0443_),
    .B1(net513));
 sg13g2_o21ai_1 _2562_ (.B1(_0443_),
    .Y(_0150_),
    .A1(_0722_),
    .A2(net403));
 sg13g2_nand2b_1 _2563_ (.Y(_0444_),
    .B(_0383_),
    .A_N(_0049_));
 sg13g2_nand2b_1 _2564_ (.Y(_0445_),
    .B(_0049_),
    .A_N(net411));
 sg13g2_nand3_1 _2565_ (.B(_0444_),
    .C(_0445_),
    .A(net443),
    .Y(_0446_));
 sg13g2_nand2_1 _2566_ (.Y(_0447_),
    .A(\pqn_inst.n[2] ),
    .B(\pqn_inst.multi.result[2] ));
 sg13g2_xnor2_1 _2567_ (.Y(_0448_),
    .A(\pqn_inst.n[2] ),
    .B(\pqn_inst.multi.result[2] ));
 sg13g2_nor2_1 _2568_ (.A(\pqn_inst.n[1] ),
    .B(net507),
    .Y(_0449_));
 sg13g2_a22oi_1 _2569_ (.Y(_0450_),
    .B1(\pqn_inst.multi.result[0] ),
    .B2(\pqn_inst.n[0] ),
    .A2(net507),
    .A1(\pqn_inst.n[1] ));
 sg13g2_or3_1 _2570_ (.A(_0448_),
    .B(_0449_),
    .C(_0450_),
    .X(_0451_));
 sg13g2_o21ai_1 _2571_ (.B1(_0448_),
    .Y(_0452_),
    .A1(_0449_),
    .A2(_0450_));
 sg13g2_nand3_1 _2572_ (.B(_0451_),
    .C(_0452_),
    .A(net444),
    .Y(_0453_));
 sg13g2_nand3_1 _2573_ (.B(_1176_),
    .C(net408),
    .A(_1173_),
    .Y(_0454_));
 sg13g2_nand4_1 _2574_ (.B(_1189_),
    .C(_1199_),
    .A(_0816_),
    .Y(_0455_),
    .D(_0454_));
 sg13g2_nor2_2 _2575_ (.A(_1172_),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_nand2b_2 _2576_ (.Y(_0457_),
    .B(_1173_),
    .A_N(_0455_));
 sg13g2_xor2_1 _2577_ (.B(net507),
    .A(\pqn_inst.n[1] ),
    .X(_0458_));
 sg13g2_nor2b_1 _2578_ (.A(\pqn_inst.n[0] ),
    .B_N(\pqn_inst.multi.result[0] ),
    .Y(_0459_));
 sg13g2_nand2b_1 _2579_ (.Y(_0460_),
    .B(\pqn_inst.n[1] ),
    .A_N(net507));
 sg13g2_o21ai_1 _2580_ (.B1(_0460_),
    .Y(_0461_),
    .A1(_0458_),
    .A2(_0459_));
 sg13g2_xor2_1 _2581_ (.B(_0461_),
    .A(_0448_),
    .X(_0462_));
 sg13g2_a21o_1 _2582_ (.A2(_0453_),
    .A1(_0446_),
    .B1(net433),
    .X(_0463_));
 sg13g2_a21oi_1 _2583_ (.A1(net433),
    .A2(_0462_),
    .Y(_0464_),
    .B1(_0457_));
 sg13g2_a221oi_1 _2584_ (.B2(_0464_),
    .C1(net515),
    .B1(_0463_),
    .A1(_0721_),
    .Y(_0151_),
    .A2(net400));
 sg13g2_nand2b_2 _2585_ (.Y(_0465_),
    .B(_0394_),
    .A_N(net411));
 sg13g2_nand2_1 _2586_ (.Y(_0466_),
    .A(_0444_),
    .B(_0465_));
 sg13g2_or2_1 _2587_ (.X(_0467_),
    .B(_0466_),
    .A(_0052_));
 sg13g2_a21oi_1 _2588_ (.A1(_0052_),
    .A2(_0466_),
    .Y(_0468_),
    .B1(net444));
 sg13g2_and2_1 _2589_ (.A(\pqn_inst.n[3] ),
    .B(\pqn_inst.multi.result[3] ),
    .X(_0469_));
 sg13g2_xnor2_1 _2590_ (.Y(_0470_),
    .A(\pqn_inst.n[3] ),
    .B(\pqn_inst.multi.result[3] ));
 sg13g2_inv_1 _2591_ (.Y(_0471_),
    .A(_0470_));
 sg13g2_nand2_1 _2592_ (.Y(_0472_),
    .A(_0447_),
    .B(_0451_));
 sg13g2_a21oi_1 _2593_ (.A1(_0447_),
    .A2(_0451_),
    .Y(_0473_),
    .B1(_0470_));
 sg13g2_xnor2_1 _2594_ (.Y(_0474_),
    .A(_0471_),
    .B(_0472_));
 sg13g2_a221oi_1 _2595_ (.B2(net445),
    .C1(net432),
    .B1(_0474_),
    .A1(_0467_),
    .Y(_0475_),
    .A2(_0468_));
 sg13g2_nor2_1 _2596_ (.A(_0721_),
    .B(\pqn_inst.multi.result[2] ),
    .Y(_0476_));
 sg13g2_a21oi_2 _2597_ (.B1(_0476_),
    .Y(_0477_),
    .A2(_0461_),
    .A1(_0448_));
 sg13g2_a21oi_1 _2598_ (.A1(_0471_),
    .A2(_0477_),
    .Y(_0478_),
    .B1(net425));
 sg13g2_o21ai_1 _2599_ (.B1(_0478_),
    .Y(_0479_),
    .A1(_0471_),
    .A2(_0477_));
 sg13g2_nand3b_1 _2600_ (.B(_0479_),
    .C(_0456_),
    .Y(_0480_),
    .A_N(_0475_));
 sg13g2_o21ai_1 _2601_ (.B1(_0480_),
    .Y(_0481_),
    .A1(net249),
    .A2(_0456_));
 sg13g2_nor2_1 _2602_ (.A(net515),
    .B(_0481_),
    .Y(_0152_));
 sg13g2_or4_1 _2603_ (.A(net523),
    .B(_0049_),
    .C(_0052_),
    .D(_0381_),
    .X(_0482_));
 sg13g2_nand3b_1 _2604_ (.B(_0394_),
    .C(\pqn_inst.n[3] ),
    .Y(_0483_),
    .A_N(net411));
 sg13g2_o21ai_1 _2605_ (.B1(\pqn_inst.n[4] ),
    .Y(_0484_),
    .A1(net411),
    .A2(_0393_));
 sg13g2_or3_1 _2606_ (.A(\pqn_inst.n[4] ),
    .B(net411),
    .C(_0393_),
    .X(_0485_));
 sg13g2_a22oi_1 _2607_ (.Y(_0486_),
    .B1(_0484_),
    .B2(_0485_),
    .A2(_0483_),
    .A1(_0482_));
 sg13g2_nand4_1 _2608_ (.B(_0483_),
    .C(_0484_),
    .A(_0482_),
    .Y(_0487_),
    .D(_0485_));
 sg13g2_nor2b_1 _2609_ (.A(_0486_),
    .B_N(_0487_),
    .Y(_0488_));
 sg13g2_nand2_1 _2610_ (.Y(_0489_),
    .A(\pqn_inst.n[4] ),
    .B(net506));
 sg13g2_xor2_1 _2611_ (.B(net506),
    .A(\pqn_inst.n[4] ),
    .X(_0490_));
 sg13g2_xnor2_1 _2612_ (.Y(_0491_),
    .A(\pqn_inst.n[4] ),
    .B(net506));
 sg13g2_nor3_1 _2613_ (.A(_0469_),
    .B(_0473_),
    .C(_0490_),
    .Y(_0492_));
 sg13g2_o21ai_1 _2614_ (.B1(_0490_),
    .Y(_0493_),
    .A1(_0469_),
    .A2(_0473_));
 sg13g2_nor2_1 _2615_ (.A(net443),
    .B(_0492_),
    .Y(_0494_));
 sg13g2_a221oi_1 _2616_ (.B2(_0494_),
    .C1(net432),
    .B1(_0493_),
    .A1(net443),
    .Y(_0495_),
    .A2(_0488_));
 sg13g2_nand2_1 _2617_ (.Y(_0496_),
    .A(\pqn_inst.n[3] ),
    .B(_0772_));
 sg13g2_o21ai_1 _2618_ (.B1(_0496_),
    .Y(_0497_),
    .A1(_0471_),
    .A2(_0477_));
 sg13g2_xnor2_1 _2619_ (.Y(_0498_),
    .A(_0491_),
    .B(_0497_));
 sg13g2_a21oi_1 _2620_ (.A1(net432),
    .A2(_0498_),
    .Y(_0499_),
    .B1(_0495_));
 sg13g2_o21ai_1 _2621_ (.B1(net529),
    .Y(_0500_),
    .A1(net400),
    .A2(_0499_));
 sg13g2_a21oi_1 _2622_ (.A1(_0720_),
    .A2(net400),
    .Y(_0153_),
    .B1(_0500_));
 sg13g2_nand2_1 _2623_ (.Y(_0501_),
    .A(\pqn_inst.n[5] ),
    .B(_0778_));
 sg13g2_xnor2_1 _2624_ (.Y(_0502_),
    .A(\pqn_inst.n[5] ),
    .B(net524));
 sg13g2_nor2_1 _2625_ (.A(_0053_),
    .B(_0465_),
    .Y(_0503_));
 sg13g2_nor2_1 _2626_ (.A(_0486_),
    .B(_0503_),
    .Y(_0504_));
 sg13g2_o21ai_1 _2627_ (.B1(_0502_),
    .Y(_0505_),
    .A1(_0486_),
    .A2(_0503_));
 sg13g2_nor2_1 _2628_ (.A(_0719_),
    .B(_0771_),
    .Y(_0506_));
 sg13g2_xnor2_1 _2629_ (.Y(_0507_),
    .A(\pqn_inst.n[5] ),
    .B(\pqn_inst.multi.result[5] ));
 sg13g2_nand2_1 _2630_ (.Y(_0508_),
    .A(_0489_),
    .B(_0493_));
 sg13g2_xnor2_1 _2631_ (.Y(_0509_),
    .A(_0502_),
    .B(_0504_));
 sg13g2_xor2_1 _2632_ (.B(_0508_),
    .A(_0507_),
    .X(_0510_));
 sg13g2_a21oi_1 _2633_ (.A1(net444),
    .A2(_0510_),
    .Y(_0511_),
    .B1(net432));
 sg13g2_o21ai_1 _2634_ (.B1(_0511_),
    .Y(_0512_),
    .A1(net444),
    .A2(_0509_));
 sg13g2_nor2_1 _2635_ (.A(_0720_),
    .B(net506),
    .Y(_0513_));
 sg13g2_a21o_1 _2636_ (.A2(_0497_),
    .A1(_0491_),
    .B1(_0513_),
    .X(_0514_));
 sg13g2_xor2_1 _2637_ (.B(_0514_),
    .A(_0507_),
    .X(_0515_));
 sg13g2_a21oi_1 _2638_ (.A1(net432),
    .A2(_0515_),
    .Y(_0516_),
    .B1(net400));
 sg13g2_a221oi_1 _2639_ (.B2(_0516_),
    .C1(net517),
    .B1(_0512_),
    .A1(_0719_),
    .Y(_0154_),
    .A2(net400));
 sg13g2_nand2_1 _2640_ (.Y(_0517_),
    .A(\pqn_inst.n[6] ),
    .B(\pqn_inst.multi.result[6] ));
 sg13g2_xor2_1 _2641_ (.B(\pqn_inst.multi.result[6] ),
    .A(\pqn_inst.n[6] ),
    .X(_0518_));
 sg13g2_a22oi_1 _2642_ (.Y(_0519_),
    .B1(_0489_),
    .B2(_0493_),
    .A2(_0771_),
    .A1(_0719_));
 sg13g2_nor3_1 _2643_ (.A(_0506_),
    .B(_0518_),
    .C(_0519_),
    .Y(_0520_));
 sg13g2_o21ai_1 _2644_ (.B1(_0518_),
    .Y(_0521_),
    .A1(_0506_),
    .A2(_0519_));
 sg13g2_nor2_1 _2645_ (.A(net443),
    .B(_0520_),
    .Y(_0522_));
 sg13g2_xnor2_1 _2646_ (.Y(_0523_),
    .A(\pqn_inst.n[6] ),
    .B(_0465_));
 sg13g2_a21oi_2 _2647_ (.B1(_0523_),
    .Y(_0524_),
    .A2(_0505_),
    .A1(_0501_));
 sg13g2_and3_1 _2648_ (.X(_0525_),
    .A(_0501_),
    .B(_0505_),
    .C(_0523_));
 sg13g2_nor3_1 _2649_ (.A(net444),
    .B(_0524_),
    .C(_0525_),
    .Y(_0526_));
 sg13g2_a21o_1 _2650_ (.A2(_0522_),
    .A1(_0521_),
    .B1(_0526_),
    .X(_0527_));
 sg13g2_nor2_1 _2651_ (.A(\pqn_inst.n[5] ),
    .B(_0771_),
    .Y(_0528_));
 sg13g2_a221oi_1 _2652_ (.B2(_0497_),
    .C1(_0513_),
    .B1(_0491_),
    .A1(\pqn_inst.n[5] ),
    .Y(_0529_),
    .A2(_0771_));
 sg13g2_o21ai_1 _2653_ (.B1(_0518_),
    .Y(_0530_),
    .A1(_0528_),
    .A2(_0529_));
 sg13g2_nor3_2 _2654_ (.A(_0518_),
    .B(_0528_),
    .C(_0529_),
    .Y(_0531_));
 sg13g2_nor2_1 _2655_ (.A(net425),
    .B(_0531_),
    .Y(_0532_));
 sg13g2_a221oi_1 _2656_ (.B2(_0532_),
    .C1(net400),
    .B1(_0530_),
    .A1(net425),
    .Y(_0533_),
    .A2(_0527_));
 sg13g2_o21ai_1 _2657_ (.B1(net529),
    .Y(_0534_),
    .A1(net283),
    .A2(_0456_));
 sg13g2_nor2_1 _2658_ (.A(_0533_),
    .B(_0534_),
    .Y(_0155_));
 sg13g2_nand2b_2 _2659_ (.Y(_0535_),
    .B(_0393_),
    .A_N(\pqn_inst.n[7] ));
 sg13g2_nand2_1 _2660_ (.Y(_0536_),
    .A(\pqn_inst.n[7] ),
    .B(_0394_));
 sg13g2_nand2_1 _2661_ (.Y(_0537_),
    .A(_0535_),
    .B(_0536_));
 sg13g2_a21oi_1 _2662_ (.A1(\pqn_inst.n[6] ),
    .A2(_0465_),
    .Y(_0538_),
    .B1(_0524_));
 sg13g2_xnor2_1 _2663_ (.Y(_0539_),
    .A(_0537_),
    .B(_0538_));
 sg13g2_nand2_1 _2664_ (.Y(_0540_),
    .A(net443),
    .B(_0539_));
 sg13g2_and2_1 _2665_ (.A(\pqn_inst.n[7] ),
    .B(\pqn_inst.multi.result[7] ),
    .X(_0541_));
 sg13g2_xnor2_1 _2666_ (.Y(_0542_),
    .A(\pqn_inst.n[7] ),
    .B(\pqn_inst.multi.result[7] ));
 sg13g2_and3_1 _2667_ (.X(_0543_),
    .A(_0517_),
    .B(_0521_),
    .C(_0542_));
 sg13g2_a21oi_2 _2668_ (.B1(_0542_),
    .Y(_0544_),
    .A2(_0521_),
    .A1(_0517_));
 sg13g2_o21ai_1 _2669_ (.B1(net444),
    .Y(_0545_),
    .A1(_0543_),
    .A2(_0544_));
 sg13g2_nand3_1 _2670_ (.B(_0540_),
    .C(_0545_),
    .A(net425),
    .Y(_0546_));
 sg13g2_nor2b_1 _2671_ (.A(\pqn_inst.multi.result[6] ),
    .B_N(\pqn_inst.n[6] ),
    .Y(_0547_));
 sg13g2_nor3_1 _2672_ (.A(_0531_),
    .B(_0542_),
    .C(_0547_),
    .Y(_0548_));
 sg13g2_o21ai_1 _2673_ (.B1(_0542_),
    .Y(_0549_),
    .A1(_0531_),
    .A2(_0547_));
 sg13g2_nor2_1 _2674_ (.A(net425),
    .B(_0548_),
    .Y(_0550_));
 sg13g2_a21oi_1 _2675_ (.A1(_0549_),
    .A2(_0550_),
    .Y(_0551_),
    .B1(net400));
 sg13g2_o21ai_1 _2676_ (.B1(net529),
    .Y(_0552_),
    .A1(net257),
    .A2(_0456_));
 sg13g2_a21oi_1 _2677_ (.A1(_0546_),
    .A2(_0551_),
    .Y(_0156_),
    .B1(_0552_));
 sg13g2_nand2_1 _2678_ (.Y(_0553_),
    .A(\pqn_inst.n[8] ),
    .B(net411));
 sg13g2_xnor2_1 _2679_ (.Y(_0554_),
    .A(\pqn_inst.n[8] ),
    .B(net411));
 sg13g2_inv_1 _2680_ (.Y(_0555_),
    .A(_0554_));
 sg13g2_nand3_1 _2681_ (.B(_0465_),
    .C(_0535_),
    .A(\pqn_inst.n[6] ),
    .Y(_0556_));
 sg13g2_nand2_1 _2682_ (.Y(_0557_),
    .A(_0536_),
    .B(_0556_));
 sg13g2_o21ai_1 _2683_ (.B1(_0555_),
    .Y(_0558_),
    .A1(_0524_),
    .A2(_0557_));
 sg13g2_nor3_1 _2684_ (.A(_0524_),
    .B(_0555_),
    .C(_0557_),
    .Y(_0559_));
 sg13g2_nor2_1 _2685_ (.A(net444),
    .B(_0559_),
    .Y(_0560_));
 sg13g2_nand2_1 _2686_ (.Y(_0561_),
    .A(\pqn_inst.n[8] ),
    .B(\pqn_inst.multi.result[8] ));
 sg13g2_xnor2_1 _2687_ (.Y(_0562_),
    .A(\pqn_inst.n[8] ),
    .B(\pqn_inst.multi.result[8] ));
 sg13g2_inv_1 _2688_ (.Y(_0563_),
    .A(_0562_));
 sg13g2_o21ai_1 _2689_ (.B1(_0563_),
    .Y(_0564_),
    .A1(_0541_),
    .A2(_0544_));
 sg13g2_nor3_1 _2690_ (.A(_0541_),
    .B(_0544_),
    .C(_0563_),
    .Y(_0565_));
 sg13g2_nor2_1 _2691_ (.A(net442),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_a22oi_1 _2692_ (.Y(_0567_),
    .B1(_0564_),
    .B2(_0566_),
    .A2(_0560_),
    .A1(_0558_));
 sg13g2_nand2_1 _2693_ (.Y(_0568_),
    .A(\pqn_inst.n[7] ),
    .B(_0769_));
 sg13g2_a21oi_2 _2694_ (.B1(_0563_),
    .Y(_0569_),
    .A2(_0568_),
    .A1(_0549_));
 sg13g2_nand3_1 _2695_ (.B(_0563_),
    .C(_0568_),
    .A(_0549_),
    .Y(_0570_));
 sg13g2_nor2_1 _2696_ (.A(net426),
    .B(_0569_),
    .Y(_0571_));
 sg13g2_a21oi_1 _2697_ (.A1(_0570_),
    .A2(_0571_),
    .Y(_0572_),
    .B1(net400));
 sg13g2_o21ai_1 _2698_ (.B1(_0572_),
    .Y(_0573_),
    .A1(net431),
    .A2(_0567_));
 sg13g2_o21ai_1 _2699_ (.B1(_0573_),
    .Y(_0574_),
    .A1(net276),
    .A2(_0456_));
 sg13g2_nor2_1 _2700_ (.A(net517),
    .B(_0574_),
    .Y(_0157_));
 sg13g2_nor2_2 _2701_ (.A(net519),
    .B(_0381_),
    .Y(_0575_));
 sg13g2_nand2_2 _2702_ (.Y(_0576_),
    .A(net521),
    .B(_0382_));
 sg13g2_xnor2_1 _2703_ (.Y(_0577_),
    .A(\pqn_inst.n[9] ),
    .B(_0575_));
 sg13g2_nand2_1 _2704_ (.Y(_0578_),
    .A(_0553_),
    .B(_0558_));
 sg13g2_xor2_1 _2705_ (.B(_0578_),
    .A(_0577_),
    .X(_0579_));
 sg13g2_and2_1 _2706_ (.A(_0561_),
    .B(_0564_),
    .X(_0580_));
 sg13g2_nand2_1 _2707_ (.Y(_0581_),
    .A(_0718_),
    .B(net464));
 sg13g2_nand2_1 _2708_ (.Y(_0582_),
    .A(\pqn_inst.n[9] ),
    .B(\pqn_inst.multi.result[9] ));
 sg13g2_and2_1 _2709_ (.A(_0581_),
    .B(_0582_),
    .X(_0583_));
 sg13g2_o21ai_1 _2710_ (.B1(net445),
    .Y(_0584_),
    .A1(_0580_),
    .A2(_0583_));
 sg13g2_a21oi_1 _2711_ (.A1(_0580_),
    .A2(_0583_),
    .Y(_0585_),
    .B1(_0584_));
 sg13g2_nor2_1 _2712_ (.A(net430),
    .B(_0585_),
    .Y(_0586_));
 sg13g2_o21ai_1 _2713_ (.B1(_0586_),
    .Y(_0587_),
    .A1(net445),
    .A2(_0579_));
 sg13g2_a21oi_2 _2714_ (.B1(_0569_),
    .Y(_0588_),
    .A2(_0768_),
    .A1(\pqn_inst.n[8] ));
 sg13g2_o21ai_1 _2715_ (.B1(net430),
    .Y(_0589_),
    .A1(_0583_),
    .A2(_0588_));
 sg13g2_a21oi_1 _2716_ (.A1(_0583_),
    .A2(_0588_),
    .Y(_0590_),
    .B1(_0589_));
 sg13g2_nor2_1 _2717_ (.A(net399),
    .B(_0590_),
    .Y(_0591_));
 sg13g2_a221oi_1 _2718_ (.B2(_0591_),
    .C1(net511),
    .B1(_0587_),
    .A1(_0718_),
    .Y(_0158_),
    .A2(net399));
 sg13g2_nor2_1 _2719_ (.A(_0717_),
    .B(_0575_),
    .Y(_0592_));
 sg13g2_xnor2_1 _2720_ (.Y(_0593_),
    .A(\pqn_inst.n[10] ),
    .B(_0575_));
 sg13g2_nand2_1 _2721_ (.Y(_0594_),
    .A(_0535_),
    .B(_0577_));
 sg13g2_o21ai_1 _2722_ (.B1(_0553_),
    .Y(_0595_),
    .A1(_0718_),
    .A2(_0575_));
 sg13g2_inv_1 _2723_ (.Y(_0596_),
    .A(_0595_));
 sg13g2_o21ai_1 _2724_ (.B1(_0596_),
    .Y(_0597_),
    .A1(_0558_),
    .A2(_0594_));
 sg13g2_o21ai_1 _2725_ (.B1(net442),
    .Y(_0598_),
    .A1(_0593_),
    .A2(_0597_));
 sg13g2_a21o_1 _2726_ (.A2(_0597_),
    .A1(_0593_),
    .B1(_0598_),
    .X(_0599_));
 sg13g2_and2_1 _2727_ (.A(\pqn_inst.n[10] ),
    .B(\pqn_inst.multi.result[10] ),
    .X(_0600_));
 sg13g2_xor2_1 _2728_ (.B(\pqn_inst.multi.result[10] ),
    .A(\pqn_inst.n[10] ),
    .X(_0601_));
 sg13g2_xnor2_1 _2729_ (.Y(_0602_),
    .A(\pqn_inst.n[10] ),
    .B(\pqn_inst.multi.result[10] ));
 sg13g2_nand3_1 _2730_ (.B(_0564_),
    .C(_0582_),
    .A(_0561_),
    .Y(_0603_));
 sg13g2_a21o_1 _2731_ (.A2(_0603_),
    .A1(_0581_),
    .B1(_0601_),
    .X(_0604_));
 sg13g2_and3_1 _2732_ (.X(_0605_),
    .A(_0581_),
    .B(_0601_),
    .C(_0603_));
 sg13g2_nor2_1 _2733_ (.A(net442),
    .B(_0605_),
    .Y(_0606_));
 sg13g2_a21oi_1 _2734_ (.A1(_0604_),
    .A2(_0606_),
    .Y(_0607_),
    .B1(net428));
 sg13g2_nand2_1 _2735_ (.Y(_0608_),
    .A(\pqn_inst.n[9] ),
    .B(net464));
 sg13g2_nor2_1 _2736_ (.A(\pqn_inst.n[9] ),
    .B(net464),
    .Y(_0609_));
 sg13g2_a21oi_2 _2737_ (.B1(_0609_),
    .Y(_0610_),
    .A2(_0608_),
    .A1(_0588_));
 sg13g2_xnor2_1 _2738_ (.Y(_0611_),
    .A(_0602_),
    .B(_0610_));
 sg13g2_a221oi_1 _2739_ (.B2(net428),
    .C1(net399),
    .B1(_0611_),
    .A1(_0599_),
    .Y(_0612_),
    .A2(_0607_));
 sg13g2_a21oi_1 _2740_ (.A1(net261),
    .A2(net398),
    .Y(_0613_),
    .B1(net509));
 sg13g2_nand2b_1 _2741_ (.Y(_0159_),
    .B(_0613_),
    .A_N(_0612_));
 sg13g2_a21oi_1 _2742_ (.A1(_0593_),
    .A2(_0597_),
    .Y(_0614_),
    .B1(_0592_));
 sg13g2_nor2_1 _2743_ (.A(net484),
    .B(_0576_),
    .Y(_0615_));
 sg13g2_xnor2_1 _2744_ (.Y(_0616_),
    .A(\pqn_inst.n[11] ),
    .B(_0575_));
 sg13g2_xnor2_1 _2745_ (.Y(_0617_),
    .A(_0614_),
    .B(_0616_));
 sg13g2_or2_1 _2746_ (.X(_0618_),
    .B(\pqn_inst.multi.result[11] ),
    .A(net484));
 sg13g2_nand2_1 _2747_ (.Y(_0619_),
    .A(net484),
    .B(\pqn_inst.multi.result[11] ));
 sg13g2_nand2_1 _2748_ (.Y(_0620_),
    .A(_0618_),
    .B(_0619_));
 sg13g2_nor2_1 _2749_ (.A(_0600_),
    .B(_0605_),
    .Y(_0621_));
 sg13g2_xor2_1 _2750_ (.B(_0621_),
    .A(_0620_),
    .X(_0622_));
 sg13g2_mux2_1 _2751_ (.A0(_0617_),
    .A1(_0622_),
    .S(net445),
    .X(_0623_));
 sg13g2_nor2_1 _2752_ (.A(net429),
    .B(_0623_),
    .Y(_0624_));
 sg13g2_nor2_1 _2753_ (.A(_0717_),
    .B(net505),
    .Y(_0625_));
 sg13g2_a21oi_2 _2754_ (.B1(_0625_),
    .Y(_0626_),
    .A2(_0610_),
    .A1(_0602_));
 sg13g2_o21ai_1 _2755_ (.B1(net428),
    .Y(_0627_),
    .A1(_0620_),
    .A2(_0626_));
 sg13g2_a21oi_1 _2756_ (.A1(_0620_),
    .A2(_0626_),
    .Y(_0628_),
    .B1(_0627_));
 sg13g2_nor3_1 _2757_ (.A(net399),
    .B(_0624_),
    .C(_0628_),
    .Y(_0629_));
 sg13g2_a21oi_1 _2758_ (.A1(net484),
    .A2(net399),
    .Y(_0630_),
    .B1(_0629_));
 sg13g2_nand2_1 _2759_ (.Y(_0160_),
    .A(net526),
    .B(_0630_));
 sg13g2_a221oi_1 _2760_ (.B2(_0597_),
    .C1(_0592_),
    .B1(_0593_),
    .A1(net484),
    .Y(_0631_),
    .A2(_0576_));
 sg13g2_xnor2_1 _2761_ (.Y(_0632_),
    .A(\pqn_inst.n[12] ),
    .B(_0576_));
 sg13g2_nor3_2 _2762_ (.A(_0615_),
    .B(_0631_),
    .C(_0632_),
    .Y(_0633_));
 sg13g2_o21ai_1 _2763_ (.B1(_0632_),
    .Y(_0634_),
    .A1(_0615_),
    .A2(_0631_));
 sg13g2_nand2_1 _2764_ (.Y(_0635_),
    .A(net442),
    .B(_0634_));
 sg13g2_and2_1 _2765_ (.A(\pqn_inst.n[12] ),
    .B(\pqn_inst.multi.result[12] ),
    .X(_0636_));
 sg13g2_xor2_1 _2766_ (.B(net504),
    .A(\pqn_inst.n[12] ),
    .X(_0637_));
 sg13g2_xnor2_1 _2767_ (.Y(_0638_),
    .A(\pqn_inst.n[12] ),
    .B(net504));
 sg13g2_o21ai_1 _2768_ (.B1(_0618_),
    .Y(_0639_),
    .A1(_0600_),
    .A2(_0605_));
 sg13g2_nand3_1 _2769_ (.B(_0638_),
    .C(_0639_),
    .A(_0619_),
    .Y(_0640_));
 sg13g2_a21oi_2 _2770_ (.B1(_0638_),
    .Y(_0641_),
    .A2(_0639_),
    .A1(_0619_));
 sg13g2_nand3b_1 _2771_ (.B(net445),
    .C(_0640_),
    .Y(_0642_),
    .A_N(_0641_));
 sg13g2_o21ai_1 _2772_ (.B1(_0642_),
    .Y(_0643_),
    .A1(_0633_),
    .A2(_0635_));
 sg13g2_nand2_1 _2773_ (.Y(_0644_),
    .A(net484),
    .B(_0766_));
 sg13g2_nor2_1 _2774_ (.A(net484),
    .B(_0766_),
    .Y(_0645_));
 sg13g2_a21o_1 _2775_ (.A2(_0644_),
    .A1(_0626_),
    .B1(_0645_),
    .X(_0646_));
 sg13g2_a21oi_1 _2776_ (.A1(_0626_),
    .A2(_0644_),
    .Y(_0647_),
    .B1(_0645_));
 sg13g2_nand2_1 _2777_ (.Y(_0648_),
    .A(_0638_),
    .B(_0647_));
 sg13g2_a21oi_1 _2778_ (.A1(_0637_),
    .A2(_0646_),
    .Y(_0649_),
    .B1(net427));
 sg13g2_a221oi_1 _2779_ (.B2(_0649_),
    .C1(net398),
    .B1(_0648_),
    .A1(net427),
    .Y(_0650_),
    .A2(_0643_));
 sg13g2_o21ai_1 _2780_ (.B1(net527),
    .Y(_0651_),
    .A1(net269),
    .A2(_0456_));
 sg13g2_nor2_1 _2781_ (.A(_0650_),
    .B(_0651_),
    .Y(_0161_));
 sg13g2_or2_1 _2782_ (.X(_0652_),
    .B(\pqn_inst.multi.result[13] ),
    .A(\pqn_inst.n[13] ));
 sg13g2_nand2_1 _2783_ (.Y(_0653_),
    .A(\pqn_inst.n[13] ),
    .B(\pqn_inst.multi.result[13] ));
 sg13g2_and2_1 _2784_ (.A(_0652_),
    .B(_0653_),
    .X(_0654_));
 sg13g2_nor2_1 _2785_ (.A(_0636_),
    .B(_0641_),
    .Y(_0655_));
 sg13g2_a21oi_1 _2786_ (.A1(_0654_),
    .A2(_0655_),
    .Y(_0656_),
    .B1(net442));
 sg13g2_o21ai_1 _2787_ (.B1(_0656_),
    .Y(_0657_),
    .A1(_0654_),
    .A2(_0655_));
 sg13g2_a21oi_1 _2788_ (.A1(_0779_),
    .A2(_0576_),
    .Y(_0658_),
    .B1(_0633_));
 sg13g2_xnor2_1 _2789_ (.Y(_0659_),
    .A(\pqn_inst.n[13] ),
    .B(_0576_));
 sg13g2_xnor2_1 _2790_ (.Y(_0660_),
    .A(_0658_),
    .B(_0659_));
 sg13g2_a21oi_1 _2791_ (.A1(net442),
    .A2(_0660_),
    .Y(_0661_),
    .B1(net429));
 sg13g2_nor2b_1 _2792_ (.A(net504),
    .B_N(\pqn_inst.n[12] ),
    .Y(_0662_));
 sg13g2_a21oi_2 _2793_ (.B1(_0662_),
    .Y(_0663_),
    .A2(_0647_),
    .A1(_0638_));
 sg13g2_o21ai_1 _2794_ (.B1(net429),
    .Y(_0664_),
    .A1(_0654_),
    .A2(_0663_));
 sg13g2_a21oi_1 _2795_ (.A1(_0654_),
    .A2(_0663_),
    .Y(_0665_),
    .B1(_0664_));
 sg13g2_a21oi_1 _2796_ (.A1(_0657_),
    .A2(_0661_),
    .Y(_0666_),
    .B1(_0665_));
 sg13g2_a21oi_1 _2797_ (.A1(net256),
    .A2(net398),
    .Y(_0667_),
    .B1(net513));
 sg13g2_o21ai_1 _2798_ (.B1(_0667_),
    .Y(_0162_),
    .A1(net398),
    .A2(_0666_));
 sg13g2_nand2_1 _2799_ (.Y(_0668_),
    .A(\pqn_inst.n[14] ),
    .B(net503));
 sg13g2_xnor2_1 _2800_ (.Y(_0669_),
    .A(\pqn_inst.n[14] ),
    .B(net503));
 sg13g2_nor2_1 _2801_ (.A(\pqn_inst.n[13] ),
    .B(_0765_),
    .Y(_0670_));
 sg13g2_nand2_1 _2802_ (.Y(_0671_),
    .A(\pqn_inst.n[13] ),
    .B(_0765_));
 sg13g2_o21ai_1 _2803_ (.B1(_0671_),
    .Y(_0672_),
    .A1(_0663_),
    .A2(_0670_));
 sg13g2_xnor2_1 _2804_ (.Y(_0673_),
    .A(_0669_),
    .B(_0672_));
 sg13g2_o21ai_1 _2805_ (.B1(_0652_),
    .Y(_0674_),
    .A1(_0636_),
    .A2(_0641_));
 sg13g2_nand3_1 _2806_ (.B(_0669_),
    .C(_0674_),
    .A(_0653_),
    .Y(_0675_));
 sg13g2_a21o_1 _2807_ (.A2(_0674_),
    .A1(_0653_),
    .B1(_0669_),
    .X(_0676_));
 sg13g2_nand3_1 _2808_ (.B(_0675_),
    .C(_0676_),
    .A(net445),
    .Y(_0677_));
 sg13g2_or4_1 _2809_ (.A(_0615_),
    .B(_0631_),
    .C(_0632_),
    .D(_0659_),
    .X(_0678_));
 sg13g2_o21ai_1 _2810_ (.B1(_0001_),
    .Y(_0679_),
    .A1(\pqn_inst.n[13] ),
    .A2(_0000_));
 sg13g2_nand2_1 _2811_ (.Y(_0680_),
    .A(_0576_),
    .B(_0679_));
 sg13g2_nand2_1 _2812_ (.Y(_0681_),
    .A(_0678_),
    .B(_0680_));
 sg13g2_xnor2_1 _2813_ (.Y(_0682_),
    .A(\pqn_inst.n[14] ),
    .B(_0576_));
 sg13g2_a21oi_1 _2814_ (.A1(_0678_),
    .A2(_0680_),
    .Y(_0683_),
    .B1(_0682_));
 sg13g2_xnor2_1 _2815_ (.Y(_0684_),
    .A(_0681_),
    .B(_0682_));
 sg13g2_a21oi_1 _2816_ (.A1(net442),
    .A2(_0684_),
    .Y(_0685_),
    .B1(net429));
 sg13g2_a221oi_1 _2817_ (.B2(_0685_),
    .C1(net398),
    .B1(_0677_),
    .A1(net429),
    .Y(_0686_),
    .A2(_0673_));
 sg13g2_a21oi_1 _2818_ (.A1(net250),
    .A2(net398),
    .Y(_0687_),
    .B1(net510));
 sg13g2_nand2b_1 _2819_ (.Y(_0163_),
    .B(_0687_),
    .A_N(_0686_));
 sg13g2_xor2_1 _2820_ (.B(\pqn_inst.multi.result[15] ),
    .A(\pqn_inst.n[15] ),
    .X(_0688_));
 sg13g2_a21o_1 _2821_ (.A2(_0676_),
    .A1(_0668_),
    .B1(_0688_),
    .X(_0689_));
 sg13g2_nand3_1 _2822_ (.B(_0676_),
    .C(_0688_),
    .A(_0668_),
    .Y(_0690_));
 sg13g2_nand3_1 _2823_ (.B(_0689_),
    .C(_0690_),
    .A(net445),
    .Y(_0691_));
 sg13g2_nand2_1 _2824_ (.Y(_0692_),
    .A(_0002_),
    .B(_0576_));
 sg13g2_nand4_1 _2825_ (.B(\pqn_inst.n[13] ),
    .C(_0575_),
    .A(\pqn_inst.n[14] ),
    .Y(_0693_),
    .D(_0633_));
 sg13g2_o21ai_1 _2826_ (.B1(_0693_),
    .Y(_0694_),
    .A1(_0683_),
    .A2(_0692_));
 sg13g2_xnor2_1 _2827_ (.Y(_0695_),
    .A(\pqn_inst.n[15] ),
    .B(_0694_));
 sg13g2_a21oi_1 _2828_ (.A1(net442),
    .A2(_0695_),
    .Y(_0696_),
    .B1(net429));
 sg13g2_nor2b_1 _2829_ (.A(net503),
    .B_N(\pqn_inst.n[14] ),
    .Y(_0697_));
 sg13g2_a21oi_1 _2830_ (.A1(_0669_),
    .A2(_0672_),
    .Y(_0698_),
    .B1(_0697_));
 sg13g2_or2_1 _2831_ (.X(_0699_),
    .B(_0698_),
    .A(_0688_));
 sg13g2_a21oi_1 _2832_ (.A1(_0688_),
    .A2(_0698_),
    .Y(_0700_),
    .B1(net427));
 sg13g2_a22oi_1 _2833_ (.Y(_0701_),
    .B1(_0699_),
    .B2(_0700_),
    .A2(_0696_),
    .A1(_0691_));
 sg13g2_a21oi_1 _2834_ (.A1(net207),
    .A2(net398),
    .Y(_0702_),
    .B1(net510));
 sg13g2_o21ai_1 _2835_ (.B1(_0702_),
    .Y(_0164_),
    .A1(net398),
    .A2(_0701_));
 sg13g2_xnor2_1 _2836_ (.Y(_0703_),
    .A(net483),
    .B(_1168_));
 sg13g2_nor2_1 _2837_ (.A(net514),
    .B(_0703_),
    .Y(_0165_));
 sg13g2_o21ai_1 _2838_ (.B1(_1166_),
    .Y(_0704_),
    .A1(_1170_),
    .A2(_1175_));
 sg13g2_o21ai_1 _2839_ (.B1(_0704_),
    .Y(_0705_),
    .A1(net213),
    .A2(_1166_));
 sg13g2_nor2_1 _2840_ (.A(net516),
    .B(_0705_),
    .Y(_0166_));
 sg13g2_and2_1 _2841_ (.A(_1168_),
    .B(_1175_),
    .X(_0706_));
 sg13g2_o21ai_1 _2842_ (.B1(net526),
    .Y(_0707_),
    .A1(net173),
    .A2(_0706_));
 sg13g2_a21oi_1 _2843_ (.A1(net173),
    .A2(_0706_),
    .Y(_0167_),
    .B1(_0707_));
 sg13g2_and2_1 _2844_ (.A(net526),
    .B(_0426_),
    .X(_0168_));
 sg13g2_nor2_2 _2845_ (.A(_1170_),
    .B(_0455_),
    .Y(_0708_));
 sg13g2_a21oi_1 _2846_ (.A1(\pqn_inst.multi.result[0] ),
    .A2(_0708_),
    .Y(_0709_),
    .B1(net162));
 sg13g2_and3_1 _2847_ (.X(_0710_),
    .A(net162),
    .B(\pqn_inst.multi.result[0] ),
    .C(_0708_));
 sg13g2_nor3_1 _2848_ (.A(net515),
    .B(net163),
    .C(_0710_),
    .Y(_0169_));
 sg13g2_nand2_1 _2849_ (.Y(_0711_),
    .A(net293),
    .B(net426));
 sg13g2_xnor2_1 _2850_ (.Y(_0712_),
    .A(_0458_),
    .B(_0459_));
 sg13g2_xnor2_1 _2851_ (.Y(_0713_),
    .A(_0711_),
    .B(_0712_));
 sg13g2_o21ai_1 _2852_ (.B1(net528),
    .Y(_0714_),
    .A1(net235),
    .A2(_0708_));
 sg13g2_a21oi_1 _2853_ (.A1(_0708_),
    .A2(_0713_),
    .Y(_0170_),
    .B1(_0714_));
 sg13g2_dfrbp_1 _2854_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net120),
    .D(_0055_),
    .Q_N(_1426_),
    .Q(\pqn_inst.multi.temp[0] ));
 sg13g2_dfrbp_1 _2855_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net104),
    .D(_0056_),
    .Q_N(_1425_),
    .Q(\pqn_inst.multi.temp[1] ));
 sg13g2_dfrbp_1 _2856_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net102),
    .D(net139),
    .Q_N(_0034_),
    .Q(\pqn_inst.multi.temp[2] ));
 sg13g2_dfrbp_1 _2857_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net100),
    .D(net223),
    .Q_N(_1424_),
    .Q(\pqn_inst.multi.temp[3] ));
 sg13g2_dfrbp_1 _2858_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net98),
    .D(net161),
    .Q_N(_0037_),
    .Q(\pqn_inst.multi.temp[4] ));
 sg13g2_dfrbp_1 _2859_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net96),
    .D(net204),
    .Q_N(_1423_),
    .Q(\pqn_inst.multi.temp[5] ));
 sg13g2_dfrbp_1 _2860_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net94),
    .D(_0061_),
    .Q_N(_1422_),
    .Q(\pqn_inst.multi.temp[6] ));
 sg13g2_dfrbp_1 _2861_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net92),
    .D(net226),
    .Q_N(_1421_),
    .Q(\pqn_inst.multi.temp[7] ));
 sg13g2_dfrbp_1 _2862_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net90),
    .D(net172),
    .Q_N(_1420_),
    .Q(\pqn_inst.multi.temp[8] ));
 sg13g2_dfrbp_1 _2863_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net88),
    .D(_0064_),
    .Q_N(_1419_),
    .Q(\pqn_inst.multi.temp[9] ));
 sg13g2_dfrbp_1 _2864_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net86),
    .D(_0065_),
    .Q_N(_0017_),
    .Q(\pqn_inst.multi.result[0] ));
 sg13g2_dfrbp_1 _2865_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net84),
    .D(_0066_),
    .Q_N(_0019_),
    .Q(\pqn_inst.multi.result[1] ));
 sg13g2_dfrbp_1 _2866_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net82),
    .D(_0067_),
    .Q_N(_0020_),
    .Q(\pqn_inst.multi.result[2] ));
 sg13g2_dfrbp_1 _2867_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net80),
    .D(_0068_),
    .Q_N(_0021_),
    .Q(\pqn_inst.multi.result[3] ));
 sg13g2_dfrbp_1 _2868_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net78),
    .D(_0069_),
    .Q_N(_0023_),
    .Q(\pqn_inst.multi.result[4] ));
 sg13g2_dfrbp_1 _2869_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net76),
    .D(_0070_),
    .Q_N(_1418_),
    .Q(\pqn_inst.multi.result[5] ));
 sg13g2_dfrbp_1 _2870_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net74),
    .D(_0071_),
    .Q_N(_1417_),
    .Q(\pqn_inst.multi.result[6] ));
 sg13g2_dfrbp_1 _2871_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net72),
    .D(_0072_),
    .Q_N(_1416_),
    .Q(\pqn_inst.multi.result[7] ));
 sg13g2_dfrbp_1 _2872_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net70),
    .D(_0073_),
    .Q_N(_1415_),
    .Q(\pqn_inst.multi.result[8] ));
 sg13g2_dfrbp_1 _2873_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net68),
    .D(net159),
    .Q_N(_1414_),
    .Q(\pqn_inst.multi.result[9] ));
 sg13g2_dfrbp_1 _2874_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net66),
    .D(_0075_),
    .Q_N(_1413_),
    .Q(\pqn_inst.multi.result[10] ));
 sg13g2_dfrbp_1 _2875_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net64),
    .D(_0076_),
    .Q_N(_1412_),
    .Q(\pqn_inst.multi.result[11] ));
 sg13g2_dfrbp_1 _2876_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net62),
    .D(_0077_),
    .Q_N(_0024_),
    .Q(\pqn_inst.multi.result[12] ));
 sg13g2_dfrbp_1 _2877_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net60),
    .D(net288),
    .Q_N(_0025_),
    .Q(\pqn_inst.multi.result[13] ));
 sg13g2_dfrbp_1 _2878_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net58),
    .D(_0079_),
    .Q_N(_0026_),
    .Q(\pqn_inst.multi.result[14] ));
 sg13g2_dfrbp_1 _2879_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net56),
    .D(net228),
    .Q_N(_0028_),
    .Q(\pqn_inst.multi.result[15] ));
 sg13g2_dfrbp_1 _2880_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net54),
    .D(_0081_),
    .Q_N(_0054_),
    .Q(\pqn_inst.multi.stage[0] ));
 sg13g2_dfrbp_1 _2881_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net52),
    .D(_0082_),
    .Q_N(_0032_),
    .Q(\pqn_inst.multi.stage[1] ));
 sg13g2_dfrbp_1 _2882_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net50),
    .D(_0083_),
    .Q_N(_0029_),
    .Q(\pqn_inst.multi.stage[2] ));
 sg13g2_dfrbp_1 _2883_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net48),
    .D(_0084_),
    .Q_N(_0031_),
    .Q(\pqn_inst.multi.stage[3] ));
 sg13g2_dfrbp_1 _2884_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net46),
    .D(_0085_),
    .Q_N(_1411_),
    .Q(\pqn_inst.multi.start ));
 sg13g2_dfrbp_1 _2885_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net45),
    .D(_0086_),
    .Q_N(_1410_),
    .Q(\pqn_inst.b[0] ));
 sg13g2_dfrbp_1 _2886_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net43),
    .D(net136),
    .Q_N(_1409_),
    .Q(\pqn_inst.b[1] ));
 sg13g2_dfrbp_1 _2887_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net41),
    .D(_0088_),
    .Q_N(_1408_),
    .Q(\pqn_inst.b[2] ));
 sg13g2_dfrbp_1 _2888_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net39),
    .D(_0089_),
    .Q_N(_1407_),
    .Q(\pqn_inst.b[3] ));
 sg13g2_dfrbp_1 _2889_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net37),
    .D(_0090_),
    .Q_N(_1406_),
    .Q(\pqn_inst.b[4] ));
 sg13g2_dfrbp_1 _2890_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net35),
    .D(_0091_),
    .Q_N(_1405_),
    .Q(\pqn_inst.b[5] ));
 sg13g2_dfrbp_1 _2891_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net33),
    .D(_0092_),
    .Q_N(_1404_),
    .Q(\pqn_inst.b[6] ));
 sg13g2_dfrbp_1 _2892_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net31),
    .D(_0093_),
    .Q_N(_1403_),
    .Q(\pqn_inst.b[7] ));
 sg13g2_dfrbp_1 _2893_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net29),
    .D(_0094_),
    .Q_N(_1402_),
    .Q(\pqn_inst.b[8] ));
 sg13g2_dfrbp_1 _2894_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net27),
    .D(_0095_),
    .Q_N(_1401_),
    .Q(\pqn_inst.b[9] ));
 sg13g2_dfrbp_1 _2895_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net25),
    .D(_0096_),
    .Q_N(_1400_),
    .Q(\pqn_inst.b[10] ));
 sg13g2_dfrbp_1 _2896_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net23),
    .D(_0097_),
    .Q_N(_1399_),
    .Q(\pqn_inst.b[11] ));
 sg13g2_dfrbp_1 _2897_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net21),
    .D(_0098_),
    .Q_N(_1398_),
    .Q(\pqn_inst.b[12] ));
 sg13g2_dfrbp_1 _2898_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net19),
    .D(net180),
    .Q_N(_1397_),
    .Q(\pqn_inst.b[13] ));
 sg13g2_dfrbp_1 _2899_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net17),
    .D(net182),
    .Q_N(_1396_),
    .Q(\pqn_inst.b[14] ));
 sg13g2_dfrbp_1 _2900_ (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net15),
    .D(net196),
    .Q_N(_1395_),
    .Q(\pqn_inst.b[15] ));
 sg13g2_dfrbp_1 _2901_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net13),
    .D(_0102_),
    .Q_N(_1394_),
    .Q(\pqn_inst.v[0] ));
 sg13g2_dfrbp_1 _2902_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net11),
    .D(_0103_),
    .Q_N(_1393_),
    .Q(\pqn_inst.v[1] ));
 sg13g2_dfrbp_1 _2903_ (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net9),
    .D(_0104_),
    .Q_N(_1392_),
    .Q(\pqn_inst.v[2] ));
 sg13g2_dfrbp_1 _2904_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net123),
    .D(_0105_),
    .Q_N(_1391_),
    .Q(\pqn_inst.v[3] ));
 sg13g2_dfrbp_1 _2905_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net121),
    .D(_0106_),
    .Q_N(_1390_),
    .Q(\pqn_inst.v[4] ));
 sg13g2_dfrbp_1 _2906_ (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net119),
    .D(_0107_),
    .Q_N(_1389_),
    .Q(\pqn_inst.v[5] ));
 sg13g2_dfrbp_1 _2907_ (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net117),
    .D(_0108_),
    .Q_N(_1388_),
    .Q(\pqn_inst.v[6] ));
 sg13g2_dfrbp_1 _2908_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net115),
    .D(_0109_),
    .Q_N(_1387_),
    .Q(\pqn_inst.v[7] ));
 sg13g2_dfrbp_1 _2909_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net113),
    .D(_0110_),
    .Q_N(_1386_),
    .Q(\pqn_inst.v[8] ));
 sg13g2_dfrbp_1 _2910_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net111),
    .D(_0111_),
    .Q_N(_1385_),
    .Q(\pqn_inst.v[9] ));
 sg13g2_dfrbp_1 _2911_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net109),
    .D(_0112_),
    .Q_N(_1384_),
    .Q(\pqn_inst.v[10] ));
 sg13g2_dfrbp_1 _2912_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net107),
    .D(_0113_),
    .Q_N(_1383_),
    .Q(\pqn_inst.v[11] ));
 sg13g2_dfrbp_1 _2913_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net105),
    .D(_0114_),
    .Q_N(_1382_),
    .Q(\pqn_inst.v[12] ));
 sg13g2_dfrbp_1 _2914_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net101),
    .D(_0115_),
    .Q_N(_1381_),
    .Q(\pqn_inst.v[13] ));
 sg13g2_dfrbp_1 _2915_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net97),
    .D(_0116_),
    .Q_N(_1380_),
    .Q(\pqn_inst.v[14] ));
 sg13g2_dfrbp_1 _2916_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net93),
    .D(_0117_),
    .Q_N(_1379_),
    .Q(\pqn_inst.v[15] ));
 sg13g2_dfrbp_1 _2917_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net89),
    .D(net186),
    .Q_N(_0033_),
    .Q(\pqn_inst.a[0] ));
 sg13g2_dfrbp_1 _2918_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net85),
    .D(net176),
    .Q_N(_0030_),
    .Q(\pqn_inst.a[1] ));
 sg13g2_dfrbp_1 _2919_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net81),
    .D(net192),
    .Q_N(_0035_),
    .Q(\pqn_inst.a[2] ));
 sg13g2_dfrbp_1 _2920_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net77),
    .D(_0121_),
    .Q_N(_0036_),
    .Q(\pqn_inst.a[3] ));
 sg13g2_dfrbp_1 _2921_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net73),
    .D(_0122_),
    .Q_N(_0038_),
    .Q(\pqn_inst.a[4] ));
 sg13g2_dfrbp_1 _2922_ (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net69),
    .D(net190),
    .Q_N(_0039_),
    .Q(\pqn_inst.a[5] ));
 sg13g2_dfrbp_1 _2923_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net65),
    .D(net134),
    .Q_N(_0040_),
    .Q(\pqn_inst.a[6] ));
 sg13g2_dfrbp_1 _2924_ (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net61),
    .D(net198),
    .Q_N(_0041_),
    .Q(\pqn_inst.a[7] ));
 sg13g2_dfrbp_1 _2925_ (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net57),
    .D(_0126_),
    .Q_N(_0042_),
    .Q(\pqn_inst.a[8] ));
 sg13g2_dfrbp_1 _2926_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net53),
    .D(_0127_),
    .Q_N(_0043_),
    .Q(\pqn_inst.a[9] ));
 sg13g2_dfrbp_1 _2927_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net49),
    .D(_0128_),
    .Q_N(_0044_),
    .Q(\pqn_inst.a[10] ));
 sg13g2_dfrbp_1 _2928_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net44),
    .D(_0129_),
    .Q_N(_0045_),
    .Q(\pqn_inst.a[11] ));
 sg13g2_dfrbp_1 _2929_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net40),
    .D(_0130_),
    .Q_N(_0046_),
    .Q(\pqn_inst.a[12] ));
 sg13g2_dfrbp_1 _2930_ (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net36),
    .D(_0131_),
    .Q_N(_0047_),
    .Q(\pqn_inst.a[13] ));
 sg13g2_dfrbp_1 _2931_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net32),
    .D(_0132_),
    .Q_N(_0048_),
    .Q(\pqn_inst.a[14] ));
 sg13g2_dfrbp_1 _2932_ (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net28),
    .D(_0133_),
    .Q_N(_1378_),
    .Q(\pqn_inst.a[15] ));
 sg13g2_dfrbp_1 _2933_ (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net24),
    .D(_0134_),
    .Q_N(_1377_),
    .Q(\pqn_inst.done ));
 sg13g2_dfrbp_1 _2934_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net22),
    .D(_0135_),
    .Q_N(_0003_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _2935_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net18),
    .D(net217),
    .Q_N(_0004_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _2936_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net14),
    .D(net215),
    .Q_N(_0006_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _2937_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net10),
    .D(net209),
    .Q_N(_0007_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _2938_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net122),
    .D(net252),
    .Q_N(_0022_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _2939_ (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net118),
    .D(net241),
    .Q_N(_0008_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _2940_ (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net114),
    .D(net246),
    .Q_N(_0009_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _2941_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net110),
    .D(net248),
    .Q_N(_0010_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _2942_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net106),
    .D(_0143_),
    .Q_N(_0011_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _2943_ (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net99),
    .D(net244),
    .Q_N(_0051_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _2944_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net91),
    .D(_0145_),
    .Q_N(_0012_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _2945_ (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net83),
    .D(net237),
    .Q_N(_0013_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _2946_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net75),
    .D(net206),
    .Q_N(_0014_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _2947_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net67),
    .D(net212),
    .Q_N(_0015_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _2948_ (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net59),
    .D(net202),
    .Q_N(_0005_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _2949_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net51),
    .D(_0150_),
    .Q_N(_0050_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _2950_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net42),
    .D(_0151_),
    .Q_N(_0049_),
    .Q(\pqn_inst.n[2] ));
 sg13g2_dfrbp_1 _2951_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net34),
    .D(_0152_),
    .Q_N(_0052_),
    .Q(\pqn_inst.n[3] ));
 sg13g2_dfrbp_1 _2952_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net26),
    .D(_0153_),
    .Q_N(_0053_),
    .Q(\pqn_inst.n[4] ));
 sg13g2_dfrbp_1 _2953_ (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net16),
    .D(_0154_),
    .Q_N(_1376_),
    .Q(\pqn_inst.n[5] ));
 sg13g2_dfrbp_1 _2954_ (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net124),
    .D(_0155_),
    .Q_N(_1375_),
    .Q(\pqn_inst.n[6] ));
 sg13g2_dfrbp_1 _2955_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net116),
    .D(_0156_),
    .Q_N(_1374_),
    .Q(\pqn_inst.n[7] ));
 sg13g2_dfrbp_1 _2956_ (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net108),
    .D(_0157_),
    .Q_N(_1373_),
    .Q(\pqn_inst.n[8] ));
 sg13g2_dfrbp_1 _2957_ (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net95),
    .D(_0158_),
    .Q_N(_1372_),
    .Q(\pqn_inst.n[9] ));
 sg13g2_dfrbp_1 _2958_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net79),
    .D(_0159_),
    .Q_N(_1371_),
    .Q(\pqn_inst.n[10] ));
 sg13g2_dfrbp_1 _2959_ (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net63),
    .D(_0160_),
    .Q_N(_1370_),
    .Q(\pqn_inst.n[11] ));
 sg13g2_dfrbp_1 _2960_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net47),
    .D(_0161_),
    .Q_N(_0000_),
    .Q(\pqn_inst.n[12] ));
 sg13g2_dfrbp_1 _2961_ (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net30),
    .D(_0162_),
    .Q_N(_0001_),
    .Q(\pqn_inst.n[13] ));
 sg13g2_dfrbp_1 _2962_ (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net12),
    .D(_0163_),
    .Q_N(_0002_),
    .Q(\pqn_inst.n[14] ));
 sg13g2_dfrbp_1 _2963_ (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net112),
    .D(_0164_),
    .Q_N(_0027_),
    .Q(\pqn_inst.n[15] ));
 sg13g2_dfrbp_1 _2964_ (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net87),
    .D(_0165_),
    .Q_N(_1369_),
    .Q(\pqn_inst.stage[0] ));
 sg13g2_dfrbp_1 _2965_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net55),
    .D(_0166_),
    .Q_N(_1368_),
    .Q(\pqn_inst.stage[1] ));
 sg13g2_dfrbp_1 _2966_ (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net20),
    .D(_0167_),
    .Q_N(_1367_),
    .Q(\pqn_inst.stage[2] ));
 sg13g2_dfrbp_1 _2967_ (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net103),
    .D(_0168_),
    .Q_N(_1366_),
    .Q(\pqn_inst.stage[3] ));
 sg13g2_dfrbp_1 _2968_ (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net38),
    .D(net164),
    .Q_N(_0016_),
    .Q(\pqn_inst.n[0] ));
 sg13g2_dfrbp_1 _2969_ (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net71),
    .D(_0170_),
    .Q_N(_0018_),
    .Q(\pqn_inst.n[1] ));
 sg13g2_tiehi _2937__10 (.L_HI(net10));
 sg13g2_tiehi _2902__11 (.L_HI(net11));
 sg13g2_tiehi _2962__12 (.L_HI(net12));
 sg13g2_tiehi _2901__13 (.L_HI(net13));
 sg13g2_tiehi _2936__14 (.L_HI(net14));
 sg13g2_tiehi _2900__15 (.L_HI(net15));
 sg13g2_tiehi _2953__16 (.L_HI(net16));
 sg13g2_tiehi _2899__17 (.L_HI(net17));
 sg13g2_tiehi _2935__18 (.L_HI(net18));
 sg13g2_tiehi _2898__19 (.L_HI(net19));
 sg13g2_tiehi _2966__20 (.L_HI(net20));
 sg13g2_tiehi _2897__21 (.L_HI(net21));
 sg13g2_tiehi _2934__22 (.L_HI(net22));
 sg13g2_tiehi _2896__23 (.L_HI(net23));
 sg13g2_tiehi _2933__24 (.L_HI(net24));
 sg13g2_tiehi _2895__25 (.L_HI(net25));
 sg13g2_tiehi _2952__26 (.L_HI(net26));
 sg13g2_tiehi _2894__27 (.L_HI(net27));
 sg13g2_tiehi _2932__28 (.L_HI(net28));
 sg13g2_tiehi _2893__29 (.L_HI(net29));
 sg13g2_tiehi _2961__30 (.L_HI(net30));
 sg13g2_tiehi _2892__31 (.L_HI(net31));
 sg13g2_tiehi _2931__32 (.L_HI(net32));
 sg13g2_tiehi _2891__33 (.L_HI(net33));
 sg13g2_tiehi _2951__34 (.L_HI(net34));
 sg13g2_tiehi _2890__35 (.L_HI(net35));
 sg13g2_tiehi _2930__36 (.L_HI(net36));
 sg13g2_tiehi _2889__37 (.L_HI(net37));
 sg13g2_tiehi _2968__38 (.L_HI(net38));
 sg13g2_tiehi _2888__39 (.L_HI(net39));
 sg13g2_tiehi _2929__40 (.L_HI(net40));
 sg13g2_tiehi _2887__41 (.L_HI(net41));
 sg13g2_tiehi _2950__42 (.L_HI(net42));
 sg13g2_tiehi _2886__43 (.L_HI(net43));
 sg13g2_tiehi _2928__44 (.L_HI(net44));
 sg13g2_tiehi _2885__45 (.L_HI(net45));
 sg13g2_tiehi _2884__46 (.L_HI(net46));
 sg13g2_tiehi _2960__47 (.L_HI(net47));
 sg13g2_tiehi _2883__48 (.L_HI(net48));
 sg13g2_tiehi _2927__49 (.L_HI(net49));
 sg13g2_tiehi _2882__50 (.L_HI(net50));
 sg13g2_tiehi _2949__51 (.L_HI(net51));
 sg13g2_tiehi _2881__52 (.L_HI(net52));
 sg13g2_tiehi _2926__53 (.L_HI(net53));
 sg13g2_tiehi _2880__54 (.L_HI(net54));
 sg13g2_tiehi _2965__55 (.L_HI(net55));
 sg13g2_tiehi _2879__56 (.L_HI(net56));
 sg13g2_tiehi _2925__57 (.L_HI(net57));
 sg13g2_tiehi _2878__58 (.L_HI(net58));
 sg13g2_tiehi _2948__59 (.L_HI(net59));
 sg13g2_tiehi _2877__60 (.L_HI(net60));
 sg13g2_tiehi _2924__61 (.L_HI(net61));
 sg13g2_tiehi _2876__62 (.L_HI(net62));
 sg13g2_tiehi _2959__63 (.L_HI(net63));
 sg13g2_tiehi _2875__64 (.L_HI(net64));
 sg13g2_tiehi _2923__65 (.L_HI(net65));
 sg13g2_tiehi _2874__66 (.L_HI(net66));
 sg13g2_tiehi _2947__67 (.L_HI(net67));
 sg13g2_tiehi _2873__68 (.L_HI(net68));
 sg13g2_tiehi _2922__69 (.L_HI(net69));
 sg13g2_tiehi _2872__70 (.L_HI(net70));
 sg13g2_tiehi _2969__71 (.L_HI(net71));
 sg13g2_tiehi _2871__72 (.L_HI(net72));
 sg13g2_tiehi _2921__73 (.L_HI(net73));
 sg13g2_tiehi _2870__74 (.L_HI(net74));
 sg13g2_tiehi _2946__75 (.L_HI(net75));
 sg13g2_tiehi _2869__76 (.L_HI(net76));
 sg13g2_tiehi _2920__77 (.L_HI(net77));
 sg13g2_tiehi _2868__78 (.L_HI(net78));
 sg13g2_tiehi _2958__79 (.L_HI(net79));
 sg13g2_tiehi _2867__80 (.L_HI(net80));
 sg13g2_tiehi _2919__81 (.L_HI(net81));
 sg13g2_tiehi _2866__82 (.L_HI(net82));
 sg13g2_tiehi _2945__83 (.L_HI(net83));
 sg13g2_tiehi _2865__84 (.L_HI(net84));
 sg13g2_tiehi _2918__85 (.L_HI(net85));
 sg13g2_tiehi _2864__86 (.L_HI(net86));
 sg13g2_tiehi _2964__87 (.L_HI(net87));
 sg13g2_tiehi _2863__88 (.L_HI(net88));
 sg13g2_tiehi _2917__89 (.L_HI(net89));
 sg13g2_tiehi _2862__90 (.L_HI(net90));
 sg13g2_tiehi _2944__91 (.L_HI(net91));
 sg13g2_tiehi _2861__92 (.L_HI(net92));
 sg13g2_tiehi _2916__93 (.L_HI(net93));
 sg13g2_tiehi _2860__94 (.L_HI(net94));
 sg13g2_tiehi _2957__95 (.L_HI(net95));
 sg13g2_tiehi _2859__96 (.L_HI(net96));
 sg13g2_tiehi _2915__97 (.L_HI(net97));
 sg13g2_tiehi _2858__98 (.L_HI(net98));
 sg13g2_tiehi _2943__99 (.L_HI(net99));
 sg13g2_tiehi _2857__100 (.L_HI(net100));
 sg13g2_tiehi _2914__101 (.L_HI(net101));
 sg13g2_tiehi _2856__102 (.L_HI(net102));
 sg13g2_tiehi _2967__103 (.L_HI(net103));
 sg13g2_tiehi _2855__104 (.L_HI(net104));
 sg13g2_tiehi _2913__105 (.L_HI(net105));
 sg13g2_tiehi _2942__106 (.L_HI(net106));
 sg13g2_tiehi _2912__107 (.L_HI(net107));
 sg13g2_tiehi _2956__108 (.L_HI(net108));
 sg13g2_tiehi _2911__109 (.L_HI(net109));
 sg13g2_tiehi _2941__110 (.L_HI(net110));
 sg13g2_tiehi _2910__111 (.L_HI(net111));
 sg13g2_tiehi _2963__112 (.L_HI(net112));
 sg13g2_tiehi _2909__113 (.L_HI(net113));
 sg13g2_tiehi _2940__114 (.L_HI(net114));
 sg13g2_tiehi _2908__115 (.L_HI(net115));
 sg13g2_tiehi _2955__116 (.L_HI(net116));
 sg13g2_tiehi _2907__117 (.L_HI(net117));
 sg13g2_tiehi _2939__118 (.L_HI(net118));
 sg13g2_tiehi _2906__119 (.L_HI(net119));
 sg13g2_tiehi _2854__120 (.L_HI(net120));
 sg13g2_tiehi _2905__121 (.L_HI(net121));
 sg13g2_tiehi _2938__122 (.L_HI(net122));
 sg13g2_tiehi _2904__123 (.L_HI(net123));
 sg13g2_tiehi _2954__124 (.L_HI(net124));
 sg13g2_tiehi tt_um_pqn_125 (.L_HI(net125));
 sg13g2_tiehi tt_um_pqn_126 (.L_HI(net126));
 sg13g2_tiehi tt_um_pqn_127 (.L_HI(net127));
 sg13g2_tiehi tt_um_pqn_128 (.L_HI(net128));
 sg13g2_tiehi tt_um_pqn_129 (.L_HI(net129));
 sg13g2_tiehi tt_um_pqn_130 (.L_HI(net130));
 sg13g2_tiehi tt_um_pqn_131 (.L_HI(net131));
 sg13g2_tiehi tt_um_pqn_132 (.L_HI(net132));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 fanout398 (.A(net399),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_0457_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_0457_),
    .X(net400));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(_1184_));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(_1184_));
 sg13g2_buf_2 fanout403 (.A(_0427_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_0427_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(net406),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(net407),
    .X(net406));
 sg13g2_buf_1 fanout407 (.A(_0427_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_1196_),
    .X(net408));
 sg13g2_buf_4 fanout409 (.X(net409),
    .A(_1179_));
 sg13g2_buf_2 fanout410 (.A(_1179_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_0383_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_1289_),
    .X(net412));
 sg13g2_buf_1 fanout413 (.A(_1289_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(net415),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_1289_),
    .X(net415));
 sg13g2_buf_4 fanout416 (.X(net416),
    .A(_1200_));
 sg13g2_buf_4 fanout417 (.X(net417),
    .A(_1195_));
 sg13g2_buf_2 fanout418 (.A(_1178_),
    .X(net418));
 sg13g2_buf_1 fanout419 (.A(net420),
    .X(net419));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(_1178_));
 sg13g2_buf_2 fanout421 (.A(net422),
    .X(net421));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(_1299_));
 sg13g2_buf_1 fanout423 (.A(_1299_),
    .X(net423));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(_1298_));
 sg13g2_buf_2 fanout425 (.A(net426),
    .X(net425));
 sg13g2_buf_4 fanout426 (.X(net426),
    .A(net427));
 sg13g2_buf_4 fanout427 (.X(net427),
    .A(_1188_));
 sg13g2_buf_2 fanout428 (.A(net429),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(net430),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(net433),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(net432),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(net433),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_1187_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(net435),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_0803_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_0803_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(net439),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_0798_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(net441),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_0798_),
    .X(net441));
 sg13g2_buf_4 fanout442 (.X(net442),
    .A(_1191_));
 sg13g2_buf_2 fanout443 (.A(_1191_),
    .X(net443));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(net445));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(_1190_));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(_1186_));
 sg13g2_buf_4 fanout447 (.X(net447),
    .A(_1185_));
 sg13g2_buf_4 fanout448 (.X(net448),
    .A(_1183_));
 sg13g2_buf_2 fanout449 (.A(_1182_),
    .X(net449));
 sg13g2_buf_1 fanout450 (.A(_1182_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(net452),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_1182_),
    .X(net452));
 sg13g2_buf_4 fanout453 (.X(net453),
    .A(_0816_));
 sg13g2_buf_2 fanout454 (.A(net456),
    .X(net454));
 sg13g2_buf_1 fanout455 (.A(net456),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_0788_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(net458),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_0788_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(net461),
    .X(net459));
 sg13g2_buf_1 fanout460 (.A(net461),
    .X(net460));
 sg13g2_buf_1 fanout461 (.A(_0788_),
    .X(net461));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(_0831_));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(_0817_));
 sg13g2_buf_2 fanout464 (.A(_0767_),
    .X(net464));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(net466));
 sg13g2_buf_4 fanout466 (.X(net466),
    .A(_0762_));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(_0762_));
 sg13g2_buf_2 fanout468 (.A(_0762_),
    .X(net468));
 sg13g2_buf_4 fanout469 (.X(net469),
    .A(net472));
 sg13g2_buf_4 fanout470 (.X(net470),
    .A(net472));
 sg13g2_buf_2 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_0761_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(net474),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net476),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_0760_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(net479),
    .X(net477));
 sg13g2_buf_1 fanout478 (.A(net479),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_0759_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(\pqn_inst.stage[1] ),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(net483),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(net262),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(net282),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(net489),
    .X(net485));
 sg13g2_buf_4 fanout486 (.X(net486),
    .A(net488));
 sg13g2_buf_1 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(net489),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(\pqn_inst.done ),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(net278),
    .X(net490));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net158));
 sg13g2_buf_4 fanout492 (.X(net492),
    .A(net493));
 sg13g2_buf_4 fanout493 (.X(net493),
    .A(net158));
 sg13g2_buf_2 fanout494 (.A(_0031_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(net253),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(\pqn_inst.multi.stage[3] ),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_4 fanout498 (.X(net498),
    .A(\pqn_inst.multi.stage[2] ));
 sg13g2_buf_4 fanout499 (.X(net499),
    .A(net500));
 sg13g2_buf_4 fanout500 (.X(net500),
    .A(net280));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(net502));
 sg13g2_buf_4 fanout502 (.X(net502),
    .A(\pqn_inst.multi.stage[0] ));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(net277));
 sg13g2_buf_4 fanout504 (.X(net504),
    .A(net266));
 sg13g2_buf_4 fanout505 (.X(net505),
    .A(net292));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(net274));
 sg13g2_buf_4 fanout507 (.X(net507),
    .A(net281));
 sg13g2_buf_1 fanout508 (.A(\pqn_inst.multi.result[1] ),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net511),
    .X(net509));
 sg13g2_buf_1 fanout510 (.A(net511),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net518),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(net514),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(net518),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(net516),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(net518),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(net518),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_0786_),
    .X(net518));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(_0778_));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(net521));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(net522));
 sg13g2_buf_2 fanout522 (.A(net525),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(net524),
    .X(net523));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(net525));
 sg13g2_buf_2 fanout525 (.A(ui_in[0]),
    .X(net525));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(net527));
 sg13g2_buf_4 fanout527 (.X(net527),
    .A(net1));
 sg13g2_buf_4 fanout528 (.X(net528),
    .A(net529));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(net1));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tiehi _2903__9 (.L_HI(net9));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\pqn_inst.a[6] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0124_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold3 (.A(\pqn_inst.b[1] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0087_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold5 (.A(\pqn_inst.multi.temp[0] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold6 (.A(\pqn_inst.multi.temp[2] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0057_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold8 (.A(\pqn_inst.a[10] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0418_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold10 (.A(\pqn_inst.a[11] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0420_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold12 (.A(\pqn_inst.a[9] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0416_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold14 (.A(\pqn_inst.b[4] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold15 (.A(_1227_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold16 (.A(\pqn_inst.b[0] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold17 (.A(_1206_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold18 (.A(\pqn_inst.a[12] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0421_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold20 (.A(\pqn_inst.b[3] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold21 (.A(_1222_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold22 (.A(\pqn_inst.a[13] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0422_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold24 (.A(\pqn_inst.a[14] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0423_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold26 (.A(\pqn_inst.multi.start ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0074_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold28 (.A(\pqn_inst.multi.temp[4] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0059_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold30 (.A(\pqn_inst.n[0] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0709_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0169_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold33 (.A(\pqn_inst.multi.temp[6] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold34 (.A(\pqn_inst.b[12] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold35 (.A(_1270_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold36 (.A(\pqn_inst.a[3] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0371_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold38 (.A(\pqn_inst.a[4] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold39 (.A(\pqn_inst.multi.temp[8] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0063_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold41 (.A(\pqn_inst.stage[2] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold42 (.A(\pqn_inst.multi.temp[1] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold43 (.A(\pqn_inst.a[1] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0119_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0054_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold46 (.A(_1158_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold47 (.A(\pqn_inst.b[13] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0099_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold49 (.A(\pqn_inst.b[14] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0100_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold51 (.A(\pqn_inst.a[8] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0413_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold53 (.A(\pqn_inst.a[0] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0118_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold55 (.A(\pqn_inst.a[15] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0424_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold57 (.A(\pqn_inst.a[5] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0123_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold59 (.A(\pqn_inst.a[2] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0120_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold61 (.A(\pqn_inst.b[2] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold62 (.A(_1216_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold63 (.A(\pqn_inst.b[15] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0101_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold65 (.A(\pqn_inst.a[7] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0125_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold67 (.A(\pqn_inst.multi.temp[9] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold68 (.A(\pqn_inst.v[0] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold69 (.A(uio_out[6]),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0149_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold71 (.A(\pqn_inst.multi.temp[5] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0060_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold73 (.A(uio_out[4]),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0147_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold75 (.A(\pqn_inst.n[15] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold76 (.A(uo_out[3]),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0138_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold78 (.A(uo_out[0]),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold79 (.A(uio_out[5]),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0148_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold81 (.A(\pqn_inst.stage[1] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold82 (.A(uo_out[2]),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0137_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold84 (.A(uo_out[1]),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0136_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold86 (.A(\pqn_inst.n[2] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold87 (.A(\pqn_inst.b[11] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold88 (.A(\pqn_inst.b[8] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold89 (.A(\pqn_inst.b[7] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold90 (.A(\pqn_inst.multi.temp[3] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0058_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold92 (.A(\pqn_inst.b[10] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold93 (.A(\pqn_inst.multi.temp[7] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0062_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold95 (.A(\pqn_inst.multi.result[15] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0080_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold97 (.A(\pqn_inst.v[8] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold98 (.A(\pqn_inst.v[15] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold99 (.A(uio_out[7]),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold100 (.A(\pqn_inst.b[6] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold101 (.A(\pqn_inst.b[5] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold102 (.A(\pqn_inst.b[9] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold103 (.A(\pqn_inst.n[1] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold104 (.A(uio_out[3]),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0146_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold106 (.A(\pqn_inst.v[10] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold107 (.A(\pqn_inst.n[4] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold108 (.A(uo_out[5]),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0140_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold110 (.A(uio_out[0]),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold111 (.A(uio_out[1]),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0144_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold113 (.A(uo_out[6]),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0141_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold115 (.A(uo_out[7]),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0142_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold117 (.A(\pqn_inst.n[3] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold118 (.A(\pqn_inst.n[14] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold119 (.A(\pqn_inst.v[4] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0139_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold121 (.A(\pqn_inst.multi.stage[3] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold122 (.A(_1165_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold123 (.A(\pqn_inst.multi.result[2] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold124 (.A(\pqn_inst.n[13] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold125 (.A(\pqn_inst.n[7] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold126 (.A(uio_out[2]),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0029_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold128 (.A(\pqn_inst.v[12] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold129 (.A(\pqn_inst.n[10] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold130 (.A(\pqn_inst.stage[0] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold131 (.A(\pqn_inst.v[11] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold132 (.A(\pqn_inst.v[14] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold133 (.A(\pqn_inst.multi.result[8] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold134 (.A(\pqn_inst.multi.result[12] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold135 (.A(\pqn_inst.v[7] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold136 (.A(\pqn_inst.n[9] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold137 (.A(\pqn_inst.n[12] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold138 (.A(\pqn_inst.v[3] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold139 (.A(\pqn_inst.v[1] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0023_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold141 (.A(\pqn_inst.v[9] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold142 (.A(\pqn_inst.multi.result[4] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold143 (.A(\pqn_inst.v[2] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold144 (.A(\pqn_inst.n[8] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold145 (.A(\pqn_inst.multi.result[14] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold146 (.A(\pqn_inst.v[13] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold147 (.A(\pqn_inst.multi.result[11] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold148 (.A(\pqn_inst.multi.stage[1] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold149 (.A(\pqn_inst.multi.result[1] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold150 (.A(\pqn_inst.n[11] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold151 (.A(\pqn_inst.n[6] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold152 (.A(\pqn_inst.multi.result[0] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold153 (.A(\pqn_inst.multi.result[6] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold154 (.A(\pqn_inst.multi.result[3] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0024_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0078_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold157 (.A(\pqn_inst.n[5] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold158 (.A(\pqn_inst.v[5] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold159 (.A(\pqn_inst.v[6] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold160 (.A(\pqn_inst.multi.result[10] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold161 (.A(\pqn_inst.multi.result[0] ),
    .X(net293));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_4 FILLER_0_63 ();
 sg13g2_fill_2 FILLER_0_67 ();
 sg13g2_decap_8 FILLER_0_73 ();
 sg13g2_decap_8 FILLER_0_80 ();
 sg13g2_decap_8 FILLER_0_87 ();
 sg13g2_decap_8 FILLER_0_94 ();
 sg13g2_decap_8 FILLER_0_101 ();
 sg13g2_decap_8 FILLER_0_108 ();
 sg13g2_fill_2 FILLER_0_119 ();
 sg13g2_fill_1 FILLER_0_121 ();
 sg13g2_decap_4 FILLER_0_152 ();
 sg13g2_fill_2 FILLER_0_156 ();
 sg13g2_decap_8 FILLER_0_162 ();
 sg13g2_decap_8 FILLER_0_169 ();
 sg13g2_decap_8 FILLER_0_181 ();
 sg13g2_decap_8 FILLER_0_188 ();
 sg13g2_decap_4 FILLER_0_195 ();
 sg13g2_fill_1 FILLER_0_199 ();
 sg13g2_decap_4 FILLER_0_204 ();
 sg13g2_decap_4 FILLER_0_268 ();
 sg13g2_fill_2 FILLER_0_272 ();
 sg13g2_fill_1 FILLER_0_300 ();
 sg13g2_fill_2 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_4 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_fill_1 FILLER_1_83 ();
 sg13g2_decap_8 FILLER_1_93 ();
 sg13g2_decap_4 FILLER_1_100 ();
 sg13g2_fill_1 FILLER_1_135 ();
 sg13g2_fill_1 FILLER_1_146 ();
 sg13g2_fill_2 FILLER_1_215 ();
 sg13g2_fill_1 FILLER_1_217 ();
 sg13g2_fill_2 FILLER_1_246 ();
 sg13g2_fill_1 FILLER_1_248 ();
 sg13g2_decap_8 FILLER_1_271 ();
 sg13g2_fill_2 FILLER_1_278 ();
 sg13g2_fill_1 FILLER_1_280 ();
 sg13g2_fill_2 FILLER_1_295 ();
 sg13g2_fill_1 FILLER_1_297 ();
 sg13g2_decap_4 FILLER_1_315 ();
 sg13g2_fill_2 FILLER_1_345 ();
 sg13g2_fill_1 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_383 ();
 sg13g2_decap_8 FILLER_1_390 ();
 sg13g2_decap_8 FILLER_1_397 ();
 sg13g2_decap_4 FILLER_1_404 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_4 FILLER_2_42 ();
 sg13g2_decap_4 FILLER_2_94 ();
 sg13g2_fill_1 FILLER_2_133 ();
 sg13g2_fill_1 FILLER_2_190 ();
 sg13g2_fill_1 FILLER_2_199 ();
 sg13g2_decap_8 FILLER_2_250 ();
 sg13g2_fill_2 FILLER_2_257 ();
 sg13g2_fill_2 FILLER_2_286 ();
 sg13g2_fill_1 FILLER_2_288 ();
 sg13g2_fill_1 FILLER_2_294 ();
 sg13g2_fill_2 FILLER_2_303 ();
 sg13g2_fill_1 FILLER_2_305 ();
 sg13g2_fill_1 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_28 ();
 sg13g2_fill_1 FILLER_3_30 ();
 sg13g2_fill_1 FILLER_3_35 ();
 sg13g2_fill_1 FILLER_3_74 ();
 sg13g2_fill_2 FILLER_3_101 ();
 sg13g2_fill_1 FILLER_3_103 ();
 sg13g2_fill_2 FILLER_3_135 ();
 sg13g2_fill_1 FILLER_3_137 ();
 sg13g2_fill_1 FILLER_3_147 ();
 sg13g2_fill_1 FILLER_3_152 ();
 sg13g2_fill_1 FILLER_3_162 ();
 sg13g2_fill_2 FILLER_3_193 ();
 sg13g2_fill_1 FILLER_3_195 ();
 sg13g2_decap_4 FILLER_3_217 ();
 sg13g2_fill_1 FILLER_3_221 ();
 sg13g2_fill_1 FILLER_3_226 ();
 sg13g2_decap_8 FILLER_3_248 ();
 sg13g2_fill_2 FILLER_3_255 ();
 sg13g2_fill_1 FILLER_3_257 ();
 sg13g2_decap_8 FILLER_3_271 ();
 sg13g2_decap_8 FILLER_3_278 ();
 sg13g2_fill_1 FILLER_3_285 ();
 sg13g2_fill_1 FILLER_3_305 ();
 sg13g2_fill_1 FILLER_3_321 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_4 FILLER_4_14 ();
 sg13g2_fill_2 FILLER_4_18 ();
 sg13g2_fill_1 FILLER_4_46 ();
 sg13g2_fill_2 FILLER_4_81 ();
 sg13g2_fill_2 FILLER_4_98 ();
 sg13g2_fill_1 FILLER_4_100 ();
 sg13g2_fill_1 FILLER_4_136 ();
 sg13g2_decap_8 FILLER_4_185 ();
 sg13g2_decap_8 FILLER_4_192 ();
 sg13g2_fill_1 FILLER_4_199 ();
 sg13g2_decap_4 FILLER_4_221 ();
 sg13g2_fill_2 FILLER_4_283 ();
 sg13g2_decap_8 FILLER_4_307 ();
 sg13g2_fill_2 FILLER_4_314 ();
 sg13g2_fill_2 FILLER_4_353 ();
 sg13g2_fill_2 FILLER_4_360 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_4 FILLER_5_21 ();
 sg13g2_fill_2 FILLER_5_25 ();
 sg13g2_fill_1 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_111 ();
 sg13g2_decap_4 FILLER_5_118 ();
 sg13g2_fill_2 FILLER_5_122 ();
 sg13g2_fill_2 FILLER_5_138 ();
 sg13g2_fill_2 FILLER_5_169 ();
 sg13g2_fill_1 FILLER_5_171 ();
 sg13g2_decap_8 FILLER_5_193 ();
 sg13g2_decap_4 FILLER_5_221 ();
 sg13g2_fill_1 FILLER_5_225 ();
 sg13g2_decap_4 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_4 FILLER_5_252 ();
 sg13g2_decap_4 FILLER_5_277 ();
 sg13g2_fill_2 FILLER_5_289 ();
 sg13g2_decap_4 FILLER_5_322 ();
 sg13g2_fill_2 FILLER_5_326 ();
 sg13g2_fill_1 FILLER_5_363 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_fill_1 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_55 ();
 sg13g2_fill_1 FILLER_6_77 ();
 sg13g2_fill_2 FILLER_6_97 ();
 sg13g2_decap_8 FILLER_6_120 ();
 sg13g2_fill_1 FILLER_6_127 ();
 sg13g2_decap_8 FILLER_6_145 ();
 sg13g2_fill_1 FILLER_6_152 ();
 sg13g2_fill_1 FILLER_6_158 ();
 sg13g2_fill_2 FILLER_6_163 ();
 sg13g2_fill_1 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_171 ();
 sg13g2_fill_2 FILLER_6_178 ();
 sg13g2_decap_8 FILLER_6_190 ();
 sg13g2_decap_4 FILLER_6_218 ();
 sg13g2_fill_1 FILLER_6_222 ();
 sg13g2_fill_2 FILLER_6_233 ();
 sg13g2_fill_1 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_282 ();
 sg13g2_fill_2 FILLER_6_289 ();
 sg13g2_fill_2 FILLER_6_319 ();
 sg13g2_fill_1 FILLER_6_321 ();
 sg13g2_fill_2 FILLER_6_332 ();
 sg13g2_fill_1 FILLER_6_334 ();
 sg13g2_fill_2 FILLER_6_345 ();
 sg13g2_fill_1 FILLER_6_347 ();
 sg13g2_fill_2 FILLER_6_375 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_14 ();
 sg13g2_fill_1 FILLER_7_16 ();
 sg13g2_fill_2 FILLER_7_32 ();
 sg13g2_fill_2 FILLER_7_44 ();
 sg13g2_fill_1 FILLER_7_46 ();
 sg13g2_fill_1 FILLER_7_82 ();
 sg13g2_fill_2 FILLER_7_96 ();
 sg13g2_fill_2 FILLER_7_171 ();
 sg13g2_fill_1 FILLER_7_215 ();
 sg13g2_fill_2 FILLER_7_220 ();
 sg13g2_fill_1 FILLER_7_222 ();
 sg13g2_decap_4 FILLER_7_249 ();
 sg13g2_fill_1 FILLER_7_253 ();
 sg13g2_fill_2 FILLER_7_258 ();
 sg13g2_fill_2 FILLER_7_281 ();
 sg13g2_fill_1 FILLER_7_283 ();
 sg13g2_decap_8 FILLER_7_296 ();
 sg13g2_fill_1 FILLER_7_303 ();
 sg13g2_decap_4 FILLER_7_324 ();
 sg13g2_fill_1 FILLER_8_64 ();
 sg13g2_decap_4 FILLER_8_114 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_144 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_4 FILLER_8_188 ();
 sg13g2_fill_1 FILLER_8_192 ();
 sg13g2_decap_4 FILLER_8_208 ();
 sg13g2_fill_1 FILLER_8_227 ();
 sg13g2_fill_2 FILLER_8_262 ();
 sg13g2_decap_4 FILLER_8_282 ();
 sg13g2_fill_2 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_4 FILLER_8_312 ();
 sg13g2_fill_1 FILLER_8_316 ();
 sg13g2_decap_4 FILLER_8_325 ();
 sg13g2_fill_2 FILLER_8_329 ();
 sg13g2_fill_2 FILLER_8_336 ();
 sg13g2_fill_1 FILLER_8_338 ();
 sg13g2_fill_1 FILLER_8_343 ();
 sg13g2_fill_2 FILLER_8_365 ();
 sg13g2_fill_2 FILLER_8_381 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_5 ();
 sg13g2_fill_1 FILLER_9_38 ();
 sg13g2_fill_1 FILLER_9_43 ();
 sg13g2_fill_1 FILLER_9_58 ();
 sg13g2_decap_4 FILLER_9_95 ();
 sg13g2_fill_2 FILLER_9_131 ();
 sg13g2_fill_1 FILLER_9_160 ();
 sg13g2_decap_4 FILLER_9_234 ();
 sg13g2_fill_2 FILLER_9_238 ();
 sg13g2_decap_4 FILLER_9_255 ();
 sg13g2_fill_1 FILLER_9_270 ();
 sg13g2_fill_2 FILLER_9_310 ();
 sg13g2_decap_4 FILLER_9_343 ();
 sg13g2_fill_2 FILLER_9_347 ();
 sg13g2_fill_2 FILLER_9_363 ();
 sg13g2_decap_4 FILLER_9_389 ();
 sg13g2_fill_1 FILLER_9_393 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_39 ();
 sg13g2_fill_1 FILLER_10_92 ();
 sg13g2_fill_1 FILLER_10_97 ();
 sg13g2_decap_4 FILLER_10_109 ();
 sg13g2_decap_4 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_fill_2 FILLER_10_208 ();
 sg13g2_decap_4 FILLER_10_230 ();
 sg13g2_fill_2 FILLER_10_234 ();
 sg13g2_fill_2 FILLER_10_239 ();
 sg13g2_fill_1 FILLER_10_241 ();
 sg13g2_decap_4 FILLER_10_257 ();
 sg13g2_fill_2 FILLER_10_268 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_fill_1 FILLER_10_284 ();
 sg13g2_fill_2 FILLER_10_314 ();
 sg13g2_fill_1 FILLER_10_316 ();
 sg13g2_fill_1 FILLER_10_344 ();
 sg13g2_fill_2 FILLER_10_349 ();
 sg13g2_fill_2 FILLER_10_369 ();
 sg13g2_fill_1 FILLER_10_371 ();
 sg13g2_fill_1 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_fill_2 FILLER_11_13 ();
 sg13g2_fill_1 FILLER_11_25 ();
 sg13g2_fill_2 FILLER_11_36 ();
 sg13g2_fill_1 FILLER_11_63 ();
 sg13g2_fill_2 FILLER_11_137 ();
 sg13g2_fill_1 FILLER_11_139 ();
 sg13g2_fill_2 FILLER_11_154 ();
 sg13g2_fill_2 FILLER_11_165 ();
 sg13g2_fill_1 FILLER_11_167 ();
 sg13g2_decap_4 FILLER_11_183 ();
 sg13g2_decap_8 FILLER_11_206 ();
 sg13g2_decap_4 FILLER_11_213 ();
 sg13g2_fill_2 FILLER_11_279 ();
 sg13g2_fill_2 FILLER_11_305 ();
 sg13g2_decap_4 FILLER_11_321 ();
 sg13g2_fill_1 FILLER_11_325 ();
 sg13g2_fill_1 FILLER_11_363 ();
 sg13g2_fill_1 FILLER_11_382 ();
 sg13g2_fill_1 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_4 ();
 sg13g2_fill_1 FILLER_12_26 ();
 sg13g2_fill_1 FILLER_12_81 ();
 sg13g2_fill_2 FILLER_12_99 ();
 sg13g2_fill_1 FILLER_12_101 ();
 sg13g2_fill_1 FILLER_12_133 ();
 sg13g2_fill_2 FILLER_12_148 ();
 sg13g2_decap_4 FILLER_12_190 ();
 sg13g2_fill_1 FILLER_12_194 ();
 sg13g2_decap_8 FILLER_12_198 ();
 sg13g2_fill_2 FILLER_12_205 ();
 sg13g2_decap_4 FILLER_12_212 ();
 sg13g2_fill_1 FILLER_12_265 ();
 sg13g2_fill_1 FILLER_12_279 ();
 sg13g2_fill_2 FILLER_12_302 ();
 sg13g2_fill_1 FILLER_12_304 ();
 sg13g2_fill_1 FILLER_12_318 ();
 sg13g2_fill_2 FILLER_12_347 ();
 sg13g2_fill_1 FILLER_12_349 ();
 sg13g2_fill_1 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_4 ();
 sg13g2_decap_4 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_54 ();
 sg13g2_fill_1 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_75 ();
 sg13g2_fill_2 FILLER_13_85 ();
 sg13g2_fill_1 FILLER_13_113 ();
 sg13g2_fill_2 FILLER_13_127 ();
 sg13g2_fill_1 FILLER_13_142 ();
 sg13g2_fill_1 FILLER_13_166 ();
 sg13g2_fill_1 FILLER_13_267 ();
 sg13g2_fill_2 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_306 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_fill_2 FILLER_13_337 ();
 sg13g2_fill_1 FILLER_13_339 ();
 sg13g2_fill_2 FILLER_13_380 ();
 sg13g2_fill_1 FILLER_13_382 ();
 sg13g2_fill_2 FILLER_14_43 ();
 sg13g2_fill_2 FILLER_14_50 ();
 sg13g2_fill_2 FILLER_14_61 ();
 sg13g2_fill_2 FILLER_14_116 ();
 sg13g2_fill_2 FILLER_14_240 ();
 sg13g2_fill_2 FILLER_14_251 ();
 sg13g2_fill_2 FILLER_14_279 ();
 sg13g2_fill_1 FILLER_14_360 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_15_100 ();
 sg13g2_fill_1 FILLER_15_149 ();
 sg13g2_fill_2 FILLER_15_176 ();
 sg13g2_decap_4 FILLER_15_308 ();
 sg13g2_fill_2 FILLER_15_312 ();
 sg13g2_decap_4 FILLER_15_319 ();
 sg13g2_fill_1 FILLER_15_323 ();
 sg13g2_fill_1 FILLER_15_333 ();
 sg13g2_fill_2 FILLER_15_347 ();
 sg13g2_fill_1 FILLER_15_349 ();
 sg13g2_fill_1 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_63 ();
 sg13g2_fill_2 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_147 ();
 sg13g2_fill_1 FILLER_16_232 ();
 sg13g2_decap_4 FILLER_16_334 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_decap_4 FILLER_16_369 ();
 sg13g2_fill_1 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_4 ();
 sg13g2_fill_1 FILLER_17_36 ();
 sg13g2_fill_2 FILLER_17_45 ();
 sg13g2_fill_1 FILLER_17_57 ();
 sg13g2_fill_2 FILLER_17_92 ();
 sg13g2_fill_1 FILLER_17_120 ();
 sg13g2_fill_1 FILLER_17_126 ();
 sg13g2_fill_1 FILLER_17_136 ();
 sg13g2_fill_1 FILLER_17_176 ();
 sg13g2_fill_2 FILLER_17_214 ();
 sg13g2_fill_2 FILLER_17_228 ();
 sg13g2_fill_1 FILLER_17_250 ();
 sg13g2_fill_1 FILLER_17_285 ();
 sg13g2_fill_2 FILLER_17_299 ();
 sg13g2_fill_2 FILLER_17_329 ();
 sg13g2_fill_1 FILLER_17_331 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_100 ();
 sg13g2_fill_2 FILLER_18_111 ();
 sg13g2_fill_1 FILLER_18_117 ();
 sg13g2_fill_2 FILLER_18_161 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_fill_1 FILLER_18_174 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_fill_2 FILLER_18_252 ();
 sg13g2_fill_1 FILLER_18_254 ();
 sg13g2_fill_2 FILLER_18_274 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_fill_2 FILLER_18_325 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_fill_2 FILLER_18_341 ();
 sg13g2_fill_2 FILLER_18_357 ();
 sg13g2_fill_1 FILLER_18_359 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_2 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_23 ();
 sg13g2_fill_1 FILLER_19_29 ();
 sg13g2_decap_8 FILLER_19_38 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_fill_2 FILLER_19_59 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_2 FILLER_19_92 ();
 sg13g2_fill_1 FILLER_19_94 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_184 ();
 sg13g2_fill_1 FILLER_19_186 ();
 sg13g2_fill_2 FILLER_19_192 ();
 sg13g2_decap_4 FILLER_19_199 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_248 ();
 sg13g2_fill_2 FILLER_19_264 ();
 sg13g2_fill_1 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_293 ();
 sg13g2_fill_1 FILLER_19_304 ();
 sg13g2_fill_2 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_317 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_decap_4 FILLER_19_332 ();
 sg13g2_fill_1 FILLER_19_343 ();
 sg13g2_fill_2 FILLER_19_358 ();
 sg13g2_fill_2 FILLER_19_381 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_25 ();
 sg13g2_fill_1 FILLER_20_36 ();
 sg13g2_fill_2 FILLER_20_68 ();
 sg13g2_fill_1 FILLER_20_77 ();
 sg13g2_fill_2 FILLER_20_91 ();
 sg13g2_fill_1 FILLER_20_93 ();
 sg13g2_decap_8 FILLER_20_114 ();
 sg13g2_decap_8 FILLER_20_121 ();
 sg13g2_decap_8 FILLER_20_128 ();
 sg13g2_fill_1 FILLER_20_135 ();
 sg13g2_decap_4 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_166 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_decap_4 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_281 ();
 sg13g2_fill_1 FILLER_20_288 ();
 sg13g2_decap_8 FILLER_20_330 ();
 sg13g2_decap_4 FILLER_20_337 ();
 sg13g2_fill_1 FILLER_20_341 ();
 sg13g2_fill_2 FILLER_20_346 ();
 sg13g2_fill_1 FILLER_20_362 ();
 sg13g2_fill_2 FILLER_20_384 ();
 sg13g2_fill_1 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_decap_4 FILLER_21_21 ();
 sg13g2_decap_4 FILLER_21_38 ();
 sg13g2_fill_1 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_4 FILLER_21_63 ();
 sg13g2_fill_2 FILLER_21_67 ();
 sg13g2_decap_8 FILLER_21_74 ();
 sg13g2_fill_1 FILLER_21_81 ();
 sg13g2_fill_1 FILLER_21_96 ();
 sg13g2_fill_1 FILLER_21_136 ();
 sg13g2_fill_1 FILLER_21_153 ();
 sg13g2_decap_4 FILLER_21_178 ();
 sg13g2_fill_1 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_4 FILLER_21_231 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_fill_1 FILLER_21_241 ();
 sg13g2_fill_2 FILLER_21_251 ();
 sg13g2_fill_2 FILLER_21_258 ();
 sg13g2_fill_2 FILLER_21_284 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_fill_1 FILLER_21_333 ();
 sg13g2_decap_4 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_358 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_9 ();
 sg13g2_fill_2 FILLER_22_27 ();
 sg13g2_fill_1 FILLER_22_29 ();
 sg13g2_fill_1 FILLER_22_52 ();
 sg13g2_fill_2 FILLER_22_106 ();
 sg13g2_fill_1 FILLER_22_108 ();
 sg13g2_fill_2 FILLER_22_134 ();
 sg13g2_decap_4 FILLER_22_150 ();
 sg13g2_fill_1 FILLER_22_154 ();
 sg13g2_fill_2 FILLER_22_173 ();
 sg13g2_fill_2 FILLER_22_187 ();
 sg13g2_fill_1 FILLER_22_199 ();
 sg13g2_fill_2 FILLER_22_218 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_256 ();
 sg13g2_fill_1 FILLER_22_258 ();
 sg13g2_fill_1 FILLER_22_297 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_fill_2 FILLER_22_357 ();
 sg13g2_fill_1 FILLER_22_359 ();
 sg13g2_fill_1 FILLER_22_372 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_2 FILLER_23_17 ();
 sg13g2_fill_1 FILLER_23_19 ();
 sg13g2_decap_4 FILLER_23_34 ();
 sg13g2_fill_2 FILLER_23_38 ();
 sg13g2_fill_2 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_62 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_fill_1 FILLER_23_119 ();
 sg13g2_decap_4 FILLER_23_133 ();
 sg13g2_fill_2 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_4 FILLER_23_175 ();
 sg13g2_fill_2 FILLER_23_184 ();
 sg13g2_fill_2 FILLER_23_202 ();
 sg13g2_decap_4 FILLER_23_213 ();
 sg13g2_fill_2 FILLER_23_234 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_260 ();
 sg13g2_decap_4 FILLER_23_267 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_decap_4 FILLER_23_276 ();
 sg13g2_decap_4 FILLER_23_303 ();
 sg13g2_fill_2 FILLER_23_313 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_fill_2 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_24 ();
 sg13g2_fill_2 FILLER_24_47 ();
 sg13g2_fill_1 FILLER_24_49 ();
 sg13g2_fill_2 FILLER_24_73 ();
 sg13g2_fill_1 FILLER_24_75 ();
 sg13g2_fill_2 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_150 ();
 sg13g2_fill_1 FILLER_24_152 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_decap_4 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_234 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_256 ();
 sg13g2_fill_2 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_decap_8 FILLER_24_290 ();
 sg13g2_decap_8 FILLER_24_297 ();
 sg13g2_fill_2 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_24_311 ();
 sg13g2_fill_1 FILLER_24_313 ();
 sg13g2_fill_1 FILLER_24_348 ();
 sg13g2_fill_2 FILLER_24_358 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_4 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_68 ();
 sg13g2_fill_2 FILLER_25_78 ();
 sg13g2_fill_1 FILLER_25_92 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_fill_2 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_fill_2 FILLER_25_127 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_decap_4 FILLER_25_173 ();
 sg13g2_fill_2 FILLER_25_202 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_fill_1 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_fill_1 FILLER_25_278 ();
 sg13g2_fill_2 FILLER_25_287 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_decap_4 FILLER_25_318 ();
 sg13g2_fill_2 FILLER_25_322 ();
 sg13g2_fill_1 FILLER_25_341 ();
 sg13g2_fill_1 FILLER_25_358 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_57 ();
 sg13g2_fill_1 FILLER_26_61 ();
 sg13g2_decap_8 FILLER_26_82 ();
 sg13g2_decap_8 FILLER_26_93 ();
 sg13g2_fill_2 FILLER_26_100 ();
 sg13g2_fill_1 FILLER_26_102 ();
 sg13g2_fill_2 FILLER_26_142 ();
 sg13g2_decap_4 FILLER_26_170 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_decap_8 FILLER_26_220 ();
 sg13g2_decap_8 FILLER_26_227 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_decap_4 FILLER_26_247 ();
 sg13g2_fill_2 FILLER_26_251 ();
 sg13g2_decap_4 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_260 ();
 sg13g2_fill_2 FILLER_26_286 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_304 ();
 sg13g2_decap_4 FILLER_26_349 ();
 sg13g2_fill_2 FILLER_26_358 ();
 sg13g2_fill_2 FILLER_26_385 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_decap_4 FILLER_27_66 ();
 sg13g2_fill_1 FILLER_27_70 ();
 sg13g2_fill_2 FILLER_27_75 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_decap_4 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_148 ();
 sg13g2_decap_4 FILLER_27_195 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_2 FILLER_27_236 ();
 sg13g2_decap_4 FILLER_27_252 ();
 sg13g2_decap_4 FILLER_27_266 ();
 sg13g2_fill_2 FILLER_27_270 ();
 sg13g2_fill_2 FILLER_27_277 ();
 sg13g2_fill_1 FILLER_27_279 ();
 sg13g2_decap_4 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_321 ();
 sg13g2_decap_4 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_330 ();
 sg13g2_fill_1 FILLER_27_336 ();
 sg13g2_fill_1 FILLER_28_26 ();
 sg13g2_fill_2 FILLER_28_32 ();
 sg13g2_fill_2 FILLER_28_39 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_decap_4 FILLER_28_157 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_194 ();
 sg13g2_fill_2 FILLER_28_233 ();
 sg13g2_fill_1 FILLER_28_235 ();
 sg13g2_fill_1 FILLER_28_245 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_337 ();
 sg13g2_fill_2 FILLER_28_371 ();
 sg13g2_fill_1 FILLER_28_373 ();
 sg13g2_fill_1 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_39 ();
 sg13g2_fill_2 FILLER_29_108 ();
 sg13g2_fill_1 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_decap_4 FILLER_29_195 ();
 sg13g2_fill_2 FILLER_29_199 ();
 sg13g2_fill_2 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_236 ();
 sg13g2_fill_2 FILLER_29_301 ();
 sg13g2_fill_2 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_352 ();
 sg13g2_fill_1 FILLER_29_386 ();
 sg13g2_decap_4 FILLER_30_13 ();
 sg13g2_fill_2 FILLER_30_23 ();
 sg13g2_fill_1 FILLER_30_25 ();
 sg13g2_fill_1 FILLER_30_75 ();
 sg13g2_fill_1 FILLER_30_103 ();
 sg13g2_fill_1 FILLER_30_109 ();
 sg13g2_fill_2 FILLER_30_115 ();
 sg13g2_fill_1 FILLER_30_117 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_fill_2 FILLER_30_141 ();
 sg13g2_fill_1 FILLER_30_143 ();
 sg13g2_decap_8 FILLER_30_162 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_176 ();
 sg13g2_fill_1 FILLER_30_181 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_fill_1 FILLER_30_220 ();
 sg13g2_fill_2 FILLER_30_230 ();
 sg13g2_fill_2 FILLER_30_241 ();
 sg13g2_fill_2 FILLER_30_262 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_340 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_15 ();
 sg13g2_fill_1 FILLER_31_17 ();
 sg13g2_fill_1 FILLER_31_23 ();
 sg13g2_fill_2 FILLER_31_43 ();
 sg13g2_fill_1 FILLER_31_45 ();
 sg13g2_fill_2 FILLER_31_50 ();
 sg13g2_fill_2 FILLER_31_64 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_fill_2 FILLER_31_80 ();
 sg13g2_decap_4 FILLER_31_141 ();
 sg13g2_fill_2 FILLER_31_157 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_fill_2 FILLER_31_292 ();
 sg13g2_fill_1 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_decap_8 FILLER_31_317 ();
 sg13g2_fill_2 FILLER_31_345 ();
 sg13g2_decap_4 FILLER_31_360 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_fill_2 FILLER_31_387 ();
 sg13g2_fill_1 FILLER_31_389 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_2 ();
 sg13g2_fill_2 FILLER_32_16 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_fill_1 FILLER_32_37 ();
 sg13g2_fill_1 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_128 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_fill_1 FILLER_32_147 ();
 sg13g2_fill_2 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_fill_1 FILLER_32_269 ();
 sg13g2_fill_2 FILLER_32_284 ();
 sg13g2_fill_2 FILLER_32_309 ();
 sg13g2_fill_2 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_346 ();
 sg13g2_fill_2 FILLER_32_358 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_13 ();
 sg13g2_fill_2 FILLER_33_46 ();
 sg13g2_fill_2 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_104 ();
 sg13g2_fill_2 FILLER_33_110 ();
 sg13g2_decap_4 FILLER_33_145 ();
 sg13g2_fill_2 FILLER_33_149 ();
 sg13g2_fill_1 FILLER_33_200 ();
 sg13g2_fill_2 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_362 ();
 sg13g2_fill_2 FILLER_33_366 ();
 sg13g2_fill_1 FILLER_33_384 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_22 ();
 sg13g2_fill_2 FILLER_34_36 ();
 sg13g2_fill_2 FILLER_34_63 ();
 sg13g2_fill_2 FILLER_34_109 ();
 sg13g2_fill_1 FILLER_34_111 ();
 sg13g2_decap_8 FILLER_34_115 ();
 sg13g2_fill_1 FILLER_34_122 ();
 sg13g2_fill_1 FILLER_34_140 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_decap_4 FILLER_34_176 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_fill_2 FILLER_34_195 ();
 sg13g2_fill_1 FILLER_34_197 ();
 sg13g2_decap_8 FILLER_34_202 ();
 sg13g2_decap_4 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_302 ();
 sg13g2_fill_2 FILLER_34_308 ();
 sg13g2_fill_1 FILLER_34_329 ();
 sg13g2_decap_4 FILLER_34_343 ();
 sg13g2_fill_1 FILLER_34_347 ();
 sg13g2_fill_2 FILLER_34_361 ();
 sg13g2_fill_2 FILLER_34_378 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_36 ();
 sg13g2_fill_2 FILLER_35_141 ();
 sg13g2_fill_1 FILLER_35_143 ();
 sg13g2_fill_2 FILLER_35_155 ();
 sg13g2_fill_2 FILLER_35_162 ();
 sg13g2_decap_4 FILLER_35_179 ();
 sg13g2_decap_4 FILLER_35_193 ();
 sg13g2_fill_2 FILLER_35_197 ();
 sg13g2_decap_4 FILLER_35_225 ();
 sg13g2_fill_2 FILLER_35_292 ();
 sg13g2_fill_2 FILLER_35_303 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_fill_2 FILLER_35_358 ();
 sg13g2_fill_1 FILLER_35_368 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_15 ();
 sg13g2_decap_4 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_decap_8 FILLER_36_177 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_fill_2 FILLER_36_193 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_fill_1 FILLER_36_210 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_fill_2 FILLER_36_379 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_fill_1 FILLER_37_71 ();
 sg13g2_fill_1 FILLER_37_81 ();
 sg13g2_fill_1 FILLER_37_86 ();
 sg13g2_fill_1 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_117 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_141 ();
 sg13g2_decap_4 FILLER_37_148 ();
 sg13g2_fill_2 FILLER_37_165 ();
 sg13g2_fill_2 FILLER_37_172 ();
 sg13g2_fill_2 FILLER_37_192 ();
 sg13g2_fill_1 FILLER_37_194 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_335 ();
 sg13g2_fill_1 FILLER_37_350 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_11 ();
 sg13g2_fill_2 FILLER_38_43 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_137 ();
 sg13g2_fill_1 FILLER_38_139 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_fill_1 FILLER_38_194 ();
 sg13g2_fill_1 FILLER_38_280 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_399 ();
 assign uio_oe[0] = net125;
 assign uio_oe[1] = net126;
 assign uio_oe[2] = net127;
 assign uio_oe[3] = net128;
 assign uio_oe[4] = net129;
 assign uio_oe[5] = net130;
 assign uio_oe[6] = net131;
 assign uio_oe[7] = net132;
endmodule
