module tt_um_rte_eink_driver (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clk_regs;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire csb;
 wire \data_out[0] ;
 wire \data_out[1] ;
 wire \data_out[2] ;
 wire \data_out[3] ;
 wire \data_out[4] ;
 wire \data_out[5] ;
 wire \data_out[6] ;
 wire \data_out[7] ;
 wire dcb;
 wire \inbuf[0] ;
 wire \inbuf[1] ;
 wire \inbuf[2] ;
 wire \inbuf[3] ;
 wire \inbuf[4] ;
 wire \inbuf[5] ;
 wire \inbuf[6] ;
 wire \inbuf[7] ;
 wire \inval[0] ;
 wire \inval[1] ;
 wire \inval[2] ;
 wire \inval[3] ;
 wire \inval[4] ;
 wire \inval[5] ;
 wire \inval[6] ;
 wire \inval[7] ;
 wire maskcsb;
 wire mosi;
 wire mosienb;
 wire passthru;
 wire resetb;
 wire sck;
 wire \spi.count[0] ;
 wire \spi.count[1] ;
 wire \spi.count[2] ;
 wire \spi.count[3] ;
 wire \spi.count[4] ;
 wire \spi.count[5] ;
 wire \spi.count[6] ;
 wire \spi.count[7] ;
 wire \spi.d_latched[0] ;
 wire \spi.d_latched[1] ;
 wire \spi.d_latched[2] ;
 wire \spi.d_latched[3] ;
 wire \spi.d_latched[4] ;
 wire \spi.d_latched[5] ;
 wire \spi.d_latched[6] ;
 wire \spi.d_latched[7] ;
 wire \spi.done ;
 wire \spi.hsck ;
 wire \spi.isck ;
 wire \spi.mosi ;
 wire \spi.nbit[0] ;
 wire \spi.nbit[1] ;
 wire \spi.nbit[2] ;
 wire \spi.reg_dat_we ;
 wire \spi.rreg[0] ;
 wire \spi.rreg[1] ;
 wire \spi.rreg[2] ;
 wire \spi.rreg[3] ;
 wire \spi.rreg[4] ;
 wire \spi.rreg[5] ;
 wire \spi.rreg[6] ;
 wire \spi.rreg[7] ;
 wire \spi.state[0] ;
 wire \spi.state[1] ;
 wire \spi.state[2] ;
 wire \spi.state[3] ;
 wire \spi.stream ;
 wire \spi.treg[0] ;
 wire \spi.treg[1] ;
 wire \spi.treg[2] ;
 wire \spi.treg[3] ;
 wire \spi.treg[4] ;
 wire \spi.treg[5] ;
 wire \spi.treg[6] ;
 wire \spi.treg[7] ;
 wire \spi.w_latched ;
 wire sramcsb;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire stream;
 wire \timer[0] ;
 wire \timer[1] ;
 wire \timer[2] ;
 wire \timer[3] ;
 wire net23;
 wire net12;
 wire net24;
 wire net25;
 wire net26;
 wire net13;
 wire net27;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;

 sg13g2_inv_1 _0719_ (.Y(_0128_),
    .A(net56));
 sg13g2_inv_1 _0720_ (.Y(_0129_),
    .A(net92));
 sg13g2_inv_1 _0721_ (.Y(_0130_),
    .A(net88));
 sg13g2_inv_1 _0722_ (.Y(_0131_),
    .A(_0036_));
 sg13g2_inv_1 _0723_ (.Y(_0132_),
    .A(net59));
 sg13g2_inv_1 _0724_ (.Y(_0133_),
    .A(net197));
 sg13g2_inv_1 _0725_ (.Y(_0134_),
    .A(\spi.state[0] ));
 sg13g2_inv_1 _0726_ (.Y(_0135_),
    .A(\spi.state[1] ));
 sg13g2_inv_1 _0727_ (.Y(_0136_),
    .A(net217));
 sg13g2_inv_2 _0728_ (.Y(_0137_),
    .A(net213));
 sg13g2_inv_2 _0729_ (.Y(_0138_),
    .A(net105));
 sg13g2_inv_1 _0730_ (.Y(_0139_),
    .A(net212));
 sg13g2_inv_1 _0731_ (.Y(_0140_),
    .A(net206));
 sg13g2_inv_1 _0732_ (.Y(_0141_),
    .A(\counter[13] ));
 sg13g2_inv_1 _0733_ (.Y(_0142_),
    .A(net74));
 sg13g2_inv_2 _0734_ (.Y(_0143_),
    .A(\spi.done ));
 sg13g2_inv_1 _0735_ (.Y(_0144_),
    .A(\inbuf[5] ));
 sg13g2_inv_1 _0736_ (.Y(_0145_),
    .A(\inbuf[6] ));
 sg13g2_inv_1 _0737_ (.Y(_0146_),
    .A(\inbuf[7] ));
 sg13g2_inv_1 _0738_ (.Y(_0147_),
    .A(\inbuf[1] ));
 sg13g2_inv_1 _0739_ (.Y(_0148_),
    .A(\inbuf[3] ));
 sg13g2_inv_1 _0740_ (.Y(_0149_),
    .A(\inval[1] ));
 sg13g2_inv_1 _0741_ (.Y(_0150_),
    .A(\inval[3] ));
 sg13g2_inv_1 _0742_ (.Y(_0151_),
    .A(\inval[5] ));
 sg13g2_inv_1 _0743_ (.Y(_0152_),
    .A(\inval[6] ));
 sg13g2_inv_1 _0744_ (.Y(_0153_),
    .A(\inval[7] ));
 sg13g2_inv_1 _0745_ (.Y(_0154_),
    .A(resetb));
 sg13g2_inv_1 _0746_ (.Y(_0155_),
    .A(net85));
 sg13g2_inv_1 _0747_ (.Y(_0156_),
    .A(_0016_));
 sg13g2_inv_1 _0748_ (.Y(_0157_),
    .A(_0020_));
 sg13g2_inv_2 _0749_ (.Y(uio_oe[1]),
    .A(mosienb));
 sg13g2_inv_1 _1332__2 (.Y(net28),
    .A(clknet_1_0__leaf_clk));
 sg13g2_nor2_2 _0751_ (.A(\spi.state[1] ),
    .B(\spi.state[2] ),
    .Y(_0158_));
 sg13g2_a21oi_1 _0752_ (.A1(net197),
    .A2(_0143_),
    .Y(_0159_),
    .B1(_0014_));
 sg13g2_nand2_2 _0753_ (.Y(_0160_),
    .A(_0158_),
    .B(_0159_));
 sg13g2_nor2_1 _0754_ (.A(\data_out[7] ),
    .B(net191),
    .Y(_0161_));
 sg13g2_a21oi_1 _0755_ (.A1(_0128_),
    .A2(_0160_),
    .Y(_0127_),
    .B1(_0161_));
 sg13g2_mux2_1 _0756_ (.A0(\data_out[6] ),
    .A1(net87),
    .S(_0160_),
    .X(_0126_));
 sg13g2_mux2_1 _0757_ (.A0(\data_out[5] ),
    .A1(net84),
    .S(net191),
    .X(_0125_));
 sg13g2_mux2_1 _0758_ (.A0(\data_out[4] ),
    .A1(net76),
    .S(net191),
    .X(_0124_));
 sg13g2_mux2_1 _0759_ (.A0(\data_out[3] ),
    .A1(net83),
    .S(_0160_),
    .X(_0123_));
 sg13g2_mux2_1 _0760_ (.A0(\data_out[2] ),
    .A1(net82),
    .S(net191),
    .X(_0122_));
 sg13g2_nand2_1 _0761_ (.Y(_0162_),
    .A(net52),
    .B(net191));
 sg13g2_o21ai_1 _0762_ (.B1(_0162_),
    .Y(_0121_),
    .A1(_0129_),
    .A2(net191));
 sg13g2_nand2_1 _0763_ (.Y(_0163_),
    .A(net64),
    .B(net191));
 sg13g2_o21ai_1 _0764_ (.B1(_0163_),
    .Y(_0120_),
    .A1(_0130_),
    .A2(net191));
 sg13g2_o21ai_1 _0765_ (.B1(_0158_),
    .Y(_0164_),
    .A1(net197),
    .A2(\spi.reg_dat_we ));
 sg13g2_o21ai_1 _0766_ (.B1(_0164_),
    .Y(_0056_),
    .A1(_0133_),
    .A2(_0014_));
 sg13g2_a21oi_1 _0767_ (.A1(_0133_),
    .A2(\spi.state[0] ),
    .Y(_0045_),
    .B1(\spi.state[3] ));
 sg13g2_nand2_1 _0768_ (.Y(_0165_),
    .A(\spi.nbit[0] ),
    .B(\spi.nbit[1] ));
 sg13g2_o21ai_1 _0769_ (.B1(\spi.state[1] ),
    .Y(_0166_),
    .A1(_0013_),
    .A2(_0165_));
 sg13g2_nand2_1 _0770_ (.Y(_0167_),
    .A(net196),
    .B(\spi.state[0] ));
 sg13g2_nand2_1 _0771_ (.Y(_0001_),
    .A(_0166_),
    .B(_0167_));
 sg13g2_nor4_1 _0772_ (.A(\spi.count[5] ),
    .B(\spi.count[4] ),
    .C(net61),
    .D(net77),
    .Y(_0168_));
 sg13g2_nand3b_1 _0773_ (.B(_0168_),
    .C(net96),
    .Y(_0169_),
    .A_N(\spi.count[2] ));
 sg13g2_nor3_2 _0774_ (.A(net89),
    .B(net85),
    .C(_0169_),
    .Y(_0170_));
 sg13g2_nor2_1 _0775_ (.A(net89),
    .B(_0170_),
    .Y(_0002_));
 sg13g2_xnor2_1 _0776_ (.Y(_0171_),
    .A(net89),
    .B(net96));
 sg13g2_nor2_1 _0777_ (.A(_0170_),
    .B(_0171_),
    .Y(_0003_));
 sg13g2_nand3_1 _0778_ (.B(net96),
    .C(net107),
    .A(net89),
    .Y(_0172_));
 sg13g2_a21o_1 _0779_ (.A2(net96),
    .A1(net89),
    .B1(net107),
    .X(_0173_));
 sg13g2_and2_1 _0780_ (.A(_0172_),
    .B(_0173_),
    .X(_0004_));
 sg13g2_nor2_2 _0781_ (.A(_0155_),
    .B(_0172_),
    .Y(_0174_));
 sg13g2_xnor2_1 _0782_ (.Y(_0005_),
    .A(net85),
    .B(_0172_));
 sg13g2_xor2_1 _0783_ (.B(_0174_),
    .A(net94),
    .X(_0006_));
 sg13g2_nand3_1 _0784_ (.B(net94),
    .C(_0174_),
    .A(net110),
    .Y(_0175_));
 sg13g2_a21o_1 _0785_ (.A2(_0174_),
    .A1(net94),
    .B1(net110),
    .X(_0176_));
 sg13g2_and2_1 _0786_ (.A(_0175_),
    .B(_0176_),
    .X(_0007_));
 sg13g2_nand4_1 _0787_ (.B(\spi.count[4] ),
    .C(\spi.count[6] ),
    .A(\spi.count[5] ),
    .Y(_0177_),
    .D(_0174_));
 sg13g2_xnor2_1 _0788_ (.Y(_0008_),
    .A(net77),
    .B(_0175_));
 sg13g2_xnor2_1 _0789_ (.Y(_0009_),
    .A(net61),
    .B(_0177_));
 sg13g2_nor3_1 _0790_ (.A(\spi.state[0] ),
    .B(\spi.state[3] ),
    .C(_0156_),
    .Y(_0010_));
 sg13g2_mux2_1 _0791_ (.A0(\spi.mosi ),
    .A1(net2),
    .S(passthru),
    .X(mosi));
 sg13g2_mux2_1 _0792_ (.A0(\spi.isck ),
    .A1(net1),
    .S(passthru),
    .X(sck));
 sg13g2_nor3_1 _0793_ (.A(_0135_),
    .B(_0013_),
    .C(_0165_),
    .Y(_0000_));
 sg13g2_or2_1 _0794_ (.X(csb),
    .B(maskcsb),
    .A(mosienb));
 sg13g2_nor2_1 _0795_ (.A(net196),
    .B(_0024_),
    .Y(_0178_));
 sg13g2_a21oi_1 _0796_ (.A1(\spi.d_latched[0] ),
    .A2(net196),
    .Y(_0055_),
    .B1(_0178_));
 sg13g2_nor2_2 _0797_ (.A(\counter[5] ),
    .B(\counter[4] ),
    .Y(_0179_));
 sg13g2_or2_2 _0798_ (.X(_0180_),
    .B(\counter[4] ),
    .A(\counter[5] ));
 sg13g2_nand2_2 _0799_ (.Y(_0181_),
    .A(\counter[3] ),
    .B(net215));
 sg13g2_nand2b_2 _0800_ (.Y(_0182_),
    .B(net216),
    .A_N(net217));
 sg13g2_or2_1 _0801_ (.X(_0183_),
    .B(_0182_),
    .A(_0181_));
 sg13g2_nor2_1 _0802_ (.A(net199),
    .B(_0183_),
    .Y(_0184_));
 sg13g2_nand2b_2 _0803_ (.Y(_0185_),
    .B(net215),
    .A_N(net213));
 sg13g2_nor2_2 _0804_ (.A(net216),
    .B(net217),
    .Y(_0186_));
 sg13g2_nor2b_2 _0805_ (.A(\counter[5] ),
    .B_N(\counter[4] ),
    .Y(_0187_));
 sg13g2_nand2b_2 _0806_ (.Y(_0188_),
    .B(\counter[4] ),
    .A_N(\counter[5] ));
 sg13g2_and2_1 _0807_ (.A(_0186_),
    .B(_0187_),
    .X(_0189_));
 sg13g2_and2_1 _0808_ (.A(net214),
    .B(_0186_),
    .X(_0190_));
 sg13g2_nor2_1 _0809_ (.A(_0185_),
    .B(_0188_),
    .Y(_0191_));
 sg13g2_a21oi_1 _0810_ (.A1(_0186_),
    .A2(_0191_),
    .Y(_0192_),
    .B1(_0184_));
 sg13g2_nor2_2 _0811_ (.A(net213),
    .B(net215),
    .Y(_0193_));
 sg13g2_nand2b_2 _0812_ (.Y(_0194_),
    .B(net218),
    .A_N(\counter[1] ));
 sg13g2_nand3b_1 _0813_ (.B(net218),
    .C(_0193_),
    .Y(_0195_),
    .A_N(net216));
 sg13g2_o21ai_1 _0814_ (.B1(_0192_),
    .Y(_0196_),
    .A1(_0188_),
    .A2(_0195_));
 sg13g2_nor2_1 _0815_ (.A(net216),
    .B(_0185_),
    .Y(_0197_));
 sg13g2_nor3_2 _0816_ (.A(net216),
    .B(_0180_),
    .C(_0185_),
    .Y(_0198_));
 sg13g2_and2_2 _0817_ (.A(_0136_),
    .B(_0198_),
    .X(_0199_));
 sg13g2_nor2_1 _0818_ (.A(_0137_),
    .B(net214),
    .Y(_0200_));
 sg13g2_nand2b_2 _0819_ (.Y(_0201_),
    .B(net213),
    .A_N(net215));
 sg13g2_nor2_2 _0820_ (.A(_0194_),
    .B(_0201_),
    .Y(_0202_));
 sg13g2_nor4_2 _0821_ (.A(net218),
    .B(net213),
    .C(net214),
    .Y(_0203_),
    .D(net199));
 sg13g2_nor2_1 _0822_ (.A(_0181_),
    .B(_0194_),
    .Y(_0204_));
 sg13g2_nor3_2 _0823_ (.A(_0181_),
    .B(_0188_),
    .C(_0194_),
    .Y(_0205_));
 sg13g2_nor3_1 _0824_ (.A(_0137_),
    .B(_0188_),
    .C(_0194_),
    .Y(_0206_));
 sg13g2_nor4_1 _0825_ (.A(_0196_),
    .B(_0199_),
    .C(_0203_),
    .D(_0206_),
    .Y(_0207_));
 sg13g2_inv_1 _0826_ (.Y(_0208_),
    .A(_0207_));
 sg13g2_nor4_2 _0827_ (.A(net216),
    .B(net218),
    .C(_0137_),
    .Y(_0209_),
    .D(net199));
 sg13g2_nor2_1 _0828_ (.A(net213),
    .B(_0182_),
    .Y(_0210_));
 sg13g2_nor3_1 _0829_ (.A(_0180_),
    .B(_0182_),
    .C(_0185_),
    .Y(_0211_));
 sg13g2_nor3_1 _0830_ (.A(_0208_),
    .B(_0209_),
    .C(_0211_),
    .Y(_0212_));
 sg13g2_and2_1 _0831_ (.A(net216),
    .B(net217),
    .X(_0213_));
 sg13g2_nand2_2 _0832_ (.Y(_0214_),
    .A(\counter[1] ),
    .B(net217));
 sg13g2_nor2_1 _0833_ (.A(_0201_),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_nor3_2 _0834_ (.A(net199),
    .B(_0201_),
    .C(_0214_),
    .Y(_0216_));
 sg13g2_a221oi_1 _0835_ (.B2(_0179_),
    .C1(_0216_),
    .B1(_0204_),
    .A1(_0185_),
    .Y(_0217_),
    .A2(_0189_));
 sg13g2_nand2_2 _0836_ (.Y(_0218_),
    .A(_0193_),
    .B(_0213_));
 sg13g2_nor2_2 _0837_ (.A(\counter[5] ),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_nand2_2 _0838_ (.Y(_0220_),
    .A(net224),
    .B(net226));
 sg13g2_and3_1 _0839_ (.X(_0221_),
    .A(net224),
    .B(net226),
    .C(_0012_));
 sg13g2_nor2b_2 _0840_ (.A(net223),
    .B_N(\state[3] ),
    .Y(_0222_));
 sg13g2_nand2b_1 _0841_ (.Y(_0223_),
    .B(\state[3] ),
    .A_N(net223));
 sg13g2_nand2_2 _0842_ (.Y(_0224_),
    .A(_0012_),
    .B(_0222_));
 sg13g2_nor2_2 _0843_ (.A(_0220_),
    .B(_0224_),
    .Y(_0225_));
 sg13g2_nor2_2 _0844_ (.A(_0180_),
    .B(_0218_),
    .Y(_0226_));
 sg13g2_nor2_2 _0845_ (.A(net199),
    .B(_0195_),
    .Y(_0227_));
 sg13g2_nor2_1 _0846_ (.A(_0226_),
    .B(_0227_),
    .Y(_0228_));
 sg13g2_nor3_2 _0847_ (.A(_0136_),
    .B(net199),
    .C(_0185_),
    .Y(_0229_));
 sg13g2_nand3b_1 _0848_ (.B(_0225_),
    .C(_0217_),
    .Y(_0230_),
    .A_N(_0229_));
 sg13g2_nor3_1 _0849_ (.A(_0219_),
    .B(_0227_),
    .C(_0230_),
    .Y(_0231_));
 sg13g2_nand2_1 _0850_ (.Y(_0232_),
    .A(_0212_),
    .B(_0231_));
 sg13g2_nor2b_1 _0851_ (.A(net224),
    .B_N(net226),
    .Y(_0233_));
 sg13g2_nand2b_2 _0852_ (.Y(_0234_),
    .B(\state[0] ),
    .A_N(net225));
 sg13g2_nor2b_2 _0853_ (.A(net222),
    .B_N(\state[2] ),
    .Y(_0235_));
 sg13g2_nand2b_2 _0854_ (.Y(_0236_),
    .B(\state[2] ),
    .A_N(net222));
 sg13g2_nand2_2 _0855_ (.Y(_0237_),
    .A(net221),
    .B(_0235_));
 sg13g2_nor2_2 _0856_ (.A(_0234_),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_nand3_1 _0857_ (.B(_0233_),
    .C(_0235_),
    .A(net221),
    .Y(_0239_));
 sg13g2_nor2_1 _0858_ (.A(_0136_),
    .B(net214),
    .Y(_0240_));
 sg13g2_nor3_1 _0859_ (.A(_0190_),
    .B(_0239_),
    .C(_0240_),
    .Y(_0241_));
 sg13g2_a21oi_1 _0860_ (.A1(_0136_),
    .A2(_0015_),
    .Y(_0242_),
    .B1(_0190_));
 sg13g2_nand3_1 _0861_ (.B(_0241_),
    .C(_0242_),
    .A(\spi.done ),
    .Y(_0243_));
 sg13g2_nor2_2 _0862_ (.A(net222),
    .B(net223),
    .Y(_0244_));
 sg13g2_or2_1 _0863_ (.X(_0245_),
    .B(net223),
    .A(net222));
 sg13g2_nand2_2 _0864_ (.Y(_0246_),
    .A(_0221_),
    .B(_0244_));
 sg13g2_nor2b_1 _0865_ (.A(net226),
    .B_N(net224),
    .Y(_0247_));
 sg13g2_nand2b_2 _0866_ (.Y(_0248_),
    .B(net224),
    .A_N(net226));
 sg13g2_nand2_2 _0867_ (.Y(_0249_),
    .A(net221),
    .B(_0244_));
 sg13g2_nand3_1 _0868_ (.B(_0244_),
    .C(_0247_),
    .A(net220),
    .Y(_0250_));
 sg13g2_nor2_2 _0869_ (.A(net224),
    .B(net226),
    .Y(_0251_));
 sg13g2_nand3_1 _0870_ (.B(_0222_),
    .C(_0251_),
    .A(_0012_),
    .Y(_0252_));
 sg13g2_nand2_1 _0871_ (.Y(_0253_),
    .A(_0250_),
    .B(_0252_));
 sg13g2_and2_1 _0872_ (.A(_0246_),
    .B(_0252_),
    .X(_0254_));
 sg13g2_nand2_1 _0873_ (.Y(_0255_),
    .A(_0250_),
    .B(_0254_));
 sg13g2_nand2_2 _0874_ (.Y(_0256_),
    .A(net222),
    .B(net223));
 sg13g2_nor3_1 _0875_ (.A(net220),
    .B(_0234_),
    .C(_0256_),
    .Y(_0257_));
 sg13g2_nor2_1 _0876_ (.A(_0255_),
    .B(_0257_),
    .Y(_0258_));
 sg13g2_nor2_1 _0877_ (.A(_0225_),
    .B(_0238_),
    .Y(_0259_));
 sg13g2_o21ai_1 _0878_ (.B1(_0258_),
    .Y(_0260_),
    .A1(_0143_),
    .A2(_0259_));
 sg13g2_nand3_1 _0879_ (.B(_0243_),
    .C(_0260_),
    .A(_0232_),
    .Y(_0261_));
 sg13g2_nor3_1 _0880_ (.A(_0212_),
    .B(_0238_),
    .C(_0255_),
    .Y(_0262_));
 sg13g2_and2_2 _0881_ (.A(_0012_),
    .B(_0233_),
    .X(_0263_));
 sg13g2_nand2_1 _0882_ (.Y(_0264_),
    .A(_0012_),
    .B(_0233_));
 sg13g2_nand2b_2 _0883_ (.Y(_0265_),
    .B(_0263_),
    .A_N(_0256_));
 sg13g2_o21ai_1 _0884_ (.B1(_0265_),
    .Y(_0266_),
    .A1(_0239_),
    .A2(_0242_));
 sg13g2_nor2_1 _0885_ (.A(_0262_),
    .B(_0266_),
    .Y(_0267_));
 sg13g2_mux2_1 _0886_ (.A0(_0267_),
    .A1(net70),
    .S(_0261_),
    .X(_0057_));
 sg13g2_nand2_2 _0887_ (.Y(_0268_),
    .A(_0244_),
    .B(_0263_));
 sg13g2_nand2_2 _0888_ (.Y(_0269_),
    .A(_0012_),
    .B(_0247_));
 sg13g2_nor2_1 _0889_ (.A(\state[2] ),
    .B(_0269_),
    .Y(_0270_));
 sg13g2_nor2_1 _0890_ (.A(_0245_),
    .B(_0269_),
    .Y(_0271_));
 sg13g2_nand2_1 _0891_ (.Y(_0272_),
    .A(net65),
    .B(net79));
 sg13g2_nand4_1 _0892_ (.B(\timer[0] ),
    .C(\timer[2] ),
    .A(\timer[1] ),
    .Y(_0273_),
    .D(\timer[3] ));
 sg13g2_nor2_2 _0893_ (.A(_0181_),
    .B(_0214_),
    .Y(_0274_));
 sg13g2_nand4_1 _0894_ (.B(\counter[4] ),
    .C(\counter[6] ),
    .A(\counter[5] ),
    .Y(_0275_),
    .D(_0274_));
 sg13g2_nand2_1 _0895_ (.Y(_0276_),
    .A(net212),
    .B(net211));
 sg13g2_nand4_1 _0896_ (.B(net210),
    .C(\counter[9] ),
    .A(net212),
    .Y(_0277_),
    .D(net208));
 sg13g2_nor2_2 _0897_ (.A(_0275_),
    .B(_0277_),
    .Y(_0278_));
 sg13g2_nand3_1 _0898_ (.B(net74),
    .C(_0278_),
    .A(net207),
    .Y(_0279_));
 sg13g2_nor2_1 _0899_ (.A(_0141_),
    .B(_0279_),
    .Y(_0280_));
 sg13g2_nand3b_1 _0900_ (.B(_0280_),
    .C(\counter[14] ),
    .Y(_0281_),
    .A_N(\counter[15] ));
 sg13g2_nor4_1 _0901_ (.A(_0245_),
    .B(_0269_),
    .C(_0273_),
    .D(_0281_),
    .Y(_0282_));
 sg13g2_nand2_1 _0902_ (.Y(_0283_),
    .A(net72),
    .B(_0280_));
 sg13g2_nor2_1 _0903_ (.A(\counter[15] ),
    .B(_0283_),
    .Y(_0284_));
 sg13g2_o21ai_1 _0904_ (.B1(_0268_),
    .Y(_0058_),
    .A1(_0132_),
    .A2(_0282_));
 sg13g2_nand3_1 _0905_ (.B(_0235_),
    .C(_0251_),
    .A(net103),
    .Y(_0285_));
 sg13g2_and2_2 _0906_ (.A(net220),
    .B(_0251_),
    .X(_0286_));
 sg13g2_nand2_1 _0907_ (.Y(_0287_),
    .A(_0235_),
    .B(_0286_));
 sg13g2_nand4_1 _0908_ (.B(net226),
    .C(net220),
    .A(net224),
    .Y(_0288_),
    .D(_0222_));
 sg13g2_and3_1 _0909_ (.X(_0289_),
    .A(net222),
    .B(net223),
    .C(_0221_));
 sg13g2_nand2_1 _0910_ (.Y(_0290_),
    .A(_0285_),
    .B(_0288_));
 sg13g2_o21ai_1 _0911_ (.B1(_0287_),
    .Y(_0291_),
    .A1(_0223_),
    .A2(_0269_));
 sg13g2_nor3_1 _0912_ (.A(_0289_),
    .B(_0290_),
    .C(_0291_),
    .Y(_0292_));
 sg13g2_nand2_1 _0913_ (.Y(_0293_),
    .A(net91),
    .B(_0292_));
 sg13g2_nand2b_1 _0914_ (.Y(_0294_),
    .B(\spi.done ),
    .A_N(_0292_));
 sg13g2_nor2_2 _0915_ (.A(_0236_),
    .B(_0264_),
    .Y(_0295_));
 sg13g2_nand2_1 _0916_ (.Y(_0296_),
    .A(_0244_),
    .B(_0286_));
 sg13g2_nor2b_1 _0917_ (.A(_0256_),
    .B_N(_0286_),
    .Y(_0297_));
 sg13g2_nand2b_1 _0918_ (.Y(_0298_),
    .B(_0286_),
    .A_N(_0256_));
 sg13g2_and3_1 _0919_ (.X(_0299_),
    .A(_0259_),
    .B(_0296_),
    .C(_0298_));
 sg13g2_nand3_1 _0920_ (.B(_0296_),
    .C(_0298_),
    .A(_0259_),
    .Y(_0300_));
 sg13g2_a221oi_1 _0921_ (.B2(_0294_),
    .C1(_0300_),
    .B1(_0293_),
    .A1(_0235_),
    .Y(_0059_),
    .A2(_0263_));
 sg13g2_o21ai_1 _0922_ (.B1(_0143_),
    .Y(_0301_),
    .A1(_0295_),
    .A2(_0300_));
 sg13g2_nor2_1 _0923_ (.A(_0234_),
    .B(_0249_),
    .Y(_0302_));
 sg13g2_nor2_2 _0924_ (.A(_0237_),
    .B(_0248_),
    .Y(_0303_));
 sg13g2_nor3_1 _0925_ (.A(net220),
    .B(_0220_),
    .C(_0223_),
    .Y(_0304_));
 sg13g2_o21ai_1 _0926_ (.B1(_0239_),
    .Y(_0305_),
    .A1(_0236_),
    .A2(_0264_));
 sg13g2_nor4_1 _0927_ (.A(_0302_),
    .B(_0303_),
    .C(_0304_),
    .D(_0305_),
    .Y(_0306_));
 sg13g2_nor3_1 _0928_ (.A(_0231_),
    .B(_0241_),
    .C(_0306_),
    .Y(_0307_));
 sg13g2_nand2_1 _0929_ (.Y(_0308_),
    .A(_0301_),
    .B(_0307_));
 sg13g2_nand2_1 _0930_ (.Y(_0309_),
    .A(net50),
    .B(_0308_));
 sg13g2_nand3b_1 _0931_ (.B(_0222_),
    .C(_0247_),
    .Y(_0310_),
    .A_N(net221));
 sg13g2_nor2_2 _0932_ (.A(_0220_),
    .B(_0249_),
    .Y(_0311_));
 sg13g2_or2_2 _0933_ (.X(_0312_),
    .B(_0249_),
    .A(_0220_));
 sg13g2_nand4_1 _0934_ (.B(_0309_),
    .C(_0310_),
    .A(_0285_),
    .Y(_0060_),
    .D(_0312_));
 sg13g2_nor2_2 _0935_ (.A(_0256_),
    .B(_0269_),
    .Y(_0313_));
 sg13g2_or2_1 _0936_ (.X(_0314_),
    .B(\inval[3] ),
    .A(\inval[2] ));
 sg13g2_nand2_1 _0937_ (.Y(_0315_),
    .A(\inval[2] ),
    .B(_0019_));
 sg13g2_nand3b_1 _0938_ (.B(\inval[3] ),
    .C(_0018_),
    .Y(_0316_),
    .A_N(\inval[2] ));
 sg13g2_nand3_1 _0939_ (.B(_0315_),
    .C(_0316_),
    .A(_0022_),
    .Y(_0317_));
 sg13g2_o21ai_1 _0940_ (.B1(net204),
    .Y(_0318_),
    .A1(net219),
    .A2(_0138_));
 sg13g2_a21o_2 _0941_ (.A2(_0138_),
    .A1(net219),
    .B1(_0318_),
    .X(_0319_));
 sg13g2_nor2b_1 _0942_ (.A(\counter[10] ),
    .B_N(\counter[9] ),
    .Y(_0320_));
 sg13g2_nand3b_1 _0943_ (.B(net206),
    .C(net209),
    .Y(_0321_),
    .A_N(net208));
 sg13g2_nand2b_1 _0944_ (.Y(_0322_),
    .B(net212),
    .A_N(net210));
 sg13g2_nor2_1 _0945_ (.A(_0321_),
    .B(_0322_),
    .Y(_0323_));
 sg13g2_nor3_1 _0946_ (.A(net213),
    .B(net214),
    .C(_0182_),
    .Y(_0324_));
 sg13g2_nor2b_1 _0947_ (.A(net209),
    .B_N(net208),
    .Y(_0325_));
 sg13g2_nand2b_1 _0948_ (.Y(_0326_),
    .B(net208),
    .A_N(net209));
 sg13g2_nand4_1 _0949_ (.B(net211),
    .C(_0140_),
    .A(net212),
    .Y(_0327_),
    .D(_0325_));
 sg13g2_o21ai_1 _0950_ (.B1(_0327_),
    .Y(_0328_),
    .A1(_0204_),
    .A2(_0324_));
 sg13g2_nand4_1 _0951_ (.B(net211),
    .C(_0020_),
    .A(net212),
    .Y(_0329_),
    .D(_0325_));
 sg13g2_nor2_1 _0952_ (.A(net206),
    .B(_0020_),
    .Y(_0330_));
 sg13g2_or2_1 _0953_ (.X(_0331_),
    .B(net210),
    .A(\counter[7] ));
 sg13g2_nor2_1 _0954_ (.A(_0330_),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_or3_1 _0955_ (.A(_0326_),
    .B(_0330_),
    .C(_0331_),
    .X(_0333_));
 sg13g2_nand3_1 _0956_ (.B(_0329_),
    .C(_0333_),
    .A(_0202_),
    .Y(_0334_));
 sg13g2_a21oi_1 _0957_ (.A1(_0328_),
    .A2(_0334_),
    .Y(_0335_),
    .B1(_0323_));
 sg13g2_a21o_1 _0958_ (.A2(_0193_),
    .A1(_0186_),
    .B1(_0274_),
    .X(_0336_));
 sg13g2_nor2b_1 _0959_ (.A(net212),
    .B_N(net210),
    .Y(_0337_));
 sg13g2_nand3_1 _0960_ (.B(net208),
    .C(_0020_),
    .A(net209),
    .Y(_0338_));
 sg13g2_nand4_1 _0961_ (.B(net208),
    .C(_0020_),
    .A(net209),
    .Y(_0339_),
    .D(_0337_));
 sg13g2_nor2_2 _0962_ (.A(net209),
    .B(net208),
    .Y(_0340_));
 sg13g2_nand3_1 _0963_ (.B(_0337_),
    .C(_0340_),
    .A(net206),
    .Y(_0341_));
 sg13g2_nand4_1 _0964_ (.B(_0210_),
    .C(_0339_),
    .A(net214),
    .Y(_0342_),
    .D(_0341_));
 sg13g2_nor2_1 _0965_ (.A(_0185_),
    .B(_0214_),
    .Y(_0343_));
 sg13g2_a21oi_1 _0966_ (.A1(_0186_),
    .A2(_0200_),
    .Y(_0344_),
    .B1(_0343_));
 sg13g2_a22oi_1 _0967_ (.Y(_0345_),
    .B1(_0342_),
    .B2(_0344_),
    .A2(_0332_),
    .A1(_0325_));
 sg13g2_nand3_1 _0968_ (.B(_0339_),
    .C(_0341_),
    .A(_0197_),
    .Y(_0346_));
 sg13g2_a21oi_1 _0969_ (.A1(_0321_),
    .A2(_0338_),
    .Y(_0347_),
    .B1(_0331_));
 sg13g2_nor2_1 _0970_ (.A(net218),
    .B(_0201_),
    .Y(_0348_));
 sg13g2_nor2_1 _0971_ (.A(_0182_),
    .B(_0201_),
    .Y(_0349_));
 sg13g2_nand2b_1 _0972_ (.Y(_0350_),
    .B(_0349_),
    .A_N(_0347_));
 sg13g2_nor3_1 _0973_ (.A(net206),
    .B(_0322_),
    .C(_0326_),
    .Y(_0351_));
 sg13g2_nor2_1 _0974_ (.A(_0020_),
    .B(_0276_),
    .Y(_0352_));
 sg13g2_a221oi_1 _0975_ (.B2(_0320_),
    .C1(_0351_),
    .B1(_0352_),
    .A1(_0346_),
    .Y(_0353_),
    .A2(_0350_));
 sg13g2_nor4_1 _0976_ (.A(_0335_),
    .B(_0336_),
    .C(_0345_),
    .D(_0353_),
    .Y(_0354_));
 sg13g2_a21o_1 _0977_ (.A2(_0195_),
    .A1(_0183_),
    .B1(_0347_),
    .X(_0355_));
 sg13g2_or2_1 _0978_ (.X(_0356_),
    .B(_0321_),
    .A(_0276_));
 sg13g2_nand4_1 _0979_ (.B(_0339_),
    .C(_0341_),
    .A(_0215_),
    .Y(_0357_),
    .D(_0356_));
 sg13g2_o21ai_1 _0980_ (.B1(_0355_),
    .Y(_0358_),
    .A1(_0351_),
    .A2(_0357_));
 sg13g2_nand4_1 _0981_ (.B(net211),
    .C(net206),
    .A(net212),
    .Y(_0359_),
    .D(_0340_));
 sg13g2_o21ai_1 _0982_ (.B1(_0359_),
    .Y(_0360_),
    .A1(_0322_),
    .A2(_0338_));
 sg13g2_inv_1 _0983_ (.Y(_0361_),
    .A(_0360_));
 sg13g2_and2_1 _0984_ (.A(_0140_),
    .B(_0277_),
    .X(_0362_));
 sg13g2_nand3b_1 _0985_ (.B(net206),
    .C(_0340_),
    .Y(_0363_),
    .A_N(net210));
 sg13g2_a21oi_1 _0986_ (.A1(_0157_),
    .A2(_0363_),
    .Y(_0364_),
    .B1(_0362_));
 sg13g2_nand2_1 _0987_ (.Y(_0365_),
    .A(net213),
    .B(_0190_));
 sg13g2_o21ai_1 _0988_ (.B1(_0218_),
    .Y(_0366_),
    .A1(_0364_),
    .A2(_0365_));
 sg13g2_o21ai_1 _0989_ (.B1(_0321_),
    .Y(_0367_),
    .A1(net206),
    .A2(_0326_));
 sg13g2_nand2_1 _0990_ (.Y(_0368_),
    .A(_0337_),
    .B(_0367_));
 sg13g2_a22oi_1 _0991_ (.Y(_0369_),
    .B1(_0366_),
    .B2(_0368_),
    .A2(_0361_),
    .A1(_0358_));
 sg13g2_nand3_1 _0992_ (.B(_0341_),
    .C(_0363_),
    .A(_0157_),
    .Y(_0370_));
 sg13g2_nand2_1 _0993_ (.Y(_0371_),
    .A(_0336_),
    .B(_0370_));
 sg13g2_a21oi_1 _0994_ (.A1(_0339_),
    .A2(_0362_),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_a21o_1 _0995_ (.A2(_0369_),
    .A1(_0354_),
    .B1(_0372_),
    .X(_0373_));
 sg13g2_xor2_1 _0996_ (.B(net210),
    .A(net214),
    .X(_0374_));
 sg13g2_a21oi_1 _0997_ (.A1(\inval[6] ),
    .A2(_0374_),
    .Y(_0375_),
    .B1(\inval[5] ));
 sg13g2_o21ai_1 _0998_ (.B1(_0375_),
    .Y(_0376_),
    .A1(\inval[6] ),
    .A2(_0373_));
 sg13g2_nand2_2 _0999_ (.Y(_0377_),
    .A(\spi.done ),
    .B(\inval[5] ));
 sg13g2_or2_1 _1000_ (.X(_0378_),
    .B(_0377_),
    .A(\spi.rreg[0] ));
 sg13g2_a21o_1 _1001_ (.A2(_0378_),
    .A1(_0376_),
    .B1(net204),
    .X(_0379_));
 sg13g2_a21oi_1 _1002_ (.A1(_0319_),
    .A2(_0379_),
    .Y(_0380_),
    .B1(net198));
 sg13g2_o21ai_1 _1003_ (.B1(_0021_),
    .Y(_0381_),
    .A1(_0317_),
    .A2(_0380_));
 sg13g2_nor3_1 _1004_ (.A(net199),
    .B(_0185_),
    .C(_0214_),
    .Y(_0382_));
 sg13g2_or2_1 _1005_ (.X(_0383_),
    .B(_0227_),
    .A(_0211_));
 sg13g2_o21ai_1 _1006_ (.B1(_0187_),
    .Y(_0384_),
    .A1(_0343_),
    .A2(_0349_));
 sg13g2_nand2_1 _1007_ (.Y(_0385_),
    .A(_0179_),
    .B(_0202_));
 sg13g2_o21ai_1 _1008_ (.B1(_0385_),
    .Y(_0386_),
    .A1(net199),
    .A2(_0365_));
 sg13g2_o21ai_1 _1009_ (.B1(_0179_),
    .Y(_0387_),
    .A1(_0274_),
    .A2(_0348_));
 sg13g2_nor2_2 _1010_ (.A(_0224_),
    .B(_0234_),
    .Y(_0388_));
 sg13g2_nand2_2 _1011_ (.Y(_0389_),
    .A(_0222_),
    .B(_0263_));
 sg13g2_nor3_1 _1012_ (.A(_0205_),
    .B(_0386_),
    .C(_0389_),
    .Y(_0390_));
 sg13g2_nand2_1 _1013_ (.Y(_0391_),
    .A(_0387_),
    .B(_0390_));
 sg13g2_a221oi_1 _1014_ (.B2(_0213_),
    .C1(_0210_),
    .B1(_0200_),
    .A1(net217),
    .Y(_0392_),
    .A2(_0197_));
 sg13g2_o21ai_1 _1015_ (.B1(_0217_),
    .Y(_0393_),
    .A1(_0188_),
    .A2(_0392_));
 sg13g2_and2_2 _1016_ (.A(\counter[1] ),
    .B(_0203_),
    .X(_0394_));
 sg13g2_or4_1 _1017_ (.A(_0196_),
    .B(_0198_),
    .C(_0219_),
    .D(_0394_),
    .X(_0395_));
 sg13g2_a21oi_1 _1018_ (.A1(_0187_),
    .A2(_0202_),
    .Y(_0396_),
    .B1(_0382_));
 sg13g2_nand3b_1 _1019_ (.B(_0384_),
    .C(_0396_),
    .Y(_0397_),
    .A_N(_0383_));
 sg13g2_nor4_2 _1020_ (.A(_0391_),
    .B(_0393_),
    .C(_0395_),
    .Y(_0398_),
    .D(_0397_));
 sg13g2_nand2_2 _1021_ (.Y(_0399_),
    .A(net220),
    .B(_0222_));
 sg13g2_nor2_2 _1022_ (.A(_0248_),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_a21oi_1 _1023_ (.A1(_0179_),
    .A2(_0193_),
    .Y(_0401_),
    .B1(_0199_));
 sg13g2_nand2_1 _1024_ (.Y(_0402_),
    .A(_0400_),
    .B(_0401_));
 sg13g2_or4_1 _1025_ (.A(net205),
    .B(\inval[5] ),
    .C(\inval[6] ),
    .D(\inval[7] ),
    .X(_0403_));
 sg13g2_nor4_2 _1026_ (.A(\inval[0] ),
    .B(\inval[1] ),
    .C(_0314_),
    .Y(_0404_),
    .D(_0403_));
 sg13g2_nor2_1 _1027_ (.A(_0199_),
    .B(_0394_),
    .Y(_0405_));
 sg13g2_nand3_1 _1028_ (.B(_0311_),
    .C(_0405_),
    .A(_0228_),
    .Y(_0406_));
 sg13g2_o21ai_1 _1029_ (.B1(_0402_),
    .Y(_0407_),
    .A1(_0203_),
    .A2(_0406_));
 sg13g2_a221oi_1 _1030_ (.B2(net192),
    .C1(_0407_),
    .B1(_0404_),
    .A1(_0207_),
    .Y(_0408_),
    .A2(_0398_));
 sg13g2_nor2_1 _1031_ (.A(_0311_),
    .B(net192),
    .Y(_0409_));
 sg13g2_nand3_1 _1032_ (.B(_0389_),
    .C(_0409_),
    .A(_0246_),
    .Y(_0410_));
 sg13g2_nand2_2 _1033_ (.Y(_0411_),
    .A(_0408_),
    .B(_0410_));
 sg13g2_o21ai_1 _1034_ (.B1(_0408_),
    .Y(_0412_),
    .A1(_0400_),
    .A2(_0410_));
 sg13g2_inv_1 _1035_ (.Y(_0413_),
    .A(_0412_));
 sg13g2_nand3b_1 _1036_ (.B(_0385_),
    .C(_0192_),
    .Y(_0414_),
    .A_N(_0219_));
 sg13g2_o21ai_1 _1037_ (.B1(_0388_),
    .Y(_0415_),
    .A1(_0397_),
    .A2(_0414_));
 sg13g2_a21oi_1 _1038_ (.A1(_0199_),
    .A2(_0311_),
    .Y(_0416_),
    .B1(_0398_));
 sg13g2_nand2_1 _1039_ (.Y(_0417_),
    .A(_0415_),
    .B(_0416_));
 sg13g2_a21o_1 _1040_ (.A2(_0405_),
    .A1(_0228_),
    .B1(_0394_),
    .X(_0418_));
 sg13g2_o21ai_1 _1041_ (.B1(_0411_),
    .Y(_0419_),
    .A1(net187),
    .A2(_0418_));
 sg13g2_a21oi_1 _1042_ (.A1(_0313_),
    .A2(_0381_),
    .Y(_0420_),
    .B1(_0417_));
 sg13g2_a22oi_1 _1043_ (.Y(_0061_),
    .B1(_0419_),
    .B2(_0420_),
    .A2(net187),
    .A1(_0130_));
 sg13g2_or2_1 _1044_ (.X(_0421_),
    .B(_0377_),
    .A(\spi.rreg[1] ));
 sg13g2_a21o_1 _1045_ (.A2(_0421_),
    .A1(_0376_),
    .B1(net204),
    .X(_0422_));
 sg13g2_a21oi_1 _1046_ (.A1(_0319_),
    .A2(_0422_),
    .Y(_0423_),
    .B1(net198));
 sg13g2_o21ai_1 _1047_ (.B1(_0021_),
    .Y(_0424_),
    .A1(_0317_),
    .A2(_0423_));
 sg13g2_nand2_1 _1048_ (.Y(_0425_),
    .A(_0246_),
    .B(_0406_));
 sg13g2_a221oi_1 _1049_ (.B2(\counter[4] ),
    .C1(_0184_),
    .B1(_0219_),
    .A1(net215),
    .Y(_0426_),
    .A2(_0209_));
 sg13g2_nor3_1 _1050_ (.A(_0216_),
    .B(_0229_),
    .C(_0383_),
    .Y(_0427_));
 sg13g2_nand2_1 _1051_ (.Y(_0428_),
    .A(_0426_),
    .B(_0427_));
 sg13g2_a21oi_1 _1052_ (.A1(_0313_),
    .A2(_0424_),
    .Y(_0429_),
    .B1(_0425_));
 sg13g2_a221oi_1 _1053_ (.B2(_0388_),
    .C1(net187),
    .B1(_0428_),
    .A1(_0394_),
    .Y(_0430_),
    .A2(_0411_));
 sg13g2_a22oi_1 _1054_ (.Y(_0062_),
    .B1(_0429_),
    .B2(_0430_),
    .A2(net187),
    .A1(_0129_));
 sg13g2_or2_1 _1055_ (.X(_0431_),
    .B(_0377_),
    .A(\spi.rreg[2] ));
 sg13g2_a21o_1 _1056_ (.A2(_0431_),
    .A1(_0376_),
    .B1(net204),
    .X(_0432_));
 sg13g2_a21oi_1 _1057_ (.A1(_0319_),
    .A2(_0432_),
    .Y(_0433_),
    .B1(net198));
 sg13g2_o21ai_1 _1058_ (.B1(_0021_),
    .Y(_0434_),
    .A1(_0317_),
    .A2(_0433_));
 sg13g2_nor4_1 _1059_ (.A(_0205_),
    .B(_0209_),
    .C(_0382_),
    .D(_0395_),
    .Y(_0435_));
 sg13g2_nor2_1 _1060_ (.A(_0389_),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_a221oi_1 _1061_ (.B2(_0434_),
    .C1(_0436_),
    .B1(net192),
    .A1(_0227_),
    .Y(_0437_),
    .A2(_0311_));
 sg13g2_nand2_1 _1062_ (.Y(_0438_),
    .A(net55),
    .B(_0412_));
 sg13g2_o21ai_1 _1063_ (.B1(_0438_),
    .Y(_0063_),
    .A1(_0411_),
    .A2(_0437_));
 sg13g2_nand2_1 _1064_ (.Y(_0439_),
    .A(net57),
    .B(_0412_));
 sg13g2_or2_1 _1065_ (.X(_0440_),
    .B(_0377_),
    .A(\spi.rreg[3] ));
 sg13g2_a21o_1 _1066_ (.A2(_0440_),
    .A1(_0376_),
    .B1(net204),
    .X(_0441_));
 sg13g2_a21oi_1 _1067_ (.A1(_0319_),
    .A2(_0441_),
    .Y(_0442_),
    .B1(net198));
 sg13g2_o21ai_1 _1068_ (.B1(_0021_),
    .Y(_0443_),
    .A1(_0317_),
    .A2(_0442_));
 sg13g2_nor2_1 _1069_ (.A(_0384_),
    .B(_0389_),
    .Y(_0444_));
 sg13g2_nand3_1 _1070_ (.B(_0405_),
    .C(_0426_),
    .A(_0384_),
    .Y(_0445_));
 sg13g2_a22oi_1 _1071_ (.Y(_0446_),
    .B1(_0445_),
    .B2(_0388_),
    .A2(_0443_),
    .A1(_0313_));
 sg13g2_o21ai_1 _1072_ (.B1(_0439_),
    .Y(_0064_),
    .A1(_0411_),
    .A2(_0446_));
 sg13g2_or2_1 _1073_ (.X(_0447_),
    .B(_0377_),
    .A(\spi.rreg[4] ));
 sg13g2_a21o_1 _1074_ (.A2(_0447_),
    .A1(_0376_),
    .B1(net204),
    .X(_0448_));
 sg13g2_a21oi_1 _1075_ (.A1(_0319_),
    .A2(_0448_),
    .Y(_0449_),
    .B1(net198));
 sg13g2_o21ai_1 _1076_ (.B1(_0021_),
    .Y(_0450_),
    .A1(_0317_),
    .A2(_0449_));
 sg13g2_nor3_1 _1077_ (.A(_0216_),
    .B(_0229_),
    .C(_0394_),
    .Y(_0451_));
 sg13g2_nor2_1 _1078_ (.A(_0389_),
    .B(_0451_),
    .Y(_0452_));
 sg13g2_o21ai_1 _1079_ (.B1(_0246_),
    .Y(_0453_),
    .A1(_0228_),
    .A2(_0312_));
 sg13g2_or4_1 _1080_ (.A(_0398_),
    .B(_0444_),
    .C(_0452_),
    .D(_0453_),
    .X(_0454_));
 sg13g2_a21oi_1 _1081_ (.A1(net192),
    .A2(_0450_),
    .Y(_0455_),
    .B1(_0454_));
 sg13g2_nand2_1 _1082_ (.Y(_0456_),
    .A(net53),
    .B(net187));
 sg13g2_o21ai_1 _1083_ (.B1(_0456_),
    .Y(_0065_),
    .A1(_0411_),
    .A2(_0455_));
 sg13g2_or2_1 _1084_ (.X(_0457_),
    .B(_0377_),
    .A(\spi.rreg[5] ));
 sg13g2_a21o_1 _1085_ (.A2(_0457_),
    .A1(_0376_),
    .B1(net205),
    .X(_0458_));
 sg13g2_a21oi_1 _1086_ (.A1(_0319_),
    .A2(_0458_),
    .Y(_0459_),
    .B1(net198));
 sg13g2_o21ai_1 _1087_ (.B1(_0021_),
    .Y(_0460_),
    .A1(_0317_),
    .A2(_0459_));
 sg13g2_nor4_1 _1088_ (.A(_0198_),
    .B(_0205_),
    .C(_0216_),
    .D(_0394_),
    .Y(_0461_));
 sg13g2_nor3_1 _1089_ (.A(_0199_),
    .B(_0226_),
    .C(_0312_),
    .Y(_0462_));
 sg13g2_nor2_1 _1090_ (.A(_0444_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_o21ai_1 _1091_ (.B1(_0463_),
    .Y(_0464_),
    .A1(_0389_),
    .A2(_0461_));
 sg13g2_a21oi_1 _1092_ (.A1(net192),
    .A2(_0460_),
    .Y(_0465_),
    .B1(_0464_));
 sg13g2_nand2_1 _1093_ (.Y(_0466_),
    .A(net46),
    .B(net187));
 sg13g2_o21ai_1 _1094_ (.B1(_0466_),
    .Y(_0066_),
    .A1(_0411_),
    .A2(_0465_));
 sg13g2_nand2_1 _1095_ (.Y(_0467_),
    .A(net48),
    .B(net187));
 sg13g2_or2_1 _1096_ (.X(_0468_),
    .B(_0377_),
    .A(\spi.rreg[6] ));
 sg13g2_a21o_1 _1097_ (.A2(_0468_),
    .A1(_0376_),
    .B1(net204),
    .X(_0469_));
 sg13g2_a21oi_1 _1098_ (.A1(_0319_),
    .A2(_0469_),
    .Y(_0470_),
    .B1(net198));
 sg13g2_o21ai_1 _1099_ (.B1(_0021_),
    .Y(_0471_),
    .A1(_0317_),
    .A2(_0470_));
 sg13g2_o21ai_1 _1100_ (.B1(_0388_),
    .Y(_0472_),
    .A1(_0196_),
    .A2(_0386_));
 sg13g2_a21oi_1 _1101_ (.A1(_0227_),
    .A2(_0311_),
    .Y(_0473_),
    .B1(_0444_));
 sg13g2_nand3_1 _1102_ (.B(_0472_),
    .C(_0473_),
    .A(_0410_),
    .Y(_0474_));
 sg13g2_a21oi_1 _1103_ (.A1(net192),
    .A2(_0471_),
    .Y(_0475_),
    .B1(_0474_));
 sg13g2_o21ai_1 _1104_ (.B1(_0413_),
    .Y(_0476_),
    .A1(_0227_),
    .A2(_0410_));
 sg13g2_o21ai_1 _1105_ (.B1(_0467_),
    .Y(_0067_),
    .A1(_0475_),
    .A2(_0476_));
 sg13g2_or2_1 _1106_ (.X(_0477_),
    .B(_0377_),
    .A(\spi.rreg[7] ));
 sg13g2_a21o_1 _1107_ (.A2(_0477_),
    .A1(_0376_),
    .B1(net204),
    .X(_0478_));
 sg13g2_a21oi_1 _1108_ (.A1(_0319_),
    .A2(_0478_),
    .Y(_0479_),
    .B1(net198));
 sg13g2_o21ai_1 _1109_ (.B1(_0021_),
    .Y(_0480_),
    .A1(_0317_),
    .A2(_0479_));
 sg13g2_a221oi_1 _1110_ (.B2(_0480_),
    .C1(_0444_),
    .B1(net192),
    .A1(_0227_),
    .Y(_0481_),
    .A2(_0311_));
 sg13g2_nand2_1 _1111_ (.Y(_0482_),
    .A(net58),
    .B(net187));
 sg13g2_o21ai_1 _1112_ (.B1(_0482_),
    .Y(_0068_),
    .A1(_0411_),
    .A2(_0481_));
 sg13g2_nand2_1 _1113_ (.Y(_0483_),
    .A(_0221_),
    .B(_0235_));
 sg13g2_nor2b_2 _1114_ (.A(_0271_),
    .B_N(_0483_),
    .Y(_0484_));
 sg13g2_inv_1 _1115_ (.Y(_0485_),
    .A(_0484_));
 sg13g2_o21ai_1 _1116_ (.B1(_0485_),
    .Y(_0486_),
    .A1(_0273_),
    .A2(_0281_));
 sg13g2_nor4_1 _1117_ (.A(\inbuf[1] ),
    .B(\inbuf[0] ),
    .C(\inbuf[3] ),
    .D(\inbuf[2] ),
    .Y(_0487_));
 sg13g2_nor4_1 _1118_ (.A(\inbuf[4] ),
    .B(\inbuf[5] ),
    .C(\inbuf[6] ),
    .D(\inbuf[7] ),
    .Y(_0488_));
 sg13g2_nand2_1 _1119_ (.Y(_0489_),
    .A(_0487_),
    .B(_0488_));
 sg13g2_xnor2_1 _1120_ (.Y(_0490_),
    .A(\inbuf[4] ),
    .B(net205));
 sg13g2_a22oi_1 _1121_ (.Y(_0491_),
    .B1(_0151_),
    .B2(\inbuf[5] ),
    .A2(\inval[1] ),
    .A1(_0147_));
 sg13g2_xnor2_1 _1122_ (.Y(_0492_),
    .A(\inbuf[2] ),
    .B(\inval[2] ));
 sg13g2_a22oi_1 _1123_ (.Y(_0493_),
    .B1(_0153_),
    .B2(\inbuf[7] ),
    .A2(_0149_),
    .A1(\inbuf[1] ));
 sg13g2_a22oi_1 _1124_ (.Y(_0494_),
    .B1(\inval[7] ),
    .B2(_0146_),
    .A2(\inval[3] ),
    .A1(_0148_));
 sg13g2_xnor2_1 _1125_ (.Y(_0495_),
    .A(\inbuf[0] ),
    .B(\inval[0] ));
 sg13g2_a22oi_1 _1126_ (.Y(_0496_),
    .B1(\inval[6] ),
    .B2(_0145_),
    .A2(_0150_),
    .A1(\inbuf[3] ));
 sg13g2_nand4_1 _1127_ (.B(_0494_),
    .C(_0495_),
    .A(_0490_),
    .Y(_0497_),
    .D(_0496_));
 sg13g2_a22oi_1 _1128_ (.Y(_0498_),
    .B1(_0152_),
    .B2(\inbuf[6] ),
    .A2(\inval[5] ),
    .A1(_0144_));
 sg13g2_nand4_1 _1129_ (.B(_0492_),
    .C(_0493_),
    .A(_0491_),
    .Y(_0499_),
    .D(_0498_));
 sg13g2_o21ai_1 _1130_ (.B1(_0489_),
    .Y(_0500_),
    .A1(_0497_),
    .A2(_0499_));
 sg13g2_nand3_1 _1131_ (.B(_0244_),
    .C(_0251_),
    .A(_0012_),
    .Y(_0501_));
 sg13g2_nand4_1 _1132_ (.B(\inbuf[5] ),
    .C(\inbuf[6] ),
    .A(\inbuf[4] ),
    .Y(_0502_),
    .D(\inbuf[7] ));
 sg13g2_nand2b_2 _1133_ (.Y(_0503_),
    .B(_0502_),
    .A_N(_0501_));
 sg13g2_nor2b_1 _1134_ (.A(_0503_),
    .B_N(_0500_),
    .Y(_0504_));
 sg13g2_nor2_1 _1135_ (.A(_0236_),
    .B(_0269_),
    .Y(_0505_));
 sg13g2_o21ai_1 _1136_ (.B1(net10),
    .Y(_0506_),
    .A1(_0303_),
    .A2(_0505_));
 sg13g2_nor2_2 _1137_ (.A(_0220_),
    .B(_0237_),
    .Y(_0507_));
 sg13g2_nand2_1 _1138_ (.Y(_0508_),
    .A(_0489_),
    .B(_0507_));
 sg13g2_and3_1 _1139_ (.X(_0509_),
    .A(_0294_),
    .B(_0506_),
    .C(_0508_));
 sg13g2_a21oi_1 _1140_ (.A1(_0154_),
    .A2(_0271_),
    .Y(_0510_),
    .B1(_0504_));
 sg13g2_nand4_1 _1141_ (.B(_0486_),
    .C(_0509_),
    .A(_0301_),
    .Y(_0511_),
    .D(_0510_));
 sg13g2_or4_2 _1142_ (.A(\counter[13] ),
    .B(\counter[12] ),
    .C(\counter[14] ),
    .D(\counter[15] ),
    .X(_0512_));
 sg13g2_nand3_1 _1143_ (.B(_0140_),
    .C(_0340_),
    .A(_0138_),
    .Y(_0513_));
 sg13g2_nor3_2 _1144_ (.A(_0331_),
    .B(_0512_),
    .C(_0513_),
    .Y(_0514_));
 sg13g2_nand2_1 _1145_ (.Y(_0515_),
    .A(_0226_),
    .B(_0514_));
 sg13g2_and2_1 _1146_ (.A(_0199_),
    .B(_0514_),
    .X(_0516_));
 sg13g2_nor2_1 _1147_ (.A(_0239_),
    .B(_0516_),
    .Y(_0517_));
 sg13g2_nor2_1 _1148_ (.A(_0501_),
    .B(_0502_),
    .Y(_0518_));
 sg13g2_nor4_1 _1149_ (.A(_0225_),
    .B(_0253_),
    .C(_0297_),
    .D(_0518_),
    .Y(_0519_));
 sg13g2_nand4_1 _1150_ (.B(net207),
    .C(_0187_),
    .A(_0138_),
    .Y(_0520_),
    .D(_0274_));
 sg13g2_nor3_2 _1151_ (.A(_0277_),
    .B(_0512_),
    .C(_0520_),
    .Y(_0521_));
 sg13g2_nand2b_1 _1152_ (.Y(_0522_),
    .B(_0521_),
    .A_N(_0296_));
 sg13g2_nor2_1 _1153_ (.A(net226),
    .B(_0399_),
    .Y(_0523_));
 sg13g2_nor2_1 _1154_ (.A(_0303_),
    .B(_0523_),
    .Y(_0524_));
 sg13g2_and4_1 _1155_ (.A(_0269_),
    .B(_0285_),
    .C(_0287_),
    .D(_0524_),
    .X(_0525_));
 sg13g2_a21oi_1 _1156_ (.A1(_0237_),
    .A2(_0249_),
    .Y(_0526_),
    .B1(_0248_));
 sg13g2_nand3_1 _1157_ (.B(_0522_),
    .C(_0525_),
    .A(_0519_),
    .Y(_0527_));
 sg13g2_a21oi_1 _1158_ (.A1(_0515_),
    .A2(_0517_),
    .Y(_0528_),
    .B1(_0527_));
 sg13g2_nand2_1 _1159_ (.Y(_0529_),
    .A(net81),
    .B(_0511_));
 sg13g2_o21ai_1 _1160_ (.B1(_0529_),
    .Y(_0069_),
    .A1(_0511_),
    .A2(_0528_));
 sg13g2_nor3_1 _1161_ (.A(_0302_),
    .B(_0517_),
    .C(_0526_),
    .Y(_0530_));
 sg13g2_nor2_1 _1162_ (.A(_0296_),
    .B(_0521_),
    .Y(_0531_));
 sg13g2_nor2_1 _1163_ (.A(net192),
    .B(_0531_),
    .Y(_0532_));
 sg13g2_inv_1 _1164_ (.Y(_0533_),
    .A(_0532_));
 sg13g2_nor4_2 _1165_ (.A(_0295_),
    .B(_0505_),
    .C(_0518_),
    .Y(_0534_),
    .D(_0533_));
 sg13g2_a21oi_1 _1166_ (.A1(_0224_),
    .A2(_0399_),
    .Y(_0535_),
    .B1(_0234_));
 sg13g2_nand2_1 _1167_ (.Y(_0536_),
    .A(_0265_),
    .B(_0268_));
 sg13g2_nor4_1 _1168_ (.A(_0270_),
    .B(_0400_),
    .C(_0535_),
    .D(_0536_),
    .Y(_0537_));
 sg13g2_nand3_1 _1169_ (.B(_0534_),
    .C(_0537_),
    .A(_0530_),
    .Y(_0538_));
 sg13g2_mux2_1 _1170_ (.A0(_0538_),
    .A1(net224),
    .S(_0511_),
    .X(_0070_));
 sg13g2_a22oi_1 _1171_ (.Y(_0539_),
    .B1(_0226_),
    .B2(_0238_),
    .A2(_0225_),
    .A1(_0205_));
 sg13g2_nand2b_1 _1172_ (.Y(_0540_),
    .B(_0514_),
    .A_N(_0539_));
 sg13g2_nor2b_1 _1173_ (.A(_0290_),
    .B_N(_0265_),
    .Y(_0541_));
 sg13g2_and4_1 _1174_ (.A(_0246_),
    .B(_0287_),
    .C(_0312_),
    .D(_0541_),
    .X(_0542_));
 sg13g2_nand3_1 _1175_ (.B(_0540_),
    .C(_0542_),
    .A(_0534_),
    .Y(_0543_));
 sg13g2_mux2_1 _1176_ (.A0(_0543_),
    .A1(net223),
    .S(_0511_),
    .X(_0071_));
 sg13g2_nor2_1 _1177_ (.A(_0298_),
    .B(_0516_),
    .Y(_0544_));
 sg13g2_nor2_1 _1178_ (.A(_0251_),
    .B(_0399_),
    .Y(_0545_));
 sg13g2_nor2_1 _1179_ (.A(_0544_),
    .B(_0545_),
    .Y(_0546_));
 sg13g2_nand2_2 _1180_ (.Y(_0547_),
    .A(_0222_),
    .B(_0286_));
 sg13g2_and4_1 _1181_ (.A(_0224_),
    .B(_0265_),
    .C(_0483_),
    .D(_0547_),
    .X(_0548_));
 sg13g2_nand4_1 _1182_ (.B(_0532_),
    .C(_0546_),
    .A(_0503_),
    .Y(_0549_),
    .D(_0548_));
 sg13g2_mux2_1 _1183_ (.A0(_0549_),
    .A1(net222),
    .S(_0511_),
    .X(_0072_));
 sg13g2_nor2b_1 _1184_ (.A(_0289_),
    .B_N(_0501_),
    .Y(_0550_));
 sg13g2_and4_1 _1185_ (.A(_0287_),
    .B(_0312_),
    .C(_0547_),
    .D(_0550_),
    .X(_0551_));
 sg13g2_nand4_1 _1186_ (.B(_0530_),
    .C(_0546_),
    .A(_0522_),
    .Y(_0552_),
    .D(_0551_));
 sg13g2_mux2_1 _1187_ (.A0(_0552_),
    .A1(net220),
    .S(_0511_),
    .X(_0073_));
 sg13g2_and3_1 _1188_ (.X(_0553_),
    .A(_0254_),
    .B(_0268_),
    .C(_0547_));
 sg13g2_nand3_1 _1189_ (.B(_0268_),
    .C(_0547_),
    .A(_0254_),
    .Y(_0554_));
 sg13g2_nand2_2 _1190_ (.Y(_0555_),
    .A(_0258_),
    .B(_0553_));
 sg13g2_inv_2 _1191_ (.Y(_0556_),
    .A(_0555_));
 sg13g2_nor2_1 _1192_ (.A(_0300_),
    .B(_0555_),
    .Y(_0557_));
 sg13g2_a22oi_1 _1193_ (.Y(_0558_),
    .B1(_0484_),
    .B2(_0557_),
    .A2(_0300_),
    .A1(_0143_));
 sg13g2_nand3_1 _1194_ (.B(_0281_),
    .C(_0557_),
    .A(net116),
    .Y(_0559_));
 sg13g2_o21ai_1 _1195_ (.B1(_0559_),
    .Y(_0560_),
    .A1(net217),
    .A2(_0299_));
 sg13g2_mux2_1 _1196_ (.A0(net217),
    .A1(_0560_),
    .S(net190),
    .X(_0074_));
 sg13g2_nor2b_1 _1197_ (.A(net190),
    .B_N(net216),
    .Y(_0561_));
 sg13g2_nand2_1 _1198_ (.Y(_0562_),
    .A(_0556_),
    .B(net188));
 sg13g2_nor3_1 _1199_ (.A(_0186_),
    .B(_0213_),
    .C(_0562_),
    .Y(_0563_));
 sg13g2_or2_1 _1200_ (.X(_0075_),
    .B(_0563_),
    .A(_0561_));
 sg13g2_nand2_1 _1201_ (.Y(_0564_),
    .A(_0213_),
    .B(net190));
 sg13g2_xor2_1 _1202_ (.B(_0564_),
    .A(net214),
    .X(_0565_));
 sg13g2_nor2_1 _1203_ (.A(_0555_),
    .B(_0565_),
    .Y(_0076_));
 sg13g2_or2_1 _1204_ (.X(_0566_),
    .B(_0564_),
    .A(net104));
 sg13g2_a21oi_2 _1205_ (.B1(_0555_),
    .Y(_0567_),
    .A2(_0299_),
    .A1(_0284_));
 sg13g2_nor2b_2 _1206_ (.A(_0567_),
    .B_N(net189),
    .Y(_0568_));
 sg13g2_xnor2_1 _1207_ (.Y(_0569_),
    .A(_0137_),
    .B(_0566_));
 sg13g2_nor2_1 _1208_ (.A(_0568_),
    .B(_0569_),
    .Y(_0077_));
 sg13g2_a21oi_1 _1209_ (.A1(_0274_),
    .A2(net190),
    .Y(_0570_),
    .B1(net108));
 sg13g2_and3_1 _1210_ (.X(_0571_),
    .A(\counter[4] ),
    .B(_0274_),
    .C(net190));
 sg13g2_nor3_1 _1211_ (.A(_0555_),
    .B(net109),
    .C(_0571_),
    .Y(_0078_));
 sg13g2_nand2_1 _1212_ (.Y(_0572_),
    .A(\counter[5] ),
    .B(_0571_));
 sg13g2_o21ai_1 _1213_ (.B1(_0556_),
    .Y(_0573_),
    .A1(net117),
    .A2(_0571_));
 sg13g2_nor2b_1 _1214_ (.A(_0573_),
    .B_N(_0572_),
    .Y(_0079_));
 sg13g2_nand2_1 _1215_ (.Y(_0574_),
    .A(_0275_),
    .B(_0556_));
 sg13g2_a22oi_1 _1216_ (.Y(_0080_),
    .B1(_0574_),
    .B2(net190),
    .A2(_0572_),
    .A1(_0138_));
 sg13g2_xor2_1 _1217_ (.B(_0275_),
    .A(net114),
    .X(_0575_));
 sg13g2_nand3_1 _1218_ (.B(_0567_),
    .C(_0575_),
    .A(net188),
    .Y(_0576_));
 sg13g2_o21ai_1 _1219_ (.B1(_0576_),
    .Y(_0081_),
    .A1(_0139_),
    .A2(net189));
 sg13g2_nor2_1 _1220_ (.A(_0139_),
    .B(_0275_),
    .Y(_0577_));
 sg13g2_a21oi_1 _1221_ (.A1(net188),
    .A2(_0577_),
    .Y(_0578_),
    .B1(net210));
 sg13g2_and3_1 _1222_ (.X(_0579_),
    .A(net210),
    .B(net188),
    .C(_0577_));
 sg13g2_nor3_1 _1223_ (.A(_0555_),
    .B(_0578_),
    .C(_0579_),
    .Y(_0082_));
 sg13g2_and2_1 _1224_ (.A(net209),
    .B(_0579_),
    .X(_0580_));
 sg13g2_o21ai_1 _1225_ (.B1(_0556_),
    .Y(_0581_),
    .A1(net209),
    .A2(_0579_));
 sg13g2_nor2_1 _1226_ (.A(_0580_),
    .B(_0581_),
    .Y(_0083_));
 sg13g2_o21ai_1 _1227_ (.B1(net188),
    .Y(_0582_),
    .A1(_0278_),
    .A2(_0555_));
 sg13g2_o21ai_1 _1228_ (.B1(_0582_),
    .Y(_0583_),
    .A1(net208),
    .A2(_0580_));
 sg13g2_inv_1 _1229_ (.Y(_0084_),
    .A(_0583_));
 sg13g2_o21ai_1 _1230_ (.B1(net188),
    .Y(_0584_),
    .A1(net111),
    .A2(_0278_));
 sg13g2_a21oi_1 _1231_ (.A1(net111),
    .A2(_0278_),
    .Y(_0585_),
    .B1(_0584_));
 sg13g2_nor2_1 _1232_ (.A(net207),
    .B(net188),
    .Y(_0586_));
 sg13g2_nor3_1 _1233_ (.A(_0568_),
    .B(_0585_),
    .C(_0586_),
    .Y(_0085_));
 sg13g2_nand2_1 _1234_ (.Y(_0587_),
    .A(_0279_),
    .B(_0556_));
 sg13g2_nand2_1 _1235_ (.Y(_0588_),
    .A(net189),
    .B(_0587_));
 sg13g2_nand3_1 _1236_ (.B(_0278_),
    .C(net188),
    .A(net207),
    .Y(_0589_));
 sg13g2_a22oi_1 _1237_ (.Y(_0086_),
    .B1(_0589_),
    .B2(_0142_),
    .A2(_0587_),
    .A1(net189));
 sg13g2_nor3_1 _1238_ (.A(net93),
    .B(_0279_),
    .C(_0562_),
    .Y(_0590_));
 sg13g2_a21o_1 _1239_ (.A2(_0588_),
    .A1(net93),
    .B1(_0590_),
    .X(_0087_));
 sg13g2_a21oi_1 _1240_ (.A1(_0280_),
    .A2(net189),
    .Y(_0591_),
    .B1(net72));
 sg13g2_nor2b_1 _1241_ (.A(_0283_),
    .B_N(net189),
    .Y(_0592_));
 sg13g2_nor3_1 _1242_ (.A(_0555_),
    .B(net73),
    .C(_0592_),
    .Y(_0088_));
 sg13g2_xnor2_1 _1243_ (.Y(_0593_),
    .A(net98),
    .B(_0592_));
 sg13g2_nor2_1 _1244_ (.A(_0568_),
    .B(_0593_),
    .Y(_0089_));
 sg13g2_o21ai_1 _1245_ (.B1(_0553_),
    .Y(_0594_),
    .A1(_0281_),
    .A2(_0484_));
 sg13g2_a21oi_1 _1246_ (.A1(_0284_),
    .A2(_0485_),
    .Y(_0595_),
    .B1(net79));
 sg13g2_a21oi_1 _1247_ (.A1(net79),
    .A2(_0594_),
    .Y(_0090_),
    .B1(_0595_));
 sg13g2_a21oi_1 _1248_ (.A1(\timer[0] ),
    .A2(_0594_),
    .Y(_0596_),
    .B1(net65));
 sg13g2_nor3_1 _1249_ (.A(_0272_),
    .B(_0281_),
    .C(_0484_),
    .Y(_0597_));
 sg13g2_nor3_1 _1250_ (.A(_0554_),
    .B(net66),
    .C(_0597_),
    .Y(_0091_));
 sg13g2_and2_1 _1251_ (.A(net101),
    .B(_0597_),
    .X(_0598_));
 sg13g2_o21ai_1 _1252_ (.B1(_0553_),
    .Y(_0599_),
    .A1(net101),
    .A2(_0597_));
 sg13g2_nor2_1 _1253_ (.A(_0598_),
    .B(_0599_),
    .Y(_0092_));
 sg13g2_a21oi_1 _1254_ (.A1(net102),
    .A2(_0598_),
    .Y(_0600_),
    .B1(_0554_));
 sg13g2_o21ai_1 _1255_ (.B1(_0600_),
    .Y(_0601_),
    .A1(net102),
    .A2(_0598_));
 sg13g2_inv_1 _1256_ (.Y(_0093_),
    .A(_0601_));
 sg13g2_nor2_1 _1257_ (.A(_0500_),
    .B(_0503_),
    .Y(_0602_));
 sg13g2_a21oi_1 _1258_ (.A1(\spi.done ),
    .A2(_0227_),
    .Y(_0603_),
    .B1(_0298_));
 sg13g2_or2_1 _1259_ (.X(_0604_),
    .B(_0507_),
    .A(_0297_));
 sg13g2_o21ai_1 _1260_ (.B1(_0501_),
    .Y(_0605_),
    .A1(_0234_),
    .A2(_0399_));
 sg13g2_o21ai_1 _1261_ (.B1(_0508_),
    .Y(_0606_),
    .A1(_0604_),
    .A2(_0605_));
 sg13g2_nor3_1 _1262_ (.A(_0602_),
    .B(_0603_),
    .C(_0606_),
    .Y(_0607_));
 sg13g2_nor2_1 _1263_ (.A(net63),
    .B(_0607_),
    .Y(_0608_));
 sg13g2_o21ai_1 _1264_ (.B1(_0502_),
    .Y(_0609_),
    .A1(_0234_),
    .A2(_0399_));
 sg13g2_nand2b_1 _1265_ (.Y(_0610_),
    .B(_0609_),
    .A_N(_0604_));
 sg13g2_a21oi_1 _1266_ (.A1(_0607_),
    .A2(_0610_),
    .Y(_0094_),
    .B1(_0608_));
 sg13g2_nor4_1 _1267_ (.A(net225),
    .B(\state[0] ),
    .C(net220),
    .D(_0245_),
    .Y(_0611_));
 sg13g2_o21ai_1 _1268_ (.B1(_0503_),
    .Y(_0612_),
    .A1(_0507_),
    .A2(_0611_));
 sg13g2_nor2b_1 _1269_ (.A(_0612_),
    .B_N(_0508_),
    .Y(_0613_));
 sg13g2_nor2_1 _1270_ (.A(net99),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_a21oi_1 _1271_ (.A1(net225),
    .A2(_0613_),
    .Y(_0095_),
    .B1(_0614_));
 sg13g2_nand2_1 _1272_ (.Y(_0615_),
    .A(net223),
    .B(_0143_));
 sg13g2_nand3_1 _1273_ (.B(_0286_),
    .C(_0615_),
    .A(net222),
    .Y(_0616_));
 sg13g2_o21ai_1 _1274_ (.B1(net68),
    .Y(_0617_),
    .A1(_0544_),
    .A2(_0616_));
 sg13g2_nand2_1 _1275_ (.Y(_0096_),
    .A(_0547_),
    .B(_0617_));
 sg13g2_mux2_1 _1276_ (.A0(net200),
    .A1(net44),
    .S(_0170_),
    .X(_0097_));
 sg13g2_o21ai_1 _1277_ (.B1(_0016_),
    .Y(_0618_),
    .A1(\spi.state[1] ),
    .A2(\spi.state[2] ));
 sg13g2_nand2_1 _1278_ (.Y(_0619_),
    .A(_0028_),
    .B(net195));
 sg13g2_o21ai_1 _1279_ (.B1(_0619_),
    .Y(_0098_),
    .A1(net9),
    .A2(net195));
 sg13g2_nand2_1 _1280_ (.Y(_0620_),
    .A(_0029_),
    .B(net195));
 sg13g2_o21ai_1 _1281_ (.B1(_0620_),
    .Y(_0099_),
    .A1(\spi.rreg[0] ),
    .A2(net195));
 sg13g2_nand2_1 _1282_ (.Y(_0621_),
    .A(_0030_),
    .B(net194));
 sg13g2_o21ai_1 _1283_ (.B1(_0621_),
    .Y(_0100_),
    .A1(\spi.rreg[1] ),
    .A2(net193));
 sg13g2_nand2_1 _1284_ (.Y(_0622_),
    .A(_0031_),
    .B(net194));
 sg13g2_o21ai_1 _1285_ (.B1(_0622_),
    .Y(_0101_),
    .A1(\spi.rreg[2] ),
    .A2(net193));
 sg13g2_nand2_1 _1286_ (.Y(_0623_),
    .A(_0032_),
    .B(net194));
 sg13g2_o21ai_1 _1287_ (.B1(_0623_),
    .Y(_0102_),
    .A1(\spi.rreg[3] ),
    .A2(net194));
 sg13g2_nand2_1 _1288_ (.Y(_0624_),
    .A(_0033_),
    .B(net193));
 sg13g2_o21ai_1 _1289_ (.B1(_0624_),
    .Y(_0103_),
    .A1(\spi.rreg[4] ),
    .A2(net193));
 sg13g2_nand2_1 _1290_ (.Y(_0625_),
    .A(_0034_),
    .B(net193));
 sg13g2_o21ai_1 _1291_ (.B1(_0625_),
    .Y(_0104_),
    .A1(\spi.rreg[5] ),
    .A2(net193));
 sg13g2_nand2_1 _1292_ (.Y(_0626_),
    .A(_0035_),
    .B(net193));
 sg13g2_o21ai_1 _1293_ (.B1(_0626_),
    .Y(_0105_),
    .A1(\spi.rreg[6] ),
    .A2(net193));
 sg13g2_nor2_1 _1294_ (.A(\spi.state[1] ),
    .B(\spi.state[3] ),
    .Y(_0627_));
 sg13g2_nor3_1 _1295_ (.A(\spi.state[0] ),
    .B(\spi.state[2] ),
    .C(_0627_),
    .Y(_0628_));
 sg13g2_a22oi_1 _1296_ (.Y(_0106_),
    .B1(_0628_),
    .B2(_0166_),
    .A2(_0167_),
    .A1(_0131_));
 sg13g2_nor2b_2 _1297_ (.A(net196),
    .B_N(\spi.isck ),
    .Y(_0629_));
 sg13g2_or2_2 _1298_ (.X(_0630_),
    .B(\spi.isck ),
    .A(net196));
 sg13g2_nor2_1 _1299_ (.A(_0037_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_a221oi_1 _1300_ (.B2(_0629_),
    .C1(_0631_),
    .B1(\spi.treg[0] ),
    .A1(\spi.d_latched[0] ),
    .Y(_0107_),
    .A2(net196));
 sg13g2_nor2_1 _1301_ (.A(_0038_),
    .B(_0630_),
    .Y(_0632_));
 sg13g2_a221oi_1 _1302_ (.B2(_0629_),
    .C1(_0632_),
    .B1(\spi.treg[1] ),
    .A1(\spi.d_latched[1] ),
    .Y(_0108_),
    .A2(net196));
 sg13g2_nor2_1 _1303_ (.A(_0039_),
    .B(_0630_),
    .Y(_0633_));
 sg13g2_a221oi_1 _1304_ (.B2(_0629_),
    .C1(_0633_),
    .B1(\spi.treg[2] ),
    .A1(\spi.d_latched[2] ),
    .Y(_0109_),
    .A2(\spi.w_latched ));
 sg13g2_nor2_1 _1305_ (.A(_0040_),
    .B(_0630_),
    .Y(_0634_));
 sg13g2_a221oi_1 _1306_ (.B2(_0629_),
    .C1(_0634_),
    .B1(\spi.treg[3] ),
    .A1(\spi.d_latched[3] ),
    .Y(_0110_),
    .A2(\spi.w_latched ));
 sg13g2_nor2_1 _1307_ (.A(_0041_),
    .B(_0630_),
    .Y(_0635_));
 sg13g2_a221oi_1 _1308_ (.B2(_0629_),
    .C1(_0635_),
    .B1(\spi.treg[4] ),
    .A1(\spi.d_latched[4] ),
    .Y(_0111_),
    .A2(net197));
 sg13g2_nor2_1 _1309_ (.A(_0042_),
    .B(_0630_),
    .Y(_0636_));
 sg13g2_a221oi_1 _1310_ (.B2(_0629_),
    .C1(_0636_),
    .B1(\spi.treg[5] ),
    .A1(\spi.d_latched[5] ),
    .Y(_0112_),
    .A2(net197));
 sg13g2_nor2_1 _1311_ (.A(_0043_),
    .B(_0630_),
    .Y(_0637_));
 sg13g2_a221oi_1 _1312_ (.B2(_0629_),
    .C1(_0637_),
    .B1(\spi.treg[6] ),
    .A1(\spi.d_latched[6] ),
    .Y(_0113_),
    .A2(net197));
 sg13g2_nand2b_1 _1313_ (.Y(_0638_),
    .B(_0629_),
    .A_N(\spi.treg[7] ));
 sg13g2_o21ai_1 _1314_ (.B1(_0638_),
    .Y(_0639_),
    .A1(\spi.mosi ),
    .A2(_0630_));
 sg13g2_a21oi_1 _1315_ (.A1(_0128_),
    .A2(net197),
    .Y(_0114_),
    .B1(_0639_));
 sg13g2_a21oi_1 _1316_ (.A1(\spi.state[3] ),
    .A2(_0158_),
    .Y(_0640_),
    .B1(\spi.state[0] ));
 sg13g2_nor3_1 _1317_ (.A(net196),
    .B(_0134_),
    .C(\spi.stream ),
    .Y(_0641_));
 sg13g2_a21oi_1 _1318_ (.A1(_0134_),
    .A2(_0017_),
    .Y(_0642_),
    .B1(_0641_));
 sg13g2_mux2_1 _1319_ (.A0(_0642_),
    .A1(_0044_),
    .S(_0640_),
    .X(_0115_));
 sg13g2_nand2b_1 _1320_ (.Y(_0643_),
    .B(\spi.done ),
    .A_N(\spi.stream ));
 sg13g2_and2_1 _1321_ (.A(net50),
    .B(_0643_),
    .X(_0116_));
 sg13g2_or3_1 _1322_ (.A(\spi.state[0] ),
    .B(_0135_),
    .C(\spi.state[2] ),
    .X(_0644_));
 sg13g2_and2_1 _1323_ (.A(_0167_),
    .B(_0644_),
    .X(_0645_));
 sg13g2_nand2_1 _1324_ (.Y(_0646_),
    .A(\spi.nbit[0] ),
    .B(_0645_));
 sg13g2_o21ai_1 _1325_ (.B1(_0646_),
    .Y(_0117_),
    .A1(\spi.nbit[0] ),
    .A2(_0644_));
 sg13g2_nand2_1 _1326_ (.Y(_0647_),
    .A(\spi.nbit[1] ),
    .B(_0645_));
 sg13g2_xnor2_1 _1327_ (.Y(_0648_),
    .A(\spi.nbit[0] ),
    .B(\spi.nbit[1] ));
 sg13g2_o21ai_1 _1328_ (.B1(_0647_),
    .Y(_0118_),
    .A1(_0644_),
    .A2(_0648_));
 sg13g2_and2_1 _1329_ (.A(_0013_),
    .B(_0165_),
    .X(_0649_));
 sg13g2_nor4_1 _1330_ (.A(\spi.state[0] ),
    .B(\spi.state[2] ),
    .C(_0166_),
    .D(_0649_),
    .Y(_0650_));
 sg13g2_a21o_1 _1331_ (.A2(_0645_),
    .A1(\spi.nbit[2] ),
    .B1(_0650_),
    .X(_0119_));
 sg13g2_inv_1 _1333__3 (.Y(net29),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _1334__4 (.Y(net30),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _1335__5 (.Y(net31),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _1336__6 (.Y(net32),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _1337__7 (.Y(net33),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _1338__8 (.Y(net34),
    .A(clknet_1_1__leaf_clk));
 sg13g2_inv_1 _1339__9 (.Y(net35),
    .A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbp_1 _1340_ (.CLK(net201),
    .RESET_B(net235),
    .D(_0045_),
    .Q_N(\spi.state[0] ),
    .Q(_0023_));
 sg13g2_dfrbp_1 _1341_ (.CLK(net201),
    .RESET_B(net234),
    .D(\spi.state[2] ),
    .Q_N(_0695_),
    .Q(\spi.state[1] ));
 sg13g2_dfrbp_1 _1342_ (.CLK(net200),
    .RESET_B(net234),
    .D(_0001_),
    .Q_N(_0696_),
    .Q(\spi.state[2] ));
 sg13g2_dfrbp_1 _1343_ (.CLK(net200),
    .RESET_B(net234),
    .D(_0000_),
    .Q_N(_0694_),
    .Q(\spi.state[3] ));
 sg13g2_dfrbp_1 _1344_ (.CLK(net201),
    .RESET_B(net234),
    .D(_0055_),
    .Q_N(\spi.treg[0] ),
    .Q(_0024_));
 sg13g2_dfrbp_1 _1345_ (.CLK(net27),
    .RESET_B(net235),
    .D(_0056_),
    .Q_N(_0693_),
    .Q(\spi.w_latched ));
 sg13g2_dfrbp_1 _1346_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net232),
    .D(net71),
    .Q_N(dcb),
    .Q(_0025_));
 sg13g2_dfrbp_1 _1347_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net231),
    .D(net60),
    .Q_N(resetb),
    .Q(_0026_));
 sg13g2_dfrbp_1 _1348_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net240),
    .D(_0059_),
    .Q_N(_0014_),
    .Q(\spi.reg_dat_we ));
 sg13g2_dfrbp_1 _1349_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net240),
    .D(_0060_),
    .Q_N(_0692_),
    .Q(stream));
 sg13g2_dfrbp_1 _1350_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net235),
    .D(_0061_),
    .Q_N(_0691_),
    .Q(\data_out[0] ));
 sg13g2_dfrbp_1 _1351_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net235),
    .D(_0062_),
    .Q_N(_0690_),
    .Q(\data_out[1] ));
 sg13g2_dfrbp_1 _1352_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net235),
    .D(_0063_),
    .Q_N(_0689_),
    .Q(\data_out[2] ));
 sg13g2_dfrbp_1 _1353_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net236),
    .D(_0064_),
    .Q_N(_0688_),
    .Q(\data_out[3] ));
 sg13g2_dfrbp_1 _1354_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net236),
    .D(net54),
    .Q_N(_0687_),
    .Q(\data_out[4] ));
 sg13g2_dfrbp_1 _1355_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net238),
    .D(net47),
    .Q_N(_0686_),
    .Q(\data_out[5] ));
 sg13g2_dfrbp_1 _1356_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net238),
    .D(net49),
    .Q_N(_0685_),
    .Q(\data_out[6] ));
 sg13g2_dfrbp_1 _1357_ (.CLK(clknet_4_10_0_clk_regs),
    .RESET_B(net239),
    .D(_0068_),
    .Q_N(_0684_),
    .Q(\data_out[7] ));
 sg13g2_dfrbp_1 _1358_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net244),
    .D(_0069_),
    .Q_N(_0683_),
    .Q(\state[0] ));
 sg13g2_dfrbp_1 _1359_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net240),
    .D(_0070_),
    .Q_N(_0682_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 _1360_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net233),
    .D(_0071_),
    .Q_N(_0681_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 _1361_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net233),
    .D(_0072_),
    .Q_N(_0680_),
    .Q(\state[3] ));
 sg13g2_dfrbp_1 _1362_ (.CLK(clknet_4_9_0_clk_regs),
    .RESET_B(net240),
    .D(_0073_),
    .Q_N(_0012_),
    .Q(\state[4] ));
 sg13g2_dfrbp_1 _1363_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net231),
    .D(_0074_),
    .Q_N(_0018_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _1364_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net229),
    .D(_0075_),
    .Q_N(_0679_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _1365_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net233),
    .D(_0076_),
    .Q_N(_0015_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _1366_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net231),
    .D(_0077_),
    .Q_N(_0678_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _1367_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net229),
    .D(_0078_),
    .Q_N(_0677_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _1368_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net229),
    .D(net118),
    .Q_N(_0676_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _1369_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net228),
    .D(net106),
    .Q_N(_0675_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _1370_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net231),
    .D(net115),
    .Q_N(_0019_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _1371_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net228),
    .D(_0082_),
    .Q_N(_0674_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _1372_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net227),
    .D(_0083_),
    .Q_N(_0673_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _1373_ (.CLK(clknet_4_1_0_clk_regs),
    .RESET_B(net227),
    .D(_0084_),
    .Q_N(_0672_),
    .Q(\counter[10] ));
 sg13g2_dfrbp_1 _1374_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net228),
    .D(net112),
    .Q_N(_0020_),
    .Q(\counter[11] ));
 sg13g2_dfrbp_1 _1375_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net228),
    .D(net75),
    .Q_N(_0671_),
    .Q(\counter[12] ));
 sg13g2_dfrbp_1 _1376_ (.CLK(clknet_4_4_0_clk_regs),
    .RESET_B(net231),
    .D(_0087_),
    .Q_N(_0670_),
    .Q(\counter[13] ));
 sg13g2_dfrbp_1 _1377_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net231),
    .D(_0088_),
    .Q_N(_0669_),
    .Q(\counter[14] ));
 sg13g2_dfrbp_1 _1378_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net231),
    .D(_0089_),
    .Q_N(_0668_),
    .Q(\counter[15] ));
 sg13g2_dfrbp_1 _1379_ (.CLK(clknet_4_6_0_clk_regs),
    .RESET_B(net231),
    .D(net80),
    .Q_N(_0667_),
    .Q(\timer[0] ));
 sg13g2_dfrbp_1 _1380_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net232),
    .D(net67),
    .Q_N(_0666_),
    .Q(\timer[1] ));
 sg13g2_dfrbp_1 _1381_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net232),
    .D(_0092_),
    .Q_N(_0665_),
    .Q(\timer[2] ));
 sg13g2_dfrbp_1 _1382_ (.CLK(clknet_4_5_0_clk_regs),
    .RESET_B(net232),
    .D(_0093_),
    .Q_N(_0664_),
    .Q(\timer[3] ));
 sg13g2_dfrbp_1 _1383_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net233),
    .D(_0094_),
    .Q_N(sramcsb),
    .Q(_0027_));
 sg13g2_dfrbp_1 _1384_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net240),
    .D(net100),
    .Q_N(_0697_),
    .Q(passthru));
 sg13g2_dfrbp_1 _1385_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net241),
    .D(net1),
    .Q_N(_0698_),
    .Q(\inbuf[0] ));
 sg13g2_dfrbp_1 _1386_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net241),
    .D(net2),
    .Q_N(_0699_),
    .Q(\inbuf[1] ));
 sg13g2_dfrbp_1 _1387_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net242),
    .D(net3),
    .Q_N(_0700_),
    .Q(\inbuf[2] ));
 sg13g2_dfrbp_1 _1388_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net242),
    .D(net4),
    .Q_N(_0701_),
    .Q(\inbuf[3] ));
 sg13g2_dfrbp_1 _1389_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net242),
    .D(net5),
    .Q_N(_0702_),
    .Q(\inbuf[4] ));
 sg13g2_dfrbp_1 _1390_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net241),
    .D(net6),
    .Q_N(_0703_),
    .Q(\inbuf[5] ));
 sg13g2_dfrbp_1 _1391_ (.CLK(clknet_4_13_0_clk_regs),
    .RESET_B(net241),
    .D(net7),
    .Q_N(_0704_),
    .Q(\inbuf[6] ));
 sg13g2_dfrbp_1 _1392_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net241),
    .D(net8),
    .Q_N(_0705_),
    .Q(\inbuf[7] ));
 sg13g2_dfrbp_1 _1393_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net243),
    .D(net38),
    .Q_N(_0021_),
    .Q(\inval[0] ));
 sg13g2_dfrbp_1 _1394_ (.CLK(clknet_4_15_0_clk_regs),
    .RESET_B(net241),
    .D(net36),
    .Q_N(_0022_),
    .Q(\inval[1] ));
 sg13g2_dfrbp_1 _1395_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net242),
    .D(net39),
    .Q_N(_0706_),
    .Q(\inval[2] ));
 sg13g2_dfrbp_1 _1396_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net242),
    .D(net37),
    .Q_N(_0707_),
    .Q(\inval[3] ));
 sg13g2_dfrbp_1 _1397_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net242),
    .D(net43),
    .Q_N(_0708_),
    .Q(\inval[4] ));
 sg13g2_dfrbp_1 _1398_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net241),
    .D(net40),
    .Q_N(_0709_),
    .Q(\inval[5] ));
 sg13g2_dfrbp_1 _1399_ (.CLK(clknet_4_12_0_clk_regs),
    .RESET_B(net241),
    .D(net41),
    .Q_N(_0710_),
    .Q(\inval[6] ));
 sg13g2_dfrbp_1 _1400_ (.CLK(clknet_4_14_0_clk_regs),
    .RESET_B(net242),
    .D(net42),
    .Q_N(_0663_),
    .Q(\inval[7] ));
 sg13g2_dfrbp_1 _1401_ (.CLK(clknet_4_7_0_clk_regs),
    .RESET_B(net233),
    .D(net69),
    .Q_N(_0662_),
    .Q(maskcsb));
 sg13g2_dfrbp_1 _1402_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net229),
    .D(net45),
    .Q_N(_0011_),
    .Q(\spi.hsck ));
 sg13g2_dfrbp_1 _1403_ (.CLK(net202),
    .RESET_B(net240),
    .D(_0098_),
    .Q_N(\spi.rreg[0] ),
    .Q(_0028_));
 sg13g2_dfrbp_1 _1404_ (.CLK(net202),
    .RESET_B(net243),
    .D(_0099_),
    .Q_N(\spi.rreg[1] ),
    .Q(_0029_));
 sg13g2_dfrbp_1 _1405_ (.CLK(net202),
    .RESET_B(net243),
    .D(_0100_),
    .Q_N(\spi.rreg[2] ),
    .Q(_0030_));
 sg13g2_dfrbp_1 _1406_ (.CLK(net202),
    .RESET_B(net243),
    .D(_0101_),
    .Q_N(\spi.rreg[3] ),
    .Q(_0031_));
 sg13g2_dfrbp_1 _1407_ (.CLK(net202),
    .RESET_B(net243),
    .D(_0102_),
    .Q_N(\spi.rreg[4] ),
    .Q(_0032_));
 sg13g2_dfrbp_1 _1408_ (.CLK(net202),
    .RESET_B(net243),
    .D(_0103_),
    .Q_N(\spi.rreg[5] ),
    .Q(_0033_));
 sg13g2_dfrbp_1 _1409_ (.CLK(net202),
    .RESET_B(net238),
    .D(_0104_),
    .Q_N(\spi.rreg[6] ),
    .Q(_0034_));
 sg13g2_dfrbp_1 _1410_ (.CLK(net202),
    .RESET_B(net238),
    .D(_0105_),
    .Q_N(\spi.rreg[7] ),
    .Q(_0035_));
 sg13g2_dfrbp_1 _1411_ (.CLK(net200),
    .RESET_B(net230),
    .D(_0106_),
    .Q_N(\spi.done ),
    .Q(_0036_));
 sg13g2_dfrbp_1 _1412_ (.CLK(net200),
    .RESET_B(net234),
    .D(_0010_),
    .Q_N(_0016_),
    .Q(\spi.isck ));
 sg13g2_dfrbp_1 _1413_ (.CLK(net203),
    .RESET_B(net234),
    .D(_0107_),
    .Q_N(\spi.treg[1] ),
    .Q(_0037_));
 sg13g2_dfrbp_1 _1414_ (.CLK(net203),
    .RESET_B(net236),
    .D(_0108_),
    .Q_N(\spi.treg[2] ),
    .Q(_0038_));
 sg13g2_dfrbp_1 _1415_ (.CLK(net203),
    .RESET_B(net236),
    .D(_0109_),
    .Q_N(\spi.treg[3] ),
    .Q(_0039_));
 sg13g2_dfrbp_1 _1416_ (.CLK(net203),
    .RESET_B(net237),
    .D(_0110_),
    .Q_N(\spi.treg[4] ),
    .Q(_0040_));
 sg13g2_dfrbp_1 _1417_ (.CLK(net203),
    .RESET_B(net237),
    .D(_0111_),
    .Q_N(\spi.treg[5] ),
    .Q(_0041_));
 sg13g2_dfrbp_1 _1418_ (.CLK(net203),
    .RESET_B(net237),
    .D(_0112_),
    .Q_N(\spi.treg[6] ),
    .Q(_0042_));
 sg13g2_dfrbp_1 _1419_ (.CLK(net203),
    .RESET_B(net236),
    .D(_0113_),
    .Q_N(\spi.treg[7] ),
    .Q(_0043_));
 sg13g2_dfrbp_1 _1420_ (.CLK(\spi.hsck ),
    .RESET_B(net238),
    .D(_0114_),
    .Q_N(_0661_),
    .Q(\spi.mosi ));
 sg13g2_dfrbp_1 _1421_ (.CLK(net201),
    .RESET_B(net240),
    .D(_0115_),
    .Q_N(mosienb),
    .Q(_0044_));
 sg13g2_dfrbp_1 _1422_ (.CLK(clknet_4_8_0_clk_regs),
    .RESET_B(net240),
    .D(net51),
    .Q_N(_0017_),
    .Q(\spi.stream ));
 sg13g2_dfrbp_1 _1423_ (.CLK(net200),
    .RESET_B(net229),
    .D(_0117_),
    .Q_N(_0660_),
    .Q(\spi.nbit[0] ));
 sg13g2_dfrbp_1 _1424_ (.CLK(net200),
    .RESET_B(net229),
    .D(_0118_),
    .Q_N(_0659_),
    .Q(\spi.nbit[1] ));
 sg13g2_dfrbp_1 _1425_ (.CLK(net200),
    .RESET_B(net230),
    .D(_0119_),
    .Q_N(_0013_),
    .Q(\spi.nbit[2] ));
 sg13g2_dfrbp_1 _1426_ (.CLK(net28),
    .RESET_B(net234),
    .D(_0120_),
    .Q_N(_0658_),
    .Q(\spi.d_latched[0] ));
 sg13g2_dfrbp_1 _1427_ (.CLK(net29),
    .RESET_B(net234),
    .D(_0121_),
    .Q_N(_0657_),
    .Q(\spi.d_latched[1] ));
 sg13g2_dfrbp_1 _1428_ (.CLK(net30),
    .RESET_B(net236),
    .D(_0122_),
    .Q_N(_0656_),
    .Q(\spi.d_latched[2] ));
 sg13g2_dfrbp_1 _1429_ (.CLK(net31),
    .RESET_B(net237),
    .D(_0123_),
    .Q_N(_0655_),
    .Q(\spi.d_latched[3] ));
 sg13g2_dfrbp_1 _1430_ (.CLK(net32),
    .RESET_B(net236),
    .D(_0124_),
    .Q_N(_0654_),
    .Q(\spi.d_latched[4] ));
 sg13g2_dfrbp_1 _1431_ (.CLK(net33),
    .RESET_B(net236),
    .D(_0125_),
    .Q_N(_0653_),
    .Q(\spi.d_latched[5] ));
 sg13g2_dfrbp_1 _1432_ (.CLK(net34),
    .RESET_B(net238),
    .D(_0126_),
    .Q_N(_0652_),
    .Q(\spi.d_latched[6] ));
 sg13g2_dfrbp_1 _1433_ (.CLK(net35),
    .RESET_B(net239),
    .D(_0127_),
    .Q_N(_0711_),
    .Q(\spi.d_latched[7] ));
 sg13g2_dfrbp_1 _1434_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net229),
    .D(net90),
    .Q_N(_0712_),
    .Q(\spi.count[0] ));
 sg13g2_dfrbp_1 _1435_ (.CLK(clknet_4_3_0_clk_regs),
    .RESET_B(net229),
    .D(net97),
    .Q_N(_0713_),
    .Q(\spi.count[1] ));
 sg13g2_dfrbp_1 _1436_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net227),
    .D(_0004_),
    .Q_N(_0714_),
    .Q(\spi.count[2] ));
 sg13g2_dfrbp_1 _1437_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net227),
    .D(net86),
    .Q_N(_0715_),
    .Q(\spi.count[3] ));
 sg13g2_dfrbp_1 _1438_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net227),
    .D(net95),
    .Q_N(_0716_),
    .Q(\spi.count[4] ));
 sg13g2_dfrbp_1 _1439_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net227),
    .D(_0007_),
    .Q_N(_0717_),
    .Q(\spi.count[5] ));
 sg13g2_dfrbp_1 _1440_ (.CLK(clknet_4_0_0_clk_regs),
    .RESET_B(net227),
    .D(net78),
    .Q_N(_0718_),
    .Q(\spi.count[6] ));
 sg13g2_dfrbp_1 _1441_ (.CLK(clknet_4_2_0_clk_regs),
    .RESET_B(net227),
    .D(net62),
    .Q_N(_0651_),
    .Q(\spi.count[7] ));
 sg13g2_tiehi tt_um_rte_eink_driver_23 (.L_HI(net23));
 sg13g2_tiehi tt_um_rte_eink_driver_24 (.L_HI(net24));
 sg13g2_tiehi tt_um_rte_eink_driver_25 (.L_HI(net25));
 sg13g2_tiehi tt_um_rte_eink_driver_26 (.L_HI(net26));
 sg13g2_inv_1 _0750__1 (.Y(net27),
    .A(clknet_1_0__leaf_clk));
 sg13g2_tielo tt_um_rte_eink_driver_12 (.L_LO(net12));
 sg13g2_tielo tt_um_rte_eink_driver_13 (.L_LO(net13));
 sg13g2_tielo tt_um_rte_eink_driver_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rte_eink_driver_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rte_eink_driver_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rte_eink_driver_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rte_eink_driver_18 (.L_LO(net18));
 sg13g2_tielo tt_um_rte_eink_driver_19 (.L_LO(net19));
 sg13g2_tielo tt_um_rte_eink_driver_20 (.L_LO(net20));
 sg13g2_tielo tt_um_rte_eink_driver_21 (.L_LO(net21));
 sg13g2_tiehi tt_um_rte_eink_driver_22 (.L_HI(net22));
 sg13g2_buf_1 _1458_ (.A(csb),
    .X(uio_out[0]));
 sg13g2_buf_1 _1459_ (.A(mosi),
    .X(uio_out[1]));
 sg13g2_buf_1 _1460_ (.A(sck),
    .X(uio_out[3]));
 sg13g2_buf_1 _1461_ (.A(sramcsb),
    .X(uio_out[4]));
 sg13g2_buf_1 _1462_ (.A(resetb),
    .X(uio_out[5]));
 sg13g2_buf_1 _1463_ (.A(dcb),
    .X(uio_out[7]));
 sg13g2_buf_1 _1464_ (.A(net9),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout187 (.A(_0412_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(net190),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(net190),
    .X(net189));
 sg13g2_buf_4 fanout190 (.X(net190),
    .A(_0558_));
 sg13g2_buf_4 fanout191 (.X(net191),
    .A(_0160_));
 sg13g2_buf_2 fanout192 (.A(_0313_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net195),
    .X(net193));
 sg13g2_buf_1 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_0618_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(net197),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(net124),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_0314_),
    .X(net198));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(_0180_));
 sg13g2_buf_2 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(\spi.hsck ),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(net203),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(\spi.hsck ),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(net205),
    .X(net204));
 sg13g2_buf_1 fanout205 (.A(\inval[4] ),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(net207),
    .X(net206));
 sg13g2_buf_1 fanout207 (.A(\counter[11] ),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(net121),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(net123),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(net113),
    .X(net210));
 sg13g2_buf_1 fanout211 (.A(\counter[8] ),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(\counter[7] ),
    .X(net212));
 sg13g2_buf_4 fanout213 (.X(net213),
    .A(\counter[3] ));
 sg13g2_buf_2 fanout214 (.A(net120),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(\counter[2] ),
    .X(net215));
 sg13g2_buf_4 fanout216 (.X(net216),
    .A(\counter[1] ));
 sg13g2_buf_4 fanout217 (.X(net217),
    .A(net219));
 sg13g2_buf_2 fanout218 (.A(net219),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(\counter[0] ),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(net119),
    .X(net220));
 sg13g2_buf_1 fanout221 (.A(\state[4] ),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(net122),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(net125),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(net225),
    .X(net224));
 sg13g2_buf_1 fanout225 (.A(\state[1] ),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(\state[0] ),
    .X(net226));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(net228));
 sg13g2_buf_4 fanout228 (.X(net228),
    .A(net230));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(net230));
 sg13g2_buf_2 fanout230 (.A(rst_n),
    .X(net230));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(net233));
 sg13g2_buf_2 fanout232 (.A(net233),
    .X(net232));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(rst_n));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(net239));
 sg13g2_buf_2 fanout235 (.A(net239),
    .X(net235));
 sg13g2_buf_4 fanout236 (.X(net236),
    .A(net238));
 sg13g2_buf_2 fanout237 (.A(net238),
    .X(net237));
 sg13g2_buf_4 fanout238 (.X(net238),
    .A(net239));
 sg13g2_buf_2 fanout239 (.A(net244),
    .X(net239));
 sg13g2_buf_4 fanout240 (.X(net240),
    .A(net244));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(net243));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(net243));
 sg13g2_buf_4 fanout243 (.X(net243),
    .A(net244));
 sg13g2_buf_2 fanout244 (.A(rst_n),
    .X(net244));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[6]),
    .X(net10));
 sg13g2_tielo tt_um_rte_eink_driver_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_4_1_0_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_4_2_0_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_4_3_0_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_4_4_0_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_4_5_0_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_4_6_0_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_4_7_0_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_4_9_0_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_4_10_0_clk_regs));
 sg13g2_inv_1 clkload10 (.A(clknet_4_11_0_clk_regs));
 sg13g2_inv_1 clkload11 (.A(clknet_4_12_0_clk_regs));
 sg13g2_inv_1 clkload12 (.A(clknet_4_13_0_clk_regs));
 sg13g2_inv_1 clkload13 (.A(clknet_4_14_0_clk_regs));
 sg13g2_inv_1 clkload14 (.A(clknet_4_15_0_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\inbuf[1] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold2 (.A(\inbuf[3] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold3 (.A(\inbuf[0] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold4 (.A(\inbuf[2] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold5 (.A(\inbuf[5] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold6 (.A(\inbuf[6] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold7 (.A(\inbuf[7] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold8 (.A(\inbuf[4] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0011_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0097_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold11 (.A(\data_out[5] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0066_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold13 (.A(\data_out[6] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0067_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold15 (.A(stream),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0116_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold17 (.A(\spi.d_latched[1] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold18 (.A(\data_out[4] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0065_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold20 (.A(\data_out[2] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold21 (.A(\spi.d_latched[7] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold22 (.A(\data_out[3] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold23 (.A(\data_out[7] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0026_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0058_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold26 (.A(\spi.count[7] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0009_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0027_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold29 (.A(\spi.d_latched[0] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold30 (.A(\timer[1] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0596_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0091_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold33 (.A(maskcsb),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0096_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0025_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0057_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold37 (.A(\counter[14] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0591_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold39 (.A(\counter[12] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0086_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold41 (.A(\spi.d_latched[4] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold42 (.A(\spi.count[6] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0008_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold44 (.A(\timer[0] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0090_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold46 (.A(\state[0] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold47 (.A(\spi.d_latched[2] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold48 (.A(\spi.d_latched[3] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold49 (.A(\spi.d_latched[5] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold50 (.A(\spi.count[3] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0005_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold52 (.A(\spi.d_latched[6] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold53 (.A(\data_out[0] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold54 (.A(\spi.count[0] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0002_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold56 (.A(\spi.reg_dat_we ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold57 (.A(\data_out[1] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold58 (.A(\counter[13] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold59 (.A(\spi.count[4] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0006_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold61 (.A(\spi.count[1] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0003_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold63 (.A(\counter[15] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold64 (.A(passthru),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0095_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold66 (.A(\timer[2] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold67 (.A(\timer[3] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0012_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0015_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold70 (.A(\counter[6] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0080_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold72 (.A(\spi.count[2] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold73 (.A(\counter[4] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0570_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold75 (.A(\spi.count[5] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0020_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0085_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold78 (.A(\counter[8] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0019_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0081_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0018_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold82 (.A(\counter[5] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0079_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold84 (.A(\state[4] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold85 (.A(\counter[2] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold86 (.A(\counter[10] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold87 (.A(\state[3] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold88 (.A(\counter[9] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold89 (.A(\spi.w_latched ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold90 (.A(\state[2] ),
    .X(net125));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_243 ();
 sg13g2_fill_2 FILLER_10_250 ();
 sg13g2_decap_8 FILLER_10_260 ();
 sg13g2_decap_8 FILLER_10_267 ();
 sg13g2_decap_4 FILLER_10_274 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_289 ();
 sg13g2_decap_8 FILLER_10_296 ();
 sg13g2_decap_8 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_19 ();
 sg13g2_decap_8 FILLER_11_26 ();
 sg13g2_decap_8 FILLER_11_33 ();
 sg13g2_decap_8 FILLER_11_40 ();
 sg13g2_decap_8 FILLER_11_47 ();
 sg13g2_decap_4 FILLER_11_54 ();
 sg13g2_fill_1 FILLER_11_58 ();
 sg13g2_decap_8 FILLER_11_68 ();
 sg13g2_decap_8 FILLER_11_75 ();
 sg13g2_decap_8 FILLER_11_82 ();
 sg13g2_decap_8 FILLER_11_89 ();
 sg13g2_decap_8 FILLER_11_96 ();
 sg13g2_decap_8 FILLER_11_103 ();
 sg13g2_decap_8 FILLER_11_110 ();
 sg13g2_decap_8 FILLER_11_117 ();
 sg13g2_decap_8 FILLER_11_124 ();
 sg13g2_decap_8 FILLER_11_131 ();
 sg13g2_decap_8 FILLER_11_138 ();
 sg13g2_decap_8 FILLER_11_145 ();
 sg13g2_decap_8 FILLER_11_152 ();
 sg13g2_decap_8 FILLER_11_159 ();
 sg13g2_decap_8 FILLER_11_166 ();
 sg13g2_decap_8 FILLER_11_173 ();
 sg13g2_decap_8 FILLER_11_180 ();
 sg13g2_decap_8 FILLER_11_187 ();
 sg13g2_decap_8 FILLER_11_194 ();
 sg13g2_decap_4 FILLER_11_201 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_fill_1 FILLER_11_224 ();
 sg13g2_fill_2 FILLER_11_255 ();
 sg13g2_decap_8 FILLER_11_309 ();
 sg13g2_decap_4 FILLER_11_316 ();
 sg13g2_decap_8 FILLER_11_372 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_9 ();
 sg13g2_decap_4 FILLER_12_36 ();
 sg13g2_fill_1 FILLER_12_40 ();
 sg13g2_decap_8 FILLER_12_80 ();
 sg13g2_fill_2 FILLER_12_87 ();
 sg13g2_fill_1 FILLER_12_89 ();
 sg13g2_decap_4 FILLER_12_102 ();
 sg13g2_fill_2 FILLER_12_106 ();
 sg13g2_decap_4 FILLER_12_117 ();
 sg13g2_fill_1 FILLER_12_121 ();
 sg13g2_decap_8 FILLER_12_148 ();
 sg13g2_decap_4 FILLER_12_155 ();
 sg13g2_decap_8 FILLER_12_167 ();
 sg13g2_decap_8 FILLER_12_226 ();
 sg13g2_decap_4 FILLER_12_233 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_fill_2 FILLER_12_256 ();
 sg13g2_fill_1 FILLER_12_258 ();
 sg13g2_decap_8 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_274 ();
 sg13g2_decap_8 FILLER_12_288 ();
 sg13g2_decap_4 FILLER_12_295 ();
 sg13g2_fill_1 FILLER_12_299 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_fill_2 FILLER_12_315 ();
 sg13g2_fill_1 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_fill_2 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_fill_2 FILLER_12_361 ();
 sg13g2_fill_1 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_decap_8 FILLER_13_61 ();
 sg13g2_fill_1 FILLER_13_93 ();
 sg13g2_decap_4 FILLER_13_120 ();
 sg13g2_decap_4 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_180 ();
 sg13g2_decap_8 FILLER_13_187 ();
 sg13g2_decap_8 FILLER_13_194 ();
 sg13g2_decap_8 FILLER_13_201 ();
 sg13g2_decap_8 FILLER_13_208 ();
 sg13g2_decap_8 FILLER_13_215 ();
 sg13g2_decap_4 FILLER_13_222 ();
 sg13g2_fill_1 FILLER_13_226 ();
 sg13g2_fill_2 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_290 ();
 sg13g2_fill_2 FILLER_13_297 ();
 sg13g2_fill_1 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_334 ();
 sg13g2_decap_4 FILLER_13_341 ();
 sg13g2_fill_2 FILLER_13_345 ();
 sg13g2_fill_2 FILLER_13_350 ();
 sg13g2_decap_4 FILLER_13_361 ();
 sg13g2_fill_2 FILLER_13_365 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_47 ();
 sg13g2_fill_1 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_92 ();
 sg13g2_decap_8 FILLER_14_103 ();
 sg13g2_fill_2 FILLER_14_110 ();
 sg13g2_fill_1 FILLER_14_112 ();
 sg13g2_decap_4 FILLER_14_123 ();
 sg13g2_fill_1 FILLER_14_127 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_fill_1 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_220 ();
 sg13g2_decap_8 FILLER_14_235 ();
 sg13g2_decap_4 FILLER_14_242 ();
 sg13g2_fill_1 FILLER_14_246 ();
 sg13g2_fill_1 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_279 ();
 sg13g2_decap_8 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_307 ();
 sg13g2_decap_4 FILLER_14_314 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_decap_4 FILLER_14_327 ();
 sg13g2_fill_1 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_fill_1 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_20 ();
 sg13g2_decap_4 FILLER_15_30 ();
 sg13g2_decap_4 FILLER_15_51 ();
 sg13g2_fill_2 FILLER_15_64 ();
 sg13g2_fill_1 FILLER_15_66 ();
 sg13g2_decap_8 FILLER_15_72 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_fill_2 FILLER_15_116 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_4 FILLER_15_151 ();
 sg13g2_fill_1 FILLER_15_155 ();
 sg13g2_fill_2 FILLER_15_163 ();
 sg13g2_decap_4 FILLER_15_192 ();
 sg13g2_fill_1 FILLER_15_200 ();
 sg13g2_decap_4 FILLER_15_241 ();
 sg13g2_fill_2 FILLER_15_245 ();
 sg13g2_fill_2 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_4 FILLER_15_266 ();
 sg13g2_fill_1 FILLER_15_314 ();
 sg13g2_fill_2 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_351 ();
 sg13g2_decap_4 FILLER_15_358 ();
 sg13g2_fill_2 FILLER_15_362 ();
 sg13g2_fill_2 FILLER_15_369 ();
 sg13g2_fill_1 FILLER_15_371 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_9 ();
 sg13g2_decap_4 FILLER_16_36 ();
 sg13g2_fill_2 FILLER_16_40 ();
 sg13g2_fill_2 FILLER_16_108 ();
 sg13g2_fill_1 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_130 ();
 sg13g2_fill_2 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_decap_4 FILLER_16_172 ();
 sg13g2_fill_2 FILLER_16_176 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_decap_4 FILLER_16_221 ();
 sg13g2_decap_4 FILLER_16_236 ();
 sg13g2_fill_2 FILLER_16_240 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_fill_1 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_296 ();
 sg13g2_fill_1 FILLER_16_307 ();
 sg13g2_fill_2 FILLER_16_341 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_fill_2 FILLER_16_388 ();
 sg13g2_fill_1 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_11 ();
 sg13g2_decap_8 FILLER_17_22 ();
 sg13g2_decap_8 FILLER_17_29 ();
 sg13g2_fill_2 FILLER_17_36 ();
 sg13g2_fill_1 FILLER_17_38 ();
 sg13g2_fill_2 FILLER_17_43 ();
 sg13g2_fill_2 FILLER_17_58 ();
 sg13g2_fill_1 FILLER_17_60 ();
 sg13g2_fill_2 FILLER_17_67 ();
 sg13g2_fill_2 FILLER_17_113 ();
 sg13g2_decap_8 FILLER_17_146 ();
 sg13g2_decap_8 FILLER_17_153 ();
 sg13g2_decap_8 FILLER_17_160 ();
 sg13g2_fill_1 FILLER_17_167 ();
 sg13g2_decap_8 FILLER_17_176 ();
 sg13g2_decap_8 FILLER_17_183 ();
 sg13g2_decap_8 FILLER_17_190 ();
 sg13g2_fill_2 FILLER_17_197 ();
 sg13g2_fill_1 FILLER_17_199 ();
 sg13g2_decap_4 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_230 ();
 sg13g2_decap_4 FILLER_17_240 ();
 sg13g2_fill_1 FILLER_17_244 ();
 sg13g2_decap_4 FILLER_17_251 ();
 sg13g2_fill_2 FILLER_17_255 ();
 sg13g2_decap_4 FILLER_17_260 ();
 sg13g2_fill_2 FILLER_17_264 ();
 sg13g2_fill_1 FILLER_17_347 ();
 sg13g2_fill_2 FILLER_17_378 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_4 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_32 ();
 sg13g2_fill_1 FILLER_18_79 ();
 sg13g2_fill_1 FILLER_18_94 ();
 sg13g2_decap_4 FILLER_18_115 ();
 sg13g2_decap_8 FILLER_18_124 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_152 ();
 sg13g2_fill_1 FILLER_18_154 ();
 sg13g2_decap_4 FILLER_18_172 ();
 sg13g2_fill_1 FILLER_18_176 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_217 ();
 sg13g2_fill_1 FILLER_18_245 ();
 sg13g2_fill_2 FILLER_18_274 ();
 sg13g2_fill_2 FILLER_18_284 ();
 sg13g2_fill_1 FILLER_18_290 ();
 sg13g2_fill_2 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_369 ();
 sg13g2_fill_2 FILLER_18_383 ();
 sg13g2_fill_1 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_24 ();
 sg13g2_decap_8 FILLER_19_31 ();
 sg13g2_decap_8 FILLER_19_48 ();
 sg13g2_decap_8 FILLER_19_55 ();
 sg13g2_fill_1 FILLER_19_76 ();
 sg13g2_fill_2 FILLER_19_90 ();
 sg13g2_fill_1 FILLER_19_92 ();
 sg13g2_decap_8 FILLER_19_100 ();
 sg13g2_decap_4 FILLER_19_107 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_decap_4 FILLER_19_117 ();
 sg13g2_fill_2 FILLER_19_121 ();
 sg13g2_decap_8 FILLER_19_142 ();
 sg13g2_fill_1 FILLER_19_149 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_190 ();
 sg13g2_fill_2 FILLER_19_197 ();
 sg13g2_decap_8 FILLER_19_213 ();
 sg13g2_decap_8 FILLER_19_229 ();
 sg13g2_decap_8 FILLER_19_249 ();
 sg13g2_fill_1 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_fill_2 FILLER_19_304 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_fill_2 FILLER_19_333 ();
 sg13g2_fill_2 FILLER_19_340 ();
 sg13g2_fill_2 FILLER_19_359 ();
 sg13g2_decap_4 FILLER_19_365 ();
 sg13g2_fill_2 FILLER_19_369 ();
 sg13g2_fill_2 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_37 ();
 sg13g2_fill_1 FILLER_20_39 ();
 sg13g2_decap_4 FILLER_20_49 ();
 sg13g2_fill_2 FILLER_20_60 ();
 sg13g2_fill_1 FILLER_20_62 ();
 sg13g2_decap_4 FILLER_20_92 ();
 sg13g2_decap_4 FILLER_20_121 ();
 sg13g2_fill_1 FILLER_20_125 ();
 sg13g2_fill_2 FILLER_20_143 ();
 sg13g2_fill_1 FILLER_20_145 ();
 sg13g2_fill_2 FILLER_20_166 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_fill_2 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_225 ();
 sg13g2_fill_2 FILLER_20_242 ();
 sg13g2_fill_1 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_276 ();
 sg13g2_decap_8 FILLER_20_282 ();
 sg13g2_decap_8 FILLER_20_289 ();
 sg13g2_fill_2 FILLER_20_296 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_fill_2 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_310 ();
 sg13g2_fill_1 FILLER_20_316 ();
 sg13g2_decap_4 FILLER_20_322 ();
 sg13g2_fill_2 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_367 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_15 ();
 sg13g2_decap_8 FILLER_21_22 ();
 sg13g2_fill_2 FILLER_21_29 ();
 sg13g2_decap_8 FILLER_21_40 ();
 sg13g2_decap_8 FILLER_21_47 ();
 sg13g2_fill_1 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_89 ();
 sg13g2_fill_2 FILLER_21_95 ();
 sg13g2_fill_1 FILLER_21_97 ();
 sg13g2_decap_8 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_116 ();
 sg13g2_fill_2 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_125 ();
 sg13g2_fill_2 FILLER_21_135 ();
 sg13g2_decap_8 FILLER_21_145 ();
 sg13g2_decap_8 FILLER_21_152 ();
 sg13g2_decap_8 FILLER_21_159 ();
 sg13g2_decap_8 FILLER_21_166 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_4 FILLER_21_189 ();
 sg13g2_fill_2 FILLER_21_212 ();
 sg13g2_decap_4 FILLER_21_219 ();
 sg13g2_fill_2 FILLER_21_223 ();
 sg13g2_fill_2 FILLER_21_233 ();
 sg13g2_decap_4 FILLER_21_245 ();
 sg13g2_fill_1 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_decap_4 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_fill_2 FILLER_21_329 ();
 sg13g2_decap_4 FILLER_21_336 ();
 sg13g2_decap_4 FILLER_21_354 ();
 sg13g2_fill_2 FILLER_21_358 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_45 ();
 sg13g2_fill_2 FILLER_22_52 ();
 sg13g2_fill_1 FILLER_22_59 ();
 sg13g2_fill_2 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_67 ();
 sg13g2_fill_1 FILLER_22_77 ();
 sg13g2_fill_2 FILLER_22_88 ();
 sg13g2_fill_1 FILLER_22_90 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_4 FILLER_22_142 ();
 sg13g2_fill_1 FILLER_22_163 ();
 sg13g2_decap_4 FILLER_22_169 ();
 sg13g2_decap_4 FILLER_22_178 ();
 sg13g2_decap_8 FILLER_22_193 ();
 sg13g2_fill_2 FILLER_22_200 ();
 sg13g2_fill_2 FILLER_22_207 ();
 sg13g2_decap_4 FILLER_22_214 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_decap_4 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_234 ();
 sg13g2_decap_4 FILLER_22_251 ();
 sg13g2_decap_4 FILLER_22_259 ();
 sg13g2_fill_2 FILLER_22_263 ();
 sg13g2_fill_2 FILLER_22_274 ();
 sg13g2_fill_1 FILLER_22_276 ();
 sg13g2_decap_8 FILLER_22_282 ();
 sg13g2_decap_8 FILLER_22_289 ();
 sg13g2_decap_8 FILLER_22_296 ();
 sg13g2_decap_8 FILLER_22_303 ();
 sg13g2_fill_1 FILLER_22_335 ();
 sg13g2_fill_2 FILLER_22_351 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_fill_2 FILLER_22_385 ();
 sg13g2_fill_1 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_14 ();
 sg13g2_fill_1 FILLER_23_16 ();
 sg13g2_decap_4 FILLER_23_26 ();
 sg13g2_fill_2 FILLER_23_40 ();
 sg13g2_fill_1 FILLER_23_48 ();
 sg13g2_fill_2 FILLER_23_66 ();
 sg13g2_fill_2 FILLER_23_74 ();
 sg13g2_fill_1 FILLER_23_76 ();
 sg13g2_decap_4 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_87 ();
 sg13g2_decap_8 FILLER_23_92 ();
 sg13g2_fill_2 FILLER_23_99 ();
 sg13g2_decap_8 FILLER_23_110 ();
 sg13g2_decap_8 FILLER_23_117 ();
 sg13g2_fill_1 FILLER_23_124 ();
 sg13g2_decap_8 FILLER_23_131 ();
 sg13g2_decap_8 FILLER_23_138 ();
 sg13g2_decap_4 FILLER_23_145 ();
 sg13g2_fill_2 FILLER_23_156 ();
 sg13g2_fill_1 FILLER_23_158 ();
 sg13g2_decap_4 FILLER_23_171 ();
 sg13g2_fill_1 FILLER_23_195 ();
 sg13g2_decap_4 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_205 ();
 sg13g2_fill_1 FILLER_23_215 ();
 sg13g2_fill_1 FILLER_23_225 ();
 sg13g2_fill_2 FILLER_23_234 ();
 sg13g2_fill_2 FILLER_23_240 ();
 sg13g2_decap_8 FILLER_23_247 ();
 sg13g2_decap_8 FILLER_23_254 ();
 sg13g2_fill_2 FILLER_23_261 ();
 sg13g2_fill_2 FILLER_23_273 ();
 sg13g2_fill_1 FILLER_23_275 ();
 sg13g2_decap_8 FILLER_23_307 ();
 sg13g2_decap_4 FILLER_23_314 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_decap_4 FILLER_23_334 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_356 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_decap_4 FILLER_24_43 ();
 sg13g2_decap_8 FILLER_24_51 ();
 sg13g2_fill_1 FILLER_24_58 ();
 sg13g2_fill_2 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_97 ();
 sg13g2_fill_1 FILLER_24_111 ();
 sg13g2_fill_2 FILLER_24_153 ();
 sg13g2_fill_1 FILLER_24_160 ();
 sg13g2_decap_8 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_decap_8 FILLER_24_191 ();
 sg13g2_decap_8 FILLER_24_198 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_fill_2 FILLER_24_219 ();
 sg13g2_decap_4 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_235 ();
 sg13g2_decap_4 FILLER_24_241 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_decap_4 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_fill_2 FILLER_24_321 ();
 sg13g2_fill_1 FILLER_24_330 ();
 sg13g2_decap_4 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_4 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_28 ();
 sg13g2_decap_4 FILLER_25_66 ();
 sg13g2_fill_1 FILLER_25_70 ();
 sg13g2_decap_4 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_88 ();
 sg13g2_fill_2 FILLER_25_95 ();
 sg13g2_fill_1 FILLER_25_97 ();
 sg13g2_decap_8 FILLER_25_102 ();
 sg13g2_decap_8 FILLER_25_109 ();
 sg13g2_fill_2 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_135 ();
 sg13g2_decap_8 FILLER_25_142 ();
 sg13g2_decap_8 FILLER_25_149 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_fill_2 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_173 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_fill_2 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_201 ();
 sg13g2_decap_4 FILLER_25_216 ();
 sg13g2_fill_2 FILLER_25_220 ();
 sg13g2_decap_4 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_239 ();
 sg13g2_fill_2 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_4 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_307 ();
 sg13g2_decap_4 FILLER_25_314 ();
 sg13g2_decap_4 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_353 ();
 sg13g2_fill_1 FILLER_25_382 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_fill_2 FILLER_26_31 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_decap_4 FILLER_26_73 ();
 sg13g2_fill_1 FILLER_26_86 ();
 sg13g2_decap_4 FILLER_26_100 ();
 sg13g2_fill_2 FILLER_26_104 ();
 sg13g2_decap_4 FILLER_26_114 ();
 sg13g2_fill_1 FILLER_26_118 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_193 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_decap_4 FILLER_26_231 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_decap_4 FILLER_26_253 ();
 sg13g2_fill_1 FILLER_26_257 ();
 sg13g2_fill_2 FILLER_26_267 ();
 sg13g2_fill_1 FILLER_26_269 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_decap_4 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_313 ();
 sg13g2_fill_2 FILLER_26_330 ();
 sg13g2_fill_1 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_359 ();
 sg13g2_decap_4 FILLER_26_366 ();
 sg13g2_fill_1 FILLER_26_370 ();
 sg13g2_fill_1 FILLER_26_375 ();
 sg13g2_fill_2 FILLER_26_380 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_18 ();
 sg13g2_decap_4 FILLER_27_29 ();
 sg13g2_decap_4 FILLER_27_47 ();
 sg13g2_fill_2 FILLER_27_94 ();
 sg13g2_fill_1 FILLER_27_96 ();
 sg13g2_fill_1 FILLER_27_123 ();
 sg13g2_fill_2 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_138 ();
 sg13g2_decap_8 FILLER_27_148 ();
 sg13g2_fill_1 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_169 ();
 sg13g2_fill_1 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_fill_2 FILLER_27_222 ();
 sg13g2_decap_8 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_fill_2 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_decap_4 FILLER_27_266 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_291 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_fill_2 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_338 ();
 sg13g2_fill_2 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_fill_2 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_fill_1 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_41 ();
 sg13g2_decap_8 FILLER_28_52 ();
 sg13g2_fill_2 FILLER_28_59 ();
 sg13g2_fill_1 FILLER_28_66 ();
 sg13g2_decap_4 FILLER_28_90 ();
 sg13g2_decap_8 FILLER_28_115 ();
 sg13g2_decap_4 FILLER_28_122 ();
 sg13g2_decap_8 FILLER_28_134 ();
 sg13g2_decap_8 FILLER_28_141 ();
 sg13g2_decap_4 FILLER_28_148 ();
 sg13g2_fill_2 FILLER_28_152 ();
 sg13g2_decap_8 FILLER_28_159 ();
 sg13g2_decap_4 FILLER_28_202 ();
 sg13g2_decap_4 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_223 ();
 sg13g2_fill_2 FILLER_28_230 ();
 sg13g2_fill_2 FILLER_28_249 ();
 sg13g2_decap_4 FILLER_28_261 ();
 sg13g2_fill_2 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_298 ();
 sg13g2_fill_2 FILLER_28_305 ();
 sg13g2_decap_8 FILLER_28_311 ();
 sg13g2_fill_2 FILLER_28_318 ();
 sg13g2_decap_8 FILLER_28_328 ();
 sg13g2_fill_2 FILLER_28_335 ();
 sg13g2_fill_2 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_348 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_366 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_43 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_decap_4 FILLER_29_59 ();
 sg13g2_decap_4 FILLER_29_80 ();
 sg13g2_fill_2 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_162 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_decap_8 FILLER_29_176 ();
 sg13g2_decap_4 FILLER_29_183 ();
 sg13g2_fill_2 FILLER_29_187 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_fill_2 FILLER_29_205 ();
 sg13g2_fill_1 FILLER_29_207 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_270 ();
 sg13g2_fill_1 FILLER_29_272 ();
 sg13g2_fill_2 FILLER_29_289 ();
 sg13g2_fill_1 FILLER_29_291 ();
 sg13g2_decap_4 FILLER_29_298 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_fill_2 FILLER_29_352 ();
 sg13g2_fill_1 FILLER_29_354 ();
 sg13g2_decap_4 FILLER_29_375 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_25 ();
 sg13g2_fill_2 FILLER_30_57 ();
 sg13g2_decap_4 FILLER_30_68 ();
 sg13g2_fill_2 FILLER_30_72 ();
 sg13g2_fill_2 FILLER_30_82 ();
 sg13g2_fill_2 FILLER_30_101 ();
 sg13g2_fill_1 FILLER_30_103 ();
 sg13g2_decap_4 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_116 ();
 sg13g2_decap_8 FILLER_30_131 ();
 sg13g2_decap_4 FILLER_30_138 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_decap_4 FILLER_30_185 ();
 sg13g2_fill_2 FILLER_30_189 ();
 sg13g2_decap_4 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_fill_2 FILLER_30_228 ();
 sg13g2_fill_1 FILLER_30_230 ();
 sg13g2_decap_4 FILLER_30_241 ();
 sg13g2_fill_1 FILLER_30_255 ();
 sg13g2_fill_2 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_282 ();
 sg13g2_fill_2 FILLER_30_297 ();
 sg13g2_fill_1 FILLER_30_299 ();
 sg13g2_fill_2 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_316 ();
 sg13g2_fill_2 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_345 ();
 sg13g2_fill_1 FILLER_30_352 ();
 sg13g2_fill_2 FILLER_30_361 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_decap_8 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_42 ();
 sg13g2_fill_1 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_101 ();
 sg13g2_fill_1 FILLER_31_134 ();
 sg13g2_fill_2 FILLER_31_166 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_fill_2 FILLER_31_220 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_decap_4 FILLER_31_229 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_decap_8 FILLER_31_254 ();
 sg13g2_decap_8 FILLER_31_261 ();
 sg13g2_fill_2 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_4 FILLER_32_105 ();
 sg13g2_decap_4 FILLER_32_123 ();
 sg13g2_fill_2 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_185 ();
 sg13g2_fill_2 FILLER_32_192 ();
 sg13g2_fill_1 FILLER_32_194 ();
 sg13g2_fill_2 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_fill_2 FILLER_32_214 ();
 sg13g2_decap_4 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_235 ();
 sg13g2_fill_1 FILLER_32_245 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_decap_4 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_decap_8 FILLER_32_325 ();
 sg13g2_fill_2 FILLER_32_332 ();
 sg13g2_fill_1 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_fill_2 FILLER_32_350 ();
 sg13g2_fill_1 FILLER_32_352 ();
 sg13g2_fill_2 FILLER_32_356 ();
 sg13g2_decap_4 FILLER_32_376 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_fill_2 FILLER_33_84 ();
 sg13g2_fill_2 FILLER_33_112 ();
 sg13g2_fill_1 FILLER_33_114 ();
 sg13g2_fill_2 FILLER_33_149 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_decap_4 FILLER_33_193 ();
 sg13g2_fill_1 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_208 ();
 sg13g2_fill_1 FILLER_33_228 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_decap_8 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_289 ();
 sg13g2_fill_1 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_296 ();
 sg13g2_decap_8 FILLER_33_303 ();
 sg13g2_decap_4 FILLER_33_310 ();
 sg13g2_fill_1 FILLER_33_355 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_4 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_81 ();
 sg13g2_fill_2 FILLER_34_111 ();
 sg13g2_fill_1 FILLER_34_113 ();
 sg13g2_fill_2 FILLER_34_132 ();
 sg13g2_fill_2 FILLER_34_139 ();
 sg13g2_fill_1 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_decap_4 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_194 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_decap_8 FILLER_34_233 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_decap_4 FILLER_34_246 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_4 FILLER_34_266 ();
 sg13g2_fill_2 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_fill_2 FILLER_34_284 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_fill_2 FILLER_34_292 ();
 sg13g2_fill_1 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_309 ();
 sg13g2_decap_4 FILLER_34_316 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_fill_2 FILLER_34_343 ();
 sg13g2_fill_1 FILLER_34_345 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_fill_1 FILLER_34_365 ();
 sg13g2_decap_8 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_34_381 ();
 sg13g2_decap_4 FILLER_34_388 ();
 sg13g2_fill_1 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_4 FILLER_35_98 ();
 sg13g2_fill_2 FILLER_35_102 ();
 sg13g2_fill_2 FILLER_35_113 ();
 sg13g2_fill_1 FILLER_35_115 ();
 sg13g2_decap_8 FILLER_35_174 ();
 sg13g2_decap_8 FILLER_35_181 ();
 sg13g2_fill_2 FILLER_35_188 ();
 sg13g2_fill_1 FILLER_35_190 ();
 sg13g2_decap_8 FILLER_35_206 ();
 sg13g2_decap_8 FILLER_35_213 ();
 sg13g2_decap_4 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_248 ();
 sg13g2_fill_2 FILLER_35_273 ();
 sg13g2_fill_1 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_295 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_decap_8 FILLER_35_330 ();
 sg13g2_decap_4 FILLER_35_337 ();
 sg13g2_decap_4 FILLER_35_374 ();
 sg13g2_fill_2 FILLER_35_378 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_128 ();
 sg13g2_decap_8 FILLER_36_134 ();
 sg13g2_decap_8 FILLER_36_141 ();
 sg13g2_decap_8 FILLER_36_148 ();
 sg13g2_decap_8 FILLER_36_155 ();
 sg13g2_fill_1 FILLER_36_162 ();
 sg13g2_decap_8 FILLER_36_166 ();
 sg13g2_decap_4 FILLER_36_218 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_237 ();
 sg13g2_fill_2 FILLER_36_244 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_decap_8 FILLER_36_270 ();
 sg13g2_decap_8 FILLER_36_277 ();
 sg13g2_decap_4 FILLER_36_284 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_decap_4 FILLER_36_294 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_decap_4 FILLER_36_304 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_361 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_4 FILLER_36_375 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_fill_1 FILLER_37_203 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_258 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_fill_2 FILLER_37_280 ();
 sg13g2_fill_2 FILLER_37_325 ();
 sg13g2_fill_1 FILLER_37_327 ();
 sg13g2_fill_2 FILLER_37_340 ();
 sg13g2_fill_1 FILLER_37_342 ();
 sg13g2_fill_2 FILLER_37_378 ();
 sg13g2_fill_1 FILLER_37_380 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_8 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_107 ();
 sg13g2_fill_1 FILLER_38_111 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_decap_8 FILLER_38_132 ();
 sg13g2_decap_8 FILLER_38_139 ();
 sg13g2_decap_8 FILLER_38_146 ();
 sg13g2_decap_8 FILLER_38_153 ();
 sg13g2_decap_8 FILLER_38_164 ();
 sg13g2_decap_8 FILLER_38_171 ();
 sg13g2_decap_4 FILLER_38_178 ();
 sg13g2_fill_2 FILLER_38_182 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_decap_4 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_228 ();
 sg13g2_decap_4 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_240 ();
 sg13g2_fill_2 FILLER_38_249 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_fill_1 FILLER_38_308 ();
 sg13g2_fill_1 FILLER_38_321 ();
 sg13g2_decap_4 FILLER_38_386 ();
 sg13g2_fill_1 FILLER_38_399 ();
 assign uio_oe[0] = net22;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net23;
 assign uio_oe[4] = net24;
 assign uio_oe[5] = net25;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net26;
 assign uio_out[2] = net13;
 assign uio_out[6] = net14;
 assign uo_out[1] = net15;
 assign uo_out[2] = net16;
 assign uo_out[3] = net17;
 assign uo_out[4] = net18;
 assign uo_out[5] = net19;
 assign uo_out[6] = net20;
 assign uo_out[7] = net21;
endmodule
