module tt_um_ds_comp_adc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire \cic_a.decim_cnt[0] ;
 wire \cic_a.decim_cnt[1] ;
 wire \cic_a.decim_cnt[2] ;
 wire \cic_a.decim_cnt[3] ;
 wire \cic_a.decim_cnt[4] ;
 wire \cic_a.decim_cnt[5] ;
 wire \cic_a.decim_cnt[6] ;
 wire \cic_a.decim_cnt[7] ;
 wire \cic_a.delay[0][0] ;
 wire \cic_a.delay[0][10] ;
 wire \cic_a.delay[0][11] ;
 wire \cic_a.delay[0][12] ;
 wire \cic_a.delay[0][1] ;
 wire \cic_a.delay[0][2] ;
 wire \cic_a.delay[0][3] ;
 wire \cic_a.delay[0][4] ;
 wire \cic_a.delay[0][5] ;
 wire \cic_a.delay[0][6] ;
 wire \cic_a.delay[0][7] ;
 wire \cic_a.delay[0][8] ;
 wire \cic_a.delay[0][9] ;
 wire \cic_a.delay[1][0] ;
 wire \cic_a.delay[1][10] ;
 wire \cic_a.delay[1][11] ;
 wire \cic_a.delay[1][12] ;
 wire \cic_a.delay[1][1] ;
 wire \cic_a.delay[1][2] ;
 wire \cic_a.delay[1][3] ;
 wire \cic_a.delay[1][4] ;
 wire \cic_a.delay[1][5] ;
 wire \cic_a.delay[1][6] ;
 wire \cic_a.delay[1][7] ;
 wire \cic_a.delay[1][8] ;
 wire \cic_a.delay[1][9] ;
 wire \cic_a.delay[2][0] ;
 wire \cic_a.delay[2][10] ;
 wire \cic_a.delay[2][11] ;
 wire \cic_a.delay[2][12] ;
 wire \cic_a.delay[2][1] ;
 wire \cic_a.delay[2][2] ;
 wire \cic_a.delay[2][3] ;
 wire \cic_a.delay[2][4] ;
 wire \cic_a.delay[2][5] ;
 wire \cic_a.delay[2][6] ;
 wire \cic_a.delay[2][7] ;
 wire \cic_a.delay[2][8] ;
 wire \cic_a.delay[2][9] ;
 wire \cic_a.filtered_out[0] ;
 wire \cic_a.filtered_out[10] ;
 wire \cic_a.filtered_out[11] ;
 wire \cic_a.filtered_out[12] ;
 wire \cic_a.filtered_out[1] ;
 wire \cic_a.filtered_out[2] ;
 wire \cic_a.filtered_out[3] ;
 wire \cic_a.filtered_out[4] ;
 wire \cic_a.filtered_out[5] ;
 wire \cic_a.filtered_out[6] ;
 wire \cic_a.filtered_out[7] ;
 wire \cic_a.filtered_out[8] ;
 wire \cic_a.filtered_out[9] ;
 wire \cic_a.integrator[0][0] ;
 wire \cic_a.integrator[0][10] ;
 wire \cic_a.integrator[0][11] ;
 wire \cic_a.integrator[0][12] ;
 wire \cic_a.integrator[0][1] ;
 wire \cic_a.integrator[0][2] ;
 wire \cic_a.integrator[0][3] ;
 wire \cic_a.integrator[0][4] ;
 wire \cic_a.integrator[0][5] ;
 wire \cic_a.integrator[0][6] ;
 wire \cic_a.integrator[0][7] ;
 wire \cic_a.integrator[0][8] ;
 wire \cic_a.integrator[0][9] ;
 wire \cic_a.integrator[1][0] ;
 wire \cic_a.integrator[1][10] ;
 wire \cic_a.integrator[1][11] ;
 wire \cic_a.integrator[1][12] ;
 wire \cic_a.integrator[1][1] ;
 wire \cic_a.integrator[1][2] ;
 wire \cic_a.integrator[1][3] ;
 wire \cic_a.integrator[1][4] ;
 wire \cic_a.integrator[1][5] ;
 wire \cic_a.integrator[1][6] ;
 wire \cic_a.integrator[1][7] ;
 wire \cic_a.integrator[1][8] ;
 wire \cic_a.integrator[1][9] ;
 wire \cic_a.integrator[2][0] ;
 wire \cic_a.integrator[2][10] ;
 wire \cic_a.integrator[2][11] ;
 wire \cic_a.integrator[2][12] ;
 wire \cic_a.integrator[2][1] ;
 wire \cic_a.integrator[2][2] ;
 wire \cic_a.integrator[2][3] ;
 wire \cic_a.integrator[2][4] ;
 wire \cic_a.integrator[2][5] ;
 wire \cic_a.integrator[2][6] ;
 wire \cic_a.integrator[2][7] ;
 wire \cic_a.integrator[2][8] ;
 wire \cic_a.integrator[2][9] ;
 wire \cic_a.pdm_in ;
 wire \cic_a.temp_comb[0][0] ;
 wire \cic_a.temp_comb[0][10] ;
 wire \cic_a.temp_comb[0][11] ;
 wire \cic_a.temp_comb[0][12] ;
 wire \cic_a.temp_comb[0][1] ;
 wire \cic_a.temp_comb[0][2] ;
 wire \cic_a.temp_comb[0][3] ;
 wire \cic_a.temp_comb[0][4] ;
 wire \cic_a.temp_comb[0][5] ;
 wire \cic_a.temp_comb[0][6] ;
 wire \cic_a.temp_comb[0][7] ;
 wire \cic_a.temp_comb[0][8] ;
 wire \cic_a.temp_comb[0][9] ;
 wire \cic_a.temp_comb[1][0] ;
 wire \cic_a.temp_comb[1][10] ;
 wire \cic_a.temp_comb[1][11] ;
 wire \cic_a.temp_comb[1][12] ;
 wire \cic_a.temp_comb[1][1] ;
 wire \cic_a.temp_comb[1][2] ;
 wire \cic_a.temp_comb[1][3] ;
 wire \cic_a.temp_comb[1][4] ;
 wire \cic_a.temp_comb[1][5] ;
 wire \cic_a.temp_comb[1][6] ;
 wire \cic_a.temp_comb[1][7] ;
 wire \cic_a.temp_comb[1][8] ;
 wire \cic_a.temp_comb[1][9] ;
 wire \cic_a.temp_comb[2][0] ;
 wire \cic_a.temp_comb[2][10] ;
 wire \cic_a.temp_comb[2][11] ;
 wire \cic_a.temp_comb[2][12] ;
 wire \cic_a.temp_comb[2][1] ;
 wire \cic_a.temp_comb[2][2] ;
 wire \cic_a.temp_comb[2][3] ;
 wire \cic_a.temp_comb[2][4] ;
 wire \cic_a.temp_comb[2][5] ;
 wire \cic_a.temp_comb[2][6] ;
 wire \cic_a.temp_comb[2][7] ;
 wire \cic_a.temp_comb[2][8] ;
 wire \cic_a.temp_comb[2][9] ;
 wire \cic_a.temp_delay[0][0] ;
 wire \cic_a.temp_delay[0][10] ;
 wire \cic_a.temp_delay[0][11] ;
 wire \cic_a.temp_delay[0][12] ;
 wire \cic_a.temp_delay[0][1] ;
 wire \cic_a.temp_delay[0][2] ;
 wire \cic_a.temp_delay[0][3] ;
 wire \cic_a.temp_delay[0][4] ;
 wire \cic_a.temp_delay[0][5] ;
 wire \cic_a.temp_delay[0][6] ;
 wire \cic_a.temp_delay[0][7] ;
 wire \cic_a.temp_delay[0][8] ;
 wire \cic_a.temp_delay[0][9] ;
 wire \cic_a.temp_delay[1][0] ;
 wire \cic_a.temp_delay[1][10] ;
 wire \cic_a.temp_delay[1][11] ;
 wire \cic_a.temp_delay[1][12] ;
 wire \cic_a.temp_delay[1][1] ;
 wire \cic_a.temp_delay[1][2] ;
 wire \cic_a.temp_delay[1][3] ;
 wire \cic_a.temp_delay[1][4] ;
 wire \cic_a.temp_delay[1][5] ;
 wire \cic_a.temp_delay[1][6] ;
 wire \cic_a.temp_delay[1][7] ;
 wire \cic_a.temp_delay[1][8] ;
 wire \cic_a.temp_delay[1][9] ;
 wire \cic_a.temp_delay[2][0] ;
 wire \cic_a.temp_delay[2][10] ;
 wire \cic_a.temp_delay[2][11] ;
 wire \cic_a.temp_delay[2][12] ;
 wire \cic_a.temp_delay[2][1] ;
 wire \cic_a.temp_delay[2][2] ;
 wire \cic_a.temp_delay[2][3] ;
 wire \cic_a.temp_delay[2][4] ;
 wire \cic_a.temp_delay[2][5] ;
 wire \cic_a.temp_delay[2][6] ;
 wire \cic_a.temp_delay[2][7] ;
 wire \cic_a.temp_delay[2][8] ;
 wire \cic_a.temp_delay[2][9] ;
 wire \cic_b.decim_cnt[0] ;
 wire \cic_b.decim_cnt[1] ;
 wire \cic_b.decim_cnt[2] ;
 wire \cic_b.decim_cnt[3] ;
 wire \cic_b.decim_cnt[4] ;
 wire \cic_b.decim_cnt[5] ;
 wire \cic_b.decim_cnt[6] ;
 wire \cic_b.decim_cnt[7] ;
 wire \cic_b.delay[0][0] ;
 wire \cic_b.delay[0][10] ;
 wire \cic_b.delay[0][11] ;
 wire \cic_b.delay[0][12] ;
 wire \cic_b.delay[0][1] ;
 wire \cic_b.delay[0][2] ;
 wire \cic_b.delay[0][3] ;
 wire \cic_b.delay[0][4] ;
 wire \cic_b.delay[0][5] ;
 wire \cic_b.delay[0][6] ;
 wire \cic_b.delay[0][7] ;
 wire \cic_b.delay[0][8] ;
 wire \cic_b.delay[0][9] ;
 wire \cic_b.delay[1][0] ;
 wire \cic_b.delay[1][10] ;
 wire \cic_b.delay[1][11] ;
 wire \cic_b.delay[1][12] ;
 wire \cic_b.delay[1][1] ;
 wire \cic_b.delay[1][2] ;
 wire \cic_b.delay[1][3] ;
 wire \cic_b.delay[1][4] ;
 wire \cic_b.delay[1][5] ;
 wire \cic_b.delay[1][6] ;
 wire \cic_b.delay[1][7] ;
 wire \cic_b.delay[1][8] ;
 wire \cic_b.delay[1][9] ;
 wire \cic_b.delay[2][0] ;
 wire \cic_b.delay[2][10] ;
 wire \cic_b.delay[2][11] ;
 wire \cic_b.delay[2][12] ;
 wire \cic_b.delay[2][1] ;
 wire \cic_b.delay[2][2] ;
 wire \cic_b.delay[2][3] ;
 wire \cic_b.delay[2][4] ;
 wire \cic_b.delay[2][5] ;
 wire \cic_b.delay[2][6] ;
 wire \cic_b.delay[2][7] ;
 wire \cic_b.delay[2][8] ;
 wire \cic_b.delay[2][9] ;
 wire \cic_b.filtered_out[0] ;
 wire \cic_b.filtered_out[10] ;
 wire \cic_b.filtered_out[11] ;
 wire \cic_b.filtered_out[12] ;
 wire \cic_b.filtered_out[1] ;
 wire \cic_b.filtered_out[2] ;
 wire \cic_b.filtered_out[3] ;
 wire \cic_b.filtered_out[4] ;
 wire \cic_b.filtered_out[5] ;
 wire \cic_b.filtered_out[6] ;
 wire \cic_b.filtered_out[7] ;
 wire \cic_b.filtered_out[8] ;
 wire \cic_b.filtered_out[9] ;
 wire \cic_b.integrator[0][0] ;
 wire \cic_b.integrator[0][10] ;
 wire \cic_b.integrator[0][11] ;
 wire \cic_b.integrator[0][12] ;
 wire \cic_b.integrator[0][1] ;
 wire \cic_b.integrator[0][2] ;
 wire \cic_b.integrator[0][3] ;
 wire \cic_b.integrator[0][4] ;
 wire \cic_b.integrator[0][5] ;
 wire \cic_b.integrator[0][6] ;
 wire \cic_b.integrator[0][7] ;
 wire \cic_b.integrator[0][8] ;
 wire \cic_b.integrator[0][9] ;
 wire \cic_b.integrator[1][0] ;
 wire \cic_b.integrator[1][10] ;
 wire \cic_b.integrator[1][11] ;
 wire \cic_b.integrator[1][12] ;
 wire \cic_b.integrator[1][1] ;
 wire \cic_b.integrator[1][2] ;
 wire \cic_b.integrator[1][3] ;
 wire \cic_b.integrator[1][4] ;
 wire \cic_b.integrator[1][5] ;
 wire \cic_b.integrator[1][6] ;
 wire \cic_b.integrator[1][7] ;
 wire \cic_b.integrator[1][8] ;
 wire \cic_b.integrator[1][9] ;
 wire \cic_b.integrator[2][0] ;
 wire \cic_b.integrator[2][10] ;
 wire \cic_b.integrator[2][11] ;
 wire \cic_b.integrator[2][12] ;
 wire \cic_b.integrator[2][1] ;
 wire \cic_b.integrator[2][2] ;
 wire \cic_b.integrator[2][3] ;
 wire \cic_b.integrator[2][4] ;
 wire \cic_b.integrator[2][5] ;
 wire \cic_b.integrator[2][6] ;
 wire \cic_b.integrator[2][7] ;
 wire \cic_b.integrator[2][8] ;
 wire \cic_b.integrator[2][9] ;
 wire \cic_b.pdm_in ;
 wire \cic_b.temp_comb[0][0] ;
 wire \cic_b.temp_comb[0][10] ;
 wire \cic_b.temp_comb[0][11] ;
 wire \cic_b.temp_comb[0][12] ;
 wire \cic_b.temp_comb[0][1] ;
 wire \cic_b.temp_comb[0][2] ;
 wire \cic_b.temp_comb[0][3] ;
 wire \cic_b.temp_comb[0][4] ;
 wire \cic_b.temp_comb[0][5] ;
 wire \cic_b.temp_comb[0][6] ;
 wire \cic_b.temp_comb[0][7] ;
 wire \cic_b.temp_comb[0][8] ;
 wire \cic_b.temp_comb[0][9] ;
 wire \cic_b.temp_comb[1][0] ;
 wire \cic_b.temp_comb[1][10] ;
 wire \cic_b.temp_comb[1][11] ;
 wire \cic_b.temp_comb[1][12] ;
 wire \cic_b.temp_comb[1][1] ;
 wire \cic_b.temp_comb[1][2] ;
 wire \cic_b.temp_comb[1][3] ;
 wire \cic_b.temp_comb[1][4] ;
 wire \cic_b.temp_comb[1][5] ;
 wire \cic_b.temp_comb[1][6] ;
 wire \cic_b.temp_comb[1][7] ;
 wire \cic_b.temp_comb[1][8] ;
 wire \cic_b.temp_comb[1][9] ;
 wire \cic_b.temp_comb[2][0] ;
 wire \cic_b.temp_comb[2][10] ;
 wire \cic_b.temp_comb[2][11] ;
 wire \cic_b.temp_comb[2][12] ;
 wire \cic_b.temp_comb[2][1] ;
 wire \cic_b.temp_comb[2][2] ;
 wire \cic_b.temp_comb[2][3] ;
 wire \cic_b.temp_comb[2][4] ;
 wire \cic_b.temp_comb[2][5] ;
 wire \cic_b.temp_comb[2][6] ;
 wire \cic_b.temp_comb[2][7] ;
 wire \cic_b.temp_comb[2][8] ;
 wire \cic_b.temp_comb[2][9] ;
 wire \cic_b.temp_delay[0][0] ;
 wire \cic_b.temp_delay[0][10] ;
 wire \cic_b.temp_delay[0][11] ;
 wire \cic_b.temp_delay[0][12] ;
 wire \cic_b.temp_delay[0][1] ;
 wire \cic_b.temp_delay[0][2] ;
 wire \cic_b.temp_delay[0][3] ;
 wire \cic_b.temp_delay[0][4] ;
 wire \cic_b.temp_delay[0][5] ;
 wire \cic_b.temp_delay[0][6] ;
 wire \cic_b.temp_delay[0][7] ;
 wire \cic_b.temp_delay[0][8] ;
 wire \cic_b.temp_delay[0][9] ;
 wire \cic_b.temp_delay[1][0] ;
 wire \cic_b.temp_delay[1][10] ;
 wire \cic_b.temp_delay[1][11] ;
 wire \cic_b.temp_delay[1][12] ;
 wire \cic_b.temp_delay[1][1] ;
 wire \cic_b.temp_delay[1][2] ;
 wire \cic_b.temp_delay[1][3] ;
 wire \cic_b.temp_delay[1][4] ;
 wire \cic_b.temp_delay[1][5] ;
 wire \cic_b.temp_delay[1][6] ;
 wire \cic_b.temp_delay[1][7] ;
 wire \cic_b.temp_delay[1][8] ;
 wire \cic_b.temp_delay[1][9] ;
 wire \cic_b.temp_delay[2][0] ;
 wire \cic_b.temp_delay[2][10] ;
 wire \cic_b.temp_delay[2][11] ;
 wire \cic_b.temp_delay[2][12] ;
 wire \cic_b.temp_delay[2][1] ;
 wire \cic_b.temp_delay[2][2] ;
 wire \cic_b.temp_delay[2][3] ;
 wire \cic_b.temp_delay[2][4] ;
 wire \cic_b.temp_delay[2][5] ;
 wire \cic_b.temp_delay[2][6] ;
 wire \cic_b.temp_delay[2][7] ;
 wire \cic_b.temp_delay[2][8] ;
 wire \cic_b.temp_delay[2][9] ;
 wire pdm_a;
 wire pdm_b;
 wire \serializer_a.bit_cnt[0] ;
 wire \serializer_a.bit_cnt[1] ;
 wire \serializer_a.bit_cnt[2] ;
 wire \serializer_a.bit_cnt[3] ;
 wire \serializer_a.sending ;
 wire \serializer_a.serial_out ;
 wire \serializer_a.shift_reg[0] ;
 wire \serializer_a.shift_reg[10] ;
 wire \serializer_a.shift_reg[11] ;
 wire \serializer_a.shift_reg[1] ;
 wire \serializer_a.shift_reg[2] ;
 wire \serializer_a.shift_reg[3] ;
 wire \serializer_a.shift_reg[4] ;
 wire \serializer_a.shift_reg[5] ;
 wire \serializer_a.shift_reg[6] ;
 wire \serializer_a.shift_reg[7] ;
 wire \serializer_a.shift_reg[8] ;
 wire \serializer_a.shift_reg[9] ;
 wire \serializer_a.valid ;
 wire \serializer_ab_subtr.bit_cnt[0] ;
 wire \serializer_ab_subtr.bit_cnt[1] ;
 wire \serializer_ab_subtr.bit_cnt[2] ;
 wire \serializer_ab_subtr.bit_cnt[3] ;
 wire \serializer_ab_subtr.sending ;
 wire \serializer_ab_subtr.serial_out ;
 wire \serializer_ab_subtr.shift_reg[0] ;
 wire \serializer_ab_subtr.shift_reg[10] ;
 wire \serializer_ab_subtr.shift_reg[11] ;
 wire \serializer_ab_subtr.shift_reg[1] ;
 wire \serializer_ab_subtr.shift_reg[2] ;
 wire \serializer_ab_subtr.shift_reg[3] ;
 wire \serializer_ab_subtr.shift_reg[4] ;
 wire \serializer_ab_subtr.shift_reg[5] ;
 wire \serializer_ab_subtr.shift_reg[6] ;
 wire \serializer_ab_subtr.shift_reg[7] ;
 wire \serializer_ab_subtr.shift_reg[8] ;
 wire \serializer_ab_subtr.shift_reg[9] ;
 wire \serializer_ab_subtr.valid ;
 wire \serializer_b.bit_cnt[0] ;
 wire \serializer_b.bit_cnt[1] ;
 wire \serializer_b.bit_cnt[2] ;
 wire \serializer_b.bit_cnt[3] ;
 wire \serializer_b.sending ;
 wire \serializer_b.serial_out ;
 wire \serializer_b.shift_reg[0] ;
 wire \serializer_b.shift_reg[10] ;
 wire \serializer_b.shift_reg[11] ;
 wire \serializer_b.shift_reg[1] ;
 wire \serializer_b.shift_reg[2] ;
 wire \serializer_b.shift_reg[3] ;
 wire \serializer_b.shift_reg[4] ;
 wire \serializer_b.shift_reg[5] ;
 wire \serializer_b.shift_reg[6] ;
 wire \serializer_b.shift_reg[7] ;
 wire \serializer_b.shift_reg[8] ;
 wire \serializer_b.shift_reg[9] ;
 wire \serializer_b.valid ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_leaf_0_clk;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;

 sg13g2_inv_1 _1724_ (.Y(_0103_),
    .A(net2));
 sg13g2_inv_1 _1725_ (.Y(_0102_),
    .A(net1));
 sg13g2_inv_1 _1726_ (.Y(_0000_),
    .A(net29));
 sg13g2_inv_1 _1727_ (.Y(_1190_),
    .A(\cic_a.decim_cnt[6] ));
 sg13g2_inv_1 _1728_ (.Y(_0008_),
    .A(net24));
 sg13g2_inv_1 _1729_ (.Y(_1191_),
    .A(\cic_b.decim_cnt[6] ));
 sg13g2_inv_1 _1730_ (.Y(_1192_),
    .A(net117));
 sg13g2_inv_1 _1731_ (.Y(_1193_),
    .A(net86));
 sg13g2_inv_1 _1732_ (.Y(_1194_),
    .A(net45));
 sg13g2_inv_1 _1733_ (.Y(_1195_),
    .A(net356));
 sg13g2_inv_1 _1734_ (.Y(_1196_),
    .A(\cic_a.filtered_out[7] ));
 sg13g2_inv_1 _1735_ (.Y(_1197_),
    .A(net209));
 sg13g2_inv_1 _1736_ (.Y(_1198_),
    .A(net260));
 sg13g2_inv_1 _1737_ (.Y(_1199_),
    .A(net203));
 sg13g2_inv_1 _1738_ (.Y(_1200_),
    .A(net207));
 sg13g2_inv_1 _1739_ (.Y(_1201_),
    .A(net83));
 sg13g2_inv_1 _1740_ (.Y(_1202_),
    .A(\cic_b.filtered_out[5] ));
 sg13g2_inv_1 _1741_ (.Y(_1203_),
    .A(net258));
 sg13g2_inv_1 _1742_ (.Y(_1204_),
    .A(net277));
 sg13g2_inv_1 _1743_ (.Y(_1205_),
    .A(net135));
 sg13g2_inv_1 _1744_ (.Y(_1206_),
    .A(net177));
 sg13g2_inv_1 _1745_ (.Y(_1207_),
    .A(net133));
 sg13g2_inv_1 _1746_ (.Y(_1208_),
    .A(net103));
 sg13g2_inv_1 _1747_ (.Y(_1209_),
    .A(net426));
 sg13g2_inv_1 _1748_ (.Y(pdm_a),
    .A(\cic_a.pdm_in ));
 sg13g2_inv_1 _1749_ (.Y(pdm_b),
    .A(\cic_b.pdm_in ));
 sg13g2_inv_1 _1750_ (.Y(_1210_),
    .A(net437));
 sg13g2_inv_1 _1751_ (.Y(_1211_),
    .A(\cic_b.integrator[0][6] ));
 sg13g2_inv_1 _1752_ (.Y(_1212_),
    .A(net634));
 sg13g2_inv_1 _1753_ (.Y(_1213_),
    .A(\cic_a.delay[0][5] ));
 sg13g2_inv_1 _1754_ (.Y(_1214_),
    .A(\cic_a.delay[0][7] ));
 sg13g2_inv_1 _1755_ (.Y(_1215_),
    .A(\cic_a.integrator[2][9] ));
 sg13g2_inv_1 _1756_ (.Y(_1216_),
    .A(net676));
 sg13g2_inv_1 _1757_ (.Y(_1217_),
    .A(net145));
 sg13g2_inv_1 _1758_ (.Y(_1218_),
    .A(\cic_a.delay[1][9] ));
 sg13g2_inv_1 _1759_ (.Y(_1219_),
    .A(\cic_a.integrator[1][9] ));
 sg13g2_inv_1 _1760_ (.Y(_1220_),
    .A(net429));
 sg13g2_inv_1 _1761_ (.Y(_1221_),
    .A(net677));
 sg13g2_inv_1 _1762_ (.Y(_1222_),
    .A(net627));
 sg13g2_inv_1 _1763_ (.Y(_1223_),
    .A(net102));
 sg13g2_inv_1 _1764_ (.Y(_1224_),
    .A(\cic_b.delay[0][5] ));
 sg13g2_inv_1 _1765_ (.Y(_1225_),
    .A(net138));
 sg13g2_inv_1 _1766_ (.Y(_1226_),
    .A(\cic_b.delay[0][9] ));
 sg13g2_inv_1 _1767_ (.Y(_1227_),
    .A(net162));
 sg13g2_inv_1 _1768_ (.Y(_1228_),
    .A(\cic_b.delay[2][9] ));
 sg13g2_inv_1 _1769_ (.Y(_1229_),
    .A(\cic_b.delay[1][4] ));
 sg13g2_inv_1 _1770_ (.Y(_1230_),
    .A(net422));
 sg13g2_inv_1 _1771_ (.Y(_1231_),
    .A(\cic_b.delay[1][9] ));
 sg13g2_inv_1 _1772_ (.Y(_1232_),
    .A(\cic_b.integrator[1][9] ));
 sg13g2_inv_1 _1773_ (.Y(_1233_),
    .A(net125));
 sg13g2_nor2b_1 _1774_ (.A(net546),
    .B_N(net3),
    .Y(_0017_));
 sg13g2_nand2b_1 _1775_ (.Y(_1234_),
    .B(net3),
    .A_N(net540));
 sg13g2_inv_1 _1776_ (.Y(_0019_),
    .A(net537));
 sg13g2_nor2b_1 _1777_ (.A(net703),
    .B_N(net3),
    .Y(_0021_));
 sg13g2_xor2_1 _1778_ (.B(net29),
    .A(net68),
    .X(_0001_));
 sg13g2_and3_2 _1779_ (.X(_1235_),
    .A(net68),
    .B(net29),
    .C(net30));
 sg13g2_a21oi_1 _1780_ (.A1(\cic_a.decim_cnt[1] ),
    .A2(net29),
    .Y(_1236_),
    .B1(net30));
 sg13g2_nor2_1 _1781_ (.A(_1235_),
    .B(net31),
    .Y(_0002_));
 sg13g2_nand2b_1 _1782_ (.Y(_1237_),
    .B(_1235_),
    .A_N(net652));
 sg13g2_nor4_1 _1783_ (.A(\cic_a.decim_cnt[5] ),
    .B(\cic_a.decim_cnt[4] ),
    .C(\cic_a.decim_cnt[7] ),
    .D(\cic_a.decim_cnt[6] ),
    .Y(_1238_));
 sg13g2_nor2b_1 _1784_ (.A(_1237_),
    .B_N(_1238_),
    .Y(_1239_));
 sg13g2_nand2b_1 _1785_ (.Y(_1240_),
    .B(net652),
    .A_N(_1235_));
 sg13g2_a21oi_1 _1786_ (.A1(_1237_),
    .A2(_1240_),
    .Y(_0003_),
    .B1(net503));
 sg13g2_nand3_1 _1787_ (.B(net707),
    .C(_1235_),
    .A(net652),
    .Y(_1241_));
 sg13g2_a21o_1 _1788_ (.A2(_1235_),
    .A1(net652),
    .B1(net707),
    .X(_1242_));
 sg13g2_and2_1 _1789_ (.A(_1241_),
    .B(_1242_),
    .X(_0004_));
 sg13g2_nand4_1 _1790_ (.B(\cic_a.decim_cnt[5] ),
    .C(\cic_a.decim_cnt[4] ),
    .A(\cic_a.decim_cnt[3] ),
    .Y(_1243_),
    .D(_1235_));
 sg13g2_xnor2_1 _1791_ (.Y(_0005_),
    .A(net291),
    .B(_1241_));
 sg13g2_nor2_1 _1792_ (.A(_1190_),
    .B(_1243_),
    .Y(_1244_));
 sg13g2_xnor2_1 _1793_ (.Y(_0006_),
    .A(net244),
    .B(_1243_));
 sg13g2_xor2_1 _1794_ (.B(_1244_),
    .A(net56),
    .X(_0007_));
 sg13g2_xor2_1 _1795_ (.B(net24),
    .A(net116),
    .X(_0009_));
 sg13g2_and3_2 _1796_ (.X(_1245_),
    .A(net116),
    .B(net24),
    .C(net60));
 sg13g2_a21oi_1 _1797_ (.A1(\cic_b.decim_cnt[1] ),
    .A2(net24),
    .Y(_1246_),
    .B1(net60));
 sg13g2_nor2_1 _1798_ (.A(_1245_),
    .B(net61),
    .Y(_0010_));
 sg13g2_nand2b_1 _1799_ (.Y(_1247_),
    .B(_1245_),
    .A_N(net670));
 sg13g2_nor4_1 _1800_ (.A(\cic_b.decim_cnt[5] ),
    .B(\cic_b.decim_cnt[4] ),
    .C(\cic_b.decim_cnt[7] ),
    .D(\cic_b.decim_cnt[6] ),
    .Y(_1248_));
 sg13g2_nor2b_2 _1801_ (.A(_1247_),
    .B_N(_1248_),
    .Y(_1249_));
 sg13g2_nand2b_1 _1802_ (.Y(_1250_),
    .B(net670),
    .A_N(_1245_));
 sg13g2_a21oi_1 _1803_ (.A1(_1247_),
    .A2(_1250_),
    .Y(_0011_),
    .B1(net472));
 sg13g2_nand3_1 _1804_ (.B(net708),
    .C(_1245_),
    .A(net670),
    .Y(_1251_));
 sg13g2_a21o_1 _1805_ (.A2(_1245_),
    .A1(net670),
    .B1(net708),
    .X(_1252_));
 sg13g2_and2_1 _1806_ (.A(_1251_),
    .B(_1252_),
    .X(_0012_));
 sg13g2_nand4_1 _1807_ (.B(\cic_b.decim_cnt[5] ),
    .C(\cic_b.decim_cnt[4] ),
    .A(\cic_b.decim_cnt[3] ),
    .Y(_1253_),
    .D(_1245_));
 sg13g2_xnor2_1 _1808_ (.Y(_0013_),
    .A(net334),
    .B(_1251_));
 sg13g2_nor2_1 _1809_ (.A(_1191_),
    .B(_1253_),
    .Y(_1254_));
 sg13g2_xnor2_1 _1810_ (.Y(_0014_),
    .A(net192),
    .B(_1253_));
 sg13g2_xor2_1 _1811_ (.B(_1254_),
    .A(net69),
    .X(_0015_));
 sg13g2_xor2_1 _1812_ (.B(\cic_b.integrator[0][0] ),
    .A(net92),
    .X(_0061_));
 sg13g2_nand3_1 _1813_ (.B(net721),
    .C(net717),
    .A(net92),
    .Y(_1255_));
 sg13g2_a21o_1 _1814_ (.A2(net455),
    .A1(net92),
    .B1(net717),
    .X(_1256_));
 sg13g2_and2_1 _1815_ (.A(_1255_),
    .B(_1256_),
    .X(_0065_));
 sg13g2_nor2_2 _1816_ (.A(_1210_),
    .B(_1255_),
    .Y(_1257_));
 sg13g2_xnor2_1 _1817_ (.Y(_0066_),
    .A(net437),
    .B(_1255_));
 sg13g2_xor2_1 _1818_ (.B(_1257_),
    .A(net693),
    .X(_0067_));
 sg13g2_nand3_1 _1819_ (.B(net729),
    .C(_1257_),
    .A(net693),
    .Y(_1258_));
 sg13g2_a21o_1 _1820_ (.A2(_1257_),
    .A1(net693),
    .B1(net729),
    .X(_1259_));
 sg13g2_and2_1 _1821_ (.A(_1258_),
    .B(_1259_),
    .X(_0068_));
 sg13g2_nand4_1 _1822_ (.B(\cic_b.integrator[0][4] ),
    .C(net625),
    .A(\cic_b.integrator[0][3] ),
    .Y(_1260_),
    .D(_1257_));
 sg13g2_xnor2_1 _1823_ (.Y(_0069_),
    .A(net625),
    .B(_1258_));
 sg13g2_nor2_1 _1824_ (.A(_1211_),
    .B(_1260_),
    .Y(_1261_));
 sg13g2_xnor2_1 _1825_ (.Y(_0070_),
    .A(net690),
    .B(_1260_));
 sg13g2_xor2_1 _1826_ (.B(_1261_),
    .A(net653),
    .X(_0071_));
 sg13g2_nand3_1 _1827_ (.B(net727),
    .C(_1261_),
    .A(\cic_b.integrator[0][7] ),
    .Y(_1262_));
 sg13g2_a21o_1 _1828_ (.A2(_1261_),
    .A1(net653),
    .B1(net727),
    .X(_1263_));
 sg13g2_and2_1 _1829_ (.A(_1262_),
    .B(_1263_),
    .X(_0072_));
 sg13g2_nor2_2 _1830_ (.A(_1212_),
    .B(_1262_),
    .Y(_1264_));
 sg13g2_xnor2_1 _1831_ (.Y(_0073_),
    .A(net634),
    .B(_1262_));
 sg13g2_xor2_1 _1832_ (.B(_1264_),
    .A(net668),
    .X(_0062_));
 sg13g2_nand3_1 _1833_ (.B(net723),
    .C(_1264_),
    .A(net668),
    .Y(_1265_));
 sg13g2_a21o_1 _1834_ (.A2(_1264_),
    .A1(net668),
    .B1(net723),
    .X(_1266_));
 sg13g2_and2_1 _1835_ (.A(_1265_),
    .B(_1266_),
    .X(_0063_));
 sg13g2_xnor2_1 _1836_ (.Y(_0064_),
    .A(net184),
    .B(_1265_));
 sg13g2_nand2_1 _1837_ (.Y(_1267_),
    .A(net712),
    .B(net458));
 sg13g2_nand2_1 _1838_ (.Y(_1268_),
    .A(\cic_a.integrator[2][1] ),
    .B(\cic_a.integrator[1][1] ));
 sg13g2_nor2_1 _1839_ (.A(\cic_a.integrator[2][1] ),
    .B(\cic_a.integrator[1][1] ),
    .Y(_1269_));
 sg13g2_xor2_1 _1840_ (.B(\cic_a.integrator[1][1] ),
    .A(\cic_a.integrator[2][1] ),
    .X(_1270_));
 sg13g2_xnor2_1 _1841_ (.Y(_0052_),
    .A(_1267_),
    .B(_1270_));
 sg13g2_and2_1 _1842_ (.A(\cic_a.integrator[2][2] ),
    .B(net773),
    .X(_1271_));
 sg13g2_or2_1 _1843_ (.X(_1272_),
    .B(net737),
    .A(\cic_a.integrator[2][2] ));
 sg13g2_nand2b_1 _1844_ (.Y(_1273_),
    .B(_1272_),
    .A_N(_1271_));
 sg13g2_o21ai_1 _1845_ (.B1(_1268_),
    .Y(_1274_),
    .A1(_1267_),
    .A2(_1269_));
 sg13g2_xnor2_1 _1846_ (.Y(_0053_),
    .A(_1273_),
    .B(_1274_));
 sg13g2_a21oi_1 _1847_ (.A1(_1272_),
    .A2(_1274_),
    .Y(_1275_),
    .B1(_1271_));
 sg13g2_nand2_1 _1848_ (.Y(_1276_),
    .A(\cic_a.integrator[2][3] ),
    .B(net786));
 sg13g2_xnor2_1 _1849_ (.Y(_1277_),
    .A(net144),
    .B(net735));
 sg13g2_xor2_1 _1850_ (.B(_1277_),
    .A(_1275_),
    .X(_0054_));
 sg13g2_nand2_1 _1851_ (.Y(_1278_),
    .A(\cic_a.integrator[2][4] ),
    .B(net750));
 sg13g2_xor2_1 _1852_ (.B(\cic_a.integrator[1][4] ),
    .A(\cic_a.integrator[2][4] ),
    .X(_1279_));
 sg13g2_o21ai_1 _1853_ (.B1(_1276_),
    .Y(_1280_),
    .A1(_1275_),
    .A2(_1277_));
 sg13g2_nand2_1 _1854_ (.Y(_1281_),
    .A(_1279_),
    .B(_1280_));
 sg13g2_xor2_1 _1855_ (.B(_1280_),
    .A(_1279_),
    .X(_0055_));
 sg13g2_nor2_1 _1856_ (.A(\cic_a.integrator[2][5] ),
    .B(\cic_a.integrator[1][5] ),
    .Y(_1282_));
 sg13g2_nand2_1 _1857_ (.Y(_1283_),
    .A(\cic_a.integrator[2][5] ),
    .B(\cic_a.integrator[1][5] ));
 sg13g2_nor2b_1 _1858_ (.A(_1282_),
    .B_N(_1283_),
    .Y(_1284_));
 sg13g2_nand2_1 _1859_ (.Y(_1285_),
    .A(net751),
    .B(_1281_));
 sg13g2_xor2_1 _1860_ (.B(_1285_),
    .A(_1284_),
    .X(_0056_));
 sg13g2_and2_1 _1861_ (.A(net767),
    .B(net732),
    .X(_1286_));
 sg13g2_xor2_1 _1862_ (.B(net788),
    .A(\cic_a.integrator[2][6] ),
    .X(_1287_));
 sg13g2_inv_1 _1863_ (.Y(_1288_),
    .A(net789));
 sg13g2_o21ai_1 _1864_ (.B1(_1283_),
    .Y(_1289_),
    .A1(_1278_),
    .A2(_1282_));
 sg13g2_nand3_1 _1865_ (.B(_1280_),
    .C(_1284_),
    .A(_1279_),
    .Y(_1290_));
 sg13g2_nand2b_1 _1866_ (.Y(_1291_),
    .B(_1290_),
    .A_N(_1289_));
 sg13g2_xnor2_1 _1867_ (.Y(_0057_),
    .A(_1288_),
    .B(_1291_));
 sg13g2_nand2_1 _1868_ (.Y(_1292_),
    .A(\cic_a.integrator[2][7] ),
    .B(net740));
 sg13g2_xnor2_1 _1869_ (.Y(_1293_),
    .A(\cic_a.integrator[2][7] ),
    .B(net740));
 sg13g2_a21oi_1 _1870_ (.A1(_1287_),
    .A2(_1291_),
    .Y(_1294_),
    .B1(_1286_));
 sg13g2_xor2_1 _1871_ (.B(_1294_),
    .A(_1293_),
    .X(_0058_));
 sg13g2_nand2_1 _1872_ (.Y(_1295_),
    .A(\cic_a.integrator[2][8] ),
    .B(\cic_a.integrator[1][8] ));
 sg13g2_xnor2_1 _1873_ (.Y(_1296_),
    .A(\cic_a.integrator[2][8] ),
    .B(net746));
 sg13g2_o21ai_1 _1874_ (.B1(_1286_),
    .Y(_1297_),
    .A1(\cic_a.integrator[2][7] ),
    .A2(net749));
 sg13g2_nor2_1 _1875_ (.A(_1288_),
    .B(_1293_),
    .Y(_1298_));
 sg13g2_nand2_1 _1876_ (.Y(_1299_),
    .A(_1289_),
    .B(_1298_));
 sg13g2_nand4_1 _1877_ (.B(_1280_),
    .C(_1284_),
    .A(_1279_),
    .Y(_1300_),
    .D(_1298_));
 sg13g2_nand4_1 _1878_ (.B(_1297_),
    .C(_1299_),
    .A(_1292_),
    .Y(_1301_),
    .D(_1300_));
 sg13g2_nand2b_1 _1879_ (.Y(_1302_),
    .B(_1301_),
    .A_N(_1296_));
 sg13g2_xnor2_1 _1880_ (.Y(_0059_),
    .A(_1296_),
    .B(_1301_));
 sg13g2_xnor2_1 _1881_ (.Y(_1303_),
    .A(net724),
    .B(\cic_a.integrator[1][9] ));
 sg13g2_nand2_1 _1882_ (.Y(_1304_),
    .A(_1295_),
    .B(_1302_));
 sg13g2_xnor2_1 _1883_ (.Y(_0060_),
    .A(net725),
    .B(_1304_));
 sg13g2_nor2_1 _1884_ (.A(_1296_),
    .B(_1303_),
    .Y(_1305_));
 sg13g2_a21oi_1 _1885_ (.A1(_1215_),
    .A2(_1219_),
    .Y(_1306_),
    .B1(_1295_));
 sg13g2_a221oi_1 _1886_ (.B2(_1305_),
    .C1(_1306_),
    .B1(_1301_),
    .A1(net769),
    .Y(_1307_),
    .A2(\cic_a.integrator[1][9] ));
 sg13g2_nand2_1 _1887_ (.Y(_1308_),
    .A(net250),
    .B(net754));
 sg13g2_xnor2_1 _1888_ (.Y(_1309_),
    .A(net250),
    .B(net754));
 sg13g2_xor2_1 _1889_ (.B(_1309_),
    .A(_1307_),
    .X(_0049_));
 sg13g2_nor2_1 _1890_ (.A(\cic_a.integrator[2][11] ),
    .B(\cic_a.integrator[1][11] ),
    .Y(_1310_));
 sg13g2_xnor2_1 _1891_ (.Y(_1311_),
    .A(net763),
    .B(net730));
 sg13g2_o21ai_1 _1892_ (.B1(_1308_),
    .Y(_1312_),
    .A1(_1307_),
    .A2(_1309_));
 sg13g2_xnor2_1 _1893_ (.Y(_0050_),
    .A(_1311_),
    .B(_1312_));
 sg13g2_or2_1 _1894_ (.X(_0415_),
    .B(_1311_),
    .A(_1309_));
 sg13g2_nor2_1 _1895_ (.A(_1308_),
    .B(_1310_),
    .Y(_0416_));
 sg13g2_a21oi_1 _1896_ (.A1(\cic_a.integrator[2][11] ),
    .A2(\cic_a.integrator[1][11] ),
    .Y(_0417_),
    .B1(_0416_));
 sg13g2_o21ai_1 _1897_ (.B1(_0417_),
    .Y(_0418_),
    .A1(_1307_),
    .A2(_0415_));
 sg13g2_xnor2_1 _1898_ (.Y(_0419_),
    .A(net701),
    .B(net698));
 sg13g2_xnor2_1 _1899_ (.Y(_0051_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_xor2_1 _1900_ (.B(net458),
    .A(\cic_a.integrator[2][0] ),
    .X(_0048_));
 sg13g2_nand2_1 _1901_ (.Y(_0420_),
    .A(net458),
    .B(net630));
 sg13g2_nand2_1 _1902_ (.Y(_0421_),
    .A(\cic_a.integrator[1][1] ),
    .B(net705));
 sg13g2_nor2_1 _1903_ (.A(\cic_a.integrator[1][1] ),
    .B(net781),
    .Y(_0422_));
 sg13g2_xor2_1 _1904_ (.B(net705),
    .A(\cic_a.integrator[1][1] ),
    .X(_0423_));
 sg13g2_xnor2_1 _1905_ (.Y(_0039_),
    .A(_0420_),
    .B(net706));
 sg13g2_and2_1 _1906_ (.A(net737),
    .B(net429),
    .X(_0424_));
 sg13g2_or2_1 _1907_ (.X(_0425_),
    .B(net429),
    .A(net737));
 sg13g2_nand2b_1 _1908_ (.Y(_0426_),
    .B(_0425_),
    .A_N(_0424_));
 sg13g2_o21ai_1 _1909_ (.B1(_0421_),
    .Y(_0427_),
    .A1(_0420_),
    .A2(_0422_));
 sg13g2_xnor2_1 _1910_ (.Y(_0040_),
    .A(_0426_),
    .B(_0427_));
 sg13g2_a21oi_2 _1911_ (.B1(_0424_),
    .Y(_0428_),
    .A2(_0427_),
    .A1(_0425_));
 sg13g2_nand2_1 _1912_ (.Y(_0429_),
    .A(net735),
    .B(net782));
 sg13g2_xnor2_1 _1913_ (.Y(_0430_),
    .A(net735),
    .B(net683));
 sg13g2_xor2_1 _1914_ (.B(_0430_),
    .A(_0428_),
    .X(_0041_));
 sg13g2_nand2_1 _1915_ (.Y(_0431_),
    .A(net750),
    .B(net720));
 sg13g2_xor2_1 _1916_ (.B(net720),
    .A(\cic_a.integrator[1][4] ),
    .X(_0432_));
 sg13g2_o21ai_1 _1917_ (.B1(_0429_),
    .Y(_0433_),
    .A1(_0428_),
    .A2(_0430_));
 sg13g2_nand2_1 _1918_ (.Y(_0434_),
    .A(_0432_),
    .B(_0433_));
 sg13g2_xor2_1 _1919_ (.B(_0433_),
    .A(_0432_),
    .X(_0042_));
 sg13g2_nor2_1 _1920_ (.A(\cic_a.integrator[1][5] ),
    .B(\cic_a.integrator[0][5] ),
    .Y(_0435_));
 sg13g2_or2_1 _1921_ (.X(_0436_),
    .B(net765),
    .A(\cic_a.integrator[1][5] ));
 sg13g2_nand2_1 _1922_ (.Y(_0437_),
    .A(\cic_a.integrator[1][5] ),
    .B(net765));
 sg13g2_nand2_1 _1923_ (.Y(_0438_),
    .A(net766),
    .B(_0437_));
 sg13g2_nand2_1 _1924_ (.Y(_0439_),
    .A(_0431_),
    .B(_0434_));
 sg13g2_xnor2_1 _1925_ (.Y(_0043_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_nand2_1 _1926_ (.Y(_0440_),
    .A(\cic_a.integrator[1][6] ),
    .B(net677));
 sg13g2_nor2_1 _1927_ (.A(\cic_a.integrator[1][6] ),
    .B(\cic_a.integrator[0][6] ),
    .Y(_0441_));
 sg13g2_xor2_1 _1928_ (.B(net677),
    .A(net732),
    .X(_0442_));
 sg13g2_nand4_1 _1929_ (.B(_0433_),
    .C(_0436_),
    .A(_0432_),
    .Y(_0443_),
    .D(_0437_));
 sg13g2_o21ai_1 _1930_ (.B1(_0437_),
    .Y(_0444_),
    .A1(_0431_),
    .A2(_0435_));
 sg13g2_nor2b_1 _1931_ (.A(_0444_),
    .B_N(_0443_),
    .Y(_0445_));
 sg13g2_xnor2_1 _1932_ (.Y(_0044_),
    .A(_0442_),
    .B(_0445_));
 sg13g2_nand2_1 _1933_ (.Y(_0446_),
    .A(\cic_a.integrator[1][7] ),
    .B(\cic_a.integrator[0][7] ));
 sg13g2_nor2_1 _1934_ (.A(\cic_a.integrator[1][7] ),
    .B(\cic_a.integrator[0][7] ),
    .Y(_0447_));
 sg13g2_xnor2_1 _1935_ (.Y(_0448_),
    .A(net740),
    .B(net688));
 sg13g2_o21ai_1 _1936_ (.B1(_0440_),
    .Y(_0449_),
    .A1(_0441_),
    .A2(_0445_));
 sg13g2_xnor2_1 _1937_ (.Y(_0045_),
    .A(_0448_),
    .B(_0449_));
 sg13g2_o21ai_1 _1938_ (.B1(_0446_),
    .Y(_0450_),
    .A1(_0440_),
    .A2(_0447_));
 sg13g2_nor2_1 _1939_ (.A(_0444_),
    .B(_0450_),
    .Y(_0451_));
 sg13g2_a221oi_1 _1940_ (.B2(_0443_),
    .C1(_0447_),
    .B1(_0451_),
    .A1(_0441_),
    .Y(_0452_),
    .A2(_0446_));
 sg13g2_nand2_1 _1941_ (.Y(_0453_),
    .A(net746),
    .B(net715));
 sg13g2_xor2_1 _1942_ (.B(net715),
    .A(net746),
    .X(_0454_));
 sg13g2_nand2_1 _1943_ (.Y(_0455_),
    .A(_0452_),
    .B(_0454_));
 sg13g2_xor2_1 _1944_ (.B(_0454_),
    .A(_0452_),
    .X(_0046_));
 sg13g2_xor2_1 _1945_ (.B(net627),
    .A(\cic_a.integrator[1][9] ),
    .X(_0456_));
 sg13g2_nand2_1 _1946_ (.Y(_0457_),
    .A(_0453_),
    .B(_0455_));
 sg13g2_xor2_1 _1947_ (.B(_0457_),
    .A(_0456_),
    .X(_0047_));
 sg13g2_and2_1 _1948_ (.A(_0454_),
    .B(_0456_),
    .X(_0458_));
 sg13g2_a21oi_1 _1949_ (.A1(_1219_),
    .A2(_1222_),
    .Y(_0459_),
    .B1(_0453_));
 sg13g2_a221oi_1 _1950_ (.B2(_0458_),
    .C1(_0459_),
    .B1(_0452_),
    .A1(\cic_a.integrator[1][9] ),
    .Y(_0460_),
    .A2(\cic_a.integrator[0][9] ));
 sg13g2_nand2_1 _1951_ (.Y(_0461_),
    .A(\cic_a.integrator[1][10] ),
    .B(net673));
 sg13g2_xnor2_1 _1952_ (.Y(_0462_),
    .A(net754),
    .B(net673));
 sg13g2_xor2_1 _1953_ (.B(_0462_),
    .A(_0460_),
    .X(_0036_));
 sg13g2_nor2_1 _1954_ (.A(\cic_a.integrator[1][11] ),
    .B(\cic_a.integrator[0][11] ),
    .Y(_0463_));
 sg13g2_xnor2_1 _1955_ (.Y(_0464_),
    .A(net730),
    .B(net722));
 sg13g2_o21ai_1 _1956_ (.B1(_0461_),
    .Y(_0465_),
    .A1(_0460_),
    .A2(_0462_));
 sg13g2_xnor2_1 _1957_ (.Y(_0037_),
    .A(_0464_),
    .B(_0465_));
 sg13g2_or2_1 _1958_ (.X(_0466_),
    .B(_0464_),
    .A(_0462_));
 sg13g2_nor2_1 _1959_ (.A(_0461_),
    .B(_0463_),
    .Y(_0467_));
 sg13g2_a21oi_1 _1960_ (.A1(\cic_a.integrator[1][11] ),
    .A2(\cic_a.integrator[0][11] ),
    .Y(_0468_),
    .B1(_0467_));
 sg13g2_o21ai_1 _1961_ (.B1(_0468_),
    .Y(_0469_),
    .A1(_0460_),
    .A2(_0466_));
 sg13g2_xnor2_1 _1962_ (.Y(_0470_),
    .A(net698),
    .B(net100));
 sg13g2_xnor2_1 _1963_ (.Y(_0038_),
    .A(_0469_),
    .B(_0470_));
 sg13g2_xor2_1 _1964_ (.B(net630),
    .A(net458),
    .X(_0035_));
 sg13g2_nand2_1 _1965_ (.Y(_0471_),
    .A(\cic_b.integrator[2][0] ),
    .B(net452));
 sg13g2_nand2_1 _1966_ (.Y(_0472_),
    .A(net352),
    .B(net759));
 sg13g2_nor2_1 _1967_ (.A(\cic_b.integrator[2][1] ),
    .B(\cic_b.integrator[1][1] ),
    .Y(_0473_));
 sg13g2_xor2_1 _1968_ (.B(net710),
    .A(net352),
    .X(_0474_));
 sg13g2_xnor2_1 _1969_ (.Y(_0091_),
    .A(_0471_),
    .B(_0474_));
 sg13g2_and2_1 _1970_ (.A(\cic_b.integrator[2][2] ),
    .B(\cic_b.integrator[1][2] ),
    .X(_0475_));
 sg13g2_or2_1 _1971_ (.X(_0476_),
    .B(\cic_b.integrator[1][2] ),
    .A(\cic_b.integrator[2][2] ));
 sg13g2_nand2b_1 _1972_ (.Y(_0477_),
    .B(_0476_),
    .A_N(_0475_));
 sg13g2_o21ai_1 _1973_ (.B1(_0472_),
    .Y(_0478_),
    .A1(_0471_),
    .A2(_0473_));
 sg13g2_xnor2_1 _1974_ (.Y(_0092_),
    .A(_0477_),
    .B(net760));
 sg13g2_a21o_1 _1975_ (.A2(_0478_),
    .A1(_0476_),
    .B1(_0475_),
    .X(_0479_));
 sg13g2_and2_1 _1976_ (.A(\cic_b.integrator[2][3] ),
    .B(net718),
    .X(_0480_));
 sg13g2_or2_1 _1977_ (.X(_0481_),
    .B(net718),
    .A(net770));
 sg13g2_nand2b_1 _1978_ (.Y(_0482_),
    .B(_0481_),
    .A_N(_0480_));
 sg13g2_xnor2_1 _1979_ (.Y(_0093_),
    .A(_0479_),
    .B(_0482_));
 sg13g2_nand2_1 _1980_ (.Y(_0483_),
    .A(\cic_b.integrator[2][4] ),
    .B(net756));
 sg13g2_xnor2_1 _1981_ (.Y(_0484_),
    .A(net764),
    .B(net756));
 sg13g2_a21o_1 _1982_ (.A2(_0481_),
    .A1(_0479_),
    .B1(_0480_),
    .X(_0485_));
 sg13g2_nand2b_1 _1983_ (.Y(_0486_),
    .B(_0485_),
    .A_N(_0484_));
 sg13g2_xnor2_1 _1984_ (.Y(_0094_),
    .A(_0484_),
    .B(_0485_));
 sg13g2_nor2_1 _1985_ (.A(\cic_b.integrator[2][5] ),
    .B(\cic_b.integrator[1][5] ),
    .Y(_0487_));
 sg13g2_nand2_1 _1986_ (.Y(_0488_),
    .A(\cic_b.integrator[2][5] ),
    .B(\cic_b.integrator[1][5] ));
 sg13g2_nor2b_1 _1987_ (.A(_0487_),
    .B_N(_0488_),
    .Y(_0489_));
 sg13g2_nand2_1 _1988_ (.Y(_0490_),
    .A(net757),
    .B(_0486_));
 sg13g2_xor2_1 _1989_ (.B(_0490_),
    .A(_0489_),
    .X(_0095_));
 sg13g2_nand2_1 _1990_ (.Y(_0491_),
    .A(net748),
    .B(net742));
 sg13g2_nor2_1 _1991_ (.A(\cic_b.integrator[2][6] ),
    .B(net777),
    .Y(_0492_));
 sg13g2_xor2_1 _1992_ (.B(net742),
    .A(net748),
    .X(_0493_));
 sg13g2_nand3b_1 _1993_ (.B(_0485_),
    .C(_0489_),
    .Y(_0494_),
    .A_N(_0484_));
 sg13g2_o21ai_1 _1994_ (.B1(_0488_),
    .Y(_0495_),
    .A1(_0483_),
    .A2(_0487_));
 sg13g2_nor2b_1 _1995_ (.A(_0495_),
    .B_N(_0494_),
    .Y(_0496_));
 sg13g2_xnor2_1 _1996_ (.Y(_0096_),
    .A(_0493_),
    .B(_0496_));
 sg13g2_nor2_1 _1997_ (.A(\cic_b.integrator[2][7] ),
    .B(\cic_b.integrator[1][7] ),
    .Y(_0497_));
 sg13g2_nand2_1 _1998_ (.Y(_0498_),
    .A(\cic_b.integrator[2][7] ),
    .B(net752));
 sg13g2_nand2b_1 _1999_ (.Y(_0499_),
    .B(_0498_),
    .A_N(_0497_));
 sg13g2_o21ai_1 _2000_ (.B1(_0491_),
    .Y(_0500_),
    .A1(_0492_),
    .A2(_0496_));
 sg13g2_xnor2_1 _2001_ (.Y(_0097_),
    .A(_0499_),
    .B(_0500_));
 sg13g2_o21ai_1 _2002_ (.B1(_0498_),
    .Y(_0501_),
    .A1(_0491_),
    .A2(_0497_));
 sg13g2_nor2_1 _2003_ (.A(_0495_),
    .B(_0501_),
    .Y(_0502_));
 sg13g2_a221oi_1 _2004_ (.B2(_0494_),
    .C1(_0497_),
    .B1(_0502_),
    .A1(_0492_),
    .Y(_0503_),
    .A2(_0498_));
 sg13g2_nand2_1 _2005_ (.Y(_0504_),
    .A(\cic_b.integrator[2][8] ),
    .B(net744));
 sg13g2_xor2_1 _2006_ (.B(net744),
    .A(net775),
    .X(_0505_));
 sg13g2_inv_1 _2007_ (.Y(_0506_),
    .A(_0505_));
 sg13g2_nand2_1 _2008_ (.Y(_0507_),
    .A(_0503_),
    .B(_0505_));
 sg13g2_xnor2_1 _2009_ (.Y(_0098_),
    .A(_0503_),
    .B(_0506_));
 sg13g2_xnor2_1 _2010_ (.Y(_0508_),
    .A(net138),
    .B(net738));
 sg13g2_nand2_1 _2011_ (.Y(_0509_),
    .A(net745),
    .B(_0507_));
 sg13g2_xnor2_1 _2012_ (.Y(_0099_),
    .A(_0508_),
    .B(_0509_));
 sg13g2_nand2_1 _2013_ (.Y(_0510_),
    .A(net662),
    .B(net709));
 sg13g2_xnor2_1 _2014_ (.Y(_0511_),
    .A(net662),
    .B(net709));
 sg13g2_a21oi_1 _2015_ (.A1(_1225_),
    .A2(_1232_),
    .Y(_0512_),
    .B1(_0504_));
 sg13g2_nor2_1 _2016_ (.A(_0506_),
    .B(_0508_),
    .Y(_0513_));
 sg13g2_a221oi_1 _2017_ (.B2(_0513_),
    .C1(_0512_),
    .B1(_0503_),
    .A1(\cic_b.integrator[2][9] ),
    .Y(_0514_),
    .A2(\cic_b.integrator[1][9] ));
 sg13g2_xor2_1 _2018_ (.B(_0514_),
    .A(_0511_),
    .X(_0088_));
 sg13g2_nor2_1 _2019_ (.A(\cic_b.integrator[2][11] ),
    .B(\cic_b.integrator[1][11] ),
    .Y(_0515_));
 sg13g2_xnor2_1 _2020_ (.Y(_0516_),
    .A(net127),
    .B(net696));
 sg13g2_o21ai_1 _2021_ (.B1(_0510_),
    .Y(_0517_),
    .A1(_0511_),
    .A2(_0514_));
 sg13g2_xnor2_1 _2022_ (.Y(_0089_),
    .A(_0516_),
    .B(_0517_));
 sg13g2_or2_1 _2023_ (.X(_0518_),
    .B(_0516_),
    .A(_0511_));
 sg13g2_nor2_1 _2024_ (.A(_0510_),
    .B(_0515_),
    .Y(_0519_));
 sg13g2_a21oi_1 _2025_ (.A1(net127),
    .A2(net696),
    .Y(_0520_),
    .B1(_0519_));
 sg13g2_o21ai_1 _2026_ (.B1(net697),
    .Y(_0521_),
    .A1(_0514_),
    .A2(_0518_));
 sg13g2_xnor2_1 _2027_ (.Y(_0522_),
    .A(net353),
    .B(net646));
 sg13g2_xnor2_1 _2028_ (.Y(_0090_),
    .A(_0521_),
    .B(_0522_));
 sg13g2_xor2_1 _2029_ (.B(net452),
    .A(\cic_b.integrator[2][0] ),
    .X(_0087_));
 sg13g2_nand2_1 _2030_ (.Y(_0523_),
    .A(net455),
    .B(net452));
 sg13g2_nand2_1 _2031_ (.Y(_0524_),
    .A(net717),
    .B(net759));
 sg13g2_nor2_1 _2032_ (.A(\cic_b.integrator[0][1] ),
    .B(\cic_b.integrator[1][1] ),
    .Y(_0525_));
 sg13g2_xor2_1 _2033_ (.B(net710),
    .A(net717),
    .X(_0526_));
 sg13g2_xnor2_1 _2034_ (.Y(_0078_),
    .A(_0523_),
    .B(_0526_));
 sg13g2_and2_1 _2035_ (.A(net437),
    .B(\cic_b.integrator[1][2] ),
    .X(_0527_));
 sg13g2_or2_1 _2036_ (.X(_0528_),
    .B(net776),
    .A(net437));
 sg13g2_nand2b_1 _2037_ (.Y(_0529_),
    .B(_0528_),
    .A_N(_0527_));
 sg13g2_o21ai_1 _2038_ (.B1(_0524_),
    .Y(_0530_),
    .A1(_0523_),
    .A2(_0525_));
 sg13g2_xnor2_1 _2039_ (.Y(_0079_),
    .A(_0529_),
    .B(_0530_));
 sg13g2_a21oi_2 _2040_ (.B1(_0527_),
    .Y(_0531_),
    .A2(_0530_),
    .A1(_0528_));
 sg13g2_nand2_1 _2041_ (.Y(_0532_),
    .A(net784),
    .B(net718));
 sg13g2_xnor2_1 _2042_ (.Y(_0533_),
    .A(net693),
    .B(net718));
 sg13g2_xor2_1 _2043_ (.B(_0533_),
    .A(_0531_),
    .X(_0080_));
 sg13g2_nand2_1 _2044_ (.Y(_0534_),
    .A(net729),
    .B(net756));
 sg13g2_xor2_1 _2045_ (.B(net756),
    .A(\cic_b.integrator[0][4] ),
    .X(_0535_));
 sg13g2_o21ai_1 _2046_ (.B1(_0532_),
    .Y(_0536_),
    .A1(_0531_),
    .A2(_0533_));
 sg13g2_nand2_1 _2047_ (.Y(_0537_),
    .A(_0535_),
    .B(_0536_));
 sg13g2_xor2_1 _2048_ (.B(_0536_),
    .A(_0535_),
    .X(_0081_));
 sg13g2_or2_1 _2049_ (.X(_0538_),
    .B(net771),
    .A(\cic_b.integrator[0][5] ));
 sg13g2_nand2_1 _2050_ (.Y(_0539_),
    .A(net625),
    .B(net771));
 sg13g2_nand2_1 _2051_ (.Y(_0540_),
    .A(_0538_),
    .B(_0539_));
 sg13g2_nand2_1 _2052_ (.Y(_0541_),
    .A(_0534_),
    .B(_0537_));
 sg13g2_xnor2_1 _2053_ (.Y(_0082_),
    .A(net772),
    .B(_0541_));
 sg13g2_nand2_1 _2054_ (.Y(_0542_),
    .A(net690),
    .B(net742));
 sg13g2_nor2_1 _2055_ (.A(net779),
    .B(net777),
    .Y(_0543_));
 sg13g2_xor2_1 _2056_ (.B(net742),
    .A(net690),
    .X(_0544_));
 sg13g2_nand2_1 _2057_ (.Y(_0545_),
    .A(_0534_),
    .B(_0539_));
 sg13g2_nand2b_1 _2058_ (.Y(_0546_),
    .B(_0537_),
    .A_N(_0545_));
 sg13g2_nand4_1 _2059_ (.B(_0536_),
    .C(_0538_),
    .A(_0535_),
    .Y(_0547_),
    .D(_0539_));
 sg13g2_nand2_1 _2060_ (.Y(_0548_),
    .A(_0538_),
    .B(_0546_));
 sg13g2_xnor2_1 _2061_ (.Y(_0083_),
    .A(_0544_),
    .B(_0548_));
 sg13g2_nor2_1 _2062_ (.A(\cic_b.integrator[0][7] ),
    .B(\cic_b.integrator[1][7] ),
    .Y(_0549_));
 sg13g2_nand2_1 _2063_ (.Y(_0550_),
    .A(\cic_b.integrator[0][7] ),
    .B(net752));
 sg13g2_nand2b_1 _2064_ (.Y(_0551_),
    .B(_0550_),
    .A_N(net753));
 sg13g2_o21ai_1 _2065_ (.B1(_0542_),
    .Y(_0552_),
    .A1(_0543_),
    .A2(_0548_));
 sg13g2_xnor2_1 _2066_ (.Y(_0084_),
    .A(_0551_),
    .B(_0552_));
 sg13g2_nand2_1 _2067_ (.Y(_0553_),
    .A(net727),
    .B(\cic_b.integrator[1][8] ));
 sg13g2_xnor2_1 _2068_ (.Y(_0554_),
    .A(net727),
    .B(net744));
 sg13g2_o21ai_1 _2069_ (.B1(_0550_),
    .Y(_0555_),
    .A1(_0542_),
    .A2(_0549_));
 sg13g2_a21oi_1 _2070_ (.A1(_0538_),
    .A2(_0545_),
    .Y(_0556_),
    .B1(_0555_));
 sg13g2_a221oi_1 _2071_ (.B2(_0547_),
    .C1(_0549_),
    .B1(_0556_),
    .A1(_0543_),
    .Y(_0557_),
    .A2(_0550_));
 sg13g2_nand2b_1 _2072_ (.Y(_0558_),
    .B(_0557_),
    .A_N(_0554_));
 sg13g2_xnor2_1 _2073_ (.Y(_0085_),
    .A(_0554_),
    .B(_0557_));
 sg13g2_nand2_1 _2074_ (.Y(_0559_),
    .A(_0553_),
    .B(_0558_));
 sg13g2_xnor2_1 _2075_ (.Y(_0560_),
    .A(net634),
    .B(net738));
 sg13g2_xnor2_1 _2076_ (.Y(_0086_),
    .A(_0559_),
    .B(_0560_));
 sg13g2_nor2_1 _2077_ (.A(_0554_),
    .B(_0560_),
    .Y(_0561_));
 sg13g2_a21oi_1 _2078_ (.A1(_1212_),
    .A2(_1232_),
    .Y(_0562_),
    .B1(_0553_));
 sg13g2_a221oi_1 _2079_ (.B2(_0561_),
    .C1(_0562_),
    .B1(_0557_),
    .A1(net762),
    .Y(_0563_),
    .A2(\cic_b.integrator[1][9] ));
 sg13g2_nand2_1 _2080_ (.Y(_0564_),
    .A(net733),
    .B(\cic_b.integrator[1][10] ));
 sg13g2_xnor2_1 _2081_ (.Y(_0565_),
    .A(net668),
    .B(net709));
 sg13g2_xor2_1 _2082_ (.B(_0565_),
    .A(_0563_),
    .X(_0075_));
 sg13g2_o21ai_1 _2083_ (.B1(net734),
    .Y(_0566_),
    .A1(_0563_),
    .A2(_0565_));
 sg13g2_nor2_1 _2084_ (.A(\cic_b.integrator[0][11] ),
    .B(\cic_b.integrator[1][11] ),
    .Y(_0567_));
 sg13g2_xnor2_1 _2085_ (.Y(_0568_),
    .A(net723),
    .B(net696));
 sg13g2_xnor2_1 _2086_ (.Y(_0076_),
    .A(_0566_),
    .B(_0568_));
 sg13g2_or2_1 _2087_ (.X(_0569_),
    .B(_0568_),
    .A(_0565_));
 sg13g2_nor2_1 _2088_ (.A(_0564_),
    .B(_0567_),
    .Y(_0570_));
 sg13g2_a21oi_1 _2089_ (.A1(\cic_b.integrator[0][11] ),
    .A2(\cic_b.integrator[1][11] ),
    .Y(_0571_),
    .B1(_0570_));
 sg13g2_o21ai_1 _2090_ (.B1(_0571_),
    .Y(_0572_),
    .A1(_0563_),
    .A2(_0569_));
 sg13g2_xnor2_1 _2091_ (.Y(_0573_),
    .A(net184),
    .B(net646));
 sg13g2_xnor2_1 _2092_ (.Y(_0077_),
    .A(_0572_),
    .B(_0573_));
 sg13g2_xor2_1 _2093_ (.B(net452),
    .A(net455),
    .X(_0074_));
 sg13g2_nand3_1 _2094_ (.B(net705),
    .C(net714),
    .A(net39),
    .Y(_0574_));
 sg13g2_a21o_1 _2095_ (.A2(net630),
    .A1(net39),
    .B1(net705),
    .X(_0575_));
 sg13g2_and2_1 _2096_ (.A(_0574_),
    .B(_0575_),
    .X(_0026_));
 sg13g2_nor2_2 _2097_ (.A(_1220_),
    .B(_0574_),
    .Y(_0576_));
 sg13g2_xnor2_1 _2098_ (.Y(_0027_),
    .A(net429),
    .B(_0574_));
 sg13g2_xor2_1 _2099_ (.B(_0576_),
    .A(net683),
    .X(_0028_));
 sg13g2_nand3_1 _2100_ (.B(net720),
    .C(_0576_),
    .A(net683),
    .Y(_0577_));
 sg13g2_a21o_1 _2101_ (.A2(_0576_),
    .A1(net683),
    .B1(net720),
    .X(_0578_));
 sg13g2_and2_1 _2102_ (.A(_0577_),
    .B(_0578_),
    .X(_0029_));
 sg13g2_nand4_1 _2103_ (.B(\cic_a.integrator[0][4] ),
    .C(net671),
    .A(\cic_a.integrator[0][3] ),
    .Y(_0579_),
    .D(_0576_));
 sg13g2_xnor2_1 _2104_ (.Y(_0030_),
    .A(net671),
    .B(_0577_));
 sg13g2_nor2_1 _2105_ (.A(_1221_),
    .B(_0579_),
    .Y(_0580_));
 sg13g2_xnor2_1 _2106_ (.Y(_0031_),
    .A(net677),
    .B(_0579_));
 sg13g2_xor2_1 _2107_ (.B(_0580_),
    .A(net688),
    .X(_0032_));
 sg13g2_nand3_1 _2108_ (.B(net715),
    .C(_0580_),
    .A(net790),
    .Y(_0581_));
 sg13g2_a21o_1 _2109_ (.A2(_0580_),
    .A1(net688),
    .B1(net715),
    .X(_0582_));
 sg13g2_and2_1 _2110_ (.A(_0581_),
    .B(_0582_),
    .X(_0033_));
 sg13g2_nor2_2 _2111_ (.A(_1222_),
    .B(_0581_),
    .Y(_0583_));
 sg13g2_xnor2_1 _2112_ (.Y(_0034_),
    .A(net627),
    .B(_0581_));
 sg13g2_xor2_1 _2113_ (.B(_0583_),
    .A(net673),
    .X(_0023_));
 sg13g2_nand3_1 _2114_ (.B(net722),
    .C(_0583_),
    .A(net673),
    .Y(_0584_));
 sg13g2_a21o_1 _2115_ (.A2(_0583_),
    .A1(net673),
    .B1(net722),
    .X(_0585_));
 sg13g2_and2_1 _2116_ (.A(_0584_),
    .B(_0585_),
    .X(_0024_));
 sg13g2_xnor2_1 _2117_ (.Y(_0025_),
    .A(net100),
    .B(_0584_));
 sg13g2_xor2_1 _2118_ (.B(\cic_a.integrator[0][0] ),
    .A(net39),
    .X(_0022_));
 sg13g2_nor2_2 _2119_ (.A(net3),
    .B(net546),
    .Y(_0586_));
 sg13g2_inv_1 _2120_ (.Y(_0587_),
    .A(_0586_));
 sg13g2_o21ai_1 _2121_ (.B1(net546),
    .Y(_0588_),
    .A1(\serializer_a.bit_cnt[0] ),
    .A2(net151));
 sg13g2_nand4_1 _2122_ (.B(net52),
    .C(net48),
    .A(net546),
    .Y(_0589_),
    .D(_0588_));
 sg13g2_and2_1 _2123_ (.A(net531),
    .B(_0589_),
    .X(_0016_));
 sg13g2_nor2_2 _2124_ (.A(net3),
    .B(net543),
    .Y(_0590_));
 sg13g2_inv_1 _2125_ (.Y(_0591_),
    .A(_0590_));
 sg13g2_o21ai_1 _2126_ (.B1(net543),
    .Y(_0592_),
    .A1(net108),
    .A2(net232));
 sg13g2_nand4_1 _2127_ (.B(net76),
    .C(net63),
    .A(net543),
    .Y(_0593_),
    .D(_0592_));
 sg13g2_and2_1 _2128_ (.A(_0591_),
    .B(_0593_),
    .X(_0020_));
 sg13g2_nor2_1 _2129_ (.A(net3),
    .B(net540),
    .Y(_0594_));
 sg13g2_or2_2 _2130_ (.X(_0595_),
    .B(net542),
    .A(net3));
 sg13g2_o21ai_1 _2131_ (.B1(net542),
    .Y(_0596_),
    .A1(net91),
    .A2(net106));
 sg13g2_nand4_1 _2132_ (.B(net96),
    .C(net81),
    .A(net540),
    .Y(_0597_),
    .D(_0596_));
 sg13g2_and2_1 _2133_ (.A(_0595_),
    .B(_0597_),
    .X(_0018_));
 sg13g2_mux2_1 _2134_ (.A0(net293),
    .A1(net159),
    .S(net523),
    .X(_0104_));
 sg13g2_mux2_1 _2135_ (.A0(net315),
    .A1(net153),
    .S(net523),
    .X(_0105_));
 sg13g2_mux2_1 _2136_ (.A0(net181),
    .A1(net121),
    .S(net520),
    .X(_0106_));
 sg13g2_mux2_1 _2137_ (.A0(net376),
    .A1(net212),
    .S(net522),
    .X(_0107_));
 sg13g2_mux2_1 _2138_ (.A0(net387),
    .A1(net163),
    .S(net515),
    .X(_0108_));
 sg13g2_mux2_1 _2139_ (.A0(\cic_a.delay[2][5] ),
    .A1(net397),
    .S(net514),
    .X(_0109_));
 sg13g2_mux2_1 _2140_ (.A0(net137),
    .A1(net395),
    .S(net514),
    .X(_0110_));
 sg13g2_mux2_1 _2141_ (.A0(net254),
    .A1(\cic_a.temp_delay[2][7] ),
    .S(net514),
    .X(_0111_));
 sg13g2_mux2_1 _2142_ (.A0(\cic_a.delay[2][8] ),
    .A1(net71),
    .S(net512),
    .X(_0112_));
 sg13g2_mux2_1 _2143_ (.A0(net421),
    .A1(net289),
    .S(net512),
    .X(_0113_));
 sg13g2_mux2_1 _2144_ (.A0(\cic_a.delay[2][10] ),
    .A1(net246),
    .S(net513),
    .X(_0114_));
 sg13g2_mux2_1 _2145_ (.A0(net424),
    .A1(net287),
    .S(net512),
    .X(_0115_));
 sg13g2_mux2_1 _2146_ (.A0(net415),
    .A1(net221),
    .S(net504),
    .X(_0116_));
 sg13g2_nor2_1 _2147_ (.A(net667),
    .B(net523),
    .Y(_0598_));
 sg13g2_nor2b_1 _2148_ (.A(net623),
    .B_N(net196),
    .Y(_0599_));
 sg13g2_xnor2_1 _2149_ (.Y(_0600_),
    .A(net623),
    .B(net196));
 sg13g2_a21oi_1 _2150_ (.A1(net523),
    .A2(_0600_),
    .Y(_0117_),
    .B1(_0598_));
 sg13g2_nor2_1 _2151_ (.A(net700),
    .B(net521),
    .Y(_0601_));
 sg13g2_nand2b_1 _2152_ (.Y(_0602_),
    .B(\cic_a.temp_comb[0][1] ),
    .A_N(\cic_a.delay[1][1] ));
 sg13g2_xor2_1 _2153_ (.B(net325),
    .A(net663),
    .X(_0603_));
 sg13g2_xnor2_1 _2154_ (.Y(_0604_),
    .A(_0599_),
    .B(_0603_));
 sg13g2_a21oi_1 _2155_ (.A1(net521),
    .A2(_0604_),
    .Y(_0118_),
    .B1(_0601_));
 sg13g2_nor2_1 _2156_ (.A(net675),
    .B(net521),
    .Y(_0605_));
 sg13g2_nor2b_1 _2157_ (.A(net373),
    .B_N(\cic_a.temp_comb[0][2] ),
    .Y(_0606_));
 sg13g2_xnor2_1 _2158_ (.Y(_0607_),
    .A(\cic_a.temp_comb[0][2] ),
    .B(\cic_a.delay[1][2] ));
 sg13g2_o21ai_1 _2159_ (.B1(_0602_),
    .Y(_0608_),
    .A1(_0599_),
    .A2(_0603_));
 sg13g2_xnor2_1 _2160_ (.Y(_0609_),
    .A(_0607_),
    .B(_0608_));
 sg13g2_a21oi_1 _2161_ (.A1(net522),
    .A2(_0609_),
    .Y(_0119_),
    .B1(_0605_));
 sg13g2_nor2_1 _2162_ (.A(net685),
    .B(net515),
    .Y(_0610_));
 sg13g2_nand2b_1 _2163_ (.Y(_0611_),
    .B(\cic_a.temp_comb[0][3] ),
    .A_N(\cic_a.delay[1][3] ));
 sg13g2_xor2_1 _2164_ (.B(net243),
    .A(\cic_a.temp_comb[0][3] ),
    .X(_0612_));
 sg13g2_a21oi_2 _2165_ (.B1(_0606_),
    .Y(_0613_),
    .A2(_0608_),
    .A1(_0607_));
 sg13g2_xnor2_1 _2166_ (.Y(_0614_),
    .A(_0612_),
    .B(_0613_));
 sg13g2_a21oi_1 _2167_ (.A1(net515),
    .A2(_0614_),
    .Y(_0120_),
    .B1(_0610_));
 sg13g2_nor2_1 _2168_ (.A(net695),
    .B(net514),
    .Y(_0615_));
 sg13g2_o21ai_1 _2169_ (.B1(_0611_),
    .Y(_0616_),
    .A1(_0612_),
    .A2(_0613_));
 sg13g2_nor2_1 _2170_ (.A(_1216_),
    .B(net428),
    .Y(_0617_));
 sg13g2_xnor2_1 _2171_ (.Y(_0618_),
    .A(\cic_a.temp_comb[0][4] ),
    .B(\cic_a.delay[1][4] ));
 sg13g2_inv_1 _2172_ (.Y(_0619_),
    .A(_0618_));
 sg13g2_xnor2_1 _2173_ (.Y(_0620_),
    .A(_0616_),
    .B(_0618_));
 sg13g2_a21oi_1 _2174_ (.A1(net514),
    .A2(_0620_),
    .Y(_0121_),
    .B1(_0615_));
 sg13g2_nor2_1 _2175_ (.A(net409),
    .B(net511),
    .Y(_0621_));
 sg13g2_nand2b_1 _2176_ (.Y(_0622_),
    .B(\cic_a.delay[1][5] ),
    .A_N(\cic_a.temp_comb[0][5] ));
 sg13g2_nor2b_1 _2177_ (.A(\cic_a.delay[1][5] ),
    .B_N(\cic_a.temp_comb[0][5] ),
    .Y(_0623_));
 sg13g2_xor2_1 _2178_ (.B(net382),
    .A(\cic_a.temp_comb[0][5] ),
    .X(_0624_));
 sg13g2_a21oi_1 _2179_ (.A1(_0616_),
    .A2(_0618_),
    .Y(_0625_),
    .B1(_0617_));
 sg13g2_xnor2_1 _2180_ (.Y(_0626_),
    .A(net666),
    .B(_0625_));
 sg13g2_a21oi_1 _2181_ (.A1(net511),
    .A2(_0626_),
    .Y(_0122_),
    .B1(_0621_));
 sg13g2_nor2_1 _2182_ (.A(net694),
    .B(net509),
    .Y(_0627_));
 sg13g2_nand2b_1 _2183_ (.Y(_0628_),
    .B(\cic_a.temp_comb[0][6] ),
    .A_N(\cic_a.delay[1][6] ));
 sg13g2_xor2_1 _2184_ (.B(\cic_a.delay[1][6] ),
    .A(\cic_a.temp_comb[0][6] ),
    .X(_0629_));
 sg13g2_nor2_1 _2185_ (.A(_0619_),
    .B(_0624_),
    .Y(_0630_));
 sg13g2_a21o_1 _2186_ (.A2(_0622_),
    .A1(_0617_),
    .B1(_0623_),
    .X(_0631_));
 sg13g2_a21oi_1 _2187_ (.A1(_0616_),
    .A2(_0630_),
    .Y(_0632_),
    .B1(_0631_));
 sg13g2_xnor2_1 _2188_ (.Y(_0633_),
    .A(_0629_),
    .B(_0632_));
 sg13g2_a21oi_1 _2189_ (.A1(net509),
    .A2(_0633_),
    .Y(_0123_),
    .B1(_0627_));
 sg13g2_nor2_1 _2190_ (.A(net680),
    .B(net509),
    .Y(_0634_));
 sg13g2_nor2b_1 _2191_ (.A(\cic_a.temp_comb[0][7] ),
    .B_N(\cic_a.delay[1][7] ),
    .Y(_0635_));
 sg13g2_nand2b_1 _2192_ (.Y(_0636_),
    .B(\cic_a.temp_comb[0][7] ),
    .A_N(\cic_a.delay[1][7] ));
 sg13g2_nand2b_1 _2193_ (.Y(_0637_),
    .B(_0636_),
    .A_N(_0635_));
 sg13g2_o21ai_1 _2194_ (.B1(_0628_),
    .Y(_0638_),
    .A1(_0629_),
    .A2(_0632_));
 sg13g2_xor2_1 _2195_ (.B(_0638_),
    .A(_0637_),
    .X(_0639_));
 sg13g2_a21oi_1 _2196_ (.A1(net511),
    .A2(_0639_),
    .Y(_0124_),
    .B1(_0634_));
 sg13g2_nor2_1 _2197_ (.A(_0629_),
    .B(_0637_),
    .Y(_0640_));
 sg13g2_and2_1 _2198_ (.A(_0630_),
    .B(_0640_),
    .X(_0641_));
 sg13g2_o21ai_1 _2199_ (.B1(_0636_),
    .Y(_0642_),
    .A1(_0628_),
    .A2(_0635_));
 sg13g2_a221oi_1 _2200_ (.B2(_0616_),
    .C1(_0642_),
    .B1(_0641_),
    .A1(_0631_),
    .Y(_0643_),
    .A2(_0640_));
 sg13g2_nand2b_1 _2201_ (.Y(_0644_),
    .B(\cic_a.temp_comb[0][8] ),
    .A_N(\cic_a.delay[1][8] ));
 sg13g2_xor2_1 _2202_ (.B(\cic_a.delay[1][8] ),
    .A(\cic_a.temp_comb[0][8] ),
    .X(_0645_));
 sg13g2_xnor2_1 _2203_ (.Y(_0646_),
    .A(_0643_),
    .B(_0645_));
 sg13g2_nor2_1 _2204_ (.A(net338),
    .B(net507),
    .Y(_0647_));
 sg13g2_a21oi_1 _2205_ (.A1(net507),
    .A2(_0646_),
    .Y(_0125_),
    .B1(_0647_));
 sg13g2_xnor2_1 _2206_ (.Y(_0648_),
    .A(\cic_a.temp_comb[0][9] ),
    .B(\cic_a.delay[1][9] ));
 sg13g2_o21ai_1 _2207_ (.B1(_0644_),
    .Y(_0649_),
    .A1(_0643_),
    .A2(_0645_));
 sg13g2_xnor2_1 _2208_ (.Y(_0650_),
    .A(_0648_),
    .B(_0649_));
 sg13g2_nor2_1 _2209_ (.A(net631),
    .B(net507),
    .Y(_0651_));
 sg13g2_a21oi_1 _2210_ (.A1(net507),
    .A2(_0650_),
    .Y(_0126_),
    .B1(_0651_));
 sg13g2_nor2_1 _2211_ (.A(net284),
    .B(net505),
    .Y(_0652_));
 sg13g2_nand2b_1 _2212_ (.Y(_0653_),
    .B(_0648_),
    .A_N(_0645_));
 sg13g2_a21oi_1 _2213_ (.A1(_1217_),
    .A2(\cic_a.delay[1][9] ),
    .Y(_0654_),
    .B1(_0644_));
 sg13g2_a21oi_1 _2214_ (.A1(\cic_a.temp_comb[0][9] ),
    .A2(_1218_),
    .Y(_0655_),
    .B1(_0654_));
 sg13g2_o21ai_1 _2215_ (.B1(_0655_),
    .Y(_0656_),
    .A1(_0643_),
    .A2(_0653_));
 sg13g2_nor2b_1 _2216_ (.A(\cic_a.delay[1][10] ),
    .B_N(\cic_a.temp_comb[0][10] ),
    .Y(_0657_));
 sg13g2_nor2b_1 _2217_ (.A(\cic_a.temp_comb[0][10] ),
    .B_N(\cic_a.delay[1][10] ),
    .Y(_0658_));
 sg13g2_nor2_1 _2218_ (.A(_0657_),
    .B(_0658_),
    .Y(_0659_));
 sg13g2_xnor2_1 _2219_ (.Y(_0660_),
    .A(_0656_),
    .B(_0659_));
 sg13g2_a21oi_1 _2220_ (.A1(net505),
    .A2(_0660_),
    .Y(_0127_),
    .B1(_0652_));
 sg13g2_nor2_1 _2221_ (.A(net692),
    .B(net505),
    .Y(_0661_));
 sg13g2_nor2b_1 _2222_ (.A(\cic_a.delay[1][11] ),
    .B_N(\cic_a.temp_comb[0][11] ),
    .Y(_0662_));
 sg13g2_nand2b_1 _2223_ (.Y(_0663_),
    .B(\cic_a.delay[1][11] ),
    .A_N(\cic_a.temp_comb[0][11] ));
 sg13g2_nand2b_1 _2224_ (.Y(_0664_),
    .B(_0663_),
    .A_N(_0662_));
 sg13g2_a21oi_1 _2225_ (.A1(_0656_),
    .A2(_0659_),
    .Y(_0665_),
    .B1(_0657_));
 sg13g2_xnor2_1 _2226_ (.Y(_0666_),
    .A(_0664_),
    .B(_0665_));
 sg13g2_a21oi_1 _2227_ (.A1(net505),
    .A2(_0666_),
    .Y(_0128_),
    .B1(_0661_));
 sg13g2_nor2_1 _2228_ (.A(net467),
    .B(net504),
    .Y(_0667_));
 sg13g2_nor3_1 _2229_ (.A(_0657_),
    .B(_0658_),
    .C(_0664_),
    .Y(_0668_));
 sg13g2_a221oi_1 _2230_ (.B2(_0656_),
    .C1(_0662_),
    .B1(_0668_),
    .A1(_0657_),
    .Y(_0669_),
    .A2(_0663_));
 sg13g2_xor2_1 _2231_ (.B(\cic_a.delay[1][12] ),
    .A(\cic_a.temp_comb[0][12] ),
    .X(_0670_));
 sg13g2_xnor2_1 _2232_ (.Y(_0671_),
    .A(_0669_),
    .B(_0670_));
 sg13g2_a21oi_1 _2233_ (.A1(net504),
    .A2(_0671_),
    .Y(_0129_),
    .B1(_0667_));
 sg13g2_mux2_1 _2234_ (.A0(net196),
    .A1(net128),
    .S(net521),
    .X(_0130_));
 sg13g2_mux2_1 _2235_ (.A0(net325),
    .A1(net309),
    .S(net519),
    .X(_0131_));
 sg13g2_mux2_1 _2236_ (.A0(net373),
    .A1(net167),
    .S(net519),
    .X(_0132_));
 sg13g2_mux2_1 _2237_ (.A0(net243),
    .A1(net156),
    .S(net515),
    .X(_0133_));
 sg13g2_mux2_1 _2238_ (.A0(net428),
    .A1(net393),
    .S(net509),
    .X(_0134_));
 sg13g2_mux2_1 _2239_ (.A0(net382),
    .A1(net225),
    .S(net510),
    .X(_0135_));
 sg13g2_mux2_1 _2240_ (.A0(\cic_a.delay[1][6] ),
    .A1(net139),
    .S(net510),
    .X(_0136_));
 sg13g2_mux2_1 _2241_ (.A0(net389),
    .A1(net252),
    .S(net510),
    .X(_0137_));
 sg13g2_mux2_1 _2242_ (.A0(net432),
    .A1(net364),
    .S(net506),
    .X(_0138_));
 sg13g2_nand2_1 _2243_ (.Y(_0672_),
    .A(net50),
    .B(net506));
 sg13g2_o21ai_1 _2244_ (.B1(_0672_),
    .Y(_0139_),
    .A1(_1218_),
    .A2(net506));
 sg13g2_mux2_1 _2245_ (.A0(net329),
    .A1(net274),
    .S(net501),
    .X(_0140_));
 sg13g2_mux2_1 _2246_ (.A0(net295),
    .A1(net281),
    .S(net501),
    .X(_0141_));
 sg13g2_mux2_1 _2247_ (.A0(net294),
    .A1(net165),
    .S(net500),
    .X(_0142_));
 sg13g2_mux2_1 _2248_ (.A0(net390),
    .A1(net197),
    .S(net518),
    .X(_0143_));
 sg13g2_mux2_1 _2249_ (.A0(net388),
    .A1(net237),
    .S(net518),
    .X(_0144_));
 sg13g2_mux2_1 _2250_ (.A0(\cic_a.delay[0][2] ),
    .A1(net110),
    .S(net518),
    .X(_0145_));
 sg13g2_mux2_1 _2251_ (.A0(\cic_a.delay[0][3] ),
    .A1(net141),
    .S(net513),
    .X(_0146_));
 sg13g2_mux2_1 _2252_ (.A0(net414),
    .A1(net344),
    .S(net512),
    .X(_0147_));
 sg13g2_nand2_1 _2253_ (.Y(_0673_),
    .A(net22),
    .B(net508));
 sg13g2_o21ai_1 _2254_ (.B1(_0673_),
    .Y(_0148_),
    .A1(_1213_),
    .A2(net507));
 sg13g2_mux2_1 _2255_ (.A0(net370),
    .A1(net327),
    .S(net508),
    .X(_0149_));
 sg13g2_nand2_1 _2256_ (.Y(_0674_),
    .A(net41),
    .B(net508));
 sg13g2_o21ai_1 _2257_ (.B1(_0674_),
    .Y(_0150_),
    .A1(_1214_),
    .A2(net508));
 sg13g2_mux2_1 _2258_ (.A0(net217),
    .A1(net189),
    .S(net501),
    .X(_0151_));
 sg13g2_mux2_1 _2259_ (.A0(net406),
    .A1(net98),
    .S(net500),
    .X(_0152_));
 sg13g2_mux2_1 _2260_ (.A0(\cic_a.delay[0][10] ),
    .A1(net54),
    .S(net503),
    .X(_0153_));
 sg13g2_mux2_1 _2261_ (.A0(net314),
    .A1(net227),
    .S(net503),
    .X(_0154_));
 sg13g2_mux2_1 _2262_ (.A0(net362),
    .A1(net306),
    .S(net503),
    .X(_0155_));
 sg13g2_nor2_1 _2263_ (.A(net623),
    .B(net520),
    .Y(_0675_));
 sg13g2_nand2b_1 _2264_ (.Y(_0676_),
    .B(net390),
    .A_N(\cic_a.integrator[2][0] ));
 sg13g2_xnor2_1 _2265_ (.Y(_0677_),
    .A(\cic_a.integrator[2][0] ),
    .B(net390));
 sg13g2_a21oi_1 _2266_ (.A1(net520),
    .A2(_0677_),
    .Y(_0156_),
    .B1(_0675_));
 sg13g2_nor2_1 _2267_ (.A(net663),
    .B(net519),
    .Y(_0678_));
 sg13g2_nor2b_1 _2268_ (.A(net388),
    .B_N(\cic_a.integrator[2][1] ),
    .Y(_0679_));
 sg13g2_xnor2_1 _2269_ (.Y(_0680_),
    .A(\cic_a.integrator[2][1] ),
    .B(net388));
 sg13g2_xnor2_1 _2270_ (.Y(_0681_),
    .A(_0676_),
    .B(_0680_));
 sg13g2_a21oi_1 _2271_ (.A1(net519),
    .A2(_0681_),
    .Y(_0157_),
    .B1(_0678_));
 sg13g2_nor2_1 _2272_ (.A(net657),
    .B(net519),
    .Y(_0682_));
 sg13g2_nand2b_1 _2273_ (.Y(_0683_),
    .B(\cic_a.integrator[2][2] ),
    .A_N(\cic_a.delay[0][2] ));
 sg13g2_xor2_1 _2274_ (.B(\cic_a.delay[0][2] ),
    .A(\cic_a.integrator[2][2] ),
    .X(_0684_));
 sg13g2_a21oi_1 _2275_ (.A1(_0676_),
    .A2(_0680_),
    .Y(_0685_),
    .B1(_0679_));
 sg13g2_xnor2_1 _2276_ (.Y(_0686_),
    .A(_0684_),
    .B(_0685_));
 sg13g2_a21oi_1 _2277_ (.A1(net519),
    .A2(_0686_),
    .Y(_0158_),
    .B1(_0682_));
 sg13g2_nor2_1 _2278_ (.A(net648),
    .B(net515),
    .Y(_0687_));
 sg13g2_nor2b_1 _2279_ (.A(\cic_a.delay[0][3] ),
    .B_N(\cic_a.integrator[2][3] ),
    .Y(_0688_));
 sg13g2_nand2b_1 _2280_ (.Y(_0689_),
    .B(\cic_a.delay[0][3] ),
    .A_N(\cic_a.integrator[2][3] ));
 sg13g2_nor2b_1 _2281_ (.A(_0688_),
    .B_N(_0689_),
    .Y(_0690_));
 sg13g2_o21ai_1 _2282_ (.B1(_0683_),
    .Y(_0691_),
    .A1(_0684_),
    .A2(_0685_));
 sg13g2_xnor2_1 _2283_ (.Y(_0692_),
    .A(_0690_),
    .B(_0691_));
 sg13g2_a21oi_1 _2284_ (.A1(net515),
    .A2(_0692_),
    .Y(_0159_),
    .B1(_0687_));
 sg13g2_a21o_2 _2285_ (.A2(_0691_),
    .A1(_0689_),
    .B1(_0688_),
    .X(_0693_));
 sg13g2_nor2b_1 _2286_ (.A(\cic_a.delay[0][4] ),
    .B_N(\cic_a.integrator[2][4] ),
    .Y(_0694_));
 sg13g2_xor2_1 _2287_ (.B(\cic_a.delay[0][4] ),
    .A(\cic_a.integrator[2][4] ),
    .X(_0695_));
 sg13g2_nand2b_1 _2288_ (.Y(_0696_),
    .B(_0695_),
    .A_N(_0693_));
 sg13g2_nand2b_1 _2289_ (.Y(_0697_),
    .B(_0693_),
    .A_N(_0695_));
 sg13g2_nand3_1 _2290_ (.B(_0696_),
    .C(_0697_),
    .A(net507),
    .Y(_0698_));
 sg13g2_o21ai_1 _2291_ (.B1(_0698_),
    .Y(_0160_),
    .A1(_1216_),
    .A2(net509));
 sg13g2_nor2_1 _2292_ (.A(\cic_a.integrator[2][5] ),
    .B(_1213_),
    .Y(_0699_));
 sg13g2_xor2_1 _2293_ (.B(net669),
    .A(\cic_a.integrator[2][5] ),
    .X(_0700_));
 sg13g2_nor2b_1 _2294_ (.A(_0694_),
    .B_N(_0697_),
    .Y(_0701_));
 sg13g2_xnor2_1 _2295_ (.Y(_0702_),
    .A(_0700_),
    .B(_0701_));
 sg13g2_nor2_1 _2296_ (.A(net665),
    .B(net509),
    .Y(_0703_));
 sg13g2_a21oi_1 _2297_ (.A1(net509),
    .A2(_0702_),
    .Y(_0161_),
    .B1(_0703_));
 sg13g2_nor2_1 _2298_ (.A(net171),
    .B(net510),
    .Y(_0704_));
 sg13g2_nor2b_1 _2299_ (.A(\cic_a.delay[0][6] ),
    .B_N(\cic_a.integrator[2][6] ),
    .Y(_0705_));
 sg13g2_nand2b_1 _2300_ (.Y(_0706_),
    .B(\cic_a.delay[0][6] ),
    .A_N(\cic_a.integrator[2][6] ));
 sg13g2_nand2b_1 _2301_ (.Y(_0707_),
    .B(_0706_),
    .A_N(_0705_));
 sg13g2_a21oi_1 _2302_ (.A1(\cic_a.integrator[2][5] ),
    .A2(_1213_),
    .Y(_0708_),
    .B1(_0694_));
 sg13g2_a21oi_1 _2303_ (.A1(_0697_),
    .A2(_0708_),
    .Y(_0709_),
    .B1(_0699_));
 sg13g2_xor2_1 _2304_ (.B(_0709_),
    .A(_0707_),
    .X(_0710_));
 sg13g2_a21oi_1 _2305_ (.A1(net507),
    .A2(_0710_),
    .Y(_0162_),
    .B1(_0704_));
 sg13g2_nor2_1 _2306_ (.A(net620),
    .B(net506),
    .Y(_0711_));
 sg13g2_nand2_1 _2307_ (.Y(_0712_),
    .A(\cic_a.integrator[2][7] ),
    .B(_1214_));
 sg13g2_xor2_1 _2308_ (.B(\cic_a.delay[0][7] ),
    .A(\cic_a.integrator[2][7] ),
    .X(_0713_));
 sg13g2_a21oi_1 _2309_ (.A1(_0706_),
    .A2(_0709_),
    .Y(_0714_),
    .B1(_0705_));
 sg13g2_xnor2_1 _2310_ (.Y(_0715_),
    .A(_0713_),
    .B(_0714_));
 sg13g2_a21oi_1 _2311_ (.A1(net506),
    .A2(_0715_),
    .Y(_0163_),
    .B1(_0711_));
 sg13g2_nor2_1 _2312_ (.A(net659),
    .B(net505),
    .Y(_0716_));
 sg13g2_nor4_1 _2313_ (.A(_0695_),
    .B(_0700_),
    .C(_0707_),
    .D(_0713_),
    .Y(_0717_));
 sg13g2_o21ai_1 _2314_ (.B1(_0705_),
    .Y(_0718_),
    .A1(\cic_a.integrator[2][7] ),
    .A2(_1214_));
 sg13g2_or4_1 _2315_ (.A(_0699_),
    .B(_0707_),
    .C(_0708_),
    .D(_0713_),
    .X(_0719_));
 sg13g2_nand3_1 _2316_ (.B(_0718_),
    .C(_0719_),
    .A(_0712_),
    .Y(_0720_));
 sg13g2_a21oi_2 _2317_ (.B1(_0720_),
    .Y(_0721_),
    .A2(_0717_),
    .A1(_0693_));
 sg13g2_nor2b_1 _2318_ (.A(\cic_a.delay[0][8] ),
    .B_N(\cic_a.integrator[2][8] ),
    .Y(_0722_));
 sg13g2_xnor2_1 _2319_ (.Y(_0723_),
    .A(\cic_a.integrator[2][8] ),
    .B(\cic_a.delay[0][8] ));
 sg13g2_nor2b_1 _2320_ (.A(_0721_),
    .B_N(_0723_),
    .Y(_0724_));
 sg13g2_xor2_1 _2321_ (.B(_0723_),
    .A(_0721_),
    .X(_0725_));
 sg13g2_a21oi_1 _2322_ (.A1(net505),
    .A2(_0725_),
    .Y(_0164_),
    .B1(_0716_));
 sg13g2_nor2_1 _2323_ (.A(_1215_),
    .B(\cic_a.delay[0][9] ),
    .Y(_0726_));
 sg13g2_nand2_1 _2324_ (.Y(_0727_),
    .A(_1215_),
    .B(\cic_a.delay[0][9] ));
 sg13g2_nand2b_1 _2325_ (.Y(_0728_),
    .B(_0727_),
    .A_N(_0726_));
 sg13g2_nor2_1 _2326_ (.A(_0722_),
    .B(_0724_),
    .Y(_0729_));
 sg13g2_xnor2_1 _2327_ (.Y(_0730_),
    .A(_0728_),
    .B(_0729_));
 sg13g2_nor2_1 _2328_ (.A(net145),
    .B(net505),
    .Y(_0731_));
 sg13g2_a21oi_1 _2329_ (.A1(net505),
    .A2(_0730_),
    .Y(_0165_),
    .B1(_0731_));
 sg13g2_nor2_1 _2330_ (.A(net629),
    .B(net501),
    .Y(_0732_));
 sg13g2_nor2b_1 _2331_ (.A(\cic_a.delay[0][10] ),
    .B_N(\cic_a.integrator[2][10] ),
    .Y(_0733_));
 sg13g2_xnor2_1 _2332_ (.Y(_0734_),
    .A(\cic_a.integrator[2][10] ),
    .B(\cic_a.delay[0][10] ));
 sg13g2_inv_1 _2333_ (.Y(_0735_),
    .A(_0734_));
 sg13g2_nand3b_1 _2334_ (.B(_0727_),
    .C(_0723_),
    .Y(_0736_),
    .A_N(_0726_));
 sg13g2_a21oi_1 _2335_ (.A1(_0722_),
    .A2(_0727_),
    .Y(_0737_),
    .B1(_0726_));
 sg13g2_o21ai_1 _2336_ (.B1(_0737_),
    .Y(_0738_),
    .A1(_0721_),
    .A2(_0736_));
 sg13g2_xnor2_1 _2337_ (.Y(_0739_),
    .A(_0734_),
    .B(_0738_));
 sg13g2_a21oi_1 _2338_ (.A1(net501),
    .A2(_0739_),
    .Y(_0166_),
    .B1(_0732_));
 sg13g2_nor2b_1 _2339_ (.A(net314),
    .B_N(\cic_a.integrator[2][11] ),
    .Y(_0740_));
 sg13g2_nand2b_1 _2340_ (.Y(_0741_),
    .B(\cic_a.delay[0][11] ),
    .A_N(\cic_a.integrator[2][11] ));
 sg13g2_nand2b_1 _2341_ (.Y(_0742_),
    .B(_0741_),
    .A_N(_0740_));
 sg13g2_a21oi_1 _2342_ (.A1(_0734_),
    .A2(_0738_),
    .Y(_0743_),
    .B1(_0733_));
 sg13g2_xnor2_1 _2343_ (.Y(_0744_),
    .A(_0742_),
    .B(_0743_));
 sg13g2_nor2_1 _2344_ (.A(net441),
    .B(net501),
    .Y(_0745_));
 sg13g2_a21oi_1 _2345_ (.A1(net500),
    .A2(_0744_),
    .Y(_0167_),
    .B1(_0745_));
 sg13g2_nor2_1 _2346_ (.A(net660),
    .B(net500),
    .Y(_0746_));
 sg13g2_nor2_1 _2347_ (.A(_0735_),
    .B(_0742_),
    .Y(_0747_));
 sg13g2_a221oi_1 _2348_ (.B2(_0738_),
    .C1(_0740_),
    .B1(_0747_),
    .A1(_0733_),
    .Y(_0748_),
    .A2(_0741_));
 sg13g2_xor2_1 _2349_ (.B(net362),
    .A(\cic_a.integrator[2][12] ),
    .X(_0749_));
 sg13g2_xnor2_1 _2350_ (.Y(_0750_),
    .A(_0748_),
    .B(_0749_));
 sg13g2_a21oi_1 _2351_ (.A1(net500),
    .A2(_0750_),
    .Y(_0168_),
    .B1(_0746_));
 sg13g2_mux2_1 _2352_ (.A0(net451),
    .A1(net119),
    .S(net525),
    .X(_0169_));
 sg13g2_mux2_1 _2353_ (.A0(net360),
    .A1(net114),
    .S(net525),
    .X(_0170_));
 sg13g2_mux2_1 _2354_ (.A0(net465),
    .A1(net391),
    .S(net525),
    .X(_0171_));
 sg13g2_mux2_1 _2355_ (.A0(net454),
    .A1(net132),
    .S(net524),
    .X(_0172_));
 sg13g2_mux2_1 _2356_ (.A0(net450),
    .A1(net313),
    .S(net524),
    .X(_0173_));
 sg13g2_mux2_1 _2357_ (.A0(net326),
    .A1(net231),
    .S(net524),
    .X(_0174_));
 sg13g2_mux2_1 _2358_ (.A0(net436),
    .A1(net271),
    .S(net520),
    .X(_0175_));
 sg13g2_nand2_1 _2359_ (.Y(_0751_),
    .A(net94),
    .B(net524));
 sg13g2_o21ai_1 _2360_ (.B1(_0751_),
    .Y(_0176_),
    .A1(_1196_),
    .A2(net526));
 sg13g2_mux2_1 _2361_ (.A0(net435),
    .A1(net270),
    .S(net517),
    .X(_0177_));
 sg13g2_mux2_1 _2362_ (.A0(net296),
    .A1(net265),
    .S(net526),
    .X(_0178_));
 sg13g2_mux2_1 _2363_ (.A0(net460),
    .A1(net439),
    .S(net517),
    .X(_0179_));
 sg13g2_mux2_1 _2364_ (.A0(net380),
    .A1(net191),
    .S(net517),
    .X(_0180_));
 sg13g2_mux2_1 _2365_ (.A0(net431),
    .A1(net412),
    .S(net528),
    .X(_0181_));
 sg13g2_nor2_1 _2366_ (.A(net119),
    .B(net525),
    .Y(_0752_));
 sg13g2_nor2b_1 _2367_ (.A(\cic_a.temp_comb[1][0] ),
    .B_N(\cic_a.delay[2][0] ),
    .Y(_0753_));
 sg13g2_xnor2_1 _2368_ (.Y(_0754_),
    .A(\cic_a.temp_comb[1][0] ),
    .B(\cic_a.delay[2][0] ));
 sg13g2_a21oi_1 _2369_ (.A1(net526),
    .A2(_0754_),
    .Y(_0182_),
    .B1(_0752_));
 sg13g2_nor2_1 _2370_ (.A(net114),
    .B(net526),
    .Y(_0755_));
 sg13g2_nand2b_1 _2371_ (.Y(_0756_),
    .B(\cic_a.temp_comb[1][1] ),
    .A_N(\cic_a.delay[2][1] ));
 sg13g2_xor2_1 _2372_ (.B(\cic_a.delay[2][1] ),
    .A(\cic_a.temp_comb[1][1] ),
    .X(_0757_));
 sg13g2_xnor2_1 _2373_ (.Y(_0758_),
    .A(_0753_),
    .B(_0757_));
 sg13g2_a21oi_1 _2374_ (.A1(net525),
    .A2(_0758_),
    .Y(_0183_),
    .B1(_0755_));
 sg13g2_nor2_1 _2375_ (.A(net391),
    .B(net525),
    .Y(_0759_));
 sg13g2_nor2b_1 _2376_ (.A(\cic_a.delay[2][2] ),
    .B_N(\cic_a.temp_comb[1][2] ),
    .Y(_0760_));
 sg13g2_xnor2_1 _2377_ (.Y(_0761_),
    .A(\cic_a.temp_comb[1][2] ),
    .B(\cic_a.delay[2][2] ));
 sg13g2_o21ai_1 _2378_ (.B1(_0756_),
    .Y(_0762_),
    .A1(_0753_),
    .A2(_0757_));
 sg13g2_xnor2_1 _2379_ (.Y(_0763_),
    .A(_0761_),
    .B(_0762_));
 sg13g2_a21oi_1 _2380_ (.A1(net523),
    .A2(_0763_),
    .Y(_0184_),
    .B1(_0759_));
 sg13g2_nor2_1 _2381_ (.A(net132),
    .B(net523),
    .Y(_0764_));
 sg13g2_nand2b_1 _2382_ (.Y(_0765_),
    .B(\cic_a.temp_comb[1][3] ),
    .A_N(\cic_a.delay[2][3] ));
 sg13g2_xor2_1 _2383_ (.B(\cic_a.delay[2][3] ),
    .A(\cic_a.temp_comb[1][3] ),
    .X(_0766_));
 sg13g2_a21oi_2 _2384_ (.B1(_0760_),
    .Y(_0767_),
    .A2(_0762_),
    .A1(_0761_));
 sg13g2_xnor2_1 _2385_ (.Y(_0768_),
    .A(_0766_),
    .B(_0767_));
 sg13g2_a21oi_1 _2386_ (.A1(net523),
    .A2(_0768_),
    .Y(_0185_),
    .B1(_0764_));
 sg13g2_o21ai_1 _2387_ (.B1(_0765_),
    .Y(_0769_),
    .A1(_0766_),
    .A2(_0767_));
 sg13g2_nand2b_1 _2388_ (.Y(_0770_),
    .B(\cic_a.temp_comb[1][4] ),
    .A_N(\cic_a.delay[2][4] ));
 sg13g2_xor2_1 _2389_ (.B(\cic_a.delay[2][4] ),
    .A(\cic_a.temp_comb[1][4] ),
    .X(_0771_));
 sg13g2_nand2b_1 _2390_ (.Y(_0772_),
    .B(_0769_),
    .A_N(_0771_));
 sg13g2_xor2_1 _2391_ (.B(_0771_),
    .A(_0769_),
    .X(_0773_));
 sg13g2_nor2_1 _2392_ (.A(net313),
    .B(net524),
    .Y(_0774_));
 sg13g2_a21oi_1 _2393_ (.A1(net524),
    .A2(_0773_),
    .Y(_0186_),
    .B1(_0774_));
 sg13g2_nor2b_1 _2394_ (.A(\cic_a.temp_comb[1][5] ),
    .B_N(\cic_a.delay[2][5] ),
    .Y(_0775_));
 sg13g2_nand2b_1 _2395_ (.Y(_0776_),
    .B(\cic_a.temp_comb[1][5] ),
    .A_N(\cic_a.delay[2][5] ));
 sg13g2_nand2b_1 _2396_ (.Y(_0777_),
    .B(_0776_),
    .A_N(_0775_));
 sg13g2_and2_1 _2397_ (.A(_0770_),
    .B(_0772_),
    .X(_0778_));
 sg13g2_xor2_1 _2398_ (.B(_0778_),
    .A(_0777_),
    .X(_0779_));
 sg13g2_mux2_1 _2399_ (.A0(net231),
    .A1(_0779_),
    .S(net524),
    .X(_0187_));
 sg13g2_nor2_1 _2400_ (.A(net271),
    .B(net520),
    .Y(_0780_));
 sg13g2_nand2b_1 _2401_ (.Y(_0781_),
    .B(\cic_a.temp_comb[1][6] ),
    .A_N(\cic_a.delay[2][6] ));
 sg13g2_xor2_1 _2402_ (.B(\cic_a.delay[2][6] ),
    .A(\cic_a.temp_comb[1][6] ),
    .X(_0782_));
 sg13g2_nor2_1 _2403_ (.A(_0771_),
    .B(_0777_),
    .Y(_0783_));
 sg13g2_o21ai_1 _2404_ (.B1(_0776_),
    .Y(_0784_),
    .A1(_0770_),
    .A2(_0775_));
 sg13g2_a21oi_1 _2405_ (.A1(_0769_),
    .A2(_0783_),
    .Y(_0785_),
    .B1(_0784_));
 sg13g2_xnor2_1 _2406_ (.Y(_0786_),
    .A(_0782_),
    .B(_0785_));
 sg13g2_a21oi_1 _2407_ (.A1(net520),
    .A2(_0786_),
    .Y(_0188_),
    .B1(_0780_));
 sg13g2_nor2_1 _2408_ (.A(net94),
    .B(net520),
    .Y(_0787_));
 sg13g2_nor2b_1 _2409_ (.A(\cic_a.temp_comb[1][7] ),
    .B_N(\cic_a.delay[2][7] ),
    .Y(_0788_));
 sg13g2_nand2b_1 _2410_ (.Y(_0789_),
    .B(\cic_a.temp_comb[1][7] ),
    .A_N(\cic_a.delay[2][7] ));
 sg13g2_nand2b_1 _2411_ (.Y(_0790_),
    .B(_0789_),
    .A_N(_0788_));
 sg13g2_o21ai_1 _2412_ (.B1(_0781_),
    .Y(_0791_),
    .A1(_0782_),
    .A2(_0785_));
 sg13g2_xor2_1 _2413_ (.B(_0791_),
    .A(_0790_),
    .X(_0792_));
 sg13g2_a21oi_1 _2414_ (.A1(net520),
    .A2(_0792_),
    .Y(_0189_),
    .B1(_0787_));
 sg13g2_nor2_1 _2415_ (.A(_0782_),
    .B(_0790_),
    .Y(_0793_));
 sg13g2_and2_1 _2416_ (.A(_0783_),
    .B(_0793_),
    .X(_0794_));
 sg13g2_o21ai_1 _2417_ (.B1(_0789_),
    .Y(_0795_),
    .A1(_0781_),
    .A2(_0788_));
 sg13g2_a221oi_1 _2418_ (.B2(_0769_),
    .C1(_0795_),
    .B1(_0794_),
    .A1(_0784_),
    .Y(_0796_),
    .A2(_0793_));
 sg13g2_nor2b_1 _2419_ (.A(\cic_a.delay[2][8] ),
    .B_N(\cic_a.temp_comb[1][8] ),
    .Y(_0797_));
 sg13g2_xor2_1 _2420_ (.B(\cic_a.delay[2][8] ),
    .A(\cic_a.temp_comb[1][8] ),
    .X(_0798_));
 sg13g2_nor2_1 _2421_ (.A(_0796_),
    .B(_0798_),
    .Y(_0799_));
 sg13g2_xnor2_1 _2422_ (.Y(_0800_),
    .A(_0796_),
    .B(_0798_));
 sg13g2_nor2_1 _2423_ (.A(net270),
    .B(net517),
    .Y(_0801_));
 sg13g2_a21oi_1 _2424_ (.A1(net517),
    .A2(_0800_),
    .Y(_0190_),
    .B1(_0801_));
 sg13g2_nor2b_1 _2425_ (.A(\cic_a.delay[2][9] ),
    .B_N(\cic_a.temp_comb[1][9] ),
    .Y(_0802_));
 sg13g2_nand2b_1 _2426_ (.Y(_0803_),
    .B(\cic_a.delay[2][9] ),
    .A_N(\cic_a.temp_comb[1][9] ));
 sg13g2_nor2b_1 _2427_ (.A(_0802_),
    .B_N(_0803_),
    .Y(_0804_));
 sg13g2_nor2_1 _2428_ (.A(_0797_),
    .B(_0799_),
    .Y(_0805_));
 sg13g2_xnor2_1 _2429_ (.Y(_0806_),
    .A(_0804_),
    .B(_0805_));
 sg13g2_mux2_1 _2430_ (.A0(net265),
    .A1(_0806_),
    .S(net527),
    .X(_0191_));
 sg13g2_nor2_1 _2431_ (.A(net439),
    .B(net517),
    .Y(_0807_));
 sg13g2_nand2b_1 _2432_ (.Y(_0808_),
    .B(_0804_),
    .A_N(_0798_));
 sg13g2_a21oi_1 _2433_ (.A1(_0797_),
    .A2(_0803_),
    .Y(_0809_),
    .B1(_0802_));
 sg13g2_o21ai_1 _2434_ (.B1(_0809_),
    .Y(_0810_),
    .A1(_0796_),
    .A2(_0808_));
 sg13g2_nor2b_1 _2435_ (.A(\cic_a.delay[2][10] ),
    .B_N(\cic_a.temp_comb[1][10] ),
    .Y(_0811_));
 sg13g2_nor2b_1 _2436_ (.A(\cic_a.temp_comb[1][10] ),
    .B_N(\cic_a.delay[2][10] ),
    .Y(_0812_));
 sg13g2_nor2_1 _2437_ (.A(_0811_),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_xnor2_1 _2438_ (.Y(_0814_),
    .A(_0810_),
    .B(_0813_));
 sg13g2_a21oi_1 _2439_ (.A1(net517),
    .A2(_0814_),
    .Y(_0192_),
    .B1(_0807_));
 sg13g2_nor2b_1 _2440_ (.A(\cic_a.delay[2][11] ),
    .B_N(\cic_a.temp_comb[1][11] ),
    .Y(_0815_));
 sg13g2_nand2b_1 _2441_ (.Y(_0816_),
    .B(\cic_a.delay[2][11] ),
    .A_N(\cic_a.temp_comb[1][11] ));
 sg13g2_nand2b_1 _2442_ (.Y(_0817_),
    .B(_0816_),
    .A_N(_0815_));
 sg13g2_a21oi_1 _2443_ (.A1(_0810_),
    .A2(_0813_),
    .Y(_0818_),
    .B1(_0811_));
 sg13g2_xor2_1 _2444_ (.B(_0818_),
    .A(_0817_),
    .X(_0819_));
 sg13g2_mux2_1 _2445_ (.A0(net191),
    .A1(_0819_),
    .S(net517),
    .X(_0193_));
 sg13g2_nor2_1 _2446_ (.A(net412),
    .B(net518),
    .Y(_0820_));
 sg13g2_nor3_1 _2447_ (.A(_0811_),
    .B(_0812_),
    .C(_0817_),
    .Y(_0821_));
 sg13g2_a221oi_1 _2448_ (.B2(_0810_),
    .C1(_0815_),
    .B1(_0821_),
    .A1(_0811_),
    .Y(_0822_),
    .A2(_0816_));
 sg13g2_xor2_1 _2449_ (.B(\cic_a.delay[2][12] ),
    .A(\cic_a.temp_comb[1][12] ),
    .X(_0823_));
 sg13g2_xnor2_1 _2450_ (.Y(_0824_),
    .A(_0822_),
    .B(_0823_));
 sg13g2_a21oi_1 _2451_ (.A1(net528),
    .A2(_0824_),
    .Y(_0194_),
    .B1(_0820_));
 sg13g2_mux2_1 _2452_ (.A0(net197),
    .A1(\cic_a.integrator[2][0] ),
    .S(net518),
    .X(_0195_));
 sg13g2_mux2_1 _2453_ (.A0(net237),
    .A1(\cic_a.integrator[2][1] ),
    .S(net518),
    .X(_0196_));
 sg13g2_mux2_1 _2454_ (.A0(net110),
    .A1(net188),
    .S(net518),
    .X(_0197_));
 sg13g2_mux2_1 _2455_ (.A0(net141),
    .A1(net144),
    .S(net513),
    .X(_0198_));
 sg13g2_mux2_1 _2456_ (.A0(net344),
    .A1(\cic_a.integrator[2][4] ),
    .S(net512),
    .X(_0199_));
 sg13g2_mux2_1 _2457_ (.A0(net22),
    .A1(net158),
    .S(net508),
    .X(_0200_));
 sg13g2_mux2_1 _2458_ (.A0(net327),
    .A1(\cic_a.integrator[2][6] ),
    .S(net502),
    .X(_0201_));
 sg13g2_mux2_1 _2459_ (.A0(net41),
    .A1(net276),
    .S(net502),
    .X(_0202_));
 sg13g2_mux2_1 _2460_ (.A0(net189),
    .A1(\cic_a.integrator[2][8] ),
    .S(net502),
    .X(_0203_));
 sg13g2_nor2_1 _2461_ (.A(net98),
    .B(net500),
    .Y(_0825_));
 sg13g2_a21oi_1 _2462_ (.A1(_1215_),
    .A2(net500),
    .Y(_0204_),
    .B1(_0825_));
 sg13g2_mux2_1 _2463_ (.A0(net54),
    .A1(net250),
    .S(net503),
    .X(_0205_));
 sg13g2_mux2_1 _2464_ (.A0(net227),
    .A1(\cic_a.integrator[2][11] ),
    .S(net503),
    .X(_0206_));
 sg13g2_mux2_1 _2465_ (.A0(net306),
    .A1(\cic_a.integrator[2][12] ),
    .S(net503),
    .X(_0207_));
 sg13g2_mux2_1 _2466_ (.A0(net128),
    .A1(\cic_a.temp_comb[0][0] ),
    .S(net521),
    .X(_0208_));
 sg13g2_mux2_1 _2467_ (.A0(net309),
    .A1(\cic_a.temp_comb[0][1] ),
    .S(net522),
    .X(_0209_));
 sg13g2_mux2_1 _2468_ (.A0(net167),
    .A1(\cic_a.temp_comb[0][2] ),
    .S(net519),
    .X(_0210_));
 sg13g2_mux2_1 _2469_ (.A0(net156),
    .A1(\cic_a.temp_comb[0][3] ),
    .S(net515),
    .X(_0211_));
 sg13g2_mux2_1 _2470_ (.A0(net393),
    .A1(\cic_a.temp_comb[0][4] ),
    .S(net509),
    .X(_0212_));
 sg13g2_mux2_1 _2471_ (.A0(net225),
    .A1(\cic_a.temp_comb[0][5] ),
    .S(net510),
    .X(_0213_));
 sg13g2_mux2_1 _2472_ (.A0(net139),
    .A1(net171),
    .S(net510),
    .X(_0214_));
 sg13g2_mux2_1 _2473_ (.A0(net252),
    .A1(\cic_a.temp_comb[0][7] ),
    .S(net510),
    .X(_0215_));
 sg13g2_mux2_1 _2474_ (.A0(net364),
    .A1(\cic_a.temp_comb[0][8] ),
    .S(net506),
    .X(_0216_));
 sg13g2_nor2_1 _2475_ (.A(net50),
    .B(net506),
    .Y(_0826_));
 sg13g2_a21oi_1 _2476_ (.A1(_1217_),
    .A2(net506),
    .Y(_0217_),
    .B1(_0826_));
 sg13g2_mux2_1 _2477_ (.A0(net274),
    .A1(\cic_a.temp_comb[0][10] ),
    .S(net501),
    .X(_0218_));
 sg13g2_mux2_1 _2478_ (.A0(net281),
    .A1(\cic_a.temp_comb[0][11] ),
    .S(net501),
    .X(_0219_));
 sg13g2_mux2_1 _2479_ (.A0(net165),
    .A1(\cic_a.temp_comb[0][12] ),
    .S(net500),
    .X(_0220_));
 sg13g2_mux2_1 _2480_ (.A0(net216),
    .A1(net201),
    .S(net495),
    .X(_0221_));
 sg13g2_mux2_1 _2481_ (.A0(net403),
    .A1(net319),
    .S(net496),
    .X(_0222_));
 sg13g2_mux2_1 _2482_ (.A0(net312),
    .A1(net219),
    .S(net495),
    .X(_0223_));
 sg13g2_mux2_1 _2483_ (.A0(net383),
    .A1(net248),
    .S(net498),
    .X(_0224_));
 sg13g2_mux2_1 _2484_ (.A0(net161),
    .A1(net272),
    .S(net487),
    .X(_0225_));
 sg13g2_mux2_1 _2485_ (.A0(net349),
    .A1(net266),
    .S(net487),
    .X(_0226_));
 sg13g2_mux2_1 _2486_ (.A0(net384),
    .A1(net256),
    .S(net489),
    .X(_0227_));
 sg13g2_mux2_1 _2487_ (.A0(net372),
    .A1(net366),
    .S(net489),
    .X(_0228_));
 sg13g2_mux2_1 _2488_ (.A0(net341),
    .A1(net322),
    .S(net477),
    .X(_0229_));
 sg13g2_nand2_1 _2489_ (.Y(_0827_),
    .A(net37),
    .B(net477));
 sg13g2_o21ai_1 _2490_ (.B1(_0827_),
    .Y(_0230_),
    .A1(_1228_),
    .A2(net477));
 sg13g2_mux2_1 _2491_ (.A0(net251),
    .A1(net241),
    .S(net480),
    .X(_0231_));
 sg13g2_mux2_1 _2492_ (.A0(\cic_b.delay[2][11] ),
    .A1(net316),
    .S(net480),
    .X(_0232_));
 sg13g2_mux2_1 _2493_ (.A0(net363),
    .A1(net342),
    .S(net473),
    .X(_0233_));
 sg13g2_nor2_1 _2494_ (.A(net642),
    .B(net495),
    .Y(_0828_));
 sg13g2_nand2b_1 _2495_ (.Y(_0829_),
    .B(net358),
    .A_N(\cic_b.temp_comb[0][0] ));
 sg13g2_xnor2_1 _2496_ (.Y(_0830_),
    .A(\cic_b.temp_comb[0][0] ),
    .B(net358));
 sg13g2_a21oi_1 _2497_ (.A1(net496),
    .A2(_0830_),
    .Y(_0234_),
    .B1(_0828_));
 sg13g2_nor2_1 _2498_ (.A(net644),
    .B(net496),
    .Y(_0831_));
 sg13g2_nor2b_1 _2499_ (.A(\cic_b.delay[1][1] ),
    .B_N(\cic_b.temp_comb[0][1] ),
    .Y(_0832_));
 sg13g2_xnor2_1 _2500_ (.Y(_0833_),
    .A(\cic_b.temp_comb[0][1] ),
    .B(net359));
 sg13g2_xnor2_1 _2501_ (.Y(_0834_),
    .A(_0829_),
    .B(_0833_));
 sg13g2_a21oi_1 _2502_ (.A1(net495),
    .A2(_0834_),
    .Y(_0235_),
    .B1(_0831_));
 sg13g2_nor2_1 _2503_ (.A(net470),
    .B(net495),
    .Y(_0835_));
 sg13g2_nor2b_1 _2504_ (.A(\cic_b.delay[1][2] ),
    .B_N(\cic_b.temp_comb[0][2] ),
    .Y(_0836_));
 sg13g2_nand2b_1 _2505_ (.Y(_0837_),
    .B(net308),
    .A_N(\cic_b.temp_comb[0][2] ));
 sg13g2_nor2b_1 _2506_ (.A(_0836_),
    .B_N(_0837_),
    .Y(_0838_));
 sg13g2_a21o_1 _2507_ (.A2(_0833_),
    .A1(_0829_),
    .B1(_0832_),
    .X(_0839_));
 sg13g2_xnor2_1 _2508_ (.Y(_0840_),
    .A(_0838_),
    .B(_0839_));
 sg13g2_a21oi_1 _2509_ (.A1(net491),
    .A2(_0840_),
    .Y(_0236_),
    .B1(_0835_));
 sg13g2_nor2_1 _2510_ (.A(net681),
    .B(net494),
    .Y(_0841_));
 sg13g2_nand2b_1 _2511_ (.Y(_0842_),
    .B(\cic_b.temp_comb[0][3] ),
    .A_N(\cic_b.delay[1][3] ));
 sg13g2_xor2_1 _2512_ (.B(net402),
    .A(\cic_b.temp_comb[0][3] ),
    .X(_0843_));
 sg13g2_a21oi_2 _2513_ (.B1(_0836_),
    .Y(_0844_),
    .A2(_0839_),
    .A1(_0837_));
 sg13g2_xnor2_1 _2514_ (.Y(_0845_),
    .A(_0843_),
    .B(_0844_));
 sg13g2_a21oi_1 _2515_ (.A1(net494),
    .A2(_0845_),
    .Y(_0237_),
    .B1(_0841_));
 sg13g2_o21ai_1 _2516_ (.B1(_0842_),
    .Y(_0846_),
    .A1(_0843_),
    .A2(_0844_));
 sg13g2_nand2_1 _2517_ (.Y(_0847_),
    .A(\cic_b.temp_comb[0][4] ),
    .B(_1229_));
 sg13g2_xor2_1 _2518_ (.B(\cic_b.delay[1][4] ),
    .A(\cic_b.temp_comb[0][4] ),
    .X(_0848_));
 sg13g2_nand2b_1 _2519_ (.Y(_0849_),
    .B(_0846_),
    .A_N(_0848_));
 sg13g2_nor2_1 _2520_ (.A(net640),
    .B(net488),
    .Y(_0850_));
 sg13g2_xor2_1 _2521_ (.B(_0848_),
    .A(_0846_),
    .X(_0851_));
 sg13g2_a21oi_1 _2522_ (.A1(net484),
    .A2(_0851_),
    .Y(_0238_),
    .B1(_0850_));
 sg13g2_nor2_1 _2523_ (.A(net687),
    .B(net484),
    .Y(_0852_));
 sg13g2_nor2b_1 _2524_ (.A(\cic_b.temp_comb[0][5] ),
    .B_N(\cic_b.delay[1][5] ),
    .Y(_0853_));
 sg13g2_nand2b_1 _2525_ (.Y(_0854_),
    .B(\cic_b.temp_comb[0][5] ),
    .A_N(\cic_b.delay[1][5] ));
 sg13g2_nand2b_1 _2526_ (.Y(_0855_),
    .B(_0854_),
    .A_N(_0853_));
 sg13g2_and2_1 _2527_ (.A(_0847_),
    .B(_0849_),
    .X(_0856_));
 sg13g2_xnor2_1 _2528_ (.Y(_0857_),
    .A(_0855_),
    .B(_0856_));
 sg13g2_a21oi_1 _2529_ (.A1(net484),
    .A2(_0857_),
    .Y(_0239_),
    .B1(_0852_));
 sg13g2_nor2_1 _2530_ (.A(net664),
    .B(net483),
    .Y(_0858_));
 sg13g2_nand2b_1 _2531_ (.Y(_0859_),
    .B(\cic_b.temp_comb[0][6] ),
    .A_N(\cic_b.delay[1][6] ));
 sg13g2_xor2_1 _2532_ (.B(net423),
    .A(\cic_b.temp_comb[0][6] ),
    .X(_0860_));
 sg13g2_nor2_1 _2533_ (.A(_0848_),
    .B(_0855_),
    .Y(_0861_));
 sg13g2_o21ai_1 _2534_ (.B1(_0854_),
    .Y(_0862_),
    .A1(_0847_),
    .A2(_0853_));
 sg13g2_a21oi_1 _2535_ (.A1(_0846_),
    .A2(_0861_),
    .Y(_0863_),
    .B1(_0862_));
 sg13g2_xnor2_1 _2536_ (.Y(_0864_),
    .A(_0860_),
    .B(_0863_));
 sg13g2_a21oi_1 _2537_ (.A1(net483),
    .A2(_0864_),
    .Y(_0240_),
    .B1(_0858_));
 sg13g2_nor2_1 _2538_ (.A(net466),
    .B(net482),
    .Y(_0865_));
 sg13g2_nor2b_1 _2539_ (.A(\cic_b.temp_comb[0][7] ),
    .B_N(\cic_b.delay[1][7] ),
    .Y(_0866_));
 sg13g2_nand2b_1 _2540_ (.Y(_0867_),
    .B(\cic_b.temp_comb[0][7] ),
    .A_N(\cic_b.delay[1][7] ));
 sg13g2_nand2b_1 _2541_ (.Y(_0868_),
    .B(_0867_),
    .A_N(_0866_));
 sg13g2_o21ai_1 _2542_ (.B1(_0859_),
    .Y(_0869_),
    .A1(_0860_),
    .A2(_0863_));
 sg13g2_xor2_1 _2543_ (.B(_0869_),
    .A(_0868_),
    .X(_0870_));
 sg13g2_a21oi_1 _2544_ (.A1(net482),
    .A2(_0870_),
    .Y(_0241_),
    .B1(_0865_));
 sg13g2_o21ai_1 _2545_ (.B1(_0867_),
    .Y(_0871_),
    .A1(_0859_),
    .A2(_0866_));
 sg13g2_nor2_1 _2546_ (.A(_0860_),
    .B(_0868_),
    .Y(_0872_));
 sg13g2_and2_1 _2547_ (.A(_0861_),
    .B(_0872_),
    .X(_0873_));
 sg13g2_a221oi_1 _2548_ (.B2(_0846_),
    .C1(_0871_),
    .B1(_0873_),
    .A1(_0862_),
    .Y(_0874_),
    .A2(_0872_));
 sg13g2_nand2b_1 _2549_ (.Y(_0875_),
    .B(net792),
    .A_N(\cic_b.delay[1][8] ));
 sg13g2_xor2_1 _2550_ (.B(net303),
    .A(net791),
    .X(_0876_));
 sg13g2_xnor2_1 _2551_ (.Y(_0877_),
    .A(_0874_),
    .B(_0876_));
 sg13g2_nor2_1 _2552_ (.A(net639),
    .B(net479),
    .Y(_0878_));
 sg13g2_a21oi_1 _2553_ (.A1(net477),
    .A2(_0877_),
    .Y(_0242_),
    .B1(_0878_));
 sg13g2_nor2_1 _2554_ (.A(net162),
    .B(net477),
    .Y(_0879_));
 sg13g2_xor2_1 _2555_ (.B(\cic_b.delay[1][9] ),
    .A(net621),
    .X(_0880_));
 sg13g2_o21ai_1 _2556_ (.B1(_0875_),
    .Y(_0881_),
    .A1(_0874_),
    .A2(_0876_));
 sg13g2_xor2_1 _2557_ (.B(_0881_),
    .A(net622),
    .X(_0882_));
 sg13g2_a21oi_1 _2558_ (.A1(net477),
    .A2(_0882_),
    .Y(_0243_),
    .B1(_0879_));
 sg13g2_nor2_1 _2559_ (.A(net457),
    .B(net480),
    .Y(_0883_));
 sg13g2_or2_1 _2560_ (.X(_0884_),
    .B(_0880_),
    .A(_0876_));
 sg13g2_a21oi_1 _2561_ (.A1(_1230_),
    .A2(\cic_b.delay[1][9] ),
    .Y(_0885_),
    .B1(_0875_));
 sg13g2_a21oi_1 _2562_ (.A1(\cic_b.temp_comb[0][9] ),
    .A2(_1231_),
    .Y(_0886_),
    .B1(_0885_));
 sg13g2_o21ai_1 _2563_ (.B1(_0886_),
    .Y(_0887_),
    .A1(_0874_),
    .A2(_0884_));
 sg13g2_nor2b_1 _2564_ (.A(\cic_b.delay[1][10] ),
    .B_N(\cic_b.temp_comb[0][10] ),
    .Y(_0888_));
 sg13g2_xnor2_1 _2565_ (.Y(_0889_),
    .A(\cic_b.temp_comb[0][10] ),
    .B(\cic_b.delay[1][10] ));
 sg13g2_inv_1 _2566_ (.Y(_0890_),
    .A(_0889_));
 sg13g2_xnor2_1 _2567_ (.Y(_0891_),
    .A(_0887_),
    .B(_0889_));
 sg13g2_a21oi_1 _2568_ (.A1(net480),
    .A2(_0891_),
    .Y(_0244_),
    .B1(_0883_));
 sg13g2_nor2_1 _2569_ (.A(net318),
    .B(net480),
    .Y(_0892_));
 sg13g2_nor2b_1 _2570_ (.A(\cic_b.delay[1][11] ),
    .B_N(\cic_b.temp_comb[0][11] ),
    .Y(_0893_));
 sg13g2_nand2b_1 _2571_ (.Y(_0894_),
    .B(\cic_b.delay[1][11] ),
    .A_N(\cic_b.temp_comb[0][11] ));
 sg13g2_nand2b_1 _2572_ (.Y(_0895_),
    .B(_0894_),
    .A_N(_0893_));
 sg13g2_a21oi_1 _2573_ (.A1(_0887_),
    .A2(_0889_),
    .Y(_0896_),
    .B1(_0888_));
 sg13g2_xnor2_1 _2574_ (.Y(_0897_),
    .A(_0895_),
    .B(_0896_));
 sg13g2_a21oi_1 _2575_ (.A1(net480),
    .A2(_0897_),
    .Y(_0245_),
    .B1(_0892_));
 sg13g2_nor2_1 _2576_ (.A(net461),
    .B(net473),
    .Y(_0898_));
 sg13g2_nor2_1 _2577_ (.A(_0890_),
    .B(_0895_),
    .Y(_0899_));
 sg13g2_a221oi_1 _2578_ (.B2(_0887_),
    .C1(_0893_),
    .B1(_0899_),
    .A1(_0888_),
    .Y(_0900_),
    .A2(_0894_));
 sg13g2_xor2_1 _2579_ (.B(\cic_b.delay[1][12] ),
    .A(net347),
    .X(_0901_));
 sg13g2_xnor2_1 _2580_ (.Y(_0902_),
    .A(_0900_),
    .B(_0901_));
 sg13g2_a21oi_1 _2581_ (.A1(net471),
    .A2(_0902_),
    .Y(_0246_),
    .B1(_0898_));
 sg13g2_mux2_1 _2582_ (.A0(net358),
    .A1(net205),
    .S(net491),
    .X(_0247_));
 sg13g2_mux2_1 _2583_ (.A0(net359),
    .A1(net336),
    .S(net492),
    .X(_0248_));
 sg13g2_mux2_1 _2584_ (.A0(net308),
    .A1(net182),
    .S(net491),
    .X(_0249_));
 sg13g2_mux2_1 _2585_ (.A0(net402),
    .A1(net268),
    .S(net494),
    .X(_0250_));
 sg13g2_nand2_1 _2586_ (.Y(_0903_),
    .A(net27),
    .B(net486));
 sg13g2_o21ai_1 _2587_ (.B1(_0903_),
    .Y(_0251_),
    .A1(_1229_),
    .A2(net486));
 sg13g2_mux2_1 _2588_ (.A0(net333),
    .A1(net304),
    .S(net484),
    .X(_0252_));
 sg13g2_mux2_1 _2589_ (.A0(net423),
    .A1(net330),
    .S(net482),
    .X(_0253_));
 sg13g2_mux2_1 _2590_ (.A0(net332),
    .A1(net233),
    .S(net476),
    .X(_0254_));
 sg13g2_mux2_1 _2591_ (.A0(net303),
    .A1(net179),
    .S(net476),
    .X(_0255_));
 sg13g2_nand2_1 _2592_ (.Y(_0904_),
    .A(net89),
    .B(net474));
 sg13g2_o21ai_1 _2593_ (.B1(_0904_),
    .Y(_0256_),
    .A1(_1231_),
    .A2(net474));
 sg13g2_mux2_1 _2594_ (.A0(\cic_b.delay[1][10] ),
    .A1(net279),
    .S(net474),
    .X(_0257_));
 sg13g2_mux2_1 _2595_ (.A0(\cic_b.delay[1][11] ),
    .A1(net146),
    .S(net471),
    .X(_0258_));
 sg13g2_mux2_1 _2596_ (.A0(\cic_b.delay[1][12] ),
    .A1(net148),
    .S(net472),
    .X(_0259_));
 sg13g2_mux2_1 _2597_ (.A0(net311),
    .A1(net299),
    .S(net493),
    .X(_0260_));
 sg13g2_mux2_1 _2598_ (.A0(\cic_b.delay[0][1] ),
    .A1(net199),
    .S(net493),
    .X(_0261_));
 sg13g2_mux2_1 _2599_ (.A0(net399),
    .A1(net239),
    .S(net493),
    .X(_0262_));
 sg13g2_mux2_1 _2600_ (.A0(net321),
    .A1(net297),
    .S(net494),
    .X(_0263_));
 sg13g2_mux2_1 _2601_ (.A0(net425),
    .A1(net385),
    .S(net485),
    .X(_0264_));
 sg13g2_nand2_1 _2602_ (.Y(_0905_),
    .A(net43),
    .B(net485));
 sg13g2_o21ai_1 _2603_ (.B1(_0905_),
    .Y(_0265_),
    .A1(_1224_),
    .A2(net485));
 sg13g2_mux2_1 _2604_ (.A0(net434),
    .A1(net223),
    .S(net483),
    .X(_0266_));
 sg13g2_mux2_1 _2605_ (.A0(net371),
    .A1(net301),
    .S(net476),
    .X(_0267_));
 sg13g2_mux2_1 _2606_ (.A0(net324),
    .A1(net229),
    .S(net475),
    .X(_0268_));
 sg13g2_nand2_1 _2607_ (.Y(_0906_),
    .A(net58),
    .B(net475));
 sg13g2_o21ai_1 _2608_ (.B1(_0906_),
    .Y(_0269_),
    .A1(_1226_),
    .A2(net475));
 sg13g2_mux2_1 _2609_ (.A0(net416),
    .A1(net235),
    .S(net471),
    .X(_0270_));
 sg13g2_mux2_1 _2610_ (.A0(\cic_b.delay[0][11] ),
    .A1(net20),
    .S(net471),
    .X(_0271_));
 sg13g2_mux2_1 _2611_ (.A0(\cic_b.delay[0][12] ),
    .A1(net186),
    .S(net472),
    .X(_0272_));
 sg13g2_nor2_1 _2612_ (.A(net655),
    .B(net492),
    .Y(_0907_));
 sg13g2_nor2b_1 _2613_ (.A(\cic_b.integrator[2][0] ),
    .B_N(net311),
    .Y(_0908_));
 sg13g2_xnor2_1 _2614_ (.Y(_0909_),
    .A(\cic_b.integrator[2][0] ),
    .B(net311));
 sg13g2_a21oi_1 _2615_ (.A1(net491),
    .A2(_0909_),
    .Y(_0273_),
    .B1(_0907_));
 sg13g2_nor2_1 _2616_ (.A(net636),
    .B(net491),
    .Y(_0910_));
 sg13g2_nand2b_1 _2617_ (.Y(_0911_),
    .B(\cic_b.integrator[2][1] ),
    .A_N(\cic_b.delay[0][1] ));
 sg13g2_xor2_1 _2618_ (.B(\cic_b.delay[0][1] ),
    .A(\cic_b.integrator[2][1] ),
    .X(_0912_));
 sg13g2_xnor2_1 _2619_ (.Y(_0913_),
    .A(_0908_),
    .B(_0912_));
 sg13g2_a21oi_1 _2620_ (.A1(net492),
    .A2(_0913_),
    .Y(_0274_),
    .B1(_0910_));
 sg13g2_nor2_1 _2621_ (.A(net468),
    .B(net491),
    .Y(_0914_));
 sg13g2_nor2b_1 _2622_ (.A(net399),
    .B_N(\cic_b.integrator[2][2] ),
    .Y(_0915_));
 sg13g2_xnor2_1 _2623_ (.Y(_0916_),
    .A(\cic_b.integrator[2][2] ),
    .B(\cic_b.delay[0][2] ));
 sg13g2_o21ai_1 _2624_ (.B1(_0911_),
    .Y(_0917_),
    .A1(_0908_),
    .A2(_0912_));
 sg13g2_xnor2_1 _2625_ (.Y(_0918_),
    .A(_0916_),
    .B(_0917_));
 sg13g2_a21oi_1 _2626_ (.A1(net493),
    .A2(_0918_),
    .Y(_0275_),
    .B1(_0914_));
 sg13g2_nor2_1 _2627_ (.A(net679),
    .B(net494),
    .Y(_0919_));
 sg13g2_nand2b_1 _2628_ (.Y(_0920_),
    .B(\cic_b.integrator[2][3] ),
    .A_N(\cic_b.delay[0][3] ));
 sg13g2_xor2_1 _2629_ (.B(net321),
    .A(\cic_b.integrator[2][3] ),
    .X(_0921_));
 sg13g2_a21oi_2 _2630_ (.B1(_0915_),
    .Y(_0922_),
    .A2(_0917_),
    .A1(_0916_));
 sg13g2_xnor2_1 _2631_ (.Y(_0923_),
    .A(_0921_),
    .B(_0922_));
 sg13g2_a21oi_1 _2632_ (.A1(net494),
    .A2(_0923_),
    .Y(_0276_),
    .B1(_0919_));
 sg13g2_o21ai_1 _2633_ (.B1(_0920_),
    .Y(_0924_),
    .A1(_0921_),
    .A2(_0922_));
 sg13g2_nor2b_1 _2634_ (.A(\cic_b.delay[0][4] ),
    .B_N(\cic_b.integrator[2][4] ),
    .Y(_0925_));
 sg13g2_xor2_1 _2635_ (.B(\cic_b.delay[0][4] ),
    .A(\cic_b.integrator[2][4] ),
    .X(_0926_));
 sg13g2_nor2b_1 _2636_ (.A(_0926_),
    .B_N(_0924_),
    .Y(_0927_));
 sg13g2_nor2_1 _2637_ (.A(net143),
    .B(net484),
    .Y(_0928_));
 sg13g2_xor2_1 _2638_ (.B(_0926_),
    .A(_0924_),
    .X(_0929_));
 sg13g2_a21oi_1 _2639_ (.A1(net485),
    .A2(_0929_),
    .Y(_0277_),
    .B1(_0928_));
 sg13g2_nor2_1 _2640_ (.A(net633),
    .B(net484),
    .Y(_0930_));
 sg13g2_xor2_1 _2641_ (.B(\cic_b.delay[0][5] ),
    .A(\cic_b.integrator[2][5] ),
    .X(_0931_));
 sg13g2_nor2_1 _2642_ (.A(_0925_),
    .B(_0927_),
    .Y(_0932_));
 sg13g2_xnor2_1 _2643_ (.Y(_0933_),
    .A(_0931_),
    .B(_0932_));
 sg13g2_a21oi_1 _2644_ (.A1(net485),
    .A2(_0933_),
    .Y(_0278_),
    .B1(_0930_));
 sg13g2_nor2_1 _2645_ (.A(net674),
    .B(net482),
    .Y(_0934_));
 sg13g2_nand2b_1 _2646_ (.Y(_0935_),
    .B(\cic_b.integrator[2][6] ),
    .A_N(\cic_b.delay[0][6] ));
 sg13g2_xor2_1 _2647_ (.B(\cic_b.delay[0][6] ),
    .A(\cic_b.integrator[2][6] ),
    .X(_0936_));
 sg13g2_a21oi_1 _2648_ (.A1(\cic_b.integrator[2][5] ),
    .A2(_1224_),
    .Y(_0937_),
    .B1(_0925_));
 sg13g2_a21oi_1 _2649_ (.A1(_1223_),
    .A2(\cic_b.delay[0][5] ),
    .Y(_0938_),
    .B1(_0937_));
 sg13g2_nor2_1 _2650_ (.A(_0926_),
    .B(_0931_),
    .Y(_0939_));
 sg13g2_a21oi_1 _2651_ (.A1(_0924_),
    .A2(_0939_),
    .Y(_0940_),
    .B1(_0938_));
 sg13g2_xnor2_1 _2652_ (.Y(_0941_),
    .A(_0936_),
    .B(_0940_));
 sg13g2_a21oi_1 _2653_ (.A1(net483),
    .A2(_0941_),
    .Y(_0279_),
    .B1(_0934_));
 sg13g2_nor2b_1 _2654_ (.A(\cic_b.integrator[2][7] ),
    .B_N(\cic_b.delay[0][7] ),
    .Y(_0942_));
 sg13g2_nand2b_1 _2655_ (.Y(_0943_),
    .B(\cic_b.integrator[2][7] ),
    .A_N(\cic_b.delay[0][7] ));
 sg13g2_nand2b_1 _2656_ (.Y(_0944_),
    .B(_0943_),
    .A_N(_0942_));
 sg13g2_o21ai_1 _2657_ (.B1(_0935_),
    .Y(_0945_),
    .A1(_0936_),
    .A2(_0940_));
 sg13g2_xor2_1 _2658_ (.B(_0945_),
    .A(_0944_),
    .X(_0946_));
 sg13g2_nor2_1 _2659_ (.A(net638),
    .B(net482),
    .Y(_0947_));
 sg13g2_a21oi_1 _2660_ (.A1(net483),
    .A2(_0946_),
    .Y(_0280_),
    .B1(_0947_));
 sg13g2_nor2_1 _2661_ (.A(_0936_),
    .B(_0944_),
    .Y(_0948_));
 sg13g2_nor4_1 _2662_ (.A(_0926_),
    .B(_0931_),
    .C(_0936_),
    .D(_0944_),
    .Y(_0949_));
 sg13g2_o21ai_1 _2663_ (.B1(_0943_),
    .Y(_0950_),
    .A1(_0935_),
    .A2(_0942_));
 sg13g2_a221oi_1 _2664_ (.B2(_0924_),
    .C1(_0950_),
    .B1(_0949_),
    .A1(_0938_),
    .Y(_0951_),
    .A2(_0948_));
 sg13g2_nand2b_1 _2665_ (.Y(_0952_),
    .B(\cic_b.integrator[2][8] ),
    .A_N(\cic_b.delay[0][8] ));
 sg13g2_xor2_1 _2666_ (.B(net324),
    .A(\cic_b.integrator[2][8] ),
    .X(_0953_));
 sg13g2_xnor2_1 _2667_ (.Y(_0954_),
    .A(_0951_),
    .B(_0953_));
 sg13g2_nor2_1 _2668_ (.A(net651),
    .B(net476),
    .Y(_0955_));
 sg13g2_a21oi_1 _2669_ (.A1(net475),
    .A2(_0954_),
    .Y(_0281_),
    .B1(_0955_));
 sg13g2_nor2_1 _2670_ (.A(net422),
    .B(net474),
    .Y(_0956_));
 sg13g2_xnor2_1 _2671_ (.Y(_0957_),
    .A(\cic_b.integrator[2][9] ),
    .B(net650));
 sg13g2_o21ai_1 _2672_ (.B1(_0952_),
    .Y(_0958_),
    .A1(_0951_),
    .A2(_0953_));
 sg13g2_xnor2_1 _2673_ (.Y(_0959_),
    .A(_0957_),
    .B(_0958_));
 sg13g2_a21oi_1 _2674_ (.A1(net474),
    .A2(_0959_),
    .Y(_0282_),
    .B1(_0956_));
 sg13g2_nor2_1 _2675_ (.A(net283),
    .B(net471),
    .Y(_0960_));
 sg13g2_nand2b_1 _2676_ (.Y(_0961_),
    .B(_0957_),
    .A_N(_0953_));
 sg13g2_a21oi_1 _2677_ (.A1(_1225_),
    .A2(\cic_b.delay[0][9] ),
    .Y(_0962_),
    .B1(_0952_));
 sg13g2_a21oi_1 _2678_ (.A1(\cic_b.integrator[2][9] ),
    .A2(_1226_),
    .Y(_0963_),
    .B1(_0962_));
 sg13g2_o21ai_1 _2679_ (.B1(_0963_),
    .Y(_0964_),
    .A1(_0951_),
    .A2(_0961_));
 sg13g2_nor2b_1 _2680_ (.A(\cic_b.delay[0][10] ),
    .B_N(\cic_b.integrator[2][10] ),
    .Y(_0965_));
 sg13g2_nor2b_1 _2681_ (.A(\cic_b.integrator[2][10] ),
    .B_N(\cic_b.delay[0][10] ),
    .Y(_0966_));
 sg13g2_nor2_1 _2682_ (.A(_0965_),
    .B(_0966_),
    .Y(_0967_));
 sg13g2_xnor2_1 _2683_ (.Y(_0968_),
    .A(_0964_),
    .B(_0967_));
 sg13g2_a21oi_1 _2684_ (.A1(net473),
    .A2(_0968_),
    .Y(_0283_),
    .B1(_0960_));
 sg13g2_nor2b_1 _2685_ (.A(\cic_b.delay[0][11] ),
    .B_N(\cic_b.integrator[2][11] ),
    .Y(_0969_));
 sg13g2_nand2b_1 _2686_ (.Y(_0970_),
    .B(\cic_b.delay[0][11] ),
    .A_N(\cic_b.integrator[2][11] ));
 sg13g2_nand2b_1 _2687_ (.Y(_0971_),
    .B(_0970_),
    .A_N(_0969_));
 sg13g2_a21oi_1 _2688_ (.A1(_0964_),
    .A2(_0967_),
    .Y(_0972_),
    .B1(_0965_));
 sg13g2_xnor2_1 _2689_ (.Y(_0973_),
    .A(_0971_),
    .B(_0972_));
 sg13g2_nor2_1 _2690_ (.A(net218),
    .B(net473),
    .Y(_0974_));
 sg13g2_a21oi_1 _2691_ (.A1(net471),
    .A2(_0973_),
    .Y(_0284_),
    .B1(_0974_));
 sg13g2_nor2_1 _2692_ (.A(net347),
    .B(net472),
    .Y(_0975_));
 sg13g2_nor3_1 _2693_ (.A(_0965_),
    .B(_0966_),
    .C(_0971_),
    .Y(_0976_));
 sg13g2_a221oi_1 _2694_ (.B2(_0964_),
    .C1(_0969_),
    .B1(_0976_),
    .A1(_0965_),
    .Y(_0977_),
    .A2(_0970_));
 sg13g2_xor2_1 _2695_ (.B(net632),
    .A(net353),
    .X(_0978_));
 sg13g2_xnor2_1 _2696_ (.Y(_0979_),
    .A(_0977_),
    .B(_0978_));
 sg13g2_a21oi_1 _2697_ (.A1(net472),
    .A2(_0979_),
    .Y(_0285_),
    .B1(_0975_));
 sg13g2_mux2_1 _2698_ (.A0(net348),
    .A1(net339),
    .S(net497),
    .X(_0286_));
 sg13g2_mux2_1 _2699_ (.A0(net456),
    .A1(net169),
    .S(net497),
    .X(_0287_));
 sg13g2_mux2_1 _2700_ (.A0(net150),
    .A1(net346),
    .S(net499),
    .X(_0288_));
 sg13g2_mux2_1 _2701_ (.A0(net440),
    .A1(net123),
    .S(net498),
    .X(_0289_));
 sg13g2_mux2_1 _2702_ (.A0(net417),
    .A1(net174),
    .S(net488),
    .X(_0290_));
 sg13g2_nand2_1 _2703_ (.Y(_0980_),
    .A(net25),
    .B(net488));
 sg13g2_o21ai_1 _2704_ (.B1(_0980_),
    .Y(_0291_),
    .A1(_1202_),
    .A2(net488));
 sg13g2_mux2_1 _2705_ (.A0(net449),
    .A1(net130),
    .S(net488),
    .X(_0292_));
 sg13g2_mux2_1 _2706_ (.A0(net381),
    .A1(net176),
    .S(net488),
    .X(_0293_));
 sg13g2_mux2_1 _2707_ (.A0(net448),
    .A1(net112),
    .S(net489),
    .X(_0294_));
 sg13g2_mux2_1 _2708_ (.A0(net446),
    .A1(net194),
    .S(net478),
    .X(_0295_));
 sg13g2_mux2_1 _2709_ (.A0(net285),
    .A1(net433),
    .S(net478),
    .X(_0296_));
 sg13g2_mux2_1 _2710_ (.A0(net447),
    .A1(net392),
    .S(net489),
    .X(_0297_));
 sg13g2_mux2_1 _2711_ (.A0(net443),
    .A1(net264),
    .S(net498),
    .X(_0298_));
 sg13g2_nor2_1 _2712_ (.A(net339),
    .B(net497),
    .Y(_0981_));
 sg13g2_nand2b_1 _2713_ (.Y(_0982_),
    .B(\cic_b.delay[2][0] ),
    .A_N(\cic_b.temp_comb[1][0] ));
 sg13g2_xnor2_1 _2714_ (.Y(_0983_),
    .A(\cic_b.temp_comb[1][0] ),
    .B(net216));
 sg13g2_a21oi_1 _2715_ (.A1(net497),
    .A2(_0983_),
    .Y(_0299_),
    .B1(_0981_));
 sg13g2_nor2_1 _2716_ (.A(net169),
    .B(net497),
    .Y(_0984_));
 sg13g2_nor2b_1 _2717_ (.A(\cic_b.delay[2][1] ),
    .B_N(\cic_b.temp_comb[1][1] ),
    .Y(_0985_));
 sg13g2_xnor2_1 _2718_ (.Y(_0986_),
    .A(\cic_b.temp_comb[1][1] ),
    .B(\cic_b.delay[2][1] ));
 sg13g2_xnor2_1 _2719_ (.Y(_0987_),
    .A(_0982_),
    .B(_0986_));
 sg13g2_a21oi_1 _2720_ (.A1(net497),
    .A2(_0987_),
    .Y(_0300_),
    .B1(_0984_));
 sg13g2_nor2b_1 _2721_ (.A(\cic_b.delay[2][2] ),
    .B_N(\cic_b.temp_comb[1][2] ),
    .Y(_0988_));
 sg13g2_nand2b_1 _2722_ (.Y(_0989_),
    .B(\cic_b.delay[2][2] ),
    .A_N(\cic_b.temp_comb[1][2] ));
 sg13g2_nor2b_1 _2723_ (.A(_0988_),
    .B_N(_0989_),
    .Y(_0990_));
 sg13g2_a21o_1 _2724_ (.A2(_0986_),
    .A1(_0982_),
    .B1(_0985_),
    .X(_0991_));
 sg13g2_xnor2_1 _2725_ (.Y(_0992_),
    .A(_0990_),
    .B(_0991_));
 sg13g2_nor2_1 _2726_ (.A(net346),
    .B(net498),
    .Y(_0993_));
 sg13g2_a21oi_1 _2727_ (.A1(net495),
    .A2(_0992_),
    .Y(_0301_),
    .B1(_0993_));
 sg13g2_nor2_1 _2728_ (.A(net123),
    .B(net498),
    .Y(_0994_));
 sg13g2_nand2b_1 _2729_ (.Y(_0995_),
    .B(\cic_b.temp_comb[1][3] ),
    .A_N(\cic_b.delay[2][3] ));
 sg13g2_xor2_1 _2730_ (.B(\cic_b.delay[2][3] ),
    .A(\cic_b.temp_comb[1][3] ),
    .X(_0996_));
 sg13g2_a21oi_1 _2731_ (.A1(_0989_),
    .A2(_0991_),
    .Y(_0997_),
    .B1(_0988_));
 sg13g2_xnor2_1 _2732_ (.Y(_0998_),
    .A(_0996_),
    .B(_0997_));
 sg13g2_a21oi_1 _2733_ (.A1(net498),
    .A2(_0998_),
    .Y(_0302_),
    .B1(_0994_));
 sg13g2_nor2_1 _2734_ (.A(net174),
    .B(net488),
    .Y(_0999_));
 sg13g2_o21ai_1 _2735_ (.B1(_0995_),
    .Y(_1000_),
    .A1(_0996_),
    .A2(_0997_));
 sg13g2_nor2b_1 _2736_ (.A(\cic_b.delay[2][4] ),
    .B_N(\cic_b.temp_comb[1][4] ),
    .Y(_1001_));
 sg13g2_xnor2_1 _2737_ (.Y(_1002_),
    .A(\cic_b.temp_comb[1][4] ),
    .B(\cic_b.delay[2][4] ));
 sg13g2_inv_1 _2738_ (.Y(_1003_),
    .A(_1002_));
 sg13g2_xnor2_1 _2739_ (.Y(_1004_),
    .A(_1000_),
    .B(_1002_));
 sg13g2_a21oi_1 _2740_ (.A1(net487),
    .A2(_1004_),
    .Y(_0303_),
    .B1(_0999_));
 sg13g2_nand2b_1 _2741_ (.Y(_1005_),
    .B(\cic_b.delay[2][5] ),
    .A_N(\cic_b.temp_comb[1][5] ));
 sg13g2_nor2b_1 _2742_ (.A(\cic_b.delay[2][5] ),
    .B_N(\cic_b.temp_comb[1][5] ),
    .Y(_1006_));
 sg13g2_xor2_1 _2743_ (.B(\cic_b.delay[2][5] ),
    .A(\cic_b.temp_comb[1][5] ),
    .X(_1007_));
 sg13g2_a21oi_1 _2744_ (.A1(_1000_),
    .A2(_1002_),
    .Y(_1008_),
    .B1(_1001_));
 sg13g2_xor2_1 _2745_ (.B(_1008_),
    .A(_1007_),
    .X(_1009_));
 sg13g2_mux2_1 _2746_ (.A0(net25),
    .A1(_1009_),
    .S(net487),
    .X(_0304_));
 sg13g2_nor2_1 _2747_ (.A(net130),
    .B(net490),
    .Y(_1010_));
 sg13g2_nand2b_1 _2748_ (.Y(_1011_),
    .B(\cic_b.temp_comb[1][6] ),
    .A_N(\cic_b.delay[2][6] ));
 sg13g2_xor2_1 _2749_ (.B(\cic_b.delay[2][6] ),
    .A(\cic_b.temp_comb[1][6] ),
    .X(_1012_));
 sg13g2_nor2_1 _2750_ (.A(_1003_),
    .B(_1007_),
    .Y(_1013_));
 sg13g2_a21o_1 _2751_ (.A2(_1005_),
    .A1(_1001_),
    .B1(_1006_),
    .X(_1014_));
 sg13g2_a21oi_1 _2752_ (.A1(_1000_),
    .A2(_1013_),
    .Y(_1015_),
    .B1(_1014_));
 sg13g2_xnor2_1 _2753_ (.Y(_1016_),
    .A(_1012_),
    .B(_1015_));
 sg13g2_a21oi_1 _2754_ (.A1(net487),
    .A2(_1016_),
    .Y(_0305_),
    .B1(_1010_));
 sg13g2_nor2b_1 _2755_ (.A(\cic_b.temp_comb[1][7] ),
    .B_N(\cic_b.delay[2][7] ),
    .Y(_1017_));
 sg13g2_nand2b_1 _2756_ (.Y(_1018_),
    .B(\cic_b.temp_comb[1][7] ),
    .A_N(\cic_b.delay[2][7] ));
 sg13g2_nand2b_1 _2757_ (.Y(_1019_),
    .B(_1018_),
    .A_N(_1017_));
 sg13g2_o21ai_1 _2758_ (.B1(_1011_),
    .Y(_1020_),
    .A1(_1012_),
    .A2(_1015_));
 sg13g2_xnor2_1 _2759_ (.Y(_1021_),
    .A(_1019_),
    .B(_1020_));
 sg13g2_mux2_1 _2760_ (.A0(net176),
    .A1(_1021_),
    .S(net489),
    .X(_0306_));
 sg13g2_nor2_1 _2761_ (.A(_1012_),
    .B(_1019_),
    .Y(_1022_));
 sg13g2_and2_1 _2762_ (.A(_1013_),
    .B(_1022_),
    .X(_1023_));
 sg13g2_o21ai_1 _2763_ (.B1(_1018_),
    .Y(_1024_),
    .A1(_1011_),
    .A2(_1017_));
 sg13g2_a221oi_1 _2764_ (.B2(_1000_),
    .C1(_1024_),
    .B1(_1023_),
    .A1(_1014_),
    .Y(_1025_),
    .A2(_1022_));
 sg13g2_nand2b_1 _2765_ (.Y(_1026_),
    .B(\cic_b.temp_comb[1][8] ),
    .A_N(\cic_b.delay[2][8] ));
 sg13g2_xor2_1 _2766_ (.B(\cic_b.delay[2][8] ),
    .A(\cic_b.temp_comb[1][8] ),
    .X(_1027_));
 sg13g2_xnor2_1 _2767_ (.Y(_1028_),
    .A(_1025_),
    .B(_1027_));
 sg13g2_nor2_1 _2768_ (.A(net112),
    .B(net478),
    .Y(_1029_));
 sg13g2_a21oi_1 _2769_ (.A1(net478),
    .A2(_1028_),
    .Y(_0307_),
    .B1(_1029_));
 sg13g2_nor2_1 _2770_ (.A(net194),
    .B(net478),
    .Y(_1030_));
 sg13g2_xnor2_1 _2771_ (.Y(_1031_),
    .A(\cic_b.temp_comb[1][9] ),
    .B(\cic_b.delay[2][9] ));
 sg13g2_o21ai_1 _2772_ (.B1(_1026_),
    .Y(_1032_),
    .A1(_1025_),
    .A2(_1027_));
 sg13g2_xnor2_1 _2773_ (.Y(_1033_),
    .A(_1031_),
    .B(_1032_));
 sg13g2_a21oi_1 _2774_ (.A1(net479),
    .A2(_1033_),
    .Y(_0308_),
    .B1(_1030_));
 sg13g2_nor2_1 _2775_ (.A(net433),
    .B(net478),
    .Y(_1034_));
 sg13g2_nand2b_1 _2776_ (.Y(_1035_),
    .B(_1031_),
    .A_N(_1027_));
 sg13g2_a21oi_1 _2777_ (.A1(_1227_),
    .A2(\cic_b.delay[2][9] ),
    .Y(_1036_),
    .B1(_1026_));
 sg13g2_a21oi_1 _2778_ (.A1(\cic_b.temp_comb[1][9] ),
    .A2(_1228_),
    .Y(_1037_),
    .B1(_1036_));
 sg13g2_o21ai_1 _2779_ (.B1(_1037_),
    .Y(_1038_),
    .A1(_1025_),
    .A2(_1035_));
 sg13g2_nor2b_1 _2780_ (.A(\cic_b.delay[2][10] ),
    .B_N(\cic_b.temp_comb[1][10] ),
    .Y(_1039_));
 sg13g2_nor2b_1 _2781_ (.A(\cic_b.temp_comb[1][10] ),
    .B_N(\cic_b.delay[2][10] ),
    .Y(_1040_));
 sg13g2_nor2_1 _2782_ (.A(_1039_),
    .B(_1040_),
    .Y(_1041_));
 sg13g2_xnor2_1 _2783_ (.Y(_1042_),
    .A(_1038_),
    .B(_1041_));
 sg13g2_a21oi_1 _2784_ (.A1(net478),
    .A2(_1042_),
    .Y(_0309_),
    .B1(_1034_));
 sg13g2_nor2b_1 _2785_ (.A(\cic_b.delay[2][11] ),
    .B_N(\cic_b.temp_comb[1][11] ),
    .Y(_1043_));
 sg13g2_nand2b_1 _2786_ (.Y(_1044_),
    .B(\cic_b.delay[2][11] ),
    .A_N(\cic_b.temp_comb[1][11] ));
 sg13g2_nand2b_1 _2787_ (.Y(_1045_),
    .B(_1044_),
    .A_N(_1043_));
 sg13g2_a21oi_1 _2788_ (.A1(_1038_),
    .A2(_1041_),
    .Y(_1046_),
    .B1(_1039_));
 sg13g2_xnor2_1 _2789_ (.Y(_1047_),
    .A(_1045_),
    .B(_1046_));
 sg13g2_nor2_1 _2790_ (.A(net392),
    .B(net489),
    .Y(_1048_));
 sg13g2_a21oi_1 _2791_ (.A1(net489),
    .A2(_1047_),
    .Y(_0310_),
    .B1(_1048_));
 sg13g2_nor2_1 _2792_ (.A(net264),
    .B(net490),
    .Y(_1049_));
 sg13g2_nor3_1 _2793_ (.A(_1039_),
    .B(_1040_),
    .C(_1045_),
    .Y(_1050_));
 sg13g2_a221oi_1 _2794_ (.B2(_1038_),
    .C1(_1043_),
    .B1(_1050_),
    .A1(_1039_),
    .Y(_1051_),
    .A2(_1044_));
 sg13g2_xor2_1 _2795_ (.B(\cic_b.delay[2][12] ),
    .A(\cic_b.temp_comb[1][12] ),
    .X(_1052_));
 sg13g2_xnor2_1 _2796_ (.Y(_1053_),
    .A(_1051_),
    .B(_1052_));
 sg13g2_a21oi_1 _2797_ (.A1(net487),
    .A2(_1053_),
    .Y(_0311_),
    .B1(_1049_));
 sg13g2_mux2_1 _2798_ (.A0(net299),
    .A1(\cic_b.integrator[2][0] ),
    .S(net493),
    .X(_0312_));
 sg13g2_mux2_1 _2799_ (.A0(net199),
    .A1(net352),
    .S(net493),
    .X(_0313_));
 sg13g2_mux2_1 _2800_ (.A0(net239),
    .A1(\cic_b.integrator[2][2] ),
    .S(net493),
    .X(_0314_));
 sg13g2_mux2_1 _2801_ (.A0(net297),
    .A1(\cic_b.integrator[2][3] ),
    .S(net494),
    .X(_0315_));
 sg13g2_mux2_1 _2802_ (.A0(net385),
    .A1(\cic_b.integrator[2][4] ),
    .S(net485),
    .X(_0316_));
 sg13g2_nor2_1 _2803_ (.A(net43),
    .B(net485),
    .Y(_1054_));
 sg13g2_a21oi_1 _2804_ (.A1(_1223_),
    .A2(net485),
    .Y(_0317_),
    .B1(_1054_));
 sg13g2_mux2_1 _2805_ (.A0(net223),
    .A1(\cic_b.integrator[2][6] ),
    .S(net483),
    .X(_0318_));
 sg13g2_mux2_1 _2806_ (.A0(net301),
    .A1(\cic_b.integrator[2][7] ),
    .S(net476),
    .X(_0319_));
 sg13g2_mux2_1 _2807_ (.A0(net229),
    .A1(\cic_b.integrator[2][8] ),
    .S(net475),
    .X(_0320_));
 sg13g2_nor2_1 _2808_ (.A(net58),
    .B(net475),
    .Y(_1055_));
 sg13g2_a21oi_1 _2809_ (.A1(_1225_),
    .A2(net475),
    .Y(_0321_),
    .B1(_1055_));
 sg13g2_mux2_1 _2810_ (.A0(net235),
    .A1(\cic_b.integrator[2][10] ),
    .S(net471),
    .X(_0322_));
 sg13g2_mux2_1 _2811_ (.A0(net20),
    .A1(net127),
    .S(net471),
    .X(_0323_));
 sg13g2_mux2_1 _2812_ (.A0(net186),
    .A1(net353),
    .S(net472),
    .X(_0324_));
 sg13g2_mux2_1 _2813_ (.A0(net159),
    .A1(\cic_a.temp_comb[1][0] ),
    .S(net525),
    .X(_0325_));
 sg13g2_mux2_1 _2814_ (.A0(net153),
    .A1(\cic_a.temp_comb[1][1] ),
    .S(net523),
    .X(_0326_));
 sg13g2_mux2_1 _2815_ (.A0(net121),
    .A1(\cic_a.temp_comb[1][2] ),
    .S(net521),
    .X(_0327_));
 sg13g2_mux2_1 _2816_ (.A0(net212),
    .A1(\cic_a.temp_comb[1][3] ),
    .S(net519),
    .X(_0328_));
 sg13g2_mux2_1 _2817_ (.A0(net163),
    .A1(\cic_a.temp_comb[1][4] ),
    .S(net515),
    .X(_0329_));
 sg13g2_mux2_1 _2818_ (.A0(net397),
    .A1(net409),
    .S(net514),
    .X(_0330_));
 sg13g2_mux2_1 _2819_ (.A0(net395),
    .A1(\cic_a.temp_comb[1][6] ),
    .S(net514),
    .X(_0331_));
 sg13g2_mux2_1 _2820_ (.A0(net262),
    .A1(\cic_a.temp_comb[1][7] ),
    .S(net514),
    .X(_0332_));
 sg13g2_mux2_1 _2821_ (.A0(net71),
    .A1(net338),
    .S(net512),
    .X(_0333_));
 sg13g2_mux2_1 _2822_ (.A0(net289),
    .A1(\cic_a.temp_comb[1][9] ),
    .S(net507),
    .X(_0334_));
 sg13g2_mux2_1 _2823_ (.A0(net246),
    .A1(net284),
    .S(net512),
    .X(_0335_));
 sg13g2_mux2_1 _2824_ (.A0(net287),
    .A1(\cic_a.temp_comb[1][11] ),
    .S(net512),
    .X(_0336_));
 sg13g2_mux2_1 _2825_ (.A0(net221),
    .A1(\cic_a.temp_comb[1][12] ),
    .S(net504),
    .X(_0337_));
 sg13g2_mux2_1 _2826_ (.A0(net205),
    .A1(\cic_b.temp_comb[0][0] ),
    .S(net492),
    .X(_0338_));
 sg13g2_mux2_1 _2827_ (.A0(net336),
    .A1(\cic_b.temp_comb[0][1] ),
    .S(net491),
    .X(_0339_));
 sg13g2_mux2_1 _2828_ (.A0(net182),
    .A1(\cic_b.temp_comb[0][2] ),
    .S(net491),
    .X(_0340_));
 sg13g2_mux2_1 _2829_ (.A0(net268),
    .A1(\cic_b.temp_comb[0][3] ),
    .S(net494),
    .X(_0341_));
 sg13g2_mux2_1 _2830_ (.A0(net27),
    .A1(net143),
    .S(net484),
    .X(_0342_));
 sg13g2_mux2_1 _2831_ (.A0(net304),
    .A1(\cic_b.temp_comb[0][5] ),
    .S(net484),
    .X(_0343_));
 sg13g2_mux2_1 _2832_ (.A0(net330),
    .A1(\cic_b.temp_comb[0][6] ),
    .S(net482),
    .X(_0344_));
 sg13g2_mux2_1 _2833_ (.A0(net233),
    .A1(\cic_b.temp_comb[0][7] ),
    .S(net476),
    .X(_0345_));
 sg13g2_mux2_1 _2834_ (.A0(net179),
    .A1(\cic_b.temp_comb[0][8] ),
    .S(net476),
    .X(_0346_));
 sg13g2_nor2_1 _2835_ (.A(net89),
    .B(net474),
    .Y(_1056_));
 sg13g2_a21oi_1 _2836_ (.A1(_1230_),
    .A2(net474),
    .Y(_0347_),
    .B1(_1056_));
 sg13g2_mux2_1 _2837_ (.A0(net279),
    .A1(net283),
    .S(net474),
    .X(_0348_));
 sg13g2_mux2_1 _2838_ (.A0(net146),
    .A1(net218),
    .S(net473),
    .X(_0349_));
 sg13g2_mux2_1 _2839_ (.A0(net148),
    .A1(net347),
    .S(net472),
    .X(_0350_));
 sg13g2_a22oi_1 _2840_ (.Y(_1057_),
    .B1(_0586_),
    .B2(net35),
    .A2(net539),
    .A1(\cic_a.filtered_out[0] ));
 sg13g2_inv_1 _2841_ (.Y(_0351_),
    .A(net36));
 sg13g2_a22oi_1 _2842_ (.Y(_1058_),
    .B1(net360),
    .B2(net539),
    .A2(net35),
    .A1(net547));
 sg13g2_o21ai_1 _2843_ (.B1(net361),
    .Y(_0352_),
    .A1(_1192_),
    .A2(net531));
 sg13g2_a22oi_1 _2844_ (.Y(_1059_),
    .B1(\cic_a.filtered_out[2] ),
    .B2(net538),
    .A2(net117),
    .A1(net546));
 sg13g2_o21ai_1 _2845_ (.B1(net118),
    .Y(_0353_),
    .A1(_1193_),
    .A2(net531));
 sg13g2_nand2_1 _2846_ (.Y(_1060_),
    .A(net547),
    .B(net86));
 sg13g2_a22oi_1 _2847_ (.Y(_1061_),
    .B1(_0586_),
    .B2(\serializer_a.shift_reg[3] ),
    .A2(net538),
    .A1(\cic_a.filtered_out[3] ));
 sg13g2_nand2_1 _2848_ (.Y(_0354_),
    .A(net87),
    .B(_1061_));
 sg13g2_a22oi_1 _2849_ (.Y(_1062_),
    .B1(\cic_a.filtered_out[4] ),
    .B2(net538),
    .A2(net172),
    .A1(net545));
 sg13g2_o21ai_1 _2850_ (.B1(net173),
    .Y(_0355_),
    .A1(_1194_),
    .A2(net530));
 sg13g2_nand2_1 _2851_ (.Y(_1063_),
    .A(net545),
    .B(net45));
 sg13g2_a22oi_1 _2852_ (.Y(_1064_),
    .B1(_0586_),
    .B2(\serializer_a.shift_reg[5] ),
    .A2(net538),
    .A1(\cic_a.filtered_out[5] ));
 sg13g2_nand2_1 _2853_ (.Y(_0356_),
    .A(net46),
    .B(_1064_));
 sg13g2_a22oi_1 _2854_ (.Y(_1065_),
    .B1(\cic_a.filtered_out[6] ),
    .B2(net538),
    .A2(net374),
    .A1(net545));
 sg13g2_o21ai_1 _2855_ (.B1(net375),
    .Y(_0357_),
    .A1(_1195_),
    .A2(net530));
 sg13g2_a22oi_1 _2856_ (.Y(_1066_),
    .B1(\cic_a.filtered_out[7] ),
    .B2(net538),
    .A2(net356),
    .A1(net545));
 sg13g2_o21ai_1 _2857_ (.B1(net357),
    .Y(_0358_),
    .A1(_1197_),
    .A2(net530));
 sg13g2_nand2_1 _2858_ (.Y(_1067_),
    .A(net545),
    .B(net209));
 sg13g2_a22oi_1 _2859_ (.Y(_1068_),
    .B1(_0586_),
    .B2(\serializer_a.shift_reg[8] ),
    .A2(net538),
    .A1(\cic_a.filtered_out[8] ));
 sg13g2_nand2_1 _2860_ (.Y(_0359_),
    .A(net210),
    .B(_1068_));
 sg13g2_a22oi_1 _2861_ (.Y(_1069_),
    .B1(\cic_a.filtered_out[9] ),
    .B2(net538),
    .A2(\serializer_a.shift_reg[8] ),
    .A1(net545));
 sg13g2_o21ai_1 _2862_ (.B1(_1069_),
    .Y(_0360_),
    .A1(_1198_),
    .A2(net530));
 sg13g2_a22oi_1 _2863_ (.Y(_1070_),
    .B1(\cic_a.filtered_out[10] ),
    .B2(net539),
    .A2(\serializer_a.shift_reg[9] ),
    .A1(net545));
 sg13g2_o21ai_1 _2864_ (.B1(_1070_),
    .Y(_0361_),
    .A1(_1199_),
    .A2(net530));
 sg13g2_a22oi_1 _2865_ (.Y(_1071_),
    .B1(\cic_a.filtered_out[11] ),
    .B2(net539),
    .A2(net203),
    .A1(net545));
 sg13g2_o21ai_1 _2866_ (.B1(_1071_),
    .Y(_0362_),
    .A1(_1200_),
    .A2(net530));
 sg13g2_a22oi_1 _2867_ (.Y(_1072_),
    .B1(\cic_a.filtered_out[12] ),
    .B2(net539),
    .A2(\serializer_a.shift_reg[11] ),
    .A1(net546));
 sg13g2_o21ai_1 _2868_ (.B1(_1072_),
    .Y(_0363_),
    .A1(_1233_),
    .A2(net530));
 sg13g2_mux2_1 _2869_ (.A0(net201),
    .A1(\cic_b.temp_comb[1][0] ),
    .S(net496),
    .X(_0364_));
 sg13g2_mux2_1 _2870_ (.A0(net319),
    .A1(\cic_b.temp_comb[1][1] ),
    .S(net495),
    .X(_0365_));
 sg13g2_mux2_1 _2871_ (.A0(net219),
    .A1(\cic_b.temp_comb[1][2] ),
    .S(net495),
    .X(_0366_));
 sg13g2_mux2_1 _2872_ (.A0(net248),
    .A1(\cic_b.temp_comb[1][3] ),
    .S(net498),
    .X(_0367_));
 sg13g2_mux2_1 _2873_ (.A0(net272),
    .A1(\cic_b.temp_comb[1][4] ),
    .S(net487),
    .X(_0368_));
 sg13g2_mux2_1 _2874_ (.A0(net266),
    .A1(\cic_b.temp_comb[1][5] ),
    .S(net487),
    .X(_0369_));
 sg13g2_mux2_1 _2875_ (.A0(net256),
    .A1(\cic_b.temp_comb[1][6] ),
    .S(net482),
    .X(_0370_));
 sg13g2_mux2_1 _2876_ (.A0(net366),
    .A1(\cic_b.temp_comb[1][7] ),
    .S(net482),
    .X(_0371_));
 sg13g2_mux2_1 _2877_ (.A0(net322),
    .A1(\cic_b.temp_comb[1][8] ),
    .S(net477),
    .X(_0372_));
 sg13g2_nor2_1 _2878_ (.A(net37),
    .B(net478),
    .Y(_1073_));
 sg13g2_a21oi_1 _2879_ (.A1(_1227_),
    .A2(net477),
    .Y(_0373_),
    .B1(_1073_));
 sg13g2_mux2_1 _2880_ (.A0(net241),
    .A1(\cic_b.temp_comb[1][10] ),
    .S(net480),
    .X(_0374_));
 sg13g2_mux2_1 _2881_ (.A0(net316),
    .A1(net318),
    .S(net480),
    .X(_0375_));
 sg13g2_mux2_1 _2882_ (.A0(net342),
    .A1(\cic_b.temp_comb[1][12] ),
    .S(net473),
    .X(_0376_));
 sg13g2_a22oi_1 _2883_ (.Y(_1074_),
    .B1(_0590_),
    .B2(net33),
    .A2(net535),
    .A1(\cic_b.filtered_out[0] ));
 sg13g2_inv_1 _2884_ (.Y(_0377_),
    .A(net34));
 sg13g2_nand2_1 _2885_ (.Y(_1075_),
    .A(net543),
    .B(net33));
 sg13g2_a22oi_1 _2886_ (.Y(_1076_),
    .B1(_0590_),
    .B2(net73),
    .A2(net535),
    .A1(\cic_b.filtered_out[1] ));
 sg13g2_nand2_1 _2887_ (.Y(_0378_),
    .A(_1075_),
    .B(net74));
 sg13g2_a22oi_1 _2888_ (.Y(_1077_),
    .B1(net150),
    .B2(net535),
    .A2(net73),
    .A1(net704));
 sg13g2_o21ai_1 _2889_ (.B1(_1077_),
    .Y(_0379_),
    .A1(_1201_),
    .A2(net529));
 sg13g2_nand2_1 _2890_ (.Y(_1078_),
    .A(net543),
    .B(net83));
 sg13g2_a22oi_1 _2891_ (.Y(_1079_),
    .B1(_0590_),
    .B2(net78),
    .A2(net535),
    .A1(\cic_b.filtered_out[3] ));
 sg13g2_nand2_1 _2892_ (.Y(_0380_),
    .A(net84),
    .B(_1079_));
 sg13g2_nand2_1 _2893_ (.Y(_1080_),
    .A(net544),
    .B(net78));
 sg13g2_a22oi_1 _2894_ (.Y(_1081_),
    .B1(_0590_),
    .B2(net65),
    .A2(net534),
    .A1(\cic_b.filtered_out[4] ));
 sg13g2_nand2_1 _2895_ (.Y(_0381_),
    .A(net79),
    .B(_1081_));
 sg13g2_nand2_1 _2896_ (.Y(_1082_),
    .A(net544),
    .B(net65));
 sg13g2_a22oi_1 _2897_ (.Y(_1083_),
    .B1(_0590_),
    .B2(\serializer_b.shift_reg[5] ),
    .A2(net534),
    .A1(\cic_b.filtered_out[5] ));
 sg13g2_nand2_1 _2898_ (.Y(_0382_),
    .A(net66),
    .B(_1083_));
 sg13g2_a22oi_1 _2899_ (.Y(_1084_),
    .B1(\cic_b.filtered_out[6] ),
    .B2(net534),
    .A2(\serializer_b.shift_reg[5] ),
    .A1(net544));
 sg13g2_o21ai_1 _2900_ (.B1(_1084_),
    .Y(_0383_),
    .A1(_1203_),
    .A2(net529));
 sg13g2_a22oi_1 _2901_ (.Y(_1085_),
    .B1(\cic_b.filtered_out[7] ),
    .B2(net534),
    .A2(net258),
    .A1(net544));
 sg13g2_o21ai_1 _2902_ (.B1(_1085_),
    .Y(_0384_),
    .A1(_1204_),
    .A2(net529));
 sg13g2_a22oi_1 _2903_ (.Y(_1086_),
    .B1(\cic_b.filtered_out[8] ),
    .B2(net534),
    .A2(\serializer_b.shift_reg[7] ),
    .A1(net544));
 sg13g2_o21ai_1 _2904_ (.B1(_1086_),
    .Y(_0385_),
    .A1(_1205_),
    .A2(net529));
 sg13g2_a22oi_1 _2905_ (.Y(_1087_),
    .B1(\cic_b.filtered_out[9] ),
    .B2(net534),
    .A2(net135),
    .A1(net544));
 sg13g2_o21ai_1 _2906_ (.B1(_1087_),
    .Y(_0386_),
    .A1(_1206_),
    .A2(net529));
 sg13g2_a22oi_1 _2907_ (.Y(_1088_),
    .B1(net285),
    .B2(net534),
    .A2(net177),
    .A1(net544));
 sg13g2_o21ai_1 _2908_ (.B1(net286),
    .Y(_0387_),
    .A1(_1207_),
    .A2(net529));
 sg13g2_a22oi_1 _2909_ (.Y(_1089_),
    .B1(\cic_b.filtered_out[11] ),
    .B2(net534),
    .A2(net133),
    .A1(net544));
 sg13g2_o21ai_1 _2910_ (.B1(net134),
    .Y(_0388_),
    .A1(_1208_),
    .A2(_0591_));
 sg13g2_nand2_1 _2911_ (.Y(_1090_),
    .A(\serializer_b.sending ),
    .B(net103));
 sg13g2_a22oi_1 _2912_ (.Y(_1091_),
    .B1(_0590_),
    .B2(\serializer_b.serial_out ),
    .A2(net535),
    .A1(\cic_b.filtered_out[12] ));
 sg13g2_nand2_1 _2913_ (.Y(_0389_),
    .A(net104),
    .B(_1091_));
 sg13g2_nor2_1 _2914_ (.A(net540),
    .B(net91),
    .Y(_1092_));
 sg13g2_a21oi_1 _2915_ (.A1(net91),
    .A2(_0595_),
    .Y(_0390_),
    .B1(_1092_));
 sg13g2_nand2_1 _2916_ (.Y(_1093_),
    .A(net106),
    .B(net533));
 sg13g2_and2_1 _2917_ (.A(net91),
    .B(net106),
    .X(_1094_));
 sg13g2_o21ai_1 _2918_ (.B1(_1093_),
    .Y(_0391_),
    .A1(_0596_),
    .A2(_1094_));
 sg13g2_nand3_1 _2919_ (.B(net96),
    .C(_1094_),
    .A(net540),
    .Y(_1095_));
 sg13g2_nand2_1 _2920_ (.Y(_1096_),
    .A(net536),
    .B(_1095_));
 sg13g2_a21oi_1 _2921_ (.A1(_0595_),
    .A2(_1094_),
    .Y(_1097_),
    .B1(net96));
 sg13g2_nor2_1 _2922_ (.A(_1096_),
    .B(net97),
    .Y(_0392_));
 sg13g2_nor2b_1 _2923_ (.A(net81),
    .B_N(_1095_),
    .Y(_1098_));
 sg13g2_a21oi_1 _2924_ (.A1(net81),
    .A2(_1096_),
    .Y(_0393_),
    .B1(_1098_));
 sg13g2_nor2_1 _2925_ (.A(net543),
    .B(net108),
    .Y(_1099_));
 sg13g2_a21oi_1 _2926_ (.A1(net108),
    .A2(net529),
    .Y(_0394_),
    .B1(_1099_));
 sg13g2_nand2_1 _2927_ (.Y(_1100_),
    .A(net232),
    .B(_0590_));
 sg13g2_and2_1 _2928_ (.A(net108),
    .B(net232),
    .X(_1101_));
 sg13g2_o21ai_1 _2929_ (.B1(_1100_),
    .Y(_0395_),
    .A1(_0592_),
    .A2(_1101_));
 sg13g2_nand3_1 _2930_ (.B(net76),
    .C(_1101_),
    .A(net543),
    .Y(_1102_));
 sg13g2_nand2b_1 _2931_ (.Y(_1103_),
    .B(_1102_),
    .A_N(net535));
 sg13g2_a21oi_1 _2932_ (.A1(net529),
    .A2(_1101_),
    .Y(_1104_),
    .B1(net76));
 sg13g2_nor2_1 _2933_ (.A(_1103_),
    .B(net77),
    .Y(_0396_));
 sg13g2_nor2b_1 _2934_ (.A(net63),
    .B_N(_1102_),
    .Y(_1105_));
 sg13g2_a21oi_1 _2935_ (.A1(net63),
    .A2(_1103_),
    .Y(_0397_),
    .B1(_1105_));
 sg13g2_nand2b_2 _2936_ (.Y(_1106_),
    .B(net348),
    .A_N(\cic_a.filtered_out[0] ));
 sg13g2_nand2b_1 _2937_ (.Y(_1107_),
    .B(\cic_a.filtered_out[0] ),
    .A_N(\cic_b.filtered_out[0] ));
 sg13g2_a21o_1 _2938_ (.A2(_1107_),
    .A1(_1106_),
    .B1(net536),
    .X(_1108_));
 sg13g2_o21ai_1 _2939_ (.B1(_1108_),
    .Y(_0398_),
    .A1(_1209_),
    .A2(_0595_));
 sg13g2_nor2b_1 _2940_ (.A(\cic_b.filtered_out[1] ),
    .B_N(\cic_a.filtered_out[1] ),
    .Y(_1109_));
 sg13g2_xnor2_1 _2941_ (.Y(_1110_),
    .A(\cic_a.filtered_out[1] ),
    .B(\cic_b.filtered_out[1] ));
 sg13g2_xnor2_1 _2942_ (.Y(_1111_),
    .A(_1106_),
    .B(_1110_));
 sg13g2_nor2_1 _2943_ (.A(net214),
    .B(_0595_),
    .Y(_1112_));
 sg13g2_a221oi_1 _2944_ (.B2(_1111_),
    .C1(_1112_),
    .B1(_0019_),
    .A1(net540),
    .Y(_0399_),
    .A2(_1209_));
 sg13g2_a21oi_2 _2945_ (.B1(_1109_),
    .Y(_1113_),
    .A2(_1110_),
    .A1(_1106_));
 sg13g2_nor2b_1 _2946_ (.A(\cic_b.filtered_out[2] ),
    .B_N(\cic_a.filtered_out[2] ),
    .Y(_1114_));
 sg13g2_xor2_1 _2947_ (.B(\cic_b.filtered_out[2] ),
    .A(\cic_a.filtered_out[2] ),
    .X(_1115_));
 sg13g2_nor2_1 _2948_ (.A(_1113_),
    .B(_1115_),
    .Y(_1116_));
 sg13g2_a21o_1 _2949_ (.A2(_1115_),
    .A1(_1113_),
    .B1(net537),
    .X(_1117_));
 sg13g2_a22oi_1 _2950_ (.Y(_1118_),
    .B1(net418),
    .B2(net533),
    .A2(net214),
    .A1(net542));
 sg13g2_o21ai_1 _2951_ (.B1(net419),
    .Y(_0400_),
    .A1(_1116_),
    .A2(_1117_));
 sg13g2_nor2b_1 _2952_ (.A(\cic_b.filtered_out[3] ),
    .B_N(\cic_a.filtered_out[3] ),
    .Y(_1119_));
 sg13g2_nor2_1 _2953_ (.A(_1114_),
    .B(_1116_),
    .Y(_1120_));
 sg13g2_nand2b_1 _2954_ (.Y(_1121_),
    .B(\cic_b.filtered_out[3] ),
    .A_N(\cic_a.filtered_out[3] ));
 sg13g2_xnor2_1 _2955_ (.Y(_1122_),
    .A(\cic_a.filtered_out[3] ),
    .B(\cic_b.filtered_out[3] ));
 sg13g2_xor2_1 _2956_ (.B(_1122_),
    .A(_1120_),
    .X(_1123_));
 sg13g2_a22oi_1 _2957_ (.Y(_1124_),
    .B1(net444),
    .B2(net532),
    .A2(net418),
    .A1(net541));
 sg13g2_o21ai_1 _2958_ (.B1(net445),
    .Y(_0401_),
    .A1(net537),
    .A2(_1123_));
 sg13g2_nor2b_1 _2959_ (.A(\cic_b.filtered_out[4] ),
    .B_N(\cic_a.filtered_out[4] ),
    .Y(_1125_));
 sg13g2_xor2_1 _2960_ (.B(\cic_b.filtered_out[4] ),
    .A(\cic_a.filtered_out[4] ),
    .X(_1126_));
 sg13g2_a21oi_1 _2961_ (.A1(_1114_),
    .A2(_1121_),
    .Y(_1127_),
    .B1(_1119_));
 sg13g2_nand2b_1 _2962_ (.Y(_1128_),
    .B(_1122_),
    .A_N(_1115_));
 sg13g2_o21ai_1 _2963_ (.B1(_1127_),
    .Y(_1129_),
    .A1(_1113_),
    .A2(_1128_));
 sg13g2_nor2b_1 _2964_ (.A(_1126_),
    .B_N(_1129_),
    .Y(_1130_));
 sg13g2_xor2_1 _2965_ (.B(_1129_),
    .A(_1126_),
    .X(_1131_));
 sg13g2_a22oi_1 _2966_ (.Y(_1132_),
    .B1(net404),
    .B2(net532),
    .A2(\serializer_ab_subtr.shift_reg[3] ),
    .A1(net541));
 sg13g2_o21ai_1 _2967_ (.B1(net405),
    .Y(_0402_),
    .A1(net536),
    .A2(_1131_));
 sg13g2_nor2_1 _2968_ (.A(\cic_a.filtered_out[5] ),
    .B(_1202_),
    .Y(_1133_));
 sg13g2_xor2_1 _2969_ (.B(\cic_b.filtered_out[5] ),
    .A(\cic_a.filtered_out[5] ),
    .X(_1134_));
 sg13g2_nor2_1 _2970_ (.A(_1125_),
    .B(_1130_),
    .Y(_1135_));
 sg13g2_xnor2_1 _2971_ (.Y(_1136_),
    .A(_1134_),
    .B(_1135_));
 sg13g2_a22oi_1 _2972_ (.Y(_1137_),
    .B1(net377),
    .B2(net532),
    .A2(\serializer_ab_subtr.shift_reg[4] ),
    .A1(net541));
 sg13g2_o21ai_1 _2973_ (.B1(net378),
    .Y(_0403_),
    .A1(net536),
    .A2(_1136_));
 sg13g2_nand2b_1 _2974_ (.Y(_1138_),
    .B(\cic_a.filtered_out[6] ),
    .A_N(\cic_b.filtered_out[6] ));
 sg13g2_xor2_1 _2975_ (.B(\cic_b.filtered_out[6] ),
    .A(\cic_a.filtered_out[6] ),
    .X(_1139_));
 sg13g2_a21oi_1 _2976_ (.A1(\cic_a.filtered_out[5] ),
    .A2(_1202_),
    .Y(_1140_),
    .B1(_1125_));
 sg13g2_nor2b_1 _2977_ (.A(_1130_),
    .B_N(_1140_),
    .Y(_1141_));
 sg13g2_or2_1 _2978_ (.X(_1142_),
    .B(_1141_),
    .A(_1133_));
 sg13g2_xnor2_1 _2979_ (.Y(_1143_),
    .A(_1139_),
    .B(_1142_));
 sg13g2_a22oi_1 _2980_ (.Y(_1144_),
    .B1(net368),
    .B2(net532),
    .A2(\serializer_ab_subtr.shift_reg[5] ),
    .A1(net541));
 sg13g2_o21ai_1 _2981_ (.B1(net369),
    .Y(_0404_),
    .A1(net536),
    .A2(_1143_));
 sg13g2_nand2_1 _2982_ (.Y(_1145_),
    .A(_1196_),
    .B(\cic_b.filtered_out[7] ));
 sg13g2_xor2_1 _2983_ (.B(\cic_b.filtered_out[7] ),
    .A(\cic_a.filtered_out[7] ),
    .X(_1146_));
 sg13g2_o21ai_1 _2984_ (.B1(_1138_),
    .Y(_1147_),
    .A1(_1139_),
    .A2(_1142_));
 sg13g2_xor2_1 _2985_ (.B(_1147_),
    .A(_1146_),
    .X(_1148_));
 sg13g2_a22oi_1 _2986_ (.Y(_1149_),
    .B1(net410),
    .B2(net532),
    .A2(net368),
    .A1(net541));
 sg13g2_o21ai_1 _2987_ (.B1(net411),
    .Y(_0405_),
    .A1(net536),
    .A2(_1148_));
 sg13g2_nor4_1 _2988_ (.A(_1126_),
    .B(_1134_),
    .C(_1139_),
    .D(_1146_),
    .Y(_1150_));
 sg13g2_nor4_1 _2989_ (.A(_1133_),
    .B(_1139_),
    .C(_1140_),
    .D(_1146_),
    .Y(_1151_));
 sg13g2_o21ai_1 _2990_ (.B1(_1138_),
    .Y(_1152_),
    .A1(_1196_),
    .A2(\cic_b.filtered_out[7] ));
 sg13g2_a221oi_1 _2991_ (.B2(_1145_),
    .C1(_1151_),
    .B1(_1152_),
    .A1(_1129_),
    .Y(_1153_),
    .A2(_1150_));
 sg13g2_nor2b_1 _2992_ (.A(\cic_b.filtered_out[8] ),
    .B_N(\cic_a.filtered_out[8] ),
    .Y(_1154_));
 sg13g2_xor2_1 _2993_ (.B(\cic_b.filtered_out[8] ),
    .A(\cic_a.filtered_out[8] ),
    .X(_1155_));
 sg13g2_nor2_1 _2994_ (.A(_1153_),
    .B(_1155_),
    .Y(_1156_));
 sg13g2_a21o_1 _2995_ (.A2(_1155_),
    .A1(_1153_),
    .B1(net536),
    .X(_1157_));
 sg13g2_a22oi_1 _2996_ (.Y(_1158_),
    .B1(net407),
    .B2(net532),
    .A2(\serializer_ab_subtr.shift_reg[7] ),
    .A1(net541));
 sg13g2_o21ai_1 _2997_ (.B1(net408),
    .Y(_0406_),
    .A1(_1156_),
    .A2(_1157_));
 sg13g2_nor2b_1 _2998_ (.A(\cic_b.filtered_out[9] ),
    .B_N(\cic_a.filtered_out[9] ),
    .Y(_1159_));
 sg13g2_nand2b_1 _2999_ (.Y(_1160_),
    .B(\cic_b.filtered_out[9] ),
    .A_N(\cic_a.filtered_out[9] ));
 sg13g2_nand2b_1 _3000_ (.Y(_1161_),
    .B(_1160_),
    .A_N(_1159_));
 sg13g2_nor2_1 _3001_ (.A(_1154_),
    .B(_1156_),
    .Y(_1162_));
 sg13g2_xnor2_1 _3002_ (.Y(_1163_),
    .A(_1161_),
    .B(_1162_));
 sg13g2_a22oi_1 _3003_ (.Y(_1164_),
    .B1(net463),
    .B2(net532),
    .A2(net407),
    .A1(net541));
 sg13g2_o21ai_1 _3004_ (.B1(net464),
    .Y(_0407_),
    .A1(net536),
    .A2(_1163_));
 sg13g2_nor2b_1 _3005_ (.A(\cic_b.filtered_out[10] ),
    .B_N(\cic_a.filtered_out[10] ),
    .Y(_1165_));
 sg13g2_xnor2_1 _3006_ (.Y(_1166_),
    .A(\cic_a.filtered_out[10] ),
    .B(\cic_b.filtered_out[10] ));
 sg13g2_or2_1 _3007_ (.X(_1167_),
    .B(_1161_),
    .A(_1155_));
 sg13g2_a21oi_1 _3008_ (.A1(_1154_),
    .A2(_1160_),
    .Y(_1168_),
    .B1(_1159_));
 sg13g2_o21ai_1 _3009_ (.B1(_1168_),
    .Y(_1169_),
    .A1(_1153_),
    .A2(_1167_));
 sg13g2_and2_1 _3010_ (.A(_1166_),
    .B(_1169_),
    .X(_1170_));
 sg13g2_o21ai_1 _3011_ (.B1(_0019_),
    .Y(_1171_),
    .A1(_1166_),
    .A2(_1169_));
 sg13g2_a22oi_1 _3012_ (.Y(_1172_),
    .B1(net354),
    .B2(net532),
    .A2(\serializer_ab_subtr.shift_reg[9] ),
    .A1(net541));
 sg13g2_o21ai_1 _3013_ (.B1(net355),
    .Y(_0408_),
    .A1(_1170_),
    .A2(_1171_));
 sg13g2_nor2b_1 _3014_ (.A(\cic_a.filtered_out[11] ),
    .B_N(\cic_b.filtered_out[11] ),
    .Y(_1173_));
 sg13g2_nand2b_1 _3015_ (.Y(_1174_),
    .B(\cic_a.filtered_out[11] ),
    .A_N(\cic_b.filtered_out[11] ));
 sg13g2_nand2b_1 _3016_ (.Y(_1175_),
    .B(_1174_),
    .A_N(_1173_));
 sg13g2_a21oi_1 _3017_ (.A1(_1166_),
    .A2(_1169_),
    .Y(_1176_),
    .B1(_1165_));
 sg13g2_xnor2_1 _3018_ (.Y(_1177_),
    .A(_1175_),
    .B(_1176_));
 sg13g2_a22oi_1 _3019_ (.Y(_1178_),
    .B1(net350),
    .B2(net533),
    .A2(\serializer_ab_subtr.shift_reg[10] ),
    .A1(net540));
 sg13g2_o21ai_1 _3020_ (.B1(net351),
    .Y(_0409_),
    .A1(net537),
    .A2(_1177_));
 sg13g2_xnor2_1 _3021_ (.Y(_1179_),
    .A(\cic_a.filtered_out[12] ),
    .B(\cic_b.filtered_out[12] ));
 sg13g2_o21ai_1 _3022_ (.B1(_1174_),
    .Y(_1180_),
    .A1(_1173_),
    .A2(_1176_));
 sg13g2_xnor2_1 _3023_ (.Y(_1181_),
    .A(_1179_),
    .B(_1180_));
 sg13g2_a22oi_1 _3024_ (.Y(_1182_),
    .B1(net400),
    .B2(net533),
    .A2(net350),
    .A1(net540));
 sg13g2_o21ai_1 _3025_ (.B1(_1182_),
    .Y(_0410_),
    .A1(net537),
    .A2(_1181_));
 sg13g2_nor2_1 _3026_ (.A(net546),
    .B(net155),
    .Y(_1183_));
 sg13g2_a21oi_1 _3027_ (.A1(net155),
    .A2(net531),
    .Y(_0411_),
    .B1(_1183_));
 sg13g2_nand2_1 _3028_ (.Y(_1184_),
    .A(net151),
    .B(_0586_));
 sg13g2_and2_1 _3029_ (.A(\serializer_a.bit_cnt[0] ),
    .B(net151),
    .X(_1185_));
 sg13g2_o21ai_1 _3030_ (.B1(_1184_),
    .Y(_0412_),
    .A1(_0588_),
    .A2(_1185_));
 sg13g2_nand3_1 _3031_ (.B(net52),
    .C(_1185_),
    .A(net546),
    .Y(_1186_));
 sg13g2_nand2b_1 _3032_ (.Y(_1187_),
    .B(_1186_),
    .A_N(net539));
 sg13g2_a21oi_1 _3033_ (.A1(net530),
    .A2(_1185_),
    .Y(_1188_),
    .B1(net52));
 sg13g2_nor2_1 _3034_ (.A(_1187_),
    .B(net53),
    .Y(_0413_));
 sg13g2_nor2b_1 _3035_ (.A(net48),
    .B_N(_1186_),
    .Y(_1189_));
 sg13g2_a21oi_1 _3036_ (.A1(net48),
    .A2(_1187_),
    .Y(_0414_),
    .B1(_1189_));
 sg13g2_dfrbp_1 _3037_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net612),
    .D(_0102_),
    .Q_N(\cic_a.pdm_in ),
    .Q(_0100_));
 sg13g2_dfrbp_1 _3038_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net595),
    .D(_0103_),
    .Q_N(\cic_b.pdm_in ),
    .Q(_0101_));
 sg13g2_dfrbp_1 _3039_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net605),
    .D(_0104_),
    .Q_N(_1623_),
    .Q(\cic_a.delay[2][0] ));
 sg13g2_dfrbp_1 _3040_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net605),
    .D(_0105_),
    .Q_N(_1622_),
    .Q(\cic_a.delay[2][1] ));
 sg13g2_dfrbp_1 _3041_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net603),
    .D(_0106_),
    .Q_N(_1621_),
    .Q(\cic_a.delay[2][2] ));
 sg13g2_dfrbp_1 _3042_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net577),
    .D(_0107_),
    .Q_N(_1620_),
    .Q(\cic_a.delay[2][3] ));
 sg13g2_dfrbp_1 _3043_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net575),
    .D(_0108_),
    .Q_N(_1619_),
    .Q(\cic_a.delay[2][4] ));
 sg13g2_dfrbp_1 _3044_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net576),
    .D(net398),
    .Q_N(_1618_),
    .Q(\cic_a.delay[2][5] ));
 sg13g2_dfrbp_1 _3045_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net575),
    .D(_0110_),
    .Q_N(_1617_),
    .Q(\cic_a.delay[2][6] ));
 sg13g2_dfrbp_1 _3046_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net570),
    .D(net255),
    .Q_N(_1616_),
    .Q(\cic_a.delay[2][7] ));
 sg13g2_dfrbp_1 _3047_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net575),
    .D(net72),
    .Q_N(_1615_),
    .Q(\cic_a.delay[2][8] ));
 sg13g2_dfrbp_1 _3048_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net569),
    .D(_0113_),
    .Q_N(_1614_),
    .Q(\cic_a.delay[2][9] ));
 sg13g2_dfrbp_1 _3049_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net572),
    .D(net247),
    .Q_N(_1613_),
    .Q(\cic_a.delay[2][10] ));
 sg13g2_dfrbp_1 _3050_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net572),
    .D(_0115_),
    .Q_N(_1612_),
    .Q(\cic_a.delay[2][11] ));
 sg13g2_dfrbp_1 _3051_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net572),
    .D(_0116_),
    .Q_N(_1611_),
    .Q(\cic_a.delay[2][12] ));
 sg13g2_dfrbp_1 _3052_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net606),
    .D(_0117_),
    .Q_N(_1610_),
    .Q(\cic_a.temp_comb[1][0] ));
 sg13g2_dfrbp_1 _3053_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net603),
    .D(_0118_),
    .Q_N(_1609_),
    .Q(\cic_a.temp_comb[1][1] ));
 sg13g2_dfrbp_1 _3054_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net603),
    .D(_0119_),
    .Q_N(_1608_),
    .Q(\cic_a.temp_comb[1][2] ));
 sg13g2_dfrbp_1 _3055_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net577),
    .D(net686),
    .Q_N(_1607_),
    .Q(\cic_a.temp_comb[1][3] ));
 sg13g2_dfrbp_1 _3056_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net576),
    .D(_0121_),
    .Q_N(_1606_),
    .Q(\cic_a.temp_comb[1][4] ));
 sg13g2_dfrbp_1 _3057_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net570),
    .D(_0122_),
    .Q_N(_1605_),
    .Q(\cic_a.temp_comb[1][5] ));
 sg13g2_dfrbp_1 _3058_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net570),
    .D(_0123_),
    .Q_N(_1604_),
    .Q(\cic_a.temp_comb[1][6] ));
 sg13g2_dfrbp_1 _3059_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net570),
    .D(_0124_),
    .Q_N(_1603_),
    .Q(\cic_a.temp_comb[1][7] ));
 sg13g2_dfrbp_1 _3060_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net569),
    .D(_0125_),
    .Q_N(_1602_),
    .Q(\cic_a.temp_comb[1][8] ));
 sg13g2_dfrbp_1 _3061_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net569),
    .D(_0126_),
    .Q_N(_1601_),
    .Q(\cic_a.temp_comb[1][9] ));
 sg13g2_dfrbp_1 _3062_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net564),
    .D(_0127_),
    .Q_N(_1600_),
    .Q(\cic_a.temp_comb[1][10] ));
 sg13g2_dfrbp_1 _3063_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net564),
    .D(_0128_),
    .Q_N(_1599_),
    .Q(\cic_a.temp_comb[1][11] ));
 sg13g2_dfrbp_1 _3064_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net572),
    .D(_0129_),
    .Q_N(_1598_),
    .Q(\cic_a.temp_comb[1][12] ));
 sg13g2_dfrbp_1 _3065_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net607),
    .D(_0130_),
    .Q_N(_1597_),
    .Q(\cic_a.delay[1][0] ));
 sg13g2_dfrbp_1 _3066_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net603),
    .D(_0131_),
    .Q_N(_1596_),
    .Q(\cic_a.delay[1][1] ));
 sg13g2_dfrbp_1 _3067_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net578),
    .D(_0132_),
    .Q_N(_1595_),
    .Q(\cic_a.delay[1][2] ));
 sg13g2_dfrbp_1 _3068_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net576),
    .D(_0133_),
    .Q_N(_1594_),
    .Q(\cic_a.delay[1][3] ));
 sg13g2_dfrbp_1 _3069_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net569),
    .D(_0134_),
    .Q_N(_1593_),
    .Q(\cic_a.delay[1][4] ));
 sg13g2_dfrbp_1 _3070_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net568),
    .D(_0135_),
    .Q_N(_1592_),
    .Q(\cic_a.delay[1][5] ));
 sg13g2_dfrbp_1 _3071_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net567),
    .D(net140),
    .Q_N(_1591_),
    .Q(\cic_a.delay[1][6] ));
 sg13g2_dfrbp_1 _3072_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net567),
    .D(_0137_),
    .Q_N(_1590_),
    .Q(\cic_a.delay[1][7] ));
 sg13g2_dfrbp_1 _3073_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net567),
    .D(_0138_),
    .Q_N(_1589_),
    .Q(\cic_a.delay[1][8] ));
 sg13g2_dfrbp_1 _3074_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net567),
    .D(net51),
    .Q_N(_1588_),
    .Q(\cic_a.delay[1][9] ));
 sg13g2_dfrbp_1 _3075_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net564),
    .D(_0140_),
    .Q_N(_1587_),
    .Q(\cic_a.delay[1][10] ));
 sg13g2_dfrbp_1 _3076_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net563),
    .D(_0141_),
    .Q_N(_1586_),
    .Q(\cic_a.delay[1][11] ));
 sg13g2_dfrbp_1 _3077_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net563),
    .D(_0142_),
    .Q_N(_1585_),
    .Q(\cic_a.delay[1][12] ));
 sg13g2_dfrbp_1 _3078_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net604),
    .D(_0143_),
    .Q_N(_1584_),
    .Q(\cic_a.delay[0][0] ));
 sg13g2_dfrbp_1 _3079_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net577),
    .D(_0144_),
    .Q_N(_1583_),
    .Q(\cic_a.delay[0][1] ));
 sg13g2_dfrbp_1 _3080_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net577),
    .D(net111),
    .Q_N(_1582_),
    .Q(\cic_a.delay[0][2] ));
 sg13g2_dfrbp_1 _3081_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net573),
    .D(net142),
    .Q_N(_1581_),
    .Q(\cic_a.delay[0][3] ));
 sg13g2_dfrbp_1 _3082_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net566),
    .D(_0147_),
    .Q_N(_1580_),
    .Q(\cic_a.delay[0][4] ));
 sg13g2_dfrbp_1 _3083_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net566),
    .D(net23),
    .Q_N(_1579_),
    .Q(\cic_a.delay[0][5] ));
 sg13g2_dfrbp_1 _3084_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net566),
    .D(_0149_),
    .Q_N(_1578_),
    .Q(\cic_a.delay[0][6] ));
 sg13g2_dfrbp_1 _3085_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net566),
    .D(net42),
    .Q_N(_1577_),
    .Q(\cic_a.delay[0][7] ));
 sg13g2_dfrbp_1 _3086_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net563),
    .D(_0151_),
    .Q_N(_1576_),
    .Q(\cic_a.delay[0][8] ));
 sg13g2_dfrbp_1 _3087_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net564),
    .D(_0152_),
    .Q_N(_1575_),
    .Q(\cic_a.delay[0][9] ));
 sg13g2_dfrbp_1 _3088_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net552),
    .D(net55),
    .Q_N(_1574_),
    .Q(\cic_a.delay[0][10] ));
 sg13g2_dfrbp_1 _3089_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net552),
    .D(_0154_),
    .Q_N(_1573_),
    .Q(\cic_a.delay[0][11] ));
 sg13g2_dfrbp_1 _3090_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net551),
    .D(_0155_),
    .Q_N(_1572_),
    .Q(\cic_a.delay[0][12] ));
 sg13g2_dfrbp_1 _3091_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net603),
    .D(net624),
    .Q_N(_1571_),
    .Q(\cic_a.temp_comb[0][0] ));
 sg13g2_dfrbp_1 _3092_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net604),
    .D(_0157_),
    .Q_N(_1570_),
    .Q(\cic_a.temp_comb[0][1] ));
 sg13g2_dfrbp_1 _3093_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net577),
    .D(net658),
    .Q_N(_1569_),
    .Q(\cic_a.temp_comb[0][2] ));
 sg13g2_dfrbp_1 _3094_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net575),
    .D(net649),
    .Q_N(_1568_),
    .Q(\cic_a.temp_comb[0][3] ));
 sg13g2_dfrbp_1 _3095_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net569),
    .D(_0160_),
    .Q_N(_1567_),
    .Q(\cic_a.temp_comb[0][4] ));
 sg13g2_dfrbp_1 _3096_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net569),
    .D(_0161_),
    .Q_N(_1566_),
    .Q(\cic_a.temp_comb[0][5] ));
 sg13g2_dfrbp_1 _3097_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net568),
    .D(_0162_),
    .Q_N(_1565_),
    .Q(\cic_a.temp_comb[0][6] ));
 sg13g2_dfrbp_1 _3098_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net567),
    .D(_0163_),
    .Q_N(_1564_),
    .Q(\cic_a.temp_comb[0][7] ));
 sg13g2_dfrbp_1 _3099_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net564),
    .D(_0164_),
    .Q_N(_1563_),
    .Q(\cic_a.temp_comb[0][8] ));
 sg13g2_dfrbp_1 _3100_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net564),
    .D(_0165_),
    .Q_N(_1562_),
    .Q(\cic_a.temp_comb[0][9] ));
 sg13g2_dfrbp_1 _3101_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net563),
    .D(_0166_),
    .Q_N(_1561_),
    .Q(\cic_a.temp_comb[0][10] ));
 sg13g2_dfrbp_1 _3102_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net563),
    .D(net442),
    .Q_N(_1560_),
    .Q(\cic_a.temp_comb[0][11] ));
 sg13g2_dfrbp_1 _3103_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net552),
    .D(net661),
    .Q_N(_1559_),
    .Q(\cic_a.temp_comb[0][12] ));
 sg13g2_dfrbp_1 _3104_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net613),
    .D(_0169_),
    .Q_N(_1558_),
    .Q(\cic_a.filtered_out[0] ));
 sg13g2_dfrbp_1 _3105_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net613),
    .D(_0170_),
    .Q_N(_1557_),
    .Q(\cic_a.filtered_out[1] ));
 sg13g2_dfrbp_1 _3106_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net613),
    .D(_0171_),
    .Q_N(_1556_),
    .Q(\cic_a.filtered_out[2] ));
 sg13g2_dfrbp_1 _3107_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net605),
    .D(_0172_),
    .Q_N(_1555_),
    .Q(\cic_a.filtered_out[3] ));
 sg13g2_dfrbp_1 _3108_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net606),
    .D(_0173_),
    .Q_N(_1554_),
    .Q(\cic_a.filtered_out[4] ));
 sg13g2_dfrbp_1 _3109_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net606),
    .D(_0174_),
    .Q_N(_1553_),
    .Q(\cic_a.filtered_out[5] ));
 sg13g2_dfrbp_1 _3110_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net604),
    .D(_0175_),
    .Q_N(_1552_),
    .Q(\cic_a.filtered_out[6] ));
 sg13g2_dfrbp_1 _3111_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net606),
    .D(net95),
    .Q_N(_1551_),
    .Q(\cic_a.filtered_out[7] ));
 sg13g2_dfrbp_1 _3112_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net606),
    .D(_0177_),
    .Q_N(_1550_),
    .Q(\cic_a.filtered_out[8] ));
 sg13g2_dfrbp_1 _3113_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net602),
    .D(_0178_),
    .Q_N(_1549_),
    .Q(\cic_a.filtered_out[9] ));
 sg13g2_dfrbp_1 _3114_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net600),
    .D(_0179_),
    .Q_N(_1548_),
    .Q(\cic_a.filtered_out[10] ));
 sg13g2_dfrbp_1 _3115_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net600),
    .D(_0180_),
    .Q_N(_1547_),
    .Q(\cic_a.filtered_out[11] ));
 sg13g2_dfrbp_1 _3116_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net600),
    .D(_0181_),
    .Q_N(_1546_),
    .Q(\cic_a.filtered_out[12] ));
 sg13g2_dfrbp_1 _3117_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net617),
    .D(net120),
    .Q_N(_1545_),
    .Q(\cic_a.temp_comb[2][0] ));
 sg13g2_dfrbp_1 _3118_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net613),
    .D(net115),
    .Q_N(_1544_),
    .Q(\cic_a.temp_comb[2][1] ));
 sg13g2_dfrbp_1 _3119_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net606),
    .D(_0184_),
    .Q_N(_1543_),
    .Q(\cic_a.temp_comb[2][2] ));
 sg13g2_dfrbp_1 _3120_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net605),
    .D(_0185_),
    .Q_N(_1542_),
    .Q(\cic_a.temp_comb[2][3] ));
 sg13g2_dfrbp_1 _3121_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net605),
    .D(_0186_),
    .Q_N(_1541_),
    .Q(\cic_a.temp_comb[2][4] ));
 sg13g2_dfrbp_1 _3122_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net605),
    .D(_0187_),
    .Q_N(_1540_),
    .Q(\cic_a.temp_comb[2][5] ));
 sg13g2_dfrbp_1 _3123_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net604),
    .D(_0188_),
    .Q_N(_1539_),
    .Q(\cic_a.temp_comb[2][6] ));
 sg13g2_dfrbp_1 _3124_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net606),
    .D(_0189_),
    .Q_N(_1538_),
    .Q(\cic_a.temp_comb[2][7] ));
 sg13g2_dfrbp_1 _3125_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net604),
    .D(_0190_),
    .Q_N(_1537_),
    .Q(\cic_a.temp_comb[2][8] ));
 sg13g2_dfrbp_1 _3126_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net604),
    .D(_0191_),
    .Q_N(_1536_),
    .Q(\cic_a.temp_comb[2][9] ));
 sg13g2_dfrbp_1 _3127_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net600),
    .D(_0192_),
    .Q_N(_1535_),
    .Q(\cic_a.temp_comb[2][10] ));
 sg13g2_dfrbp_1 _3128_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net600),
    .D(_0193_),
    .Q_N(_1534_),
    .Q(\cic_a.temp_comb[2][11] ));
 sg13g2_dfrbp_1 _3129_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net599),
    .D(net413),
    .Q_N(_1624_),
    .Q(\cic_a.temp_comb[2][12] ));
 sg13g2_dfrbp_1 _3130_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net604),
    .D(net459),
    .Q_N(_1625_),
    .Q(\cic_a.integrator[2][0] ));
 sg13g2_dfrbp_1 _3131_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net574),
    .D(net713),
    .Q_N(_1626_),
    .Q(\cic_a.integrator[2][1] ));
 sg13g2_dfrbp_1 _3132_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net574),
    .D(net774),
    .Q_N(_1627_),
    .Q(\cic_a.integrator[2][2] ));
 sg13g2_dfrbp_1 _3133_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net573),
    .D(net736),
    .Q_N(_1628_),
    .Q(\cic_a.integrator[2][3] ));
 sg13g2_dfrbp_1 _3134_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net565),
    .D(net787),
    .Q_N(_1629_),
    .Q(\cic_a.integrator[2][4] ));
 sg13g2_dfrbp_1 _3135_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net565),
    .D(_0056_),
    .Q_N(_1630_),
    .Q(\cic_a.integrator[2][5] ));
 sg13g2_dfrbp_1 _3136_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net565),
    .D(_0057_),
    .Q_N(_1631_),
    .Q(\cic_a.integrator[2][6] ));
 sg13g2_dfrbp_1 _3137_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net565),
    .D(net768),
    .Q_N(_1632_),
    .Q(\cic_a.integrator[2][7] ));
 sg13g2_dfrbp_1 _3138_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net554),
    .D(_0059_),
    .Q_N(_1633_),
    .Q(\cic_a.integrator[2][8] ));
 sg13g2_dfrbp_1 _3139_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net554),
    .D(net726),
    .Q_N(_1634_),
    .Q(\cic_a.integrator[2][9] ));
 sg13g2_dfrbp_1 _3140_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net554),
    .D(_0049_),
    .Q_N(_1635_),
    .Q(\cic_a.integrator[2][10] ));
 sg13g2_dfrbp_1 _3141_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net551),
    .D(_0050_),
    .Q_N(_1636_),
    .Q(\cic_a.integrator[2][11] ));
 sg13g2_dfrbp_1 _3142_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net551),
    .D(net702),
    .Q_N(_1637_),
    .Q(\cic_a.integrator[2][12] ));
 sg13g2_dfrbp_1 _3143_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net600),
    .D(_0035_),
    .Q_N(_1638_),
    .Q(\cic_a.integrator[1][0] ));
 sg13g2_dfrbp_1 _3144_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net574),
    .D(_0039_),
    .Q_N(_1639_),
    .Q(\cic_a.integrator[1][1] ));
 sg13g2_dfrbp_1 _3145_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net574),
    .D(_0040_),
    .Q_N(_1640_),
    .Q(\cic_a.integrator[1][2] ));
 sg13g2_dfrbp_1 _3146_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net579),
    .D(_0041_),
    .Q_N(_1641_),
    .Q(\cic_a.integrator[1][3] ));
 sg13g2_dfrbp_1 _3147_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net572),
    .D(net783),
    .Q_N(_1642_),
    .Q(\cic_a.integrator[1][4] ));
 sg13g2_dfrbp_1 _3148_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net572),
    .D(_0043_),
    .Q_N(_1643_),
    .Q(\cic_a.integrator[1][5] ));
 sg13g2_dfrbp_1 _3149_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net565),
    .D(_0044_),
    .Q_N(_1644_),
    .Q(\cic_a.integrator[1][6] ));
 sg13g2_dfrbp_1 _3150_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net565),
    .D(net741),
    .Q_N(_1645_),
    .Q(\cic_a.integrator[1][7] ));
 sg13g2_dfrbp_1 _3151_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net553),
    .D(_0046_),
    .Q_N(_1646_),
    .Q(\cic_a.integrator[1][8] ));
 sg13g2_dfrbp_1 _3152_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net553),
    .D(net747),
    .Q_N(_1647_),
    .Q(\cic_a.integrator[1][9] ));
 sg13g2_dfrbp_1 _3153_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net552),
    .D(net755),
    .Q_N(_1648_),
    .Q(\cic_a.integrator[1][10] ));
 sg13g2_dfrbp_1 _3154_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net551),
    .D(net731),
    .Q_N(_1649_),
    .Q(\cic_a.integrator[1][11] ));
 sg13g2_dfrbp_1 _3155_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net551),
    .D(net699),
    .Q_N(_1650_),
    .Q(\cic_a.integrator[1][12] ));
 sg13g2_dfrbp_1 _3156_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net600),
    .D(net40),
    .Q_N(_1651_),
    .Q(\cic_a.integrator[0][0] ));
 sg13g2_dfrbp_1 _3157_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net599),
    .D(_0026_),
    .Q_N(_1652_),
    .Q(\cic_a.integrator[0][1] ));
 sg13g2_dfrbp_1 _3158_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net574),
    .D(net430),
    .Q_N(_1653_),
    .Q(\cic_a.integrator[0][2] ));
 sg13g2_dfrbp_1 _3159_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net579),
    .D(net684),
    .Q_N(_1654_),
    .Q(\cic_a.integrator[0][3] ));
 sg13g2_dfrbp_1 _3160_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net561),
    .D(_0029_),
    .Q_N(_1655_),
    .Q(\cic_a.integrator[0][4] ));
 sg13g2_dfrbp_1 _3161_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net561),
    .D(net672),
    .Q_N(_1656_),
    .Q(\cic_a.integrator[0][5] ));
 sg13g2_dfrbp_1 _3162_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net561),
    .D(net678),
    .Q_N(_1657_),
    .Q(\cic_a.integrator[0][6] ));
 sg13g2_dfrbp_1 _3163_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net554),
    .D(net689),
    .Q_N(_1658_),
    .Q(\cic_a.integrator[0][7] ));
 sg13g2_dfrbp_1 _3164_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net553),
    .D(net716),
    .Q_N(_1659_),
    .Q(\cic_a.integrator[0][8] ));
 sg13g2_dfrbp_1 _3165_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net553),
    .D(net628),
    .Q_N(_1660_),
    .Q(\cic_a.integrator[0][9] ));
 sg13g2_dfrbp_1 _3166_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net553),
    .D(_0023_),
    .Q_N(_1661_),
    .Q(\cic_a.integrator[0][10] ));
 sg13g2_dfrbp_1 _3167_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net553),
    .D(_0024_),
    .Q_N(_1662_),
    .Q(\cic_a.integrator[0][11] ));
 sg13g2_dfrbp_1 _3168_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net551),
    .D(net101),
    .Q_N(_1533_),
    .Q(\cic_a.integrator[0][12] ));
 sg13g2_dfrbp_1 _3169_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net604),
    .D(net198),
    .Q_N(_1532_),
    .Q(\cic_a.temp_delay[0][0] ));
 sg13g2_dfrbp_1 _3170_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net577),
    .D(net238),
    .Q_N(_1531_),
    .Q(\cic_a.temp_delay[0][1] ));
 sg13g2_dfrbp_1 _3171_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net574),
    .D(_0197_),
    .Q_N(_1530_),
    .Q(\cic_a.temp_delay[0][2] ));
 sg13g2_dfrbp_1 _3172_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net573),
    .D(_0198_),
    .Q_N(_1529_),
    .Q(\cic_a.temp_delay[0][3] ));
 sg13g2_dfrbp_1 _3173_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net566),
    .D(net345),
    .Q_N(_1528_),
    .Q(\cic_a.temp_delay[0][4] ));
 sg13g2_dfrbp_1 _3174_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net566),
    .D(_0200_),
    .Q_N(_1527_),
    .Q(\cic_a.temp_delay[0][5] ));
 sg13g2_dfrbp_1 _3175_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net565),
    .D(net328),
    .Q_N(_1526_),
    .Q(\cic_a.temp_delay[0][6] ));
 sg13g2_dfrbp_1 _3176_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net565),
    .D(_0202_),
    .Q_N(_1525_),
    .Q(\cic_a.temp_delay[0][7] ));
 sg13g2_dfrbp_1 _3177_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net563),
    .D(net190),
    .Q_N(_1524_),
    .Q(\cic_a.temp_delay[0][8] ));
 sg13g2_dfrbp_1 _3178_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net552),
    .D(net99),
    .Q_N(_1523_),
    .Q(\cic_a.temp_delay[0][9] ));
 sg13g2_dfrbp_1 _3179_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net552),
    .D(_0205_),
    .Q_N(_1522_),
    .Q(\cic_a.temp_delay[0][10] ));
 sg13g2_dfrbp_1 _3180_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net551),
    .D(net228),
    .Q_N(_1521_),
    .Q(\cic_a.temp_delay[0][11] ));
 sg13g2_dfrbp_1 _3181_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net551),
    .D(net307),
    .Q_N(_1663_),
    .Q(\cic_a.temp_delay[0][12] ));
 sg13g2_dfrbp_1 _3182_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net550),
    .D(_0000_),
    .Q_N(_1664_),
    .Q(\cic_a.decim_cnt[0] ));
 sg13g2_dfrbp_1 _3183_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net548),
    .D(_0001_),
    .Q_N(_1665_),
    .Q(\cic_a.decim_cnt[1] ));
 sg13g2_dfrbp_1 _3184_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net548),
    .D(net32),
    .Q_N(_1666_),
    .Q(\cic_a.decim_cnt[2] ));
 sg13g2_dfrbp_1 _3185_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net550),
    .D(_0003_),
    .Q_N(_1667_),
    .Q(\cic_a.decim_cnt[3] ));
 sg13g2_dfrbp_1 _3186_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net550),
    .D(_0004_),
    .Q_N(_1668_),
    .Q(\cic_a.decim_cnt[4] ));
 sg13g2_dfrbp_1 _3187_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net548),
    .D(net292),
    .Q_N(_1669_),
    .Q(\cic_a.decim_cnt[5] ));
 sg13g2_dfrbp_1 _3188_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net548),
    .D(net245),
    .Q_N(_1670_),
    .Q(\cic_a.decim_cnt[6] ));
 sg13g2_dfrbp_1 _3189_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net548),
    .D(net57),
    .Q_N(_1520_),
    .Q(\cic_a.decim_cnt[7] ));
 sg13g2_dfrbp_1 _3190_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net603),
    .D(net129),
    .Q_N(_1519_),
    .Q(\cic_a.temp_delay[1][0] ));
 sg13g2_dfrbp_1 _3191_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net603),
    .D(net310),
    .Q_N(_1518_),
    .Q(\cic_a.temp_delay[1][1] ));
 sg13g2_dfrbp_1 _3192_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net577),
    .D(net168),
    .Q_N(_1517_),
    .Q(\cic_a.temp_delay[1][2] ));
 sg13g2_dfrbp_1 _3193_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net575),
    .D(net157),
    .Q_N(_1516_),
    .Q(\cic_a.temp_delay[1][3] ));
 sg13g2_dfrbp_1 _3194_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net569),
    .D(net394),
    .Q_N(_1515_),
    .Q(\cic_a.temp_delay[1][4] ));
 sg13g2_dfrbp_1 _3195_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net568),
    .D(net226),
    .Q_N(_1514_),
    .Q(\cic_a.temp_delay[1][5] ));
 sg13g2_dfrbp_1 _3196_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net567),
    .D(_0214_),
    .Q_N(_1513_),
    .Q(\cic_a.temp_delay[1][6] ));
 sg13g2_dfrbp_1 _3197_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net567),
    .D(net253),
    .Q_N(_1512_),
    .Q(\cic_a.temp_delay[1][7] ));
 sg13g2_dfrbp_1 _3198_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net564),
    .D(net365),
    .Q_N(_1511_),
    .Q(\cic_a.temp_delay[1][8] ));
 sg13g2_dfrbp_1 _3199_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net567),
    .D(_0217_),
    .Q_N(_1510_),
    .Q(\cic_a.temp_delay[1][9] ));
 sg13g2_dfrbp_1 _3200_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net563),
    .D(net275),
    .Q_N(_1509_),
    .Q(\cic_a.temp_delay[1][10] ));
 sg13g2_dfrbp_1 _3201_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net563),
    .D(net282),
    .Q_N(_1508_),
    .Q(\cic_a.temp_delay[1][11] ));
 sg13g2_dfrbp_1 _3202_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net552),
    .D(net166),
    .Q_N(_1507_),
    .Q(\cic_a.temp_delay[1][12] ));
 sg13g2_dfrbp_1 _3203_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net596),
    .D(_0221_),
    .Q_N(_1506_),
    .Q(\cic_b.delay[2][0] ));
 sg13g2_dfrbp_1 _3204_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net595),
    .D(_0222_),
    .Q_N(_1505_),
    .Q(\cic_b.delay[2][1] ));
 sg13g2_dfrbp_1 _3205_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net595),
    .D(_0223_),
    .Q_N(_1504_),
    .Q(\cic_b.delay[2][2] ));
 sg13g2_dfrbp_1 _3206_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net597),
    .D(_0224_),
    .Q_N(_1503_),
    .Q(\cic_b.delay[2][3] ));
 sg13g2_dfrbp_1 _3207_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net597),
    .D(_0225_),
    .Q_N(_1502_),
    .Q(\cic_b.delay[2][4] ));
 sg13g2_dfrbp_1 _3208_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net587),
    .D(_0226_),
    .Q_N(_1501_),
    .Q(\cic_b.delay[2][5] ));
 sg13g2_dfrbp_1 _3209_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net587),
    .D(_0227_),
    .Q_N(_1500_),
    .Q(\cic_b.delay[2][6] ));
 sg13g2_dfrbp_1 _3210_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net587),
    .D(_0228_),
    .Q_N(_1499_),
    .Q(\cic_b.delay[2][7] ));
 sg13g2_dfrbp_1 _3211_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net589),
    .D(_0229_),
    .Q_N(_1498_),
    .Q(\cic_b.delay[2][8] ));
 sg13g2_dfrbp_1 _3212_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net589),
    .D(net38),
    .Q_N(_1497_),
    .Q(\cic_b.delay[2][9] ));
 sg13g2_dfrbp_1 _3213_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net562),
    .D(_0231_),
    .Q_N(_1496_),
    .Q(\cic_b.delay[2][10] ));
 sg13g2_dfrbp_1 _3214_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net560),
    .D(net317),
    .Q_N(_1495_),
    .Q(\cic_b.delay[2][11] ));
 sg13g2_dfrbp_1 _3215_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net561),
    .D(_0233_),
    .Q_N(_1494_),
    .Q(\cic_b.delay[2][12] ));
 sg13g2_dfrbp_1 _3216_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net594),
    .D(net643),
    .Q_N(_1493_),
    .Q(\cic_b.temp_comb[1][0] ));
 sg13g2_dfrbp_1 _3217_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net594),
    .D(net645),
    .Q_N(_1492_),
    .Q(\cic_b.temp_comb[1][1] ));
 sg13g2_dfrbp_1 _3218_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net594),
    .D(_0236_),
    .Q_N(_1491_),
    .Q(\cic_b.temp_comb[1][2] ));
 sg13g2_dfrbp_1 _3219_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net597),
    .D(net682),
    .Q_N(_1490_),
    .Q(\cic_b.temp_comb[1][3] ));
 sg13g2_dfrbp_1 _3220_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net587),
    .D(net641),
    .Q_N(_1489_),
    .Q(\cic_b.temp_comb[1][4] ));
 sg13g2_dfrbp_1 _3221_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net587),
    .D(_0239_),
    .Q_N(_1488_),
    .Q(\cic_b.temp_comb[1][5] ));
 sg13g2_dfrbp_1 _3222_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net587),
    .D(_0240_),
    .Q_N(_1487_),
    .Q(\cic_b.temp_comb[1][6] ));
 sg13g2_dfrbp_1 _3223_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net586),
    .D(_0241_),
    .Q_N(_1486_),
    .Q(\cic_b.temp_comb[1][7] ));
 sg13g2_dfrbp_1 _3224_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net586),
    .D(_0242_),
    .Q_N(_1485_),
    .Q(\cic_b.temp_comb[1][8] ));
 sg13g2_dfrbp_1 _3225_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net586),
    .D(_0243_),
    .Q_N(_1484_),
    .Q(\cic_b.temp_comb[1][9] ));
 sg13g2_dfrbp_1 _3226_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net560),
    .D(_0244_),
    .Q_N(_1483_),
    .Q(\cic_b.temp_comb[1][10] ));
 sg13g2_dfrbp_1 _3227_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net560),
    .D(_0245_),
    .Q_N(_1482_),
    .Q(\cic_b.temp_comb[1][11] ));
 sg13g2_dfrbp_1 _3228_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net561),
    .D(net462),
    .Q_N(_1481_),
    .Q(\cic_b.temp_comb[1][12] ));
 sg13g2_dfrbp_1 _3229_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net596),
    .D(_0247_),
    .Q_N(_1480_),
    .Q(\cic_b.delay[1][0] ));
 sg13g2_dfrbp_1 _3230_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net594),
    .D(_0248_),
    .Q_N(_1479_),
    .Q(\cic_b.delay[1][1] ));
 sg13g2_dfrbp_1 _3231_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net594),
    .D(_0249_),
    .Q_N(_1478_),
    .Q(\cic_b.delay[1][2] ));
 sg13g2_dfrbp_1 _3232_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net593),
    .D(_0250_),
    .Q_N(_1477_),
    .Q(\cic_b.delay[1][3] ));
 sg13g2_dfrbp_1 _3233_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net585),
    .D(net28),
    .Q_N(_1476_),
    .Q(\cic_b.delay[1][4] ));
 sg13g2_dfrbp_1 _3234_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net583),
    .D(_0252_),
    .Q_N(_1475_),
    .Q(\cic_b.delay[1][5] ));
 sg13g2_dfrbp_1 _3235_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net586),
    .D(_0253_),
    .Q_N(_1474_),
    .Q(\cic_b.delay[1][6] ));
 sg13g2_dfrbp_1 _3236_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net582),
    .D(_0254_),
    .Q_N(_1473_),
    .Q(\cic_b.delay[1][7] ));
 sg13g2_dfrbp_1 _3237_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net560),
    .D(_0255_),
    .Q_N(_1472_),
    .Q(\cic_b.delay[1][8] ));
 sg13g2_dfrbp_1 _3238_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net560),
    .D(net90),
    .Q_N(_1471_),
    .Q(\cic_b.delay[1][9] ));
 sg13g2_dfrbp_1 _3239_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net560),
    .D(net280),
    .Q_N(_1470_),
    .Q(\cic_b.delay[1][10] ));
 sg13g2_dfrbp_1 _3240_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net561),
    .D(net147),
    .Q_N(_1469_),
    .Q(\cic_b.delay[1][11] ));
 sg13g2_dfrbp_1 _3241_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net553),
    .D(net149),
    .Q_N(_1468_),
    .Q(\cic_b.delay[1][12] ));
 sg13g2_dfrbp_1 _3242_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net591),
    .D(_0260_),
    .Q_N(_1467_),
    .Q(\cic_b.delay[0][0] ));
 sg13g2_dfrbp_1 _3243_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net591),
    .D(net200),
    .Q_N(_1466_),
    .Q(\cic_b.delay[0][1] ));
 sg13g2_dfrbp_1 _3244_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net590),
    .D(_0262_),
    .Q_N(_1465_),
    .Q(\cic_b.delay[0][2] ));
 sg13g2_dfrbp_1 _3245_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net593),
    .D(_0263_),
    .Q_N(_1464_),
    .Q(\cic_b.delay[0][3] ));
 sg13g2_dfrbp_1 _3246_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net583),
    .D(_0264_),
    .Q_N(_1463_),
    .Q(\cic_b.delay[0][4] ));
 sg13g2_dfrbp_1 _3247_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net583),
    .D(net44),
    .Q_N(_1462_),
    .Q(\cic_b.delay[0][5] ));
 sg13g2_dfrbp_1 _3248_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net582),
    .D(_0266_),
    .Q_N(_1461_),
    .Q(\cic_b.delay[0][6] ));
 sg13g2_dfrbp_1 _3249_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net581),
    .D(_0267_),
    .Q_N(_1460_),
    .Q(\cic_b.delay[0][7] ));
 sg13g2_dfrbp_1 _3250_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net558),
    .D(_0268_),
    .Q_N(_1459_),
    .Q(\cic_b.delay[0][8] ));
 sg13g2_dfrbp_1 _3251_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net558),
    .D(net59),
    .Q_N(_1458_),
    .Q(\cic_b.delay[0][9] ));
 sg13g2_dfrbp_1 _3252_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net556),
    .D(_0270_),
    .Q_N(_1457_),
    .Q(\cic_b.delay[0][10] ));
 sg13g2_dfrbp_1 _3253_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net556),
    .D(net21),
    .Q_N(_1456_),
    .Q(\cic_b.delay[0][11] ));
 sg13g2_dfrbp_1 _3254_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net550),
    .D(net187),
    .Q_N(_1455_),
    .Q(\cic_b.delay[0][12] ));
 sg13g2_dfrbp_1 _3255_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net591),
    .D(net656),
    .Q_N(_1454_),
    .Q(\cic_b.temp_comb[0][0] ));
 sg13g2_dfrbp_1 _3256_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net592),
    .D(net637),
    .Q_N(_1453_),
    .Q(\cic_b.temp_comb[0][1] ));
 sg13g2_dfrbp_1 _3257_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net592),
    .D(net469),
    .Q_N(_1452_),
    .Q(\cic_b.temp_comb[0][2] ));
 sg13g2_dfrbp_1 _3258_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net593),
    .D(_0276_),
    .Q_N(_1451_),
    .Q(\cic_b.temp_comb[0][3] ));
 sg13g2_dfrbp_1 _3259_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net583),
    .D(_0277_),
    .Q_N(_1450_),
    .Q(\cic_b.temp_comb[0][4] ));
 sg13g2_dfrbp_1 _3260_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net583),
    .D(_0278_),
    .Q_N(_1449_),
    .Q(\cic_b.temp_comb[0][5] ));
 sg13g2_dfrbp_1 _3261_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net582),
    .D(_0279_),
    .Q_N(_1448_),
    .Q(\cic_b.temp_comb[0][6] ));
 sg13g2_dfrbp_1 _3262_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net582),
    .D(_0280_),
    .Q_N(_1447_),
    .Q(\cic_b.temp_comb[0][7] ));
 sg13g2_dfrbp_1 _3263_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net558),
    .D(_0281_),
    .Q_N(_1446_),
    .Q(\cic_b.temp_comb[0][8] ));
 sg13g2_dfrbp_1 _3264_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net558),
    .D(_0282_),
    .Q_N(_1445_),
    .Q(\cic_b.temp_comb[0][9] ));
 sg13g2_dfrbp_1 _3265_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net555),
    .D(_0283_),
    .Q_N(_1444_),
    .Q(\cic_b.temp_comb[0][10] ));
 sg13g2_dfrbp_1 _3266_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net555),
    .D(_0284_),
    .Q_N(_1443_),
    .Q(\cic_b.temp_comb[0][11] ));
 sg13g2_dfrbp_1 _3267_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net549),
    .D(_0285_),
    .Q_N(_1442_),
    .Q(\cic_b.temp_comb[0][12] ));
 sg13g2_dfrbp_1 _3268_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net611),
    .D(_0286_),
    .Q_N(_1441_),
    .Q(\cic_b.filtered_out[0] ));
 sg13g2_dfrbp_1 _3269_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net611),
    .D(_0287_),
    .Q_N(_1440_),
    .Q(\cic_b.filtered_out[1] ));
 sg13g2_dfrbp_1 _3270_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net611),
    .D(_0288_),
    .Q_N(_1439_),
    .Q(\cic_b.filtered_out[2] ));
 sg13g2_dfrbp_1 _3271_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net608),
    .D(_0289_),
    .Q_N(_1438_),
    .Q(\cic_b.filtered_out[3] ));
 sg13g2_dfrbp_1 _3272_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net601),
    .D(_0290_),
    .Q_N(_1437_),
    .Q(\cic_b.filtered_out[4] ));
 sg13g2_dfrbp_1 _3273_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net601),
    .D(net26),
    .Q_N(_1436_),
    .Q(\cic_b.filtered_out[5] ));
 sg13g2_dfrbp_1 _3274_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net601),
    .D(_0292_),
    .Q_N(_1435_),
    .Q(\cic_b.filtered_out[6] ));
 sg13g2_dfrbp_1 _3275_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net601),
    .D(_0293_),
    .Q_N(_1434_),
    .Q(\cic_b.filtered_out[7] ));
 sg13g2_dfrbp_1 _3276_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net599),
    .D(_0294_),
    .Q_N(_1433_),
    .Q(\cic_b.filtered_out[8] ));
 sg13g2_dfrbp_1 _3277_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net599),
    .D(_0295_),
    .Q_N(_1432_),
    .Q(\cic_b.filtered_out[9] ));
 sg13g2_dfrbp_1 _3278_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net599),
    .D(_0296_),
    .Q_N(_1431_),
    .Q(\cic_b.filtered_out[10] ));
 sg13g2_dfrbp_1 _3279_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net601),
    .D(_0297_),
    .Q_N(_1430_),
    .Q(\cic_b.filtered_out[11] ));
 sg13g2_dfrbp_1 _3280_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net609),
    .D(_0298_),
    .Q_N(_1429_),
    .Q(\cic_b.filtered_out[12] ));
 sg13g2_dfrbp_1 _3281_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net612),
    .D(net340),
    .Q_N(_1428_),
    .Q(\cic_b.temp_comb[2][0] ));
 sg13g2_dfrbp_1 _3282_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net612),
    .D(net170),
    .Q_N(_1427_),
    .Q(\cic_b.temp_comb[2][1] ));
 sg13g2_dfrbp_1 _3283_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net595),
    .D(_0301_),
    .Q_N(_1426_),
    .Q(\cic_b.temp_comb[2][2] ));
 sg13g2_dfrbp_1 _3284_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net597),
    .D(net124),
    .Q_N(_1425_),
    .Q(\cic_b.temp_comb[2][3] ));
 sg13g2_dfrbp_1 _3285_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net588),
    .D(net175),
    .Q_N(_1424_),
    .Q(\cic_b.temp_comb[2][4] ));
 sg13g2_dfrbp_1 _3286_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net588),
    .D(_0304_),
    .Q_N(_1423_),
    .Q(\cic_b.temp_comb[2][5] ));
 sg13g2_dfrbp_1 _3287_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net588),
    .D(net131),
    .Q_N(_1422_),
    .Q(\cic_b.temp_comb[2][6] ));
 sg13g2_dfrbp_1 _3288_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net588),
    .D(_0306_),
    .Q_N(_1421_),
    .Q(\cic_b.temp_comb[2][7] ));
 sg13g2_dfrbp_1 _3289_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net599),
    .D(net113),
    .Q_N(_1420_),
    .Q(\cic_b.temp_comb[2][8] ));
 sg13g2_dfrbp_1 _3290_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net599),
    .D(net195),
    .Q_N(_1419_),
    .Q(\cic_b.temp_comb[2][9] ));
 sg13g2_dfrbp_1 _3291_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net599),
    .D(_0309_),
    .Q_N(_1418_),
    .Q(\cic_b.temp_comb[2][10] ));
 sg13g2_dfrbp_1 _3292_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net586),
    .D(_0310_),
    .Q_N(_1417_),
    .Q(\cic_b.temp_comb[2][11] ));
 sg13g2_dfrbp_1 _3293_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net597),
    .D(_0311_),
    .Q_N(_1671_),
    .Q(\cic_b.temp_comb[2][12] ));
 sg13g2_dfrbp_1 _3294_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net591),
    .D(net453),
    .Q_N(_1672_),
    .Q(\cic_b.integrator[2][0] ));
 sg13g2_dfrbp_1 _3295_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net591),
    .D(net711),
    .Q_N(_1673_),
    .Q(\cic_b.integrator[2][1] ));
 sg13g2_dfrbp_1 _3296_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net590),
    .D(net761),
    .Q_N(_1674_),
    .Q(\cic_b.integrator[2][2] ));
 sg13g2_dfrbp_1 _3297_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net593),
    .D(_0093_),
    .Q_N(_1675_),
    .Q(\cic_b.integrator[2][3] ));
 sg13g2_dfrbp_1 _3298_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net584),
    .D(_0094_),
    .Q_N(_1676_),
    .Q(\cic_b.integrator[2][4] ));
 sg13g2_dfrbp_1 _3299_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net584),
    .D(net758),
    .Q_N(_1677_),
    .Q(\cic_b.integrator[2][5] ));
 sg13g2_dfrbp_1 _3300_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net581),
    .D(_0096_),
    .Q_N(_1678_),
    .Q(\cic_b.integrator[2][6] ));
 sg13g2_dfrbp_1 _3301_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net581),
    .D(net778),
    .Q_N(_1679_),
    .Q(\cic_b.integrator[2][7] ));
 sg13g2_dfrbp_1 _3302_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net557),
    .D(_0098_),
    .Q_N(_1680_),
    .Q(\cic_b.integrator[2][8] ));
 sg13g2_dfrbp_1 _3303_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net557),
    .D(_0099_),
    .Q_N(_1681_),
    .Q(\cic_b.integrator[2][9] ));
 sg13g2_dfrbp_1 _3304_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net555),
    .D(_0088_),
    .Q_N(_1682_),
    .Q(\cic_b.integrator[2][10] ));
 sg13g2_dfrbp_1 _3305_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net556),
    .D(_0089_),
    .Q_N(_1683_),
    .Q(\cic_b.integrator[2][11] ));
 sg13g2_dfrbp_1 _3306_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net549),
    .D(_0090_),
    .Q_N(_1684_),
    .Q(\cic_b.integrator[2][12] ));
 sg13g2_dfrbp_1 _3307_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net591),
    .D(_0074_),
    .Q_N(_1685_),
    .Q(\cic_b.integrator[1][0] ));
 sg13g2_dfrbp_1 _3308_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net590),
    .D(_0078_),
    .Q_N(_1686_),
    .Q(\cic_b.integrator[1][1] ));
 sg13g2_dfrbp_1 _3309_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net590),
    .D(_0079_),
    .Q_N(_1687_),
    .Q(\cic_b.integrator[1][2] ));
 sg13g2_dfrbp_1 _3310_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net593),
    .D(net719),
    .Q_N(_1688_),
    .Q(\cic_b.integrator[1][3] ));
 sg13g2_dfrbp_1 _3311_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net584),
    .D(net785),
    .Q_N(_1689_),
    .Q(\cic_b.integrator[1][4] ));
 sg13g2_dfrbp_1 _3312_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net584),
    .D(_0082_),
    .Q_N(_1690_),
    .Q(\cic_b.integrator[1][5] ));
 sg13g2_dfrbp_1 _3313_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net581),
    .D(net743),
    .Q_N(_1691_),
    .Q(\cic_b.integrator[1][6] ));
 sg13g2_dfrbp_1 _3314_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net581),
    .D(net780),
    .Q_N(_1692_),
    .Q(\cic_b.integrator[1][7] ));
 sg13g2_dfrbp_1 _3315_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net557),
    .D(_0085_),
    .Q_N(_1693_),
    .Q(\cic_b.integrator[1][8] ));
 sg13g2_dfrbp_1 _3316_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net557),
    .D(net739),
    .Q_N(_1694_),
    .Q(\cic_b.integrator[1][9] ));
 sg13g2_dfrbp_1 _3317_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net555),
    .D(_0075_),
    .Q_N(_1695_),
    .Q(\cic_b.integrator[1][10] ));
 sg13g2_dfrbp_1 _3318_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net555),
    .D(_0076_),
    .Q_N(_1696_),
    .Q(\cic_b.integrator[1][11] ));
 sg13g2_dfrbp_1 _3319_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net549),
    .D(net647),
    .Q_N(_1697_),
    .Q(\cic_b.integrator[1][12] ));
 sg13g2_dfrbp_1 _3320_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net590),
    .D(net93),
    .Q_N(_1698_),
    .Q(\cic_b.integrator[0][0] ));
 sg13g2_dfrbp_1 _3321_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net590),
    .D(_0065_),
    .Q_N(_1699_),
    .Q(\cic_b.integrator[0][1] ));
 sg13g2_dfrbp_1 _3322_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net590),
    .D(net438),
    .Q_N(_1700_),
    .Q(\cic_b.integrator[0][2] ));
 sg13g2_dfrbp_1 _3323_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net593),
    .D(_0067_),
    .Q_N(_1701_),
    .Q(\cic_b.integrator[0][3] ));
 sg13g2_dfrbp_1 _3324_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net584),
    .D(_0068_),
    .Q_N(_1702_),
    .Q(\cic_b.integrator[0][4] ));
 sg13g2_dfrbp_1 _3325_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net584),
    .D(net626),
    .Q_N(_1703_),
    .Q(\cic_b.integrator[0][5] ));
 sg13g2_dfrbp_1 _3326_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net581),
    .D(net691),
    .Q_N(_1704_),
    .Q(\cic_b.integrator[0][6] ));
 sg13g2_dfrbp_1 _3327_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net557),
    .D(net654),
    .Q_N(_1705_),
    .Q(\cic_b.integrator[0][7] ));
 sg13g2_dfrbp_1 _3328_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net557),
    .D(net728),
    .Q_N(_1706_),
    .Q(\cic_b.integrator[0][8] ));
 sg13g2_dfrbp_1 _3329_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net557),
    .D(net635),
    .Q_N(_1707_),
    .Q(\cic_b.integrator[0][9] ));
 sg13g2_dfrbp_1 _3330_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net555),
    .D(_0062_),
    .Q_N(_1708_),
    .Q(\cic_b.integrator[0][10] ));
 sg13g2_dfrbp_1 _3331_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net555),
    .D(_0063_),
    .Q_N(_1709_),
    .Q(\cic_b.integrator[0][11] ));
 sg13g2_dfrbp_1 _3332_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net555),
    .D(net185),
    .Q_N(_1416_),
    .Q(\cic_b.integrator[0][12] ));
 sg13g2_dfrbp_1 _3333_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net591),
    .D(net300),
    .Q_N(_1415_),
    .Q(\cic_b.temp_delay[0][0] ));
 sg13g2_dfrbp_1 _3334_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net592),
    .D(_0313_),
    .Q_N(_1414_),
    .Q(\cic_b.temp_delay[0][1] ));
 sg13g2_dfrbp_1 _3335_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net590),
    .D(net240),
    .Q_N(_1413_),
    .Q(\cic_b.temp_delay[0][2] ));
 sg13g2_dfrbp_1 _3336_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net593),
    .D(net298),
    .Q_N(_1412_),
    .Q(\cic_b.temp_delay[0][3] ));
 sg13g2_dfrbp_1 _3337_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net584),
    .D(net386),
    .Q_N(_1411_),
    .Q(\cic_b.temp_delay[0][4] ));
 sg13g2_dfrbp_1 _3338_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net583),
    .D(_0317_),
    .Q_N(_1410_),
    .Q(\cic_b.temp_delay[0][5] ));
 sg13g2_dfrbp_1 _3339_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net581),
    .D(net224),
    .Q_N(_1409_),
    .Q(\cic_b.temp_delay[0][6] ));
 sg13g2_dfrbp_1 _3340_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net581),
    .D(net302),
    .Q_N(_1408_),
    .Q(\cic_b.temp_delay[0][7] ));
 sg13g2_dfrbp_1 _3341_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net557),
    .D(net230),
    .Q_N(_1407_),
    .Q(\cic_b.temp_delay[0][8] ));
 sg13g2_dfrbp_1 _3342_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net558),
    .D(_0321_),
    .Q_N(_1406_),
    .Q(\cic_b.temp_delay[0][9] ));
 sg13g2_dfrbp_1 _3343_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net556),
    .D(net236),
    .Q_N(_1405_),
    .Q(\cic_b.temp_delay[0][10] ));
 sg13g2_dfrbp_1 _3344_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net556),
    .D(_0323_),
    .Q_N(_1404_),
    .Q(\cic_b.temp_delay[0][11] ));
 sg13g2_dfrbp_1 _3345_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net550),
    .D(_0324_),
    .Q_N(_1710_),
    .Q(\cic_b.temp_delay[0][12] ));
 sg13g2_dfrbp_1 _3346_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net548),
    .D(_0008_),
    .Q_N(_1711_),
    .Q(\cic_b.decim_cnt[0] ));
 sg13g2_dfrbp_1 _3347_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net548),
    .D(_0009_),
    .Q_N(_1712_),
    .Q(\cic_b.decim_cnt[1] ));
 sg13g2_dfrbp_1 _3348_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net548),
    .D(net62),
    .Q_N(_1713_),
    .Q(\cic_b.decim_cnt[2] ));
 sg13g2_dfrbp_1 _3349_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net549),
    .D(_0011_),
    .Q_N(_1714_),
    .Q(\cic_b.decim_cnt[3] ));
 sg13g2_dfrbp_1 _3350_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net549),
    .D(_0012_),
    .Q_N(_1715_),
    .Q(\cic_b.decim_cnt[4] ));
 sg13g2_dfrbp_1 _3351_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net549),
    .D(net335),
    .Q_N(_1716_),
    .Q(\cic_b.decim_cnt[5] ));
 sg13g2_dfrbp_1 _3352_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net549),
    .D(net193),
    .Q_N(_1717_),
    .Q(\cic_b.decim_cnt[6] ));
 sg13g2_dfrbp_1 _3353_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net549),
    .D(net70),
    .Q_N(_1403_),
    .Q(\cic_b.decim_cnt[7] ));
 sg13g2_dfrbp_1 _3354_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net605),
    .D(net160),
    .Q_N(_1402_),
    .Q(\cic_a.temp_delay[2][0] ));
 sg13g2_dfrbp_1 _3355_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net605),
    .D(net154),
    .Q_N(_1401_),
    .Q(\cic_a.temp_delay[2][1] ));
 sg13g2_dfrbp_1 _3356_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net603),
    .D(net122),
    .Q_N(_1400_),
    .Q(\cic_a.temp_delay[2][2] ));
 sg13g2_dfrbp_1 _3357_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net577),
    .D(net213),
    .Q_N(_1399_),
    .Q(\cic_a.temp_delay[2][3] ));
 sg13g2_dfrbp_1 _3358_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net575),
    .D(net164),
    .Q_N(_1398_),
    .Q(\cic_a.temp_delay[2][4] ));
 sg13g2_dfrbp_1 _3359_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net576),
    .D(_0330_),
    .Q_N(_1397_),
    .Q(\cic_a.temp_delay[2][5] ));
 sg13g2_dfrbp_1 _3360_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net575),
    .D(net396),
    .Q_N(_1396_),
    .Q(\cic_a.temp_delay[2][6] ));
 sg13g2_dfrbp_1 _3361_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net570),
    .D(net263),
    .Q_N(_1395_),
    .Q(\cic_a.temp_delay[2][7] ));
 sg13g2_dfrbp_1 _3362_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net575),
    .D(_0333_),
    .Q_N(_1394_),
    .Q(\cic_a.temp_delay[2][8] ));
 sg13g2_dfrbp_1 _3363_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net569),
    .D(net290),
    .Q_N(_1393_),
    .Q(\cic_a.temp_delay[2][9] ));
 sg13g2_dfrbp_1 _3364_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net573),
    .D(_0335_),
    .Q_N(_1392_),
    .Q(\cic_a.temp_delay[2][10] ));
 sg13g2_dfrbp_1 _3365_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net572),
    .D(net288),
    .Q_N(_1391_),
    .Q(\cic_a.temp_delay[2][11] ));
 sg13g2_dfrbp_1 _3366_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net572),
    .D(net222),
    .Q_N(_1390_),
    .Q(\cic_a.temp_delay[2][12] ));
 sg13g2_dfrbp_1 _3367_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net594),
    .D(net206),
    .Q_N(_1389_),
    .Q(\cic_b.temp_delay[1][0] ));
 sg13g2_dfrbp_1 _3368_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net594),
    .D(net337),
    .Q_N(_1388_),
    .Q(\cic_b.temp_delay[1][1] ));
 sg13g2_dfrbp_1 _3369_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net592),
    .D(net183),
    .Q_N(_1387_),
    .Q(\cic_b.temp_delay[1][2] ));
 sg13g2_dfrbp_1 _3370_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net593),
    .D(net269),
    .Q_N(_1386_),
    .Q(\cic_b.temp_delay[1][3] ));
 sg13g2_dfrbp_1 _3371_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net583),
    .D(_0342_),
    .Q_N(_1385_),
    .Q(\cic_b.temp_delay[1][4] ));
 sg13g2_dfrbp_1 _3372_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net583),
    .D(net305),
    .Q_N(_1384_),
    .Q(\cic_b.temp_delay[1][5] ));
 sg13g2_dfrbp_1 _3373_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net586),
    .D(net331),
    .Q_N(_1383_),
    .Q(\cic_b.temp_delay[1][6] ));
 sg13g2_dfrbp_1 _3374_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net582),
    .D(net234),
    .Q_N(_1382_),
    .Q(\cic_b.temp_delay[1][7] ));
 sg13g2_dfrbp_1 _3375_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net558),
    .D(net180),
    .Q_N(_1381_),
    .Q(\cic_b.temp_delay[1][8] ));
 sg13g2_dfrbp_1 _3376_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net558),
    .D(_0347_),
    .Q_N(_1380_),
    .Q(\cic_b.temp_delay[1][9] ));
 sg13g2_dfrbp_1 _3377_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net560),
    .D(_0348_),
    .Q_N(_1379_),
    .Q(\cic_b.temp_delay[1][10] ));
 sg13g2_dfrbp_1 _3378_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net561),
    .D(_0349_),
    .Q_N(_1378_),
    .Q(\cic_b.temp_delay[1][11] ));
 sg13g2_dfrbp_1 _3379_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net553),
    .D(_0350_),
    .Q_N(_1377_),
    .Q(\cic_b.temp_delay[1][12] ));
 sg13g2_dfrbp_1 _3380_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net616),
    .D(_0351_),
    .Q_N(_1376_),
    .Q(\serializer_a.shift_reg[0] ));
 sg13g2_dfrbp_1 _3381_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net616),
    .D(_0352_),
    .Q_N(_1375_),
    .Q(\serializer_a.shift_reg[1] ));
 sg13g2_dfrbp_1 _3382_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net613),
    .D(_0353_),
    .Q_N(_1374_),
    .Q(\serializer_a.shift_reg[2] ));
 sg13g2_dfrbp_1 _3383_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net613),
    .D(net88),
    .Q_N(_1373_),
    .Q(\serializer_a.shift_reg[3] ));
 sg13g2_dfrbp_1 _3384_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net613),
    .D(_0355_),
    .Q_N(_1372_),
    .Q(\serializer_a.shift_reg[4] ));
 sg13g2_dfrbp_1 _3385_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net613),
    .D(net47),
    .Q_N(_1371_),
    .Q(\serializer_a.shift_reg[5] ));
 sg13g2_dfrbp_1 _3386_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net614),
    .D(_0357_),
    .Q_N(_1370_),
    .Q(\serializer_a.shift_reg[6] ));
 sg13g2_dfrbp_1 _3387_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net614),
    .D(_0358_),
    .Q_N(_1369_),
    .Q(\serializer_a.shift_reg[7] ));
 sg13g2_dfrbp_1 _3388_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net614),
    .D(net211),
    .Q_N(_1368_),
    .Q(\serializer_a.shift_reg[8] ));
 sg13g2_dfrbp_1 _3389_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net610),
    .D(net261),
    .Q_N(_1367_),
    .Q(\serializer_a.shift_reg[9] ));
 sg13g2_dfrbp_1 _3390_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net610),
    .D(net204),
    .Q_N(_1366_),
    .Q(\serializer_a.shift_reg[10] ));
 sg13g2_dfrbp_1 _3391_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net612),
    .D(net208),
    .Q_N(_1365_),
    .Q(\serializer_a.shift_reg[11] ));
 sg13g2_dfrbp_1 _3392_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net611),
    .D(net126),
    .Q_N(_1718_),
    .Q(\serializer_a.serial_out ));
 sg13g2_dfrbp_1 _3393_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net616),
    .D(_0016_),
    .Q_N(_1364_),
    .Q(\serializer_a.sending ));
 sg13g2_dfrbp_1 _3394_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net595),
    .D(net202),
    .Q_N(_1363_),
    .Q(\cic_b.temp_delay[2][0] ));
 sg13g2_dfrbp_1 _3395_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net595),
    .D(net320),
    .Q_N(_1362_),
    .Q(\cic_b.temp_delay[2][1] ));
 sg13g2_dfrbp_1 _3396_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net594),
    .D(net220),
    .Q_N(_1361_),
    .Q(\cic_b.temp_delay[2][2] ));
 sg13g2_dfrbp_1 _3397_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net597),
    .D(net249),
    .Q_N(_1360_),
    .Q(\cic_b.temp_delay[2][3] ));
 sg13g2_dfrbp_1 _3398_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net597),
    .D(net273),
    .Q_N(_1359_),
    .Q(\cic_b.temp_delay[2][4] ));
 sg13g2_dfrbp_1 _3399_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net587),
    .D(net267),
    .Q_N(_1358_),
    .Q(\cic_b.temp_delay[2][5] ));
 sg13g2_dfrbp_1 _3400_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net587),
    .D(net257),
    .Q_N(_1357_),
    .Q(\cic_b.temp_delay[2][6] ));
 sg13g2_dfrbp_1 _3401_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net586),
    .D(net367),
    .Q_N(_1356_),
    .Q(\cic_b.temp_delay[2][7] ));
 sg13g2_dfrbp_1 _3402_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net589),
    .D(net323),
    .Q_N(_1355_),
    .Q(\cic_b.temp_delay[2][8] ));
 sg13g2_dfrbp_1 _3403_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net586),
    .D(_0373_),
    .Q_N(_1354_),
    .Q(\cic_b.temp_delay[2][9] ));
 sg13g2_dfrbp_1 _3404_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net562),
    .D(net242),
    .Q_N(_1353_),
    .Q(\cic_b.temp_delay[2][10] ));
 sg13g2_dfrbp_1 _3405_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net560),
    .D(_0375_),
    .Q_N(_1352_),
    .Q(\cic_b.temp_delay[2][11] ));
 sg13g2_dfrbp_1 _3406_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net561),
    .D(net343),
    .Q_N(_1719_),
    .Q(\cic_b.temp_delay[2][12] ));
 sg13g2_dfrbp_1 _3407_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net611),
    .D(net539),
    .Q_N(_1351_),
    .Q(\serializer_a.valid ));
 sg13g2_dfrbp_1 _3408_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net611),
    .D(_0377_),
    .Q_N(_1350_),
    .Q(\serializer_b.shift_reg[0] ));
 sg13g2_dfrbp_1 _3409_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net611),
    .D(net75),
    .Q_N(_1349_),
    .Q(\serializer_b.shift_reg[1] ));
 sg13g2_dfrbp_1 _3410_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net609),
    .D(_0379_),
    .Q_N(_1348_),
    .Q(\serializer_b.shift_reg[2] ));
 sg13g2_dfrbp_1 _3411_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net608),
    .D(net85),
    .Q_N(_1347_),
    .Q(\serializer_b.shift_reg[3] ));
 sg13g2_dfrbp_1 _3412_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net610),
    .D(net80),
    .Q_N(_1346_),
    .Q(\serializer_b.shift_reg[4] ));
 sg13g2_dfrbp_1 _3413_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net610),
    .D(net67),
    .Q_N(_1345_),
    .Q(\serializer_b.shift_reg[5] ));
 sg13g2_dfrbp_1 _3414_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net601),
    .D(net259),
    .Q_N(_1344_),
    .Q(\serializer_b.shift_reg[6] ));
 sg13g2_dfrbp_1 _3415_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net601),
    .D(net278),
    .Q_N(_1343_),
    .Q(\serializer_b.shift_reg[7] ));
 sg13g2_dfrbp_1 _3416_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net601),
    .D(net136),
    .Q_N(_1342_),
    .Q(\serializer_b.shift_reg[8] ));
 sg13g2_dfrbp_1 _3417_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net609),
    .D(net178),
    .Q_N(_1341_),
    .Q(\serializer_b.shift_reg[9] ));
 sg13g2_dfrbp_1 _3418_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net609),
    .D(_0387_),
    .Q_N(_1340_),
    .Q(\serializer_b.shift_reg[10] ));
 sg13g2_dfrbp_1 _3419_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net608),
    .D(_0388_),
    .Q_N(_1339_),
    .Q(\serializer_b.shift_reg[11] ));
 sg13g2_dfrbp_1 _3420_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net611),
    .D(net105),
    .Q_N(_1720_),
    .Q(\serializer_b.serial_out ));
 sg13g2_dfrbp_1 _3421_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net608),
    .D(_0020_),
    .Q_N(_1338_),
    .Q(\serializer_b.sending ));
 sg13g2_dfrbp_1 _3422_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net615),
    .D(_0390_),
    .Q_N(_1337_),
    .Q(\serializer_ab_subtr.bit_cnt[0] ));
 sg13g2_dfrbp_1 _3423_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net615),
    .D(net107),
    .Q_N(_1336_),
    .Q(\serializer_ab_subtr.bit_cnt[1] ));
 sg13g2_dfrbp_1 _3424_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net615),
    .D(_0392_),
    .Q_N(_1335_),
    .Q(\serializer_ab_subtr.bit_cnt[2] ));
 sg13g2_dfrbp_1 _3425_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net615),
    .D(net82),
    .Q_N(_1721_),
    .Q(\serializer_ab_subtr.bit_cnt[3] ));
 sg13g2_dfrbp_1 _3426_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net595),
    .D(net535),
    .Q_N(_1334_),
    .Q(\serializer_b.valid ));
 sg13g2_dfrbp_1 _3427_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net608),
    .D(net109),
    .Q_N(_1333_),
    .Q(\serializer_b.bit_cnt[0] ));
 sg13g2_dfrbp_1 _3428_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net608),
    .D(_0395_),
    .Q_N(_1332_),
    .Q(\serializer_b.bit_cnt[1] ));
 sg13g2_dfrbp_1 _3429_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net608),
    .D(_0396_),
    .Q_N(_1331_),
    .Q(\serializer_b.bit_cnt[2] ));
 sg13g2_dfrbp_1 _3430_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net608),
    .D(net64),
    .Q_N(_1330_),
    .Q(\serializer_b.bit_cnt[3] ));
 sg13g2_dfrbp_1 _3431_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net615),
    .D(net427),
    .Q_N(_1329_),
    .Q(\serializer_ab_subtr.shift_reg[0] ));
 sg13g2_dfrbp_1 _3432_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net615),
    .D(net215),
    .Q_N(_1328_),
    .Q(\serializer_ab_subtr.shift_reg[1] ));
 sg13g2_dfrbp_1 _3433_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net615),
    .D(net420),
    .Q_N(_1327_),
    .Q(\serializer_ab_subtr.shift_reg[2] ));
 sg13g2_dfrbp_1 _3434_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net614),
    .D(_0401_),
    .Q_N(_1326_),
    .Q(\serializer_ab_subtr.shift_reg[3] ));
 sg13g2_dfrbp_1 _3435_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net614),
    .D(_0402_),
    .Q_N(_1325_),
    .Q(\serializer_ab_subtr.shift_reg[4] ));
 sg13g2_dfrbp_1 _3436_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net614),
    .D(net379),
    .Q_N(_1324_),
    .Q(\serializer_ab_subtr.shift_reg[5] ));
 sg13g2_dfrbp_1 _3437_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net614),
    .D(_0404_),
    .Q_N(_1323_),
    .Q(\serializer_ab_subtr.shift_reg[6] ));
 sg13g2_dfrbp_1 _3438_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net614),
    .D(_0405_),
    .Q_N(_1322_),
    .Q(\serializer_ab_subtr.shift_reg[7] ));
 sg13g2_dfrbp_1 _3439_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net610),
    .D(_0406_),
    .Q_N(_1321_),
    .Q(\serializer_ab_subtr.shift_reg[8] ));
 sg13g2_dfrbp_1 _3440_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net610),
    .D(_0407_),
    .Q_N(_1320_),
    .Q(\serializer_ab_subtr.shift_reg[9] ));
 sg13g2_dfrbp_1 _3441_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net610),
    .D(_0408_),
    .Q_N(_1319_),
    .Q(\serializer_ab_subtr.shift_reg[10] ));
 sg13g2_dfrbp_1 _3442_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net612),
    .D(_0409_),
    .Q_N(_1318_),
    .Q(\serializer_ab_subtr.shift_reg[11] ));
 sg13g2_dfrbp_1 _3443_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net612),
    .D(net401),
    .Q_N(_1722_),
    .Q(\serializer_ab_subtr.serial_out ));
 sg13g2_dfrbp_1 _3444_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net615),
    .D(_0018_),
    .Q_N(_1317_),
    .Q(\serializer_ab_subtr.sending ));
 sg13g2_dfrbp_1 _3445_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net616),
    .D(_0411_),
    .Q_N(_1316_),
    .Q(\serializer_a.bit_cnt[0] ));
 sg13g2_dfrbp_1 _3446_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net616),
    .D(net152),
    .Q_N(_1315_),
    .Q(\serializer_a.bit_cnt[1] ));
 sg13g2_dfrbp_1 _3447_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net616),
    .D(_0413_),
    .Q_N(_1314_),
    .Q(\serializer_a.bit_cnt[2] ));
 sg13g2_dfrbp_1 _3448_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net616),
    .D(net49),
    .Q_N(_1723_),
    .Q(\serializer_a.bit_cnt[3] ));
 sg13g2_dfrbp_1 _3449_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net595),
    .D(_0019_),
    .Q_N(_1313_),
    .Q(\serializer_ab_subtr.valid ));
 sg13g2_tielo tt_um_ds_comp_adc_5 (.L_LO(net5));
 sg13g2_tielo tt_um_ds_comp_adc_6 (.L_LO(net6));
 sg13g2_tielo tt_um_ds_comp_adc_7 (.L_LO(net7));
 sg13g2_tielo tt_um_ds_comp_adc_8 (.L_LO(net8));
 sg13g2_tielo tt_um_ds_comp_adc_9 (.L_LO(net9));
 sg13g2_tielo tt_um_ds_comp_adc_10 (.L_LO(net10));
 sg13g2_tielo tt_um_ds_comp_adc_11 (.L_LO(net11));
 sg13g2_tielo tt_um_ds_comp_adc_12 (.L_LO(net12));
 sg13g2_tielo tt_um_ds_comp_adc_13 (.L_LO(net13));
 sg13g2_tielo tt_um_ds_comp_adc_14 (.L_LO(net14));
 sg13g2_tielo tt_um_ds_comp_adc_15 (.L_LO(net15));
 sg13g2_tielo tt_um_ds_comp_adc_16 (.L_LO(net16));
 sg13g2_tielo tt_um_ds_comp_adc_17 (.L_LO(net17));
 sg13g2_tielo tt_um_ds_comp_adc_18 (.L_LO(net18));
 sg13g2_tielo tt_um_ds_comp_adc_19 (.L_LO(net19));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_2 _3466_ (.A(pdm_a),
    .X(uo_out[0]));
 sg13g2_buf_2 _3467_ (.A(pdm_b),
    .X(uo_out[1]));
 sg13g2_buf_2 _3468_ (.A(\serializer_a.serial_out ),
    .X(uo_out[2]));
 sg13g2_buf_1 _3469_ (.A(\serializer_b.serial_out ),
    .X(uo_out[3]));
 sg13g2_buf_1 _3470_ (.A(\serializer_ab_subtr.serial_out ),
    .X(uo_out[4]));
 sg13g2_buf_1 _3471_ (.A(\serializer_a.valid ),
    .X(uo_out[5]));
 sg13g2_buf_1 _3472_ (.A(\serializer_b.valid ),
    .X(uo_out[6]));
 sg13g2_buf_1 _3473_ (.A(\serializer_ab_subtr.valid ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout471 (.X(net471),
    .A(net472));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(net473));
 sg13g2_buf_2 fanout473 (.A(net481),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_4 fanout476 (.X(net476),
    .A(net481));
 sg13g2_buf_2 fanout477 (.A(net479),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(net479),
    .X(net478));
 sg13g2_buf_1 fanout479 (.A(net481),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(net481),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_1249_),
    .X(net481));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(net483));
 sg13g2_buf_2 fanout483 (.A(net486),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(net486),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(net490),
    .X(net486));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(net488));
 sg13g2_buf_4 fanout488 (.X(net488),
    .A(net489));
 sg13g2_buf_4 fanout489 (.X(net489),
    .A(net490));
 sg13g2_buf_2 fanout490 (.A(_1249_),
    .X(net490));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net499));
 sg13g2_buf_1 fanout492 (.A(net493),
    .X(net492));
 sg13g2_buf_4 fanout493 (.X(net493),
    .A(net499));
 sg13g2_buf_2 fanout494 (.A(net499),
    .X(net494));
 sg13g2_buf_4 fanout495 (.X(net495),
    .A(net497));
 sg13g2_buf_1 fanout496 (.A(net497),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(net499),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_1249_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net502),
    .X(net500));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(net502));
 sg13g2_buf_2 fanout502 (.A(net503),
    .X(net502));
 sg13g2_buf_4 fanout503 (.X(net503),
    .A(net504));
 sg13g2_buf_2 fanout504 (.A(net528),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(net511),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(net511),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(net508),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net511),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_4 fanout510 (.X(net510),
    .A(net511));
 sg13g2_buf_2 fanout511 (.A(net516),
    .X(net511));
 sg13g2_buf_4 fanout512 (.X(net512),
    .A(net513));
 sg13g2_buf_2 fanout513 (.A(net516),
    .X(net513));
 sg13g2_buf_4 fanout514 (.X(net514),
    .A(net516));
 sg13g2_buf_2 fanout515 (.A(net516),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(net528),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(net518),
    .X(net517));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(net527));
 sg13g2_buf_2 fanout519 (.A(net522),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(net522),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(net522),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(net527),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(net524),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(net525),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(net526),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(net527),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_4 fanout528 (.X(net528),
    .A(_1239_));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(_0591_));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(_0587_));
 sg13g2_buf_1 fanout531 (.A(_0587_),
    .X(net531));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(_0594_));
 sg13g2_buf_2 fanout533 (.A(_0594_),
    .X(net533));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(net535));
 sg13g2_buf_2 fanout535 (.A(_0021_),
    .X(net535));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(_1234_));
 sg13g2_buf_1 fanout537 (.A(_1234_),
    .X(net537));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(net539));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(_0017_));
 sg13g2_buf_2 fanout540 (.A(net542),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(\serializer_ab_subtr.sending ),
    .X(net541));
 sg13g2_buf_1 fanout542 (.A(\serializer_ab_subtr.sending ),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(\serializer_b.sending ),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(\serializer_b.sending ),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(net547),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(\serializer_a.sending ),
    .X(net547));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(net550));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(net550));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(net580));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(net552));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(net554));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(net554));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(net580));
 sg13g2_buf_4 fanout555 (.X(net555),
    .A(net559));
 sg13g2_buf_2 fanout556 (.A(net559),
    .X(net556));
 sg13g2_buf_4 fanout557 (.X(net557),
    .A(net559));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(net559));
 sg13g2_buf_2 fanout559 (.A(net562),
    .X(net559));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(net562));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(net562));
 sg13g2_buf_2 fanout562 (.A(net580),
    .X(net562));
 sg13g2_buf_4 fanout563 (.X(net563),
    .A(net564));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(net571));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(net571));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(net571));
 sg13g2_buf_4 fanout567 (.X(net567),
    .A(net568));
 sg13g2_buf_2 fanout568 (.A(net571),
    .X(net568));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(net571));
 sg13g2_buf_2 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(net580),
    .X(net571));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(net574));
 sg13g2_buf_2 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(net579));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(net578));
 sg13g2_buf_2 fanout576 (.A(net578),
    .X(net576));
 sg13g2_buf_4 fanout577 (.X(net577),
    .A(net578));
 sg13g2_buf_2 fanout578 (.A(net579),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_4 fanout580 (.X(net580),
    .A(rst_n));
 sg13g2_buf_4 fanout581 (.X(net581),
    .A(net585));
 sg13g2_buf_2 fanout582 (.A(net585),
    .X(net582));
 sg13g2_buf_4 fanout583 (.X(net583),
    .A(net584));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(net585));
 sg13g2_buf_2 fanout585 (.A(net619),
    .X(net585));
 sg13g2_buf_4 fanout586 (.X(net586),
    .A(net589));
 sg13g2_buf_4 fanout587 (.X(net587),
    .A(net589));
 sg13g2_buf_2 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_4 fanout589 (.X(net589),
    .A(net619));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(net591));
 sg13g2_buf_4 fanout591 (.X(net591),
    .A(net598));
 sg13g2_buf_2 fanout592 (.A(net598),
    .X(net592));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(net598));
 sg13g2_buf_4 fanout594 (.X(net594),
    .A(net596));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(net596));
 sg13g2_buf_2 fanout596 (.A(net597),
    .X(net596));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(net598));
 sg13g2_buf_2 fanout598 (.A(net619),
    .X(net598));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(net602));
 sg13g2_buf_4 fanout600 (.X(net600),
    .A(net602));
 sg13g2_buf_4 fanout601 (.X(net601),
    .A(net602));
 sg13g2_buf_2 fanout602 (.A(net618),
    .X(net602));
 sg13g2_buf_4 fanout603 (.X(net603),
    .A(net607));
 sg13g2_buf_4 fanout604 (.X(net604),
    .A(net607));
 sg13g2_buf_4 fanout605 (.X(net605),
    .A(net606));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(net607));
 sg13g2_buf_2 fanout607 (.A(net618),
    .X(net607));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(net609));
 sg13g2_buf_2 fanout609 (.A(net610),
    .X(net609));
 sg13g2_buf_4 fanout610 (.X(net610),
    .A(net618));
 sg13g2_buf_8 fanout611 (.A(net612),
    .X(net611));
 sg13g2_buf_8 fanout612 (.A(net618),
    .X(net612));
 sg13g2_buf_4 fanout613 (.X(net613),
    .A(net617));
 sg13g2_buf_4 fanout614 (.X(net614),
    .A(net617));
 sg13g2_buf_4 fanout615 (.X(net615),
    .A(net617));
 sg13g2_buf_4 fanout616 (.X(net616),
    .A(net617));
 sg13g2_buf_2 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(net619),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(rst_n),
    .X(net619));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[7]),
    .X(net3));
 sg13g2_tielo tt_um_ds_comp_adc_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload2 (.A(clknet_leaf_52_clk));
 sg13g2_inv_4 clkload3 (.A(clknet_leaf_53_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_leaf_4_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_46_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_39_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_41_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_33_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_34_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_9_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_18_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\cic_b.temp_delay[0][11] ),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0271_),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold3 (.A(\cic_a.temp_delay[0][5] ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0148_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cic_b.decim_cnt[0] ),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold6 (.A(\cic_b.temp_comb[2][5] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0291_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold8 (.A(\cic_b.temp_delay[1][4] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0251_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cic_a.decim_cnt[0] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cic_a.decim_cnt[2] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold12 (.A(_1236_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0002_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold14 (.A(\serializer_b.shift_reg[0] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold15 (.A(_1074_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold16 (.A(\serializer_a.shift_reg[0] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold17 (.A(_1057_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold18 (.A(\cic_b.temp_delay[2][9] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0230_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold20 (.A(\cic_a.pdm_in ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0022_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold22 (.A(\cic_a.temp_delay[0][7] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0150_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cic_b.temp_delay[0][5] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0265_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold26 (.A(\serializer_a.shift_reg[4] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold27 (.A(_1063_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0356_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold29 (.A(\serializer_a.bit_cnt[3] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0414_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cic_a.temp_delay[1][9] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0139_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold33 (.A(\serializer_a.bit_cnt[2] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold34 (.A(_1188_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold35 (.A(\cic_a.temp_delay[0][10] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0153_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold37 (.A(\cic_a.decim_cnt[7] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0007_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold39 (.A(\cic_b.temp_delay[0][9] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0269_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold41 (.A(\cic_b.decim_cnt[2] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold42 (.A(_1246_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0010_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold44 (.A(\serializer_b.bit_cnt[3] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0397_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold46 (.A(\serializer_b.shift_reg[4] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold47 (.A(_1082_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0382_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold49 (.A(\cic_a.decim_cnt[1] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold50 (.A(\cic_b.decim_cnt[7] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0015_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold52 (.A(\cic_a.temp_delay[2][8] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0112_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold54 (.A(\serializer_b.shift_reg[1] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold55 (.A(_1076_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0378_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold57 (.A(\serializer_b.bit_cnt[2] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold58 (.A(_1104_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold59 (.A(\serializer_b.shift_reg[3] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold60 (.A(_1080_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0381_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold62 (.A(\serializer_ab_subtr.bit_cnt[3] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0393_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold64 (.A(\serializer_b.shift_reg[2] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold65 (.A(_1078_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0380_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold67 (.A(\serializer_a.shift_reg[2] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold68 (.A(_1060_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0354_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold70 (.A(\cic_b.temp_delay[1][9] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0256_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold72 (.A(\serializer_ab_subtr.bit_cnt[0] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cic_b.pdm_in ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0061_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cic_a.temp_comb[2][7] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0176_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold77 (.A(\serializer_ab_subtr.bit_cnt[2] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold78 (.A(_1097_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold79 (.A(\cic_a.temp_delay[0][9] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0204_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold81 (.A(\cic_a.integrator[0][12] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0025_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold83 (.A(\cic_b.integrator[2][5] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold84 (.A(\serializer_b.shift_reg[11] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold85 (.A(_1090_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0389_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold87 (.A(\serializer_ab_subtr.bit_cnt[1] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0391_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold89 (.A(\serializer_b.bit_cnt[0] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0394_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold91 (.A(\cic_a.temp_delay[0][2] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0145_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cic_b.temp_comb[2][8] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0307_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cic_a.temp_comb[2][1] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0183_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cic_b.decim_cnt[1] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold98 (.A(\serializer_a.shift_reg[1] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold99 (.A(_1059_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cic_a.temp_comb[2][0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0182_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cic_a.temp_delay[2][2] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0327_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cic_b.temp_comb[2][3] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0302_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold106 (.A(\serializer_a.serial_out ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0363_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cic_b.integrator[2][11] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cic_a.temp_delay[1][0] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0208_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold111 (.A(\cic_b.temp_comb[2][6] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0305_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold113 (.A(\cic_a.temp_comb[2][3] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold114 (.A(\serializer_b.shift_reg[10] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold115 (.A(_1089_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold116 (.A(\serializer_b.shift_reg[8] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0385_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cic_a.delay[2][6] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold119 (.A(\cic_b.integrator[2][9] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cic_a.temp_delay[1][6] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0136_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cic_a.temp_delay[0][3] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0146_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cic_b.temp_comb[0][4] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cic_a.integrator[2][3] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cic_a.temp_comb[0][9] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold127 (.A(\cic_b.temp_delay[1][11] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0258_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold129 (.A(\cic_b.temp_delay[1][12] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0259_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold131 (.A(\cic_b.filtered_out[2] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold132 (.A(\serializer_a.bit_cnt[1] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0412_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cic_a.temp_delay[2][1] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0326_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold136 (.A(\serializer_a.bit_cnt[0] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold137 (.A(\cic_a.temp_delay[1][3] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0211_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold139 (.A(\cic_a.integrator[2][5] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cic_a.temp_delay[2][0] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0325_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cic_b.delay[2][4] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cic_b.temp_comb[1][9] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cic_a.temp_delay[2][4] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0329_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold146 (.A(\cic_a.temp_delay[1][12] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0220_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold148 (.A(\cic_a.temp_delay[1][2] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0210_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold150 (.A(\cic_b.temp_comb[2][1] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0300_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cic_a.temp_comb[0][6] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold153 (.A(\serializer_a.shift_reg[3] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold154 (.A(_1062_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cic_b.temp_comb[2][4] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0303_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold157 (.A(\cic_b.temp_comb[2][7] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold158 (.A(\serializer_b.shift_reg[9] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0386_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold160 (.A(\cic_b.temp_delay[1][8] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0346_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold162 (.A(\cic_a.delay[2][2] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold163 (.A(\cic_b.temp_delay[1][2] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0340_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold165 (.A(\cic_b.integrator[0][12] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0064_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold167 (.A(\cic_b.temp_delay[0][12] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0272_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cic_a.integrator[2][2] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold170 (.A(\cic_a.temp_delay[0][8] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0203_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold172 (.A(\cic_a.temp_comb[2][11] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cic_b.decim_cnt[6] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0014_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold175 (.A(\cic_b.temp_comb[2][9] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0308_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold177 (.A(\cic_a.delay[1][0] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold178 (.A(\cic_a.temp_delay[0][0] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0195_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cic_b.temp_delay[0][1] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0261_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cic_b.temp_delay[2][0] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0364_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold184 (.A(\serializer_a.shift_reg[10] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0361_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold186 (.A(\cic_b.temp_delay[1][0] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0338_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold188 (.A(\serializer_a.shift_reg[11] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0362_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold190 (.A(\serializer_a.shift_reg[7] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold191 (.A(_1067_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0359_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold193 (.A(\cic_a.temp_delay[2][3] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0328_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold195 (.A(\serializer_ab_subtr.shift_reg[1] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0399_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold197 (.A(\cic_b.delay[2][0] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold198 (.A(\cic_a.delay[0][8] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold199 (.A(\cic_b.temp_comb[0][11] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold200 (.A(\cic_b.temp_delay[2][2] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0366_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold202 (.A(\cic_a.temp_delay[2][12] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0337_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold204 (.A(\cic_b.temp_delay[0][6] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0318_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold206 (.A(\cic_a.temp_delay[1][5] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0213_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold208 (.A(\cic_a.temp_delay[0][11] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0206_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold210 (.A(\cic_b.temp_delay[0][8] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0320_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold212 (.A(\cic_a.temp_comb[2][5] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold213 (.A(\serializer_b.bit_cnt[1] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold214 (.A(\cic_b.temp_delay[1][7] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0345_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold216 (.A(\cic_b.temp_delay[0][10] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0322_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold218 (.A(\cic_a.temp_delay[0][1] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0196_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold220 (.A(\cic_b.temp_delay[0][2] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0314_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold222 (.A(\cic_b.temp_delay[2][10] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0374_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold224 (.A(\cic_a.delay[1][3] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold225 (.A(\cic_a.decim_cnt[6] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0006_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold227 (.A(\cic_a.temp_delay[2][10] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0114_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold229 (.A(\cic_b.temp_delay[2][3] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0367_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold231 (.A(\cic_a.integrator[2][10] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold232 (.A(\cic_b.delay[2][10] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold233 (.A(\cic_a.temp_delay[1][7] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0215_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold235 (.A(\cic_a.delay[2][7] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0111_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold237 (.A(\cic_b.temp_delay[2][6] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0370_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold239 (.A(\serializer_b.shift_reg[6] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0383_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold241 (.A(\serializer_a.shift_reg[9] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0360_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold243 (.A(\cic_a.temp_delay[2][7] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0332_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold245 (.A(\cic_b.temp_comb[2][12] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold246 (.A(\cic_a.temp_comb[2][9] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold247 (.A(\cic_b.temp_delay[2][5] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0369_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold249 (.A(\cic_b.temp_delay[1][3] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0341_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold251 (.A(\cic_a.temp_comb[2][8] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold252 (.A(\cic_a.temp_comb[2][6] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold253 (.A(\cic_b.temp_delay[2][4] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0368_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold255 (.A(\cic_a.temp_delay[1][10] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0218_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold257 (.A(\cic_a.integrator[2][7] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold258 (.A(\serializer_b.shift_reg[7] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0384_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold260 (.A(\cic_b.temp_delay[1][10] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0257_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold262 (.A(\cic_a.temp_delay[1][11] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0219_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold264 (.A(\cic_b.temp_comb[0][10] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold265 (.A(\cic_a.temp_comb[1][10] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold266 (.A(\cic_b.filtered_out[10] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold267 (.A(_1088_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold268 (.A(\cic_a.temp_delay[2][11] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0336_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold270 (.A(\cic_a.temp_delay[2][9] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0334_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold272 (.A(\cic_a.decim_cnt[5] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0005_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold274 (.A(\cic_a.delay[2][0] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold275 (.A(\cic_a.delay[1][12] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold276 (.A(\cic_a.delay[1][11] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold277 (.A(\cic_a.filtered_out[9] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold278 (.A(\cic_b.temp_delay[0][3] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0315_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold280 (.A(\cic_b.temp_delay[0][0] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0312_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold282 (.A(\cic_b.temp_delay[0][7] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0319_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold284 (.A(\cic_b.delay[1][8] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold285 (.A(\cic_b.temp_delay[1][5] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold286 (.A(_0343_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold287 (.A(\cic_a.temp_delay[0][12] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0207_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold289 (.A(\cic_b.delay[1][2] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold290 (.A(\cic_a.temp_delay[1][1] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0209_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold292 (.A(\cic_b.delay[0][0] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold293 (.A(\cic_b.delay[2][2] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold294 (.A(\cic_a.temp_comb[2][4] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold295 (.A(\cic_a.delay[0][11] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold296 (.A(\cic_a.delay[2][1] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold297 (.A(\cic_b.temp_delay[2][11] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0232_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold299 (.A(\cic_b.temp_comb[1][11] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold300 (.A(\cic_b.temp_delay[2][1] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0365_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold302 (.A(\cic_b.delay[0][3] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold303 (.A(\cic_b.temp_delay[2][8] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0372_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold305 (.A(\cic_b.delay[0][8] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold306 (.A(\cic_a.delay[1][1] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold307 (.A(\cic_a.filtered_out[5] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold308 (.A(\cic_a.temp_delay[0][6] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0201_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold310 (.A(\cic_a.delay[1][10] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold311 (.A(\cic_b.temp_delay[1][6] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0344_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold313 (.A(\cic_b.delay[1][7] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold314 (.A(\cic_b.delay[1][5] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold315 (.A(\cic_b.decim_cnt[5] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0013_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold317 (.A(\cic_b.temp_delay[1][1] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0339_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold319 (.A(\cic_a.temp_comb[1][8] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold320 (.A(\cic_b.temp_comb[2][0] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0299_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold322 (.A(\cic_b.delay[2][8] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold323 (.A(\cic_b.temp_delay[2][12] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0376_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold325 (.A(\cic_a.temp_delay[0][4] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0199_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold327 (.A(\cic_b.temp_comb[2][2] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold328 (.A(\cic_b.temp_comb[0][12] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold329 (.A(\cic_b.filtered_out[0] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold330 (.A(\cic_b.delay[2][5] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold331 (.A(\serializer_ab_subtr.shift_reg[11] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold332 (.A(_1178_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold333 (.A(\cic_b.integrator[2][1] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold334 (.A(\cic_b.integrator[2][12] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold335 (.A(\serializer_ab_subtr.shift_reg[10] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold336 (.A(_1172_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold337 (.A(\serializer_a.shift_reg[6] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold338 (.A(_1066_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold339 (.A(\cic_b.delay[1][0] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold340 (.A(\cic_b.delay[1][1] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold341 (.A(\cic_a.filtered_out[1] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold342 (.A(_1058_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold343 (.A(\cic_a.delay[0][12] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold344 (.A(\cic_b.delay[2][12] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold345 (.A(\cic_a.temp_delay[1][8] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0216_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold347 (.A(\cic_b.temp_delay[2][7] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0371_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold349 (.A(\serializer_ab_subtr.shift_reg[6] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold350 (.A(_1144_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold351 (.A(\cic_a.delay[0][6] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold352 (.A(\cic_b.delay[0][7] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold353 (.A(\cic_b.delay[2][7] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold354 (.A(\cic_a.delay[1][2] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold355 (.A(\serializer_a.shift_reg[5] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold356 (.A(_1065_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold357 (.A(\cic_a.delay[2][3] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold358 (.A(\serializer_ab_subtr.shift_reg[5] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold359 (.A(_1137_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0403_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold361 (.A(\cic_a.filtered_out[11] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold362 (.A(\cic_b.filtered_out[7] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold363 (.A(\cic_a.delay[1][5] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold364 (.A(\cic_b.delay[2][3] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold365 (.A(\cic_b.delay[2][6] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold366 (.A(\cic_b.temp_delay[0][4] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0316_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold368 (.A(\cic_a.delay[2][4] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold369 (.A(\cic_a.delay[0][1] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold370 (.A(\cic_a.delay[1][7] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold371 (.A(\cic_a.delay[0][0] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold372 (.A(\cic_a.temp_comb[2][2] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold373 (.A(\cic_b.temp_comb[2][11] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold374 (.A(\cic_a.temp_delay[1][4] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0212_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold376 (.A(\cic_a.temp_delay[2][6] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0331_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold378 (.A(\cic_a.temp_delay[2][5] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0109_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold380 (.A(\cic_b.delay[0][2] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold381 (.A(\serializer_ab_subtr.serial_out ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0410_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold383 (.A(\cic_b.delay[1][3] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold384 (.A(\cic_b.delay[2][1] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold385 (.A(\serializer_ab_subtr.shift_reg[4] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold386 (.A(_1132_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold387 (.A(\cic_a.delay[0][9] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold388 (.A(\serializer_ab_subtr.shift_reg[8] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold389 (.A(_1158_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold390 (.A(\cic_a.temp_comb[1][5] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold391 (.A(\serializer_ab_subtr.shift_reg[7] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold392 (.A(_1149_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold393 (.A(\cic_a.temp_comb[2][12] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0194_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold395 (.A(\cic_a.delay[0][4] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold396 (.A(\cic_a.delay[2][12] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold397 (.A(\cic_b.delay[0][10] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold398 (.A(\cic_b.filtered_out[4] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold399 (.A(\serializer_ab_subtr.shift_reg[2] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold400 (.A(_1118_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0400_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold402 (.A(\cic_a.delay[2][9] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold403 (.A(\cic_b.temp_comb[0][9] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold404 (.A(\cic_b.delay[1][6] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold405 (.A(\cic_a.delay[2][11] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold406 (.A(\cic_b.delay[0][4] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold407 (.A(\serializer_ab_subtr.shift_reg[0] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0398_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold409 (.A(\cic_a.delay[1][4] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold410 (.A(\cic_a.integrator[0][2] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0027_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold412 (.A(\cic_a.filtered_out[12] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold413 (.A(\cic_a.delay[1][8] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold414 (.A(\cic_b.temp_comb[2][10] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold415 (.A(\cic_b.delay[0][6] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold416 (.A(\cic_a.filtered_out[8] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold417 (.A(\cic_a.filtered_out[6] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold418 (.A(\cic_b.integrator[0][2] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0066_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold420 (.A(\cic_a.temp_comb[2][10] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold421 (.A(\cic_b.filtered_out[3] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold422 (.A(\cic_a.temp_comb[0][11] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0167_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold424 (.A(\cic_b.filtered_out[12] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold425 (.A(\serializer_ab_subtr.shift_reg[3] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold426 (.A(_1124_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold427 (.A(\cic_b.filtered_out[9] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold428 (.A(\cic_b.filtered_out[11] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold429 (.A(\cic_b.filtered_out[8] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold430 (.A(\cic_b.filtered_out[6] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold431 (.A(\cic_a.filtered_out[4] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold432 (.A(\cic_a.filtered_out[0] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold433 (.A(\cic_b.integrator[1][0] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0087_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold435 (.A(\cic_a.filtered_out[3] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold436 (.A(\cic_b.integrator[0][0] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold437 (.A(\cic_b.filtered_out[1] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold438 (.A(\cic_b.temp_comb[1][10] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold439 (.A(\cic_a.integrator[1][0] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold440 (.A(_0048_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold441 (.A(\cic_a.filtered_out[10] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold442 (.A(\cic_b.temp_comb[1][12] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0246_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold444 (.A(\serializer_ab_subtr.shift_reg[9] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold445 (.A(_1164_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold446 (.A(\cic_a.filtered_out[2] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold447 (.A(\cic_b.temp_comb[1][7] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold448 (.A(\cic_a.temp_comb[1][12] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold449 (.A(\cic_b.temp_comb[0][2] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0275_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold451 (.A(\cic_b.temp_comb[1][2] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold452 (.A(\cic_a.temp_comb[0][7] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold453 (.A(\cic_b.temp_comb[0][9] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0880_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold455 (.A(\cic_a.temp_comb[0][0] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0156_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold457 (.A(\cic_b.integrator[0][5] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0069_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold459 (.A(\cic_a.integrator[0][9] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0034_),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold461 (.A(\cic_a.temp_comb[0][10] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold462 (.A(\cic_a.integrator[0][0] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold463 (.A(\cic_a.temp_comb[1][9] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold464 (.A(\cic_b.delay[0][12] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold465 (.A(\cic_b.temp_comb[0][5] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold466 (.A(\cic_b.integrator[0][9] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold467 (.A(_0073_),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold468 (.A(\cic_b.temp_comb[0][1] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold469 (.A(_0274_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold470 (.A(\cic_b.temp_comb[0][7] ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold471 (.A(\cic_b.temp_comb[1][8] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold472 (.A(\cic_b.temp_comb[1][4] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0238_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold474 (.A(\cic_b.temp_comb[1][0] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0234_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold476 (.A(\cic_b.temp_comb[1][1] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold477 (.A(_0235_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold478 (.A(\cic_b.integrator[1][12] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0077_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold480 (.A(\cic_a.temp_comb[0][3] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold481 (.A(_0159_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold482 (.A(\cic_b.delay[0][9] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold483 (.A(\cic_b.temp_comb[0][8] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold484 (.A(\cic_a.decim_cnt[3] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold485 (.A(\cic_b.integrator[0][7] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold486 (.A(_0071_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold487 (.A(\cic_b.temp_comb[0][0] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold488 (.A(_0273_),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold489 (.A(\cic_a.temp_comb[0][2] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold490 (.A(_0158_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold491 (.A(\cic_a.temp_comb[0][8] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold492 (.A(\cic_a.temp_comb[0][12] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0168_),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold494 (.A(\cic_b.integrator[2][10] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold495 (.A(\cic_a.temp_comb[0][1] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold496 (.A(\cic_b.temp_comb[1][6] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold497 (.A(\cic_a.temp_comb[0][5] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0624_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold499 (.A(\cic_a.temp_comb[1][0] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold500 (.A(\cic_b.integrator[0][10] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold501 (.A(\cic_a.delay[0][5] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold502 (.A(\cic_b.decim_cnt[3] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold503 (.A(\cic_a.integrator[0][5] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold504 (.A(_0030_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold505 (.A(\cic_a.integrator[0][10] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold506 (.A(\cic_b.temp_comb[0][6] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold507 (.A(\cic_a.temp_comb[1][2] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold508 (.A(\cic_a.temp_comb[0][4] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold509 (.A(\cic_a.integrator[0][6] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold510 (.A(_0031_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold511 (.A(\cic_b.temp_comb[0][3] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold512 (.A(\cic_a.temp_comb[1][7] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold513 (.A(\cic_b.temp_comb[1][3] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold514 (.A(_0237_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold515 (.A(\cic_a.integrator[0][3] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0028_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold517 (.A(\cic_a.temp_comb[1][3] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold518 (.A(_0120_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold519 (.A(\cic_b.temp_comb[1][5] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold520 (.A(\cic_a.integrator[0][7] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold521 (.A(_0032_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold522 (.A(\cic_b.integrator[0][6] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0070_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold524 (.A(\cic_a.temp_comb[1][11] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold525 (.A(\cic_b.integrator[0][3] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold526 (.A(\cic_a.temp_comb[1][6] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold527 (.A(\cic_a.temp_comb[1][4] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold528 (.A(\cic_b.integrator[1][11] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold529 (.A(_0520_),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold530 (.A(\cic_a.integrator[1][12] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0038_),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold532 (.A(\cic_a.temp_comb[1][1] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold533 (.A(\cic_a.integrator[2][12] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold534 (.A(_0051_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold535 (.A(\serializer_b.sending ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold536 (.A(net543),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold537 (.A(\cic_a.integrator[0][1] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold538 (.A(_0423_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold539 (.A(\cic_a.decim_cnt[4] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold540 (.A(\cic_b.decim_cnt[4] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold541 (.A(\cic_b.integrator[1][10] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold542 (.A(\cic_b.integrator[1][1] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold543 (.A(_0091_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold544 (.A(\cic_a.integrator[2][0] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold545 (.A(_0052_),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold546 (.A(\cic_a.integrator[0][0] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold547 (.A(\cic_a.integrator[0][8] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0033_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold549 (.A(\cic_b.integrator[0][1] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold550 (.A(\cic_b.integrator[1][3] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold551 (.A(_0080_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold552 (.A(\cic_a.integrator[0][4] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold553 (.A(\cic_b.integrator[0][0] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold554 (.A(\cic_a.integrator[0][11] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold555 (.A(\cic_b.integrator[0][11] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold556 (.A(\cic_a.integrator[2][9] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold557 (.A(_1303_),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold558 (.A(_0060_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold559 (.A(\cic_b.integrator[0][8] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold560 (.A(_0072_),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold561 (.A(\cic_b.integrator[0][4] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold562 (.A(\cic_a.integrator[1][11] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold563 (.A(_0037_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold564 (.A(\cic_a.integrator[1][6] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold565 (.A(\cic_b.integrator[0][10] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold566 (.A(_0564_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold567 (.A(\cic_a.integrator[1][3] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold568 (.A(_0054_),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold569 (.A(\cic_a.integrator[1][2] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold570 (.A(\cic_b.integrator[1][9] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold571 (.A(_0086_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold572 (.A(\cic_a.integrator[1][7] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0045_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold574 (.A(\cic_b.integrator[1][6] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold575 (.A(_0083_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold576 (.A(\cic_b.integrator[1][8] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold577 (.A(_0504_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold578 (.A(\cic_a.integrator[1][8] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold579 (.A(_0047_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold580 (.A(\cic_b.integrator[2][6] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold581 (.A(\cic_a.integrator[1][7] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold582 (.A(\cic_a.integrator[1][4] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold583 (.A(_1278_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold584 (.A(\cic_b.integrator[1][7] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold585 (.A(_0549_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold586 (.A(\cic_a.integrator[1][10] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold587 (.A(_0036_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold588 (.A(\cic_b.integrator[1][4] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold589 (.A(_0483_),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold590 (.A(_0095_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold591 (.A(\cic_b.integrator[1][1] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold592 (.A(_0478_),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold593 (.A(_0092_),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold594 (.A(\cic_b.integrator[0][9] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold595 (.A(\cic_a.integrator[2][11] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold596 (.A(\cic_b.integrator[2][4] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold597 (.A(\cic_a.integrator[0][5] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold598 (.A(_0436_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold599 (.A(\cic_a.integrator[2][6] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold600 (.A(_0058_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold601 (.A(\cic_a.integrator[2][9] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold602 (.A(\cic_b.integrator[2][3] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold603 (.A(\cic_b.integrator[1][5] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold604 (.A(_0540_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold605 (.A(\cic_a.integrator[1][2] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold606 (.A(_0053_),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold607 (.A(\cic_b.integrator[2][8] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold608 (.A(\cic_b.integrator[1][2] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold609 (.A(\cic_b.integrator[1][6] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold610 (.A(_0097_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold611 (.A(\cic_b.integrator[0][6] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold612 (.A(_0084_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold613 (.A(\cic_a.integrator[0][1] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold614 (.A(\cic_a.integrator[0][3] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold615 (.A(_0042_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold616 (.A(\cic_b.integrator[0][3] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold617 (.A(_0081_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold618 (.A(\cic_a.integrator[1][3] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold619 (.A(_0055_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold620 (.A(\cic_a.integrator[1][6] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold621 (.A(_1287_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold622 (.A(\cic_a.integrator[0][7] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold623 (.A(\cic_b.temp_comb[0][8] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold624 (.A(\cic_b.temp_comb[0][8] ),
    .X(net792));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_fill_1 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_108 ();
 sg13g2_decap_4 FILLER_0_115 ();
 sg13g2_fill_1 FILLER_0_119 ();
 sg13g2_decap_4 FILLER_0_137 ();
 sg13g2_fill_2 FILLER_0_141 ();
 sg13g2_decap_4 FILLER_0_169 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_4 FILLER_0_217 ();
 sg13g2_fill_2 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_244 ();
 sg13g2_decap_8 FILLER_0_251 ();
 sg13g2_decap_8 FILLER_0_258 ();
 sg13g2_decap_8 FILLER_0_265 ();
 sg13g2_decap_8 FILLER_0_272 ();
 sg13g2_decap_8 FILLER_0_279 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_293 ();
 sg13g2_decap_8 FILLER_0_300 ();
 sg13g2_decap_8 FILLER_0_307 ();
 sg13g2_decap_8 FILLER_0_314 ();
 sg13g2_decap_8 FILLER_0_321 ();
 sg13g2_decap_8 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_4 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_fill_1 FILLER_1_84 ();
 sg13g2_fill_1 FILLER_1_140 ();
 sg13g2_decap_4 FILLER_1_201 ();
 sg13g2_fill_1 FILLER_1_205 ();
 sg13g2_decap_4 FILLER_1_232 ();
 sg13g2_fill_1 FILLER_1_236 ();
 sg13g2_fill_1 FILLER_1_263 ();
 sg13g2_decap_8 FILLER_1_290 ();
 sg13g2_fill_2 FILLER_1_297 ();
 sg13g2_decap_8 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_342 ();
 sg13g2_decap_8 FILLER_1_349 ();
 sg13g2_decap_8 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_8 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_fill_1 FILLER_2_77 ();
 sg13g2_decap_4 FILLER_2_166 ();
 sg13g2_fill_2 FILLER_2_170 ();
 sg13g2_fill_1 FILLER_2_206 ();
 sg13g2_decap_8 FILLER_2_341 ();
 sg13g2_decap_8 FILLER_2_348 ();
 sg13g2_decap_8 FILLER_2_355 ();
 sg13g2_decap_8 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_376 ();
 sg13g2_decap_8 FILLER_2_383 ();
 sg13g2_decap_8 FILLER_2_390 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_4 FILLER_2_404 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_fill_2 FILLER_3_70 ();
 sg13g2_fill_1 FILLER_3_72 ();
 sg13g2_fill_1 FILLER_3_117 ();
 sg13g2_fill_1 FILLER_3_135 ();
 sg13g2_fill_1 FILLER_3_154 ();
 sg13g2_decap_4 FILLER_3_164 ();
 sg13g2_fill_2 FILLER_3_168 ();
 sg13g2_fill_2 FILLER_3_242 ();
 sg13g2_fill_1 FILLER_3_244 ();
 sg13g2_fill_1 FILLER_3_285 ();
 sg13g2_decap_8 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_356 ();
 sg13g2_decap_8 FILLER_3_363 ();
 sg13g2_decap_8 FILLER_3_370 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_fill_2 FILLER_4_70 ();
 sg13g2_fill_1 FILLER_4_72 ();
 sg13g2_decap_8 FILLER_4_78 ();
 sg13g2_fill_2 FILLER_4_85 ();
 sg13g2_fill_1 FILLER_4_87 ();
 sg13g2_fill_2 FILLER_4_97 ();
 sg13g2_fill_1 FILLER_4_99 ();
 sg13g2_decap_4 FILLER_4_109 ();
 sg13g2_fill_2 FILLER_4_113 ();
 sg13g2_fill_1 FILLER_4_141 ();
 sg13g2_decap_8 FILLER_4_177 ();
 sg13g2_fill_1 FILLER_4_229 ();
 sg13g2_fill_2 FILLER_4_311 ();
 sg13g2_fill_1 FILLER_4_313 ();
 sg13g2_decap_8 FILLER_4_337 ();
 sg13g2_decap_4 FILLER_4_344 ();
 sg13g2_decap_8 FILLER_4_374 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_fill_2 FILLER_5_35 ();
 sg13g2_fill_1 FILLER_5_37 ();
 sg13g2_fill_2 FILLER_5_64 ();
 sg13g2_decap_4 FILLER_5_73 ();
 sg13g2_fill_1 FILLER_5_92 ();
 sg13g2_decap_4 FILLER_5_102 ();
 sg13g2_decap_4 FILLER_5_131 ();
 sg13g2_decap_4 FILLER_5_144 ();
 sg13g2_decap_4 FILLER_5_157 ();
 sg13g2_fill_2 FILLER_5_179 ();
 sg13g2_fill_1 FILLER_5_181 ();
 sg13g2_decap_4 FILLER_5_191 ();
 sg13g2_decap_4 FILLER_5_251 ();
 sg13g2_decap_4 FILLER_5_274 ();
 sg13g2_fill_2 FILLER_5_283 ();
 sg13g2_fill_1 FILLER_5_285 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_4 FILLER_6_42 ();
 sg13g2_fill_1 FILLER_6_55 ();
 sg13g2_fill_2 FILLER_6_91 ();
 sg13g2_fill_1 FILLER_6_93 ();
 sg13g2_fill_2 FILLER_6_171 ();
 sg13g2_fill_1 FILLER_6_173 ();
 sg13g2_fill_1 FILLER_6_196 ();
 sg13g2_decap_4 FILLER_6_206 ();
 sg13g2_fill_1 FILLER_6_215 ();
 sg13g2_fill_2 FILLER_6_229 ();
 sg13g2_fill_2 FILLER_6_284 ();
 sg13g2_decap_4 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_369 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_8 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_fill_1 FILLER_7_42 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_58 ();
 sg13g2_fill_2 FILLER_7_129 ();
 sg13g2_fill_1 FILLER_7_131 ();
 sg13g2_fill_2 FILLER_7_146 ();
 sg13g2_decap_4 FILLER_7_156 ();
 sg13g2_decap_8 FILLER_7_173 ();
 sg13g2_decap_8 FILLER_7_206 ();
 sg13g2_fill_2 FILLER_7_213 ();
 sg13g2_fill_1 FILLER_7_215 ();
 sg13g2_fill_2 FILLER_7_240 ();
 sg13g2_fill_2 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_338 ();
 sg13g2_fill_1 FILLER_7_345 ();
 sg13g2_decap_8 FILLER_7_355 ();
 sg13g2_decap_8 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_369 ();
 sg13g2_decap_8 FILLER_7_376 ();
 sg13g2_decap_8 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_4 FILLER_8_49 ();
 sg13g2_fill_1 FILLER_8_86 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_fill_2 FILLER_8_168 ();
 sg13g2_decap_4 FILLER_8_212 ();
 sg13g2_fill_2 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_fill_1 FILLER_8_275 ();
 sg13g2_fill_2 FILLER_8_285 ();
 sg13g2_fill_1 FILLER_8_287 ();
 sg13g2_fill_2 FILLER_8_306 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_4 FILLER_9_35 ();
 sg13g2_fill_1 FILLER_9_39 ();
 sg13g2_fill_1 FILLER_9_70 ();
 sg13g2_decap_4 FILLER_9_79 ();
 sg13g2_fill_2 FILLER_9_83 ();
 sg13g2_fill_2 FILLER_9_93 ();
 sg13g2_fill_1 FILLER_9_95 ();
 sg13g2_fill_2 FILLER_9_122 ();
 sg13g2_fill_1 FILLER_9_143 ();
 sg13g2_decap_8 FILLER_9_149 ();
 sg13g2_fill_1 FILLER_9_156 ();
 sg13g2_fill_1 FILLER_9_183 ();
 sg13g2_fill_1 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_195 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_fill_1 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_247 ();
 sg13g2_decap_8 FILLER_9_254 ();
 sg13g2_decap_8 FILLER_9_261 ();
 sg13g2_fill_1 FILLER_9_268 ();
 sg13g2_decap_8 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_281 ();
 sg13g2_fill_2 FILLER_9_288 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_fill_2 FILLER_9_301 ();
 sg13g2_fill_1 FILLER_9_303 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_381 ();
 sg13g2_decap_8 FILLER_9_388 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_fill_2 FILLER_10_42 ();
 sg13g2_fill_1 FILLER_10_44 ();
 sg13g2_fill_1 FILLER_10_80 ();
 sg13g2_fill_1 FILLER_10_90 ();
 sg13g2_decap_4 FILLER_10_96 ();
 sg13g2_fill_2 FILLER_10_100 ();
 sg13g2_fill_2 FILLER_10_105 ();
 sg13g2_fill_2 FILLER_10_186 ();
 sg13g2_fill_1 FILLER_10_188 ();
 sg13g2_fill_1 FILLER_10_194 ();
 sg13g2_fill_1 FILLER_10_231 ();
 sg13g2_decap_4 FILLER_10_242 ();
 sg13g2_fill_1 FILLER_10_256 ();
 sg13g2_fill_1 FILLER_10_274 ();
 sg13g2_fill_2 FILLER_10_311 ();
 sg13g2_decap_8 FILLER_10_339 ();
 sg13g2_decap_4 FILLER_10_346 ();
 sg13g2_fill_1 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_4 FILLER_11_42 ();
 sg13g2_fill_1 FILLER_11_46 ();
 sg13g2_fill_1 FILLER_11_59 ();
 sg13g2_decap_8 FILLER_11_104 ();
 sg13g2_decap_4 FILLER_11_111 ();
 sg13g2_fill_2 FILLER_11_115 ();
 sg13g2_decap_8 FILLER_11_121 ();
 sg13g2_decap_8 FILLER_11_128 ();
 sg13g2_decap_8 FILLER_11_135 ();
 sg13g2_decap_4 FILLER_11_142 ();
 sg13g2_fill_2 FILLER_11_146 ();
 sg13g2_fill_1 FILLER_11_152 ();
 sg13g2_fill_1 FILLER_11_185 ();
 sg13g2_fill_2 FILLER_11_194 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_fill_1 FILLER_11_216 ();
 sg13g2_fill_2 FILLER_11_226 ();
 sg13g2_fill_1 FILLER_11_228 ();
 sg13g2_decap_4 FILLER_11_325 ();
 sg13g2_fill_2 FILLER_11_329 ();
 sg13g2_fill_2 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_395 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_4 FILLER_12_49 ();
 sg13g2_fill_1 FILLER_12_53 ();
 sg13g2_fill_1 FILLER_12_107 ();
 sg13g2_decap_8 FILLER_12_113 ();
 sg13g2_decap_8 FILLER_12_120 ();
 sg13g2_decap_8 FILLER_12_127 ();
 sg13g2_decap_8 FILLER_12_134 ();
 sg13g2_decap_8 FILLER_12_141 ();
 sg13g2_decap_4 FILLER_12_148 ();
 sg13g2_fill_2 FILLER_12_152 ();
 sg13g2_decap_4 FILLER_12_204 ();
 sg13g2_fill_1 FILLER_12_208 ();
 sg13g2_decap_8 FILLER_12_218 ();
 sg13g2_decap_4 FILLER_12_225 ();
 sg13g2_fill_2 FILLER_12_229 ();
 sg13g2_decap_4 FILLER_12_240 ();
 sg13g2_fill_2 FILLER_12_244 ();
 sg13g2_decap_4 FILLER_12_255 ();
 sg13g2_fill_2 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_4 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_fill_2 FILLER_13_42 ();
 sg13g2_fill_1 FILLER_13_44 ();
 sg13g2_fill_2 FILLER_13_71 ();
 sg13g2_decap_4 FILLER_13_83 ();
 sg13g2_decap_4 FILLER_13_131 ();
 sg13g2_fill_1 FILLER_13_135 ();
 sg13g2_fill_2 FILLER_13_144 ();
 sg13g2_fill_1 FILLER_13_146 ();
 sg13g2_decap_8 FILLER_13_162 ();
 sg13g2_fill_1 FILLER_13_169 ();
 sg13g2_decap_4 FILLER_13_179 ();
 sg13g2_fill_2 FILLER_13_183 ();
 sg13g2_fill_1 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_225 ();
 sg13g2_fill_2 FILLER_13_230 ();
 sg13g2_fill_1 FILLER_13_250 ();
 sg13g2_fill_1 FILLER_13_268 ();
 sg13g2_decap_4 FILLER_13_279 ();
 sg13g2_decap_8 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_306 ();
 sg13g2_decap_4 FILLER_13_313 ();
 sg13g2_fill_2 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_fill_1 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_decap_4 FILLER_13_367 ();
 sg13g2_fill_2 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_fill_1 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_55 ();
 sg13g2_decap_4 FILLER_14_71 ();
 sg13g2_fill_1 FILLER_14_75 ();
 sg13g2_fill_2 FILLER_14_132 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_8 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_decap_4 FILLER_14_207 ();
 sg13g2_fill_2 FILLER_14_237 ();
 sg13g2_fill_1 FILLER_14_239 ();
 sg13g2_decap_4 FILLER_14_266 ();
 sg13g2_fill_1 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_279 ();
 sg13g2_decap_8 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_305 ();
 sg13g2_fill_1 FILLER_14_312 ();
 sg13g2_fill_1 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_64 ();
 sg13g2_decap_4 FILLER_15_71 ();
 sg13g2_fill_1 FILLER_15_75 ();
 sg13g2_decap_8 FILLER_15_129 ();
 sg13g2_fill_2 FILLER_15_136 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_fill_1 FILLER_15_165 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_decap_8 FILLER_15_204 ();
 sg13g2_fill_2 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_216 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_fill_2 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_317 ();
 sg13g2_decap_4 FILLER_15_324 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_22 ();
 sg13g2_decap_4 FILLER_16_29 ();
 sg13g2_decap_8 FILLER_16_72 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_decap_8 FILLER_16_85 ();
 sg13g2_decap_8 FILLER_16_92 ();
 sg13g2_decap_4 FILLER_16_99 ();
 sg13g2_fill_1 FILLER_16_103 ();
 sg13g2_decap_8 FILLER_16_113 ();
 sg13g2_fill_1 FILLER_16_120 ();
 sg13g2_fill_2 FILLER_16_125 ();
 sg13g2_decap_8 FILLER_16_136 ();
 sg13g2_decap_8 FILLER_16_143 ();
 sg13g2_decap_8 FILLER_16_150 ();
 sg13g2_fill_2 FILLER_16_157 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_fill_1 FILLER_16_224 ();
 sg13g2_fill_2 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_fill_2 FILLER_16_332 ();
 sg13g2_fill_1 FILLER_16_348 ();
 sg13g2_fill_1 FILLER_16_359 ();
 sg13g2_fill_1 FILLER_16_374 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_2 FILLER_17_41 ();
 sg13g2_fill_1 FILLER_17_43 ();
 sg13g2_decap_8 FILLER_17_80 ();
 sg13g2_fill_2 FILLER_17_103 ();
 sg13g2_fill_1 FILLER_17_127 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_decap_8 FILLER_17_240 ();
 sg13g2_fill_1 FILLER_17_273 ();
 sg13g2_fill_1 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_332 ();
 sg13g2_fill_1 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_fill_2 FILLER_17_357 ();
 sg13g2_fill_1 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_83 ();
 sg13g2_decap_8 FILLER_18_90 ();
 sg13g2_decap_8 FILLER_18_97 ();
 sg13g2_fill_2 FILLER_18_104 ();
 sg13g2_fill_2 FILLER_18_158 ();
 sg13g2_decap_4 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_182 ();
 sg13g2_fill_1 FILLER_18_184 ();
 sg13g2_fill_2 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_4 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_240 ();
 sg13g2_fill_1 FILLER_18_247 ();
 sg13g2_fill_2 FILLER_18_257 ();
 sg13g2_fill_2 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_312 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_329 ();
 sg13g2_decap_4 FILLER_18_356 ();
 sg13g2_fill_2 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_34 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_118 ();
 sg13g2_fill_1 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_187 ();
 sg13g2_fill_1 FILLER_19_238 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_fill_2 FILLER_19_294 ();
 sg13g2_fill_1 FILLER_19_339 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_fill_1 FILLER_19_372 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_19_392 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_31 ();
 sg13g2_fill_1 FILLER_20_33 ();
 sg13g2_decap_4 FILLER_20_133 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_decap_4 FILLER_20_147 ();
 sg13g2_fill_2 FILLER_20_151 ();
 sg13g2_fill_2 FILLER_20_162 ();
 sg13g2_decap_8 FILLER_20_208 ();
 sg13g2_decap_4 FILLER_20_215 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_decap_8 FILLER_20_279 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_fill_1 FILLER_20_320 ();
 sg13g2_fill_2 FILLER_20_331 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_fill_2 FILLER_21_43 ();
 sg13g2_fill_1 FILLER_21_45 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_fill_2 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_77 ();
 sg13g2_fill_2 FILLER_21_94 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_fill_2 FILLER_21_126 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_fill_2 FILLER_21_138 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_fill_2 FILLER_21_163 ();
 sg13g2_decap_8 FILLER_21_173 ();
 sg13g2_decap_4 FILLER_21_180 ();
 sg13g2_decap_4 FILLER_21_192 ();
 sg13g2_fill_2 FILLER_21_196 ();
 sg13g2_decap_4 FILLER_21_210 ();
 sg13g2_decap_4 FILLER_21_218 ();
 sg13g2_fill_1 FILLER_21_245 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_fill_2 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_277 ();
 sg13g2_fill_2 FILLER_21_327 ();
 sg13g2_fill_2 FILLER_21_342 ();
 sg13g2_fill_1 FILLER_21_344 ();
 sg13g2_fill_2 FILLER_21_371 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_fill_2 FILLER_22_98 ();
 sg13g2_decap_4 FILLER_22_136 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_2 FILLER_22_147 ();
 sg13g2_fill_1 FILLER_22_149 ();
 sg13g2_fill_1 FILLER_22_164 ();
 sg13g2_fill_2 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_197 ();
 sg13g2_fill_1 FILLER_22_230 ();
 sg13g2_fill_1 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_307 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_fill_2 FILLER_22_352 ();
 sg13g2_decap_4 FILLER_22_364 ();
 sg13g2_fill_1 FILLER_22_377 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_2 FILLER_23_33 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_81 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_decap_8 FILLER_23_120 ();
 sg13g2_fill_2 FILLER_23_127 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_fill_1 FILLER_23_139 ();
 sg13g2_fill_2 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_fill_1 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_fill_2 FILLER_23_305 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_decap_4 FILLER_23_333 ();
 sg13g2_fill_1 FILLER_23_337 ();
 sg13g2_decap_4 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_351 ();
 sg13g2_decap_4 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_365 ();
 sg13g2_decap_4 FILLER_23_384 ();
 sg13g2_fill_1 FILLER_23_388 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_1 FILLER_24_26 ();
 sg13g2_fill_1 FILLER_24_32 ();
 sg13g2_fill_1 FILLER_24_59 ();
 sg13g2_fill_2 FILLER_24_70 ();
 sg13g2_fill_1 FILLER_24_72 ();
 sg13g2_decap_8 FILLER_24_82 ();
 sg13g2_fill_2 FILLER_24_89 ();
 sg13g2_decap_8 FILLER_24_99 ();
 sg13g2_decap_4 FILLER_24_106 ();
 sg13g2_fill_1 FILLER_24_110 ();
 sg13g2_fill_2 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_157 ();
 sg13g2_fill_1 FILLER_24_184 ();
 sg13g2_fill_1 FILLER_24_194 ();
 sg13g2_fill_2 FILLER_24_242 ();
 sg13g2_fill_1 FILLER_24_244 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_4 FILLER_24_285 ();
 sg13g2_fill_1 FILLER_24_289 ();
 sg13g2_decap_4 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_304 ();
 sg13g2_fill_2 FILLER_24_379 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_57 ();
 sg13g2_decap_8 FILLER_25_64 ();
 sg13g2_fill_2 FILLER_25_79 ();
 sg13g2_fill_2 FILLER_25_117 ();
 sg13g2_decap_4 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_169 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_fill_1 FILLER_25_222 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_decap_8 FILLER_25_271 ();
 sg13g2_fill_2 FILLER_25_278 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_4 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_decap_4 FILLER_25_359 ();
 sg13g2_fill_2 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_42 ();
 sg13g2_fill_1 FILLER_26_46 ();
 sg13g2_decap_8 FILLER_26_55 ();
 sg13g2_decap_8 FILLER_26_62 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_121 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_4 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_189 ();
 sg13g2_fill_1 FILLER_26_195 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_260 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_decap_4 FILLER_26_320 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_fill_2 FILLER_26_356 ();
 sg13g2_fill_2 FILLER_26_366 ();
 sg13g2_fill_1 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_27_26 ();
 sg13g2_decap_4 FILLER_27_33 ();
 sg13g2_decap_4 FILLER_27_72 ();
 sg13g2_fill_1 FILLER_27_76 ();
 sg13g2_fill_1 FILLER_27_121 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_decap_8 FILLER_27_132 ();
 sg13g2_decap_8 FILLER_27_148 ();
 sg13g2_decap_8 FILLER_27_165 ();
 sg13g2_decap_8 FILLER_27_172 ();
 sg13g2_decap_4 FILLER_27_179 ();
 sg13g2_decap_8 FILLER_27_186 ();
 sg13g2_decap_4 FILLER_27_193 ();
 sg13g2_fill_2 FILLER_27_197 ();
 sg13g2_decap_8 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_decap_4 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_258 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_fill_2 FILLER_27_308 ();
 sg13g2_fill_1 FILLER_27_310 ();
 sg13g2_decap_8 FILLER_27_320 ();
 sg13g2_fill_1 FILLER_27_327 ();
 sg13g2_decap_8 FILLER_27_333 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_8 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_354 ();
 sg13g2_fill_2 FILLER_27_361 ();
 sg13g2_fill_1 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_374 ();
 sg13g2_fill_2 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_fill_2 FILLER_28_44 ();
 sg13g2_fill_1 FILLER_28_46 ();
 sg13g2_decap_4 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_85 ();
 sg13g2_decap_8 FILLER_28_114 ();
 sg13g2_fill_2 FILLER_28_121 ();
 sg13g2_decap_8 FILLER_28_127 ();
 sg13g2_decap_8 FILLER_28_134 ();
 sg13g2_decap_8 FILLER_28_141 ();
 sg13g2_decap_8 FILLER_28_148 ();
 sg13g2_decap_4 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_fill_2 FILLER_28_310 ();
 sg13g2_fill_2 FILLER_28_317 ();
 sg13g2_decap_4 FILLER_28_359 ();
 sg13g2_fill_2 FILLER_28_363 ();
 sg13g2_decap_4 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_28_388 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_fill_1 FILLER_29_33 ();
 sg13g2_fill_1 FILLER_29_43 ();
 sg13g2_decap_4 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_4 FILLER_29_98 ();
 sg13g2_fill_2 FILLER_29_102 ();
 sg13g2_fill_2 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_199 ();
 sg13g2_decap_4 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_261 ();
 sg13g2_fill_2 FILLER_29_268 ();
 sg13g2_fill_1 FILLER_29_270 ();
 sg13g2_fill_1 FILLER_29_280 ();
 sg13g2_decap_4 FILLER_29_310 ();
 sg13g2_fill_1 FILLER_29_359 ();
 sg13g2_decap_4 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_6 ();
 sg13g2_decap_8 FILLER_30_32 ();
 sg13g2_decap_8 FILLER_30_39 ();
 sg13g2_decap_4 FILLER_30_46 ();
 sg13g2_fill_1 FILLER_30_50 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_fill_1 FILLER_30_71 ();
 sg13g2_decap_8 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_88 ();
 sg13g2_decap_4 FILLER_30_93 ();
 sg13g2_decap_4 FILLER_30_102 ();
 sg13g2_fill_2 FILLER_30_106 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_decap_4 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_fill_1 FILLER_30_216 ();
 sg13g2_decap_8 FILLER_30_230 ();
 sg13g2_decap_4 FILLER_30_237 ();
 sg13g2_fill_2 FILLER_30_241 ();
 sg13g2_fill_2 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_decap_4 FILLER_30_345 ();
 sg13g2_fill_1 FILLER_30_375 ();
 sg13g2_fill_2 FILLER_30_384 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_fill_1 FILLER_31_15 ();
 sg13g2_fill_2 FILLER_31_25 ();
 sg13g2_fill_1 FILLER_31_51 ();
 sg13g2_decap_4 FILLER_31_66 ();
 sg13g2_fill_1 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_fill_1 FILLER_31_119 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_fill_2 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_decap_8 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_fill_2 FILLER_31_291 ();
 sg13g2_fill_1 FILLER_31_293 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_fill_2 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_368 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_18 ();
 sg13g2_decap_4 FILLER_32_118 ();
 sg13g2_fill_1 FILLER_32_122 ();
 sg13g2_decap_8 FILLER_32_144 ();
 sg13g2_fill_2 FILLER_32_156 ();
 sg13g2_decap_4 FILLER_32_163 ();
 sg13g2_fill_2 FILLER_32_167 ();
 sg13g2_fill_2 FILLER_32_173 ();
 sg13g2_fill_1 FILLER_32_179 ();
 sg13g2_fill_2 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_decap_8 FILLER_32_201 ();
 sg13g2_decap_8 FILLER_32_208 ();
 sg13g2_decap_8 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_229 ();
 sg13g2_decap_8 FILLER_32_236 ();
 sg13g2_fill_2 FILLER_32_243 ();
 sg13g2_decap_8 FILLER_32_316 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_decap_4 FILLER_32_328 ();
 sg13g2_decap_8 FILLER_32_337 ();
 sg13g2_decap_4 FILLER_32_344 ();
 sg13g2_decap_8 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_360 ();
 sg13g2_decap_8 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_fill_2 FILLER_32_386 ();
 sg13g2_fill_1 FILLER_32_388 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_30 ();
 sg13g2_fill_2 FILLER_33_52 ();
 sg13g2_fill_1 FILLER_33_54 ();
 sg13g2_fill_2 FILLER_33_73 ();
 sg13g2_fill_2 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_86 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_fill_1 FILLER_33_130 ();
 sg13g2_decap_8 FILLER_33_136 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_161 ();
 sg13g2_fill_2 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_179 ();
 sg13g2_decap_4 FILLER_33_206 ();
 sg13g2_fill_2 FILLER_33_210 ();
 sg13g2_fill_1 FILLER_33_225 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_fill_2 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_decap_8 FILLER_33_265 ();
 sg13g2_decap_4 FILLER_33_272 ();
 sg13g2_fill_1 FILLER_33_276 ();
 sg13g2_decap_8 FILLER_33_285 ();
 sg13g2_decap_8 FILLER_33_292 ();
 sg13g2_decap_8 FILLER_33_299 ();
 sg13g2_decap_8 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_313 ();
 sg13g2_decap_8 FILLER_33_320 ();
 sg13g2_fill_1 FILLER_33_327 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_343 ();
 sg13g2_fill_1 FILLER_33_355 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_decap_4 FILLER_33_385 ();
 sg13g2_fill_2 FILLER_33_389 ();
 sg13g2_fill_2 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_16 ();
 sg13g2_fill_2 FILLER_34_30 ();
 sg13g2_fill_1 FILLER_34_54 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_4 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_95 ();
 sg13g2_fill_2 FILLER_34_184 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_fill_2 FILLER_34_248 ();
 sg13g2_fill_1 FILLER_34_250 ();
 sg13g2_decap_4 FILLER_34_277 ();
 sg13g2_fill_2 FILLER_34_281 ();
 sg13g2_decap_8 FILLER_34_288 ();
 sg13g2_fill_2 FILLER_34_295 ();
 sg13g2_fill_1 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_324 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_55 ();
 sg13g2_fill_1 FILLER_35_57 ();
 sg13g2_fill_2 FILLER_35_71 ();
 sg13g2_fill_1 FILLER_35_73 ();
 sg13g2_fill_1 FILLER_35_78 ();
 sg13g2_fill_1 FILLER_35_83 ();
 sg13g2_decap_4 FILLER_35_93 ();
 sg13g2_decap_4 FILLER_35_106 ();
 sg13g2_fill_1 FILLER_35_110 ();
 sg13g2_decap_8 FILLER_35_116 ();
 sg13g2_decap_4 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_132 ();
 sg13g2_decap_8 FILLER_35_138 ();
 sg13g2_decap_8 FILLER_35_145 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_193 ();
 sg13g2_fill_1 FILLER_35_195 ();
 sg13g2_fill_2 FILLER_35_214 ();
 sg13g2_decap_8 FILLER_35_234 ();
 sg13g2_decap_8 FILLER_35_241 ();
 sg13g2_fill_2 FILLER_35_267 ();
 sg13g2_decap_4 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_382 ();
 sg13g2_fill_2 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_60 ();
 sg13g2_fill_1 FILLER_36_92 ();
 sg13g2_fill_1 FILLER_36_115 ();
 sg13g2_decap_8 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_192 ();
 sg13g2_fill_1 FILLER_36_214 ();
 sg13g2_fill_1 FILLER_36_223 ();
 sg13g2_decap_4 FILLER_36_250 ();
 sg13g2_fill_1 FILLER_36_262 ();
 sg13g2_decap_8 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_297 ();
 sg13g2_fill_2 FILLER_36_335 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_2 FILLER_36_371 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_28 ();
 sg13g2_decap_4 FILLER_37_118 ();
 sg13g2_fill_2 FILLER_37_122 ();
 sg13g2_decap_4 FILLER_37_128 ();
 sg13g2_fill_2 FILLER_37_156 ();
 sg13g2_fill_1 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_195 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_decap_4 FILLER_37_233 ();
 sg13g2_decap_8 FILLER_37_292 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_fill_1 FILLER_37_315 ();
 sg13g2_fill_2 FILLER_37_336 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_356 ();
 sg13g2_decap_4 FILLER_37_363 ();
 sg13g2_fill_2 FILLER_37_375 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_4 ();
 sg13g2_decap_4 FILLER_38_13 ();
 sg13g2_fill_2 FILLER_38_17 ();
 sg13g2_decap_8 FILLER_38_37 ();
 sg13g2_fill_1 FILLER_38_44 ();
 sg13g2_fill_2 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_57 ();
 sg13g2_fill_2 FILLER_38_67 ();
 sg13g2_decap_4 FILLER_38_98 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_decap_8 FILLER_38_122 ();
 sg13g2_decap_8 FILLER_38_129 ();
 sg13g2_fill_1 FILLER_38_136 ();
 sg13g2_fill_2 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_240 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_decap_4 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_256 ();
 sg13g2_fill_2 FILLER_38_281 ();
 sg13g2_fill_2 FILLER_38_302 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_decap_4 FILLER_38_369 ();
 sg13g2_fill_1 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_382 ();
 sg13g2_fill_1 FILLER_38_397 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_19 ();
 sg13g2_decap_8 FILLER_39_26 ();
 sg13g2_decap_8 FILLER_39_33 ();
 sg13g2_decap_8 FILLER_39_40 ();
 sg13g2_decap_4 FILLER_39_47 ();
 sg13g2_fill_2 FILLER_39_51 ();
 sg13g2_fill_2 FILLER_39_81 ();
 sg13g2_decap_4 FILLER_39_109 ();
 sg13g2_fill_1 FILLER_39_113 ();
 sg13g2_decap_4 FILLER_39_140 ();
 sg13g2_fill_2 FILLER_39_144 ();
 sg13g2_decap_8 FILLER_39_180 ();
 sg13g2_fill_2 FILLER_39_187 ();
 sg13g2_fill_1 FILLER_39_189 ();
 sg13g2_decap_4 FILLER_39_235 ();
 sg13g2_fill_1 FILLER_39_239 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_fill_1 FILLER_40_0 ();
 sg13g2_decap_4 FILLER_40_30 ();
 sg13g2_fill_1 FILLER_40_34 ();
 sg13g2_decap_8 FILLER_40_39 ();
 sg13g2_fill_1 FILLER_40_46 ();
 sg13g2_fill_2 FILLER_40_73 ();
 sg13g2_fill_1 FILLER_40_75 ();
 sg13g2_fill_2 FILLER_40_102 ();
 sg13g2_fill_1 FILLER_40_104 ();
 sg13g2_decap_4 FILLER_40_141 ();
 sg13g2_fill_1 FILLER_40_155 ();
 sg13g2_fill_2 FILLER_40_170 ();
 sg13g2_decap_4 FILLER_40_224 ();
 sg13g2_fill_2 FILLER_40_228 ();
 sg13g2_fill_1 FILLER_40_235 ();
 sg13g2_fill_1 FILLER_40_266 ();
 sg13g2_fill_1 FILLER_40_279 ();
 sg13g2_decap_4 FILLER_40_297 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_decap_4 FILLER_40_312 ();
 sg13g2_fill_1 FILLER_40_316 ();
 sg13g2_fill_1 FILLER_41_48 ();
 sg13g2_fill_2 FILLER_41_75 ();
 sg13g2_fill_1 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_124 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_4 FILLER_41_161 ();
 sg13g2_fill_1 FILLER_41_165 ();
 sg13g2_decap_4 FILLER_41_200 ();
 sg13g2_fill_2 FILLER_41_204 ();
 sg13g2_decap_8 FILLER_41_214 ();
 sg13g2_decap_4 FILLER_41_221 ();
 sg13g2_fill_1 FILLER_41_225 ();
 sg13g2_decap_4 FILLER_41_231 ();
 sg13g2_fill_1 FILLER_41_243 ();
 sg13g2_decap_4 FILLER_41_369 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_9 ();
 sg13g2_fill_2 FILLER_42_33 ();
 sg13g2_fill_2 FILLER_42_61 ();
 sg13g2_decap_4 FILLER_42_73 ();
 sg13g2_fill_1 FILLER_42_77 ();
 sg13g2_decap_4 FILLER_42_87 ();
 sg13g2_decap_4 FILLER_42_101 ();
 sg13g2_fill_2 FILLER_42_114 ();
 sg13g2_fill_1 FILLER_42_116 ();
 sg13g2_fill_2 FILLER_42_131 ();
 sg13g2_fill_1 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_138 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_4 FILLER_42_182 ();
 sg13g2_fill_2 FILLER_42_186 ();
 sg13g2_decap_4 FILLER_42_198 ();
 sg13g2_fill_1 FILLER_42_202 ();
 sg13g2_fill_2 FILLER_42_212 ();
 sg13g2_fill_1 FILLER_42_270 ();
 sg13g2_decap_8 FILLER_42_288 ();
 sg13g2_decap_8 FILLER_42_295 ();
 sg13g2_fill_2 FILLER_42_302 ();
 sg13g2_fill_1 FILLER_42_313 ();
 sg13g2_fill_2 FILLER_42_324 ();
 sg13g2_fill_1 FILLER_42_326 ();
 sg13g2_fill_2 FILLER_42_345 ();
 sg13g2_fill_1 FILLER_42_360 ();
 sg13g2_fill_2 FILLER_42_370 ();
 sg13g2_fill_2 FILLER_42_380 ();
 sg13g2_fill_1 FILLER_42_382 ();
 sg13g2_fill_1 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_402 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_23 ();
 sg13g2_fill_1 FILLER_43_34 ();
 sg13g2_decap_4 FILLER_43_49 ();
 sg13g2_fill_1 FILLER_43_53 ();
 sg13g2_decap_4 FILLER_43_78 ();
 sg13g2_fill_1 FILLER_43_82 ();
 sg13g2_fill_2 FILLER_43_109 ();
 sg13g2_fill_1 FILLER_43_111 ();
 sg13g2_fill_1 FILLER_43_120 ();
 sg13g2_fill_2 FILLER_43_126 ();
 sg13g2_fill_1 FILLER_43_128 ();
 sg13g2_fill_2 FILLER_43_165 ();
 sg13g2_fill_1 FILLER_43_167 ();
 sg13g2_decap_4 FILLER_43_173 ();
 sg13g2_fill_2 FILLER_43_185 ();
 sg13g2_decap_8 FILLER_43_309 ();
 sg13g2_decap_8 FILLER_43_324 ();
 sg13g2_decap_4 FILLER_43_331 ();
 sg13g2_fill_2 FILLER_43_353 ();
 sg13g2_fill_1 FILLER_43_355 ();
 sg13g2_decap_4 FILLER_43_365 ();
 sg13g2_fill_2 FILLER_43_369 ();
 sg13g2_decap_4 FILLER_43_394 ();
 sg13g2_fill_1 FILLER_43_398 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_2 ();
 sg13g2_fill_2 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_53 ();
 sg13g2_decap_8 FILLER_44_60 ();
 sg13g2_decap_4 FILLER_44_67 ();
 sg13g2_decap_8 FILLER_44_76 ();
 sg13g2_decap_8 FILLER_44_83 ();
 sg13g2_decap_8 FILLER_44_90 ();
 sg13g2_fill_1 FILLER_44_97 ();
 sg13g2_fill_2 FILLER_44_102 ();
 sg13g2_fill_2 FILLER_44_118 ();
 sg13g2_fill_1 FILLER_44_190 ();
 sg13g2_decap_8 FILLER_44_204 ();
 sg13g2_fill_2 FILLER_44_211 ();
 sg13g2_decap_4 FILLER_44_216 ();
 sg13g2_fill_2 FILLER_44_220 ();
 sg13g2_fill_2 FILLER_44_265 ();
 sg13g2_fill_1 FILLER_44_267 ();
 sg13g2_fill_2 FILLER_44_273 ();
 sg13g2_fill_1 FILLER_44_275 ();
 sg13g2_fill_1 FILLER_44_334 ();
 sg13g2_fill_2 FILLER_44_349 ();
 sg13g2_fill_1 FILLER_44_351 ();
 sg13g2_fill_2 FILLER_44_381 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_fill_2 FILLER_45_24 ();
 sg13g2_fill_1 FILLER_45_26 ();
 sg13g2_decap_8 FILLER_45_57 ();
 sg13g2_fill_1 FILLER_45_64 ();
 sg13g2_fill_2 FILLER_45_75 ();
 sg13g2_fill_1 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_fill_2 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_129 ();
 sg13g2_fill_2 FILLER_45_194 ();
 sg13g2_fill_2 FILLER_45_225 ();
 sg13g2_decap_8 FILLER_45_253 ();
 sg13g2_decap_8 FILLER_45_260 ();
 sg13g2_fill_2 FILLER_45_267 ();
 sg13g2_fill_1 FILLER_45_269 ();
 sg13g2_fill_1 FILLER_45_302 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_decap_4 FILLER_45_388 ();
 sg13g2_decap_4 FILLER_45_405 ();
 sg13g2_fill_2 FILLER_46_60 ();
 sg13g2_fill_1 FILLER_46_75 ();
 sg13g2_fill_2 FILLER_46_102 ();
 sg13g2_decap_4 FILLER_46_108 ();
 sg13g2_fill_1 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_131 ();
 sg13g2_decap_4 FILLER_46_138 ();
 sg13g2_fill_1 FILLER_46_142 ();
 sg13g2_fill_1 FILLER_46_161 ();
 sg13g2_decap_4 FILLER_46_167 ();
 sg13g2_fill_1 FILLER_46_171 ();
 sg13g2_fill_2 FILLER_46_177 ();
 sg13g2_decap_8 FILLER_46_184 ();
 sg13g2_decap_8 FILLER_46_191 ();
 sg13g2_decap_8 FILLER_46_198 ();
 sg13g2_fill_1 FILLER_46_205 ();
 sg13g2_decap_8 FILLER_46_215 ();
 sg13g2_fill_2 FILLER_46_222 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_4 FILLER_46_290 ();
 sg13g2_decap_4 FILLER_46_299 ();
 sg13g2_fill_1 FILLER_46_303 ();
 sg13g2_decap_8 FILLER_46_314 ();
 sg13g2_fill_2 FILLER_46_347 ();
 sg13g2_fill_1 FILLER_46_349 ();
 sg13g2_fill_1 FILLER_46_376 ();
 sg13g2_fill_2 FILLER_46_391 ();
 sg13g2_fill_1 FILLER_46_393 ();
 sg13g2_fill_2 FILLER_46_407 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_22 ();
 sg13g2_fill_2 FILLER_47_87 ();
 sg13g2_fill_2 FILLER_47_129 ();
 sg13g2_fill_2 FILLER_47_145 ();
 sg13g2_decap_8 FILLER_47_155 ();
 sg13g2_decap_4 FILLER_47_162 ();
 sg13g2_fill_1 FILLER_47_166 ();
 sg13g2_fill_2 FILLER_47_172 ();
 sg13g2_fill_2 FILLER_47_183 ();
 sg13g2_fill_1 FILLER_47_185 ();
 sg13g2_decap_8 FILLER_47_222 ();
 sg13g2_decap_8 FILLER_47_229 ();
 sg13g2_fill_2 FILLER_47_236 ();
 sg13g2_fill_1 FILLER_47_238 ();
 sg13g2_fill_2 FILLER_47_247 ();
 sg13g2_fill_2 FILLER_47_275 ();
 sg13g2_fill_1 FILLER_47_277 ();
 sg13g2_decap_4 FILLER_47_313 ();
 sg13g2_fill_2 FILLER_47_317 ();
 sg13g2_fill_2 FILLER_47_333 ();
 sg13g2_fill_1 FILLER_47_335 ();
 sg13g2_decap_8 FILLER_47_344 ();
 sg13g2_fill_1 FILLER_47_351 ();
 sg13g2_decap_8 FILLER_47_361 ();
 sg13g2_decap_8 FILLER_47_393 ();
 sg13g2_decap_8 FILLER_47_400 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_13 ();
 sg13g2_decap_8 FILLER_48_18 ();
 sg13g2_decap_4 FILLER_48_25 ();
 sg13g2_fill_1 FILLER_48_29 ();
 sg13g2_decap_8 FILLER_48_38 ();
 sg13g2_decap_4 FILLER_48_45 ();
 sg13g2_fill_1 FILLER_48_77 ();
 sg13g2_fill_2 FILLER_48_92 ();
 sg13g2_fill_1 FILLER_48_94 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_fill_2 FILLER_48_120 ();
 sg13g2_fill_1 FILLER_48_158 ();
 sg13g2_decap_4 FILLER_48_208 ();
 sg13g2_fill_2 FILLER_48_212 ();
 sg13g2_fill_1 FILLER_48_240 ();
 sg13g2_decap_8 FILLER_48_302 ();
 sg13g2_decap_8 FILLER_48_309 ();
 sg13g2_decap_8 FILLER_48_316 ();
 sg13g2_decap_8 FILLER_48_323 ();
 sg13g2_decap_4 FILLER_48_330 ();
 sg13g2_fill_2 FILLER_48_334 ();
 sg13g2_decap_8 FILLER_48_341 ();
 sg13g2_decap_8 FILLER_48_348 ();
 sg13g2_decap_8 FILLER_48_355 ();
 sg13g2_decap_8 FILLER_48_362 ();
 sg13g2_decap_4 FILLER_48_369 ();
 sg13g2_fill_1 FILLER_48_373 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_26 ();
 sg13g2_decap_8 FILLER_49_33 ();
 sg13g2_decap_8 FILLER_49_40 ();
 sg13g2_fill_2 FILLER_49_47 ();
 sg13g2_fill_1 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_58 ();
 sg13g2_decap_4 FILLER_49_65 ();
 sg13g2_fill_1 FILLER_49_82 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_98 ();
 sg13g2_fill_1 FILLER_49_100 ();
 sg13g2_decap_8 FILLER_49_106 ();
 sg13g2_decap_4 FILLER_49_113 ();
 sg13g2_fill_2 FILLER_49_126 ();
 sg13g2_fill_2 FILLER_49_138 ();
 sg13g2_fill_1 FILLER_49_191 ();
 sg13g2_decap_8 FILLER_49_237 ();
 sg13g2_decap_4 FILLER_49_244 ();
 sg13g2_decap_4 FILLER_49_256 ();
 sg13g2_fill_2 FILLER_49_260 ();
 sg13g2_fill_2 FILLER_49_266 ();
 sg13g2_fill_1 FILLER_49_268 ();
 sg13g2_decap_8 FILLER_49_279 ();
 sg13g2_fill_1 FILLER_49_286 ();
 sg13g2_fill_1 FILLER_49_305 ();
 sg13g2_decap_8 FILLER_49_311 ();
 sg13g2_fill_1 FILLER_49_318 ();
 sg13g2_fill_1 FILLER_49_365 ();
 sg13g2_fill_2 FILLER_49_371 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_45 ();
 sg13g2_fill_1 FILLER_50_47 ();
 sg13g2_fill_2 FILLER_50_56 ();
 sg13g2_fill_1 FILLER_50_58 ();
 sg13g2_decap_8 FILLER_50_71 ();
 sg13g2_decap_8 FILLER_50_78 ();
 sg13g2_decap_8 FILLER_50_85 ();
 sg13g2_fill_2 FILLER_50_92 ();
 sg13g2_decap_8 FILLER_50_103 ();
 sg13g2_fill_2 FILLER_50_110 ();
 sg13g2_decap_8 FILLER_50_117 ();
 sg13g2_fill_2 FILLER_50_124 ();
 sg13g2_fill_2 FILLER_50_165 ();
 sg13g2_fill_1 FILLER_50_167 ();
 sg13g2_decap_4 FILLER_50_189 ();
 sg13g2_fill_2 FILLER_50_198 ();
 sg13g2_fill_1 FILLER_50_200 ();
 sg13g2_decap_4 FILLER_50_211 ();
 sg13g2_fill_2 FILLER_50_215 ();
 sg13g2_decap_8 FILLER_50_231 ();
 sg13g2_decap_8 FILLER_50_238 ();
 sg13g2_decap_4 FILLER_50_245 ();
 sg13g2_decap_8 FILLER_50_268 ();
 sg13g2_decap_8 FILLER_50_275 ();
 sg13g2_decap_4 FILLER_50_282 ();
 sg13g2_fill_2 FILLER_50_386 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_2 ();
 sg13g2_fill_2 FILLER_51_58 ();
 sg13g2_fill_2 FILLER_51_77 ();
 sg13g2_fill_1 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_141 ();
 sg13g2_decap_8 FILLER_51_151 ();
 sg13g2_decap_8 FILLER_51_158 ();
 sg13g2_fill_2 FILLER_51_165 ();
 sg13g2_fill_1 FILLER_51_167 ();
 sg13g2_fill_2 FILLER_51_173 ();
 sg13g2_fill_1 FILLER_51_175 ();
 sg13g2_decap_8 FILLER_51_202 ();
 sg13g2_fill_2 FILLER_51_209 ();
 sg13g2_fill_1 FILLER_51_211 ();
 sg13g2_decap_8 FILLER_51_230 ();
 sg13g2_fill_1 FILLER_51_237 ();
 sg13g2_fill_2 FILLER_51_248 ();
 sg13g2_fill_1 FILLER_51_250 ();
 sg13g2_decap_8 FILLER_51_276 ();
 sg13g2_decap_4 FILLER_51_283 ();
 sg13g2_fill_2 FILLER_51_323 ();
 sg13g2_fill_1 FILLER_51_325 ();
 sg13g2_decap_4 FILLER_51_331 ();
 sg13g2_fill_2 FILLER_51_335 ();
 sg13g2_fill_2 FILLER_51_368 ();
 sg13g2_fill_1 FILLER_51_370 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_8 ();
 sg13g2_fill_2 FILLER_52_17 ();
 sg13g2_fill_1 FILLER_52_46 ();
 sg13g2_fill_2 FILLER_52_83 ();
 sg13g2_fill_1 FILLER_52_85 ();
 sg13g2_decap_8 FILLER_52_136 ();
 sg13g2_decap_8 FILLER_52_143 ();
 sg13g2_decap_4 FILLER_52_150 ();
 sg13g2_decap_8 FILLER_52_159 ();
 sg13g2_decap_8 FILLER_52_166 ();
 sg13g2_fill_1 FILLER_52_191 ();
 sg13g2_decap_4 FILLER_52_244 ();
 sg13g2_fill_2 FILLER_52_248 ();
 sg13g2_fill_2 FILLER_52_255 ();
 sg13g2_fill_1 FILLER_52_257 ();
 sg13g2_fill_1 FILLER_52_266 ();
 sg13g2_decap_8 FILLER_52_321 ();
 sg13g2_decap_8 FILLER_52_328 ();
 sg13g2_decap_8 FILLER_52_335 ();
 sg13g2_fill_2 FILLER_52_342 ();
 sg13g2_fill_1 FILLER_52_344 ();
 sg13g2_decap_4 FILLER_52_404 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_37 ();
 sg13g2_fill_1 FILLER_53_39 ();
 sg13g2_fill_1 FILLER_53_88 ();
 sg13g2_fill_1 FILLER_53_94 ();
 sg13g2_fill_2 FILLER_53_124 ();
 sg13g2_decap_8 FILLER_53_178 ();
 sg13g2_fill_2 FILLER_53_185 ();
 sg13g2_fill_2 FILLER_53_216 ();
 sg13g2_decap_8 FILLER_53_244 ();
 sg13g2_decap_4 FILLER_53_251 ();
 sg13g2_fill_1 FILLER_53_264 ();
 sg13g2_decap_4 FILLER_53_314 ();
 sg13g2_fill_1 FILLER_53_318 ();
 sg13g2_decap_4 FILLER_53_328 ();
 sg13g2_fill_2 FILLER_53_350 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_22 ();
 sg13g2_fill_2 FILLER_54_53 ();
 sg13g2_fill_1 FILLER_54_55 ();
 sg13g2_decap_8 FILLER_54_85 ();
 sg13g2_fill_2 FILLER_54_92 ();
 sg13g2_fill_1 FILLER_54_112 ();
 sg13g2_fill_1 FILLER_54_176 ();
 sg13g2_fill_2 FILLER_54_209 ();
 sg13g2_decap_8 FILLER_54_253 ();
 sg13g2_decap_8 FILLER_54_260 ();
 sg13g2_fill_1 FILLER_54_305 ();
 sg13g2_fill_2 FILLER_54_358 ();
 sg13g2_fill_1 FILLER_54_360 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_4 ();
 sg13g2_fill_2 FILLER_55_35 ();
 sg13g2_fill_1 FILLER_55_37 ();
 sg13g2_fill_1 FILLER_55_71 ();
 sg13g2_fill_2 FILLER_55_85 ();
 sg13g2_fill_2 FILLER_55_100 ();
 sg13g2_fill_1 FILLER_55_160 ();
 sg13g2_decap_4 FILLER_55_170 ();
 sg13g2_decap_8 FILLER_55_187 ();
 sg13g2_fill_1 FILLER_55_194 ();
 sg13g2_fill_1 FILLER_55_219 ();
 sg13g2_fill_2 FILLER_55_243 ();
 sg13g2_fill_1 FILLER_55_245 ();
 sg13g2_fill_2 FILLER_55_272 ();
 sg13g2_fill_1 FILLER_55_274 ();
 sg13g2_fill_1 FILLER_55_286 ();
 sg13g2_fill_1 FILLER_55_307 ();
 sg13g2_fill_1 FILLER_55_348 ();
 sg13g2_fill_2 FILLER_55_380 ();
 sg13g2_fill_1 FILLER_55_382 ();
 sg13g2_fill_1 FILLER_55_392 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_4 FILLER_56_14 ();
 sg13g2_fill_1 FILLER_56_27 ();
 sg13g2_fill_2 FILLER_56_116 ();
 sg13g2_fill_1 FILLER_56_118 ();
 sg13g2_fill_2 FILLER_56_138 ();
 sg13g2_decap_8 FILLER_56_149 ();
 sg13g2_decap_4 FILLER_56_199 ();
 sg13g2_fill_1 FILLER_56_203 ();
 sg13g2_decap_8 FILLER_56_235 ();
 sg13g2_fill_1 FILLER_56_242 ();
 sg13g2_fill_2 FILLER_56_310 ();
 sg13g2_decap_8 FILLER_56_321 ();
 sg13g2_decap_8 FILLER_56_328 ();
 sg13g2_decap_4 FILLER_56_335 ();
 sg13g2_fill_2 FILLER_56_339 ();
 sg13g2_decap_8 FILLER_56_349 ();
 sg13g2_fill_2 FILLER_56_356 ();
 sg13g2_decap_8 FILLER_56_371 ();
 sg13g2_decap_8 FILLER_56_378 ();
 sg13g2_fill_2 FILLER_56_402 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_2 ();
 sg13g2_fill_2 FILLER_57_29 ();
 sg13g2_fill_1 FILLER_57_31 ();
 sg13g2_fill_1 FILLER_57_127 ();
 sg13g2_decap_8 FILLER_57_137 ();
 sg13g2_decap_8 FILLER_57_144 ();
 sg13g2_fill_2 FILLER_57_151 ();
 sg13g2_fill_2 FILLER_57_182 ();
 sg13g2_fill_1 FILLER_57_220 ();
 sg13g2_fill_2 FILLER_57_237 ();
 sg13g2_fill_1 FILLER_57_239 ();
 sg13g2_decap_4 FILLER_57_265 ();
 sg13g2_decap_8 FILLER_57_318 ();
 sg13g2_decap_4 FILLER_57_325 ();
 sg13g2_fill_1 FILLER_57_329 ();
 sg13g2_fill_2 FILLER_57_335 ();
 sg13g2_fill_2 FILLER_57_351 ();
 sg13g2_fill_1 FILLER_57_353 ();
 sg13g2_fill_1 FILLER_57_373 ();
 sg13g2_fill_1 FILLER_57_378 ();
 sg13g2_decap_8 FILLER_57_389 ();
 sg13g2_decap_4 FILLER_57_405 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_2 ();
 sg13g2_decap_4 FILLER_58_38 ();
 sg13g2_fill_1 FILLER_58_51 ();
 sg13g2_fill_1 FILLER_58_67 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_4 FILLER_58_84 ();
 sg13g2_fill_1 FILLER_58_88 ();
 sg13g2_fill_2 FILLER_58_109 ();
 sg13g2_decap_4 FILLER_58_120 ();
 sg13g2_fill_2 FILLER_58_124 ();
 sg13g2_fill_2 FILLER_58_188 ();
 sg13g2_fill_2 FILLER_58_221 ();
 sg13g2_fill_1 FILLER_58_223 ();
 sg13g2_fill_2 FILLER_58_239 ();
 sg13g2_fill_2 FILLER_58_249 ();
 sg13g2_fill_1 FILLER_58_251 ();
 sg13g2_decap_4 FILLER_58_260 ();
 sg13g2_fill_1 FILLER_58_279 ();
 sg13g2_decap_4 FILLER_58_289 ();
 sg13g2_decap_8 FILLER_58_302 ();
 sg13g2_fill_1 FILLER_58_309 ();
 sg13g2_fill_1 FILLER_58_382 ();
 sg13g2_decap_4 FILLER_59_13 ();
 sg13g2_fill_1 FILLER_59_26 ();
 sg13g2_fill_1 FILLER_59_32 ();
 sg13g2_decap_8 FILLER_59_38 ();
 sg13g2_decap_8 FILLER_59_45 ();
 sg13g2_decap_8 FILLER_59_52 ();
 sg13g2_decap_8 FILLER_59_59 ();
 sg13g2_decap_8 FILLER_59_66 ();
 sg13g2_decap_8 FILLER_59_73 ();
 sg13g2_decap_8 FILLER_59_80 ();
 sg13g2_fill_1 FILLER_59_87 ();
 sg13g2_decap_8 FILLER_59_97 ();
 sg13g2_decap_8 FILLER_59_104 ();
 sg13g2_fill_2 FILLER_59_111 ();
 sg13g2_fill_2 FILLER_59_126 ();
 sg13g2_fill_2 FILLER_59_173 ();
 sg13g2_fill_1 FILLER_59_175 ();
 sg13g2_fill_2 FILLER_59_190 ();
 sg13g2_fill_2 FILLER_59_206 ();
 sg13g2_fill_1 FILLER_59_248 ();
 sg13g2_decap_8 FILLER_59_253 ();
 sg13g2_decap_8 FILLER_59_296 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_decap_4 FILLER_60_58 ();
 sg13g2_fill_2 FILLER_60_62 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_fill_1 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_111 ();
 sg13g2_fill_1 FILLER_60_118 ();
 sg13g2_decap_8 FILLER_60_124 ();
 sg13g2_decap_4 FILLER_60_131 ();
 sg13g2_fill_1 FILLER_60_135 ();
 sg13g2_fill_1 FILLER_60_153 ();
 sg13g2_fill_2 FILLER_60_180 ();
 sg13g2_fill_2 FILLER_60_237 ();
 sg13g2_fill_1 FILLER_60_243 ();
 sg13g2_decap_4 FILLER_60_252 ();
 sg13g2_fill_1 FILLER_60_264 ();
 sg13g2_decap_4 FILLER_60_285 ();
 sg13g2_fill_1 FILLER_60_312 ();
 sg13g2_decap_8 FILLER_60_358 ();
 sg13g2_decap_4 FILLER_60_365 ();
 sg13g2_fill_1 FILLER_60_369 ();
 sg13g2_decap_4 FILLER_60_404 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_89 ();
 sg13g2_fill_2 FILLER_61_108 ();
 sg13g2_fill_1 FILLER_61_110 ();
 sg13g2_decap_8 FILLER_61_121 ();
 sg13g2_decap_8 FILLER_61_128 ();
 sg13g2_decap_8 FILLER_61_135 ();
 sg13g2_decap_8 FILLER_61_142 ();
 sg13g2_decap_8 FILLER_61_149 ();
 sg13g2_fill_2 FILLER_61_156 ();
 sg13g2_decap_4 FILLER_61_193 ();
 sg13g2_fill_1 FILLER_61_197 ();
 sg13g2_fill_2 FILLER_61_244 ();
 sg13g2_fill_2 FILLER_61_264 ();
 sg13g2_decap_8 FILLER_61_351 ();
 sg13g2_decap_8 FILLER_61_358 ();
 sg13g2_decap_4 FILLER_61_365 ();
 sg13g2_fill_2 FILLER_61_369 ();
 sg13g2_decap_4 FILLER_61_380 ();
 sg13g2_decap_4 FILLER_61_393 ();
 sg13g2_fill_2 FILLER_61_397 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_fill_1 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_44 ();
 sg13g2_fill_1 FILLER_62_46 ();
 sg13g2_decap_4 FILLER_62_109 ();
 sg13g2_decap_8 FILLER_62_139 ();
 sg13g2_decap_8 FILLER_62_146 ();
 sg13g2_decap_8 FILLER_62_153 ();
 sg13g2_decap_8 FILLER_62_160 ();
 sg13g2_decap_4 FILLER_62_167 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_4 FILLER_62_182 ();
 sg13g2_fill_2 FILLER_62_186 ();
 sg13g2_fill_2 FILLER_62_249 ();
 sg13g2_fill_2 FILLER_62_256 ();
 sg13g2_decap_4 FILLER_62_344 ();
 sg13g2_fill_2 FILLER_62_357 ();
 sg13g2_fill_1 FILLER_62_359 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_18 ();
 sg13g2_decap_4 FILLER_63_25 ();
 sg13g2_fill_1 FILLER_63_29 ();
 sg13g2_fill_1 FILLER_63_66 ();
 sg13g2_fill_2 FILLER_63_76 ();
 sg13g2_fill_1 FILLER_63_78 ();
 sg13g2_fill_1 FILLER_63_243 ();
 sg13g2_fill_2 FILLER_63_254 ();
 sg13g2_fill_1 FILLER_63_256 ();
 sg13g2_fill_1 FILLER_63_277 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_7 ();
 sg13g2_fill_1 FILLER_64_11 ();
 sg13g2_fill_2 FILLER_64_17 ();
 sg13g2_decap_8 FILLER_64_24 ();
 sg13g2_fill_2 FILLER_64_31 ();
 sg13g2_fill_1 FILLER_64_33 ();
 sg13g2_fill_2 FILLER_64_39 ();
 sg13g2_fill_1 FILLER_64_41 ();
 sg13g2_decap_8 FILLER_64_47 ();
 sg13g2_fill_2 FILLER_64_54 ();
 sg13g2_fill_1 FILLER_64_56 ();
 sg13g2_decap_4 FILLER_64_66 ();
 sg13g2_fill_1 FILLER_64_110 ();
 sg13g2_decap_8 FILLER_64_169 ();
 sg13g2_decap_4 FILLER_64_176 ();
 sg13g2_fill_1 FILLER_64_180 ();
 sg13g2_fill_1 FILLER_64_186 ();
 sg13g2_fill_2 FILLER_64_196 ();
 sg13g2_fill_2 FILLER_64_208 ();
 sg13g2_fill_1 FILLER_64_242 ();
 sg13g2_fill_2 FILLER_64_264 ();
 sg13g2_fill_1 FILLER_64_266 ();
 sg13g2_decap_8 FILLER_64_291 ();
 sg13g2_fill_2 FILLER_64_298 ();
 sg13g2_fill_2 FILLER_64_380 ();
 sg13g2_fill_1 FILLER_64_382 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_19 ();
 sg13g2_decap_8 FILLER_65_50 ();
 sg13g2_decap_4 FILLER_65_57 ();
 sg13g2_fill_1 FILLER_65_61 ();
 sg13g2_fill_2 FILLER_65_75 ();
 sg13g2_fill_1 FILLER_65_77 ();
 sg13g2_decap_4 FILLER_65_87 ();
 sg13g2_fill_1 FILLER_65_91 ();
 sg13g2_fill_1 FILLER_65_101 ();
 sg13g2_decap_4 FILLER_65_124 ();
 sg13g2_fill_2 FILLER_65_147 ();
 sg13g2_fill_1 FILLER_65_154 ();
 sg13g2_decap_4 FILLER_65_198 ();
 sg13g2_fill_2 FILLER_65_206 ();
 sg13g2_fill_1 FILLER_65_208 ();
 sg13g2_fill_2 FILLER_65_218 ();
 sg13g2_fill_1 FILLER_65_246 ();
 sg13g2_fill_1 FILLER_65_255 ();
 sg13g2_fill_1 FILLER_65_320 ();
 sg13g2_fill_1 FILLER_65_359 ();
 sg13g2_fill_1 FILLER_65_379 ();
 sg13g2_fill_2 FILLER_65_389 ();
 sg13g2_fill_1 FILLER_65_391 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_62 ();
 sg13g2_fill_1 FILLER_66_64 ();
 sg13g2_decap_8 FILLER_66_82 ();
 sg13g2_fill_2 FILLER_66_89 ();
 sg13g2_decap_4 FILLER_66_109 ();
 sg13g2_decap_8 FILLER_66_135 ();
 sg13g2_decap_8 FILLER_66_142 ();
 sg13g2_fill_1 FILLER_66_172 ();
 sg13g2_fill_1 FILLER_66_208 ();
 sg13g2_decap_8 FILLER_66_238 ();
 sg13g2_decap_8 FILLER_66_245 ();
 sg13g2_fill_2 FILLER_66_252 ();
 sg13g2_fill_1 FILLER_66_280 ();
 sg13g2_decap_4 FILLER_66_290 ();
 sg13g2_fill_1 FILLER_66_320 ();
 sg13g2_fill_2 FILLER_66_358 ();
 sg13g2_fill_1 FILLER_66_377 ();
 sg13g2_fill_1 FILLER_66_392 ();
 sg13g2_fill_2 FILLER_66_401 ();
 sg13g2_fill_1 FILLER_66_403 ();
 sg13g2_fill_2 FILLER_67_26 ();
 sg13g2_fill_1 FILLER_67_28 ();
 sg13g2_fill_1 FILLER_67_43 ();
 sg13g2_fill_2 FILLER_67_70 ();
 sg13g2_fill_2 FILLER_67_114 ();
 sg13g2_fill_1 FILLER_67_116 ();
 sg13g2_decap_4 FILLER_67_145 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_4 FILLER_67_161 ();
 sg13g2_fill_2 FILLER_67_165 ();
 sg13g2_fill_2 FILLER_67_181 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_245 ();
 sg13g2_decap_4 FILLER_67_252 ();
 sg13g2_fill_1 FILLER_67_256 ();
 sg13g2_decap_4 FILLER_67_266 ();
 sg13g2_fill_1 FILLER_67_270 ();
 sg13g2_decap_4 FILLER_67_297 ();
 sg13g2_fill_1 FILLER_67_330 ();
 sg13g2_fill_2 FILLER_67_365 ();
 sg13g2_fill_2 FILLER_67_381 ();
 sg13g2_decap_4 FILLER_68_0 ();
 sg13g2_decap_4 FILLER_68_13 ();
 sg13g2_decap_8 FILLER_68_26 ();
 sg13g2_fill_1 FILLER_68_33 ();
 sg13g2_decap_8 FILLER_68_41 ();
 sg13g2_decap_8 FILLER_68_48 ();
 sg13g2_fill_2 FILLER_68_65 ();
 sg13g2_fill_2 FILLER_68_107 ();
 sg13g2_fill_1 FILLER_68_109 ();
 sg13g2_fill_2 FILLER_68_118 ();
 sg13g2_fill_1 FILLER_68_120 ();
 sg13g2_fill_2 FILLER_68_165 ();
 sg13g2_fill_1 FILLER_68_167 ();
 sg13g2_decap_8 FILLER_68_172 ();
 sg13g2_decap_4 FILLER_68_179 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_decap_8 FILLER_68_256 ();
 sg13g2_fill_1 FILLER_68_263 ();
 sg13g2_decap_4 FILLER_68_284 ();
 sg13g2_fill_2 FILLER_68_307 ();
 sg13g2_fill_2 FILLER_68_323 ();
 sg13g2_fill_2 FILLER_68_381 ();
 sg13g2_decap_4 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_4 ();
 sg13g2_fill_1 FILLER_69_18 ();
 sg13g2_decap_8 FILLER_69_24 ();
 sg13g2_decap_4 FILLER_69_31 ();
 sg13g2_fill_2 FILLER_69_35 ();
 sg13g2_decap_4 FILLER_69_46 ();
 sg13g2_fill_2 FILLER_69_50 ();
 sg13g2_decap_8 FILLER_69_62 ();
 sg13g2_decap_4 FILLER_69_192 ();
 sg13g2_fill_2 FILLER_69_226 ();
 sg13g2_fill_1 FILLER_69_228 ();
 sg13g2_decap_4 FILLER_69_235 ();
 sg13g2_decap_8 FILLER_69_267 ();
 sg13g2_decap_4 FILLER_69_274 ();
 sg13g2_fill_2 FILLER_69_278 ();
 sg13g2_fill_1 FILLER_69_286 ();
 sg13g2_decap_4 FILLER_69_300 ();
 sg13g2_fill_1 FILLER_69_304 ();
 sg13g2_decap_4 FILLER_69_310 ();
 sg13g2_fill_1 FILLER_69_314 ();
 sg13g2_fill_1 FILLER_69_340 ();
 sg13g2_fill_1 FILLER_69_380 ();
 sg13g2_decap_8 FILLER_69_401 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_4 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_4 ();
 sg13g2_fill_1 FILLER_70_72 ();
 sg13g2_fill_2 FILLER_70_102 ();
 sg13g2_fill_1 FILLER_70_104 ();
 sg13g2_fill_1 FILLER_70_164 ();
 sg13g2_decap_8 FILLER_70_201 ();
 sg13g2_decap_8 FILLER_70_227 ();
 sg13g2_fill_1 FILLER_70_234 ();
 sg13g2_fill_2 FILLER_70_263 ();
 sg13g2_decap_4 FILLER_70_277 ();
 sg13g2_fill_2 FILLER_70_291 ();
 sg13g2_decap_8 FILLER_70_297 ();
 sg13g2_fill_2 FILLER_70_304 ();
 sg13g2_fill_1 FILLER_70_306 ();
 sg13g2_fill_2 FILLER_70_320 ();
 sg13g2_decap_8 FILLER_70_364 ();
 sg13g2_decap_4 FILLER_70_371 ();
 sg13g2_fill_2 FILLER_70_406 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_fill_2 FILLER_71_43 ();
 sg13g2_decap_8 FILLER_71_58 ();
 sg13g2_decap_8 FILLER_71_65 ();
 sg13g2_fill_1 FILLER_71_81 ();
 sg13g2_fill_2 FILLER_71_91 ();
 sg13g2_decap_4 FILLER_71_102 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_fill_2 FILLER_71_133 ();
 sg13g2_fill_1 FILLER_71_135 ();
 sg13g2_decap_8 FILLER_71_145 ();
 sg13g2_fill_2 FILLER_71_152 ();
 sg13g2_decap_8 FILLER_71_159 ();
 sg13g2_decap_8 FILLER_71_166 ();
 sg13g2_decap_8 FILLER_71_173 ();
 sg13g2_decap_8 FILLER_71_180 ();
 sg13g2_decap_8 FILLER_71_187 ();
 sg13g2_fill_2 FILLER_71_194 ();
 sg13g2_fill_1 FILLER_71_216 ();
 sg13g2_fill_1 FILLER_71_245 ();
 sg13g2_decap_4 FILLER_71_284 ();
 sg13g2_decap_8 FILLER_71_314 ();
 sg13g2_fill_1 FILLER_71_321 ();
 sg13g2_fill_2 FILLER_71_334 ();
 sg13g2_decap_8 FILLER_71_360 ();
 sg13g2_fill_2 FILLER_71_367 ();
 sg13g2_fill_1 FILLER_71_369 ();
 sg13g2_fill_1 FILLER_71_384 ();
 sg13g2_fill_2 FILLER_71_395 ();
 sg13g2_fill_2 FILLER_71_406 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_30 ();
 sg13g2_fill_1 FILLER_72_58 ();
 sg13g2_decap_8 FILLER_72_117 ();
 sg13g2_decap_8 FILLER_72_124 ();
 sg13g2_fill_1 FILLER_72_131 ();
 sg13g2_fill_1 FILLER_72_140 ();
 sg13g2_decap_4 FILLER_72_151 ();
 sg13g2_fill_1 FILLER_72_155 ();
 sg13g2_fill_2 FILLER_72_165 ();
 sg13g2_fill_1 FILLER_72_167 ();
 sg13g2_decap_4 FILLER_72_173 ();
 sg13g2_fill_1 FILLER_72_177 ();
 sg13g2_fill_2 FILLER_72_204 ();
 sg13g2_fill_1 FILLER_72_206 ();
 sg13g2_decap_4 FILLER_72_246 ();
 sg13g2_fill_1 FILLER_72_250 ();
 sg13g2_decap_4 FILLER_72_321 ();
 sg13g2_fill_2 FILLER_72_325 ();
 sg13g2_fill_2 FILLER_72_348 ();
 sg13g2_fill_2 FILLER_72_381 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_92 ();
 sg13g2_fill_1 FILLER_73_119 ();
 sg13g2_fill_2 FILLER_73_128 ();
 sg13g2_fill_1 FILLER_73_130 ();
 sg13g2_decap_8 FILLER_73_245 ();
 sg13g2_decap_8 FILLER_73_252 ();
 sg13g2_fill_1 FILLER_73_259 ();
 sg13g2_fill_1 FILLER_73_273 ();
 sg13g2_fill_1 FILLER_73_285 ();
 sg13g2_fill_2 FILLER_73_300 ();
 sg13g2_fill_1 FILLER_73_302 ();
 sg13g2_fill_2 FILLER_73_376 ();
 sg13g2_fill_2 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_33 ();
 sg13g2_fill_2 FILLER_74_71 ();
 sg13g2_fill_1 FILLER_74_151 ();
 sg13g2_fill_2 FILLER_74_210 ();
 sg13g2_fill_1 FILLER_74_212 ();
 sg13g2_fill_1 FILLER_74_218 ();
 sg13g2_fill_2 FILLER_74_259 ();
 sg13g2_fill_1 FILLER_74_261 ();
 sg13g2_decap_4 FILLER_74_279 ();
 sg13g2_decap_8 FILLER_74_312 ();
 sg13g2_fill_2 FILLER_74_351 ();
 sg13g2_decap_4 FILLER_74_361 ();
 sg13g2_fill_1 FILLER_74_365 ();
 sg13g2_fill_2 FILLER_74_381 ();
 sg13g2_fill_2 FILLER_75_26 ();
 sg13g2_decap_8 FILLER_75_44 ();
 sg13g2_decap_8 FILLER_75_51 ();
 sg13g2_decap_4 FILLER_75_58 ();
 sg13g2_fill_1 FILLER_75_62 ();
 sg13g2_fill_1 FILLER_75_72 ();
 sg13g2_fill_1 FILLER_75_87 ();
 sg13g2_decap_4 FILLER_75_108 ();
 sg13g2_fill_2 FILLER_75_112 ();
 sg13g2_fill_1 FILLER_75_139 ();
 sg13g2_decap_4 FILLER_75_164 ();
 sg13g2_fill_2 FILLER_75_168 ();
 sg13g2_fill_2 FILLER_75_186 ();
 sg13g2_fill_1 FILLER_75_207 ();
 sg13g2_decap_8 FILLER_75_213 ();
 sg13g2_fill_1 FILLER_75_220 ();
 sg13g2_decap_4 FILLER_75_252 ();
 sg13g2_fill_2 FILLER_75_256 ();
 sg13g2_fill_2 FILLER_75_319 ();
 sg13g2_fill_1 FILLER_75_321 ();
 sg13g2_fill_1 FILLER_75_328 ();
 sg13g2_fill_2 FILLER_75_359 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_fill_2 FILLER_75_380 ();
 sg13g2_fill_1 FILLER_75_382 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_decap_4 FILLER_76_34 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_fill_2 FILLER_76_60 ();
 sg13g2_fill_1 FILLER_76_62 ();
 sg13g2_fill_2 FILLER_76_93 ();
 sg13g2_fill_1 FILLER_76_95 ();
 sg13g2_decap_4 FILLER_76_114 ();
 sg13g2_fill_2 FILLER_76_118 ();
 sg13g2_decap_4 FILLER_76_141 ();
 sg13g2_decap_8 FILLER_76_149 ();
 sg13g2_fill_1 FILLER_76_156 ();
 sg13g2_fill_2 FILLER_76_161 ();
 sg13g2_fill_1 FILLER_76_163 ();
 sg13g2_decap_8 FILLER_76_180 ();
 sg13g2_fill_1 FILLER_76_187 ();
 sg13g2_fill_1 FILLER_76_193 ();
 sg13g2_decap_4 FILLER_76_213 ();
 sg13g2_fill_2 FILLER_76_239 ();
 sg13g2_fill_2 FILLER_76_318 ();
 sg13g2_fill_2 FILLER_76_334 ();
 sg13g2_fill_2 FILLER_76_345 ();
 sg13g2_fill_1 FILLER_76_356 ();
 sg13g2_fill_2 FILLER_76_366 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_7 ();
 sg13g2_decap_4 FILLER_77_16 ();
 sg13g2_fill_1 FILLER_77_77 ();
 sg13g2_fill_2 FILLER_77_104 ();
 sg13g2_fill_1 FILLER_77_106 ();
 sg13g2_fill_2 FILLER_77_125 ();
 sg13g2_fill_2 FILLER_77_213 ();
 sg13g2_fill_1 FILLER_77_215 ();
 sg13g2_fill_2 FILLER_77_251 ();
 sg13g2_fill_1 FILLER_77_253 ();
 sg13g2_fill_1 FILLER_77_258 ();
 sg13g2_fill_2 FILLER_77_266 ();
 sg13g2_fill_1 FILLER_77_268 ();
 sg13g2_fill_1 FILLER_77_283 ();
 sg13g2_fill_2 FILLER_77_310 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_fill_1 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_fill_1 FILLER_78_35 ();
 sg13g2_fill_1 FILLER_78_93 ();
 sg13g2_fill_1 FILLER_78_125 ();
 sg13g2_fill_2 FILLER_78_304 ();
 sg13g2_fill_1 FILLER_78_306 ();
 sg13g2_decap_8 FILLER_78_373 ();
 sg13g2_decap_8 FILLER_78_380 ();
 sg13g2_decap_8 FILLER_78_387 ();
 sg13g2_decap_8 FILLER_78_394 ();
 sg13g2_decap_8 FILLER_78_401 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_4 FILLER_79_28 ();
 sg13g2_fill_1 FILLER_79_32 ();
 sg13g2_fill_1 FILLER_79_71 ();
 sg13g2_fill_2 FILLER_79_104 ();
 sg13g2_fill_1 FILLER_79_106 ();
 sg13g2_decap_4 FILLER_79_169 ();
 sg13g2_fill_2 FILLER_79_209 ();
 sg13g2_fill_1 FILLER_79_211 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_fill_1 FILLER_79_245 ();
 sg13g2_fill_2 FILLER_79_347 ();
 sg13g2_decap_8 FILLER_79_375 ();
 sg13g2_decap_8 FILLER_79_382 ();
 sg13g2_decap_8 FILLER_79_389 ();
 sg13g2_decap_8 FILLER_79_396 ();
 sg13g2_decap_4 FILLER_79_403 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_4 FILLER_80_21 ();
 sg13g2_fill_2 FILLER_80_25 ();
 sg13g2_fill_1 FILLER_80_81 ();
 sg13g2_fill_1 FILLER_80_121 ();
 sg13g2_fill_1 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_187 ();
 sg13g2_fill_2 FILLER_80_195 ();
 sg13g2_fill_1 FILLER_80_197 ();
 sg13g2_decap_8 FILLER_80_211 ();
 sg13g2_decap_4 FILLER_80_218 ();
 sg13g2_decap_8 FILLER_80_240 ();
 sg13g2_decap_8 FILLER_80_247 ();
 sg13g2_decap_8 FILLER_80_254 ();
 sg13g2_decap_8 FILLER_80_261 ();
 sg13g2_decap_8 FILLER_80_268 ();
 sg13g2_fill_1 FILLER_80_275 ();
 sg13g2_fill_2 FILLER_80_279 ();
 sg13g2_decap_4 FILLER_80_308 ();
 sg13g2_decap_4 FILLER_80_317 ();
 sg13g2_fill_1 FILLER_80_321 ();
 sg13g2_decap_8 FILLER_80_326 ();
 sg13g2_decap_4 FILLER_80_333 ();
 sg13g2_decap_8 FILLER_80_375 ();
 sg13g2_decap_8 FILLER_80_382 ();
 sg13g2_decap_8 FILLER_80_389 ();
 sg13g2_decap_8 FILLER_80_396 ();
 sg13g2_decap_4 FILLER_80_403 ();
 sg13g2_fill_2 FILLER_80_407 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
endmodule
