VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_pwm_block
  CLASS BLOCK ;
  FOREIGN tt_um_pwm_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 202.080 BY 313.740 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 21.580 3.560 23.780 310.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 60.450 3.560 62.650 310.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 99.320 3.560 101.520 310.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 138.190 3.560 140.390 310.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 177.060 3.560 179.260 310.180 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 15.380 3.560 17.580 310.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 54.250 3.560 56.450 310.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 93.120 3.560 95.320 310.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 131.990 3.560 134.190 310.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 170.860 3.560 173.060 310.180 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.646800 ;
    ANTENNADIFFAREA 8.061600 ;
    PORT
      LAYER Metal5 ;
        RECT 187.050 312.740 187.350 313.740 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 190.890 312.740 191.190 313.740 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.314600 ;
    PORT
      LAYER Metal5 ;
        RECT 183.210 312.740 183.510 313.740 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 179.370 312.740 179.670 313.740 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.530 312.740 175.830 313.740 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 171.690 312.740 171.990 313.740 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 167.850 312.740 168.150 313.740 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 164.010 312.740 164.310 313.740 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 160.170 312.740 160.470 313.740 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 156.330 312.740 156.630 313.740 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 152.490 312.740 152.790 313.740 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 148.650 312.740 148.950 313.740 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 144.810 312.740 145.110 313.740 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 140.970 312.740 141.270 313.740 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 137.130 312.740 137.430 313.740 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal5 ;
        RECT 133.290 312.740 133.590 313.740 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 129.450 312.740 129.750 313.740 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal5 ;
        RECT 125.610 312.740 125.910 313.740 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495300 ;
    PORT
      LAYER Metal5 ;
        RECT 121.770 312.740 122.070 313.740 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal5 ;
        RECT 56.490 312.740 56.790 313.740 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal5 ;
        RECT 52.650 312.740 52.950 313.740 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal5 ;
        RECT 48.810 312.740 49.110 313.740 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal5 ;
        RECT 44.970 312.740 45.270 313.740 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 41.130 312.740 41.430 313.740 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal5 ;
        RECT 37.290 312.740 37.590 313.740 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 33.450 312.740 33.750 313.740 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 29.610 312.740 29.910 313.740 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 87.210 312.740 87.510 313.740 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 83.370 312.740 83.670 313.740 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 79.530 312.740 79.830 313.740 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 75.690 312.740 75.990 313.740 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 71.850 312.740 72.150 313.740 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 68.010 312.740 68.310 313.740 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 64.170 312.740 64.470 313.740 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 60.330 312.740 60.630 313.740 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal5 ;
        RECT 117.930 312.740 118.230 313.740 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal5 ;
        RECT 114.090 312.740 114.390 313.740 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal5 ;
        RECT 110.250 312.740 110.550 313.740 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 106.410 312.740 106.710 313.740 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 102.570 312.740 102.870 313.740 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 98.730 312.740 99.030 313.740 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 94.890 312.740 95.190 313.740 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal5 ;
        RECT 91.050 312.740 91.350 313.740 ;
    END
  END uo_out[7]
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 199.200 310.110 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 199.200 310.180 ;
      LAYER Metal2 ;
        RECT 2.605 2.840 200.785 310.060 ;
      LAYER Metal3 ;
        RECT 3.260 2.795 200.740 312.625 ;
      LAYER Metal4 ;
        RECT 6.575 3.680 198.865 312.580 ;
      LAYER Metal5 ;
        RECT 14.780 312.530 29.400 312.740 ;
        RECT 30.120 312.530 33.240 312.740 ;
        RECT 33.960 312.530 37.080 312.740 ;
        RECT 37.800 312.530 40.920 312.740 ;
        RECT 41.640 312.530 44.760 312.740 ;
        RECT 45.480 312.530 48.600 312.740 ;
        RECT 49.320 312.530 52.440 312.740 ;
        RECT 53.160 312.530 56.280 312.740 ;
        RECT 57.000 312.530 60.120 312.740 ;
        RECT 60.840 312.530 63.960 312.740 ;
        RECT 64.680 312.530 67.800 312.740 ;
        RECT 68.520 312.530 71.640 312.740 ;
        RECT 72.360 312.530 75.480 312.740 ;
        RECT 76.200 312.530 79.320 312.740 ;
        RECT 80.040 312.530 83.160 312.740 ;
        RECT 83.880 312.530 87.000 312.740 ;
        RECT 87.720 312.530 90.840 312.740 ;
        RECT 91.560 312.530 94.680 312.740 ;
        RECT 95.400 312.530 98.520 312.740 ;
        RECT 99.240 312.530 102.360 312.740 ;
        RECT 103.080 312.530 106.200 312.740 ;
        RECT 106.920 312.530 110.040 312.740 ;
        RECT 110.760 312.530 113.880 312.740 ;
        RECT 114.600 312.530 117.720 312.740 ;
        RECT 118.440 312.530 121.560 312.740 ;
        RECT 122.280 312.530 125.400 312.740 ;
        RECT 126.120 312.530 129.240 312.740 ;
        RECT 129.960 312.530 133.080 312.740 ;
        RECT 133.800 312.530 136.920 312.740 ;
        RECT 137.640 312.530 140.760 312.740 ;
        RECT 141.480 312.530 144.600 312.740 ;
        RECT 145.320 312.530 148.440 312.740 ;
        RECT 149.160 312.530 152.280 312.740 ;
        RECT 153.000 312.530 156.120 312.740 ;
        RECT 156.840 312.530 159.960 312.740 ;
        RECT 160.680 312.530 163.800 312.740 ;
        RECT 164.520 312.530 167.640 312.740 ;
        RECT 168.360 312.530 171.480 312.740 ;
        RECT 172.200 312.530 175.320 312.740 ;
        RECT 176.040 312.530 179.160 312.740 ;
        RECT 179.880 312.530 183.000 312.740 ;
        RECT 183.720 312.530 186.840 312.740 ;
        RECT 187.560 312.530 190.680 312.740 ;
        RECT 191.400 312.530 196.420 312.740 ;
        RECT 14.780 310.390 196.420 312.530 ;
        RECT 14.780 5.735 15.170 310.390 ;
        RECT 17.790 5.735 21.370 310.390 ;
        RECT 23.990 5.735 54.040 310.390 ;
        RECT 56.660 5.735 60.240 310.390 ;
        RECT 62.860 5.735 92.910 310.390 ;
        RECT 95.530 5.735 99.110 310.390 ;
        RECT 101.730 5.735 131.780 310.390 ;
        RECT 134.400 5.735 137.980 310.390 ;
        RECT 140.600 5.735 170.650 310.390 ;
        RECT 173.270 5.735 176.850 310.390 ;
        RECT 179.470 5.735 196.420 310.390 ;
  END
END tt_um_pwm_block
END LIBRARY

