module tt_um_abhinav8prasad_dds (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire \accum.PHASE_INC[0] ;
 wire \accum.PHASE_INC[1] ;
 wire \accum.PHASE_INC[2] ;
 wire \accum.PHASE_INC[3] ;
 wire \accum.PHASE_INC[4] ;
 wire \accum.PHASE_INC[5] ;
 wire \accum.PHASE_INC[6] ;
 wire \accum.PHASE_INC[7] ;
 wire \accum.addr[0] ;
 wire \accum.addr[1] ;
 wire \accum.addr[2] ;
 wire \accum.addr[3] ;
 wire \accum.addr[4] ;
 wire \accum.addr[5] ;
 wire \accum.addr[6] ;
 wire \accum.addr[7] ;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire clknet_0_clk;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;

 sg13g2_inv_2 _328_ (.Y(_280_),
    .A(\accum.addr[7] ));
 sg13g2_inv_1 _329_ (.Y(_281_),
    .A(net142));
 sg13g2_inv_2 _330_ (.Y(_282_),
    .A(net159));
 sg13g2_inv_1 _331_ (.Y(_283_),
    .A(net164));
 sg13g2_inv_2 _332_ (.Y(_284_),
    .A(net162));
 sg13g2_inv_1 _333_ (.Y(_285_),
    .A(net157));
 sg13g2_inv_1 _334_ (.Y(_286_),
    .A(_003_));
 sg13g2_nor2_2 _335_ (.A(net137),
    .B(net140),
    .Y(_287_));
 sg13g2_nand2_1 _336_ (.Y(_288_),
    .A(net159),
    .B(_007_));
 sg13g2_nor2_2 _337_ (.A(net158),
    .B(net164),
    .Y(_289_));
 sg13g2_nor2b_2 _338_ (.A(net165),
    .B_N(net163),
    .Y(_290_));
 sg13g2_a21oi_1 _339_ (.A1(net162),
    .A2(_289_),
    .Y(_291_),
    .B1(net153));
 sg13g2_nand2_1 _340_ (.Y(_292_),
    .A(net153),
    .B(net159));
 sg13g2_nand2_1 _341_ (.Y(_293_),
    .A(net164),
    .B(_284_));
 sg13g2_nand2_2 _342_ (.Y(_294_),
    .A(net155),
    .B(net165));
 sg13g2_inv_1 _343_ (.Y(_295_),
    .A(_294_));
 sg13g2_o21ai_1 _344_ (.B1(_292_),
    .Y(_296_),
    .A1(net162),
    .A2(_294_));
 sg13g2_nand2_2 _345_ (.Y(_297_),
    .A(net158),
    .B(net162));
 sg13g2_o21ai_1 _346_ (.B1(_296_),
    .Y(_298_),
    .A1(net165),
    .A2(_297_));
 sg13g2_nand2_1 _347_ (.Y(_299_),
    .A(net132),
    .B(_298_));
 sg13g2_a21oi_1 _348_ (.A1(_288_),
    .A2(_291_),
    .Y(_300_),
    .B1(_299_));
 sg13g2_xor2_1 _349_ (.B(\accum.addr[1] ),
    .A(net166),
    .X(_301_));
 sg13g2_and2_2 _350_ (.A(net147),
    .B(net156),
    .X(_302_));
 sg13g2_nand2_2 _351_ (.Y(_303_),
    .A(net142),
    .B(net150));
 sg13g2_nand2_2 _352_ (.Y(_304_),
    .A(net159),
    .B(net165));
 sg13g2_nand3b_1 _353_ (.B(_302_),
    .C(_304_),
    .Y(_305_),
    .A_N(_301_));
 sg13g2_nor2_2 _354_ (.A(net133),
    .B(net155),
    .Y(_306_));
 sg13g2_nand2b_2 _355_ (.Y(_307_),
    .B(net142),
    .A_N(net150));
 sg13g2_nor2_1 _356_ (.A(_282_),
    .B(_290_),
    .Y(_308_));
 sg13g2_nor2b_1 _357_ (.A(net159),
    .B_N(_007_),
    .Y(_309_));
 sg13g2_nand2_1 _358_ (.Y(_310_),
    .A(_282_),
    .B(_007_));
 sg13g2_nor2_1 _359_ (.A(_308_),
    .B(_309_),
    .Y(_311_));
 sg13g2_nand2_1 _360_ (.Y(_312_),
    .A(net164),
    .B(net162));
 sg13g2_nor2_1 _361_ (.A(net158),
    .B(net130),
    .Y(_313_));
 sg13g2_nor2_1 _362_ (.A(net164),
    .B(net162),
    .Y(_314_));
 sg13g2_nand2_2 _363_ (.Y(_315_),
    .A(_283_),
    .B(_284_));
 sg13g2_o21ai_1 _364_ (.B1(_305_),
    .Y(_316_),
    .A1(_307_),
    .A2(_311_));
 sg13g2_o21ai_1 _365_ (.B1(_287_),
    .Y(_317_),
    .A1(_300_),
    .A2(_316_));
 sg13g2_or2_2 _366_ (.X(_318_),
    .B(net163),
    .A(net160));
 sg13g2_nand2_2 _367_ (.Y(_319_),
    .A(_282_),
    .B(_301_));
 sg13g2_nand2b_1 _368_ (.Y(_320_),
    .B(_319_),
    .A_N(_308_));
 sg13g2_nor2b_2 _369_ (.A(net158),
    .B_N(net151),
    .Y(_025_));
 sg13g2_nor2b_1 _370_ (.A(net130),
    .B_N(_025_),
    .Y(_026_));
 sg13g2_a21oi_1 _371_ (.A1(_294_),
    .A2(_320_),
    .Y(_027_),
    .B1(_026_));
 sg13g2_nor2_1 _372_ (.A(net146),
    .B(net149),
    .Y(_028_));
 sg13g2_nor2b_1 _373_ (.A(net135),
    .B_N(net139),
    .Y(_029_));
 sg13g2_nand2b_1 _374_ (.Y(_030_),
    .B(net140),
    .A_N(net136));
 sg13g2_a221oi_1 _375_ (.B2(_301_),
    .C1(_030_),
    .B1(_028_),
    .A1(net146),
    .Y(_031_),
    .A2(_027_));
 sg13g2_nor2_1 _376_ (.A(_292_),
    .B(_293_),
    .Y(_032_));
 sg13g2_nand2_1 _377_ (.Y(_033_),
    .A(net159),
    .B(net131));
 sg13g2_a21oi_1 _378_ (.A1(_294_),
    .A2(_033_),
    .Y(_034_),
    .B1(_032_));
 sg13g2_nor2_1 _379_ (.A(net145),
    .B(_034_),
    .Y(_035_));
 sg13g2_nor2b_2 _380_ (.A(net141),
    .B_N(net136),
    .Y(_036_));
 sg13g2_nand2b_2 _381_ (.Y(_037_),
    .B(net136),
    .A_N(net140));
 sg13g2_nand2_2 _382_ (.Y(_038_),
    .A(net158),
    .B(_006_));
 sg13g2_o21ai_1 _383_ (.B1(_038_),
    .Y(_039_),
    .A1(_283_),
    .A2(_318_));
 sg13g2_o21ai_1 _384_ (.B1(_036_),
    .Y(_040_),
    .A1(_307_),
    .A2(_039_));
 sg13g2_nor2_1 _385_ (.A(net159),
    .B(_290_),
    .Y(_041_));
 sg13g2_o21ai_1 _386_ (.B1(_288_),
    .Y(_042_),
    .A1(net159),
    .A2(_290_));
 sg13g2_and2_1 _387_ (.A(net155),
    .B(_042_),
    .X(_043_));
 sg13g2_nor2_1 _388_ (.A(net154),
    .B(net158),
    .Y(_044_));
 sg13g2_nor2_1 _389_ (.A(net164),
    .B(_318_),
    .Y(_045_));
 sg13g2_nand2_2 _390_ (.Y(_046_),
    .A(_284_),
    .B(_289_));
 sg13g2_nor2_1 _391_ (.A(net152),
    .B(_046_),
    .Y(_047_));
 sg13g2_nor2_1 _392_ (.A(net144),
    .B(_047_),
    .Y(_048_));
 sg13g2_o21ai_1 _393_ (.B1(net133),
    .Y(_049_),
    .A1(net154),
    .A2(_046_));
 sg13g2_nor2_1 _394_ (.A(net153),
    .B(_282_),
    .Y(_050_));
 sg13g2_nor2_1 _395_ (.A(net152),
    .B(_038_),
    .Y(_051_));
 sg13g2_nor3_1 _396_ (.A(_043_),
    .B(_049_),
    .C(_051_),
    .Y(_052_));
 sg13g2_and2_2 _397_ (.A(net137),
    .B(net140),
    .X(_053_));
 sg13g2_nand2_2 _398_ (.Y(_054_),
    .A(net135),
    .B(net139));
 sg13g2_o21ai_1 _399_ (.B1(_053_),
    .Y(_055_),
    .A1(_007_),
    .A2(_303_));
 sg13g2_nor2_1 _400_ (.A(_314_),
    .B(_033_),
    .Y(_056_));
 sg13g2_nand2_2 _401_ (.Y(_057_),
    .A(net160),
    .B(_301_));
 sg13g2_nor3_1 _402_ (.A(_307_),
    .B(_309_),
    .C(_056_),
    .Y(_058_));
 sg13g2_nor3_1 _403_ (.A(_052_),
    .B(_055_),
    .C(_058_),
    .Y(_059_));
 sg13g2_o21ai_1 _404_ (.B1(net134),
    .Y(_060_),
    .A1(_035_),
    .A2(_040_));
 sg13g2_nor3_1 _405_ (.A(_031_),
    .B(_059_),
    .C(_060_),
    .Y(_061_));
 sg13g2_nand2b_2 _406_ (.Y(_062_),
    .B(_006_),
    .A_N(net160));
 sg13g2_nand3_1 _407_ (.B(_304_),
    .C(_062_),
    .A(_297_),
    .Y(_063_));
 sg13g2_a22oi_1 _408_ (.Y(_064_),
    .B1(_063_),
    .B2(_302_),
    .A2(_028_),
    .A1(_301_));
 sg13g2_o21ai_1 _409_ (.B1(_064_),
    .Y(_065_),
    .A1(_307_),
    .A2(_320_));
 sg13g2_nor2b_2 _410_ (.A(_289_),
    .B_N(_304_),
    .Y(_066_));
 sg13g2_nand2b_2 _411_ (.Y(_067_),
    .B(net143),
    .A_N(net138));
 sg13g2_nor3_1 _412_ (.A(net129),
    .B(_026_),
    .C(_067_),
    .Y(_068_));
 sg13g2_o21ai_1 _413_ (.B1(_068_),
    .Y(_069_),
    .A1(net153),
    .A2(_066_));
 sg13g2_nand2b_1 _414_ (.Y(_070_),
    .B(net164),
    .A_N(net150));
 sg13g2_or2_2 _415_ (.X(_071_),
    .B(net143),
    .A(net138));
 sg13g2_a21oi_1 _416_ (.A1(_298_),
    .A2(_070_),
    .Y(_072_),
    .B1(_071_));
 sg13g2_a21oi_1 _417_ (.A1(net139),
    .A2(_065_),
    .Y(_073_),
    .B1(_072_));
 sg13g2_a21oi_1 _418_ (.A1(_069_),
    .A2(_073_),
    .Y(_074_),
    .B1(net135));
 sg13g2_nand2_2 _419_ (.Y(_075_),
    .A(net150),
    .B(_318_));
 sg13g2_nor2_1 _420_ (.A(_066_),
    .B(_075_),
    .Y(_076_));
 sg13g2_nor2_1 _421_ (.A(net145),
    .B(_076_),
    .Y(_077_));
 sg13g2_nor2b_1 _422_ (.A(net129),
    .B_N(_044_),
    .Y(_078_));
 sg13g2_nor2_1 _423_ (.A(net151),
    .B(_297_),
    .Y(_079_));
 sg13g2_nor4_1 _424_ (.A(net144),
    .B(_076_),
    .C(_078_),
    .D(_079_),
    .Y(_080_));
 sg13g2_nor2_1 _425_ (.A(net150),
    .B(_289_),
    .Y(_081_));
 sg13g2_a221oi_1 _426_ (.B2(_081_),
    .C1(net132),
    .B1(_057_),
    .A1(net153),
    .Y(_082_),
    .A2(net164));
 sg13g2_nor3_1 _427_ (.A(_054_),
    .B(_080_),
    .C(_082_),
    .Y(_083_));
 sg13g2_o21ai_1 _428_ (.B1(_306_),
    .Y(_084_),
    .A1(net162),
    .A2(_289_));
 sg13g2_nor2_2 _429_ (.A(net150),
    .B(net157),
    .Y(_085_));
 sg13g2_nand2_1 _430_ (.Y(_086_),
    .A(net130),
    .B(_085_));
 sg13g2_a22oi_1 _431_ (.Y(_087_),
    .B1(net131),
    .B2(_085_),
    .A2(_310_),
    .A1(net153));
 sg13g2_o21ai_1 _432_ (.B1(net132),
    .Y(_088_),
    .A1(_032_),
    .A2(_087_));
 sg13g2_a21oi_1 _433_ (.A1(_084_),
    .A2(_088_),
    .Y(_089_),
    .B1(_037_));
 sg13g2_nor4_1 _434_ (.A(net134),
    .B(_074_),
    .C(_083_),
    .D(_089_),
    .Y(_090_));
 sg13g2_a21oi_2 _435_ (.B1(_090_),
    .Y(uo_out[0]),
    .A2(_061_),
    .A1(_317_));
 sg13g2_nand2b_1 _436_ (.Y(_091_),
    .B(_284_),
    .A_N(_070_));
 sg13g2_nand4_1 _437_ (.B(_075_),
    .C(_086_),
    .A(net142),
    .Y(_092_),
    .D(_091_));
 sg13g2_nor2b_2 _438_ (.A(net147),
    .B_N(net155),
    .Y(_093_));
 sg13g2_nand2_1 _439_ (.Y(_094_),
    .A(net132),
    .B(net150));
 sg13g2_xnor2_1 _440_ (.Y(_095_),
    .A(net160),
    .B(_290_));
 sg13g2_nor2_1 _441_ (.A(_094_),
    .B(_095_),
    .Y(_096_));
 sg13g2_o21ai_1 _442_ (.B1(_092_),
    .Y(_097_),
    .A1(net142),
    .A2(_070_));
 sg13g2_o21ai_1 _443_ (.B1(_029_),
    .Y(_098_),
    .A1(_096_),
    .A2(_097_));
 sg13g2_nand2_1 _444_ (.Y(_099_),
    .A(_057_),
    .B(_062_));
 sg13g2_nor2_2 _445_ (.A(net147),
    .B(net156),
    .Y(_100_));
 sg13g2_inv_2 _446_ (.Y(_101_),
    .A(_100_));
 sg13g2_nor3_1 _447_ (.A(_005_),
    .B(net131),
    .C(_101_),
    .Y(_102_));
 sg13g2_a21o_1 _448_ (.A2(_042_),
    .A1(_306_),
    .B1(_102_),
    .X(_103_));
 sg13g2_a221oi_1 _449_ (.B2(_099_),
    .C1(_103_),
    .B1(_093_),
    .A1(net146),
    .Y(_104_),
    .A2(_295_));
 sg13g2_nor3_1 _450_ (.A(_041_),
    .B(_056_),
    .C(_101_),
    .Y(_105_));
 sg13g2_mux2_1 _451_ (.A0(_006_),
    .A1(net129),
    .S(_050_),
    .X(_106_));
 sg13g2_nand2_1 _452_ (.Y(_107_),
    .A(_319_),
    .B(_038_));
 sg13g2_a221oi_1 _453_ (.B2(_093_),
    .C1(_105_),
    .B1(_107_),
    .A1(net148),
    .Y(_108_),
    .A2(_106_));
 sg13g2_o21ai_1 _454_ (.B1(_288_),
    .Y(_109_),
    .A1(_283_),
    .A2(_318_));
 sg13g2_nand2_1 _455_ (.Y(_110_),
    .A(_291_),
    .B(_293_));
 sg13g2_nand2_1 _456_ (.Y(_111_),
    .A(net145),
    .B(_110_));
 sg13g2_nand3_1 _457_ (.B(net166),
    .C(\accum.addr[1] ),
    .A(net160),
    .Y(_112_));
 sg13g2_nor3_1 _458_ (.A(net144),
    .B(net129),
    .C(_044_),
    .Y(_113_));
 sg13g2_nand2_2 _459_ (.Y(_114_),
    .A(_282_),
    .B(net131));
 sg13g2_a21oi_1 _460_ (.A1(net166),
    .A2(net163),
    .Y(_115_),
    .B1(net160));
 sg13g2_nor2_1 _461_ (.A(_101_),
    .B(_114_),
    .Y(_116_));
 sg13g2_a21oi_1 _462_ (.A1(_112_),
    .A2(_113_),
    .Y(_117_),
    .B1(_116_));
 sg13g2_a22oi_1 _463_ (.Y(_118_),
    .B1(_111_),
    .B2(_117_),
    .A2(_109_),
    .A1(_302_));
 sg13g2_nand2b_1 _464_ (.Y(_119_),
    .B(_287_),
    .A_N(_118_));
 sg13g2_o21ai_1 _465_ (.B1(\accum.addr[7] ),
    .Y(_120_),
    .A1(_037_),
    .A2(_104_));
 sg13g2_o21ai_1 _466_ (.B1(_098_),
    .Y(_121_),
    .A1(_054_),
    .A2(_108_));
 sg13g2_nor2_1 _467_ (.A(_120_),
    .B(_121_),
    .Y(_122_));
 sg13g2_nor2_1 _468_ (.A(net130),
    .B(_025_),
    .Y(_123_));
 sg13g2_nor3_1 _469_ (.A(net129),
    .B(_071_),
    .C(_123_),
    .Y(_124_));
 sg13g2_o21ai_1 _470_ (.B1(_081_),
    .Y(_125_),
    .A1(_283_),
    .A2(_006_));
 sg13g2_nand3_1 _471_ (.B(_075_),
    .C(_125_),
    .A(net145),
    .Y(_126_));
 sg13g2_o21ai_1 _472_ (.B1(net139),
    .Y(_127_),
    .A1(_007_),
    .A2(_101_));
 sg13g2_nor2_1 _473_ (.A(_096_),
    .B(_127_),
    .Y(_128_));
 sg13g2_nand3_1 _474_ (.B(_057_),
    .C(_093_),
    .A(_318_),
    .Y(_129_));
 sg13g2_nand2_2 _475_ (.Y(_130_),
    .A(net142),
    .B(_318_));
 sg13g2_nor3_1 _476_ (.A(net155),
    .B(_066_),
    .C(_130_),
    .Y(_131_));
 sg13g2_a221oi_1 _477_ (.B2(_112_),
    .C1(_131_),
    .B1(_100_),
    .A1(_007_),
    .Y(_132_),
    .A2(_302_));
 sg13g2_a21oi_1 _478_ (.A1(_129_),
    .A2(_132_),
    .Y(_133_),
    .B1(_037_));
 sg13g2_o21ai_1 _479_ (.B1(_100_),
    .Y(_134_),
    .A1(_041_),
    .A2(_056_));
 sg13g2_a21oi_1 _480_ (.A1(_284_),
    .A2(_070_),
    .Y(_135_),
    .B1(_130_));
 sg13g2_xnor2_1 _481_ (.Y(_136_),
    .A(_284_),
    .B(_289_));
 sg13g2_a21oi_1 _482_ (.A1(_093_),
    .A2(_136_),
    .Y(_137_),
    .B1(_135_));
 sg13g2_a21oi_1 _483_ (.A1(_134_),
    .A2(_137_),
    .Y(_138_),
    .B1(_054_));
 sg13g2_a21oi_1 _484_ (.A1(_296_),
    .A2(_304_),
    .Y(_139_),
    .B1(_067_));
 sg13g2_a221oi_1 _485_ (.B2(_110_),
    .C1(_124_),
    .B1(_139_),
    .A1(_126_),
    .Y(_140_),
    .A2(_128_));
 sg13g2_nor2_1 _486_ (.A(net135),
    .B(_140_),
    .Y(_141_));
 sg13g2_nor4_1 _487_ (.A(net134),
    .B(_133_),
    .C(_138_),
    .D(_141_),
    .Y(_142_));
 sg13g2_a21oi_2 _488_ (.B1(_142_),
    .Y(uo_out[1]),
    .A2(_122_),
    .A1(_119_));
 sg13g2_nand2_1 _489_ (.Y(_143_),
    .A(_062_),
    .B(_112_));
 sg13g2_nand3_1 _490_ (.B(_033_),
    .C(_093_),
    .A(_318_),
    .Y(_144_));
 sg13g2_a22oi_1 _491_ (.Y(_145_),
    .B1(_143_),
    .B2(net147),
    .A2(_100_),
    .A1(_301_));
 sg13g2_nand3_1 _492_ (.B(_144_),
    .C(_145_),
    .A(net140),
    .Y(_146_));
 sg13g2_nor2b_1 _493_ (.A(net141),
    .B_N(_095_),
    .Y(_147_));
 sg13g2_nand2b_1 _494_ (.Y(_148_),
    .B(_095_),
    .A_N(net141));
 sg13g2_a21oi_1 _495_ (.A1(_146_),
    .A2(_148_),
    .Y(_149_),
    .B1(_302_));
 sg13g2_nor2_1 _496_ (.A(net140),
    .B(_303_),
    .Y(_150_));
 sg13g2_nor2b_1 _497_ (.A(_136_),
    .B_N(_150_),
    .Y(_151_));
 sg13g2_nor3_1 _498_ (.A(net136),
    .B(_149_),
    .C(_151_),
    .Y(_152_));
 sg13g2_o21ai_1 _499_ (.B1(net133),
    .Y(_153_),
    .A1(_004_),
    .A2(_143_));
 sg13g2_a22oi_1 _500_ (.Y(_154_),
    .B1(_306_),
    .B2(_099_),
    .A2(_302_),
    .A1(net163));
 sg13g2_nand2_1 _501_ (.Y(_155_),
    .A(_153_),
    .B(_154_));
 sg13g2_o21ai_1 _502_ (.B1(net146),
    .Y(_156_),
    .A1(net155),
    .A2(net149));
 sg13g2_nand2b_1 _503_ (.Y(_157_),
    .B(_066_),
    .A_N(_156_));
 sg13g2_a21oi_2 _504_ (.B1(net155),
    .Y(_158_),
    .A2(net163),
    .A1(net160));
 sg13g2_a21oi_1 _505_ (.A1(_301_),
    .A2(_158_),
    .Y(_159_),
    .B1(_043_));
 sg13g2_o21ai_1 _506_ (.B1(_157_),
    .Y(_160_),
    .A1(net146),
    .A2(_159_));
 sg13g2_a221oi_1 _507_ (.B2(_053_),
    .C1(_152_),
    .B1(_160_),
    .A1(_036_),
    .Y(_161_),
    .A2(_155_));
 sg13g2_nor2_1 _508_ (.A(net133),
    .B(net149),
    .Y(_162_));
 sg13g2_a21oi_1 _509_ (.A1(net129),
    .A2(_100_),
    .Y(_163_),
    .B1(_302_));
 sg13g2_a22oi_1 _510_ (.Y(_164_),
    .B1(_163_),
    .B2(_147_),
    .A2(_150_),
    .A1(_107_));
 sg13g2_o21ai_1 _511_ (.B1(_164_),
    .Y(_165_),
    .A1(_146_),
    .A2(_162_));
 sg13g2_nand2b_1 _512_ (.Y(_166_),
    .B(_165_),
    .A_N(net136));
 sg13g2_nor2_1 _513_ (.A(net155),
    .B(_130_),
    .Y(_167_));
 sg13g2_nand3_1 _514_ (.B(_093_),
    .C(_112_),
    .A(_062_),
    .Y(_168_));
 sg13g2_a22oi_1 _515_ (.Y(_169_),
    .B1(_057_),
    .B2(_167_),
    .A2(_302_),
    .A1(_006_));
 sg13g2_a21oi_1 _516_ (.A1(_168_),
    .A2(_169_),
    .Y(_170_),
    .B1(_037_));
 sg13g2_a221oi_1 _517_ (.B2(_110_),
    .C1(_054_),
    .B1(_077_),
    .A1(net145),
    .Y(_171_),
    .A2(_066_));
 sg13g2_nor3_1 _518_ (.A(_280_),
    .B(_170_),
    .C(_171_),
    .Y(_172_));
 sg13g2_a22oi_1 _519_ (.Y(uo_out[2]),
    .B1(_166_),
    .B2(_172_),
    .A2(_161_),
    .A1(_280_));
 sg13g2_nor2b_2 _520_ (.A(_313_),
    .B_N(_038_),
    .Y(_173_));
 sg13g2_nand2_1 _521_ (.Y(_174_),
    .A(net150),
    .B(_173_));
 sg13g2_a221oi_1 _522_ (.B2(net151),
    .C1(_071_),
    .B1(_173_),
    .A1(_319_),
    .Y(_175_),
    .A2(_158_));
 sg13g2_nand3_1 _523_ (.B(_303_),
    .C(_130_),
    .A(net138),
    .Y(_176_));
 sg13g2_a21oi_1 _524_ (.A1(net151),
    .A2(net158),
    .Y(_177_),
    .B1(net143));
 sg13g2_nand3_1 _525_ (.B(_081_),
    .C(_112_),
    .A(_318_),
    .Y(_178_));
 sg13g2_a21oi_1 _526_ (.A1(_177_),
    .A2(_178_),
    .Y(_179_),
    .B1(_176_));
 sg13g2_and2_1 _527_ (.A(net157),
    .B(net130),
    .X(_180_));
 sg13g2_nand2_2 _528_ (.Y(_181_),
    .A(net157),
    .B(net130));
 sg13g2_a221oi_1 _529_ (.B2(_181_),
    .C1(_067_),
    .B1(_158_),
    .A1(_315_),
    .Y(_182_),
    .A2(_025_));
 sg13g2_nor3_1 _530_ (.A(_175_),
    .B(_179_),
    .C(_182_),
    .Y(_183_));
 sg13g2_a21oi_1 _531_ (.A1(net129),
    .A2(_050_),
    .Y(_184_),
    .B1(_078_));
 sg13g2_nor2_1 _532_ (.A(net142),
    .B(_184_),
    .Y(_185_));
 sg13g2_a21oi_1 _533_ (.A1(_297_),
    .A2(_319_),
    .Y(_186_),
    .B1(_303_));
 sg13g2_a21oi_1 _534_ (.A1(_046_),
    .A2(_173_),
    .Y(_187_),
    .B1(_307_));
 sg13g2_nand3_1 _535_ (.B(net158),
    .C(net162),
    .A(net153),
    .Y(_188_));
 sg13g2_a21oi_1 _536_ (.A1(_297_),
    .A2(_181_),
    .Y(_189_),
    .B1(_094_));
 sg13g2_or4_1 _537_ (.A(_185_),
    .B(_186_),
    .C(_187_),
    .D(_189_),
    .X(_190_));
 sg13g2_nor2b_1 _538_ (.A(_075_),
    .B_N(_297_),
    .Y(_191_));
 sg13g2_a21oi_1 _539_ (.A1(_285_),
    .A2(_315_),
    .Y(_192_),
    .B1(net152));
 sg13g2_or3_1 _540_ (.A(net132),
    .B(_191_),
    .C(_192_),
    .X(_193_));
 sg13g2_or3_1 _541_ (.A(net149),
    .B(_005_),
    .C(net130),
    .X(_194_));
 sg13g2_a21oi_1 _542_ (.A1(net132),
    .A2(_194_),
    .Y(_195_),
    .B1(_037_));
 sg13g2_o21ai_1 _543_ (.B1(net134),
    .Y(_196_),
    .A1(net135),
    .A2(_183_));
 sg13g2_a221oi_1 _544_ (.B2(_195_),
    .C1(_196_),
    .B1(_193_),
    .A1(_053_),
    .Y(_197_),
    .A2(_190_));
 sg13g2_nand3_1 _545_ (.B(_315_),
    .C(_025_),
    .A(net143),
    .Y(_198_));
 sg13g2_o21ai_1 _546_ (.B1(_198_),
    .Y(_199_),
    .A1(net151),
    .A2(_173_));
 sg13g2_nor3_1 _547_ (.A(net138),
    .B(_189_),
    .C(_199_),
    .Y(_200_));
 sg13g2_xnor2_1 _548_ (.Y(_201_),
    .A(net157),
    .B(net130));
 sg13g2_a221oi_1 _549_ (.B2(_201_),
    .C1(_176_),
    .B1(_100_),
    .A1(net157),
    .Y(_202_),
    .A2(_093_));
 sg13g2_nor3_1 _550_ (.A(net135),
    .B(_200_),
    .C(_202_),
    .Y(_203_));
 sg13g2_o21ai_1 _551_ (.B1(net132),
    .Y(_204_),
    .A1(net149),
    .A2(_112_));
 sg13g2_nand2_1 _552_ (.Y(_205_),
    .A(_193_),
    .B(_204_));
 sg13g2_a21oi_1 _553_ (.A1(net142),
    .A2(_045_),
    .Y(_206_),
    .B1(_174_));
 sg13g2_nand3_1 _554_ (.B(_319_),
    .C(_158_),
    .A(net143),
    .Y(_207_));
 sg13g2_nor3_1 _555_ (.A(_054_),
    .B(_185_),
    .C(_206_),
    .Y(_208_));
 sg13g2_a221oi_1 _556_ (.B2(_208_),
    .C1(_203_),
    .B1(_207_),
    .A1(_036_),
    .Y(_209_),
    .A2(_205_));
 sg13g2_a21oi_2 _557_ (.B1(_197_),
    .Y(uo_out[3]),
    .A2(_209_),
    .A1(_280_));
 sg13g2_a22oi_1 _558_ (.Y(_210_),
    .B1(_100_),
    .B2(_114_),
    .A2(_093_),
    .A1(net157));
 sg13g2_nor2b_1 _559_ (.A(_210_),
    .B_N(net138),
    .Y(_211_));
 sg13g2_nor2_1 _560_ (.A(_289_),
    .B(_075_),
    .Y(_212_));
 sg13g2_nor3_1 _561_ (.A(_051_),
    .B(_078_),
    .C(_212_),
    .Y(_213_));
 sg13g2_nor2_1 _562_ (.A(_071_),
    .B(_213_),
    .Y(_214_));
 sg13g2_nor2b_1 _563_ (.A(net157),
    .B_N(net152),
    .Y(_215_));
 sg13g2_nor3_1 _564_ (.A(_067_),
    .B(_158_),
    .C(_215_),
    .Y(_216_));
 sg13g2_nor3_1 _565_ (.A(_211_),
    .B(_214_),
    .C(_216_),
    .Y(_217_));
 sg13g2_nand3_1 _566_ (.B(_286_),
    .C(_188_),
    .A(net135),
    .Y(_218_));
 sg13g2_o21ai_1 _567_ (.B1(_054_),
    .Y(_219_),
    .A1(_192_),
    .A2(_218_));
 sg13g2_a22oi_1 _568_ (.Y(_220_),
    .B1(_180_),
    .B2(net151),
    .A2(_085_),
    .A1(_315_));
 sg13g2_nor2_1 _569_ (.A(net132),
    .B(_213_),
    .Y(_221_));
 sg13g2_o21ai_1 _570_ (.B1(net138),
    .Y(_222_),
    .A1(net143),
    .A2(_220_));
 sg13g2_o21ai_1 _571_ (.B1(_219_),
    .Y(_223_),
    .A1(_221_),
    .A2(_222_));
 sg13g2_o21ai_1 _572_ (.B1(_223_),
    .Y(_224_),
    .A1(net135),
    .A2(_217_));
 sg13g2_nand2_1 _573_ (.Y(_225_),
    .A(net153),
    .B(_181_));
 sg13g2_a21oi_1 _574_ (.A1(net151),
    .A2(_180_),
    .Y(_226_),
    .B1(_079_));
 sg13g2_nand3b_1 _575_ (.B(_226_),
    .C(net143),
    .Y(_227_),
    .A_N(_047_));
 sg13g2_or3_1 _576_ (.A(net143),
    .B(_192_),
    .C(_212_),
    .X(_228_));
 sg13g2_nand3_1 _577_ (.B(_227_),
    .C(_228_),
    .A(net138),
    .Y(_229_));
 sg13g2_o21ai_1 _578_ (.B1(_177_),
    .Y(_230_),
    .A1(net151),
    .A2(_181_));
 sg13g2_nand2_1 _579_ (.Y(_231_),
    .A(net138),
    .B(_230_));
 sg13g2_nor2_1 _580_ (.A(_071_),
    .B(_226_),
    .Y(_232_));
 sg13g2_nor3_1 _581_ (.A(_025_),
    .B(_067_),
    .C(_079_),
    .Y(_233_));
 sg13g2_nor3_1 _582_ (.A(net137),
    .B(_232_),
    .C(_233_),
    .Y(_234_));
 sg13g2_a221oi_1 _583_ (.B2(_234_),
    .C1(net134),
    .B1(_231_),
    .A1(_219_),
    .Y(_235_),
    .A2(_229_));
 sg13g2_a21o_1 _584_ (.A2(_224_),
    .A1(net134),
    .B1(_235_),
    .X(uo_out[4]));
 sg13g2_nand2_1 _585_ (.Y(_236_),
    .A(_003_),
    .B(_225_));
 sg13g2_o21ai_1 _586_ (.B1(_236_),
    .Y(_237_),
    .A1(_003_),
    .A2(_158_));
 sg13g2_o21ai_1 _587_ (.B1(_287_),
    .Y(_238_),
    .A1(_049_),
    .A2(_225_));
 sg13g2_a21o_1 _588_ (.A2(_158_),
    .A1(_049_),
    .B1(_238_),
    .X(_239_));
 sg13g2_nor2_1 _589_ (.A(_037_),
    .B(_188_),
    .Y(_240_));
 sg13g2_nand3_1 _590_ (.B(_003_),
    .C(_029_),
    .A(net149),
    .Y(_241_));
 sg13g2_and3_1 _591_ (.X(_242_),
    .A(net145),
    .B(net149),
    .C(_297_));
 sg13g2_a21oi_1 _592_ (.A1(_028_),
    .A2(_114_),
    .Y(_243_),
    .B1(_242_));
 sg13g2_nand3_1 _593_ (.B(_037_),
    .C(_243_),
    .A(_030_),
    .Y(_244_));
 sg13g2_a22oi_1 _594_ (.Y(_245_),
    .B1(_240_),
    .B2(_286_),
    .A2(_116_),
    .A1(_029_));
 sg13g2_a21oi_1 _595_ (.A1(_244_),
    .A2(_245_),
    .Y(_246_),
    .B1(net134));
 sg13g2_o21ai_1 _596_ (.B1(net134),
    .Y(_247_),
    .A1(_181_),
    .A2(_241_));
 sg13g2_a221oi_1 _597_ (.B2(net145),
    .C1(_247_),
    .B1(_240_),
    .A1(_053_),
    .Y(_248_),
    .A2(_237_));
 sg13g2_a21oi_1 _598_ (.A1(_239_),
    .A2(_248_),
    .Y(uo_out[5]),
    .B1(_246_));
 sg13g2_o21ai_1 _599_ (.B1(_287_),
    .Y(_249_),
    .A1(_048_),
    .A2(_242_));
 sg13g2_o21ai_1 _600_ (.B1(_003_),
    .Y(_250_),
    .A1(net149),
    .A2(_115_));
 sg13g2_nand3b_1 _601_ (.B(_236_),
    .C(net136),
    .Y(_251_),
    .A_N(_002_));
 sg13g2_o21ai_1 _602_ (.B1(_287_),
    .Y(_252_),
    .A1(_003_),
    .A2(_158_));
 sg13g2_nand2_1 _603_ (.Y(_253_),
    .A(_251_),
    .B(_252_));
 sg13g2_a21oi_1 _604_ (.A1(_053_),
    .A2(_250_),
    .Y(_254_),
    .B1(_280_));
 sg13g2_a22oi_1 _605_ (.Y(uo_out[6]),
    .B1(_254_),
    .B2(_249_),
    .A2(_253_),
    .A1(_280_));
 sg13g2_nand2_1 _606_ (.Y(_255_),
    .A(_001_),
    .B(net129));
 sg13g2_nor4_1 _607_ (.A(net152),
    .B(_285_),
    .C(_071_),
    .D(_255_),
    .Y(_256_));
 sg13g2_or2_1 _608_ (.X(uo_out[7]),
    .B(_256_),
    .A(_000_));
 sg13g2_and2_1 _609_ (.A(net166),
    .B(net27),
    .X(_257_));
 sg13g2_xor2_1 _610_ (.B(net27),
    .A(net166),
    .X(_008_));
 sg13g2_and2_1 _611_ (.A(net163),
    .B(net32),
    .X(_258_));
 sg13g2_xor2_1 _612_ (.B(net32),
    .A(net163),
    .X(_259_));
 sg13g2_xor2_1 _613_ (.B(_259_),
    .A(_257_),
    .X(_009_));
 sg13g2_nand2_1 _614_ (.Y(_260_),
    .A(net160),
    .B(net34));
 sg13g2_xnor2_1 _615_ (.Y(_261_),
    .A(net161),
    .B(net34));
 sg13g2_a21oi_1 _616_ (.A1(_257_),
    .A2(_259_),
    .Y(_262_),
    .B1(_258_));
 sg13g2_xor2_1 _617_ (.B(_262_),
    .A(_261_),
    .X(_010_));
 sg13g2_and2_1 _618_ (.A(net156),
    .B(net31),
    .X(_263_));
 sg13g2_xor2_1 _619_ (.B(net31),
    .A(net156),
    .X(_264_));
 sg13g2_o21ai_1 _620_ (.B1(_260_),
    .Y(_265_),
    .A1(_261_),
    .A2(_262_));
 sg13g2_xor2_1 _621_ (.B(_265_),
    .A(_264_),
    .X(_011_));
 sg13g2_nand2_1 _622_ (.Y(_266_),
    .A(net146),
    .B(net36));
 sg13g2_xnor2_1 _623_ (.Y(_267_),
    .A(net146),
    .B(net36));
 sg13g2_a21o_1 _624_ (.A2(_265_),
    .A1(_264_),
    .B1(_263_),
    .X(_268_));
 sg13g2_nand2b_1 _625_ (.Y(_269_),
    .B(_268_),
    .A_N(_267_));
 sg13g2_xnor2_1 _626_ (.Y(_012_),
    .A(_267_),
    .B(_268_));
 sg13g2_nor2_1 _627_ (.A(net141),
    .B(net35),
    .Y(_270_));
 sg13g2_xor2_1 _628_ (.B(net35),
    .A(net140),
    .X(_271_));
 sg13g2_and2_1 _629_ (.A(_266_),
    .B(_269_),
    .X(_272_));
 sg13g2_xnor2_1 _630_ (.Y(_013_),
    .A(_271_),
    .B(_272_));
 sg13g2_and2_1 _631_ (.A(net136),
    .B(net33),
    .X(_273_));
 sg13g2_xor2_1 _632_ (.B(net33),
    .A(net136),
    .X(_274_));
 sg13g2_a22oi_1 _633_ (.Y(_275_),
    .B1(net35),
    .B2(net140),
    .A2(net39),
    .A1(net146));
 sg13g2_a21oi_1 _634_ (.A1(_269_),
    .A2(_275_),
    .Y(_276_),
    .B1(_270_));
 sg13g2_xor2_1 _635_ (.B(_276_),
    .A(_274_),
    .X(_014_));
 sg13g2_a21oi_1 _636_ (.A1(_274_),
    .A2(_276_),
    .Y(_277_),
    .B1(_273_));
 sg13g2_xor2_1 _637_ (.B(net30),
    .A(net37),
    .X(_278_));
 sg13g2_xnor2_1 _638_ (.Y(_015_),
    .A(_277_),
    .B(_278_));
 sg13g2_nor2_1 _639_ (.A(net29),
    .B(net10),
    .Y(_279_));
 sg13g2_a21oi_1 _640_ (.A1(net2),
    .A2(net167),
    .Y(_017_),
    .B1(_279_));
 sg13g2_mux2_1 _641_ (.A0(net32),
    .A1(net3),
    .S(net167),
    .X(_018_));
 sg13g2_mux2_1 _642_ (.A0(net34),
    .A1(net4),
    .S(net167),
    .X(_019_));
 sg13g2_mux2_1 _643_ (.A0(net31),
    .A1(net5),
    .S(net167),
    .X(_020_));
 sg13g2_mux2_1 _644_ (.A0(net36),
    .A1(net6),
    .S(net167),
    .X(_021_));
 sg13g2_mux2_1 _645_ (.A0(net35),
    .A1(net7),
    .S(net167),
    .X(_022_));
 sg13g2_mux2_1 _646_ (.A0(net33),
    .A1(net8),
    .S(net167),
    .X(_023_));
 sg13g2_mux2_1 _647_ (.A0(net30),
    .A1(net9),
    .S(net167),
    .X(_024_));
 sg13g2_dfrbp_1 _648_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net168),
    .D(_017_),
    .Q_N(\accum.PHASE_INC[0] ),
    .Q(_016_));
 sg13g2_dfrbp_1 _649_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net169),
    .D(_018_),
    .Q_N(_326_),
    .Q(\accum.PHASE_INC[1] ));
 sg13g2_dfrbp_1 _650_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net168),
    .D(_019_),
    .Q_N(_325_),
    .Q(\accum.PHASE_INC[2] ));
 sg13g2_dfrbp_1 _651_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net168),
    .D(_020_),
    .Q_N(_324_),
    .Q(\accum.PHASE_INC[3] ));
 sg13g2_dfrbp_1 _652_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net168),
    .D(_021_),
    .Q_N(_323_),
    .Q(\accum.PHASE_INC[4] ));
 sg13g2_dfrbp_1 _653_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net1),
    .D(_022_),
    .Q_N(_322_),
    .Q(\accum.PHASE_INC[5] ));
 sg13g2_dfrbp_1 _654_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net169),
    .D(_023_),
    .Q_N(_321_),
    .Q(\accum.PHASE_INC[6] ));
 sg13g2_dfrbp_1 _655_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net169),
    .D(_024_),
    .Q_N(_327_),
    .Q(\accum.PHASE_INC[7] ));
 sg13g2_dfrbp_1 _656_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net168),
    .D(net28),
    .Q_N(_007_),
    .Q(\accum.addr[0] ));
 sg13g2_dfrbp_1 _657_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net168),
    .D(_009_),
    .Q_N(_006_),
    .Q(\accum.addr[1] ));
 sg13g2_dfrbp_1 _658_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net168),
    .D(_010_),
    .Q_N(_005_),
    .Q(\accum.addr[2] ));
 sg13g2_dfrbp_1 _659_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net168),
    .D(_011_),
    .Q_N(_004_),
    .Q(\accum.addr[3] ));
 sg13g2_dfrbp_1 _660_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net169),
    .D(_012_),
    .Q_N(_003_),
    .Q(\accum.addr[4] ));
 sg13g2_dfrbp_1 _661_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net169),
    .D(_013_),
    .Q_N(_002_),
    .Q(\accum.addr[5] ));
 sg13g2_dfrbp_1 _662_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net169),
    .D(_014_),
    .Q_N(_001_),
    .Q(\accum.addr[6] ));
 sg13g2_dfrbp_1 _663_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net169),
    .D(_015_),
    .Q_N(_000_),
    .Q(\accum.addr[7] ));
 sg13g2_tielo tt_um_abhinav8prasad_dds_12 (.L_LO(net12));
 sg13g2_tielo tt_um_abhinav8prasad_dds_13 (.L_LO(net13));
 sg13g2_tielo tt_um_abhinav8prasad_dds_14 (.L_LO(net14));
 sg13g2_tielo tt_um_abhinav8prasad_dds_15 (.L_LO(net15));
 sg13g2_tielo tt_um_abhinav8prasad_dds_16 (.L_LO(net16));
 sg13g2_tielo tt_um_abhinav8prasad_dds_17 (.L_LO(net17));
 sg13g2_tielo tt_um_abhinav8prasad_dds_18 (.L_LO(net18));
 sg13g2_tielo tt_um_abhinav8prasad_dds_19 (.L_LO(net19));
 sg13g2_tielo tt_um_abhinav8prasad_dds_20 (.L_LO(net20));
 sg13g2_tielo tt_um_abhinav8prasad_dds_21 (.L_LO(net21));
 sg13g2_tielo tt_um_abhinav8prasad_dds_22 (.L_LO(net22));
 sg13g2_tielo tt_um_abhinav8prasad_dds_23 (.L_LO(net23));
 sg13g2_tielo tt_um_abhinav8prasad_dds_24 (.L_LO(net24));
 sg13g2_tielo tt_um_abhinav8prasad_dds_25 (.L_LO(net25));
 sg13g2_tielo tt_um_abhinav8prasad_dds_26 (.L_LO(net26));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 fanout129 (.A(_314_),
    .X(net129));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(_312_));
 sg13g2_buf_2 fanout131 (.A(_312_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(net133),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_281_),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(\accum.addr[7] ));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net137));
 sg13g2_buf_2 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(\accum.addr[6] ),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(\accum.addr[5] ),
    .X(net139));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(\accum.addr[5] ));
 sg13g2_buf_2 fanout141 (.A(\accum.addr[5] ),
    .X(net141));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net144));
 sg13g2_buf_2 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_1 fanout144 (.A(net145),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(net148),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(net148),
    .X(net146));
 sg13g2_buf_1 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(\accum.addr[4] ),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_004_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(net154),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(net154),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(\accum.addr[3] ),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(\accum.addr[3] ),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(\accum.addr[3] ),
    .X(net156));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(_005_));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(net161));
 sg13g2_buf_2 fanout159 (.A(net161),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(net161),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(net38),
    .X(net161));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(net163));
 sg13g2_buf_2 fanout163 (.A(\accum.addr[1] ),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(net165),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(\accum.addr[0] ),
    .X(net166));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(net10));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(net169));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(net1));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_tielo tt_um_abhinav8prasad_dds_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\accum.PHASE_INC[0] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold2 (.A(_008_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold3 (.A(_016_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold4 (.A(\accum.PHASE_INC[7] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold5 (.A(\accum.PHASE_INC[3] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold6 (.A(\accum.PHASE_INC[1] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold7 (.A(\accum.PHASE_INC[6] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold8 (.A(\accum.PHASE_INC[2] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold9 (.A(\accum.PHASE_INC[5] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold10 (.A(\accum.PHASE_INC[4] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold11 (.A(\accum.addr[7] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold12 (.A(\accum.addr[2] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold13 (.A(\accum.PHASE_INC[4] ),
    .X(net39));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_4 FILLER_23_182 ();
 sg13g2_fill_2 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_209 ();
 sg13g2_decap_4 FILLER_23_220 ();
 sg13g2_fill_2 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_230 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_fill_1 FILLER_23_239 ();
 sg13g2_decap_8 FILLER_23_248 ();
 sg13g2_decap_8 FILLER_23_255 ();
 sg13g2_decap_8 FILLER_23_262 ();
 sg13g2_decap_8 FILLER_23_269 ();
 sg13g2_decap_8 FILLER_23_276 ();
 sg13g2_decap_8 FILLER_23_283 ();
 sg13g2_decap_8 FILLER_23_290 ();
 sg13g2_decap_8 FILLER_23_297 ();
 sg13g2_decap_8 FILLER_23_304 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_decap_8 FILLER_23_318 ();
 sg13g2_decap_8 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_8 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_decap_8 FILLER_24_163 ();
 sg13g2_fill_2 FILLER_24_170 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_fill_2 FILLER_24_177 ();
 sg13g2_decap_8 FILLER_24_187 ();
 sg13g2_fill_2 FILLER_24_194 ();
 sg13g2_fill_1 FILLER_24_196 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_223 ();
 sg13g2_fill_2 FILLER_24_233 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_241 ();
 sg13g2_fill_2 FILLER_24_247 ();
 sg13g2_fill_2 FILLER_24_259 ();
 sg13g2_fill_2 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_293 ();
 sg13g2_decap_8 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_314 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_decap_8 FILLER_24_328 ();
 sg13g2_decap_8 FILLER_24_335 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_4 FILLER_25_140 ();
 sg13g2_fill_1 FILLER_25_144 ();
 sg13g2_fill_2 FILLER_25_159 ();
 sg13g2_fill_1 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_167 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_decap_8 FILLER_25_208 ();
 sg13g2_decap_4 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_228 ();
 sg13g2_decap_8 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_247 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_fill_2 FILLER_25_265 ();
 sg13g2_fill_1 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_284 ();
 sg13g2_decap_8 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_321 ();
 sg13g2_decap_4 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_4 FILLER_26_152 ();
 sg13g2_fill_2 FILLER_26_156 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_decap_4 FILLER_26_235 ();
 sg13g2_fill_2 FILLER_26_268 ();
 sg13g2_fill_1 FILLER_26_270 ();
 sg13g2_decap_4 FILLER_26_288 ();
 sg13g2_fill_1 FILLER_26_292 ();
 sg13g2_fill_2 FILLER_26_317 ();
 sg13g2_fill_1 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_132 ();
 sg13g2_decap_8 FILLER_27_139 ();
 sg13g2_fill_1 FILLER_27_146 ();
 sg13g2_fill_2 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_fill_1 FILLER_27_168 ();
 sg13g2_decap_4 FILLER_27_178 ();
 sg13g2_fill_2 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_decap_4 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_228 ();
 sg13g2_decap_8 FILLER_27_237 ();
 sg13g2_decap_4 FILLER_27_244 ();
 sg13g2_fill_2 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_decap_8 FILLER_27_262 ();
 sg13g2_decap_4 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_296 ();
 sg13g2_fill_1 FILLER_27_303 ();
 sg13g2_decap_4 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_314 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_decap_8 FILLER_27_330 ();
 sg13g2_decap_8 FILLER_27_337 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_fill_2 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_370 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_decap_8 FILLER_27_384 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_4 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_128 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_fill_2 FILLER_28_150 ();
 sg13g2_decap_8 FILLER_28_162 ();
 sg13g2_fill_2 FILLER_28_169 ();
 sg13g2_decap_4 FILLER_28_192 ();
 sg13g2_decap_8 FILLER_28_206 ();
 sg13g2_fill_2 FILLER_28_222 ();
 sg13g2_decap_8 FILLER_28_244 ();
 sg13g2_decap_8 FILLER_28_267 ();
 sg13g2_decap_4 FILLER_28_274 ();
 sg13g2_fill_2 FILLER_28_278 ();
 sg13g2_decap_4 FILLER_28_289 ();
 sg13g2_fill_2 FILLER_28_293 ();
 sg13g2_fill_2 FILLER_28_305 ();
 sg13g2_decap_8 FILLER_28_325 ();
 sg13g2_fill_1 FILLER_28_332 ();
 sg13g2_fill_2 FILLER_28_337 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_4 FILLER_29_168 ();
 sg13g2_fill_2 FILLER_29_179 ();
 sg13g2_fill_2 FILLER_29_201 ();
 sg13g2_fill_1 FILLER_29_203 ();
 sg13g2_fill_1 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_219 ();
 sg13g2_decap_8 FILLER_29_225 ();
 sg13g2_fill_2 FILLER_29_232 ();
 sg13g2_fill_2 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_250 ();
 sg13g2_decap_4 FILLER_29_269 ();
 sg13g2_fill_2 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_293 ();
 sg13g2_fill_1 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_decap_4 FILLER_29_323 ();
 sg13g2_decap_4 FILLER_29_348 ();
 sg13g2_decap_4 FILLER_29_360 ();
 sg13g2_fill_2 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_134 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_fill_2 FILLER_30_156 ();
 sg13g2_fill_1 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_167 ();
 sg13g2_decap_4 FILLER_30_179 ();
 sg13g2_fill_2 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_4 FILLER_30_196 ();
 sg13g2_fill_2 FILLER_30_200 ();
 sg13g2_fill_2 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_decap_8 FILLER_30_258 ();
 sg13g2_decap_8 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_decap_8 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_fill_1 FILLER_30_354 ();
 sg13g2_fill_2 FILLER_30_373 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_fill_2 FILLER_30_392 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_4 FILLER_31_105 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_decap_8 FILLER_31_128 ();
 sg13g2_decap_8 FILLER_31_135 ();
 sg13g2_decap_8 FILLER_31_142 ();
 sg13g2_fill_2 FILLER_31_170 ();
 sg13g2_fill_1 FILLER_31_172 ();
 sg13g2_decap_4 FILLER_31_178 ();
 sg13g2_decap_4 FILLER_31_186 ();
 sg13g2_decap_8 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_decap_8 FILLER_31_209 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_decap_8 FILLER_31_221 ();
 sg13g2_decap_4 FILLER_31_228 ();
 sg13g2_fill_2 FILLER_31_232 ();
 sg13g2_decap_8 FILLER_31_265 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_decap_8 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_304 ();
 sg13g2_fill_2 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_fill_2 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_124 ();
 sg13g2_fill_2 FILLER_32_131 ();
 sg13g2_decap_4 FILLER_32_153 ();
 sg13g2_fill_1 FILLER_32_157 ();
 sg13g2_fill_2 FILLER_32_163 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_decap_4 FILLER_32_175 ();
 sg13g2_decap_4 FILLER_32_197 ();
 sg13g2_fill_2 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_207 ();
 sg13g2_fill_2 FILLER_32_216 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_decap_4 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_244 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_fill_1 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_265 ();
 sg13g2_fill_2 FILLER_32_305 ();
 sg13g2_decap_4 FILLER_32_319 ();
 sg13g2_decap_8 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_346 ();
 sg13g2_decap_8 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_360 ();
 sg13g2_decap_4 FILLER_32_367 ();
 sg13g2_fill_2 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_fill_2 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_4 FILLER_33_133 ();
 sg13g2_fill_2 FILLER_33_137 ();
 sg13g2_decap_8 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_157 ();
 sg13g2_fill_1 FILLER_33_159 ();
 sg13g2_decap_4 FILLER_33_176 ();
 sg13g2_fill_2 FILLER_33_180 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_decap_4 FILLER_33_213 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_233 ();
 sg13g2_fill_2 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_271 ();
 sg13g2_fill_1 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_283 ();
 sg13g2_decap_4 FILLER_33_290 ();
 sg13g2_fill_2 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_318 ();
 sg13g2_fill_2 FILLER_33_325 ();
 sg13g2_decap_8 FILLER_33_339 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_fill_2 FILLER_33_364 ();
 sg13g2_fill_1 FILLER_33_366 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_112 ();
 sg13g2_decap_4 FILLER_34_133 ();
 sg13g2_fill_2 FILLER_34_137 ();
 sg13g2_decap_8 FILLER_34_153 ();
 sg13g2_fill_1 FILLER_34_160 ();
 sg13g2_decap_4 FILLER_34_169 ();
 sg13g2_fill_2 FILLER_34_173 ();
 sg13g2_decap_4 FILLER_34_184 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_decap_4 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_198 ();
 sg13g2_fill_1 FILLER_34_219 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_246 ();
 sg13g2_decap_8 FILLER_34_257 ();
 sg13g2_decap_4 FILLER_34_264 ();
 sg13g2_fill_2 FILLER_34_274 ();
 sg13g2_decap_8 FILLER_34_299 ();
 sg13g2_decap_4 FILLER_34_306 ();
 sg13g2_fill_2 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_320 ();
 sg13g2_decap_8 FILLER_34_327 ();
 sg13g2_decap_8 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_fill_2 FILLER_34_347 ();
 sg13g2_fill_1 FILLER_34_349 ();
 sg13g2_decap_8 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_383 ();
 sg13g2_fill_2 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_114 ();
 sg13g2_fill_2 FILLER_35_121 ();
 sg13g2_fill_2 FILLER_35_143 ();
 sg13g2_fill_1 FILLER_35_145 ();
 sg13g2_fill_2 FILLER_35_158 ();
 sg13g2_fill_2 FILLER_35_172 ();
 sg13g2_fill_1 FILLER_35_179 ();
 sg13g2_decap_8 FILLER_35_194 ();
 sg13g2_fill_2 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_decap_4 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_243 ();
 sg13g2_fill_1 FILLER_35_249 ();
 sg13g2_fill_2 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_264 ();
 sg13g2_decap_8 FILLER_35_281 ();
 sg13g2_decap_8 FILLER_35_288 ();
 sg13g2_fill_2 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_342 ();
 sg13g2_decap_4 FILLER_35_360 ();
 sg13g2_fill_2 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_402 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_4 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_127 ();
 sg13g2_decap_4 FILLER_36_134 ();
 sg13g2_fill_2 FILLER_36_138 ();
 sg13g2_decap_8 FILLER_36_149 ();
 sg13g2_fill_2 FILLER_36_156 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_179 ();
 sg13g2_decap_4 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_190 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_4 FILLER_36_231 ();
 sg13g2_fill_2 FILLER_36_235 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_decap_4 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_decap_8 FILLER_36_271 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_fill_2 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_fill_1 FILLER_36_333 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_fill_2 FILLER_37_189 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_decap_8 FILLER_37_197 ();
 sg13g2_decap_8 FILLER_37_235 ();
 sg13g2_fill_2 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_fill_1 FILLER_37_284 ();
 sg13g2_decap_4 FILLER_37_301 ();
 sg13g2_fill_2 FILLER_37_313 ();
 sg13g2_fill_1 FILLER_37_334 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_fill_2 FILLER_38_215 ();
 sg13g2_fill_1 FILLER_38_217 ();
 sg13g2_decap_4 FILLER_38_244 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_4 FILLER_38_271 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_fill_1 FILLER_38_308 ();
 sg13g2_fill_1 FILLER_38_339 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net11;
 assign uio_oe[1] = net12;
 assign uio_oe[2] = net13;
 assign uio_oe[3] = net14;
 assign uio_oe[4] = net15;
 assign uio_oe[5] = net16;
 assign uio_oe[6] = net17;
 assign uio_oe[7] = net18;
 assign uio_out[0] = net19;
 assign uio_out[1] = net20;
 assign uio_out[2] = net21;
 assign uio_out[3] = net22;
 assign uio_out[4] = net23;
 assign uio_out[5] = net24;
 assign uio_out[6] = net25;
 assign uio_out[7] = net26;
endmodule
