module tt_um_rodald_cpr (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire net207;
 wire net208;
 wire clk_regs;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire \crp.controller.aluDec.aluRtypeDec.func[0] ;
 wire \crp.controller.aluDec.aluRtypeDec.func[1] ;
 wire \crp.controller.aluDec.aluRtypeDec.func[2] ;
 wire \crp.controller.aluDec.aluRtypeDec.func[3] ;
 wire \crp.controller.aluDec.aluRtypeDec.state[0] ;
 wire \crp.controller.aluDec.aluRtypeDec.state[1] ;
 wire \crp.controller.aluDec.aluRtypeDec.state[2] ;
 wire \crp.controller.aluDec.opcode[0] ;
 wire \crp.controller.aluDec.opcode[1] ;
 wire \crp.controller.aluDec.opcode[2] ;
 wire \crp.controller.aluDec.opcode[3] ;
 wire \crp.controller.flags[0] ;
 wire \crp.controller.flags[1] ;
 wire \crp.controller.flags[2] ;
 wire \crp.controller.flags[3] ;
 wire \crp.controller.mainDecoder.memWriteReq ;
 wire \crp.datapath.aluSrc1SelMux.d0[0] ;
 wire \crp.datapath.aluSrc1SelMux.d0[10] ;
 wire \crp.datapath.aluSrc1SelMux.d0[11] ;
 wire \crp.datapath.aluSrc1SelMux.d0[12] ;
 wire \crp.datapath.aluSrc1SelMux.d0[13] ;
 wire \crp.datapath.aluSrc1SelMux.d0[14] ;
 wire \crp.datapath.aluSrc1SelMux.d0[1] ;
 wire \crp.datapath.aluSrc1SelMux.d0[2] ;
 wire \crp.datapath.aluSrc1SelMux.d0[3] ;
 wire \crp.datapath.aluSrc1SelMux.d0[4] ;
 wire \crp.datapath.aluSrc1SelMux.d0[5] ;
 wire \crp.datapath.aluSrc1SelMux.d0[6] ;
 wire \crp.datapath.aluSrc1SelMux.d0[7] ;
 wire \crp.datapath.aluSrc1SelMux.d0[8] ;
 wire \crp.datapath.aluSrc1SelMux.d0[9] ;
 wire \crp.datapath.aluSrc1SelMux.d1[0] ;
 wire \crp.datapath.aluSrc1SelMux.d1[10] ;
 wire \crp.datapath.aluSrc1SelMux.d1[11] ;
 wire \crp.datapath.aluSrc1SelMux.d1[12] ;
 wire \crp.datapath.aluSrc1SelMux.d1[13] ;
 wire \crp.datapath.aluSrc1SelMux.d1[14] ;
 wire \crp.datapath.aluSrc1SelMux.d1[1] ;
 wire \crp.datapath.aluSrc1SelMux.d1[2] ;
 wire \crp.datapath.aluSrc1SelMux.d1[3] ;
 wire \crp.datapath.aluSrc1SelMux.d1[4] ;
 wire \crp.datapath.aluSrc1SelMux.d1[5] ;
 wire \crp.datapath.aluSrc1SelMux.d1[6] ;
 wire \crp.datapath.aluSrc1SelMux.d1[7] ;
 wire \crp.datapath.aluSrc1SelMux.d1[8] ;
 wire \crp.datapath.aluSrc1SelMux.d1[9] ;
 wire \crp.datapath.aluSrc2SelMux.d2[4] ;
 wire \crp.datapath.aluSrc2SelMux.d2[5] ;
 wire \crp.datapath.aluSrc2SelMux.d2[6] ;
 wire \crp.datapath.aluSrc2SelMux.d2[7] ;
 wire \crp.datapath.aluSrc2SelMux.d3[10] ;
 wire \crp.datapath.aluSrc2SelMux.d3[11] ;
 wire \crp.datapath.aluSrc2SelMux.d3[12] ;
 wire \crp.datapath.aluSrc2SelMux.d3[9] ;
 wire \crp.datapath.memReadData[0] ;
 wire \crp.datapath.memReadData[1] ;
 wire \crp.datapath.memReadData[2] ;
 wire \crp.datapath.memReadData[3] ;
 wire \crp.datapath.memReadData[4] ;
 wire \crp.datapath.memReadData[5] ;
 wire \crp.datapath.memReadData[6] ;
 wire \crp.datapath.memReadData[7] ;
 wire \crp.datapath.registerFile.regs[0][0] ;
 wire \crp.datapath.registerFile.regs[0][1] ;
 wire \crp.datapath.registerFile.regs[0][2] ;
 wire \crp.datapath.registerFile.regs[0][3] ;
 wire \crp.datapath.registerFile.regs[0][4] ;
 wire \crp.datapath.registerFile.regs[0][5] ;
 wire \crp.datapath.registerFile.regs[0][6] ;
 wire \crp.datapath.registerFile.regs[0][7] ;
 wire \crp.datapath.registerFile.regs[10][0] ;
 wire \crp.datapath.registerFile.regs[10][1] ;
 wire \crp.datapath.registerFile.regs[10][2] ;
 wire \crp.datapath.registerFile.regs[10][3] ;
 wire \crp.datapath.registerFile.regs[10][4] ;
 wire \crp.datapath.registerFile.regs[10][5] ;
 wire \crp.datapath.registerFile.regs[10][6] ;
 wire \crp.datapath.registerFile.regs[10][7] ;
 wire \crp.datapath.registerFile.regs[11][0] ;
 wire \crp.datapath.registerFile.regs[11][1] ;
 wire \crp.datapath.registerFile.regs[11][2] ;
 wire \crp.datapath.registerFile.regs[11][3] ;
 wire \crp.datapath.registerFile.regs[11][4] ;
 wire \crp.datapath.registerFile.regs[11][5] ;
 wire \crp.datapath.registerFile.regs[11][6] ;
 wire \crp.datapath.registerFile.regs[11][7] ;
 wire \crp.datapath.registerFile.regs[12][0] ;
 wire \crp.datapath.registerFile.regs[12][1] ;
 wire \crp.datapath.registerFile.regs[12][2] ;
 wire \crp.datapath.registerFile.regs[12][3] ;
 wire \crp.datapath.registerFile.regs[12][4] ;
 wire \crp.datapath.registerFile.regs[12][5] ;
 wire \crp.datapath.registerFile.regs[12][6] ;
 wire \crp.datapath.registerFile.regs[12][7] ;
 wire \crp.datapath.registerFile.regs[13][0] ;
 wire \crp.datapath.registerFile.regs[13][1] ;
 wire \crp.datapath.registerFile.regs[13][2] ;
 wire \crp.datapath.registerFile.regs[13][3] ;
 wire \crp.datapath.registerFile.regs[13][4] ;
 wire \crp.datapath.registerFile.regs[13][5] ;
 wire \crp.datapath.registerFile.regs[13][6] ;
 wire \crp.datapath.registerFile.regs[13][7] ;
 wire \crp.datapath.registerFile.regs[14][0] ;
 wire \crp.datapath.registerFile.regs[14][1] ;
 wire \crp.datapath.registerFile.regs[14][2] ;
 wire \crp.datapath.registerFile.regs[14][3] ;
 wire \crp.datapath.registerFile.regs[14][4] ;
 wire \crp.datapath.registerFile.regs[14][5] ;
 wire \crp.datapath.registerFile.regs[14][6] ;
 wire \crp.datapath.registerFile.regs[14][7] ;
 wire \crp.datapath.registerFile.regs[15][0] ;
 wire \crp.datapath.registerFile.regs[15][1] ;
 wire \crp.datapath.registerFile.regs[15][2] ;
 wire \crp.datapath.registerFile.regs[15][3] ;
 wire \crp.datapath.registerFile.regs[15][4] ;
 wire \crp.datapath.registerFile.regs[15][5] ;
 wire \crp.datapath.registerFile.regs[15][6] ;
 wire \crp.datapath.registerFile.regs[15][7] ;
 wire \crp.datapath.registerFile.regs[1][0] ;
 wire \crp.datapath.registerFile.regs[1][1] ;
 wire \crp.datapath.registerFile.regs[1][2] ;
 wire \crp.datapath.registerFile.regs[1][3] ;
 wire \crp.datapath.registerFile.regs[1][4] ;
 wire \crp.datapath.registerFile.regs[1][5] ;
 wire \crp.datapath.registerFile.regs[1][6] ;
 wire \crp.datapath.registerFile.regs[1][7] ;
 wire \crp.datapath.registerFile.regs[2][0] ;
 wire \crp.datapath.registerFile.regs[2][1] ;
 wire \crp.datapath.registerFile.regs[2][2] ;
 wire \crp.datapath.registerFile.regs[2][3] ;
 wire \crp.datapath.registerFile.regs[2][4] ;
 wire \crp.datapath.registerFile.regs[2][5] ;
 wire \crp.datapath.registerFile.regs[2][6] ;
 wire \crp.datapath.registerFile.regs[2][7] ;
 wire \crp.datapath.registerFile.regs[3][0] ;
 wire \crp.datapath.registerFile.regs[3][1] ;
 wire \crp.datapath.registerFile.regs[3][2] ;
 wire \crp.datapath.registerFile.regs[3][3] ;
 wire \crp.datapath.registerFile.regs[3][4] ;
 wire \crp.datapath.registerFile.regs[3][5] ;
 wire \crp.datapath.registerFile.regs[3][6] ;
 wire \crp.datapath.registerFile.regs[3][7] ;
 wire \crp.datapath.registerFile.regs[4][0] ;
 wire \crp.datapath.registerFile.regs[4][1] ;
 wire \crp.datapath.registerFile.regs[4][2] ;
 wire \crp.datapath.registerFile.regs[4][3] ;
 wire \crp.datapath.registerFile.regs[4][4] ;
 wire \crp.datapath.registerFile.regs[4][5] ;
 wire \crp.datapath.registerFile.regs[4][6] ;
 wire \crp.datapath.registerFile.regs[4][7] ;
 wire \crp.datapath.registerFile.regs[5][0] ;
 wire \crp.datapath.registerFile.regs[5][1] ;
 wire \crp.datapath.registerFile.regs[5][2] ;
 wire \crp.datapath.registerFile.regs[5][3] ;
 wire \crp.datapath.registerFile.regs[5][4] ;
 wire \crp.datapath.registerFile.regs[5][5] ;
 wire \crp.datapath.registerFile.regs[5][6] ;
 wire \crp.datapath.registerFile.regs[5][7] ;
 wire \crp.datapath.registerFile.regs[6][0] ;
 wire \crp.datapath.registerFile.regs[6][1] ;
 wire \crp.datapath.registerFile.regs[6][2] ;
 wire \crp.datapath.registerFile.regs[6][3] ;
 wire \crp.datapath.registerFile.regs[6][4] ;
 wire \crp.datapath.registerFile.regs[6][5] ;
 wire \crp.datapath.registerFile.regs[6][6] ;
 wire \crp.datapath.registerFile.regs[6][7] ;
 wire \crp.datapath.registerFile.regs[7][0] ;
 wire \crp.datapath.registerFile.regs[7][1] ;
 wire \crp.datapath.registerFile.regs[7][2] ;
 wire \crp.datapath.registerFile.regs[7][3] ;
 wire \crp.datapath.registerFile.regs[7][4] ;
 wire \crp.datapath.registerFile.regs[7][5] ;
 wire \crp.datapath.registerFile.regs[7][6] ;
 wire \crp.datapath.registerFile.regs[7][7] ;
 wire \crp.datapath.registerFile.regs[8][0] ;
 wire \crp.datapath.registerFile.regs[8][1] ;
 wire \crp.datapath.registerFile.regs[8][2] ;
 wire \crp.datapath.registerFile.regs[8][3] ;
 wire \crp.datapath.registerFile.regs[8][4] ;
 wire \crp.datapath.registerFile.regs[8][5] ;
 wire \crp.datapath.registerFile.regs[8][6] ;
 wire \crp.datapath.registerFile.regs[8][7] ;
 wire \crp.datapath.registerFile.regs[9][0] ;
 wire \crp.datapath.registerFile.regs[9][1] ;
 wire \crp.datapath.registerFile.regs[9][2] ;
 wire \crp.datapath.registerFile.regs[9][3] ;
 wire \crp.datapath.registerFile.regs[9][4] ;
 wire \crp.datapath.registerFile.regs[9][5] ;
 wire \crp.datapath.registerFile.regs[9][6] ;
 wire \crp.datapath.registerFile.regs[9][7] ;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire delaynet_0_clk;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;

 sg13g2_inv_1 _1810_ (.Y(_1150_),
    .A(net376));
 sg13g2_inv_1 _1811_ (.Y(_1151_),
    .A(net377));
 sg13g2_inv_1 _1812_ (.Y(_1152_),
    .A(net209));
 sg13g2_inv_1 _1813_ (.Y(_1153_),
    .A(net364));
 sg13g2_inv_1 _1814_ (.Y(_1154_),
    .A(net332));
 sg13g2_inv_1 _1815_ (.Y(_1155_),
    .A(net350));
 sg13g2_inv_1 _1816_ (.Y(_1156_),
    .A(net321));
 sg13g2_inv_1 _1817_ (.Y(_1157_),
    .A(net723));
 sg13g2_inv_1 _1818_ (.Y(_1158_),
    .A(net724));
 sg13g2_inv_1 _1819_ (.Y(_1159_),
    .A(net3));
 sg13g2_inv_2 _1820_ (.Y(_1160_),
    .A(net726));
 sg13g2_inv_1 _1821_ (.Y(_1161_),
    .A(net2));
 sg13g2_inv_1 _1822_ (.Y(_1162_),
    .A(net389));
 sg13g2_inv_1 _1823_ (.Y(_1163_),
    .A(net299));
 sg13g2_inv_2 _1824_ (.Y(_1164_),
    .A(net385));
 sg13g2_inv_1 _1825_ (.Y(_1165_),
    .A(net384));
 sg13g2_inv_1 _1826_ (.Y(_1166_),
    .A(net378));
 sg13g2_inv_2 _1827_ (.Y(_1167_),
    .A(net373));
 sg13g2_inv_2 _1828_ (.Y(_1168_),
    .A(net374));
 sg13g2_inv_1 _1829_ (.Y(_1169_),
    .A(net381));
 sg13g2_inv_1 _1830_ (.Y(_1170_),
    .A(net382));
 sg13g2_inv_1 _1831_ (.Y(_1171_),
    .A(net358));
 sg13g2_inv_1 _1832_ (.Y(_1172_),
    .A(net307));
 sg13g2_inv_1 _1833_ (.Y(_1173_),
    .A(net322));
 sg13g2_inv_1 _1834_ (.Y(_1174_),
    .A(net345));
 sg13g2_inv_1 _1835_ (.Y(_1175_),
    .A(net365));
 sg13g2_inv_1 _1836_ (.Y(_1176_),
    .A(net360));
 sg13g2_inv_1 _1837_ (.Y(_1177_),
    .A(net362));
 sg13g2_inv_1 _1838_ (.Y(_1178_),
    .A(net352));
 sg13g2_inv_2 _1839_ (.Y(_1179_),
    .A(net367));
 sg13g2_inv_1 _1840_ (.Y(_1180_),
    .A(net222));
 sg13g2_inv_1 _1841_ (.Y(_1181_),
    .A(net210));
 sg13g2_inv_1 _1842_ (.Y(_1182_),
    .A(net212));
 sg13g2_inv_1 _1843_ (.Y(_1183_),
    .A(net217));
 sg13g2_inv_1 _1844_ (.Y(_1184_),
    .A(net320));
 sg13g2_inv_1 _1845_ (.Y(_1185_),
    .A(net303));
 sg13g2_inv_1 _1846_ (.Y(_1186_),
    .A(net337));
 sg13g2_inv_1 _1847_ (.Y(_1187_),
    .A(net230));
 sg13g2_inv_1 _1848_ (.Y(_1188_),
    .A(net211));
 sg13g2_inv_1 _1849_ (.Y(_1189_),
    .A(net742));
 sg13g2_inv_1 _1850_ (.Y(_1190_),
    .A(net733));
 sg13g2_inv_1 _1851_ (.Y(_1191_),
    .A(_0012_));
 sg13g2_inv_1 _1852_ (.Y(_1192_),
    .A(net223));
 sg13g2_inv_1 _1853_ (.Y(_1193_),
    .A(net224));
 sg13g2_inv_1 _1854_ (.Y(_1194_),
    .A(_0013_));
 sg13g2_inv_2 _1855_ (.Y(_1195_),
    .A(_0015_));
 sg13g2_inv_1 _1856_ (.Y(_1196_),
    .A(_0017_));
 sg13g2_inv_1 _1857_ (.Y(_1197_),
    .A(net214));
 sg13g2_inv_1 _1858_ (.Y(_1198_),
    .A(net215));
 sg13g2_inv_1 _1859_ (.Y(_1199_),
    .A(net226));
 sg13g2_inv_1 _1860_ (.Y(_1200_),
    .A(net221));
 sg13g2_inv_1 _1861_ (.Y(_1201_),
    .A(_0023_));
 sg13g2_inv_1 _1862_ (.Y(_1202_),
    .A(net216));
 sg13g2_inv_1 _1863_ (.Y(_1203_),
    .A(net218));
 sg13g2_inv_1 _1864_ (.Y(_1204_),
    .A(_0026_));
 sg13g2_inv_1 _1865_ (.Y(_1205_),
    .A(net220));
 sg13g2_inv_1 _1866_ (.Y(_1206_),
    .A(net228));
 sg13g2_inv_1 _1867_ (.Y(_1207_),
    .A(net713));
 sg13g2_inv_1 _1868_ (.Y(_1208_),
    .A(_0030_));
 sg13g2_inv_1 _1869_ (.Y(_1209_),
    .A(net227));
 sg13g2_inv_1 _1870_ (.Y(_1210_),
    .A(_0036_));
 sg13g2_inv_1 _1871_ (.Y(_1211_),
    .A(net219));
 sg13g2_inv_1 _1872_ (.Y(_1212_),
    .A(net213));
 sg13g2_inv_1 _1873_ (.Y(_1213_),
    .A(_0047_));
 sg13g2_inv_1 _1874_ (.Y(_1214_),
    .A(_0046_));
 sg13g2_inv_1 _1875_ (.Y(_1215_),
    .A(_0049_));
 sg13g2_inv_1 _1876_ (.Y(_1216_),
    .A(_0048_));
 sg13g2_inv_1 _1877_ (.Y(_1217_),
    .A(net235));
 sg13g2_inv_1 _1878_ (.Y(_1218_),
    .A(net305));
 sg13g2_inv_1 _1879_ (.Y(_1219_),
    .A(net260));
 sg13g2_inv_1 _1880_ (.Y(_1220_),
    .A(_0069_));
 sg13g2_inv_1 _1881_ (.Y(_1221_),
    .A(_0073_));
 sg13g2_inv_1 _1882_ (.Y(_1222_),
    .A(_0077_));
 sg13g2_inv_1 _1883_ (.Y(_1223_),
    .A(_0088_));
 sg13g2_inv_1 _1884_ (.Y(_1224_),
    .A(_0092_));
 sg13g2_inv_1 _1885_ (.Y(_1225_),
    .A(_0091_));
 sg13g2_inv_1 _1886_ (.Y(_1226_),
    .A(_0094_));
 sg13g2_inv_1 _1887_ (.Y(_1227_),
    .A(_0096_));
 sg13g2_inv_1 _1888_ (.Y(_1228_),
    .A(_0098_));
 sg13g2_inv_1 _1889_ (.Y(_1229_),
    .A(_0102_));
 sg13g2_inv_1 _1890_ (.Y(_1230_),
    .A(_0105_));
 sg13g2_inv_1 _1891_ (.Y(_1231_),
    .A(_0111_));
 sg13g2_inv_1 _1892_ (.Y(_1232_),
    .A(_0110_));
 sg13g2_inv_1 _1893_ (.Y(_1233_),
    .A(_0112_));
 sg13g2_inv_1 _1894_ (.Y(_1234_),
    .A(_0115_));
 sg13g2_inv_1 _1895_ (.Y(_1235_),
    .A(_0114_));
 sg13g2_inv_1 _1896_ (.Y(_1236_),
    .A(_0117_));
 sg13g2_inv_1 _1897_ (.Y(_1237_),
    .A(_0116_));
 sg13g2_inv_1 _1898_ (.Y(_1238_),
    .A(_0122_));
 sg13g2_inv_1 _1899_ (.Y(_1239_),
    .A(_0128_));
 sg13g2_inv_1 _1900_ (.Y(_1240_),
    .A(_0130_));
 sg13g2_inv_1 _1901_ (.Y(_1241_),
    .A(_0132_));
 sg13g2_inv_1 _1902_ (.Y(_1242_),
    .A(_0131_));
 sg13g2_inv_1 _1903_ (.Y(_1243_),
    .A(_0134_));
 sg13g2_inv_1 _1904_ (.Y(_1244_),
    .A(_0133_));
 sg13g2_inv_1 _1905_ (.Y(_1245_),
    .A(_0137_));
 sg13g2_inv_1 _1906_ (.Y(_1246_),
    .A(_0136_));
 sg13g2_inv_1 _1907_ (.Y(_1247_),
    .A(_0139_));
 sg13g2_inv_1 _1908_ (.Y(_1248_),
    .A(_0145_));
 sg13g2_inv_1 _1909_ (.Y(_1249_),
    .A(_0144_));
 sg13g2_inv_1 _1910_ (.Y(_1250_),
    .A(_0147_));
 sg13g2_inv_1 _1911_ (.Y(_1251_),
    .A(_0149_));
 sg13g2_inv_1 _1912_ (.Y(_1252_),
    .A(_0148_));
 sg13g2_inv_1 _1913_ (.Y(_1253_),
    .A(_0000_));
 sg13g2_inv_1 _1914_ (.Y(_1254_),
    .A(_0001_));
 sg13g2_inv_1 _1915_ (.Y(_1255_),
    .A(_0002_));
 sg13g2_inv_1 _1916_ (.Y(_1256_),
    .A(_0003_));
 sg13g2_inv_1 _1917_ (.Y(_1257_),
    .A(_0004_));
 sg13g2_inv_1 _1918_ (.Y(_1258_),
    .A(_0005_));
 sg13g2_inv_1 _1919_ (.Y(_1259_),
    .A(_0006_));
 sg13g2_inv_1 _3256__2 (.Y(net207),
    .A(clknet_1_0__leaf_clk));
 sg13g2_nor2_2 _1921_ (.A(\crp.controller.aluDec.aluRtypeDec.state[2] ),
    .B(\crp.controller.aluDec.aluRtypeDec.state[1] ),
    .Y(_1260_));
 sg13g2_nor2b_2 _1922_ (.A(net703),
    .B_N(net701),
    .Y(_1261_));
 sg13g2_nand2b_1 _1923_ (.Y(_1262_),
    .B(net390),
    .A_N(net703));
 sg13g2_and2_2 _1924_ (.A(_0007_),
    .B(_1261_),
    .X(_1263_));
 sg13g2_nand3b_1 _1925_ (.B(net701),
    .C(_0007_),
    .Y(_1264_),
    .A_N(net703));
 sg13g2_nand2_2 _1926_ (.Y(_1265_),
    .A(\crp.controller.aluDec.opcode[1] ),
    .B(\crp.controller.aluDec.opcode[0] ));
 sg13g2_nor2_2 _1927_ (.A(net728),
    .B(\crp.controller.aluDec.opcode[2] ),
    .Y(_1266_));
 sg13g2_nor4_2 _1928_ (.A(net728),
    .B(\crp.controller.aluDec.opcode[2] ),
    .C(net699),
    .Y(_1267_),
    .D(_1265_));
 sg13g2_nand2b_1 _1929_ (.Y(_1268_),
    .B(\crp.controller.aluDec.opcode[2] ),
    .A_N(\crp.controller.aluDec.opcode[1] ));
 sg13g2_nand2b_2 _1930_ (.Y(_1269_),
    .B(\crp.controller.aluDec.opcode[1] ),
    .A_N(\crp.controller.aluDec.opcode[0] ));
 sg13g2_nor2_1 _1931_ (.A(net728),
    .B(_1269_),
    .Y(_1270_));
 sg13g2_a21oi_1 _1932_ (.A1(_1268_),
    .A2(_1269_),
    .Y(_1271_),
    .B1(net728));
 sg13g2_a21oi_2 _1933_ (.B1(_1267_),
    .Y(_1272_),
    .A2(_1271_),
    .A1(_1263_));
 sg13g2_nand2b_2 _1934_ (.Y(_1273_),
    .B(\crp.controller.aluDec.opcode[0] ),
    .A_N(\crp.controller.aluDec.opcode[1] ));
 sg13g2_nor2_1 _1935_ (.A(net699),
    .B(_1273_),
    .Y(_1274_));
 sg13g2_and2_1 _1936_ (.A(_1266_),
    .B(_1274_),
    .X(_1275_));
 sg13g2_a221oi_1 _1937_ (.B2(_1266_),
    .C1(_1267_),
    .B1(_1274_),
    .A1(_1263_),
    .Y(_1276_),
    .A2(_1271_));
 sg13g2_nand2b_2 _1938_ (.Y(_1277_),
    .B(_1272_),
    .A_N(_1275_));
 sg13g2_nor2_2 _1939_ (.A(\crp.controller.aluDec.opcode[1] ),
    .B(\crp.controller.aluDec.opcode[0] ),
    .Y(_1278_));
 sg13g2_and2_1 _1940_ (.A(_1266_),
    .B(_1278_),
    .X(_1279_));
 sg13g2_nand2_2 _1941_ (.Y(_1280_),
    .A(_1266_),
    .B(_1278_));
 sg13g2_nand2b_2 _1942_ (.Y(_1281_),
    .B(net725),
    .A_N(net723));
 sg13g2_nand2b_1 _1943_ (.Y(_1282_),
    .B(net726),
    .A_N(\crp.controller.aluDec.aluRtypeDec.func[0] ));
 sg13g2_nor2_1 _1944_ (.A(net722),
    .B(\crp.controller.aluDec.aluRtypeDec.func[0] ),
    .Y(_1283_));
 sg13g2_nor2_1 _1945_ (.A(_1281_),
    .B(_1282_),
    .Y(_1284_));
 sg13g2_nor2_1 _1946_ (.A(_1160_),
    .B(_1162_),
    .Y(_1285_));
 sg13g2_nand2_2 _1947_ (.Y(_1286_),
    .A(net726),
    .B(net727));
 sg13g2_nor2_1 _1948_ (.A(net722),
    .B(net724),
    .Y(_1287_));
 sg13g2_or2_1 _1949_ (.X(_1288_),
    .B(net727),
    .A(net726));
 sg13g2_a22oi_1 _1950_ (.Y(_1289_),
    .B1(_1287_),
    .B2(_1288_),
    .A2(_1286_),
    .A1(net724));
 sg13g2_nor2_1 _1951_ (.A(_1284_),
    .B(_1289_),
    .Y(_1290_));
 sg13g2_or3_1 _1952_ (.A(_1263_),
    .B(_1284_),
    .C(_1289_),
    .X(_1291_));
 sg13g2_and2_1 _1953_ (.A(net694),
    .B(_1291_),
    .X(_1292_));
 sg13g2_nand3_1 _1954_ (.B(net703),
    .C(_0007_),
    .A(net701),
    .Y(_1293_));
 sg13g2_nor2_1 _1955_ (.A(net700),
    .B(_1293_),
    .Y(_1294_));
 sg13g2_nor2b_2 _1956_ (.A(net724),
    .B_N(net722),
    .Y(_1295_));
 sg13g2_nand2b_1 _1957_ (.Y(_1296_),
    .B(net722),
    .A_N(net724));
 sg13g2_nor4_2 _1958_ (.A(net700),
    .B(_1286_),
    .C(_1293_),
    .Y(_1297_),
    .D(_1296_));
 sg13g2_nand2_1 _1959_ (.Y(_1298_),
    .A(net722),
    .B(net724));
 sg13g2_or3_1 _1960_ (.A(net698),
    .B(_1286_),
    .C(_1298_),
    .X(_1299_));
 sg13g2_o21ai_1 _1961_ (.B1(_1299_),
    .Y(_1300_),
    .A1(_1284_),
    .A2(_1289_));
 sg13g2_nor2_1 _1962_ (.A(_1297_),
    .B(_1300_),
    .Y(_1301_));
 sg13g2_nor2b_1 _1963_ (.A(_1301_),
    .B_N(_1292_),
    .Y(_1302_));
 sg13g2_nor2_1 _1964_ (.A(_1277_),
    .B(_1302_),
    .Y(_1303_));
 sg13g2_nor2_2 _1965_ (.A(_1164_),
    .B(net699),
    .Y(_1304_));
 sg13g2_nor4_1 _1966_ (.A(net728),
    .B(_1164_),
    .C(net698),
    .D(_1265_),
    .Y(_1305_));
 sg13g2_nand2b_2 _1967_ (.Y(_1306_),
    .B(net728),
    .A_N(\crp.controller.aluDec.opcode[2] ));
 sg13g2_or2_1 _1968_ (.X(_1307_),
    .B(_1306_),
    .A(_1269_));
 sg13g2_nor2b_2 _1969_ (.A(net390),
    .B_N(net703),
    .Y(_1308_));
 sg13g2_inv_1 _1970_ (.Y(_1309_),
    .A(_1308_));
 sg13g2_nand2_1 _1971_ (.Y(_1310_),
    .A(\crp.controller.aluDec.aluRtypeDec.state[2] ),
    .B(_1308_));
 sg13g2_nor2_1 _1972_ (.A(_1265_),
    .B(_1306_),
    .Y(_1311_));
 sg13g2_nor2_1 _1973_ (.A(_1163_),
    .B(_1164_),
    .Y(_1312_));
 sg13g2_nor2_1 _1974_ (.A(_1311_),
    .B(_1312_),
    .Y(_1313_));
 sg13g2_o21ai_1 _1975_ (.B1(_1313_),
    .Y(_1314_),
    .A1(_1307_),
    .A2(_1310_));
 sg13g2_or2_1 _1976_ (.X(_1315_),
    .B(_1306_),
    .A(_1273_));
 sg13g2_nor3_1 _1977_ (.A(_0007_),
    .B(_1262_),
    .C(_1315_),
    .Y(_1316_));
 sg13g2_nor4_1 _1978_ (.A(\crp.controller.aluDec.opcode[1] ),
    .B(\crp.controller.aluDec.opcode[0] ),
    .C(net698),
    .D(_1306_),
    .Y(_1317_));
 sg13g2_inv_1 _1979_ (.Y(_1318_),
    .A(_1317_));
 sg13g2_nor4_1 _1980_ (.A(net693),
    .B(_1314_),
    .C(_1316_),
    .D(_1317_),
    .Y(_1319_));
 sg13g2_nor4_2 _1981_ (.A(net722),
    .B(net724),
    .C(net698),
    .Y(_1320_),
    .D(_1288_));
 sg13g2_nand2b_2 _1982_ (.Y(_1321_),
    .B(net700),
    .A_N(net701));
 sg13g2_nand2_2 _1983_ (.Y(_1322_),
    .A(net727),
    .B(_1295_));
 sg13g2_nor4_1 _1984_ (.A(\crp.controller.aluDec.aluRtypeDec.func[1] ),
    .B(net702),
    .C(_1321_),
    .D(_1322_),
    .Y(_1323_));
 sg13g2_and2_1 _1985_ (.A(_1284_),
    .B(_1294_),
    .X(_1324_));
 sg13g2_or3_1 _1986_ (.A(_1320_),
    .B(_1323_),
    .C(_1324_),
    .X(_1325_));
 sg13g2_nand2_1 _1987_ (.Y(_1326_),
    .A(_1162_),
    .B(_1295_));
 sg13g2_or2_1 _1988_ (.X(_1327_),
    .B(_1286_),
    .A(_1281_));
 sg13g2_nand2_1 _1989_ (.Y(_1328_),
    .A(_1326_),
    .B(_1327_));
 sg13g2_nor3_1 _1990_ (.A(net727),
    .B(_1293_),
    .C(_1296_),
    .Y(_1329_));
 sg13g2_nor2b_2 _1991_ (.A(net700),
    .B_N(_1329_),
    .Y(_1330_));
 sg13g2_or4_1 _1992_ (.A(net700),
    .B(_1281_),
    .C(_1293_),
    .D(_1286_),
    .X(_1331_));
 sg13g2_a21oi_1 _1993_ (.A1(_1294_),
    .A2(_1328_),
    .Y(_1332_),
    .B1(_1325_));
 sg13g2_nand2b_1 _1994_ (.Y(_1333_),
    .B(_1292_),
    .A_N(_1332_));
 sg13g2_and3_1 _1995_ (.X(_1334_),
    .A(_1303_),
    .B(_1319_),
    .C(_1333_));
 sg13g2_o21ai_1 _1996_ (.B1(net744),
    .Y(_1335_),
    .A1(_1260_),
    .A2(_1334_));
 sg13g2_a21o_1 _1997_ (.A2(net701),
    .A1(net702),
    .B1(net386),
    .X(_1336_));
 sg13g2_a21oi_1 _1998_ (.A1(_1293_),
    .A2(net387),
    .Y(_0284_),
    .B1(_1335_));
 sg13g2_a21oi_1 _1999_ (.A1(net391),
    .A2(_1309_),
    .Y(_0283_),
    .B1(_1335_));
 sg13g2_nor2_1 _2000_ (.A(_1152_),
    .B(_1335_),
    .Y(_0282_));
 sg13g2_nand2b_2 _2001_ (.Y(_1337_),
    .B(net701),
    .A_N(net700));
 sg13g2_or2_1 _2002_ (.X(_1338_),
    .B(_1337_),
    .A(net702));
 sg13g2_nor2_1 _2003_ (.A(_1307_),
    .B(_1338_),
    .Y(_1339_));
 sg13g2_o21ai_1 _2004_ (.B1(_1293_),
    .Y(_1340_),
    .A1(net702),
    .A2(_1321_));
 sg13g2_nor2b_1 _2005_ (.A(_1315_),
    .B_N(_1340_),
    .Y(_1341_));
 sg13g2_xnor2_1 _2006_ (.Y(_1342_),
    .A(net700),
    .B(\crp.controller.aluDec.aluRtypeDec.state[1] ));
 sg13g2_nor3_2 _2007_ (.A(_1269_),
    .B(_1306_),
    .C(_1342_),
    .Y(_1343_));
 sg13g2_and2_2 _2008_ (.A(net702),
    .B(_1343_),
    .X(_1344_));
 sg13g2_nor3_2 _2009_ (.A(net694),
    .B(_1341_),
    .C(_1344_),
    .Y(_1345_));
 sg13g2_nor3_2 _2010_ (.A(net726),
    .B(_1293_),
    .C(_1322_),
    .Y(_1346_));
 sg13g2_nor2_2 _2011_ (.A(_1297_),
    .B(_1346_),
    .Y(_1347_));
 sg13g2_or3_1 _2012_ (.A(_1281_),
    .B(_1286_),
    .C(_1337_),
    .X(_1348_));
 sg13g2_or3_2 _2013_ (.A(net698),
    .B(_1281_),
    .C(_1282_),
    .X(_1349_));
 sg13g2_nand2_1 _2014_ (.Y(_1350_),
    .A(_1348_),
    .B(_1349_));
 sg13g2_nor2_1 _2015_ (.A(_1326_),
    .B(_1337_),
    .Y(_1351_));
 sg13g2_nor3_2 _2016_ (.A(_1280_),
    .B(_1350_),
    .C(_1351_),
    .Y(_1352_));
 sg13g2_a21oi_1 _2017_ (.A1(_1347_),
    .A2(_1352_),
    .Y(_1353_),
    .B1(_1345_));
 sg13g2_a21o_1 _2018_ (.A2(_1352_),
    .A1(_1347_),
    .B1(_1345_),
    .X(_1354_));
 sg13g2_nor4_2 _2019_ (.A(_1280_),
    .B(_1297_),
    .C(_1330_),
    .Y(_1355_),
    .D(_1346_));
 sg13g2_nor2_1 _2020_ (.A(_1345_),
    .B(net665),
    .Y(_1356_));
 sg13g2_or2_2 _2021_ (.X(_1357_),
    .B(net665),
    .A(_1345_));
 sg13g2_o21ai_1 _2022_ (.B1(net695),
    .Y(_1358_),
    .A1(net699),
    .A2(_1322_));
 sg13g2_nor2_2 _2023_ (.A(_1330_),
    .B(_1358_),
    .Y(_1359_));
 sg13g2_or2_1 _2024_ (.X(_1360_),
    .B(_1358_),
    .A(_1330_));
 sg13g2_nand2_1 _2025_ (.Y(_1361_),
    .A(\crp.controller.flags[0] ),
    .B(_1311_));
 sg13g2_mux2_1 _2026_ (.A0(\crp.controller.aluDec.opcode[0] ),
    .A1(\crp.controller.aluDec.opcode[1] ),
    .S(\crp.controller.flags[2] ),
    .X(_1362_));
 sg13g2_a21oi_1 _2027_ (.A1(\crp.controller.flags[0] ),
    .A2(_1278_),
    .Y(_1363_),
    .B1(_1362_));
 sg13g2_nor2_1 _2028_ (.A(\crp.controller.flags[3] ),
    .B(\crp.controller.flags[1] ),
    .Y(_1364_));
 sg13g2_and2_1 _2029_ (.A(\crp.controller.flags[3] ),
    .B(\crp.controller.flags[1] ),
    .X(_1365_));
 sg13g2_nor3_1 _2030_ (.A(_1265_),
    .B(_1364_),
    .C(_1365_),
    .Y(_1366_));
 sg13g2_o21ai_1 _2031_ (.B1(_1312_),
    .Y(_1367_),
    .A1(_1363_),
    .A2(_1366_));
 sg13g2_a21o_1 _2032_ (.A2(_1367_),
    .A1(_1361_),
    .B1(_1338_),
    .X(_1368_));
 sg13g2_o21ai_1 _2033_ (.B1(net700),
    .Y(_1369_),
    .A1(_1261_),
    .A2(_1308_));
 sg13g2_nand2b_1 _2034_ (.Y(_1370_),
    .B(_1369_),
    .A_N(_1340_));
 sg13g2_o21ai_1 _2035_ (.B1(_1280_),
    .Y(_1371_),
    .A1(_1315_),
    .A2(_1337_));
 sg13g2_a21oi_1 _2036_ (.A1(_1343_),
    .A2(_1370_),
    .Y(_1372_),
    .B1(_1371_));
 sg13g2_nand3_1 _2037_ (.B(_1368_),
    .C(_1372_),
    .A(_1318_),
    .Y(_1373_));
 sg13g2_a21o_1 _2038_ (.A2(_1373_),
    .A1(_1360_),
    .B1(_1260_),
    .X(_1374_));
 sg13g2_inv_2 _2039_ (.Y(_1375_),
    .A(net613));
 sg13g2_nor3_2 _2040_ (.A(_1273_),
    .B(_1306_),
    .C(_1321_),
    .Y(_1376_));
 sg13g2_or2_1 _2041_ (.X(_1377_),
    .B(_1376_),
    .A(net695));
 sg13g2_nor2_1 _2042_ (.A(net702),
    .B(net694),
    .Y(_1378_));
 sg13g2_a21oi_1 _2043_ (.A1(net702),
    .A2(_1376_),
    .Y(_1379_),
    .B1(net695));
 sg13g2_and2_1 _2044_ (.A(_1276_),
    .B(_1379_),
    .X(_1380_));
 sg13g2_nand4_1 _2045_ (.B(_0007_),
    .C(_1261_),
    .A(_1162_),
    .Y(_1381_),
    .D(_1295_));
 sg13g2_nand3_1 _2046_ (.B(_1349_),
    .C(_1381_),
    .A(_1348_),
    .Y(_1382_));
 sg13g2_o21ai_1 _2047_ (.B1(_1291_),
    .Y(_1383_),
    .A1(_1300_),
    .A2(_1382_));
 sg13g2_a21oi_2 _2048_ (.B1(_1380_),
    .Y(_1384_),
    .A2(_1383_),
    .A1(net695));
 sg13g2_a21o_1 _2049_ (.A2(_1383_),
    .A1(net695),
    .B1(_1380_),
    .X(_1385_));
 sg13g2_nor2_2 _2050_ (.A(_1344_),
    .B(_1371_),
    .Y(_1386_));
 sg13g2_nand2_1 _2051_ (.Y(_1387_),
    .A(_1160_),
    .B(_1330_));
 sg13g2_a21oi_1 _2052_ (.A1(net726),
    .A2(_1351_),
    .Y(_1388_),
    .B1(_1358_));
 sg13g2_a21oi_2 _2053_ (.B1(_1386_),
    .Y(_1389_),
    .A2(_1388_),
    .A1(_1387_));
 sg13g2_a21o_1 _2054_ (.A2(_1388_),
    .A1(_1387_),
    .B1(_1386_),
    .X(_1390_));
 sg13g2_nor2_1 _2055_ (.A(net626),
    .B(_1389_),
    .Y(_1391_));
 sg13g2_nor2_2 _2056_ (.A(_1384_),
    .B(net622),
    .Y(_1392_));
 sg13g2_nor3_1 _2057_ (.A(\crp.datapath.aluSrc1SelMux.d1[0] ),
    .B(net626),
    .C(net622),
    .Y(_1393_));
 sg13g2_a21oi_1 _2058_ (.A1(\crp.controller.flags[0] ),
    .A2(_1389_),
    .Y(_1394_),
    .B1(net625));
 sg13g2_or2_1 _2059_ (.X(_1395_),
    .B(_1394_),
    .A(_1393_));
 sg13g2_nand2_2 _2060_ (.Y(_1396_),
    .A(_1331_),
    .B(_1349_));
 sg13g2_a21oi_2 _2061_ (.B1(_1280_),
    .Y(_1397_),
    .A2(_1331_),
    .A1(_1349_));
 sg13g2_a21o_1 _2062_ (.A2(_1349_),
    .A1(_1331_),
    .B1(_1280_),
    .X(_1398_));
 sg13g2_nor2_2 _2063_ (.A(net680),
    .B(net730),
    .Y(_1399_));
 sg13g2_nand2_2 _2064_ (.Y(_1400_),
    .A(net709),
    .B(net670));
 sg13g2_nor3_1 _2065_ (.A(net734),
    .B(_0028_),
    .C(net683),
    .Y(_1401_));
 sg13g2_nor2_1 _2066_ (.A(_1195_),
    .B(net682),
    .Y(_1402_));
 sg13g2_nand2_1 _2067_ (.Y(_1403_),
    .A(_0015_),
    .B(net675));
 sg13g2_a21o_1 _2068_ (.A2(net676),
    .A1(net711),
    .B1(_0027_),
    .X(_1404_));
 sg13g2_nand3b_1 _2069_ (.B(net653),
    .C(_1404_),
    .Y(_1405_),
    .A_N(_1401_));
 sg13g2_nor2_2 _2070_ (.A(_1191_),
    .B(net683),
    .Y(_1406_));
 sg13g2_nand2_1 _2071_ (.Y(_1407_),
    .A(_0012_),
    .B(net675));
 sg13g2_or3_1 _2072_ (.A(net734),
    .B(_0024_),
    .C(net682),
    .X(_1408_));
 sg13g2_a221oi_1 _2073_ (.B2(_1396_),
    .C1(_1195_),
    .B1(net697),
    .A1(net734),
    .Y(_1409_),
    .A2(_1201_));
 sg13g2_a21oi_1 _2074_ (.A1(_1408_),
    .A2(_1409_),
    .Y(_1410_),
    .B1(_1406_));
 sg13g2_and2_2 _2075_ (.A(_0020_),
    .B(net674),
    .X(_1411_));
 sg13g2_nand2_2 _2076_ (.Y(_1412_),
    .A(_0020_),
    .B(net674));
 sg13g2_nor2_1 _2077_ (.A(net733),
    .B(_0022_),
    .Y(_1413_));
 sg13g2_nor3_1 _2078_ (.A(_1195_),
    .B(net682),
    .C(_1413_),
    .Y(_1414_));
 sg13g2_o21ai_1 _2079_ (.B1(_1414_),
    .Y(_1415_),
    .A1(_0021_),
    .A2(_1399_));
 sg13g2_a21o_1 _2080_ (.A2(net676),
    .A1(net711),
    .B1(_0025_),
    .X(_1416_));
 sg13g2_a22oi_1 _2081_ (.Y(_1417_),
    .B1(net676),
    .B2(_0015_),
    .A2(_1204_),
    .A1(net710));
 sg13g2_a21oi_1 _2082_ (.A1(_1416_),
    .A2(_1417_),
    .Y(_1418_),
    .B1(net649));
 sg13g2_a221oi_1 _2083_ (.B2(_1418_),
    .C1(_1411_),
    .B1(_1415_),
    .A1(_1405_),
    .Y(_1419_),
    .A2(_1410_));
 sg13g2_nand2_1 _2084_ (.Y(_1420_),
    .A(net626),
    .B(net623));
 sg13g2_or3_1 _2085_ (.A(net731),
    .B(_0019_),
    .C(net679),
    .X(_1421_));
 sg13g2_a21o_1 _2086_ (.A2(net669),
    .A1(net709),
    .B1(_0018_),
    .X(_1422_));
 sg13g2_nand3_1 _2087_ (.B(_1421_),
    .C(_1422_),
    .A(net651),
    .Y(_1423_));
 sg13g2_or3_1 _2088_ (.A(net731),
    .B(_0014_),
    .C(net680),
    .X(_1424_));
 sg13g2_a221oi_1 _2089_ (.B2(_1396_),
    .C1(_1195_),
    .B1(net697),
    .A1(net731),
    .Y(_1425_),
    .A2(_1194_));
 sg13g2_a21oi_1 _2090_ (.A1(_1424_),
    .A2(_1425_),
    .Y(_1426_),
    .B1(net650));
 sg13g2_nor2_1 _2091_ (.A(net730),
    .B(_0010_),
    .Y(_1427_));
 sg13g2_nor3_1 _2092_ (.A(_1195_),
    .B(net680),
    .C(_1427_),
    .Y(_1428_));
 sg13g2_o21ai_1 _2093_ (.B1(_1428_),
    .Y(_1429_),
    .A1(_0009_),
    .A2(net663));
 sg13g2_a21o_1 _2094_ (.A2(net668),
    .A1(net709),
    .B1(_0016_),
    .X(_1430_));
 sg13g2_a22oi_1 _2095_ (.Y(_1431_),
    .B1(net669),
    .B2(_0015_),
    .A2(_1196_),
    .A1(net709));
 sg13g2_a21oi_1 _2096_ (.A1(_1430_),
    .A2(_1431_),
    .Y(_1432_),
    .B1(net648));
 sg13g2_a221oi_1 _2097_ (.B2(_1432_),
    .C1(_1412_),
    .B1(_1429_),
    .A1(_1423_),
    .Y(_1433_),
    .A2(_1426_));
 sg13g2_or3_1 _2098_ (.A(_1419_),
    .B(_1420_),
    .C(_1433_),
    .X(_1434_));
 sg13g2_a22oi_1 _2099_ (.Y(_1435_),
    .B1(_1395_),
    .B2(_1434_),
    .A2(_1391_),
    .A1(_0008_));
 sg13g2_nor2_1 _2100_ (.A(net614),
    .B(_1435_),
    .Y(_1436_));
 sg13g2_or3_1 _2101_ (.A(net702),
    .B(_1307_),
    .C(_1321_),
    .X(_1437_));
 sg13g2_and3_2 _2102_ (.X(_1438_),
    .A(_1318_),
    .B(_1368_),
    .C(_1437_));
 sg13g2_inv_1 _2103_ (.Y(_1439_),
    .A(_1438_));
 sg13g2_nand2_1 _2104_ (.Y(_1440_),
    .A(_1276_),
    .B(_1438_));
 sg13g2_inv_1 _2105_ (.Y(_1441_),
    .A(_1440_));
 sg13g2_nor2_2 _2106_ (.A(net612),
    .B(_1440_),
    .Y(_1442_));
 sg13g2_or2_1 _2107_ (.X(_1443_),
    .B(_1440_),
    .A(net612));
 sg13g2_nand2_1 _2108_ (.Y(_1444_),
    .A(_0030_),
    .B(net677));
 sg13g2_nor2_2 _2109_ (.A(net707),
    .B(net679),
    .Y(_1445_));
 sg13g2_nand2_2 _2110_ (.Y(_1446_),
    .A(net717),
    .B(net673));
 sg13g2_and2_2 _2111_ (.A(_0031_),
    .B(net675),
    .X(_1447_));
 sg13g2_nand2_1 _2112_ (.Y(_1448_),
    .A(_0031_),
    .B(net675));
 sg13g2_mux4_1 _2113_ (.S0(net639),
    .A0(\crp.datapath.registerFile.regs[12][2] ),
    .A1(\crp.datapath.registerFile.regs[13][2] ),
    .A2(\crp.datapath.registerFile.regs[14][2] ),
    .A3(\crp.datapath.registerFile.regs[15][2] ),
    .S1(net645),
    .X(_1449_));
 sg13g2_nor2_1 _2114_ (.A(_1447_),
    .B(_1449_),
    .Y(_1450_));
 sg13g2_and2_2 _2115_ (.A(_0032_),
    .B(net675),
    .X(_1451_));
 sg13g2_nand2_2 _2116_ (.Y(_1452_),
    .A(_0032_),
    .B(net677));
 sg13g2_mux2_1 _2117_ (.A0(\crp.datapath.registerFile.regs[10][2] ),
    .A1(\crp.datapath.registerFile.regs[11][2] ),
    .S(net638),
    .X(_1453_));
 sg13g2_a21oi_1 _2118_ (.A1(net708),
    .A2(_1219_),
    .Y(_1454_),
    .B1(net645));
 sg13g2_o21ai_1 _2119_ (.B1(_1454_),
    .Y(_1455_),
    .A1(\crp.datapath.registerFile.regs[8][2] ),
    .A2(net638));
 sg13g2_a21oi_1 _2120_ (.A1(net644),
    .A2(_1453_),
    .Y(_1456_),
    .B1(net637));
 sg13g2_a21oi_1 _2121_ (.A1(_1455_),
    .A2(_1456_),
    .Y(_1457_),
    .B1(_1450_));
 sg13g2_mux2_1 _2122_ (.A0(\crp.datapath.registerFile.regs[6][2] ),
    .A1(\crp.datapath.registerFile.regs[7][2] ),
    .S(net638),
    .X(_1458_));
 sg13g2_a21oi_1 _2123_ (.A1(net706),
    .A2(_1218_),
    .Y(_1459_),
    .B1(net642));
 sg13g2_o21ai_1 _2124_ (.B1(_1459_),
    .Y(_1460_),
    .A1(\crp.datapath.registerFile.regs[4][2] ),
    .A2(net638));
 sg13g2_a21oi_1 _2125_ (.A1(net642),
    .A2(_1458_),
    .Y(_1461_),
    .B1(_1447_));
 sg13g2_mux2_1 _2126_ (.A0(\crp.datapath.registerFile.regs[2][2] ),
    .A1(\crp.datapath.registerFile.regs[3][2] ),
    .S(net638),
    .X(_1462_));
 sg13g2_a21oi_1 _2127_ (.A1(net706),
    .A2(_1217_),
    .Y(_1463_),
    .B1(net642));
 sg13g2_o21ai_1 _2128_ (.B1(_1463_),
    .Y(_1464_),
    .A1(\crp.datapath.registerFile.regs[0][2] ),
    .A2(net638));
 sg13g2_a21oi_1 _2129_ (.A1(net642),
    .A2(_1462_),
    .Y(_1465_),
    .B1(net634));
 sg13g2_a221oi_1 _2130_ (.B2(_1465_),
    .C1(net633),
    .B1(_1464_),
    .A1(_1460_),
    .Y(_1466_),
    .A2(_1461_));
 sg13g2_a21o_2 _2131_ (.A2(_1457_),
    .A1(net633),
    .B1(_1466_),
    .X(_1467_));
 sg13g2_nand2_1 _2132_ (.Y(_1468_),
    .A(net725),
    .B(_1277_));
 sg13g2_o21ai_1 _2133_ (.B1(_1468_),
    .Y(_1469_),
    .A1(_1160_),
    .A2(_1438_));
 sg13g2_a21oi_1 _2134_ (.A1(_1442_),
    .A2(_1467_),
    .Y(_1470_),
    .B1(_1469_));
 sg13g2_a21o_2 _2135_ (.A2(_1467_),
    .A1(_1442_),
    .B1(_1469_),
    .X(_1471_));
 sg13g2_mux4_1 _2136_ (.S0(net639),
    .A0(\crp.datapath.registerFile.regs[12][1] ),
    .A1(\crp.datapath.registerFile.regs[13][1] ),
    .A2(\crp.datapath.registerFile.regs[14][1] ),
    .A3(\crp.datapath.registerFile.regs[15][1] ),
    .S1(net646),
    .X(_1472_));
 sg13g2_nand2b_1 _2137_ (.Y(_1473_),
    .B(net637),
    .A_N(_1472_));
 sg13g2_and3_1 _2138_ (.X(_1474_),
    .A(net718),
    .B(\crp.datapath.registerFile.regs[10][1] ),
    .C(net674));
 sg13g2_a21oi_1 _2139_ (.A1(net718),
    .A2(net674),
    .Y(_1475_),
    .B1(_1212_));
 sg13g2_o21ai_1 _2140_ (.B1(net645),
    .Y(_1476_),
    .A1(_1474_),
    .A2(_1475_));
 sg13g2_nand3b_1 _2141_ (.B(net675),
    .C(net718),
    .Y(_1477_),
    .A_N(\crp.datapath.registerFile.regs[8][1] ));
 sg13g2_nor2_1 _2142_ (.A(net718),
    .B(\crp.datapath.registerFile.regs[9][1] ),
    .Y(_1478_));
 sg13g2_nor3_1 _2143_ (.A(net705),
    .B(net682),
    .C(_1478_),
    .Y(_1479_));
 sg13g2_a21oi_1 _2144_ (.A1(_1477_),
    .A2(_1479_),
    .Y(_1480_),
    .B1(net636));
 sg13g2_a21oi_2 _2145_ (.B1(_1451_),
    .Y(_1481_),
    .A2(_1480_),
    .A1(_1476_));
 sg13g2_a21oi_1 _2146_ (.A1(net714),
    .A2(net671),
    .Y(_1482_),
    .B1(\crp.datapath.registerFile.regs[7][1] ));
 sg13g2_a221oi_1 _2147_ (.B2(_1211_),
    .C1(_1482_),
    .B1(net640),
    .A1(_0030_),
    .Y(_1483_),
    .A2(net671));
 sg13g2_nor3_1 _2148_ (.A(net707),
    .B(\crp.datapath.registerFile.regs[4][1] ),
    .C(net681),
    .Y(_1484_));
 sg13g2_nor2_1 _2149_ (.A(net714),
    .B(\crp.datapath.registerFile.regs[5][1] ),
    .Y(_1485_));
 sg13g2_nor3_1 _2150_ (.A(net644),
    .B(_1484_),
    .C(_1485_),
    .Y(_1486_));
 sg13g2_or3_1 _2151_ (.A(_1447_),
    .B(_1483_),
    .C(_1486_),
    .X(_1487_));
 sg13g2_and3_1 _2152_ (.X(_1488_),
    .A(net716),
    .B(\crp.datapath.registerFile.regs[2][1] ),
    .C(net672));
 sg13g2_a21oi_1 _2153_ (.A1(net716),
    .A2(net672),
    .Y(_1489_),
    .B1(_1209_));
 sg13g2_o21ai_1 _2154_ (.B1(net644),
    .Y(_1490_),
    .A1(_1488_),
    .A2(_1489_));
 sg13g2_nand3b_1 _2155_ (.B(net672),
    .C(net716),
    .Y(_1491_),
    .A_N(\crp.datapath.registerFile.regs[0][1] ));
 sg13g2_nor2_1 _2156_ (.A(net716),
    .B(\crp.datapath.registerFile.regs[1][1] ),
    .Y(_1492_));
 sg13g2_nor3_1 _2157_ (.A(net704),
    .B(net681),
    .C(_1492_),
    .Y(_1493_));
 sg13g2_a21oi_1 _2158_ (.A1(_1491_),
    .A2(_1493_),
    .Y(_1494_),
    .B1(net635));
 sg13g2_a21oi_1 _2159_ (.A1(_1490_),
    .A2(_1494_),
    .Y(_1495_),
    .B1(_1452_));
 sg13g2_a22oi_1 _2160_ (.Y(_1496_),
    .B1(_1487_),
    .B2(_1495_),
    .A2(_1481_),
    .A1(_1473_));
 sg13g2_a22oi_1 _2161_ (.Y(_1497_),
    .B1(_1439_),
    .B2(net727),
    .A2(_1277_),
    .A1(net726));
 sg13g2_o21ai_1 _2162_ (.B1(_1497_),
    .Y(_1498_),
    .A1(_1443_),
    .A2(_1496_));
 sg13g2_inv_2 _2163_ (.Y(_1499_),
    .A(net590));
 sg13g2_nor3_2 _2164_ (.A(net728),
    .B(net699),
    .C(_1268_),
    .Y(_1500_));
 sg13g2_nor3_1 _2165_ (.A(net727),
    .B(net698),
    .C(_1298_),
    .Y(_1501_));
 sg13g2_nor3_1 _2166_ (.A(net698),
    .B(_1281_),
    .C(_1288_),
    .Y(_1502_));
 sg13g2_nor4_1 _2167_ (.A(net722),
    .B(net724),
    .C(net698),
    .D(_1286_),
    .Y(_1503_));
 sg13g2_or3_1 _2168_ (.A(_1501_),
    .B(_1502_),
    .C(_1503_),
    .X(_1504_));
 sg13g2_a21oi_2 _2169_ (.B1(_1500_),
    .Y(_1505_),
    .A2(_1504_),
    .A1(net694));
 sg13g2_inv_1 _2170_ (.Y(_1506_),
    .A(_1505_));
 sg13g2_nand2_1 _2171_ (.Y(_1507_),
    .A(_1263_),
    .B(net694));
 sg13g2_nor4_1 _2172_ (.A(_1158_),
    .B(_1283_),
    .C(_1285_),
    .D(_1507_),
    .Y(_1508_));
 sg13g2_a21oi_2 _2173_ (.B1(_1508_),
    .Y(_1509_),
    .A2(_1304_),
    .A1(_1270_));
 sg13g2_or2_1 _2174_ (.X(_1510_),
    .B(_1283_),
    .A(net725));
 sg13g2_nand4_1 _2175_ (.B(_1281_),
    .C(_1288_),
    .A(_1263_),
    .Y(_1511_),
    .D(_1510_));
 sg13g2_nor2_1 _2176_ (.A(_1329_),
    .B(_1502_),
    .Y(_1512_));
 sg13g2_a21oi_1 _2177_ (.A1(_1511_),
    .A2(_1512_),
    .Y(_1513_),
    .B1(_1280_));
 sg13g2_nor3_1 _2178_ (.A(net728),
    .B(net699),
    .C(_1273_),
    .Y(_1514_));
 sg13g2_nor4_2 _2179_ (.A(_1267_),
    .B(_1344_),
    .C(_1513_),
    .Y(_1515_),
    .D(_1514_));
 sg13g2_nor2_1 _2180_ (.A(net621),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_nand2_2 _2181_ (.Y(_1517_),
    .A(_1505_),
    .B(_1516_));
 sg13g2_mux4_1 _2182_ (.S0(net639),
    .A0(_1202_),
    .A1(_1203_),
    .A2(_1205_),
    .A3(_1206_),
    .S1(net646),
    .X(_1518_));
 sg13g2_nor3_1 _2183_ (.A(_1199_),
    .B(net708),
    .C(net682),
    .Y(_1519_));
 sg13g2_a21oi_1 _2184_ (.A1(net720),
    .A2(net675),
    .Y(_1520_),
    .B1(_1200_));
 sg13g2_o21ai_1 _2185_ (.B1(net645),
    .Y(_1521_),
    .A1(_1519_),
    .A2(_1520_));
 sg13g2_nand3b_1 _2186_ (.B(net720),
    .C(net677),
    .Y(_1522_),
    .A_N(\crp.datapath.registerFile.regs[8][0] ));
 sg13g2_nor2_1 _2187_ (.A(\crp.datapath.registerFile.regs[9][0] ),
    .B(net720),
    .Y(_1523_));
 sg13g2_nor3_1 _2188_ (.A(net705),
    .B(net682),
    .C(_1523_),
    .Y(_1524_));
 sg13g2_a21oi_1 _2189_ (.A1(_1522_),
    .A2(_1524_),
    .Y(_1525_),
    .B1(net637));
 sg13g2_a221oi_1 _2190_ (.B2(_1525_),
    .C1(_1451_),
    .B1(_1521_),
    .A1(_1518_),
    .Y(_1526_),
    .A2(net636));
 sg13g2_nor3_1 _2191_ (.A(_1197_),
    .B(net706),
    .C(net679),
    .Y(_1527_));
 sg13g2_a21oi_1 _2192_ (.A1(net713),
    .A2(net669),
    .Y(_1528_),
    .B1(_1198_));
 sg13g2_o21ai_1 _2193_ (.B1(net644),
    .Y(_1529_),
    .A1(_1527_),
    .A2(_1528_));
 sg13g2_nand3b_1 _2194_ (.B(net715),
    .C(net668),
    .Y(_1530_),
    .A_N(\crp.datapath.registerFile.regs[4][0] ));
 sg13g2_nor2_1 _2195_ (.A(\crp.datapath.registerFile.regs[5][0] ),
    .B(net715),
    .Y(_1531_));
 sg13g2_nor3_1 _2196_ (.A(net704),
    .B(net680),
    .C(_1531_),
    .Y(_1532_));
 sg13g2_a21oi_1 _2197_ (.A1(_1530_),
    .A2(_1532_),
    .Y(_1533_),
    .B1(_1447_));
 sg13g2_nor3_1 _2198_ (.A(_1192_),
    .B(net706),
    .C(net680),
    .Y(_1534_));
 sg13g2_a21oi_1 _2199_ (.A1(net715),
    .A2(net669),
    .Y(_1535_),
    .B1(_1193_));
 sg13g2_o21ai_1 _2200_ (.B1(net642),
    .Y(_1536_),
    .A1(_1534_),
    .A2(_1535_));
 sg13g2_nand3b_1 _2201_ (.B(net715),
    .C(net669),
    .Y(_1537_),
    .A_N(\crp.datapath.registerFile.regs[0][0] ));
 sg13g2_nor2_1 _2202_ (.A(\crp.datapath.registerFile.regs[1][0] ),
    .B(net716),
    .Y(_1538_));
 sg13g2_nor3_1 _2203_ (.A(net704),
    .B(net680),
    .C(_1538_),
    .Y(_1539_));
 sg13g2_a21oi_1 _2204_ (.A1(_1537_),
    .A2(_1539_),
    .Y(_1540_),
    .B1(net634));
 sg13g2_a221oi_1 _2205_ (.B2(_1540_),
    .C1(net633),
    .B1(_1536_),
    .A1(_1529_),
    .Y(_1541_),
    .A2(_1533_));
 sg13g2_or3_1 _2206_ (.A(_1526_),
    .B(net611),
    .C(_1541_),
    .X(_1542_));
 sg13g2_a22oi_1 _2207_ (.Y(_1543_),
    .B1(_1441_),
    .B2(_1542_),
    .A2(_1277_),
    .A1(net727));
 sg13g2_nand2_1 _2208_ (.Y(_1544_),
    .A(_1435_),
    .B(net587));
 sg13g2_nor3_2 _2209_ (.A(net591),
    .B(_1517_),
    .C(_1544_),
    .Y(_1545_));
 sg13g2_or2_1 _2210_ (.X(_1546_),
    .B(net621),
    .A(_1505_));
 sg13g2_and2_2 _2211_ (.A(_0050_),
    .B(net610),
    .X(_1547_));
 sg13g2_nand2_1 _2212_ (.Y(_1548_),
    .A(_0050_),
    .B(net610));
 sg13g2_nor2_1 _2213_ (.A(_0055_),
    .B(net663),
    .Y(_1549_));
 sg13g2_nor2_1 _2214_ (.A(net729),
    .B(_0056_),
    .Y(_1550_));
 sg13g2_o21ai_1 _2215_ (.B1(net651),
    .Y(_1551_),
    .A1(_1549_),
    .A2(_1550_));
 sg13g2_or2_1 _2216_ (.X(_1552_),
    .B(_0052_),
    .A(net729));
 sg13g2_o21ai_1 _2217_ (.B1(_1552_),
    .Y(_1553_),
    .A1(_0051_),
    .A2(net663));
 sg13g2_a21oi_1 _2218_ (.A1(net657),
    .A2(_1553_),
    .Y(_1554_),
    .B1(net648));
 sg13g2_nand2_1 _2219_ (.Y(_1555_),
    .A(_0057_),
    .B(net658));
 sg13g2_a21oi_1 _2220_ (.A1(_0058_),
    .A2(net663),
    .Y(_1556_),
    .B1(net657));
 sg13g2_nand2b_1 _2221_ (.Y(_1557_),
    .B(net729),
    .A_N(_0053_));
 sg13g2_o21ai_1 _2222_ (.B1(_1557_),
    .Y(_1558_),
    .A1(_0054_),
    .A2(net658));
 sg13g2_a22oi_1 _2223_ (.Y(_1559_),
    .B1(_1558_),
    .B2(net657),
    .A2(_1556_),
    .A1(_1555_));
 sg13g2_a221oi_1 _2224_ (.B2(net648),
    .C1(_1412_),
    .B1(_1559_),
    .A1(_1551_),
    .Y(_1560_),
    .A2(_1554_));
 sg13g2_nor2_1 _2225_ (.A(_0063_),
    .B(net664),
    .Y(_1561_));
 sg13g2_nor2_1 _2226_ (.A(net733),
    .B(_0064_),
    .Y(_1562_));
 sg13g2_o21ai_1 _2227_ (.B1(net653),
    .Y(_1563_),
    .A1(_1561_),
    .A2(_1562_));
 sg13g2_or2_1 _2228_ (.X(_1564_),
    .B(_0060_),
    .A(net733));
 sg13g2_o21ai_1 _2229_ (.B1(_1564_),
    .Y(_1565_),
    .A1(_0059_),
    .A2(net664));
 sg13g2_a21oi_1 _2230_ (.A1(net656),
    .A2(_1565_),
    .Y(_1566_),
    .B1(net649));
 sg13g2_nand2_1 _2231_ (.Y(_1567_),
    .A(_0065_),
    .B(net661));
 sg13g2_a21oi_1 _2232_ (.A1(_0066_),
    .A2(net664),
    .Y(_1568_),
    .B1(net656));
 sg13g2_nand2b_1 _2233_ (.Y(_1569_),
    .B(net733),
    .A_N(_0061_));
 sg13g2_o21ai_1 _2234_ (.B1(_1569_),
    .Y(_1570_),
    .A1(_0062_),
    .A2(net659));
 sg13g2_a221oi_1 _2235_ (.B2(net656),
    .C1(_1406_),
    .B1(_1570_),
    .A1(_1567_),
    .Y(_1571_),
    .A2(_1568_));
 sg13g2_a221oi_1 _2236_ (.B2(_1566_),
    .C1(_1571_),
    .B1(_1563_),
    .A1(_0020_),
    .Y(_1572_),
    .A2(net677));
 sg13g2_or3_1 _2237_ (.A(net624),
    .B(_1560_),
    .C(_1572_),
    .X(_1573_));
 sg13g2_nand3_1 _2238_ (.B(net626),
    .C(_1389_),
    .A(\crp.controller.flags[2] ),
    .Y(_1574_));
 sg13g2_o21ai_1 _2239_ (.B1(_1574_),
    .Y(_1575_),
    .A1(_1179_),
    .A2(net626));
 sg13g2_a21oi_2 _2240_ (.B1(_1575_),
    .Y(_1576_),
    .A2(_1573_),
    .A1(net623));
 sg13g2_a21o_1 _2241_ (.A2(_1573_),
    .A1(net623),
    .B1(_1575_),
    .X(_1577_));
 sg13g2_nor2_2 _2242_ (.A(_1547_),
    .B(_1576_),
    .Y(_1578_));
 sg13g2_o21ai_1 _2243_ (.B1(net588),
    .Y(_1579_),
    .A1(_1547_),
    .A2(_1576_));
 sg13g2_nor2_1 _2244_ (.A(_0072_),
    .B(net662),
    .Y(_1580_));
 sg13g2_nor2_1 _2245_ (.A(net729),
    .B(_0073_),
    .Y(_1581_));
 sg13g2_o21ai_1 _2246_ (.B1(net651),
    .Y(_1582_),
    .A1(_1580_),
    .A2(_1581_));
 sg13g2_nand2_1 _2247_ (.Y(_1583_),
    .A(net709),
    .B(_1220_));
 sg13g2_o21ai_1 _2248_ (.B1(_1583_),
    .Y(_1584_),
    .A1(_0068_),
    .A2(net662));
 sg13g2_a21oi_1 _2249_ (.A1(net657),
    .A2(_1584_),
    .Y(_0345_),
    .B1(net648));
 sg13g2_nand2_1 _2250_ (.Y(_0346_),
    .A(_0074_),
    .B(net658));
 sg13g2_a21oi_1 _2251_ (.A1(_0075_),
    .A2(net662),
    .Y(_0347_),
    .B1(net657));
 sg13g2_nand2b_1 _2252_ (.Y(_0348_),
    .B(net729),
    .A_N(_0070_));
 sg13g2_o21ai_1 _2253_ (.B1(_0348_),
    .Y(_0349_),
    .A1(_0071_),
    .A2(net658));
 sg13g2_a22oi_1 _2254_ (.Y(_0350_),
    .B1(_0349_),
    .B2(net657),
    .A2(_0347_),
    .A1(_0346_));
 sg13g2_a221oi_1 _2255_ (.B2(net648),
    .C1(_1412_),
    .B1(_0350_),
    .A1(_1582_),
    .Y(_0351_),
    .A2(_0345_));
 sg13g2_or2_1 _2256_ (.X(_0352_),
    .B(_0081_),
    .A(net733));
 sg13g2_o21ai_1 _2257_ (.B1(_0352_),
    .Y(_0353_),
    .A1(_0080_),
    .A2(net664));
 sg13g2_nor2_1 _2258_ (.A(_0076_),
    .B(net664),
    .Y(_0354_));
 sg13g2_nor2_1 _2259_ (.A(net733),
    .B(_0077_),
    .Y(_0355_));
 sg13g2_o21ai_1 _2260_ (.B1(net656),
    .Y(_0356_),
    .A1(_0354_),
    .A2(_0355_));
 sg13g2_a21oi_1 _2261_ (.A1(net653),
    .A2(_0353_),
    .Y(_0357_),
    .B1(net649));
 sg13g2_nand2_1 _2262_ (.Y(_0358_),
    .A(_0082_),
    .B(net661));
 sg13g2_a21oi_1 _2263_ (.A1(_0083_),
    .A2(net664),
    .Y(_0359_),
    .B1(net656));
 sg13g2_nand2b_1 _2264_ (.Y(_0360_),
    .B(net733),
    .A_N(_0078_));
 sg13g2_o21ai_1 _2265_ (.B1(_0360_),
    .Y(_0361_),
    .A1(_0079_),
    .A2(net659));
 sg13g2_a221oi_1 _2266_ (.B2(net656),
    .C1(_1406_),
    .B1(_0361_),
    .A1(_0358_),
    .Y(_0362_),
    .A2(_0359_));
 sg13g2_a221oi_1 _2267_ (.B2(_0357_),
    .C1(_0362_),
    .B1(_0356_),
    .A1(_0020_),
    .Y(_0363_),
    .A2(net677));
 sg13g2_or3_1 _2268_ (.A(net624),
    .B(_0351_),
    .C(_0363_),
    .X(_0364_));
 sg13g2_nor3_1 _2269_ (.A(_1150_),
    .B(net625),
    .C(net622),
    .Y(_0365_));
 sg13g2_a221oi_1 _2270_ (.B2(_0364_),
    .C1(_0365_),
    .B1(net623),
    .A1(\crp.datapath.aluSrc1SelMux.d1[3] ),
    .Y(_0366_),
    .A2(net625));
 sg13g2_a21oi_1 _2271_ (.A1(_0067_),
    .A2(net609),
    .Y(_0367_),
    .B1(_0366_));
 sg13g2_inv_1 _2272_ (.Y(_0368_),
    .A(net572));
 sg13g2_mux2_1 _2273_ (.A0(net572),
    .A1(_1578_),
    .S(net587),
    .X(_0369_));
 sg13g2_nor3_1 _2274_ (.A(\crp.datapath.aluSrc1SelMux.d1[1] ),
    .B(net626),
    .C(net622),
    .Y(_0370_));
 sg13g2_a21oi_1 _2275_ (.A1(\crp.controller.flags[1] ),
    .A2(_1389_),
    .Y(_0371_),
    .B1(net625));
 sg13g2_or2_1 _2276_ (.X(_0372_),
    .B(_0371_),
    .A(_0370_));
 sg13g2_a21o_1 _2277_ (.A2(net673),
    .A1(net711),
    .B1(_0044_),
    .X(_0373_));
 sg13g2_or3_1 _2278_ (.A(net734),
    .B(_0045_),
    .C(net682),
    .X(_0374_));
 sg13g2_nand3_1 _2279_ (.B(_0373_),
    .C(_0374_),
    .A(net649),
    .Y(_0375_));
 sg13g2_a21o_1 _2280_ (.A2(net675),
    .A1(net710),
    .B1(_0042_),
    .X(_0376_));
 sg13g2_nor2_1 _2281_ (.A(net734),
    .B(_0043_),
    .Y(_0377_));
 sg13g2_nor3_1 _2282_ (.A(_1191_),
    .B(net682),
    .C(_0377_),
    .Y(_0378_));
 sg13g2_a21oi_1 _2283_ (.A1(_0376_),
    .A2(_0378_),
    .Y(_0379_),
    .B1(net654));
 sg13g2_mux4_1 _2284_ (.S0(net661),
    .A0(_1213_),
    .A1(_1214_),
    .A2(_1215_),
    .A3(_1216_),
    .S1(net648),
    .X(_0380_));
 sg13g2_a221oi_1 _2285_ (.B2(net653),
    .C1(_1411_),
    .B1(_0380_),
    .A1(_0375_),
    .Y(_0381_),
    .A2(_0379_));
 sg13g2_or3_1 _2286_ (.A(net732),
    .B(_0041_),
    .C(net681),
    .X(_0382_));
 sg13g2_a21o_1 _2287_ (.A2(net672),
    .A1(net712),
    .B1(_0040_),
    .X(_0383_));
 sg13g2_nand3_1 _2288_ (.B(_0382_),
    .C(_0383_),
    .A(net652),
    .Y(_0384_));
 sg13g2_or3_1 _2289_ (.A(net731),
    .B(_0037_),
    .C(net681),
    .X(_0385_));
 sg13g2_a221oi_1 _2290_ (.B2(_1396_),
    .C1(_1195_),
    .B1(net697),
    .A1(net731),
    .Y(_0386_),
    .A2(_1210_));
 sg13g2_a21oi_1 _2291_ (.A1(_0385_),
    .A2(_0386_),
    .Y(_0387_),
    .B1(net650));
 sg13g2_a21o_1 _2292_ (.A2(net671),
    .A1(net712),
    .B1(_0038_),
    .X(_0388_));
 sg13g2_or2_1 _2293_ (.X(_0389_),
    .B(_0039_),
    .A(net731));
 sg13g2_nand3_1 _2294_ (.B(_0388_),
    .C(_0389_),
    .A(net651),
    .Y(_0390_));
 sg13g2_a21o_1 _2295_ (.A2(net671),
    .A1(net709),
    .B1(_0034_),
    .X(_0391_));
 sg13g2_nor2_1 _2296_ (.A(net731),
    .B(_0035_),
    .Y(_0392_));
 sg13g2_nor3_1 _2297_ (.A(_1195_),
    .B(net681),
    .C(_0392_),
    .Y(_0393_));
 sg13g2_a21oi_1 _2298_ (.A1(_0391_),
    .A2(_0393_),
    .Y(_0394_),
    .B1(net648));
 sg13g2_a221oi_1 _2299_ (.B2(_0394_),
    .C1(_1412_),
    .B1(_0390_),
    .A1(_0384_),
    .Y(_0395_),
    .A2(_0387_));
 sg13g2_or3_1 _2300_ (.A(_1420_),
    .B(_0381_),
    .C(_0395_),
    .X(_0396_));
 sg13g2_a22oi_1 _2301_ (.Y(_0397_),
    .B1(_0372_),
    .B2(_0396_),
    .A2(net610),
    .A1(_0033_));
 sg13g2_nor2_1 _2302_ (.A(net588),
    .B(net585),
    .Y(_0398_));
 sg13g2_nor2b_1 _2303_ (.A(_1435_),
    .B_N(net588),
    .Y(_0399_));
 sg13g2_nor3_1 _2304_ (.A(net591),
    .B(_0398_),
    .C(_0399_),
    .Y(_0400_));
 sg13g2_a21oi_1 _2305_ (.A1(net591),
    .A2(_0369_),
    .Y(_0401_),
    .B1(_0400_));
 sg13g2_nor2_1 _2306_ (.A(_1546_),
    .B(_0401_),
    .Y(_0402_));
 sg13g2_o21ai_1 _2307_ (.B1(net577),
    .Y(_0403_),
    .A1(_1545_),
    .A2(_0402_));
 sg13g2_inv_1 _2308_ (.Y(_0404_),
    .A(_0403_));
 sg13g2_nor2_1 _2309_ (.A(net577),
    .B(_1546_),
    .Y(_0405_));
 sg13g2_mux4_1 _2310_ (.S0(net661),
    .A0(_0130_),
    .A1(_0129_),
    .A2(_0134_),
    .A3(_0133_),
    .S1(net653),
    .X(_0406_));
 sg13g2_nor2_1 _2311_ (.A(net650),
    .B(_0406_),
    .Y(_0407_));
 sg13g2_a22oi_1 _2312_ (.Y(_0408_),
    .B1(_1242_),
    .B2(net661),
    .A2(_1241_),
    .A1(net711));
 sg13g2_nand2b_1 _2313_ (.Y(_0409_),
    .B(net661),
    .A_N(_0127_));
 sg13g2_a21oi_1 _2314_ (.A1(net711),
    .A2(_1239_),
    .Y(_0410_),
    .B1(net653));
 sg13g2_a221oi_1 _2315_ (.B2(_0410_),
    .C1(net649),
    .B1(_0409_),
    .A1(net653),
    .Y(_0411_),
    .A2(_0408_));
 sg13g2_o21ai_1 _2316_ (.B1(_1412_),
    .Y(_0412_),
    .A1(_0407_),
    .A2(_0411_));
 sg13g2_nor3_1 _2317_ (.A(net730),
    .B(_1238_),
    .C(net679),
    .Y(_0413_));
 sg13g2_a21oi_1 _2318_ (.A1(_0121_),
    .A2(net658),
    .Y(_0414_),
    .B1(_0413_));
 sg13g2_and3_1 _2319_ (.X(_0415_),
    .A(net709),
    .B(_0126_),
    .C(net670));
 sg13g2_a21oi_1 _2320_ (.A1(_0125_),
    .A2(net658),
    .Y(_0416_),
    .B1(_0415_));
 sg13g2_or2_1 _2321_ (.X(_0417_),
    .B(_0124_),
    .A(net729));
 sg13g2_o21ai_1 _2322_ (.B1(_0417_),
    .Y(_0418_),
    .A1(_0123_),
    .A2(net662));
 sg13g2_or2_1 _2323_ (.X(_0419_),
    .B(_0120_),
    .A(net730));
 sg13g2_o21ai_1 _2324_ (.B1(_0419_),
    .Y(_0420_),
    .A1(_0119_),
    .A2(net662));
 sg13g2_mux4_1 _2325_ (.S0(net651),
    .A0(_0414_),
    .A1(_0416_),
    .A2(_0420_),
    .A3(_0418_),
    .S1(net650),
    .X(_0421_));
 sg13g2_a21oi_1 _2326_ (.A1(_1411_),
    .A2(_0421_),
    .Y(_0422_),
    .B1(net624));
 sg13g2_a21oi_1 _2327_ (.A1(\crp.datapath.aluSrc1SelMux.d1[6] ),
    .A2(net624),
    .Y(_0423_),
    .B1(net622));
 sg13g2_a221oi_1 _2328_ (.B2(_0422_),
    .C1(_0423_),
    .B1(_0412_),
    .A1(_0118_),
    .Y(_0424_),
    .A2(net610));
 sg13g2_nor2b_1 _2329_ (.A(_0424_),
    .B_N(net586),
    .Y(_0425_));
 sg13g2_inv_1 _2330_ (.Y(_0426_),
    .A(_0425_));
 sg13g2_mux4_1 _2331_ (.S0(net660),
    .A0(_0147_),
    .A1(_0146_),
    .A2(_0151_),
    .A3(_0150_),
    .S1(net654),
    .X(_0427_));
 sg13g2_a22oi_1 _2332_ (.Y(_0428_),
    .B1(_1252_),
    .B2(net660),
    .A2(_1251_),
    .A1(net710));
 sg13g2_a22oi_1 _2333_ (.Y(_0429_),
    .B1(_1249_),
    .B2(net660),
    .A2(_1248_),
    .A1(net710));
 sg13g2_mux2_1 _2334_ (.A0(_0428_),
    .A1(_0429_),
    .S(net657),
    .X(_0430_));
 sg13g2_mux4_1 _2335_ (.S0(net659),
    .A0(_0139_),
    .A1(_0138_),
    .A2(_0143_),
    .A3(_0142_),
    .S1(net651),
    .X(_0431_));
 sg13g2_or2_1 _2336_ (.X(_0432_),
    .B(_0141_),
    .A(net732));
 sg13g2_o21ai_1 _2337_ (.B1(_0432_),
    .Y(_0433_),
    .A1(_0140_),
    .A2(net662));
 sg13g2_o21ai_1 _2338_ (.B1(_1246_),
    .Y(_0434_),
    .A1(net731),
    .A2(net679));
 sg13g2_nand2_1 _2339_ (.Y(_0435_),
    .A(net709),
    .B(_1245_));
 sg13g2_a21oi_1 _2340_ (.A1(_0434_),
    .A2(_0435_),
    .Y(_0436_),
    .B1(net652));
 sg13g2_a21oi_2 _2341_ (.B1(_0436_),
    .Y(_0437_),
    .A2(_0433_),
    .A1(net652));
 sg13g2_mux4_1 _2342_ (.S0(net650),
    .A0(_0427_),
    .A1(_0430_),
    .A2(_0431_),
    .A3(_0437_),
    .S1(_1411_),
    .X(_0438_));
 sg13g2_a21oi_1 _2343_ (.A1(\crp.datapath.aluSrc1SelMux.d1[7] ),
    .A2(net624),
    .Y(_0439_),
    .B1(net622));
 sg13g2_a221oi_1 _2344_ (.B2(net626),
    .C1(_0439_),
    .B1(_0438_),
    .A1(_0135_),
    .Y(_0440_),
    .A2(net610));
 sg13g2_o21ai_1 _2345_ (.B1(_0426_),
    .Y(_0441_),
    .A1(net587),
    .A2(net584));
 sg13g2_mux4_1 _2346_ (.S0(net660),
    .A0(_0096_),
    .A1(_0095_),
    .A2(_0100_),
    .A3(_0099_),
    .S1(net654),
    .X(_0442_));
 sg13g2_nor2_1 _2347_ (.A(net650),
    .B(_0442_),
    .Y(_0443_));
 sg13g2_nand2b_1 _2348_ (.Y(_0444_),
    .B(net660),
    .A_N(_0097_));
 sg13g2_a21oi_1 _2349_ (.A1(net710),
    .A2(_1228_),
    .Y(_0445_),
    .B1(net656));
 sg13g2_nand2b_1 _2350_ (.Y(_0446_),
    .B(net660),
    .A_N(_0093_));
 sg13g2_a21oi_1 _2351_ (.A1(net710),
    .A2(_1226_),
    .Y(_0447_),
    .B1(net653));
 sg13g2_a221oi_1 _2352_ (.B2(_0446_),
    .C1(net648),
    .B1(_0447_),
    .A1(_0444_),
    .Y(_0448_),
    .A2(_0445_));
 sg13g2_o21ai_1 _2353_ (.B1(_1412_),
    .Y(_0449_),
    .A1(_0448_),
    .A2(_0443_));
 sg13g2_nor3_1 _2354_ (.A(net729),
    .B(_1223_),
    .C(net679),
    .Y(_0450_));
 sg13g2_a21oi_1 _2355_ (.A1(_0087_),
    .A2(net658),
    .Y(_0451_),
    .B1(_0450_));
 sg13g2_mux2_1 _2356_ (.A0(_1224_),
    .A1(_1225_),
    .S(net658),
    .X(_0452_));
 sg13g2_or2_1 _2357_ (.X(_0453_),
    .B(_0090_),
    .A(net729));
 sg13g2_o21ai_1 _2358_ (.B1(_0453_),
    .Y(_0454_),
    .A1(net662),
    .A2(_0089_));
 sg13g2_or2_1 _2359_ (.X(_0455_),
    .B(_0086_),
    .A(net730));
 sg13g2_o21ai_1 _2360_ (.B1(_0455_),
    .Y(_0456_),
    .A1(_0085_),
    .A2(net662));
 sg13g2_mux4_1 _2361_ (.S0(net651),
    .A0(_0451_),
    .A1(_0452_),
    .A2(_0456_),
    .A3(_0454_),
    .S1(net650),
    .X(_0457_));
 sg13g2_a21oi_2 _2362_ (.B1(net624),
    .Y(_0458_),
    .A2(_1411_),
    .A1(_0457_));
 sg13g2_a21oi_1 _2363_ (.A1(\crp.datapath.aluSrc1SelMux.d1[4] ),
    .A2(net624),
    .Y(_0459_),
    .B1(net622));
 sg13g2_a221oi_1 _2364_ (.B2(_0449_),
    .C1(_0459_),
    .B1(_0458_),
    .A1(_0084_),
    .Y(_0460_),
    .A2(net610));
 sg13g2_nand2b_1 _2365_ (.Y(_0461_),
    .B(net586),
    .A_N(_0460_));
 sg13g2_mux4_1 _2366_ (.S0(net661),
    .A0(_0113_),
    .A1(_0112_),
    .A2(_0117_),
    .A3(_0116_),
    .S1(net654),
    .X(_0462_));
 sg13g2_a22oi_1 _2367_ (.Y(_0463_),
    .B1(_1235_),
    .B2(net660),
    .A2(_1234_),
    .A1(net710));
 sg13g2_a22oi_1 _2368_ (.Y(_0464_),
    .B1(_1232_),
    .B2(net660),
    .A2(_1231_),
    .A1(net710));
 sg13g2_mux2_1 _2369_ (.A0(_0463_),
    .A1(_0464_),
    .S(net656),
    .X(_0465_));
 sg13g2_mux4_1 _2370_ (.S0(net659),
    .A0(_0105_),
    .A1(_0104_),
    .A2(_0109_),
    .A3(_0108_),
    .S1(net652),
    .X(_0466_));
 sg13g2_or2_1 _2371_ (.X(_0467_),
    .B(_0107_),
    .A(net732));
 sg13g2_o21ai_1 _2372_ (.B1(_0467_),
    .Y(_0468_),
    .A1(_0106_),
    .A2(_1399_));
 sg13g2_o21ai_1 _2373_ (.B1(_1229_),
    .Y(_0469_),
    .A1(net732),
    .A2(net683));
 sg13g2_or2_1 _2374_ (.X(_0470_),
    .B(_0103_),
    .A(net732));
 sg13g2_a21oi_1 _2375_ (.A1(_0469_),
    .A2(_0470_),
    .Y(_0471_),
    .B1(net651));
 sg13g2_a21oi_2 _2376_ (.B1(_0471_),
    .Y(_0472_),
    .A2(_0468_),
    .A1(net652));
 sg13g2_mux4_1 _2377_ (.S0(net650),
    .A0(_0462_),
    .A1(_0465_),
    .A2(_0466_),
    .A3(_0472_),
    .S1(_1411_),
    .X(_0473_));
 sg13g2_a21oi_1 _2378_ (.A1(\crp.datapath.aluSrc1SelMux.d1[5] ),
    .A2(net624),
    .Y(_0474_),
    .B1(net622));
 sg13g2_a221oi_1 _2379_ (.B2(net626),
    .C1(_0474_),
    .B1(_0473_),
    .A1(_0101_),
    .Y(_0475_),
    .A2(net610));
 sg13g2_mux2_1 _2380_ (.A0(net583),
    .A1(_0460_),
    .S(net586),
    .X(_0476_));
 sg13g2_nor2_1 _2381_ (.A(net589),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_a21o_1 _2382_ (.A2(_0441_),
    .A1(net589),
    .B1(_0477_),
    .X(_0478_));
 sg13g2_nor2b_1 _2383_ (.A(_0478_),
    .B_N(_0405_),
    .Y(_0479_));
 sg13g2_nand2b_2 _2384_ (.Y(_0480_),
    .B(_1435_),
    .A_N(net588));
 sg13g2_and2_1 _2385_ (.A(_1506_),
    .B(_1515_),
    .X(_0481_));
 sg13g2_nand2_2 _2386_ (.Y(_0482_),
    .A(net621),
    .B(_0481_));
 sg13g2_inv_1 _2387_ (.Y(_0483_),
    .A(_0482_));
 sg13g2_nor3_1 _2388_ (.A(_1516_),
    .B(_0399_),
    .C(_0481_),
    .Y(_0484_));
 sg13g2_o21ai_1 _2389_ (.B1(_0484_),
    .Y(_0485_),
    .A1(_1506_),
    .A2(_0480_));
 sg13g2_o21ai_1 _2390_ (.B1(_0485_),
    .Y(_0486_),
    .A1(_0480_),
    .A2(_0482_));
 sg13g2_nor3_2 _2391_ (.A(_0404_),
    .B(_0479_),
    .C(_0486_),
    .Y(_0487_));
 sg13g2_a21o_2 _2392_ (.A2(_0487_),
    .A1(net613),
    .B1(_1436_),
    .X(_0488_));
 sg13g2_o21ai_1 _2393_ (.B1(net632),
    .Y(_0489_),
    .A1(\crp.datapath.aluSrc1SelMux.d1[0] ),
    .A2(net665));
 sg13g2_a21oi_1 _2394_ (.A1(_1357_),
    .A2(_0488_),
    .Y(_0490_),
    .B1(_0489_));
 sg13g2_a21o_1 _2395_ (.A2(net630),
    .A1(\crp.datapath.aluSrc1SelMux.d0[0] ),
    .B1(_0490_),
    .X(_0491_));
 sg13g2_nor2_1 _2396_ (.A(net686),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_mux2_1 _2397_ (.A0(_0079_),
    .A1(_0078_),
    .S(net640),
    .X(_0493_));
 sg13g2_a21oi_1 _2398_ (.A1(net708),
    .A2(_1222_),
    .Y(_0494_),
    .B1(net645));
 sg13g2_o21ai_1 _2399_ (.B1(_0494_),
    .Y(_0495_),
    .A1(_0076_),
    .A2(net639));
 sg13g2_a21oi_1 _2400_ (.A1(net644),
    .A2(_0493_),
    .Y(_0496_),
    .B1(net637));
 sg13g2_mux4_1 _2401_ (.S0(net641),
    .A0(_0081_),
    .A1(_0080_),
    .A2(_0083_),
    .A3(_0082_),
    .S1(net645),
    .X(_0497_));
 sg13g2_o21ai_1 _2402_ (.B1(_1452_),
    .Y(_0498_),
    .A1(_1447_),
    .A2(_0497_));
 sg13g2_a21oi_1 _2403_ (.A1(_0495_),
    .A2(_0496_),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_mux2_1 _2404_ (.A0(_0071_),
    .A1(_0070_),
    .S(net640),
    .X(_0500_));
 sg13g2_a21oi_1 _2405_ (.A1(net706),
    .A2(_1220_),
    .Y(_0501_),
    .B1(net642));
 sg13g2_o21ai_1 _2406_ (.B1(_0501_),
    .Y(_0502_),
    .A1(_0068_),
    .A2(net638));
 sg13g2_a21oi_1 _2407_ (.A1(net643),
    .A2(_0500_),
    .Y(_0503_),
    .B1(net634));
 sg13g2_mux2_1 _2408_ (.A0(_0075_),
    .A1(_0074_),
    .S(net640),
    .X(_0504_));
 sg13g2_a21oi_1 _2409_ (.A1(net706),
    .A2(_1221_),
    .Y(_0505_),
    .B1(net643));
 sg13g2_o21ai_1 _2410_ (.B1(_0505_),
    .Y(_0506_),
    .A1(_0072_),
    .A2(net638));
 sg13g2_a21oi_1 _2411_ (.A1(net643),
    .A2(_0504_),
    .Y(_0507_),
    .B1(_1447_));
 sg13g2_a221oi_1 _2412_ (.B2(_0507_),
    .C1(net633),
    .B1(_0506_),
    .A1(_0502_),
    .Y(_0508_),
    .A2(_0503_));
 sg13g2_nor2_2 _2413_ (.A(_0499_),
    .B(_0508_),
    .Y(_0509_));
 sg13g2_and2_1 _2414_ (.A(_1442_),
    .B(_0509_),
    .X(_0510_));
 sg13g2_a22oi_1 _2415_ (.Y(_0511_),
    .B1(_1439_),
    .B2(net725),
    .A2(_1277_),
    .A1(net723));
 sg13g2_nor2b_1 _2416_ (.A(_0510_),
    .B_N(_0511_),
    .Y(_0512_));
 sg13g2_nand2b_2 _2417_ (.Y(_0513_),
    .B(_0511_),
    .A_N(_0510_));
 sg13g2_nor3_2 _2418_ (.A(net578),
    .B(_1547_),
    .C(_1576_),
    .Y(_0514_));
 sg13g2_a21oi_2 _2419_ (.B1(_1471_),
    .Y(_0515_),
    .A2(_1577_),
    .A1(_1548_));
 sg13g2_o21ai_1 _2420_ (.B1(net578),
    .Y(_0516_),
    .A1(_1547_),
    .A2(_1576_));
 sg13g2_nor2_2 _2421_ (.A(_0514_),
    .B(_0515_),
    .Y(_0517_));
 sg13g2_nand2_1 _2422_ (.Y(_0518_),
    .A(net592),
    .B(net585));
 sg13g2_xor2_1 _2423_ (.B(net585),
    .A(net592),
    .X(_0519_));
 sg13g2_xnor2_1 _2424_ (.Y(_0520_),
    .A(net592),
    .B(net585));
 sg13g2_nor2_2 _2425_ (.A(_1435_),
    .B(net588),
    .Y(_0521_));
 sg13g2_nand2b_1 _2426_ (.Y(_0522_),
    .B(net585),
    .A_N(net592));
 sg13g2_o21ai_1 _2427_ (.B1(_0522_),
    .Y(_0523_),
    .A1(_0519_),
    .A2(_0521_));
 sg13g2_o21ai_1 _2428_ (.B1(_0523_),
    .Y(_0524_),
    .A1(_0514_),
    .A2(_0515_));
 sg13g2_nand2_1 _2429_ (.Y(_0525_),
    .A(net578),
    .B(_1578_));
 sg13g2_a22oi_1 _2430_ (.Y(_0526_),
    .B1(net573),
    .B2(_0512_),
    .A2(_1578_),
    .A1(net578));
 sg13g2_a22oi_1 _2431_ (.Y(_0527_),
    .B1(_0524_),
    .B2(_0526_),
    .A2(_0513_),
    .A1(_0368_));
 sg13g2_a21oi_1 _2432_ (.A1(net718),
    .A2(net673),
    .Y(_0528_),
    .B1(_0113_));
 sg13g2_a221oi_1 _2433_ (.B2(_1233_),
    .C1(_0528_),
    .B1(net641),
    .A1(_0030_),
    .Y(_0529_),
    .A2(net673));
 sg13g2_a221oi_1 _2434_ (.B2(_1396_),
    .C1(net705),
    .B1(net696),
    .A1(net717),
    .Y(_0530_),
    .A2(_1232_));
 sg13g2_o21ai_1 _2435_ (.B1(_0530_),
    .Y(_0531_),
    .A1(_0111_),
    .A2(net641));
 sg13g2_nand3b_1 _2436_ (.B(_0531_),
    .C(_1447_),
    .Y(_0532_),
    .A_N(_0529_));
 sg13g2_mux4_1 _2437_ (.S0(net641),
    .A0(_1234_),
    .A1(_1235_),
    .A2(_1236_),
    .A3(_1237_),
    .S1(net646),
    .X(_0533_));
 sg13g2_a21oi_1 _2438_ (.A1(net636),
    .A2(_0533_),
    .Y(_0534_),
    .B1(_1451_));
 sg13g2_mux2_1 _2439_ (.A0(_0109_),
    .A1(_0108_),
    .S(net640),
    .X(_0535_));
 sg13g2_nor3_1 _2440_ (.A(net707),
    .B(_0106_),
    .C(net681),
    .Y(_0536_));
 sg13g2_or2_1 _2441_ (.X(_0537_),
    .B(_0107_),
    .A(net714));
 sg13g2_nand3_1 _2442_ (.B(net671),
    .C(_0537_),
    .A(_0030_),
    .Y(_0538_));
 sg13g2_o21ai_1 _2443_ (.B1(net635),
    .Y(_0539_),
    .A1(_0536_),
    .A2(_0538_));
 sg13g2_a21o_1 _2444_ (.A2(_0535_),
    .A1(net644),
    .B1(_0539_),
    .X(_0540_));
 sg13g2_and3_1 _2445_ (.X(_0541_),
    .A(net713),
    .B(_0104_),
    .C(net671));
 sg13g2_a21oi_1 _2446_ (.A1(net714),
    .A2(net671),
    .Y(_0542_),
    .B1(_1230_));
 sg13g2_o21ai_1 _2447_ (.B1(net644),
    .Y(_0543_),
    .A1(_0541_),
    .A2(_0542_));
 sg13g2_nand3_1 _2448_ (.B(_1229_),
    .C(net671),
    .A(net716),
    .Y(_0544_));
 sg13g2_nor2_1 _2449_ (.A(net716),
    .B(_0103_),
    .Y(_0545_));
 sg13g2_nor3_1 _2450_ (.A(net704),
    .B(net683),
    .C(_0545_),
    .Y(_0546_));
 sg13g2_a21oi_1 _2451_ (.A1(_0544_),
    .A2(_0546_),
    .Y(_0547_),
    .B1(net634));
 sg13g2_a21oi_2 _2452_ (.B1(_1452_),
    .Y(_0548_),
    .A2(_0547_),
    .A1(_0543_));
 sg13g2_a22oi_1 _2453_ (.Y(_0549_),
    .B1(_0540_),
    .B2(_0548_),
    .A2(_0534_),
    .A1(_0532_));
 sg13g2_nand2_1 _2454_ (.Y(_0550_),
    .A(\crp.datapath.aluSrc2SelMux.d2[5] ),
    .B(_1277_));
 sg13g2_o21ai_1 _2455_ (.B1(_0550_),
    .Y(_0551_),
    .A1(net720),
    .A2(net647));
 sg13g2_a21oi_1 _2456_ (.A1(_1442_),
    .A2(_0549_),
    .Y(_0552_),
    .B1(_0551_));
 sg13g2_a21o_2 _2457_ (.A2(_0549_),
    .A1(_1442_),
    .B1(_0551_),
    .X(_0553_));
 sg13g2_nand2_1 _2458_ (.Y(_0554_),
    .A(net583),
    .B(_0553_));
 sg13g2_nor2_1 _2459_ (.A(net583),
    .B(_0553_),
    .Y(_0555_));
 sg13g2_xnor2_1 _2460_ (.Y(_0556_),
    .A(net583),
    .B(_0553_));
 sg13g2_and3_1 _2461_ (.X(_0557_),
    .A(net713),
    .B(_0087_),
    .C(net668));
 sg13g2_a21oi_1 _2462_ (.A1(net715),
    .A2(net668),
    .Y(_0558_),
    .B1(_1223_));
 sg13g2_o21ai_1 _2463_ (.B1(net642),
    .Y(_0559_),
    .A1(_0557_),
    .A2(_0558_));
 sg13g2_a21o_1 _2464_ (.A2(net668),
    .A1(net715),
    .B1(_0086_),
    .X(_0560_));
 sg13g2_nor2_1 _2465_ (.A(net706),
    .B(_0085_),
    .Y(_0561_));
 sg13g2_nor3_1 _2466_ (.A(net704),
    .B(net679),
    .C(_0561_),
    .Y(_0562_));
 sg13g2_and3_1 _2467_ (.X(_0563_),
    .A(net717),
    .B(_0095_),
    .C(net673));
 sg13g2_a21oi_1 _2468_ (.A1(net717),
    .A2(net673),
    .Y(_0564_),
    .B1(_1227_));
 sg13g2_o21ai_1 _2469_ (.B1(net646),
    .Y(_0565_),
    .A1(_0563_),
    .A2(_0564_));
 sg13g2_nand3b_1 _2470_ (.B(net673),
    .C(net717),
    .Y(_0566_),
    .A_N(_0093_));
 sg13g2_a221oi_1 _2471_ (.B2(_1396_),
    .C1(net705),
    .B1(net696),
    .A1(net708),
    .Y(_0567_),
    .A2(_1226_));
 sg13g2_mux4_1 _2472_ (.S0(net640),
    .A0(_0090_),
    .A1(_0089_),
    .A2(_0092_),
    .A3(_0091_),
    .S1(net643),
    .X(_0568_));
 sg13g2_nand2b_2 _2473_ (.Y(_0569_),
    .B(net634),
    .A_N(_0568_));
 sg13g2_a21oi_1 _2474_ (.A1(_0560_),
    .A2(_0562_),
    .Y(_0570_),
    .B1(net634));
 sg13g2_a21oi_2 _2475_ (.B1(net633),
    .Y(_0571_),
    .A2(_0570_),
    .A1(_0559_));
 sg13g2_mux4_1 _2476_ (.S0(net641),
    .A0(_0098_),
    .A1(_0097_),
    .A2(_0100_),
    .A3(_0099_),
    .S1(net646),
    .X(_0572_));
 sg13g2_nand2b_1 _2477_ (.Y(_0573_),
    .B(net636),
    .A_N(_0572_));
 sg13g2_a21oi_1 _2478_ (.A1(_0566_),
    .A2(_0567_),
    .Y(_0574_),
    .B1(net636));
 sg13g2_a21oi_1 _2479_ (.A1(_0565_),
    .A2(_0574_),
    .Y(_0575_),
    .B1(_1451_));
 sg13g2_a22oi_1 _2480_ (.Y(_0576_),
    .B1(_0573_),
    .B2(_0575_),
    .A2(_0571_),
    .A1(_0569_));
 sg13g2_nor2_1 _2481_ (.A(_1156_),
    .B(_1276_),
    .Y(_0577_));
 sg13g2_a221oi_1 _2482_ (.B2(_0576_),
    .C1(_0577_),
    .B1(_1442_),
    .A1(net723),
    .Y(_0578_),
    .A2(_1439_));
 sg13g2_nand2b_2 _2483_ (.Y(_0579_),
    .B(_0460_),
    .A_N(_0578_));
 sg13g2_nand2b_1 _2484_ (.Y(_0580_),
    .B(_0578_),
    .A_N(_0460_));
 sg13g2_nand2_2 _2485_ (.Y(_0581_),
    .A(_0580_),
    .B(_0579_));
 sg13g2_nand2_2 _2486_ (.Y(_0582_),
    .A(_0556_),
    .B(_0581_));
 sg13g2_a221oi_1 _2487_ (.B2(_0526_),
    .C1(_0582_),
    .B1(_0524_),
    .A1(_0368_),
    .Y(_0583_),
    .A2(_0513_));
 sg13g2_and3_1 _2488_ (.X(_0584_),
    .A(net713),
    .B(_0138_),
    .C(net670));
 sg13g2_a21oi_1 _2489_ (.A1(net713),
    .A2(net670),
    .Y(_0585_),
    .B1(_1247_));
 sg13g2_o21ai_1 _2490_ (.B1(net643),
    .Y(_0586_),
    .A1(_0584_),
    .A2(_0585_));
 sg13g2_nand3_1 _2491_ (.B(_1246_),
    .C(net669),
    .A(net713),
    .Y(_0587_));
 sg13g2_a221oi_1 _2492_ (.B2(_1396_),
    .C1(net704),
    .B1(net697),
    .A1(net707),
    .Y(_0588_),
    .A2(_1245_));
 sg13g2_and3_1 _2493_ (.X(_0589_),
    .A(net717),
    .B(_0146_),
    .C(net674));
 sg13g2_a21oi_1 _2494_ (.A1(net717),
    .A2(net674),
    .Y(_0590_),
    .B1(_1250_));
 sg13g2_o21ai_1 _2495_ (.B1(net646),
    .Y(_0591_),
    .A1(_0589_),
    .A2(_0590_));
 sg13g2_nand3_1 _2496_ (.B(_1249_),
    .C(net673),
    .A(net717),
    .Y(_0592_));
 sg13g2_a221oi_1 _2497_ (.B2(_1396_),
    .C1(net705),
    .B1(net696),
    .A1(net708),
    .Y(_0593_),
    .A2(_1248_));
 sg13g2_mux4_1 _2498_ (.S0(net640),
    .A0(_0141_),
    .A1(_0140_),
    .A2(_0143_),
    .A3(_0142_),
    .S1(net643),
    .X(_0594_));
 sg13g2_nand2b_1 _2499_ (.Y(_0595_),
    .B(net635),
    .A_N(_0594_));
 sg13g2_a21oi_1 _2500_ (.A1(_0587_),
    .A2(_0588_),
    .Y(_0596_),
    .B1(net635));
 sg13g2_a21oi_1 _2501_ (.A1(_0586_),
    .A2(_0596_),
    .Y(_0597_),
    .B1(net633));
 sg13g2_mux4_1 _2502_ (.S0(net641),
    .A0(_0149_),
    .A1(_0148_),
    .A2(_0151_),
    .A3(_0150_),
    .S1(net646),
    .X(_0598_));
 sg13g2_nand2b_1 _2503_ (.Y(_0599_),
    .B(net636),
    .A_N(_0598_));
 sg13g2_a21oi_1 _2504_ (.A1(_0592_),
    .A2(_0593_),
    .Y(_0600_),
    .B1(net636));
 sg13g2_a21oi_2 _2505_ (.B1(_1451_),
    .Y(_0601_),
    .A2(_0600_),
    .A1(_0591_));
 sg13g2_a22oi_1 _2506_ (.Y(_0602_),
    .B1(_0599_),
    .B2(_0601_),
    .A2(_0597_),
    .A1(_0595_));
 sg13g2_nor2_1 _2507_ (.A(_0031_),
    .B(net647),
    .Y(_0603_));
 sg13g2_a221oi_1 _2508_ (.B2(_0602_),
    .C1(_0603_),
    .B1(_1442_),
    .A1(\crp.datapath.aluSrc2SelMux.d2[7] ),
    .Y(_0604_),
    .A2(_1277_));
 sg13g2_or2_1 _2509_ (.X(_0605_),
    .B(_0604_),
    .A(_0440_));
 sg13g2_nand2_1 _2510_ (.Y(_0606_),
    .A(_0440_),
    .B(_0604_));
 sg13g2_and3_1 _2511_ (.X(_0607_),
    .A(net713),
    .B(_0121_),
    .C(net668));
 sg13g2_a21oi_1 _2512_ (.A1(net715),
    .A2(net668),
    .Y(_0608_),
    .B1(_1238_));
 sg13g2_o21ai_1 _2513_ (.B1(net642),
    .Y(_0609_),
    .A1(_0607_),
    .A2(_0608_));
 sg13g2_a21o_1 _2514_ (.A2(net668),
    .A1(net715),
    .B1(_0120_),
    .X(_0610_));
 sg13g2_nor2_1 _2515_ (.A(net706),
    .B(_0119_),
    .Y(_0611_));
 sg13g2_nor3_1 _2516_ (.A(net704),
    .B(net679),
    .C(_0611_),
    .Y(_0612_));
 sg13g2_and3_1 _2517_ (.X(_0613_),
    .A(net719),
    .B(_0129_),
    .C(net677));
 sg13g2_a21oi_1 _2518_ (.A1(net719),
    .A2(net677),
    .Y(_0614_),
    .B1(_1240_));
 sg13g2_o21ai_1 _2519_ (.B1(net645),
    .Y(_0615_),
    .A1(_0613_),
    .A2(_0614_));
 sg13g2_nand3b_1 _2520_ (.B(net677),
    .C(net719),
    .Y(_0616_),
    .A_N(_0127_));
 sg13g2_a221oi_1 _2521_ (.B2(_1396_),
    .C1(net705),
    .B1(net696),
    .A1(net708),
    .Y(_0617_),
    .A2(_1239_));
 sg13g2_mux4_1 _2522_ (.S0(net640),
    .A0(_0124_),
    .A1(_0123_),
    .A2(_0126_),
    .A3(_0125_),
    .S1(net643),
    .X(_0618_));
 sg13g2_nand2b_1 _2523_ (.Y(_0619_),
    .B(net634),
    .A_N(_0618_));
 sg13g2_a21oi_1 _2524_ (.A1(_0610_),
    .A2(_0612_),
    .Y(_0620_),
    .B1(net634));
 sg13g2_a21oi_1 _2525_ (.A1(_0609_),
    .A2(_0620_),
    .Y(_0621_),
    .B1(net633));
 sg13g2_mux4_1 _2526_ (.S0(net641),
    .A0(_1241_),
    .A1(_1242_),
    .A2(_1243_),
    .A3(_1244_),
    .S1(net645),
    .X(_0622_));
 sg13g2_a21oi_1 _2527_ (.A1(_0616_),
    .A2(_0617_),
    .Y(_0623_),
    .B1(net636));
 sg13g2_a22oi_1 _2528_ (.Y(_0624_),
    .B1(_0623_),
    .B2(_0615_),
    .A2(_0622_),
    .A1(net637));
 sg13g2_a22oi_1 _2529_ (.Y(_0625_),
    .B1(_0624_),
    .B2(net633),
    .A2(_0621_),
    .A1(_0619_));
 sg13g2_nor2_1 _2530_ (.A(_1154_),
    .B(_1276_),
    .Y(_0626_));
 sg13g2_a221oi_1 _2531_ (.B2(_0625_),
    .C1(_0626_),
    .B1(_1442_),
    .A1(net704),
    .Y(_0627_),
    .A2(_1439_));
 sg13g2_nand2_1 _2532_ (.Y(_0628_),
    .A(_0424_),
    .B(_0627_));
 sg13g2_nand2_1 _2533_ (.Y(_0629_),
    .A(_0606_),
    .B(_0628_));
 sg13g2_nand2_1 _2534_ (.Y(_0630_),
    .A(_0605_),
    .B(_0629_));
 sg13g2_nand2_1 _2535_ (.Y(_0631_),
    .A(_0460_),
    .B(_0578_));
 sg13g2_nor2b_1 _2536_ (.A(_0631_),
    .B_N(_0556_),
    .Y(_0632_));
 sg13g2_a21oi_1 _2537_ (.A1(_0475_),
    .A2(_0552_),
    .Y(_0633_),
    .B1(_0632_));
 sg13g2_inv_1 _2538_ (.Y(_0634_),
    .A(_0633_));
 sg13g2_nand2_1 _2539_ (.Y(_0635_),
    .A(_0630_),
    .B(_0633_));
 sg13g2_nand2b_2 _2540_ (.Y(_0636_),
    .B(_0424_),
    .A_N(_0627_));
 sg13g2_nand2b_1 _2541_ (.Y(_0637_),
    .B(_0627_),
    .A_N(_0424_));
 sg13g2_and2_2 _2542_ (.A(_0636_),
    .B(_0637_),
    .X(_0638_));
 sg13g2_inv_1 _2543_ (.Y(_0639_),
    .A(_0638_));
 sg13g2_nand2b_1 _2544_ (.Y(_0640_),
    .B(net584),
    .A_N(_0604_));
 sg13g2_inv_1 _2545_ (.Y(_0641_),
    .A(_0640_));
 sg13g2_nand2b_1 _2546_ (.Y(_0642_),
    .B(_0604_),
    .A_N(net584));
 sg13g2_nand2_2 _2547_ (.Y(_0643_),
    .A(_0605_),
    .B(_0606_));
 sg13g2_o21ai_1 _2548_ (.B1(_0630_),
    .Y(_0644_),
    .A1(_0638_),
    .A2(_0643_));
 sg13g2_o21ai_1 _2549_ (.B1(_0644_),
    .Y(_0645_),
    .A1(_0635_),
    .A2(_0583_));
 sg13g2_nor2_2 _2550_ (.A(_0032_),
    .B(net647),
    .Y(_0646_));
 sg13g2_a22oi_1 _2551_ (.Y(_0647_),
    .B1(_1392_),
    .B2(\crp.datapath.aluSrc1SelMux.d1[8] ),
    .A2(net609),
    .A1(_1253_));
 sg13g2_nand2b_1 _2552_ (.Y(_0648_),
    .B(_0646_),
    .A_N(_0647_));
 sg13g2_nor2_1 _2553_ (.A(_0646_),
    .B(_0647_),
    .Y(_0649_));
 sg13g2_xnor2_1 _2554_ (.Y(_0650_),
    .A(_0646_),
    .B(_0647_));
 sg13g2_xor2_1 _2555_ (.B(_0647_),
    .A(_0646_),
    .X(_0651_));
 sg13g2_nor2b_2 _2556_ (.A(_1515_),
    .B_N(net621),
    .Y(_0652_));
 sg13g2_and2_2 _2557_ (.A(_1505_),
    .B(_0652_),
    .X(_0653_));
 sg13g2_nand2_2 _2558_ (.Y(_0654_),
    .A(_1505_),
    .B(_0652_));
 sg13g2_xnor2_1 _2559_ (.Y(_0655_),
    .A(_0651_),
    .B(_0645_));
 sg13g2_nand2_1 _2560_ (.Y(_0656_),
    .A(net572),
    .B(_0513_));
 sg13g2_o21ai_1 _2561_ (.B1(_0518_),
    .Y(_0657_),
    .A1(_0520_),
    .A2(_0480_));
 sg13g2_a21oi_2 _2562_ (.B1(_0514_),
    .Y(_0658_),
    .A2(_0516_),
    .A1(_0657_));
 sg13g2_nor2_1 _2563_ (.A(net572),
    .B(_0513_),
    .Y(_0659_));
 sg13g2_xnor2_1 _2564_ (.Y(_0660_),
    .A(net573),
    .B(_0512_));
 sg13g2_o21ai_1 _2565_ (.B1(_0656_),
    .Y(_0661_),
    .A1(_0659_),
    .A2(_0658_));
 sg13g2_nor2_1 _2566_ (.A(_0556_),
    .B(_0581_),
    .Y(_0662_));
 sg13g2_o21ai_1 _2567_ (.B1(_0554_),
    .Y(_0663_),
    .A1(_0555_),
    .A2(_0579_));
 sg13g2_nand2b_1 _2568_ (.Y(_0664_),
    .B(_0642_),
    .A_N(_0636_));
 sg13g2_nand3_1 _2569_ (.B(_0643_),
    .C(_0663_),
    .A(_0638_),
    .Y(_0665_));
 sg13g2_nand3_1 _2570_ (.B(_0664_),
    .C(_0665_),
    .A(_0640_),
    .Y(_0666_));
 sg13g2_and3_1 _2571_ (.X(_0667_),
    .A(_0638_),
    .B(_0643_),
    .C(_0662_));
 sg13g2_a21oi_2 _2572_ (.B1(_0666_),
    .Y(_0668_),
    .A2(_0661_),
    .A1(_0667_));
 sg13g2_or2_1 _2573_ (.X(_0669_),
    .B(_0668_),
    .A(_0651_));
 sg13g2_and2_2 _2574_ (.A(_1505_),
    .B(_1515_),
    .X(_0670_));
 sg13g2_and2_1 _2575_ (.A(net621),
    .B(_0670_),
    .X(_0671_));
 sg13g2_nand2_2 _2576_ (.Y(_0672_),
    .A(net621),
    .B(_0670_));
 sg13g2_a21oi_1 _2577_ (.A1(_0651_),
    .A2(_0668_),
    .Y(_0673_),
    .B1(net601));
 sg13g2_a22oi_1 _2578_ (.Y(_0674_),
    .B1(_0669_),
    .B2(_0673_),
    .A2(_0655_),
    .A1(_0653_));
 sg13g2_nand2_2 _2579_ (.Y(_0675_),
    .A(_0674_),
    .B(net612));
 sg13g2_and2_2 _2580_ (.A(_1542_),
    .B(_0675_),
    .X(_0676_));
 sg13g2_inv_4 _2581_ (.A(_0676_),
    .Y(_0677_));
 sg13g2_o21ai_1 _2582_ (.B1(net632),
    .Y(_0678_),
    .A1(\crp.datapath.aluSrc1SelMux.d1[8] ),
    .A2(net665));
 sg13g2_a21oi_2 _2583_ (.B1(_0678_),
    .Y(_0679_),
    .A2(_0677_),
    .A1(_1357_));
 sg13g2_a21oi_2 _2584_ (.B1(_0679_),
    .Y(_0680_),
    .A2(net630),
    .A1(\crp.datapath.aluSrc1SelMux.d0[8] ));
 sg13g2_a21oi_2 _2585_ (.B1(_0492_),
    .Y(uo_out[0]),
    .A2(net686),
    .A1(_0680_));
 sg13g2_xnor2_1 _2586_ (.Y(_0681_),
    .A(_0480_),
    .B(_0520_));
 sg13g2_nand2_1 _2587_ (.Y(_0682_),
    .A(net602),
    .B(_0681_));
 sg13g2_nor2b_1 _2588_ (.A(net586),
    .B_N(_0460_),
    .Y(_0683_));
 sg13g2_a21o_1 _2589_ (.A2(net572),
    .A1(net587),
    .B1(_0683_),
    .X(_0684_));
 sg13g2_nor2_1 _2590_ (.A(net587),
    .B(_1578_),
    .Y(_0685_));
 sg13g2_nor2b_1 _2591_ (.A(net585),
    .B_N(net588),
    .Y(_0686_));
 sg13g2_nor3_1 _2592_ (.A(net590),
    .B(_0685_),
    .C(_0686_),
    .Y(_0687_));
 sg13g2_a21oi_1 _2593_ (.A1(net591),
    .A2(_0684_),
    .Y(_0688_),
    .B1(_0687_));
 sg13g2_or2_1 _2594_ (.X(_0689_),
    .B(_0688_),
    .A(_1546_));
 sg13g2_or4_1 _2595_ (.A(net591),
    .B(_1517_),
    .C(_0521_),
    .D(_0686_),
    .X(_0690_));
 sg13g2_and2_1 _2596_ (.A(net577),
    .B(_0690_),
    .X(_0691_));
 sg13g2_nor2b_1 _2597_ (.A(net586),
    .B_N(_0424_),
    .Y(_0692_));
 sg13g2_and2_1 _2598_ (.A(net586),
    .B(net583),
    .X(_0693_));
 sg13g2_o21ai_1 _2599_ (.B1(_1499_),
    .Y(_0694_),
    .A1(_0692_),
    .A2(_0693_));
 sg13g2_nand2_1 _2600_ (.Y(_0695_),
    .A(net587),
    .B(net584));
 sg13g2_o21ai_1 _2601_ (.B1(_0694_),
    .Y(_0696_),
    .A1(_1499_),
    .A2(_0695_));
 sg13g2_nand2b_1 _2602_ (.Y(_0697_),
    .B(_0481_),
    .A_N(net621));
 sg13g2_nand2b_1 _2603_ (.Y(_0698_),
    .B(_0696_),
    .A_N(_0697_));
 sg13g2_nand2_1 _2604_ (.Y(_0699_),
    .A(net589),
    .B(net584));
 sg13g2_nand2_1 _2605_ (.Y(_0700_),
    .A(_0694_),
    .B(_0699_));
 sg13g2_nor3_2 _2606_ (.A(_1505_),
    .B(net621),
    .C(_1515_),
    .Y(_0701_));
 sg13g2_a21oi_1 _2607_ (.A1(_0700_),
    .A2(_0701_),
    .Y(_0702_),
    .B1(net577));
 sg13g2_a22oi_1 _2608_ (.Y(_0703_),
    .B1(_0698_),
    .B2(_0702_),
    .A2(_0691_),
    .A1(_0689_));
 sg13g2_xnor2_1 _2609_ (.Y(_0704_),
    .A(_0520_),
    .B(_0521_));
 sg13g2_or2_1 _2610_ (.X(_0705_),
    .B(_0518_),
    .A(_0482_));
 sg13g2_and2_2 _2611_ (.A(_1506_),
    .B(_0652_),
    .X(_0706_));
 sg13g2_o21ai_1 _2612_ (.B1(_0706_),
    .Y(_0707_),
    .A1(net592),
    .A2(net585));
 sg13g2_a22oi_1 _2613_ (.Y(_0708_),
    .B1(_0704_),
    .B2(_0653_),
    .A2(_0670_),
    .A1(_0519_));
 sg13g2_nand4_1 _2614_ (.B(_0705_),
    .C(_0707_),
    .A(net601),
    .Y(_0709_),
    .D(_0708_));
 sg13g2_o21ai_1 _2615_ (.B1(_0682_),
    .Y(_0710_),
    .A1(_0703_),
    .A2(_0709_));
 sg13g2_nand2_1 _2616_ (.Y(_0711_),
    .A(net612),
    .B(_0710_));
 sg13g2_o21ai_1 _2617_ (.B1(_0711_),
    .Y(_0712_),
    .A1(net611),
    .A2(_0397_));
 sg13g2_o21ai_1 _2618_ (.B1(net632),
    .Y(_0713_),
    .A1(\crp.datapath.aluSrc1SelMux.d1[1] ),
    .A2(_1355_));
 sg13g2_a21oi_1 _2619_ (.A1(_1357_),
    .A2(_0712_),
    .Y(_0714_),
    .B1(_0713_));
 sg13g2_a21oi_2 _2620_ (.B1(_0714_),
    .Y(_0715_),
    .A2(net630),
    .A1(\crp.datapath.aluSrc1SelMux.d0[1] ));
 sg13g2_nor2_1 _2621_ (.A(net734),
    .B(net647),
    .Y(_0716_));
 sg13g2_a22oi_1 _2622_ (.Y(_0717_),
    .B1(_1392_),
    .B2(\crp.datapath.aluSrc1SelMux.d1[9] ),
    .A2(net609),
    .A1(_1254_));
 sg13g2_nand2b_1 _2623_ (.Y(_0718_),
    .B(_0717_),
    .A_N(_0716_));
 sg13g2_nand2b_1 _2624_ (.Y(_0719_),
    .B(_0716_),
    .A_N(_0717_));
 sg13g2_and2_1 _2625_ (.A(_0718_),
    .B(_0719_),
    .X(_0720_));
 sg13g2_nand2_2 _2626_ (.Y(_0721_),
    .A(_0718_),
    .B(_0719_));
 sg13g2_o21ai_1 _2627_ (.B1(_0648_),
    .Y(_0722_),
    .A1(_0651_),
    .A2(_0668_));
 sg13g2_a21oi_1 _2628_ (.A1(_0720_),
    .A2(_0722_),
    .Y(_0723_),
    .B1(_0672_));
 sg13g2_o21ai_1 _2629_ (.B1(_0723_),
    .Y(_0724_),
    .A1(_0720_),
    .A2(_0722_));
 sg13g2_nor2_1 _2630_ (.A(_0649_),
    .B(_0721_),
    .Y(_0725_));
 sg13g2_o21ai_1 _2631_ (.B1(_0725_),
    .Y(_0726_),
    .A1(_0645_),
    .A2(_0650_));
 sg13g2_nand2_1 _2632_ (.Y(_0727_),
    .A(_0651_),
    .B(_0721_));
 sg13g2_a21oi_1 _2633_ (.A1(_0649_),
    .A2(_0721_),
    .Y(_0728_),
    .B1(_0654_));
 sg13g2_o21ai_1 _2634_ (.B1(_0728_),
    .Y(_0729_),
    .A1(_0727_),
    .A2(_0645_));
 sg13g2_nor2b_1 _2635_ (.A(_0729_),
    .B_N(_0726_),
    .Y(_0730_));
 sg13g2_nor2_2 _2636_ (.A(_1375_),
    .B(_0730_),
    .Y(_0731_));
 sg13g2_a22oi_1 _2637_ (.Y(_0732_),
    .B1(_0724_),
    .B2(_0731_),
    .A2(_1496_),
    .A1(_1375_));
 sg13g2_nor2_1 _2638_ (.A(\crp.datapath.aluSrc1SelMux.d1[9] ),
    .B(net666),
    .Y(_0733_));
 sg13g2_nor2_1 _2639_ (.A(net628),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_o21ai_1 _2640_ (.B1(_0734_),
    .Y(_0735_),
    .A1(_0732_),
    .A2(net627));
 sg13g2_o21ai_1 _2641_ (.B1(_0735_),
    .Y(_0736_),
    .A1(_1184_),
    .A2(net631));
 sg13g2_nand2_1 _2642_ (.Y(_0737_),
    .A(_0736_),
    .B(net686));
 sg13g2_o21ai_1 _2643_ (.B1(_0737_),
    .Y(uo_out[1]),
    .A1(net686),
    .A2(_0715_));
 sg13g2_o21ai_1 _2644_ (.B1(_1579_),
    .Y(_0738_),
    .A1(net588),
    .A2(net585));
 sg13g2_a21o_1 _2645_ (.A2(_1544_),
    .A1(net591),
    .B1(_1517_),
    .X(_0739_));
 sg13g2_a21oi_1 _2646_ (.A1(_1499_),
    .A2(_0738_),
    .Y(_0740_),
    .B1(_0739_));
 sg13g2_nor2_1 _2647_ (.A(net591),
    .B(_0369_),
    .Y(_0741_));
 sg13g2_nor2_1 _2648_ (.A(_1499_),
    .B(_0476_),
    .Y(_0742_));
 sg13g2_nor3_1 _2649_ (.A(_1546_),
    .B(_0741_),
    .C(_0742_),
    .Y(_0743_));
 sg13g2_o21ai_1 _2650_ (.B1(net578),
    .Y(_0744_),
    .A1(_0740_),
    .A2(_0743_));
 sg13g2_xnor2_1 _2651_ (.Y(_0745_),
    .A(_0517_),
    .B(_0523_));
 sg13g2_nor2b_2 _2652_ (.A(_1509_),
    .B_N(_0670_),
    .Y(_0746_));
 sg13g2_inv_1 _2653_ (.Y(_0747_),
    .A(_0746_));
 sg13g2_nor2_2 _2654_ (.A(net589),
    .B(_0441_),
    .Y(_0748_));
 sg13g2_nor2_1 _2655_ (.A(_1515_),
    .B(_0699_),
    .Y(_0749_));
 sg13g2_o21ai_1 _2656_ (.B1(_0405_),
    .Y(_0750_),
    .A1(_0748_),
    .A2(_0749_));
 sg13g2_nand2_1 _2657_ (.Y(_0751_),
    .A(_0517_),
    .B(_0746_));
 sg13g2_a221oi_1 _2658_ (.B2(_0706_),
    .C1(net602),
    .B1(_0516_),
    .A1(_0483_),
    .Y(_0752_),
    .A2(_0514_));
 sg13g2_nand3_1 _2659_ (.B(_0751_),
    .C(_0752_),
    .A(_0750_),
    .Y(_0753_));
 sg13g2_a21oi_1 _2660_ (.A1(_0653_),
    .A2(_0745_),
    .Y(_0754_),
    .B1(_0753_));
 sg13g2_xnor2_1 _2661_ (.Y(_0755_),
    .A(_0517_),
    .B(_0657_));
 sg13g2_a22oi_1 _2662_ (.Y(_0756_),
    .B1(_0755_),
    .B2(net602),
    .A2(_0754_),
    .A1(_0744_));
 sg13g2_mux2_2 _2663_ (.A0(_1578_),
    .A1(_0756_),
    .S(net612),
    .X(_0757_));
 sg13g2_nor2_1 _2664_ (.A(\crp.datapath.aluSrc1SelMux.d1[2] ),
    .B(net665),
    .Y(_0758_));
 sg13g2_nor2_1 _2665_ (.A(net630),
    .B(_0758_),
    .Y(_0759_));
 sg13g2_o21ai_1 _2666_ (.B1(_0759_),
    .Y(_0760_),
    .A1(_1356_),
    .A2(_0757_));
 sg13g2_o21ai_1 _2667_ (.B1(_0760_),
    .Y(_0761_),
    .A1(_1188_),
    .A2(net631));
 sg13g2_nor2_1 _2668_ (.A(net685),
    .B(_0761_),
    .Y(_0762_));
 sg13g2_nor2_1 _2669_ (.A(net611),
    .B(_1467_),
    .Y(_0763_));
 sg13g2_nor2_2 _2670_ (.A(_0012_),
    .B(net647),
    .Y(_0764_));
 sg13g2_a22oi_1 _2671_ (.Y(_0765_),
    .B1(_1392_),
    .B2(\crp.datapath.aluSrc1SelMux.d1[10] ),
    .A2(net609),
    .A1(_1255_));
 sg13g2_nor2_1 _2672_ (.A(_0764_),
    .B(_0765_),
    .Y(_0766_));
 sg13g2_xnor2_1 _2673_ (.Y(_0767_),
    .A(_0764_),
    .B(_0765_));
 sg13g2_inv_1 _2674_ (.Y(_0768_),
    .A(_0767_));
 sg13g2_nand2_1 _2675_ (.Y(_0769_),
    .A(_0650_),
    .B(_0720_));
 sg13g2_nand2_1 _2676_ (.Y(_0770_),
    .A(_0648_),
    .B(_0719_));
 sg13g2_nand2_1 _2677_ (.Y(_0771_),
    .A(_0718_),
    .B(_0770_));
 sg13g2_o21ai_1 _2678_ (.B1(_0771_),
    .Y(_0772_),
    .A1(_0668_),
    .A2(_0769_));
 sg13g2_nand2_1 _2679_ (.Y(_0773_),
    .A(_0767_),
    .B(_0772_));
 sg13g2_o21ai_1 _2680_ (.B1(_0671_),
    .Y(_0774_),
    .A1(_0767_),
    .A2(_0772_));
 sg13g2_nand2b_1 _2681_ (.Y(_0775_),
    .B(_0773_),
    .A_N(_0774_));
 sg13g2_nor2_1 _2682_ (.A(_0716_),
    .B(_0717_),
    .Y(_0776_));
 sg13g2_a21oi_1 _2683_ (.A1(_0649_),
    .A2(_0721_),
    .Y(_0777_),
    .B1(_0776_));
 sg13g2_o21ai_1 _2684_ (.B1(_0777_),
    .Y(_0778_),
    .A1(_0645_),
    .A2(_0727_));
 sg13g2_nand2b_1 _2685_ (.Y(_0779_),
    .B(_0767_),
    .A_N(_0778_));
 sg13g2_a21oi_1 _2686_ (.A1(_0768_),
    .A2(_0778_),
    .Y(_0780_),
    .B1(_0654_));
 sg13g2_a21oi_2 _2687_ (.B1(_1375_),
    .Y(_0781_),
    .A2(_0780_),
    .A1(_0779_));
 sg13g2_a21oi_2 _2688_ (.B1(_0763_),
    .Y(_0782_),
    .A2(_0775_),
    .A1(_0781_));
 sg13g2_or2_1 _2689_ (.X(_0783_),
    .B(net627),
    .A(_0782_));
 sg13g2_nor2_1 _2690_ (.A(\crp.datapath.aluSrc1SelMux.d1[10] ),
    .B(net666),
    .Y(_0784_));
 sg13g2_nor2_1 _2691_ (.A(net629),
    .B(_0784_),
    .Y(_0785_));
 sg13g2_a22oi_1 _2692_ (.Y(_0786_),
    .B1(_0783_),
    .B2(_0785_),
    .A2(net629),
    .A1(\crp.datapath.aluSrc1SelMux.d0[10] ));
 sg13g2_a21oi_2 _2693_ (.B1(_0762_),
    .Y(uo_out[2]),
    .A2(net685),
    .A1(_0786_));
 sg13g2_xnor2_1 _2694_ (.Y(_0787_),
    .A(_0658_),
    .B(_0660_));
 sg13g2_nor2_1 _2695_ (.A(net601),
    .B(_0787_),
    .Y(_0788_));
 sg13g2_nand2_1 _2696_ (.Y(_0789_),
    .A(_0524_),
    .B(_0525_));
 sg13g2_xnor2_1 _2697_ (.Y(_0790_),
    .A(_0660_),
    .B(_0789_));
 sg13g2_nand2_1 _2698_ (.Y(_0791_),
    .A(_0653_),
    .B(_0790_));
 sg13g2_nor3_1 _2699_ (.A(_1499_),
    .B(_0521_),
    .C(_0686_),
    .Y(_0792_));
 sg13g2_a21oi_1 _2700_ (.A1(net587),
    .A2(_0368_),
    .Y(_0793_),
    .B1(_0685_));
 sg13g2_a21o_1 _2701_ (.A2(_0793_),
    .A1(_1499_),
    .B1(_0792_),
    .X(_0794_));
 sg13g2_nor2_2 _2702_ (.A(_1471_),
    .B(_1517_),
    .Y(_0795_));
 sg13g2_o21ai_1 _2703_ (.B1(_0706_),
    .Y(_0796_),
    .A1(net572),
    .A2(_0513_));
 sg13g2_nand3_1 _2704_ (.B(_0483_),
    .C(_0513_),
    .A(net572),
    .Y(_0797_));
 sg13g2_nand2_1 _2705_ (.Y(_0798_),
    .A(_0660_),
    .B(_0670_));
 sg13g2_nand4_1 _2706_ (.B(_0796_),
    .C(_0797_),
    .A(net601),
    .Y(_0799_),
    .D(_0798_));
 sg13g2_nor2_2 _2707_ (.A(_1471_),
    .B(net589),
    .Y(_0800_));
 sg13g2_nand2b_1 _2708_ (.Y(_0801_),
    .B(_0800_),
    .A_N(_0684_));
 sg13g2_nand2_1 _2709_ (.Y(_0802_),
    .A(net577),
    .B(net589));
 sg13g2_inv_1 _2710_ (.Y(_0803_),
    .A(_0802_));
 sg13g2_nor3_1 _2711_ (.A(_0692_),
    .B(_0693_),
    .C(_0802_),
    .Y(_0804_));
 sg13g2_nor2_1 _2712_ (.A(_1471_),
    .B(_0697_),
    .Y(_0805_));
 sg13g2_and2_1 _2713_ (.A(net584),
    .B(_0701_),
    .X(_0806_));
 sg13g2_o21ai_1 _2714_ (.B1(_0701_),
    .Y(_0807_),
    .A1(net577),
    .A2(net584));
 sg13g2_nand2b_1 _2715_ (.Y(_0808_),
    .B(_0807_),
    .A_N(_0805_));
 sg13g2_nor3_1 _2716_ (.A(net589),
    .B(_0695_),
    .C(_0697_),
    .Y(_0809_));
 sg13g2_nor2_1 _2717_ (.A(_0808_),
    .B(_0809_),
    .Y(_0810_));
 sg13g2_nor2_1 _2718_ (.A(_0804_),
    .B(_0810_),
    .Y(_0811_));
 sg13g2_a221oi_1 _2719_ (.B2(_0811_),
    .C1(_0799_),
    .B1(_0801_),
    .A1(_0794_),
    .Y(_0812_),
    .A2(_0795_));
 sg13g2_a21o_2 _2720_ (.A2(_0812_),
    .A1(_0791_),
    .B1(_0788_),
    .X(_0813_));
 sg13g2_nand2_1 _2721_ (.Y(_0814_),
    .A(net613),
    .B(_0813_));
 sg13g2_o21ai_1 _2722_ (.B1(_0814_),
    .Y(_0815_),
    .A1(net613),
    .A2(net573));
 sg13g2_o21ai_1 _2723_ (.B1(net632),
    .Y(_0816_),
    .A1(\crp.datapath.aluSrc1SelMux.d1[3] ),
    .A2(net665));
 sg13g2_a21oi_1 _2724_ (.A1(_1357_),
    .A2(_0815_),
    .Y(_0817_),
    .B1(_0816_));
 sg13g2_a21o_1 _2725_ (.A2(net630),
    .A1(\crp.datapath.aluSrc1SelMux.d0[3] ),
    .B1(_0817_),
    .X(_0818_));
 sg13g2_nor2_1 _2726_ (.A(net685),
    .B(_0818_),
    .Y(_0819_));
 sg13g2_nand2_1 _2727_ (.Y(_0820_),
    .A(\crp.datapath.aluSrc1SelMux.d0[11] ),
    .B(net629));
 sg13g2_nor2_1 _2728_ (.A(net611),
    .B(_0509_),
    .Y(_0821_));
 sg13g2_nor2_1 _2729_ (.A(_0015_),
    .B(net647),
    .Y(_0822_));
 sg13g2_inv_1 _2730_ (.Y(_0823_),
    .A(_0822_));
 sg13g2_a22oi_1 _2731_ (.Y(_0824_),
    .B1(_1392_),
    .B2(\crp.datapath.aluSrc1SelMux.d1[11] ),
    .A2(net609),
    .A1(_1256_));
 sg13g2_nor2_1 _2732_ (.A(_0823_),
    .B(_0824_),
    .Y(_0825_));
 sg13g2_xnor2_1 _2733_ (.Y(_0826_),
    .A(_0822_),
    .B(_0824_));
 sg13g2_inv_1 _2734_ (.Y(_0827_),
    .A(_0826_));
 sg13g2_nand2b_1 _2735_ (.Y(_0828_),
    .B(_0764_),
    .A_N(_0765_));
 sg13g2_a21o_1 _2736_ (.A2(_0828_),
    .A1(_0773_),
    .B1(_0827_),
    .X(_0829_));
 sg13g2_nand3_1 _2737_ (.B(_0827_),
    .C(_0828_),
    .A(_0773_),
    .Y(_0830_));
 sg13g2_nand3_1 _2738_ (.B(_0829_),
    .C(_0830_),
    .A(_0671_),
    .Y(_0831_));
 sg13g2_a21oi_2 _2739_ (.B1(_0766_),
    .Y(_0832_),
    .A2(_0778_),
    .A1(_0768_));
 sg13g2_or2_1 _2740_ (.X(_0833_),
    .B(_0832_),
    .A(_0826_));
 sg13g2_a21oi_2 _2741_ (.B1(_0654_),
    .Y(_0834_),
    .A2(_0832_),
    .A1(_0826_));
 sg13g2_a21oi_2 _2742_ (.B1(_1375_),
    .Y(_0835_),
    .A2(_0834_),
    .A1(_0833_));
 sg13g2_a21oi_2 _2743_ (.B1(_0821_),
    .Y(_0836_),
    .A2(_0835_),
    .A1(_0831_));
 sg13g2_nor2_1 _2744_ (.A(\crp.datapath.aluSrc1SelMux.d1[11] ),
    .B(net666),
    .Y(_0837_));
 sg13g2_nor2_1 _2745_ (.A(net628),
    .B(_0837_),
    .Y(_0838_));
 sg13g2_o21ai_1 _2746_ (.B1(_0838_),
    .Y(_0839_),
    .A1(net627),
    .A2(_0836_));
 sg13g2_and2_1 _2747_ (.A(_0820_),
    .B(_0839_),
    .X(_0840_));
 sg13g2_a21oi_2 _2748_ (.B1(_0819_),
    .Y(uo_out[3]),
    .A2(net685),
    .A1(_0840_));
 sg13g2_nor2_1 _2749_ (.A(net611),
    .B(_0460_),
    .Y(_0841_));
 sg13g2_nand2b_1 _2750_ (.Y(_0842_),
    .B(_0661_),
    .A_N(_0581_));
 sg13g2_nand2b_1 _2751_ (.Y(_0843_),
    .B(_0581_),
    .A_N(_0661_));
 sg13g2_a21o_1 _2752_ (.A2(_0843_),
    .A1(_0842_),
    .B1(net601),
    .X(_0844_));
 sg13g2_nand2_1 _2753_ (.Y(_0845_),
    .A(_0527_),
    .B(_0581_));
 sg13g2_o21ai_1 _2754_ (.B1(_0653_),
    .Y(_0846_),
    .A1(_0527_),
    .A2(_0581_));
 sg13g2_nor2b_1 _2755_ (.A(_0846_),
    .B_N(_0845_),
    .Y(_0847_));
 sg13g2_o21ai_1 _2756_ (.B1(_0461_),
    .Y(_0848_),
    .A1(net586),
    .A2(net572));
 sg13g2_o21ai_1 _2757_ (.B1(net601),
    .Y(_0849_),
    .A1(_0482_),
    .A2(_0579_));
 sg13g2_a21oi_1 _2758_ (.A1(_0580_),
    .A2(_0706_),
    .Y(_0850_),
    .B1(_0849_));
 sg13g2_o21ai_1 _2759_ (.B1(_0850_),
    .Y(_0851_),
    .A1(_0581_),
    .A2(_0747_));
 sg13g2_nand2_1 _2760_ (.Y(_0852_),
    .A(net577),
    .B(_0478_));
 sg13g2_a21oi_1 _2761_ (.A1(_0808_),
    .A2(_0852_),
    .Y(_0853_),
    .B1(_0851_));
 sg13g2_a22oi_1 _2762_ (.Y(_0854_),
    .B1(_0848_),
    .B2(_0800_),
    .A2(_0803_),
    .A1(_0738_));
 sg13g2_o21ai_1 _2763_ (.B1(_0854_),
    .Y(_0855_),
    .A1(_1545_),
    .A2(_0795_));
 sg13g2_nand2_1 _2764_ (.Y(_0856_),
    .A(_0853_),
    .B(_0855_));
 sg13g2_o21ai_1 _2765_ (.B1(_0844_),
    .Y(_0857_),
    .A1(_0847_),
    .A2(_0856_));
 sg13g2_a21oi_2 _2766_ (.B1(_0841_),
    .Y(_0858_),
    .A2(_0857_),
    .A1(net611));
 sg13g2_nor2_1 _2767_ (.A(\crp.datapath.aluSrc1SelMux.d1[4] ),
    .B(net666),
    .Y(_0859_));
 sg13g2_nor2_1 _2768_ (.A(net628),
    .B(_0859_),
    .Y(_0860_));
 sg13g2_o21ai_1 _2769_ (.B1(_0860_),
    .Y(_0861_),
    .A1(net627),
    .A2(_0858_));
 sg13g2_o21ai_1 _2770_ (.B1(_0861_),
    .Y(_0862_),
    .A1(_1187_),
    .A2(net631));
 sg13g2_nor2_1 _2771_ (.A(net684),
    .B(_0862_),
    .Y(_0863_));
 sg13g2_nor2_1 _2772_ (.A(net613),
    .B(_0576_),
    .Y(_0864_));
 sg13g2_nor2_2 _2773_ (.A(_0020_),
    .B(net647),
    .Y(_0865_));
 sg13g2_inv_1 _2774_ (.Y(_0866_),
    .A(_0865_));
 sg13g2_a22oi_1 _2775_ (.Y(_0867_),
    .B1(_1392_),
    .B2(\crp.datapath.aluSrc1SelMux.d1[12] ),
    .A2(net609),
    .A1(_1257_));
 sg13g2_nor2_1 _2776_ (.A(_0866_),
    .B(_0867_),
    .Y(_0868_));
 sg13g2_or2_1 _2777_ (.X(_0869_),
    .B(_0867_),
    .A(_0865_));
 sg13g2_xnor2_1 _2778_ (.Y(_0870_),
    .A(_0865_),
    .B(_0867_));
 sg13g2_nand2_1 _2779_ (.Y(_0871_),
    .A(_0767_),
    .B(_0826_));
 sg13g2_or2_1 _2780_ (.X(_0872_),
    .B(_0871_),
    .A(_0769_));
 sg13g2_nor2_1 _2781_ (.A(_0771_),
    .B(_0871_),
    .Y(_0873_));
 sg13g2_a21oi_1 _2782_ (.A1(_0823_),
    .A2(_0824_),
    .Y(_0874_),
    .B1(_0828_));
 sg13g2_nor3_1 _2783_ (.A(_0825_),
    .B(_0873_),
    .C(_0874_),
    .Y(_0875_));
 sg13g2_o21ai_1 _2784_ (.B1(_0875_),
    .Y(_0876_),
    .A1(_0872_),
    .A2(_0668_));
 sg13g2_or2_1 _2785_ (.X(_0877_),
    .B(_0876_),
    .A(_0870_));
 sg13g2_a21oi_1 _2786_ (.A1(_0870_),
    .A2(_0876_),
    .Y(_0878_),
    .B1(net601));
 sg13g2_nand4_1 _2787_ (.B(_0721_),
    .C(_0768_),
    .A(_0651_),
    .Y(_0879_),
    .D(_0827_));
 sg13g2_nor2_1 _2788_ (.A(_0822_),
    .B(_0824_),
    .Y(_0880_));
 sg13g2_nand2b_1 _2789_ (.Y(_0881_),
    .B(_0777_),
    .A_N(_0766_));
 sg13g2_a21oi_1 _2790_ (.A1(_0764_),
    .A2(_0765_),
    .Y(_0882_),
    .B1(_0826_));
 sg13g2_a21oi_1 _2791_ (.A1(_0881_),
    .A2(_0882_),
    .Y(_0883_),
    .B1(_0880_));
 sg13g2_o21ai_1 _2792_ (.B1(_0883_),
    .Y(_0884_),
    .A1(_0879_),
    .A2(_0645_));
 sg13g2_inv_1 _2793_ (.Y(_0885_),
    .A(_0884_));
 sg13g2_nand2b_1 _2794_ (.Y(_0886_),
    .B(_0884_),
    .A_N(_0870_));
 sg13g2_a21oi_1 _2795_ (.A1(_0870_),
    .A2(_0885_),
    .Y(_0887_),
    .B1(_0654_));
 sg13g2_a22oi_1 _2796_ (.Y(_0888_),
    .B1(_0886_),
    .B2(_0887_),
    .A2(_0878_),
    .A1(_0877_));
 sg13g2_a21o_2 _2797_ (.A2(net613),
    .A1(_0888_),
    .B1(_0864_),
    .X(_0889_));
 sg13g2_o21ai_1 _2798_ (.B1(net631),
    .Y(_0890_),
    .A1(\crp.datapath.aluSrc1SelMux.d1[12] ),
    .A2(net665));
 sg13g2_a21oi_1 _2799_ (.A1(_1357_),
    .A2(_0889_),
    .Y(_0891_),
    .B1(_0890_));
 sg13g2_a21oi_1 _2800_ (.A1(\crp.datapath.aluSrc1SelMux.d0[12] ),
    .A2(net628),
    .Y(_0892_),
    .B1(_0891_));
 sg13g2_a21oi_2 _2801_ (.B1(_0863_),
    .Y(uo_out[4]),
    .A2(net685),
    .A1(_0892_));
 sg13g2_nand2_1 _2802_ (.Y(_0893_),
    .A(_0579_),
    .B(_0842_));
 sg13g2_xor2_1 _2803_ (.B(_0893_),
    .A(_0556_),
    .X(_0894_));
 sg13g2_nor2_1 _2804_ (.A(_0793_),
    .B(_0802_),
    .Y(_0895_));
 sg13g2_o21ai_1 _2805_ (.B1(_0690_),
    .Y(_0896_),
    .A1(_1471_),
    .A2(_1517_));
 sg13g2_nor2_1 _2806_ (.A(_0683_),
    .B(_0693_),
    .Y(_0897_));
 sg13g2_a21oi_1 _2807_ (.A1(_0800_),
    .A2(_0897_),
    .Y(_0898_),
    .B1(_0895_));
 sg13g2_or2_1 _2808_ (.X(_0899_),
    .B(_0807_),
    .A(_0694_));
 sg13g2_o21ai_1 _2809_ (.B1(_0806_),
    .Y(_0900_),
    .A1(_1471_),
    .A2(net590));
 sg13g2_o21ai_1 _2810_ (.B1(_0706_),
    .Y(_0901_),
    .A1(net583),
    .A2(_0553_));
 sg13g2_or2_1 _2811_ (.X(_0902_),
    .B(_0554_),
    .A(_0482_));
 sg13g2_nor2_1 _2812_ (.A(_0556_),
    .B(_0747_),
    .Y(_0903_));
 sg13g2_nand4_1 _2813_ (.B(_0900_),
    .C(_0901_),
    .A(_0899_),
    .Y(_0904_),
    .D(_0902_));
 sg13g2_a21oi_1 _2814_ (.A1(_0696_),
    .A2(_0805_),
    .Y(_0905_),
    .B1(_0903_));
 sg13g2_nand2b_1 _2815_ (.Y(_0906_),
    .B(_0905_),
    .A_N(_0904_));
 sg13g2_nand3b_1 _2816_ (.B(_0631_),
    .C(_0845_),
    .Y(_0907_),
    .A_N(_0556_));
 sg13g2_nor3_1 _2817_ (.A(_0583_),
    .B(_0632_),
    .C(_0654_),
    .Y(_0908_));
 sg13g2_a221oi_1 _2818_ (.B2(_0908_),
    .C1(_0906_),
    .B1(_0907_),
    .A1(_0896_),
    .Y(_0909_),
    .A2(_0898_));
 sg13g2_o21ai_1 _2819_ (.B1(_0909_),
    .Y(_0910_),
    .A1(net601),
    .A2(_0894_));
 sg13g2_inv_1 _2820_ (.Y(_0911_),
    .A(_0910_));
 sg13g2_mux2_2 _2821_ (.A0(net583),
    .A1(_0910_),
    .S(net611),
    .X(_0912_));
 sg13g2_nor2_1 _2822_ (.A(\crp.datapath.aluSrc1SelMux.d1[5] ),
    .B(net666),
    .Y(_0913_));
 sg13g2_nor2_1 _2823_ (.A(net628),
    .B(_0913_),
    .Y(_0914_));
 sg13g2_o21ai_1 _2824_ (.B1(_0914_),
    .Y(_0915_),
    .A1(net627),
    .A2(_0912_));
 sg13g2_o21ai_1 _2825_ (.B1(_0915_),
    .Y(_0916_),
    .A1(_1186_),
    .A2(net631));
 sg13g2_nor2_1 _2826_ (.A(net687),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_nor2_1 _2827_ (.A(net613),
    .B(_0549_),
    .Y(_0918_));
 sg13g2_a22oi_1 _2828_ (.Y(_0919_),
    .B1(_1392_),
    .B2(\crp.datapath.aluSrc1SelMux.d1[13] ),
    .A2(net609),
    .A1(_1258_));
 sg13g2_xnor2_1 _2829_ (.Y(_0920_),
    .A(_0865_),
    .B(_0919_));
 sg13g2_xnor2_1 _2830_ (.Y(_0921_),
    .A(_0866_),
    .B(_0919_));
 sg13g2_nand3_1 _2831_ (.B(_0869_),
    .C(_0920_),
    .A(_0886_),
    .Y(_0922_));
 sg13g2_a21o_1 _2832_ (.A2(_0886_),
    .A1(_0869_),
    .B1(_0920_),
    .X(_0923_));
 sg13g2_nand3_1 _2833_ (.B(_0923_),
    .C(_0922_),
    .A(_0653_),
    .Y(_0924_));
 sg13g2_a21oi_2 _2834_ (.B1(_0868_),
    .Y(_0925_),
    .A2(_0870_),
    .A1(_0876_));
 sg13g2_nand2b_1 _2835_ (.Y(_0926_),
    .B(_0920_),
    .A_N(_0925_));
 sg13g2_a21oi_1 _2836_ (.A1(_0921_),
    .A2(_0925_),
    .Y(_0927_),
    .B1(_0672_));
 sg13g2_a21oi_1 _2837_ (.A1(_0926_),
    .A2(_0927_),
    .Y(_0928_),
    .B1(_1375_));
 sg13g2_a21oi_2 _2838_ (.B1(_0918_),
    .Y(_0929_),
    .A2(_0924_),
    .A1(_0928_));
 sg13g2_or2_1 _2839_ (.X(_0930_),
    .B(net627),
    .A(_0929_));
 sg13g2_nor2_1 _2840_ (.A(\crp.datapath.aluSrc1SelMux.d1[13] ),
    .B(net666),
    .Y(_0931_));
 sg13g2_nor2_1 _2841_ (.A(net629),
    .B(_0931_),
    .Y(_0932_));
 sg13g2_a22oi_1 _2842_ (.Y(_0933_),
    .B1(_0930_),
    .B2(_0932_),
    .A2(net628),
    .A1(\crp.datapath.aluSrc1SelMux.d0[13] ));
 sg13g2_a21oi_2 _2843_ (.B1(_0917_),
    .Y(uo_out[5]),
    .A2(net687),
    .A1(_0933_));
 sg13g2_a21oi_1 _2844_ (.A1(_0661_),
    .A2(_0662_),
    .Y(_0934_),
    .B1(_0663_));
 sg13g2_xnor2_1 _2845_ (.Y(_0935_),
    .A(_0639_),
    .B(_0934_));
 sg13g2_nand3b_1 _2846_ (.B(_0633_),
    .C(_0638_),
    .Y(_0936_),
    .A_N(_0583_));
 sg13g2_o21ai_1 _2847_ (.B1(_0639_),
    .Y(_0937_),
    .A1(_0583_),
    .A2(_0634_));
 sg13g2_nand3_1 _2848_ (.B(_0936_),
    .C(_0937_),
    .A(_0653_),
    .Y(_0938_));
 sg13g2_o21ai_1 _2849_ (.B1(_0426_),
    .Y(_0939_),
    .A1(net586),
    .A2(net583));
 sg13g2_a22oi_1 _2850_ (.Y(_0940_),
    .B1(_0939_),
    .B2(_0800_),
    .A2(_0848_),
    .A1(_0803_));
 sg13g2_o21ai_1 _2851_ (.B1(_0940_),
    .Y(_0941_),
    .A1(_0740_),
    .A2(_0795_));
 sg13g2_a21oi_1 _2852_ (.A1(_0748_),
    .A2(_0808_),
    .Y(_0942_),
    .B1(net602));
 sg13g2_o21ai_1 _2853_ (.B1(_0900_),
    .Y(_0943_),
    .A1(_0482_),
    .A2(_0636_));
 sg13g2_a221oi_1 _2854_ (.B2(_0637_),
    .C1(_0943_),
    .B1(_0706_),
    .A1(_0638_),
    .Y(_0944_),
    .A2(_0670_));
 sg13g2_and3_1 _2855_ (.X(_0945_),
    .A(_0941_),
    .B(_0942_),
    .C(_0944_));
 sg13g2_a22oi_1 _2856_ (.Y(_0946_),
    .B1(_0938_),
    .B2(_0945_),
    .A2(_0935_),
    .A1(net602));
 sg13g2_mux2_2 _2857_ (.A0(_0424_),
    .A1(_0946_),
    .S(net611),
    .X(_0947_));
 sg13g2_nor2_1 _2858_ (.A(\crp.datapath.aluSrc1SelMux.d1[6] ),
    .B(net666),
    .Y(_0948_));
 sg13g2_nor2_1 _2859_ (.A(net628),
    .B(_0948_),
    .Y(_0949_));
 sg13g2_o21ai_1 _2860_ (.B1(_0949_),
    .Y(_0950_),
    .A1(net627),
    .A2(_0947_));
 sg13g2_o21ai_1 _2861_ (.B1(_0950_),
    .Y(_0951_),
    .A1(_1185_),
    .A2(net631));
 sg13g2_nor2_1 _2862_ (.A(net613),
    .B(_0625_),
    .Y(_0952_));
 sg13g2_a22oi_1 _2863_ (.Y(_0953_),
    .B1(_1392_),
    .B2(\crp.datapath.aluSrc1SelMux.d1[14] ),
    .A2(net609),
    .A1(_1259_));
 sg13g2_xnor2_1 _2864_ (.Y(_0954_),
    .A(_0866_),
    .B(_0953_));
 sg13g2_nand3_1 _2865_ (.B(_0920_),
    .C(_0876_),
    .A(_0870_),
    .Y(_0955_));
 sg13g2_a21o_1 _2866_ (.A2(_0919_),
    .A1(_0867_),
    .B1(_0866_),
    .X(_0956_));
 sg13g2_nand3_1 _2867_ (.B(_0955_),
    .C(_0956_),
    .A(_0954_),
    .Y(_0957_));
 sg13g2_a21o_1 _2868_ (.A2(_0955_),
    .A1(_0956_),
    .B1(_0954_),
    .X(_0958_));
 sg13g2_nand3_1 _2869_ (.B(_0957_),
    .C(_0958_),
    .A(net602),
    .Y(_0959_));
 sg13g2_nor2_1 _2870_ (.A(_0870_),
    .B(_0920_),
    .Y(_0960_));
 sg13g2_a21oi_1 _2871_ (.A1(_0867_),
    .A2(_0919_),
    .Y(_0961_),
    .B1(_0865_));
 sg13g2_a21o_1 _2872_ (.A2(_0884_),
    .A1(_0960_),
    .B1(_0961_),
    .X(_0962_));
 sg13g2_or2_1 _2873_ (.X(_0963_),
    .B(_0962_),
    .A(_0954_));
 sg13g2_a21oi_2 _2874_ (.B1(_0654_),
    .Y(_0964_),
    .A2(_0962_),
    .A1(_0954_));
 sg13g2_a21oi_2 _2875_ (.B1(_1375_),
    .Y(_0965_),
    .A2(_0963_),
    .A1(_0964_));
 sg13g2_a21oi_2 _2876_ (.B1(_0952_),
    .Y(_0966_),
    .A2(_0959_),
    .A1(_0965_));
 sg13g2_nor2_1 _2877_ (.A(\crp.datapath.aluSrc1SelMux.d1[14] ),
    .B(net666),
    .Y(_0967_));
 sg13g2_nor2_1 _2878_ (.A(net628),
    .B(_0967_),
    .Y(_0968_));
 sg13g2_o21ai_1 _2879_ (.B1(_0968_),
    .Y(_0969_),
    .A1(_0966_),
    .A2(net627));
 sg13g2_o21ai_1 _2880_ (.B1(_0969_),
    .Y(_0970_),
    .A1(_1180_),
    .A2(net631));
 sg13g2_mux2_2 _2881_ (.A0(_0951_),
    .A1(_0970_),
    .S(net684),
    .X(uo_out[6]));
 sg13g2_nand2b_1 _2882_ (.Y(_0971_),
    .B(_1375_),
    .A_N(net584));
 sg13g2_o21ai_1 _2883_ (.B1(_0636_),
    .Y(_0972_),
    .A1(_0639_),
    .A2(_0934_));
 sg13g2_xor2_1 _2884_ (.B(_0972_),
    .A(_0643_),
    .X(_0973_));
 sg13g2_nor2_1 _2885_ (.A(net578),
    .B(_1517_),
    .Y(_0974_));
 sg13g2_nand2_1 _2886_ (.Y(_0975_),
    .A(net589),
    .B(_0897_));
 sg13g2_nand3b_1 _2887_ (.B(_0695_),
    .C(_1499_),
    .Y(_0976_),
    .A_N(_0692_));
 sg13g2_nand3_1 _2888_ (.B(_0975_),
    .C(_0976_),
    .A(_0795_),
    .Y(_0977_));
 sg13g2_a22oi_1 _2889_ (.Y(_0978_),
    .B1(_0642_),
    .B2(_0706_),
    .A2(_0641_),
    .A1(_0483_));
 sg13g2_nand2b_1 _2890_ (.Y(_0979_),
    .B(_0978_),
    .A_N(_0806_));
 sg13g2_a21oi_1 _2891_ (.A1(net577),
    .A2(_0809_),
    .Y(_0980_),
    .B1(_0979_));
 sg13g2_nand2_1 _2892_ (.Y(_0981_),
    .A(_0977_),
    .B(_0980_));
 sg13g2_a221oi_1 _2893_ (.B2(_0974_),
    .C1(_0981_),
    .B1(_0794_),
    .A1(_0643_),
    .Y(_0982_),
    .A2(_0746_));
 sg13g2_nand2_1 _2894_ (.Y(_0983_),
    .A(_0628_),
    .B(_0937_));
 sg13g2_xnor2_1 _2895_ (.Y(_0984_),
    .A(_0643_),
    .B(_0983_));
 sg13g2_a22oi_1 _2896_ (.Y(_0985_),
    .B1(_0984_),
    .B2(_0653_),
    .A2(_0973_),
    .A1(net602));
 sg13g2_nand2_2 _2897_ (.Y(_0986_),
    .A(_0982_),
    .B(_0985_));
 sg13g2_inv_1 _2898_ (.Y(_0987_),
    .A(_0986_));
 sg13g2_o21ai_1 _2899_ (.B1(_0971_),
    .Y(_0988_),
    .A1(_1375_),
    .A2(_0986_));
 sg13g2_o21ai_1 _2900_ (.B1(net631),
    .Y(_0989_),
    .A1(\crp.datapath.aluSrc1SelMux.d1[7] ),
    .A2(net665));
 sg13g2_a21oi_1 _2901_ (.A1(_1357_),
    .A2(_0988_),
    .Y(_0990_),
    .B1(_0989_));
 sg13g2_a21oi_1 _2902_ (.A1(\crp.datapath.aluSrc1SelMux.d0[7] ),
    .A2(net630),
    .Y(_0991_),
    .B1(_0990_));
 sg13g2_nor2_2 _2903_ (.A(net685),
    .B(_0991_),
    .Y(uo_out[7]));
 sg13g2_nand2_1 _2904_ (.Y(_0992_),
    .A(net686),
    .B(_0491_));
 sg13g2_o21ai_1 _2905_ (.B1(_0992_),
    .Y(uio_out[0]),
    .A1(_0680_),
    .A2(net687));
 sg13g2_nor2_2 _2906_ (.A(net686),
    .B(_0736_),
    .Y(_0993_));
 sg13g2_a21oi_2 _2907_ (.B1(_0993_),
    .Y(uio_out[1]),
    .A2(_0715_),
    .A1(net685));
 sg13g2_nand2_1 _2908_ (.Y(_0994_),
    .A(net686),
    .B(_0761_));
 sg13g2_o21ai_1 _2909_ (.B1(_0994_),
    .Y(uio_out[2]),
    .A1(_0786_),
    .A2(net684));
 sg13g2_nand2_1 _2910_ (.Y(_0995_),
    .A(net685),
    .B(_0818_));
 sg13g2_o21ai_1 _2911_ (.B1(_0995_),
    .Y(uio_out[3]),
    .A1(net684),
    .A2(_0840_));
 sg13g2_nand2_1 _2912_ (.Y(_0996_),
    .A(net687),
    .B(_0862_));
 sg13g2_o21ai_1 _2913_ (.B1(_0996_),
    .Y(uio_out[4]),
    .A1(_0892_),
    .A2(net684));
 sg13g2_nand2_1 _2914_ (.Y(_0997_),
    .A(net684),
    .B(_0916_));
 sg13g2_o21ai_1 _2915_ (.B1(_0997_),
    .Y(uio_out[5]),
    .A1(_0933_),
    .A2(net684));
 sg13g2_mux2_2 _2916_ (.A0(_0970_),
    .A1(_0951_),
    .S(net684),
    .X(uio_out[6]));
 sg13g2_a21oi_1 _2917_ (.A1(_1326_),
    .A2(_1327_),
    .Y(_0998_),
    .B1(_1507_));
 sg13g2_a21o_1 _2918_ (.A2(_1378_),
    .A1(_1343_),
    .B1(_0998_),
    .X(\crp.controller.mainDecoder.memWriteReq ));
 sg13g2_o21ai_1 _2919_ (.B1(_1291_),
    .Y(_0999_),
    .A1(_1290_),
    .A2(_1325_));
 sg13g2_nor2_1 _2920_ (.A(net693),
    .B(_1377_),
    .Y(_1000_));
 sg13g2_a22oi_1 _2921_ (.Y(_1001_),
    .B1(_1000_),
    .B2(_1272_),
    .A2(_0999_),
    .A1(net694));
 sg13g2_nor2_2 _2922_ (.A(\crp.datapath.aluSrc2SelMux.d3[10] ),
    .B(\crp.datapath.aluSrc2SelMux.d3[9] ),
    .Y(_1002_));
 sg13g2_nand4_1 _2923_ (.B(_1168_),
    .C(net608),
    .A(_1167_),
    .Y(_1003_),
    .D(_1002_));
 sg13g2_o21ai_1 _2924_ (.B1(_1377_),
    .Y(_1004_),
    .A1(_1280_),
    .A2(_1325_));
 sg13g2_inv_1 _2925_ (.Y(_1005_),
    .A(_1004_));
 sg13g2_and2_1 _2926_ (.A(net694),
    .B(_1320_),
    .X(_1006_));
 sg13g2_nor3_1 _2927_ (.A(net692),
    .B(_1005_),
    .C(net667),
    .Y(_1007_));
 sg13g2_o21ai_1 _2928_ (.B1(net667),
    .Y(_1008_),
    .A1(_1526_),
    .A2(_1541_));
 sg13g2_nor3_2 _2929_ (.A(net693),
    .B(_1004_),
    .C(_1006_),
    .Y(_1009_));
 sg13g2_a221oi_1 _2930_ (.B2(\crp.datapath.memReadData[0] ),
    .C1(net600),
    .B1(_1009_),
    .A1(net727),
    .Y(_1010_),
    .A2(net692));
 sg13g2_a22oi_1 _2931_ (.Y(_1011_),
    .B1(_1008_),
    .B2(_1010_),
    .A2(net599),
    .A1(_0487_));
 sg13g2_mux2_1 _2932_ (.A0(net568),
    .A1(net325),
    .S(_1003_),
    .X(_0156_));
 sg13g2_nand2b_1 _2933_ (.Y(_1012_),
    .B(net599),
    .A_N(_0710_));
 sg13g2_nand2b_1 _2934_ (.Y(_1013_),
    .B(net667),
    .A_N(_1496_));
 sg13g2_a22oi_1 _2935_ (.Y(_1014_),
    .B1(_1009_),
    .B2(\crp.datapath.memReadData[1] ),
    .A2(net692),
    .A1(net726));
 sg13g2_nand3_1 _2936_ (.B(_1013_),
    .C(_1014_),
    .A(_1012_),
    .Y(_1015_));
 sg13g2_mux2_1 _2937_ (.A0(net564),
    .A1(net340),
    .S(_1003_),
    .X(_0157_));
 sg13g2_nand2_1 _2938_ (.Y(_1016_),
    .A(_0756_),
    .B(net600));
 sg13g2_nand2_1 _2939_ (.Y(_1017_),
    .A(net725),
    .B(net692));
 sg13g2_a22oi_1 _2940_ (.Y(_1018_),
    .B1(_1009_),
    .B2(\crp.datapath.memReadData[2] ),
    .A2(net667),
    .A1(_1467_));
 sg13g2_nand3_1 _2941_ (.B(_1017_),
    .C(_1018_),
    .A(_1016_),
    .Y(_1019_));
 sg13g2_mux2_1 _2942_ (.A0(net562),
    .A1(net346),
    .S(_1003_),
    .X(_0158_));
 sg13g2_nand2_1 _2943_ (.Y(_1020_),
    .A(_0509_),
    .B(_1006_));
 sg13g2_a22oi_1 _2944_ (.Y(_1021_),
    .B1(_1009_),
    .B2(\crp.datapath.memReadData[3] ),
    .A2(_1004_),
    .A1(net722));
 sg13g2_nand2_1 _2945_ (.Y(_1022_),
    .A(_1020_),
    .B(_1021_));
 sg13g2_nor2_1 _2946_ (.A(net600),
    .B(_1022_),
    .Y(_1023_));
 sg13g2_a21oi_2 _2947_ (.B1(_1023_),
    .Y(_1024_),
    .A2(net599),
    .A1(_0813_));
 sg13g2_mux2_1 _2948_ (.A0(net570),
    .A1(net301),
    .S(_1003_),
    .X(_0159_));
 sg13g2_nand2b_1 _2949_ (.Y(_1025_),
    .B(net599),
    .A_N(_0857_));
 sg13g2_nand2_1 _2950_ (.Y(_1026_),
    .A(\crp.datapath.aluSrc2SelMux.d2[4] ),
    .B(net692));
 sg13g2_a22oi_1 _2951_ (.Y(_1027_),
    .B1(_1009_),
    .B2(\crp.datapath.memReadData[4] ),
    .A2(net667),
    .A1(_0576_));
 sg13g2_nand3_1 _2952_ (.B(_1026_),
    .C(_1027_),
    .A(_1025_),
    .Y(_1028_));
 sg13g2_mux2_1 _2953_ (.A0(net560),
    .A1(net261),
    .S(_1003_),
    .X(_0160_));
 sg13g2_nand2_1 _2954_ (.Y(_1029_),
    .A(_0549_),
    .B(net667));
 sg13g2_a221oi_1 _2955_ (.B2(\crp.datapath.memReadData[5] ),
    .C1(net600),
    .B1(_1009_),
    .A1(\crp.datapath.aluSrc2SelMux.d2[5] ),
    .Y(_1030_),
    .A2(net692));
 sg13g2_a22oi_1 _2956_ (.Y(_1031_),
    .B1(_1029_),
    .B2(_1030_),
    .A2(net599),
    .A1(_0911_));
 sg13g2_mux2_1 _2957_ (.A0(net558),
    .A1(net253),
    .S(_1003_),
    .X(_0161_));
 sg13g2_nand2_1 _2958_ (.Y(_1032_),
    .A(_0946_),
    .B(net599));
 sg13g2_nand2_1 _2959_ (.Y(_1033_),
    .A(_0625_),
    .B(net667));
 sg13g2_a22oi_1 _2960_ (.Y(_1034_),
    .B1(_1009_),
    .B2(\crp.datapath.memReadData[6] ),
    .A2(net692),
    .A1(\crp.datapath.aluSrc2SelMux.d2[6] ));
 sg13g2_nand3_1 _2961_ (.B(_1033_),
    .C(_1034_),
    .A(_1032_),
    .Y(_1035_));
 sg13g2_mux2_1 _2962_ (.A0(net566),
    .A1(net251),
    .S(_1003_),
    .X(_0162_));
 sg13g2_nand2_1 _2963_ (.Y(_1036_),
    .A(_0602_),
    .B(net667));
 sg13g2_a221oi_1 _2964_ (.B2(\crp.datapath.memReadData[7] ),
    .C1(net599),
    .B1(_1009_),
    .A1(\crp.datapath.aluSrc2SelMux.d2[7] ),
    .Y(_1037_),
    .A2(net692));
 sg13g2_a22oi_1 _2965_ (.Y(_1038_),
    .B1(_1036_),
    .B2(_1037_),
    .A2(net599),
    .A1(_0987_));
 sg13g2_mux2_1 _2966_ (.A0(net556),
    .A1(net232),
    .S(_1003_),
    .X(_0163_));
 sg13g2_nor2_2 _2967_ (.A(_1169_),
    .B(\crp.datapath.aluSrc2SelMux.d3[9] ),
    .Y(_1039_));
 sg13g2_nand4_1 _2968_ (.B(_1168_),
    .C(net608),
    .A(_1167_),
    .Y(_1040_),
    .D(_1039_));
 sg13g2_nor2_1 _2969_ (.A(net568),
    .B(net598),
    .Y(_1041_));
 sg13g2_a21oi_1 _2970_ (.A1(_1192_),
    .A2(net598),
    .Y(_0164_),
    .B1(_1041_));
 sg13g2_mux2_1 _2971_ (.A0(net564),
    .A1(net336),
    .S(net598),
    .X(_0165_));
 sg13g2_mux2_1 _2972_ (.A0(net562),
    .A1(net319),
    .S(net598),
    .X(_0166_));
 sg13g2_mux2_1 _2973_ (.A0(net570),
    .A1(net242),
    .S(net598),
    .X(_0167_));
 sg13g2_mux2_1 _2974_ (.A0(net560),
    .A1(net264),
    .S(net598),
    .X(_0168_));
 sg13g2_mux2_1 _2975_ (.A0(net558),
    .A1(net276),
    .S(net598),
    .X(_0169_));
 sg13g2_mux2_1 _2976_ (.A0(net566),
    .A1(net313),
    .S(net598),
    .X(_0170_));
 sg13g2_mux2_1 _2977_ (.A0(net556),
    .A1(net239),
    .S(_1040_),
    .X(_0171_));
 sg13g2_nor2_2 _2978_ (.A(\crp.datapath.aluSrc2SelMux.d3[10] ),
    .B(_1170_),
    .Y(_1042_));
 sg13g2_nand4_1 _2979_ (.B(_1168_),
    .C(net608),
    .A(_1167_),
    .Y(_1043_),
    .D(_1042_));
 sg13g2_mux2_1 _2980_ (.A0(net568),
    .A1(net331),
    .S(net597),
    .X(_0172_));
 sg13g2_mux2_1 _2981_ (.A0(net564),
    .A1(net323),
    .S(net597),
    .X(_0173_));
 sg13g2_nor2_1 _2982_ (.A(net562),
    .B(net597),
    .Y(_1044_));
 sg13g2_a21oi_1 _2983_ (.A1(_1217_),
    .A2(net597),
    .Y(_0174_),
    .B1(_1044_));
 sg13g2_mux2_1 _2984_ (.A0(net570),
    .A1(net289),
    .S(net597),
    .X(_0175_));
 sg13g2_mux2_1 _2985_ (.A0(net560),
    .A1(net263),
    .S(net597),
    .X(_0176_));
 sg13g2_mux2_1 _2986_ (.A0(net558),
    .A1(net252),
    .S(net597),
    .X(_0177_));
 sg13g2_mux2_1 _2987_ (.A0(net566),
    .A1(net302),
    .S(net597),
    .X(_0178_));
 sg13g2_mux2_1 _2988_ (.A0(net556),
    .A1(net254),
    .S(_1043_),
    .X(_0179_));
 sg13g2_nor2_2 _2989_ (.A(_1167_),
    .B(net393),
    .Y(_1045_));
 sg13g2_nand3_1 _2990_ (.B(_1002_),
    .C(_1045_),
    .A(_1001_),
    .Y(_1046_));
 sg13g2_mux2_1 _2991_ (.A0(net569),
    .A1(net328),
    .S(_1046_),
    .X(_0180_));
 sg13g2_mux2_1 _2992_ (.A0(net565),
    .A1(net357),
    .S(_1046_),
    .X(_0181_));
 sg13g2_mux2_1 _2993_ (.A0(net563),
    .A1(net341),
    .S(_1046_),
    .X(_0182_));
 sg13g2_mux2_1 _2994_ (.A0(net571),
    .A1(net286),
    .S(_1046_),
    .X(_0183_));
 sg13g2_mux2_1 _2995_ (.A0(net561),
    .A1(net294),
    .S(_1046_),
    .X(_0184_));
 sg13g2_mux2_1 _2996_ (.A0(net559),
    .A1(net269),
    .S(_1046_),
    .X(_0185_));
 sg13g2_mux2_1 _2997_ (.A0(net567),
    .A1(net258),
    .S(_1046_),
    .X(_0186_));
 sg13g2_mux2_1 _2998_ (.A0(net557),
    .A1(net290),
    .S(_1046_),
    .X(_0187_));
 sg13g2_and3_2 _2999_ (.X(_1047_),
    .A(\crp.datapath.aluSrc2SelMux.d3[12] ),
    .B(\crp.datapath.aluSrc2SelMux.d3[11] ),
    .C(_1001_));
 sg13g2_nand3_1 _3000_ (.B(\crp.datapath.aluSrc2SelMux.d3[9] ),
    .C(_1047_),
    .A(\crp.datapath.aluSrc2SelMux.d3[10] ),
    .Y(_1048_));
 sg13g2_nor2_1 _3001_ (.A(net569),
    .B(net582),
    .Y(_1049_));
 sg13g2_a21oi_1 _3002_ (.A1(_1206_),
    .A2(net582),
    .Y(_0188_),
    .B1(_1049_));
 sg13g2_mux2_1 _3003_ (.A0(net565),
    .A1(net353),
    .S(net582),
    .X(_0189_));
 sg13g2_mux2_1 _3004_ (.A0(net563),
    .A1(net327),
    .S(net582),
    .X(_0190_));
 sg13g2_mux2_1 _3005_ (.A0(net571),
    .A1(net281),
    .S(net582),
    .X(_0191_));
 sg13g2_mux2_1 _3006_ (.A0(net561),
    .A1(net306),
    .S(net582),
    .X(_0192_));
 sg13g2_mux2_1 _3007_ (.A0(net559),
    .A1(net233),
    .S(net582),
    .X(_0193_));
 sg13g2_mux2_1 _3008_ (.A0(net567),
    .A1(net310),
    .S(net582),
    .X(_0194_));
 sg13g2_mux2_1 _3009_ (.A0(net557),
    .A1(net295),
    .S(_1048_),
    .X(_0195_));
 sg13g2_nand2_1 _3010_ (.Y(_1050_),
    .A(_1039_),
    .B(_1047_));
 sg13g2_nor2_1 _3011_ (.A(net569),
    .B(net581),
    .Y(_1051_));
 sg13g2_a21oi_1 _3012_ (.A1(_1205_),
    .A2(net581),
    .Y(_0196_),
    .B1(_1051_));
 sg13g2_mux2_1 _3013_ (.A0(net565),
    .A1(net348),
    .S(net581),
    .X(_0197_));
 sg13g2_mux2_1 _3014_ (.A0(net563),
    .A1(net351),
    .S(net581),
    .X(_0198_));
 sg13g2_mux2_1 _3015_ (.A0(net571),
    .A1(net272),
    .S(net581),
    .X(_0199_));
 sg13g2_mux2_1 _3016_ (.A0(net561),
    .A1(net277),
    .S(_1050_),
    .X(_0200_));
 sg13g2_mux2_1 _3017_ (.A0(net559),
    .A1(net238),
    .S(net581),
    .X(_0201_));
 sg13g2_mux2_1 _3018_ (.A0(net567),
    .A1(net262),
    .S(net581),
    .X(_0202_));
 sg13g2_mux2_1 _3019_ (.A0(net557),
    .A1(net274),
    .S(net581),
    .X(_0203_));
 sg13g2_and2_1 _3020_ (.A(net1),
    .B(net745),
    .X(_0204_));
 sg13g2_nor2_1 _3021_ (.A(_1161_),
    .B(net736),
    .Y(_0205_));
 sg13g2_nor2_1 _3022_ (.A(_1159_),
    .B(net736),
    .Y(_0206_));
 sg13g2_and2_1 _3023_ (.A(net4),
    .B(net743),
    .X(_0207_));
 sg13g2_and2_1 _3024_ (.A(net5),
    .B(net743),
    .X(_0208_));
 sg13g2_and2_1 _3025_ (.A(net6),
    .B(net743),
    .X(_0209_));
 sg13g2_and2_1 _3026_ (.A(net7),
    .B(net743),
    .X(_0210_));
 sg13g2_and2_1 _3027_ (.A(net8),
    .B(net742),
    .X(_0211_));
 sg13g2_nand2_1 _3028_ (.Y(_1052_),
    .A(_1042_),
    .B(_1047_));
 sg13g2_nor2_1 _3029_ (.A(net569),
    .B(net580),
    .Y(_1053_));
 sg13g2_a21oi_1 _3030_ (.A1(_1203_),
    .A2(net580),
    .Y(_0212_),
    .B1(_1053_));
 sg13g2_mux2_1 _3031_ (.A0(net565),
    .A1(net326),
    .S(net580),
    .X(_0213_));
 sg13g2_mux2_1 _3032_ (.A0(net563),
    .A1(net344),
    .S(net580),
    .X(_0214_));
 sg13g2_mux2_1 _3033_ (.A0(net571),
    .A1(net246),
    .S(net580),
    .X(_0215_));
 sg13g2_mux2_1 _3034_ (.A0(net561),
    .A1(net280),
    .S(_1052_),
    .X(_0216_));
 sg13g2_mux2_1 _3035_ (.A0(net559),
    .A1(net234),
    .S(net580),
    .X(_0217_));
 sg13g2_mux2_1 _3036_ (.A0(net567),
    .A1(net240),
    .S(net580),
    .X(_0218_));
 sg13g2_mux2_1 _3037_ (.A0(net557),
    .A1(net248),
    .S(net580),
    .X(_0219_));
 sg13g2_o21ai_1 _3038_ (.B1(net647),
    .Y(_1054_),
    .A1(_1315_),
    .A2(_1369_));
 sg13g2_nor2_1 _3039_ (.A(_1260_),
    .B(_1054_),
    .Y(_1055_));
 sg13g2_or2_1 _3040_ (.X(_1056_),
    .B(_1054_),
    .A(_1260_));
 sg13g2_o21ai_1 _3041_ (.B1(net742),
    .Y(_1057_),
    .A1(net361),
    .A2(net604));
 sg13g2_a21oi_1 _3042_ (.A1(_0488_),
    .A2(net604),
    .Y(_0220_),
    .B1(_1057_));
 sg13g2_o21ai_1 _3043_ (.B1(net742),
    .Y(_1058_),
    .A1(net366),
    .A2(net604));
 sg13g2_a21oi_1 _3044_ (.A1(_0712_),
    .A2(net604),
    .Y(_0221_),
    .B1(_1058_));
 sg13g2_o21ai_1 _3045_ (.B1(net742),
    .Y(_1059_),
    .A1(_0757_),
    .A2(net607));
 sg13g2_a21oi_1 _3046_ (.A1(_1188_),
    .A2(net607),
    .Y(_0222_),
    .B1(_1059_));
 sg13g2_o21ai_1 _3047_ (.B1(net740),
    .Y(_1060_),
    .A1(net354),
    .A2(net603));
 sg13g2_a21oi_1 _3048_ (.A1(_0815_),
    .A2(net603),
    .Y(_0223_),
    .B1(_1060_));
 sg13g2_o21ai_1 _3049_ (.B1(net740),
    .Y(_1061_),
    .A1(_0858_),
    .A2(net606));
 sg13g2_a21oi_1 _3050_ (.A1(_1187_),
    .A2(net606),
    .Y(_0224_),
    .B1(_1061_));
 sg13g2_o21ai_1 _3051_ (.B1(net740),
    .Y(_1062_),
    .A1(_0912_),
    .A2(net606));
 sg13g2_a21oi_1 _3052_ (.A1(_1186_),
    .A2(net606),
    .Y(_0225_),
    .B1(_1062_));
 sg13g2_o21ai_1 _3053_ (.B1(net740),
    .Y(_1063_),
    .A1(_0947_),
    .A2(net606));
 sg13g2_a21oi_1 _3054_ (.A1(_1185_),
    .A2(net606),
    .Y(_0226_),
    .B1(_1063_));
 sg13g2_o21ai_1 _3055_ (.B1(net740),
    .Y(_1064_),
    .A1(net359),
    .A2(net603));
 sg13g2_a21oi_1 _3056_ (.A1(_0988_),
    .A2(net603),
    .Y(_0227_),
    .B1(_1064_));
 sg13g2_o21ai_1 _3057_ (.B1(net740),
    .Y(_1065_),
    .A1(net372),
    .A2(net603));
 sg13g2_a21oi_1 _3058_ (.A1(_0677_),
    .A2(net603),
    .Y(_0228_),
    .B1(_1065_));
 sg13g2_o21ai_1 _3059_ (.B1(net741),
    .Y(_1066_),
    .A1(_0732_),
    .A2(net605));
 sg13g2_a21oi_1 _3060_ (.A1(_1184_),
    .A2(net607),
    .Y(_0229_),
    .B1(_1066_));
 sg13g2_o21ai_1 _3061_ (.B1(net741),
    .Y(_1067_),
    .A1(_0782_),
    .A2(net605));
 sg13g2_a21oi_1 _3062_ (.A1(_1183_),
    .A2(net605),
    .Y(_0230_),
    .B1(_1067_));
 sg13g2_o21ai_1 _3063_ (.B1(net741),
    .Y(_1068_),
    .A1(_0836_),
    .A2(net605));
 sg13g2_a21oi_1 _3064_ (.A1(_1182_),
    .A2(net605),
    .Y(_0231_),
    .B1(_1068_));
 sg13g2_o21ai_1 _3065_ (.B1(net741),
    .Y(_1069_),
    .A1(net363),
    .A2(net603));
 sg13g2_a21oi_1 _3066_ (.A1(_0889_),
    .A2(net603),
    .Y(_0232_),
    .B1(_1069_));
 sg13g2_o21ai_1 _3067_ (.B1(net740),
    .Y(_1070_),
    .A1(_0929_),
    .A2(net605));
 sg13g2_a21oi_1 _3068_ (.A1(_1181_),
    .A2(net605),
    .Y(_0233_),
    .B1(_1070_));
 sg13g2_o21ai_1 _3069_ (.B1(net740),
    .Y(_1071_),
    .A1(_0966_),
    .A2(net606));
 sg13g2_a21oi_1 _3070_ (.A1(_1180_),
    .A2(net605),
    .Y(_0234_),
    .B1(_1071_));
 sg13g2_nand2_2 _3071_ (.Y(_1072_),
    .A(_1002_),
    .B(_1047_));
 sg13g2_nor2_1 _3072_ (.A(net569),
    .B(net579),
    .Y(_1073_));
 sg13g2_a21oi_1 _3073_ (.A1(_1202_),
    .A2(net579),
    .Y(_0235_),
    .B1(_1073_));
 sg13g2_mux2_1 _3074_ (.A0(net565),
    .A1(net338),
    .S(net579),
    .X(_0236_));
 sg13g2_mux2_1 _3075_ (.A0(net563),
    .A1(net342),
    .S(net579),
    .X(_0237_));
 sg13g2_mux2_1 _3076_ (.A0(net571),
    .A1(net283),
    .S(net579),
    .X(_0238_));
 sg13g2_mux2_1 _3077_ (.A0(net561),
    .A1(net256),
    .S(_1072_),
    .X(_0239_));
 sg13g2_mux2_1 _3078_ (.A0(net559),
    .A1(net241),
    .S(net579),
    .X(_0240_));
 sg13g2_mux2_1 _3079_ (.A0(net567),
    .A1(net231),
    .S(net579),
    .X(_0241_));
 sg13g2_mux2_1 _3080_ (.A0(net557),
    .A1(net250),
    .S(net579),
    .X(_0242_));
 sg13g2_nor2_1 _3081_ (.A(_1359_),
    .B(_1386_),
    .Y(_1074_));
 sg13g2_or2_1 _3082_ (.X(_1075_),
    .B(_1386_),
    .A(_1359_));
 sg13g2_a21oi_1 _3083_ (.A1(net379),
    .A2(net617),
    .Y(_1076_),
    .B1(net737));
 sg13g2_o21ai_1 _3084_ (.B1(_1076_),
    .Y(_0243_),
    .A1(_0488_),
    .A2(net616));
 sg13g2_a21oi_1 _3085_ (.A1(net383),
    .A2(net617),
    .Y(_1077_),
    .B1(net737));
 sg13g2_o21ai_1 _3086_ (.B1(_1077_),
    .Y(_0244_),
    .A1(_0712_),
    .A2(net616));
 sg13g2_a21oi_1 _3087_ (.A1(_0757_),
    .A2(net620),
    .Y(_1078_),
    .B1(net737));
 sg13g2_o21ai_1 _3088_ (.B1(_1078_),
    .Y(_0245_),
    .A1(_1179_),
    .A2(net620));
 sg13g2_a21oi_1 _3089_ (.A1(net369),
    .A2(net616),
    .Y(_1079_),
    .B1(net736));
 sg13g2_o21ai_1 _3090_ (.B1(_1079_),
    .Y(_0246_),
    .A1(_0815_),
    .A2(net616));
 sg13g2_a21oi_1 _3091_ (.A1(_0858_),
    .A2(net619),
    .Y(_1080_),
    .B1(net738));
 sg13g2_o21ai_1 _3092_ (.B1(_1080_),
    .Y(_0247_),
    .A1(_1178_),
    .A2(net619));
 sg13g2_a21oi_1 _3093_ (.A1(_0912_),
    .A2(net619),
    .Y(_1081_),
    .B1(net738));
 sg13g2_o21ai_1 _3094_ (.B1(_1081_),
    .Y(_0248_),
    .A1(_1177_),
    .A2(net619));
 sg13g2_a21oi_1 _3095_ (.A1(_0947_),
    .A2(net619),
    .Y(_1082_),
    .B1(net738));
 sg13g2_o21ai_1 _3096_ (.B1(_1082_),
    .Y(_0249_),
    .A1(_1176_),
    .A2(net619));
 sg13g2_a21oi_1 _3097_ (.A1(net371),
    .A2(net616),
    .Y(_1083_),
    .B1(net736));
 sg13g2_o21ai_1 _3098_ (.B1(_1083_),
    .Y(_0250_),
    .A1(_0988_),
    .A2(net616));
 sg13g2_a21oi_1 _3099_ (.A1(net370),
    .A2(net617),
    .Y(_1084_),
    .B1(net737));
 sg13g2_o21ai_1 _3100_ (.B1(_1084_),
    .Y(_0251_),
    .A1(_0677_),
    .A2(net617));
 sg13g2_a21oi_1 _3101_ (.A1(_0732_),
    .A2(net618),
    .Y(_1085_),
    .B1(net738));
 sg13g2_o21ai_1 _3102_ (.B1(_1085_),
    .Y(_0252_),
    .A1(_1175_),
    .A2(net620));
 sg13g2_a21oi_1 _3103_ (.A1(_0782_),
    .A2(net618),
    .Y(_1086_),
    .B1(net738));
 sg13g2_o21ai_1 _3104_ (.B1(_1086_),
    .Y(_0253_),
    .A1(_1174_),
    .A2(net618));
 sg13g2_a21oi_1 _3105_ (.A1(_0836_),
    .A2(net618),
    .Y(_1087_),
    .B1(net738));
 sg13g2_o21ai_1 _3106_ (.B1(_1087_),
    .Y(_0254_),
    .A1(_1173_),
    .A2(net618));
 sg13g2_a21oi_1 _3107_ (.A1(net375),
    .A2(net616),
    .Y(_1088_),
    .B1(net737));
 sg13g2_o21ai_1 _3108_ (.B1(_1088_),
    .Y(_0255_),
    .A1(_0889_),
    .A2(net616));
 sg13g2_a21oi_1 _3109_ (.A1(_0929_),
    .A2(net618),
    .Y(_1089_),
    .B1(net738));
 sg13g2_o21ai_1 _3110_ (.B1(_1089_),
    .Y(_0256_),
    .A1(_1172_),
    .A2(net618));
 sg13g2_a21oi_1 _3111_ (.A1(_0966_),
    .A2(net619),
    .Y(_1090_),
    .B1(net738));
 sg13g2_o21ai_1 _3112_ (.B1(_1090_),
    .Y(_0257_),
    .A1(_1171_),
    .A2(net618));
 sg13g2_nand2_1 _3113_ (.Y(_1091_),
    .A(_0007_),
    .B(_1308_));
 sg13g2_o21ai_1 _3114_ (.B1(net739),
    .Y(_1092_),
    .A1(net1),
    .A2(net690));
 sg13g2_a21oi_1 _3115_ (.A1(_1170_),
    .A2(net690),
    .Y(_0258_),
    .B1(_1092_));
 sg13g2_o21ai_1 _3116_ (.B1(net739),
    .Y(_1093_),
    .A1(net2),
    .A2(net690));
 sg13g2_a21oi_1 _3117_ (.A1(_1169_),
    .A2(net690),
    .Y(_0259_),
    .B1(_1093_));
 sg13g2_o21ai_1 _3118_ (.B1(net739),
    .Y(_1094_),
    .A1(net3),
    .A2(net690));
 sg13g2_a21oi_1 _3119_ (.A1(_1168_),
    .A2(net690),
    .Y(_0260_),
    .B1(_1094_));
 sg13g2_o21ai_1 _3120_ (.B1(net739),
    .Y(_1095_),
    .A1(net4),
    .A2(net690));
 sg13g2_a21oi_1 _3121_ (.A1(_1167_),
    .A2(net690),
    .Y(_0261_),
    .B1(_1095_));
 sg13g2_o21ai_1 _3122_ (.B1(net742),
    .Y(_1096_),
    .A1(net5),
    .A2(net691));
 sg13g2_a21oi_1 _3123_ (.A1(_1166_),
    .A2(net691),
    .Y(_0262_),
    .B1(_1096_));
 sg13g2_o21ai_1 _3124_ (.B1(net742),
    .Y(_1097_),
    .A1(net6),
    .A2(net691));
 sg13g2_a21oi_1 _3125_ (.A1(_1165_),
    .A2(net691),
    .Y(_0263_),
    .B1(_1097_));
 sg13g2_o21ai_1 _3126_ (.B1(net743),
    .Y(_1098_),
    .A1(net7),
    .A2(net691));
 sg13g2_a21oi_1 _3127_ (.A1(_1164_),
    .A2(net691),
    .Y(_0264_),
    .B1(_1098_));
 sg13g2_o21ai_1 _3128_ (.B1(net742),
    .Y(_1099_),
    .A1(net8),
    .A2(net691));
 sg13g2_a21oi_1 _3129_ (.A1(_1163_),
    .A2(net691),
    .Y(_0265_),
    .B1(_1099_));
 sg13g2_nand3_1 _3130_ (.B(\crp.datapath.aluSrc2SelMux.d3[9] ),
    .C(net608),
    .A(\crp.datapath.aluSrc2SelMux.d3[10] ),
    .Y(_1100_));
 sg13g2_inv_2 _3131_ (.Y(_1101_),
    .A(_1100_));
 sg13g2_nand2_2 _3132_ (.Y(_1102_),
    .A(_1045_),
    .B(_1101_));
 sg13g2_nor2_1 _3133_ (.A(net569),
    .B(net576),
    .Y(_1103_));
 sg13g2_a21oi_1 _3134_ (.A1(_1200_),
    .A2(net576),
    .Y(_0266_),
    .B1(_1103_));
 sg13g2_nor2_1 _3135_ (.A(net565),
    .B(net576),
    .Y(_1104_));
 sg13g2_a21oi_1 _3136_ (.A1(_1212_),
    .A2(net576),
    .Y(_0267_),
    .B1(_1104_));
 sg13g2_mux2_1 _3137_ (.A0(net563),
    .A1(net329),
    .S(net576),
    .X(_0268_));
 sg13g2_mux2_1 _3138_ (.A0(net571),
    .A1(net257),
    .S(net576),
    .X(_0269_));
 sg13g2_mux2_1 _3139_ (.A0(net561),
    .A1(net287),
    .S(_1102_),
    .X(_0270_));
 sg13g2_mux2_1 _3140_ (.A0(net559),
    .A1(net249),
    .S(_1102_),
    .X(_0271_));
 sg13g2_mux2_1 _3141_ (.A0(net567),
    .A1(net314),
    .S(net576),
    .X(_0272_));
 sg13g2_mux2_1 _3142_ (.A0(net557),
    .A1(net278),
    .S(net576),
    .X(_0273_));
 sg13g2_nand3b_1 _3143_ (.B(_0007_),
    .C(_1260_),
    .Y(_1105_),
    .A_N(net703));
 sg13g2_o21ai_1 _3144_ (.B1(net739),
    .Y(_1106_),
    .A1(net1),
    .A2(net688));
 sg13g2_a21oi_1 _3145_ (.A1(_1162_),
    .A2(net688),
    .Y(_0274_),
    .B1(_1106_));
 sg13g2_o21ai_1 _3146_ (.B1(net739),
    .Y(_1107_),
    .A1(net2),
    .A2(net688));
 sg13g2_a21oi_1 _3147_ (.A1(_1160_),
    .A2(net688),
    .Y(_0275_),
    .B1(_1107_));
 sg13g2_o21ai_1 _3148_ (.B1(net739),
    .Y(_1108_),
    .A1(net3),
    .A2(net688));
 sg13g2_a21oi_1 _3149_ (.A1(_1158_),
    .A2(net688),
    .Y(_0276_),
    .B1(_1108_));
 sg13g2_o21ai_1 _3150_ (.B1(net739),
    .Y(_1109_),
    .A1(net4),
    .A2(net688));
 sg13g2_a21oi_1 _3151_ (.A1(_1157_),
    .A2(net688),
    .Y(_0277_),
    .B1(_1109_));
 sg13g2_o21ai_1 _3152_ (.B1(net744),
    .Y(_1110_),
    .A1(net5),
    .A2(net689));
 sg13g2_a21oi_1 _3153_ (.A1(_1156_),
    .A2(net689),
    .Y(_0278_),
    .B1(_1110_));
 sg13g2_o21ai_1 _3154_ (.B1(net744),
    .Y(_1111_),
    .A1(net6),
    .A2(net689));
 sg13g2_a21oi_1 _3155_ (.A1(_1155_),
    .A2(net689),
    .Y(_0279_),
    .B1(_1111_));
 sg13g2_o21ai_1 _3156_ (.B1(net744),
    .Y(_1112_),
    .A1(net7),
    .A2(net689));
 sg13g2_a21oi_1 _3157_ (.A1(_1154_),
    .A2(net689),
    .Y(_0280_),
    .B1(_1112_));
 sg13g2_o21ai_1 _3158_ (.B1(net745),
    .Y(_1113_),
    .A1(net8),
    .A2(net689));
 sg13g2_a21oi_1 _3159_ (.A1(_1153_),
    .A2(net689),
    .Y(_0281_),
    .B1(_1113_));
 sg13g2_nor2_2 _3160_ (.A(net392),
    .B(_1168_),
    .Y(_1114_));
 sg13g2_nand3_1 _3161_ (.B(_1002_),
    .C(_1114_),
    .A(net608),
    .Y(_1115_));
 sg13g2_mux2_1 _3162_ (.A0(net568),
    .A1(net335),
    .S(_1115_),
    .X(_0285_));
 sg13g2_mux2_1 _3163_ (.A0(net564),
    .A1(net349),
    .S(_1115_),
    .X(_0286_));
 sg13g2_mux2_1 _3164_ (.A0(net562),
    .A1(net347),
    .S(_1115_),
    .X(_0287_));
 sg13g2_mux2_1 _3165_ (.A0(net570),
    .A1(net308),
    .S(_1115_),
    .X(_0288_));
 sg13g2_mux2_1 _3166_ (.A0(net560),
    .A1(net270),
    .S(_1115_),
    .X(_0289_));
 sg13g2_mux2_1 _3167_ (.A0(net558),
    .A1(net271),
    .S(_1115_),
    .X(_0290_));
 sg13g2_mux2_1 _3168_ (.A0(net566),
    .A1(net255),
    .S(_1115_),
    .X(_0291_));
 sg13g2_mux2_1 _3169_ (.A0(net556),
    .A1(net316),
    .S(_1115_),
    .X(_0292_));
 sg13g2_nand3_1 _3170_ (.B(_1042_),
    .C(_1114_),
    .A(net608),
    .Y(_1116_));
 sg13g2_mux2_1 _3171_ (.A0(net568),
    .A1(net339),
    .S(net596),
    .X(_0293_));
 sg13g2_mux2_1 _3172_ (.A0(net564),
    .A1(net334),
    .S(net596),
    .X(_0294_));
 sg13g2_nor2_1 _3173_ (.A(net562),
    .B(net596),
    .Y(_1117_));
 sg13g2_a21oi_1 _3174_ (.A1(_1218_),
    .A2(net596),
    .Y(_0295_),
    .B1(_1117_));
 sg13g2_mux2_1 _3175_ (.A0(net570),
    .A1(net229),
    .S(net596),
    .X(_0296_));
 sg13g2_mux2_1 _3176_ (.A0(net560),
    .A1(net267),
    .S(net596),
    .X(_0297_));
 sg13g2_mux2_1 _3177_ (.A0(net558),
    .A1(net293),
    .S(net596),
    .X(_0298_));
 sg13g2_mux2_1 _3178_ (.A0(net566),
    .A1(net268),
    .S(net596),
    .X(_0299_));
 sg13g2_mux2_1 _3179_ (.A0(net556),
    .A1(net279),
    .S(_1116_),
    .X(_0300_));
 sg13g2_nand2_2 _3180_ (.Y(_1118_),
    .A(_1101_),
    .B(_1114_));
 sg13g2_nor2_1 _3181_ (.A(net568),
    .B(net575),
    .Y(_1119_));
 sg13g2_a21oi_1 _3182_ (.A1(_1198_),
    .A2(net575),
    .Y(_0301_),
    .B1(_1119_));
 sg13g2_mux2_1 _3183_ (.A0(net564),
    .A1(net333),
    .S(net575),
    .X(_0302_));
 sg13g2_mux2_1 _3184_ (.A0(net562),
    .A1(net330),
    .S(net575),
    .X(_0303_));
 sg13g2_mux2_1 _3185_ (.A0(net570),
    .A1(net243),
    .S(net575),
    .X(_0304_));
 sg13g2_mux2_1 _3186_ (.A0(net560),
    .A1(net282),
    .S(net575),
    .X(_0305_));
 sg13g2_mux2_1 _3187_ (.A0(net558),
    .A1(net312),
    .S(net575),
    .X(_0306_));
 sg13g2_mux2_1 _3188_ (.A0(net566),
    .A1(net247),
    .S(net575),
    .X(_0307_));
 sg13g2_mux2_1 _3189_ (.A0(net556),
    .A1(net275),
    .S(_1118_),
    .X(_0308_));
 sg13g2_and2_1 _3190_ (.A(net695),
    .B(_1297_),
    .X(_1120_));
 sg13g2_nand2_2 _3191_ (.Y(_1121_),
    .A(net694),
    .B(_1297_));
 sg13g2_nand2b_1 _3192_ (.Y(_1122_),
    .B(_1121_),
    .A_N(_0986_));
 sg13g2_nor2b_1 _3193_ (.A(_0756_),
    .B_N(_0487_),
    .Y(_1123_));
 sg13g2_nand4_1 _3194_ (.B(_0813_),
    .C(_0857_),
    .A(_0710_),
    .Y(_1124_),
    .D(_1123_));
 sg13g2_nor4_1 _3195_ (.A(_0910_),
    .B(_0946_),
    .C(_1122_),
    .D(_1124_),
    .Y(_1125_));
 sg13g2_nand2_1 _3196_ (.Y(_1126_),
    .A(net1),
    .B(_1120_));
 sg13g2_nor2_1 _3197_ (.A(net615),
    .B(_1125_),
    .Y(_1127_));
 sg13g2_a221oi_1 _3198_ (.B2(_1127_),
    .C1(net736),
    .B1(_1126_),
    .A1(_1151_),
    .Y(_0309_),
    .A2(net615));
 sg13g2_nand2_1 _3199_ (.Y(_1128_),
    .A(net368),
    .B(net615));
 sg13g2_a21oi_1 _3200_ (.A1(_1161_),
    .A2(_1120_),
    .Y(_1129_),
    .B1(net615));
 sg13g2_nand2_1 _3201_ (.Y(_1130_),
    .A(_1122_),
    .B(_1129_));
 sg13g2_a21oi_1 _3202_ (.A1(_1128_),
    .A2(_1130_),
    .Y(_0310_),
    .B1(net736));
 sg13g2_nand2_1 _3203_ (.Y(_1131_),
    .A(_0674_),
    .B(_1121_));
 sg13g2_a21oi_1 _3204_ (.A1(_1159_),
    .A2(_1120_),
    .Y(_1132_),
    .B1(net615));
 sg13g2_a22oi_1 _3205_ (.Y(_1133_),
    .B1(_1131_),
    .B2(_1132_),
    .A2(net615),
    .A1(net380));
 sg13g2_nor2_1 _3206_ (.A(net736),
    .B(_1133_),
    .Y(_0311_));
 sg13g2_o21ai_1 _3207_ (.B1(net602),
    .Y(_1134_),
    .A1(_0641_),
    .A2(_0986_));
 sg13g2_a21oi_1 _3208_ (.A1(_0642_),
    .A2(_0986_),
    .Y(_1135_),
    .B1(_1134_));
 sg13g2_a21o_1 _3209_ (.A2(_0986_),
    .A1(_0605_),
    .B1(_0654_),
    .X(_1136_));
 sg13g2_a21oi_1 _3210_ (.A1(_0606_),
    .A2(_0987_),
    .Y(_1137_),
    .B1(_1136_));
 sg13g2_o21ai_1 _3211_ (.B1(_1121_),
    .Y(_1138_),
    .A1(_1135_),
    .A2(_1137_));
 sg13g2_a21oi_1 _3212_ (.A1(net4),
    .A2(_1120_),
    .Y(_1139_),
    .B1(net615));
 sg13g2_a221oi_1 _3213_ (.B2(_1139_),
    .C1(net736),
    .B1(_1138_),
    .A1(_1150_),
    .Y(_0312_),
    .A2(net615));
 sg13g2_nand3_1 _3214_ (.B(_1039_),
    .C(_1045_),
    .A(net608),
    .Y(_1140_));
 sg13g2_nor2_1 _3215_ (.A(net569),
    .B(net595),
    .Y(_1141_));
 sg13g2_a21oi_1 _3216_ (.A1(_1199_),
    .A2(net595),
    .Y(_0313_),
    .B1(_1141_));
 sg13g2_mux2_1 _3217_ (.A0(net565),
    .A1(net355),
    .S(net595),
    .X(_0314_));
 sg13g2_mux2_1 _3218_ (.A0(net563),
    .A1(net318),
    .S(net595),
    .X(_0315_));
 sg13g2_mux2_1 _3219_ (.A0(net571),
    .A1(net317),
    .S(net595),
    .X(_0316_));
 sg13g2_mux2_1 _3220_ (.A0(net561),
    .A1(net273),
    .S(_1140_),
    .X(_0317_));
 sg13g2_mux2_1 _3221_ (.A0(net559),
    .A1(net245),
    .S(net595),
    .X(_0318_));
 sg13g2_mux2_1 _3222_ (.A0(net567),
    .A1(net236),
    .S(net595),
    .X(_0319_));
 sg13g2_mux2_1 _3223_ (.A0(net557),
    .A1(net298),
    .S(net595),
    .X(_0320_));
 sg13g2_nand3_1 _3224_ (.B(_1168_),
    .C(_1101_),
    .A(_1167_),
    .Y(_1142_));
 sg13g2_nor2_1 _3225_ (.A(net568),
    .B(_1142_),
    .Y(_1143_));
 sg13g2_a21oi_1 _3226_ (.A1(_1193_),
    .A2(_1142_),
    .Y(_0321_),
    .B1(_1143_));
 sg13g2_nor2_1 _3227_ (.A(net564),
    .B(net574),
    .Y(_1144_));
 sg13g2_a21oi_1 _3228_ (.A1(_1209_),
    .A2(net574),
    .Y(_0322_),
    .B1(_1144_));
 sg13g2_mux2_1 _3229_ (.A0(net562),
    .A1(net324),
    .S(net574),
    .X(_0323_));
 sg13g2_mux2_1 _3230_ (.A0(net570),
    .A1(net237),
    .S(net574),
    .X(_0324_));
 sg13g2_mux2_1 _3231_ (.A0(net560),
    .A1(net311),
    .S(net574),
    .X(_0325_));
 sg13g2_mux2_1 _3232_ (.A0(net558),
    .A1(net315),
    .S(net574),
    .X(_0326_));
 sg13g2_mux2_1 _3233_ (.A0(net566),
    .A1(net288),
    .S(net574),
    .X(_0327_));
 sg13g2_mux2_1 _3234_ (.A0(net556),
    .A1(net285),
    .S(net574),
    .X(_0328_));
 sg13g2_nand3_1 _3235_ (.B(_1042_),
    .C(_1045_),
    .A(_1001_),
    .Y(_1145_));
 sg13g2_mux2_1 _3236_ (.A0(net569),
    .A1(net343),
    .S(net594),
    .X(_0329_));
 sg13g2_mux2_1 _3237_ (.A0(net565),
    .A1(net356),
    .S(net594),
    .X(_0330_));
 sg13g2_nor2_1 _3238_ (.A(net563),
    .B(net594),
    .Y(_1146_));
 sg13g2_a21oi_1 _3239_ (.A1(_1219_),
    .A2(net594),
    .Y(_0331_),
    .B1(_1146_));
 sg13g2_mux2_1 _3240_ (.A0(net571),
    .A1(net297),
    .S(net594),
    .X(_0332_));
 sg13g2_mux2_1 _3241_ (.A0(net561),
    .A1(net291),
    .S(_1145_),
    .X(_0333_));
 sg13g2_mux2_1 _3242_ (.A0(net559),
    .A1(net266),
    .S(net594),
    .X(_0334_));
 sg13g2_mux2_1 _3243_ (.A0(net567),
    .A1(net300),
    .S(net594),
    .X(_0335_));
 sg13g2_mux2_1 _3244_ (.A0(net557),
    .A1(net265),
    .S(net594),
    .X(_0336_));
 sg13g2_nand3_1 _3245_ (.B(_1039_),
    .C(_1114_),
    .A(net608),
    .Y(_1147_));
 sg13g2_nor2_1 _3246_ (.A(net568),
    .B(net593),
    .Y(_1148_));
 sg13g2_a21oi_1 _3247_ (.A1(_1197_),
    .A2(net593),
    .Y(_0337_),
    .B1(_1148_));
 sg13g2_nor2_1 _3248_ (.A(net564),
    .B(_1147_),
    .Y(_1149_));
 sg13g2_a21oi_1 _3249_ (.A1(_1211_),
    .A2(net593),
    .Y(_0338_),
    .B1(_1149_));
 sg13g2_mux2_1 _3250_ (.A0(net562),
    .A1(net309),
    .S(net593),
    .X(_0339_));
 sg13g2_mux2_1 _3251_ (.A0(net570),
    .A1(net244),
    .S(net593),
    .X(_0340_));
 sg13g2_mux2_1 _3252_ (.A0(net560),
    .A1(net284),
    .S(net593),
    .X(_0341_));
 sg13g2_mux2_1 _3253_ (.A0(net558),
    .A1(net304),
    .S(net593),
    .X(_0342_));
 sg13g2_mux2_1 _3254_ (.A0(net566),
    .A1(net259),
    .S(net593),
    .X(_0343_));
 sg13g2_mux2_1 _3255_ (.A0(net556),
    .A1(net292),
    .S(_1147_),
    .X(_0344_));
 sg13g2_inv_1 _3257__3 (.Y(net208),
    .A(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbp_1 _3258_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net11),
    .D(_0156_),
    .Q_N(_0009_),
    .Q(\crp.datapath.registerFile.regs[0][0] ));
 sg13g2_dfrbp_1 _3259_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net121),
    .D(_0157_),
    .Q_N(_0034_),
    .Q(\crp.datapath.registerFile.regs[0][1] ));
 sg13g2_dfrbp_1 _3260_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net120),
    .D(_0158_),
    .Q_N(_0051_),
    .Q(\crp.datapath.registerFile.regs[0][2] ));
 sg13g2_dfrbp_1 _3261_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net119),
    .D(_0159_),
    .Q_N(_0068_),
    .Q(\crp.datapath.registerFile.regs[0][3] ));
 sg13g2_dfrbp_1 _3262_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net118),
    .D(_0160_),
    .Q_N(_0085_),
    .Q(\crp.datapath.registerFile.regs[0][4] ));
 sg13g2_dfrbp_1 _3263_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net117),
    .D(_0161_),
    .Q_N(_0102_),
    .Q(\crp.datapath.registerFile.regs[0][5] ));
 sg13g2_dfrbp_1 _3264_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net116),
    .D(_0162_),
    .Q_N(_0119_),
    .Q(\crp.datapath.registerFile.regs[0][6] ));
 sg13g2_dfrbp_1 _3265_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net115),
    .D(_0163_),
    .Q_N(_0136_),
    .Q(\crp.datapath.registerFile.regs[0][7] ));
 sg13g2_dfrbp_1 _3266_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net114),
    .D(_0164_),
    .Q_N(_0013_),
    .Q(\crp.datapath.registerFile.regs[2][0] ));
 sg13g2_dfrbp_1 _3267_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net113),
    .D(_0165_),
    .Q_N(_0036_),
    .Q(\crp.datapath.registerFile.regs[2][1] ));
 sg13g2_dfrbp_1 _3268_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net112),
    .D(_0166_),
    .Q_N(_0053_),
    .Q(\crp.datapath.registerFile.regs[2][2] ));
 sg13g2_dfrbp_1 _3269_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net111),
    .D(_0167_),
    .Q_N(_0070_),
    .Q(\crp.datapath.registerFile.regs[2][3] ));
 sg13g2_dfrbp_1 _3270_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net110),
    .D(_0168_),
    .Q_N(_0087_),
    .Q(\crp.datapath.registerFile.regs[2][4] ));
 sg13g2_dfrbp_1 _3271_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net109),
    .D(_0169_),
    .Q_N(_0104_),
    .Q(\crp.datapath.registerFile.regs[2][5] ));
 sg13g2_dfrbp_1 _3272_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net108),
    .D(_0170_),
    .Q_N(_0121_),
    .Q(\crp.datapath.registerFile.regs[2][6] ));
 sg13g2_dfrbp_1 _3273_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net107),
    .D(_0171_),
    .Q_N(_0138_),
    .Q(\crp.datapath.registerFile.regs[2][7] ));
 sg13g2_dfrbp_1 _3274_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net106),
    .D(_0172_),
    .Q_N(_0010_),
    .Q(\crp.datapath.registerFile.regs[1][0] ));
 sg13g2_dfrbp_1 _3275_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net105),
    .D(_0173_),
    .Q_N(_0035_),
    .Q(\crp.datapath.registerFile.regs[1][1] ));
 sg13g2_dfrbp_1 _3276_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net104),
    .D(_0174_),
    .Q_N(_0052_),
    .Q(\crp.datapath.registerFile.regs[1][2] ));
 sg13g2_dfrbp_1 _3277_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net103),
    .D(_0175_),
    .Q_N(_0069_),
    .Q(\crp.datapath.registerFile.regs[1][3] ));
 sg13g2_dfrbp_1 _3278_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net102),
    .D(_0176_),
    .Q_N(_0086_),
    .Q(\crp.datapath.registerFile.regs[1][4] ));
 sg13g2_dfrbp_1 _3279_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net101),
    .D(_0177_),
    .Q_N(_0103_),
    .Q(\crp.datapath.registerFile.regs[1][5] ));
 sg13g2_dfrbp_1 _3280_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net100),
    .D(_0178_),
    .Q_N(_0120_),
    .Q(\crp.datapath.registerFile.regs[1][6] ));
 sg13g2_dfrbp_1 _3281_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net99),
    .D(_0179_),
    .Q_N(_0137_),
    .Q(\crp.datapath.registerFile.regs[1][7] ));
 sg13g2_dfrbp_1 _3282_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net98),
    .D(_0180_),
    .Q_N(_0021_),
    .Q(\crp.datapath.registerFile.regs[8][0] ));
 sg13g2_dfrbp_1 _3283_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net97),
    .D(_0181_),
    .Q_N(_0042_),
    .Q(\crp.datapath.registerFile.regs[8][1] ));
 sg13g2_dfrbp_1 _3284_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net96),
    .D(_0182_),
    .Q_N(_0059_),
    .Q(\crp.datapath.registerFile.regs[8][2] ));
 sg13g2_dfrbp_1 _3285_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net95),
    .D(_0183_),
    .Q_N(_0076_),
    .Q(\crp.datapath.registerFile.regs[8][3] ));
 sg13g2_dfrbp_1 _3286_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net94),
    .D(_0184_),
    .Q_N(_0093_),
    .Q(\crp.datapath.registerFile.regs[8][4] ));
 sg13g2_dfrbp_1 _3287_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net93),
    .D(_0185_),
    .Q_N(_0110_),
    .Q(\crp.datapath.registerFile.regs[8][5] ));
 sg13g2_dfrbp_1 _3288_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net92),
    .D(_0186_),
    .Q_N(_0127_),
    .Q(\crp.datapath.registerFile.regs[8][6] ));
 sg13g2_dfrbp_1 _3289_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net91),
    .D(_0187_),
    .Q_N(_0144_),
    .Q(\crp.datapath.registerFile.regs[8][7] ));
 sg13g2_dfrbp_1 _3290_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net90),
    .D(_0188_),
    .Q_N(_0028_),
    .Q(\crp.datapath.registerFile.regs[15][0] ));
 sg13g2_dfrbp_1 _3291_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net89),
    .D(_0189_),
    .Q_N(_0049_),
    .Q(\crp.datapath.registerFile.regs[15][1] ));
 sg13g2_dfrbp_1 _3292_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net88),
    .D(_0190_),
    .Q_N(_0066_),
    .Q(\crp.datapath.registerFile.regs[15][2] ));
 sg13g2_dfrbp_1 _3293_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net87),
    .D(_0191_),
    .Q_N(_0083_),
    .Q(\crp.datapath.registerFile.regs[15][3] ));
 sg13g2_dfrbp_1 _3294_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net86),
    .D(_0192_),
    .Q_N(_0100_),
    .Q(\crp.datapath.registerFile.regs[15][4] ));
 sg13g2_dfrbp_1 _3295_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net85),
    .D(_0193_),
    .Q_N(_0117_),
    .Q(\crp.datapath.registerFile.regs[15][5] ));
 sg13g2_dfrbp_1 _3296_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net84),
    .D(_0194_),
    .Q_N(_0134_),
    .Q(\crp.datapath.registerFile.regs[15][6] ));
 sg13g2_dfrbp_1 _3297_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net83),
    .D(net296),
    .Q_N(_0151_),
    .Q(\crp.datapath.registerFile.regs[15][7] ));
 sg13g2_dfrbp_1 _3298_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net82),
    .D(_0196_),
    .Q_N(_0027_),
    .Q(\crp.datapath.registerFile.regs[14][0] ));
 sg13g2_dfrbp_1 _3299_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net81),
    .D(_0197_),
    .Q_N(_0048_),
    .Q(\crp.datapath.registerFile.regs[14][1] ));
 sg13g2_dfrbp_1 _3300_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net80),
    .D(_0198_),
    .Q_N(_0065_),
    .Q(\crp.datapath.registerFile.regs[14][2] ));
 sg13g2_dfrbp_1 _3301_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net79),
    .D(_0199_),
    .Q_N(_0082_),
    .Q(\crp.datapath.registerFile.regs[14][3] ));
 sg13g2_dfrbp_1 _3302_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net78),
    .D(_0200_),
    .Q_N(_0099_),
    .Q(\crp.datapath.registerFile.regs[14][4] ));
 sg13g2_dfrbp_1 _3303_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net77),
    .D(_0201_),
    .Q_N(_0116_),
    .Q(\crp.datapath.registerFile.regs[14][5] ));
 sg13g2_dfrbp_1 _3304_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net76),
    .D(_0202_),
    .Q_N(_0133_),
    .Q(\crp.datapath.registerFile.regs[14][6] ));
 sg13g2_dfrbp_1 _3305_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net75),
    .D(_0203_),
    .Q_N(_0150_),
    .Q(\crp.datapath.registerFile.regs[14][7] ));
 sg13g2_dfrbp_1 _3306_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net74),
    .D(_0204_),
    .Q_N(_1620_),
    .Q(\crp.datapath.memReadData[0] ));
 sg13g2_dfrbp_1 _3307_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net73),
    .D(_0205_),
    .Q_N(_1619_),
    .Q(\crp.datapath.memReadData[1] ));
 sg13g2_dfrbp_1 _3308_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net72),
    .D(_0206_),
    .Q_N(_1618_),
    .Q(\crp.datapath.memReadData[2] ));
 sg13g2_dfrbp_1 _3309_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net71),
    .D(_0207_),
    .Q_N(_1617_),
    .Q(\crp.datapath.memReadData[3] ));
 sg13g2_dfrbp_1 _3310_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net70),
    .D(_0208_),
    .Q_N(_1616_),
    .Q(\crp.datapath.memReadData[4] ));
 sg13g2_dfrbp_1 _3311_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net69),
    .D(_0209_),
    .Q_N(_1615_),
    .Q(\crp.datapath.memReadData[5] ));
 sg13g2_dfrbp_1 _3312_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net68),
    .D(_0210_),
    .Q_N(_1614_),
    .Q(\crp.datapath.memReadData[6] ));
 sg13g2_dfrbp_1 _3313_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net67),
    .D(_0211_),
    .Q_N(_1613_),
    .Q(\crp.datapath.memReadData[7] ));
 sg13g2_dfrbp_1 _3314_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net66),
    .D(_0212_),
    .Q_N(_0026_),
    .Q(\crp.datapath.registerFile.regs[13][0] ));
 sg13g2_dfrbp_1 _3315_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net65),
    .D(_0213_),
    .Q_N(_0047_),
    .Q(\crp.datapath.registerFile.regs[13][1] ));
 sg13g2_dfrbp_1 _3316_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net64),
    .D(_0214_),
    .Q_N(_0064_),
    .Q(\crp.datapath.registerFile.regs[13][2] ));
 sg13g2_dfrbp_1 _3317_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net63),
    .D(_0215_),
    .Q_N(_0081_),
    .Q(\crp.datapath.registerFile.regs[13][3] ));
 sg13g2_dfrbp_1 _3318_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net62),
    .D(_0216_),
    .Q_N(_0098_),
    .Q(\crp.datapath.registerFile.regs[13][4] ));
 sg13g2_dfrbp_1 _3319_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net61),
    .D(_0217_),
    .Q_N(_0115_),
    .Q(\crp.datapath.registerFile.regs[13][5] ));
 sg13g2_dfrbp_1 _3320_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net60),
    .D(_0218_),
    .Q_N(_0132_),
    .Q(\crp.datapath.registerFile.regs[13][6] ));
 sg13g2_dfrbp_1 _3321_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net59),
    .D(_0219_),
    .Q_N(_0149_),
    .Q(\crp.datapath.registerFile.regs[13][7] ));
 sg13g2_dfrbp_1 _3322_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net58),
    .D(_0220_),
    .Q_N(_0008_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[0] ));
 sg13g2_dfrbp_1 _3323_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net56),
    .D(_0221_),
    .Q_N(_0033_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[1] ));
 sg13g2_dfrbp_1 _3324_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net54),
    .D(_0222_),
    .Q_N(_0050_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[2] ));
 sg13g2_dfrbp_1 _3325_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net52),
    .D(_0223_),
    .Q_N(_0067_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[3] ));
 sg13g2_dfrbp_1 _3326_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net50),
    .D(_0224_),
    .Q_N(_0084_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[4] ));
 sg13g2_dfrbp_1 _3327_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net48),
    .D(_0225_),
    .Q_N(_0101_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[5] ));
 sg13g2_dfrbp_1 _3328_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net46),
    .D(_0226_),
    .Q_N(_0118_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[6] ));
 sg13g2_dfrbp_1 _3329_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net44),
    .D(_0227_),
    .Q_N(_0135_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[7] ));
 sg13g2_dfrbp_1 _3330_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net42),
    .D(_0228_),
    .Q_N(_0000_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[8] ));
 sg13g2_dfrbp_1 _3331_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net40),
    .D(_0229_),
    .Q_N(_0001_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[9] ));
 sg13g2_dfrbp_1 _3332_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net38),
    .D(_0230_),
    .Q_N(_0002_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[10] ));
 sg13g2_dfrbp_1 _3333_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net36),
    .D(_0231_),
    .Q_N(_0003_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[11] ));
 sg13g2_dfrbp_1 _3334_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net34),
    .D(_0232_),
    .Q_N(_0004_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[12] ));
 sg13g2_dfrbp_1 _3335_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net32),
    .D(_0233_),
    .Q_N(_0005_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[13] ));
 sg13g2_dfrbp_1 _3336_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net30),
    .D(_0234_),
    .Q_N(_0006_),
    .Q(\crp.datapath.aluSrc1SelMux.d0[14] ));
 sg13g2_dfrbp_1 _3337_ (.CLK(clknet_5_23__leaf_clk_regs),
    .RESET_B(net28),
    .D(_0235_),
    .Q_N(_0025_),
    .Q(\crp.datapath.registerFile.regs[12][0] ));
 sg13g2_dfrbp_1 _3338_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net27),
    .D(_0236_),
    .Q_N(_0046_),
    .Q(\crp.datapath.registerFile.regs[12][1] ));
 sg13g2_dfrbp_1 _3339_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net26),
    .D(_0237_),
    .Q_N(_0063_),
    .Q(\crp.datapath.registerFile.regs[12][2] ));
 sg13g2_dfrbp_1 _3340_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net25),
    .D(_0238_),
    .Q_N(_0080_),
    .Q(\crp.datapath.registerFile.regs[12][3] ));
 sg13g2_dfrbp_1 _3341_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net24),
    .D(_0239_),
    .Q_N(_0097_),
    .Q(\crp.datapath.registerFile.regs[12][4] ));
 sg13g2_dfrbp_1 _3342_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net23),
    .D(_0240_),
    .Q_N(_0114_),
    .Q(\crp.datapath.registerFile.regs[12][5] ));
 sg13g2_dfrbp_1 _3343_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net22),
    .D(_0241_),
    .Q_N(_0131_),
    .Q(\crp.datapath.registerFile.regs[12][6] ));
 sg13g2_dfrbp_1 _3344_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net21),
    .D(_0242_),
    .Q_N(_0148_),
    .Q(\crp.datapath.registerFile.regs[12][7] ));
 sg13g2_dfrbp_1 _3345_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net20),
    .D(_0243_),
    .Q_N(_1612_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[0] ));
 sg13g2_dfrbp_1 _3346_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net18),
    .D(_0244_),
    .Q_N(_1611_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[1] ));
 sg13g2_dfrbp_1 _3347_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net16),
    .D(_0245_),
    .Q_N(_1610_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[2] ));
 sg13g2_dfrbp_1 _3348_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net14),
    .D(_0246_),
    .Q_N(_1609_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[3] ));
 sg13g2_dfrbp_1 _3349_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net12),
    .D(_0247_),
    .Q_N(_1608_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[4] ));
 sg13g2_dfrbp_1 _3350_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net10),
    .D(_0248_),
    .Q_N(_1607_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[5] ));
 sg13g2_dfrbp_1 _3351_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net197),
    .D(_0249_),
    .Q_N(_1606_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[6] ));
 sg13g2_dfrbp_1 _3352_ (.CLK(clknet_5_25__leaf_clk_regs),
    .RESET_B(net195),
    .D(_0250_),
    .Q_N(_1605_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[7] ));
 sg13g2_dfrbp_1 _3353_ (.CLK(clknet_5_31__leaf_clk_regs),
    .RESET_B(net193),
    .D(_0251_),
    .Q_N(_1604_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[8] ));
 sg13g2_dfrbp_1 _3354_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net191),
    .D(_0252_),
    .Q_N(_1603_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[9] ));
 sg13g2_dfrbp_1 _3355_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net189),
    .D(_0253_),
    .Q_N(_1602_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[10] ));
 sg13g2_dfrbp_1 _3356_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net187),
    .D(_0254_),
    .Q_N(_1601_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[11] ));
 sg13g2_dfrbp_1 _3357_ (.CLK(clknet_5_29__leaf_clk_regs),
    .RESET_B(net185),
    .D(_0255_),
    .Q_N(_1600_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[12] ));
 sg13g2_dfrbp_1 _3358_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net183),
    .D(_0256_),
    .Q_N(_1599_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[13] ));
 sg13g2_dfrbp_1 _3359_ (.CLK(clknet_5_28__leaf_clk_regs),
    .RESET_B(net181),
    .D(_0257_),
    .Q_N(_1598_),
    .Q(\crp.datapath.aluSrc1SelMux.d1[14] ));
 sg13g2_dfrbp_1 _3360_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net179),
    .D(_0258_),
    .Q_N(_0011_),
    .Q(\crp.datapath.aluSrc2SelMux.d3[9] ));
 sg13g2_dfrbp_1 _3361_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net177),
    .D(_0259_),
    .Q_N(_0012_),
    .Q(\crp.datapath.aluSrc2SelMux.d3[10] ));
 sg13g2_dfrbp_1 _3362_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net175),
    .D(_0260_),
    .Q_N(_0015_),
    .Q(\crp.datapath.aluSrc2SelMux.d3[11] ));
 sg13g2_dfrbp_1 _3363_ (.CLK(clknet_5_24__leaf_clk_regs),
    .RESET_B(net173),
    .D(_0261_),
    .Q_N(_0020_),
    .Q(\crp.datapath.aluSrc2SelMux.d3[12] ));
 sg13g2_dfrbp_1 _3364_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net171),
    .D(_0262_),
    .Q_N(_1597_),
    .Q(\crp.controller.aluDec.opcode[0] ));
 sg13g2_dfrbp_1 _3365_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net169),
    .D(_0263_),
    .Q_N(_1596_),
    .Q(\crp.controller.aluDec.opcode[1] ));
 sg13g2_dfrbp_1 _3366_ (.CLK(clknet_5_27__leaf_clk_regs),
    .RESET_B(net167),
    .D(_0264_),
    .Q_N(_1595_),
    .Q(\crp.controller.aluDec.opcode[2] ));
 sg13g2_dfrbp_1 _3367_ (.CLK(clknet_5_30__leaf_clk_regs),
    .RESET_B(net165),
    .D(_0265_),
    .Q_N(_1594_),
    .Q(\crp.controller.aluDec.opcode[3] ));
 sg13g2_dfrbp_1 _3368_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net163),
    .D(_0266_),
    .Q_N(_0024_),
    .Q(\crp.datapath.registerFile.regs[11][0] ));
 sg13g2_dfrbp_1 _3369_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net162),
    .D(_0267_),
    .Q_N(_0045_),
    .Q(\crp.datapath.registerFile.regs[11][1] ));
 sg13g2_dfrbp_1 _3370_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net161),
    .D(_0268_),
    .Q_N(_0062_),
    .Q(\crp.datapath.registerFile.regs[11][2] ));
 sg13g2_dfrbp_1 _3371_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net160),
    .D(_0269_),
    .Q_N(_0079_),
    .Q(\crp.datapath.registerFile.regs[11][3] ));
 sg13g2_dfrbp_1 _3372_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net159),
    .D(_0270_),
    .Q_N(_0096_),
    .Q(\crp.datapath.registerFile.regs[11][4] ));
 sg13g2_dfrbp_1 _3373_ (.CLK(clknet_5_21__leaf_clk_regs),
    .RESET_B(net158),
    .D(_0271_),
    .Q_N(_0113_),
    .Q(\crp.datapath.registerFile.regs[11][5] ));
 sg13g2_dfrbp_1 _3374_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net157),
    .D(_0272_),
    .Q_N(_0130_),
    .Q(\crp.datapath.registerFile.regs[11][6] ));
 sg13g2_dfrbp_1 _3375_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net156),
    .D(_0273_),
    .Q_N(_0147_),
    .Q(\crp.datapath.registerFile.regs[11][7] ));
 sg13g2_dfrbp_1 _3376_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net155),
    .D(_0274_),
    .Q_N(_1593_),
    .Q(\crp.controller.aluDec.aluRtypeDec.func[0] ));
 sg13g2_dfrbp_1 _3377_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net153),
    .D(_0275_),
    .Q_N(_1592_),
    .Q(\crp.controller.aluDec.aluRtypeDec.func[1] ));
 sg13g2_dfrbp_1 _3378_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net151),
    .D(_0276_),
    .Q_N(_1591_),
    .Q(\crp.controller.aluDec.aluRtypeDec.func[2] ));
 sg13g2_dfrbp_1 _3379_ (.CLK(clknet_5_14__leaf_clk_regs),
    .RESET_B(net149),
    .D(_0277_),
    .Q_N(_1590_),
    .Q(\crp.controller.aluDec.aluRtypeDec.func[3] ));
 sg13g2_dfrbp_1 _3380_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net147),
    .D(_0278_),
    .Q_N(_0029_),
    .Q(\crp.datapath.aluSrc2SelMux.d2[4] ));
 sg13g2_dfrbp_1 _3381_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net145),
    .D(_0279_),
    .Q_N(_0030_),
    .Q(\crp.datapath.aluSrc2SelMux.d2[5] ));
 sg13g2_dfrbp_1 _3382_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net143),
    .D(_0280_),
    .Q_N(_0031_),
    .Q(\crp.datapath.aluSrc2SelMux.d2[6] ));
 sg13g2_dfrbp_1 _3383_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net141),
    .D(_0281_),
    .Q_N(_0032_),
    .Q(\crp.datapath.aluSrc2SelMux.d2[7] ));
 sg13g2_dfrbp_1 _3384_ (.CLK(net206),
    .RESET_B(net139),
    .D(_0282_),
    .Q_N(_0152_),
    .Q(\crp.controller.aluDec.aluRtypeDec.state[0] ));
 sg13g2_dfrbp_1 _3385_ (.CLK(net207),
    .RESET_B(net137),
    .D(_0283_),
    .Q_N(_1589_),
    .Q(\crp.controller.aluDec.aluRtypeDec.state[1] ));
 sg13g2_dfrbp_1 _3386_ (.CLK(net208),
    .RESET_B(net135),
    .D(_0284_),
    .Q_N(_0007_),
    .Q(\crp.controller.aluDec.aluRtypeDec.state[2] ));
 sg13g2_dfrbp_1 _3387_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net133),
    .D(_0285_),
    .Q_N(_0016_),
    .Q(\crp.datapath.registerFile.regs[4][0] ));
 sg13g2_dfrbp_1 _3388_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net132),
    .D(_0286_),
    .Q_N(_0038_),
    .Q(\crp.datapath.registerFile.regs[4][1] ));
 sg13g2_dfrbp_1 _3389_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net131),
    .D(_0287_),
    .Q_N(_0055_),
    .Q(\crp.datapath.registerFile.regs[4][2] ));
 sg13g2_dfrbp_1 _3390_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net130),
    .D(_0288_),
    .Q_N(_0072_),
    .Q(\crp.datapath.registerFile.regs[4][3] ));
 sg13g2_dfrbp_1 _3391_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net129),
    .D(_0289_),
    .Q_N(_0089_),
    .Q(\crp.datapath.registerFile.regs[4][4] ));
 sg13g2_dfrbp_1 _3392_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net128),
    .D(_0290_),
    .Q_N(_0106_),
    .Q(\crp.datapath.registerFile.regs[4][5] ));
 sg13g2_dfrbp_1 _3393_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net127),
    .D(_0291_),
    .Q_N(_0123_),
    .Q(\crp.datapath.registerFile.regs[4][6] ));
 sg13g2_dfrbp_1 _3394_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net126),
    .D(_0292_),
    .Q_N(_0140_),
    .Q(\crp.datapath.registerFile.regs[4][7] ));
 sg13g2_dfrbp_1 _3395_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net125),
    .D(_0293_),
    .Q_N(_0017_),
    .Q(\crp.datapath.registerFile.regs[5][0] ));
 sg13g2_dfrbp_1 _3396_ (.CLK(clknet_5_13__leaf_clk_regs),
    .RESET_B(net124),
    .D(_0294_),
    .Q_N(_0039_),
    .Q(\crp.datapath.registerFile.regs[5][1] ));
 sg13g2_dfrbp_1 _3397_ (.CLK(clknet_5_8__leaf_clk_regs),
    .RESET_B(net123),
    .D(_0295_),
    .Q_N(_0056_),
    .Q(\crp.datapath.registerFile.regs[5][2] ));
 sg13g2_dfrbp_1 _3398_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net122),
    .D(_0296_),
    .Q_N(_0073_),
    .Q(\crp.datapath.registerFile.regs[5][3] ));
 sg13g2_dfrbp_1 _3399_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net57),
    .D(_0297_),
    .Q_N(_0090_),
    .Q(\crp.datapath.registerFile.regs[5][4] ));
 sg13g2_dfrbp_1 _3400_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net55),
    .D(_0298_),
    .Q_N(_0107_),
    .Q(\crp.datapath.registerFile.regs[5][5] ));
 sg13g2_dfrbp_1 _3401_ (.CLK(clknet_5_2__leaf_clk_regs),
    .RESET_B(net53),
    .D(_0299_),
    .Q_N(_0124_),
    .Q(\crp.datapath.registerFile.regs[5][6] ));
 sg13g2_dfrbp_1 _3402_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net51),
    .D(_0300_),
    .Q_N(_0141_),
    .Q(\crp.datapath.registerFile.regs[5][7] ));
 sg13g2_dfrbp_1 _3403_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net49),
    .D(_0301_),
    .Q_N(_0019_),
    .Q(\crp.datapath.registerFile.regs[7][0] ));
 sg13g2_dfrbp_1 _3404_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net47),
    .D(_0302_),
    .Q_N(_0041_),
    .Q(\crp.datapath.registerFile.regs[7][1] ));
 sg13g2_dfrbp_1 _3405_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net45),
    .D(_0303_),
    .Q_N(_0058_),
    .Q(\crp.datapath.registerFile.regs[7][2] ));
 sg13g2_dfrbp_1 _3406_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net43),
    .D(_0304_),
    .Q_N(_0075_),
    .Q(\crp.datapath.registerFile.regs[7][3] ));
 sg13g2_dfrbp_1 _3407_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net41),
    .D(_0305_),
    .Q_N(_0092_),
    .Q(\crp.datapath.registerFile.regs[7][4] ));
 sg13g2_dfrbp_1 _3408_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net39),
    .D(_0306_),
    .Q_N(_0109_),
    .Q(\crp.datapath.registerFile.regs[7][5] ));
 sg13g2_dfrbp_1 _3409_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net37),
    .D(_0307_),
    .Q_N(_0126_),
    .Q(\crp.datapath.registerFile.regs[7][6] ));
 sg13g2_dfrbp_1 _3410_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net35),
    .D(_0308_),
    .Q_N(_0143_),
    .Q(\crp.datapath.registerFile.regs[7][7] ));
 sg13g2_dfrbp_1 _3411_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net33),
    .D(_0309_),
    .Q_N(_1588_),
    .Q(\crp.controller.flags[0] ));
 sg13g2_dfrbp_1 _3412_ (.CLK(clknet_5_15__leaf_clk_regs),
    .RESET_B(net29),
    .D(_0310_),
    .Q_N(_1587_),
    .Q(\crp.controller.flags[1] ));
 sg13g2_dfrbp_1 _3413_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net17),
    .D(_0311_),
    .Q_N(_1586_),
    .Q(\crp.controller.flags[2] ));
 sg13g2_dfrbp_1 _3414_ (.CLK(clknet_5_26__leaf_clk_regs),
    .RESET_B(net13),
    .D(_0312_),
    .Q_N(_1585_),
    .Q(\crp.controller.flags[3] ));
 sg13g2_dfrbp_1 _3415_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net9),
    .D(_0313_),
    .Q_N(_0023_),
    .Q(\crp.datapath.registerFile.regs[10][0] ));
 sg13g2_dfrbp_1 _3416_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net196),
    .D(_0314_),
    .Q_N(_0044_),
    .Q(\crp.datapath.registerFile.regs[10][1] ));
 sg13g2_dfrbp_1 _3417_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net194),
    .D(_0315_),
    .Q_N(_0061_),
    .Q(\crp.datapath.registerFile.regs[10][2] ));
 sg13g2_dfrbp_1 _3418_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net192),
    .D(_0316_),
    .Q_N(_0078_),
    .Q(\crp.datapath.registerFile.regs[10][3] ));
 sg13g2_dfrbp_1 _3419_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net190),
    .D(_0317_),
    .Q_N(_0095_),
    .Q(\crp.datapath.registerFile.regs[10][4] ));
 sg13g2_dfrbp_1 _3420_ (.CLK(clknet_5_20__leaf_clk_regs),
    .RESET_B(net188),
    .D(_0318_),
    .Q_N(_0112_),
    .Q(\crp.datapath.registerFile.regs[10][5] ));
 sg13g2_dfrbp_1 _3421_ (.CLK(clknet_5_16__leaf_clk_regs),
    .RESET_B(net186),
    .D(_0319_),
    .Q_N(_0129_),
    .Q(\crp.datapath.registerFile.regs[10][6] ));
 sg13g2_dfrbp_1 _3422_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net184),
    .D(_0320_),
    .Q_N(_0146_),
    .Q(\crp.datapath.registerFile.regs[10][7] ));
 sg13g2_dfrbp_1 _3423_ (.CLK(clknet_5_11__leaf_clk_regs),
    .RESET_B(net182),
    .D(net225),
    .Q_N(_0014_),
    .Q(\crp.datapath.registerFile.regs[3][0] ));
 sg13g2_dfrbp_1 _3424_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net180),
    .D(_0322_),
    .Q_N(_0037_),
    .Q(\crp.datapath.registerFile.regs[3][1] ));
 sg13g2_dfrbp_1 _3425_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net178),
    .D(_0323_),
    .Q_N(_0054_),
    .Q(\crp.datapath.registerFile.regs[3][2] ));
 sg13g2_dfrbp_1 _3426_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net176),
    .D(_0324_),
    .Q_N(_0071_),
    .Q(\crp.datapath.registerFile.regs[3][3] ));
 sg13g2_dfrbp_1 _3427_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net174),
    .D(_0325_),
    .Q_N(_0088_),
    .Q(\crp.datapath.registerFile.regs[3][4] ));
 sg13g2_dfrbp_1 _3428_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net172),
    .D(_0326_),
    .Q_N(_0105_),
    .Q(\crp.datapath.registerFile.regs[3][5] ));
 sg13g2_dfrbp_1 _3429_ (.CLK(clknet_5_10__leaf_clk_regs),
    .RESET_B(net170),
    .D(_0327_),
    .Q_N(_0122_),
    .Q(\crp.datapath.registerFile.regs[3][6] ));
 sg13g2_dfrbp_1 _3430_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net168),
    .D(_0328_),
    .Q_N(_0139_),
    .Q(\crp.datapath.registerFile.regs[3][7] ));
 sg13g2_dfrbp_1 _3431_ (.CLK(clknet_5_7__leaf_clk_regs),
    .RESET_B(net166),
    .D(_0329_),
    .Q_N(_0022_),
    .Q(\crp.datapath.registerFile.regs[9][0] ));
 sg13g2_dfrbp_1 _3432_ (.CLK(clknet_5_22__leaf_clk_regs),
    .RESET_B(net164),
    .D(_0330_),
    .Q_N(_0043_),
    .Q(\crp.datapath.registerFile.regs[9][1] ));
 sg13g2_dfrbp_1 _3433_ (.CLK(clknet_5_6__leaf_clk_regs),
    .RESET_B(net154),
    .D(_0331_),
    .Q_N(_0060_),
    .Q(\crp.datapath.registerFile.regs[9][2] ));
 sg13g2_dfrbp_1 _3434_ (.CLK(clknet_5_5__leaf_clk_regs),
    .RESET_B(net152),
    .D(_0332_),
    .Q_N(_0077_),
    .Q(\crp.datapath.registerFile.regs[9][3] ));
 sg13g2_dfrbp_1 _3435_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net150),
    .D(_0333_),
    .Q_N(_0094_),
    .Q(\crp.datapath.registerFile.regs[9][4] ));
 sg13g2_dfrbp_1 _3436_ (.CLK(clknet_5_19__leaf_clk_regs),
    .RESET_B(net148),
    .D(_0334_),
    .Q_N(_0111_),
    .Q(\crp.datapath.registerFile.regs[9][5] ));
 sg13g2_dfrbp_1 _3437_ (.CLK(clknet_5_18__leaf_clk_regs),
    .RESET_B(net146),
    .D(_0335_),
    .Q_N(_0128_),
    .Q(\crp.datapath.registerFile.regs[9][6] ));
 sg13g2_dfrbp_1 _3438_ (.CLK(clknet_5_17__leaf_clk_regs),
    .RESET_B(net144),
    .D(_0336_),
    .Q_N(_0145_),
    .Q(\crp.datapath.registerFile.regs[9][7] ));
 sg13g2_dfrbp_1 _3439_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net142),
    .D(_0337_),
    .Q_N(_0018_),
    .Q(\crp.datapath.registerFile.regs[6][0] ));
 sg13g2_dfrbp_1 _3440_ (.CLK(clknet_5_12__leaf_clk_regs),
    .RESET_B(net140),
    .D(_0338_),
    .Q_N(_0040_),
    .Q(\crp.datapath.registerFile.regs[6][1] ));
 sg13g2_dfrbp_1 _3441_ (.CLK(clknet_5_3__leaf_clk_regs),
    .RESET_B(net138),
    .D(_0339_),
    .Q_N(_0057_),
    .Q(\crp.datapath.registerFile.regs[6][2] ));
 sg13g2_dfrbp_1 _3442_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net136),
    .D(_0340_),
    .Q_N(_0074_),
    .Q(\crp.datapath.registerFile.regs[6][3] ));
 sg13g2_dfrbp_1 _3443_ (.CLK(clknet_5_1__leaf_clk_regs),
    .RESET_B(net134),
    .D(_0341_),
    .Q_N(_0091_),
    .Q(\crp.datapath.registerFile.regs[6][4] ));
 sg13g2_dfrbp_1 _3444_ (.CLK(clknet_5_4__leaf_clk_regs),
    .RESET_B(net31),
    .D(_0342_),
    .Q_N(_0108_),
    .Q(\crp.datapath.registerFile.regs[6][5] ));
 sg13g2_dfrbp_1 _3445_ (.CLK(clknet_5_0__leaf_clk_regs),
    .RESET_B(net19),
    .D(_0343_),
    .Q_N(_0125_),
    .Q(\crp.datapath.registerFile.regs[6][6] ));
 sg13g2_dfrbp_1 _3446_ (.CLK(clknet_5_9__leaf_clk_regs),
    .RESET_B(net15),
    .D(_0344_),
    .Q_N(_0142_),
    .Q(\crp.datapath.registerFile.regs[6][7] ));
 sg13g2_tiehi _3350__10 (.L_HI(net10));
 sg13g2_tiehi _3258__11 (.L_HI(net11));
 sg13g2_tiehi _3349__12 (.L_HI(net12));
 sg13g2_tiehi _3414__13 (.L_HI(net13));
 sg13g2_tiehi _3348__14 (.L_HI(net14));
 sg13g2_tiehi _3446__15 (.L_HI(net15));
 sg13g2_tiehi _3347__16 (.L_HI(net16));
 sg13g2_tiehi _3413__17 (.L_HI(net17));
 sg13g2_tiehi _3346__18 (.L_HI(net18));
 sg13g2_tiehi _3445__19 (.L_HI(net19));
 sg13g2_tiehi _3345__20 (.L_HI(net20));
 sg13g2_tiehi _3344__21 (.L_HI(net21));
 sg13g2_tiehi _3343__22 (.L_HI(net22));
 sg13g2_tiehi _3342__23 (.L_HI(net23));
 sg13g2_tiehi _3341__24 (.L_HI(net24));
 sg13g2_tiehi _3340__25 (.L_HI(net25));
 sg13g2_tiehi _3339__26 (.L_HI(net26));
 sg13g2_tiehi _3338__27 (.L_HI(net27));
 sg13g2_tiehi _3337__28 (.L_HI(net28));
 sg13g2_tiehi _3412__29 (.L_HI(net29));
 sg13g2_tiehi _3336__30 (.L_HI(net30));
 sg13g2_tiehi _3444__31 (.L_HI(net31));
 sg13g2_tiehi _3335__32 (.L_HI(net32));
 sg13g2_tiehi _3411__33 (.L_HI(net33));
 sg13g2_tiehi _3334__34 (.L_HI(net34));
 sg13g2_tiehi _3410__35 (.L_HI(net35));
 sg13g2_tiehi _3333__36 (.L_HI(net36));
 sg13g2_tiehi _3409__37 (.L_HI(net37));
 sg13g2_tiehi _3332__38 (.L_HI(net38));
 sg13g2_tiehi _3408__39 (.L_HI(net39));
 sg13g2_tiehi _3331__40 (.L_HI(net40));
 sg13g2_tiehi _3407__41 (.L_HI(net41));
 sg13g2_tiehi _3330__42 (.L_HI(net42));
 sg13g2_tiehi _3406__43 (.L_HI(net43));
 sg13g2_tiehi _3329__44 (.L_HI(net44));
 sg13g2_tiehi _3405__45 (.L_HI(net45));
 sg13g2_tiehi _3328__46 (.L_HI(net46));
 sg13g2_tiehi _3404__47 (.L_HI(net47));
 sg13g2_tiehi _3327__48 (.L_HI(net48));
 sg13g2_tiehi _3403__49 (.L_HI(net49));
 sg13g2_tiehi _3326__50 (.L_HI(net50));
 sg13g2_tiehi _3402__51 (.L_HI(net51));
 sg13g2_tiehi _3325__52 (.L_HI(net52));
 sg13g2_tiehi _3401__53 (.L_HI(net53));
 sg13g2_tiehi _3324__54 (.L_HI(net54));
 sg13g2_tiehi _3400__55 (.L_HI(net55));
 sg13g2_tiehi _3323__56 (.L_HI(net56));
 sg13g2_tiehi _3399__57 (.L_HI(net57));
 sg13g2_tiehi _3322__58 (.L_HI(net58));
 sg13g2_tiehi _3321__59 (.L_HI(net59));
 sg13g2_tiehi _3320__60 (.L_HI(net60));
 sg13g2_tiehi _3319__61 (.L_HI(net61));
 sg13g2_tiehi _3318__62 (.L_HI(net62));
 sg13g2_tiehi _3317__63 (.L_HI(net63));
 sg13g2_tiehi _3316__64 (.L_HI(net64));
 sg13g2_tiehi _3315__65 (.L_HI(net65));
 sg13g2_tiehi _3314__66 (.L_HI(net66));
 sg13g2_tiehi _3313__67 (.L_HI(net67));
 sg13g2_tiehi _3312__68 (.L_HI(net68));
 sg13g2_tiehi _3311__69 (.L_HI(net69));
 sg13g2_tiehi _3310__70 (.L_HI(net70));
 sg13g2_tiehi _3309__71 (.L_HI(net71));
 sg13g2_tiehi _3308__72 (.L_HI(net72));
 sg13g2_tiehi _3307__73 (.L_HI(net73));
 sg13g2_tiehi _3306__74 (.L_HI(net74));
 sg13g2_tiehi _3305__75 (.L_HI(net75));
 sg13g2_tiehi _3304__76 (.L_HI(net76));
 sg13g2_tiehi _3303__77 (.L_HI(net77));
 sg13g2_tiehi _3302__78 (.L_HI(net78));
 sg13g2_tiehi _3301__79 (.L_HI(net79));
 sg13g2_tiehi _3300__80 (.L_HI(net80));
 sg13g2_tiehi _3299__81 (.L_HI(net81));
 sg13g2_tiehi _3298__82 (.L_HI(net82));
 sg13g2_tiehi _3297__83 (.L_HI(net83));
 sg13g2_tiehi _3296__84 (.L_HI(net84));
 sg13g2_tiehi _3295__85 (.L_HI(net85));
 sg13g2_tiehi _3294__86 (.L_HI(net86));
 sg13g2_tiehi _3293__87 (.L_HI(net87));
 sg13g2_tiehi _3292__88 (.L_HI(net88));
 sg13g2_tiehi _3291__89 (.L_HI(net89));
 sg13g2_tiehi _3290__90 (.L_HI(net90));
 sg13g2_tiehi _3289__91 (.L_HI(net91));
 sg13g2_tiehi _3288__92 (.L_HI(net92));
 sg13g2_tiehi _3287__93 (.L_HI(net93));
 sg13g2_tiehi _3286__94 (.L_HI(net94));
 sg13g2_tiehi _3285__95 (.L_HI(net95));
 sg13g2_tiehi _3284__96 (.L_HI(net96));
 sg13g2_tiehi _3283__97 (.L_HI(net97));
 sg13g2_tiehi _3282__98 (.L_HI(net98));
 sg13g2_tiehi _3281__99 (.L_HI(net99));
 sg13g2_tiehi _3280__100 (.L_HI(net100));
 sg13g2_tiehi _3279__101 (.L_HI(net101));
 sg13g2_tiehi _3278__102 (.L_HI(net102));
 sg13g2_tiehi _3277__103 (.L_HI(net103));
 sg13g2_tiehi _3276__104 (.L_HI(net104));
 sg13g2_tiehi _3275__105 (.L_HI(net105));
 sg13g2_tiehi _3274__106 (.L_HI(net106));
 sg13g2_tiehi _3273__107 (.L_HI(net107));
 sg13g2_tiehi _3272__108 (.L_HI(net108));
 sg13g2_tiehi _3271__109 (.L_HI(net109));
 sg13g2_tiehi _3270__110 (.L_HI(net110));
 sg13g2_tiehi _3269__111 (.L_HI(net111));
 sg13g2_tiehi _3268__112 (.L_HI(net112));
 sg13g2_tiehi _3267__113 (.L_HI(net113));
 sg13g2_tiehi _3266__114 (.L_HI(net114));
 sg13g2_tiehi _3265__115 (.L_HI(net115));
 sg13g2_tiehi _3264__116 (.L_HI(net116));
 sg13g2_tiehi _3263__117 (.L_HI(net117));
 sg13g2_tiehi _3262__118 (.L_HI(net118));
 sg13g2_tiehi _3261__119 (.L_HI(net119));
 sg13g2_tiehi _3260__120 (.L_HI(net120));
 sg13g2_tiehi _3259__121 (.L_HI(net121));
 sg13g2_tiehi _3398__122 (.L_HI(net122));
 sg13g2_tiehi _3397__123 (.L_HI(net123));
 sg13g2_tiehi _3396__124 (.L_HI(net124));
 sg13g2_tiehi _3395__125 (.L_HI(net125));
 sg13g2_tiehi _3394__126 (.L_HI(net126));
 sg13g2_tiehi _3393__127 (.L_HI(net127));
 sg13g2_tiehi _3392__128 (.L_HI(net128));
 sg13g2_tiehi _3391__129 (.L_HI(net129));
 sg13g2_tiehi _3390__130 (.L_HI(net130));
 sg13g2_tiehi _3389__131 (.L_HI(net131));
 sg13g2_tiehi _3388__132 (.L_HI(net132));
 sg13g2_tiehi _3387__133 (.L_HI(net133));
 sg13g2_tiehi _3443__134 (.L_HI(net134));
 sg13g2_tiehi _3386__135 (.L_HI(net135));
 sg13g2_tiehi _3442__136 (.L_HI(net136));
 sg13g2_tiehi _3385__137 (.L_HI(net137));
 sg13g2_tiehi _3441__138 (.L_HI(net138));
 sg13g2_tiehi _3384__139 (.L_HI(net139));
 sg13g2_tiehi _3440__140 (.L_HI(net140));
 sg13g2_tiehi _3383__141 (.L_HI(net141));
 sg13g2_tiehi _3439__142 (.L_HI(net142));
 sg13g2_tiehi _3382__143 (.L_HI(net143));
 sg13g2_tiehi _3438__144 (.L_HI(net144));
 sg13g2_tiehi _3381__145 (.L_HI(net145));
 sg13g2_tiehi _3437__146 (.L_HI(net146));
 sg13g2_tiehi _3380__147 (.L_HI(net147));
 sg13g2_tiehi _3436__148 (.L_HI(net148));
 sg13g2_tiehi _3379__149 (.L_HI(net149));
 sg13g2_tiehi _3435__150 (.L_HI(net150));
 sg13g2_tiehi _3378__151 (.L_HI(net151));
 sg13g2_tiehi _3434__152 (.L_HI(net152));
 sg13g2_tiehi _3377__153 (.L_HI(net153));
 sg13g2_tiehi _3433__154 (.L_HI(net154));
 sg13g2_tiehi _3376__155 (.L_HI(net155));
 sg13g2_tiehi _3375__156 (.L_HI(net156));
 sg13g2_tiehi _3374__157 (.L_HI(net157));
 sg13g2_tiehi _3373__158 (.L_HI(net158));
 sg13g2_tiehi _3372__159 (.L_HI(net159));
 sg13g2_tiehi _3371__160 (.L_HI(net160));
 sg13g2_tiehi _3370__161 (.L_HI(net161));
 sg13g2_tiehi _3369__162 (.L_HI(net162));
 sg13g2_tiehi _3368__163 (.L_HI(net163));
 sg13g2_tiehi _3432__164 (.L_HI(net164));
 sg13g2_tiehi _3367__165 (.L_HI(net165));
 sg13g2_tiehi _3431__166 (.L_HI(net166));
 sg13g2_tiehi _3366__167 (.L_HI(net167));
 sg13g2_tiehi _3430__168 (.L_HI(net168));
 sg13g2_tiehi _3365__169 (.L_HI(net169));
 sg13g2_tiehi _3429__170 (.L_HI(net170));
 sg13g2_tiehi _3364__171 (.L_HI(net171));
 sg13g2_tiehi _3428__172 (.L_HI(net172));
 sg13g2_tiehi _3363__173 (.L_HI(net173));
 sg13g2_tiehi _3427__174 (.L_HI(net174));
 sg13g2_tiehi _3362__175 (.L_HI(net175));
 sg13g2_tiehi _3426__176 (.L_HI(net176));
 sg13g2_tiehi _3361__177 (.L_HI(net177));
 sg13g2_tiehi _3425__178 (.L_HI(net178));
 sg13g2_tiehi _3360__179 (.L_HI(net179));
 sg13g2_tiehi _3424__180 (.L_HI(net180));
 sg13g2_tiehi _3359__181 (.L_HI(net181));
 sg13g2_tiehi _3423__182 (.L_HI(net182));
 sg13g2_tiehi _3358__183 (.L_HI(net183));
 sg13g2_tiehi _3422__184 (.L_HI(net184));
 sg13g2_tiehi _3357__185 (.L_HI(net185));
 sg13g2_tiehi _3421__186 (.L_HI(net186));
 sg13g2_tiehi _3356__187 (.L_HI(net187));
 sg13g2_tiehi _3420__188 (.L_HI(net188));
 sg13g2_tiehi _3355__189 (.L_HI(net189));
 sg13g2_tiehi _3419__190 (.L_HI(net190));
 sg13g2_tiehi _3354__191 (.L_HI(net191));
 sg13g2_tiehi _3418__192 (.L_HI(net192));
 sg13g2_tiehi _3353__193 (.L_HI(net193));
 sg13g2_tiehi _3417__194 (.L_HI(net194));
 sg13g2_tiehi _3352__195 (.L_HI(net195));
 sg13g2_tiehi _3416__196 (.L_HI(net196));
 sg13g2_tiehi _3351__197 (.L_HI(net197));
 sg13g2_tiehi tt_um_rodald_cpr_198 (.L_HI(net198));
 sg13g2_tiehi tt_um_rodald_cpr_199 (.L_HI(net199));
 sg13g2_tiehi tt_um_rodald_cpr_200 (.L_HI(net200));
 sg13g2_tiehi tt_um_rodald_cpr_201 (.L_HI(net201));
 sg13g2_tiehi tt_um_rodald_cpr_202 (.L_HI(net202));
 sg13g2_tiehi tt_um_rodald_cpr_203 (.L_HI(net203));
 sg13g2_tiehi tt_um_rodald_cpr_204 (.L_HI(net204));
 sg13g2_tiehi tt_um_rodald_cpr_205 (.L_HI(net205));
 sg13g2_inv_1 _1920__1 (.Y(net206),
    .A(clknet_1_1__leaf_clk));
 sg13g2_buf_4 _3644_ (.X(uio_out[7]),
    .A(\crp.controller.mainDecoder.memWriteReq ));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(_1038_));
 sg13g2_buf_2 fanout557 (.A(_1038_),
    .X(net557));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(_1031_));
 sg13g2_buf_4 fanout559 (.X(net559),
    .A(_1031_));
 sg13g2_buf_4 fanout560 (.X(net560),
    .A(_1028_));
 sg13g2_buf_4 fanout561 (.X(net561),
    .A(_1028_));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(_1019_));
 sg13g2_buf_2 fanout563 (.A(_1019_),
    .X(net563));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(_1015_));
 sg13g2_buf_4 fanout565 (.X(net565),
    .A(_1015_));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(_1035_));
 sg13g2_buf_2 fanout567 (.A(_1035_),
    .X(net567));
 sg13g2_buf_4 fanout568 (.X(net568),
    .A(_1011_));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(_1011_));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(_1024_));
 sg13g2_buf_2 fanout571 (.A(_1024_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_0367_),
    .X(net573));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(_1142_));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(_1118_));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(_1102_));
 sg13g2_buf_2 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_1470_),
    .X(net578));
 sg13g2_buf_4 fanout579 (.X(net579),
    .A(_1072_));
 sg13g2_buf_4 fanout580 (.X(net580),
    .A(_1052_));
 sg13g2_buf_4 fanout581 (.X(net581),
    .A(_1050_));
 sg13g2_buf_4 fanout582 (.X(net582),
    .A(_1048_));
 sg13g2_buf_4 fanout583 (.X(net583),
    .A(_0475_));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(_0440_));
 sg13g2_buf_4 fanout585 (.X(net585),
    .A(_0397_));
 sg13g2_buf_2 fanout586 (.A(net587),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_8 fanout588 (.A(_1543_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_1 fanout590 (.A(net591),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_1498_),
    .X(net592));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(_1147_));
 sg13g2_buf_4 fanout594 (.X(net594),
    .A(_1145_));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(_1140_));
 sg13g2_buf_4 fanout596 (.X(net596),
    .A(_1116_));
 sg13g2_buf_4 fanout597 (.X(net597),
    .A(_1043_));
 sg13g2_buf_4 fanout598 (.X(net598),
    .A(_1040_));
 sg13g2_buf_2 fanout599 (.A(_1007_),
    .X(net599));
 sg13g2_buf_1 fanout600 (.A(_1007_),
    .X(net600));
 sg13g2_buf_4 fanout601 (.X(net601),
    .A(_0672_));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(_0671_));
 sg13g2_buf_2 fanout603 (.A(_1056_),
    .X(net603));
 sg13g2_buf_1 fanout604 (.A(_1056_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(net606),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_1055_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_1001_),
    .X(net608));
 sg13g2_buf_4 fanout609 (.X(net609),
    .A(net610));
 sg13g2_buf_4 fanout610 (.X(net610),
    .A(_1391_));
 sg13g2_buf_2 fanout611 (.A(net614),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(net614),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_1374_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_1303_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_1075_),
    .X(net616));
 sg13g2_buf_1 fanout617 (.A(_1075_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(net619),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_1074_),
    .X(net620));
 sg13g2_buf_4 fanout621 (.X(net621),
    .A(_1509_));
 sg13g2_buf_2 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_1390_),
    .X(net623));
 sg13g2_buf_4 fanout624 (.X(net624),
    .A(_1385_));
 sg13g2_buf_1 fanout625 (.A(_1385_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_1384_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_1356_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(net630),
    .X(net628));
 sg13g2_buf_1 fanout629 (.A(net630),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_1354_),
    .X(net630));
 sg13g2_buf_4 fanout631 (.X(net631),
    .A(_1353_));
 sg13g2_buf_1 fanout632 (.A(_1353_),
    .X(net632));
 sg13g2_buf_4 fanout633 (.X(net633),
    .A(_1452_));
 sg13g2_buf_4 fanout634 (.X(net634),
    .A(_1448_));
 sg13g2_buf_2 fanout635 (.A(_1448_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net637),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_1448_),
    .X(net637));
 sg13g2_buf_4 fanout638 (.X(net638),
    .A(_1446_));
 sg13g2_buf_8 fanout639 (.A(_1446_),
    .X(net639));
 sg13g2_buf_4 fanout640 (.X(net640),
    .A(_1445_));
 sg13g2_buf_4 fanout641 (.X(net641),
    .A(_1445_));
 sg13g2_buf_2 fanout642 (.A(net643),
    .X(net642));
 sg13g2_buf_4 fanout643 (.X(net643),
    .A(net644));
 sg13g2_buf_4 fanout644 (.X(net644),
    .A(_1444_));
 sg13g2_buf_4 fanout645 (.X(net645),
    .A(_1444_));
 sg13g2_buf_4 fanout646 (.X(net646),
    .A(_1444_));
 sg13g2_buf_4 fanout647 (.X(net647),
    .A(_1438_));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(_1407_));
 sg13g2_buf_2 fanout649 (.A(_1407_),
    .X(net649));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(_1406_));
 sg13g2_buf_8 fanout651 (.A(net655),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(net655),
    .X(net652));
 sg13g2_buf_8 fanout653 (.A(net655),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(net655),
    .X(net654));
 sg13g2_buf_4 fanout655 (.X(net655),
    .A(_1403_));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(net657));
 sg13g2_buf_4 fanout657 (.X(net657),
    .A(_1402_));
 sg13g2_buf_4 fanout658 (.X(net658),
    .A(net659));
 sg13g2_buf_8 fanout659 (.A(_1400_),
    .X(net659));
 sg13g2_buf_4 fanout660 (.X(net660),
    .A(net661));
 sg13g2_buf_8 fanout661 (.A(_1400_),
    .X(net661));
 sg13g2_buf_16 fanout662 (.X(net662),
    .A(net664));
 sg13g2_buf_2 fanout663 (.A(net664),
    .X(net663));
 sg13g2_buf_8 fanout664 (.A(_1399_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_1355_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_1355_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_1006_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(net670),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net670),
    .X(net669));
 sg13g2_buf_4 fanout670 (.X(net670),
    .A(net678));
 sg13g2_buf_2 fanout671 (.A(net678),
    .X(net671));
 sg13g2_buf_1 fanout672 (.A(net678),
    .X(net672));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(net674));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(net676));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(net676));
 sg13g2_buf_8 fanout676 (.A(net678),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(_1398_));
 sg13g2_buf_2 fanout679 (.A(net681),
    .X(net679));
 sg13g2_buf_16 fanout680 (.X(net680),
    .A(net681));
 sg13g2_buf_16 fanout681 (.X(net681),
    .A(net683));
 sg13g2_buf_2 fanout682 (.A(net683),
    .X(net682));
 sg13g2_buf_8 fanout683 (.A(_1397_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(net687),
    .X(net684));
 sg13g2_buf_4 fanout685 (.X(net685),
    .A(net686));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_1339_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_1105_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_1105_),
    .X(net689));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(_1091_));
 sg13g2_buf_2 fanout691 (.A(_1091_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_1305_),
    .X(net693));
 sg13g2_buf_4 fanout694 (.X(net694),
    .A(net696));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(net697),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_1279_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_1264_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_1264_),
    .X(net699));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(\crp.controller.aluDec.aluRtypeDec.state[2] ));
 sg13g2_buf_8 fanout701 (.A(\crp.controller.aluDec.aluRtypeDec.state[1] ),
    .X(net701));
 sg13g2_buf_4 fanout702 (.X(net702),
    .A(\crp.controller.aluDec.aluRtypeDec.state[0] ));
 sg13g2_buf_2 fanout703 (.A(\crp.controller.aluDec.aluRtypeDec.state[0] ),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(_1208_));
 sg13g2_buf_2 fanout705 (.A(_1208_),
    .X(net705));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(net707));
 sg13g2_buf_2 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(_1207_));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(net712));
 sg13g2_buf_2 fanout710 (.A(net711),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(net712),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(_1190_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(net721),
    .X(net713));
 sg13g2_buf_1 fanout714 (.A(net721),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(net721),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(net718),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(net719),
    .X(net718));
 sg13g2_buf_1 fanout719 (.A(net720),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(net721),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_0029_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(net723),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(net388),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(net725),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(\crp.controller.aluDec.aluRtypeDec.func[2] ),
    .X(net725));
 sg13g2_buf_4 fanout726 (.X(net726),
    .A(\crp.controller.aluDec.aluRtypeDec.func[1] ));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(\crp.controller.aluDec.aluRtypeDec.func[0] ));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(\crp.controller.aluDec.opcode[3] ));
 sg13g2_buf_4 fanout729 (.X(net729),
    .A(net735));
 sg13g2_buf_2 fanout730 (.A(net735),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(net732),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(net735),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(net735),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(net735),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_0011_),
    .X(net735));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(_1189_));
 sg13g2_buf_1 fanout737 (.A(_1189_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_1189_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(net745),
    .X(net739));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(net745));
 sg13g2_buf_1 fanout741 (.A(net745),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(net744),
    .X(net742));
 sg13g2_buf_1 fanout743 (.A(net744),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(net745),
    .X(net744));
 sg13g2_buf_4 fanout745 (.X(net745),
    .A(rst_n));
 sg13g2_buf_4 input1 (.X(net1),
    .A(ui_in[0]));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[1]));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[2]));
 sg13g2_buf_4 input4 (.X(net4),
    .A(ui_in[3]));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tiehi _3415__9 (.L_HI(net9));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_2 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0152_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold2 (.A(\crp.datapath.aluSrc1SelMux.d0[13] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold3 (.A(\crp.datapath.aluSrc1SelMux.d0[2] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold4 (.A(\crp.datapath.aluSrc1SelMux.d0[11] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold5 (.A(\crp.datapath.registerFile.regs[11][1] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold6 (.A(\crp.datapath.registerFile.regs[6][0] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold7 (.A(\crp.datapath.registerFile.regs[7][0] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold8 (.A(\crp.datapath.registerFile.regs[12][0] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold9 (.A(\crp.datapath.aluSrc1SelMux.d0[10] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold10 (.A(\crp.datapath.registerFile.regs[13][0] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold11 (.A(\crp.datapath.registerFile.regs[6][1] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold12 (.A(\crp.datapath.registerFile.regs[14][0] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold13 (.A(\crp.datapath.registerFile.regs[11][0] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold14 (.A(\crp.datapath.aluSrc1SelMux.d0[14] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold15 (.A(\crp.datapath.registerFile.regs[2][0] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold16 (.A(\crp.datapath.registerFile.regs[3][0] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0321_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold18 (.A(\crp.datapath.registerFile.regs[10][0] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold19 (.A(\crp.datapath.registerFile.regs[3][1] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold20 (.A(\crp.datapath.registerFile.regs[15][0] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold21 (.A(\crp.datapath.registerFile.regs[5][3] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold22 (.A(\crp.datapath.aluSrc1SelMux.d0[4] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold23 (.A(\crp.datapath.registerFile.regs[12][6] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold24 (.A(\crp.datapath.registerFile.regs[0][7] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold25 (.A(\crp.datapath.registerFile.regs[15][5] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold26 (.A(\crp.datapath.registerFile.regs[13][5] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold27 (.A(\crp.datapath.registerFile.regs[1][2] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold28 (.A(\crp.datapath.registerFile.regs[10][6] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold29 (.A(\crp.datapath.registerFile.regs[3][3] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold30 (.A(\crp.datapath.registerFile.regs[14][5] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold31 (.A(\crp.datapath.registerFile.regs[2][7] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold32 (.A(\crp.datapath.registerFile.regs[13][6] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold33 (.A(\crp.datapath.registerFile.regs[12][5] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold34 (.A(\crp.datapath.registerFile.regs[2][3] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold35 (.A(\crp.datapath.registerFile.regs[7][3] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold36 (.A(\crp.datapath.registerFile.regs[6][3] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold37 (.A(\crp.datapath.registerFile.regs[10][5] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold38 (.A(\crp.datapath.registerFile.regs[13][3] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold39 (.A(\crp.datapath.registerFile.regs[7][6] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold40 (.A(\crp.datapath.registerFile.regs[13][7] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold41 (.A(\crp.datapath.registerFile.regs[11][5] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold42 (.A(\crp.datapath.registerFile.regs[12][7] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold43 (.A(\crp.datapath.registerFile.regs[0][6] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold44 (.A(\crp.datapath.registerFile.regs[1][5] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold45 (.A(\crp.datapath.registerFile.regs[0][5] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold46 (.A(\crp.datapath.registerFile.regs[1][7] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold47 (.A(\crp.datapath.registerFile.regs[4][6] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold48 (.A(\crp.datapath.registerFile.regs[12][4] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold49 (.A(\crp.datapath.registerFile.regs[11][3] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold50 (.A(\crp.datapath.registerFile.regs[8][6] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold51 (.A(\crp.datapath.registerFile.regs[6][6] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold52 (.A(\crp.datapath.registerFile.regs[9][2] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold53 (.A(\crp.datapath.registerFile.regs[0][4] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold54 (.A(\crp.datapath.registerFile.regs[14][6] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold55 (.A(\crp.datapath.registerFile.regs[1][4] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold56 (.A(\crp.datapath.registerFile.regs[2][4] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold57 (.A(\crp.datapath.registerFile.regs[9][7] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold58 (.A(\crp.datapath.registerFile.regs[9][5] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold59 (.A(\crp.datapath.registerFile.regs[5][4] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold60 (.A(\crp.datapath.registerFile.regs[5][6] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold61 (.A(\crp.datapath.registerFile.regs[8][5] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold62 (.A(\crp.datapath.registerFile.regs[4][4] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold63 (.A(\crp.datapath.registerFile.regs[4][5] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold64 (.A(\crp.datapath.registerFile.regs[14][3] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold65 (.A(\crp.datapath.registerFile.regs[10][4] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold66 (.A(\crp.datapath.registerFile.regs[14][7] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold67 (.A(\crp.datapath.registerFile.regs[7][7] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold68 (.A(\crp.datapath.registerFile.regs[2][5] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold69 (.A(\crp.datapath.registerFile.regs[14][4] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold70 (.A(\crp.datapath.registerFile.regs[11][7] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold71 (.A(\crp.datapath.registerFile.regs[5][7] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold72 (.A(\crp.datapath.registerFile.regs[13][4] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold73 (.A(\crp.datapath.registerFile.regs[15][3] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold74 (.A(\crp.datapath.registerFile.regs[7][4] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold75 (.A(\crp.datapath.registerFile.regs[12][3] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold76 (.A(\crp.datapath.registerFile.regs[6][4] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold77 (.A(\crp.datapath.registerFile.regs[3][7] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold78 (.A(\crp.datapath.registerFile.regs[8][3] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold79 (.A(\crp.datapath.registerFile.regs[11][4] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold80 (.A(\crp.datapath.registerFile.regs[3][6] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold81 (.A(\crp.datapath.registerFile.regs[1][3] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold82 (.A(\crp.datapath.registerFile.regs[8][7] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold83 (.A(\crp.datapath.registerFile.regs[9][4] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold84 (.A(\crp.datapath.registerFile.regs[6][7] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold85 (.A(\crp.datapath.registerFile.regs[5][5] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold86 (.A(\crp.datapath.registerFile.regs[8][4] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold87 (.A(\crp.datapath.registerFile.regs[15][7] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0195_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold89 (.A(\crp.datapath.registerFile.regs[9][3] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold90 (.A(\crp.datapath.registerFile.regs[10][7] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold91 (.A(\crp.controller.aluDec.opcode[3] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold92 (.A(\crp.datapath.registerFile.regs[9][6] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold93 (.A(\crp.datapath.registerFile.regs[0][3] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold94 (.A(\crp.datapath.registerFile.regs[1][6] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold95 (.A(\crp.datapath.aluSrc1SelMux.d0[6] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold96 (.A(\crp.datapath.registerFile.regs[6][5] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold97 (.A(\crp.datapath.registerFile.regs[5][2] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold98 (.A(\crp.datapath.registerFile.regs[15][4] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold99 (.A(\crp.datapath.aluSrc1SelMux.d1[13] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold100 (.A(\crp.datapath.registerFile.regs[4][3] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold101 (.A(\crp.datapath.registerFile.regs[6][2] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold102 (.A(\crp.datapath.registerFile.regs[15][6] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold103 (.A(\crp.datapath.registerFile.regs[3][4] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold104 (.A(\crp.datapath.registerFile.regs[7][5] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold105 (.A(\crp.datapath.registerFile.regs[2][6] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold106 (.A(\crp.datapath.registerFile.regs[11][6] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold107 (.A(\crp.datapath.registerFile.regs[3][5] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold108 (.A(\crp.datapath.registerFile.regs[4][7] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold109 (.A(\crp.datapath.registerFile.regs[10][3] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold110 (.A(\crp.datapath.registerFile.regs[10][2] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold111 (.A(\crp.datapath.registerFile.regs[2][2] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold112 (.A(\crp.datapath.aluSrc1SelMux.d0[9] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold113 (.A(\crp.datapath.aluSrc2SelMux.d2[4] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold114 (.A(\crp.datapath.aluSrc1SelMux.d1[11] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold115 (.A(\crp.datapath.registerFile.regs[1][1] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold116 (.A(\crp.datapath.registerFile.regs[3][2] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold117 (.A(\crp.datapath.registerFile.regs[0][0] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold118 (.A(\crp.datapath.registerFile.regs[13][1] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold119 (.A(\crp.datapath.registerFile.regs[15][2] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold120 (.A(\crp.datapath.registerFile.regs[8][0] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold121 (.A(\crp.datapath.registerFile.regs[11][2] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold122 (.A(\crp.datapath.registerFile.regs[7][2] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold123 (.A(\crp.datapath.registerFile.regs[1][0] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold124 (.A(\crp.datapath.aluSrc2SelMux.d2[6] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold125 (.A(\crp.datapath.registerFile.regs[7][1] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold126 (.A(\crp.datapath.registerFile.regs[5][1] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold127 (.A(\crp.datapath.registerFile.regs[4][0] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold128 (.A(\crp.datapath.registerFile.regs[2][1] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold129 (.A(\crp.datapath.aluSrc1SelMux.d0[5] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold130 (.A(\crp.datapath.registerFile.regs[12][1] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold131 (.A(\crp.datapath.registerFile.regs[5][0] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold132 (.A(\crp.datapath.registerFile.regs[0][1] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold133 (.A(\crp.datapath.registerFile.regs[8][2] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold134 (.A(\crp.datapath.registerFile.regs[12][2] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold135 (.A(\crp.datapath.registerFile.regs[9][0] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold136 (.A(\crp.datapath.registerFile.regs[13][2] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold137 (.A(\crp.datapath.aluSrc1SelMux.d1[10] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold138 (.A(\crp.datapath.registerFile.regs[0][2] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold139 (.A(\crp.datapath.registerFile.regs[4][2] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold140 (.A(\crp.datapath.registerFile.regs[14][1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold141 (.A(\crp.datapath.registerFile.regs[4][1] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold142 (.A(\crp.datapath.aluSrc2SelMux.d2[5] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold143 (.A(\crp.datapath.registerFile.regs[14][2] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold144 (.A(\crp.datapath.aluSrc1SelMux.d1[4] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold145 (.A(\crp.datapath.registerFile.regs[15][1] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold146 (.A(\crp.datapath.aluSrc1SelMux.d0[3] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold147 (.A(\crp.datapath.registerFile.regs[10][1] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold148 (.A(\crp.datapath.registerFile.regs[9][1] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold149 (.A(\crp.datapath.registerFile.regs[8][1] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold150 (.A(\crp.datapath.aluSrc1SelMux.d1[14] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold151 (.A(\crp.datapath.aluSrc1SelMux.d0[7] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold152 (.A(\crp.datapath.aluSrc1SelMux.d1[6] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold153 (.A(\crp.datapath.aluSrc1SelMux.d0[0] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold154 (.A(\crp.datapath.aluSrc1SelMux.d1[5] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold155 (.A(\crp.datapath.aluSrc1SelMux.d0[12] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold156 (.A(\crp.datapath.aluSrc2SelMux.d2[7] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold157 (.A(\crp.datapath.aluSrc1SelMux.d1[9] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold158 (.A(\crp.datapath.aluSrc1SelMux.d0[1] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold159 (.A(\crp.datapath.aluSrc1SelMux.d1[2] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold160 (.A(\crp.controller.flags[1] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold161 (.A(\crp.datapath.aluSrc1SelMux.d1[3] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold162 (.A(\crp.datapath.aluSrc1SelMux.d1[8] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold163 (.A(\crp.datapath.aluSrc1SelMux.d1[7] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold164 (.A(\crp.datapath.aluSrc1SelMux.d0[8] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold165 (.A(\crp.datapath.aluSrc2SelMux.d3[12] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold166 (.A(\crp.datapath.aluSrc2SelMux.d3[11] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold167 (.A(\crp.datapath.aluSrc1SelMux.d1[12] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold168 (.A(\crp.controller.flags[3] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold169 (.A(\crp.controller.flags[0] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold170 (.A(\crp.controller.aluDec.opcode[0] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold171 (.A(\crp.datapath.aluSrc1SelMux.d1[0] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold172 (.A(\crp.controller.flags[2] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold173 (.A(\crp.datapath.aluSrc2SelMux.d3[10] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold174 (.A(\crp.datapath.aluSrc2SelMux.d3[9] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold175 (.A(\crp.datapath.aluSrc1SelMux.d1[1] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold176 (.A(\crp.controller.aluDec.opcode[1] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold177 (.A(\crp.controller.aluDec.opcode[2] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0007_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold179 (.A(_1336_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold180 (.A(\crp.controller.aluDec.aluRtypeDec.func[3] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold181 (.A(\crp.controller.aluDec.aluRtypeDec.func[0] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold182 (.A(net701),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold183 (.A(_1262_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold184 (.A(\crp.datapath.aluSrc2SelMux.d3[12] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold185 (.A(\crp.datapath.aluSrc2SelMux.d3[11] ),
    .X(net393));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_fill_2 FILLER_0_91 ();
 sg13g2_fill_1 FILLER_0_93 ();
 sg13g2_decap_8 FILLER_0_113 ();
 sg13g2_decap_8 FILLER_0_120 ();
 sg13g2_decap_8 FILLER_0_127 ();
 sg13g2_decap_8 FILLER_0_134 ();
 sg13g2_decap_8 FILLER_0_141 ();
 sg13g2_decap_8 FILLER_0_148 ();
 sg13g2_decap_8 FILLER_0_155 ();
 sg13g2_decap_8 FILLER_0_162 ();
 sg13g2_decap_8 FILLER_0_169 ();
 sg13g2_decap_8 FILLER_0_176 ();
 sg13g2_decap_8 FILLER_0_183 ();
 sg13g2_decap_8 FILLER_0_190 ();
 sg13g2_decap_8 FILLER_0_197 ();
 sg13g2_decap_8 FILLER_0_204 ();
 sg13g2_decap_8 FILLER_0_211 ();
 sg13g2_decap_8 FILLER_0_218 ();
 sg13g2_decap_8 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_232 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_253 ();
 sg13g2_decap_8 FILLER_0_260 ();
 sg13g2_decap_8 FILLER_0_267 ();
 sg13g2_decap_8 FILLER_0_274 ();
 sg13g2_decap_8 FILLER_0_281 ();
 sg13g2_decap_8 FILLER_0_288 ();
 sg13g2_decap_8 FILLER_0_295 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_4 FILLER_1_77 ();
 sg13g2_decap_4 FILLER_1_107 ();
 sg13g2_decap_4 FILLER_1_121 ();
 sg13g2_fill_2 FILLER_1_125 ();
 sg13g2_fill_2 FILLER_1_131 ();
 sg13g2_fill_1 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_160 ();
 sg13g2_decap_8 FILLER_1_167 ();
 sg13g2_decap_8 FILLER_1_174 ();
 sg13g2_decap_8 FILLER_1_181 ();
 sg13g2_decap_8 FILLER_1_188 ();
 sg13g2_decap_8 FILLER_1_195 ();
 sg13g2_decap_8 FILLER_1_202 ();
 sg13g2_decap_8 FILLER_1_209 ();
 sg13g2_decap_8 FILLER_1_216 ();
 sg13g2_decap_8 FILLER_1_223 ();
 sg13g2_decap_8 FILLER_1_230 ();
 sg13g2_decap_8 FILLER_1_237 ();
 sg13g2_decap_8 FILLER_1_244 ();
 sg13g2_decap_8 FILLER_1_251 ();
 sg13g2_decap_8 FILLER_1_258 ();
 sg13g2_decap_8 FILLER_1_265 ();
 sg13g2_decap_8 FILLER_1_272 ();
 sg13g2_decap_8 FILLER_1_279 ();
 sg13g2_decap_8 FILLER_1_286 ();
 sg13g2_decap_8 FILLER_1_293 ();
 sg13g2_decap_8 FILLER_1_300 ();
 sg13g2_decap_8 FILLER_1_307 ();
 sg13g2_decap_8 FILLER_1_314 ();
 sg13g2_decap_8 FILLER_1_321 ();
 sg13g2_decap_8 FILLER_1_328 ();
 sg13g2_decap_8 FILLER_1_335 ();
 sg13g2_decap_8 FILLER_1_342 ();
 sg13g2_decap_8 FILLER_1_349 ();
 sg13g2_decap_8 FILLER_1_356 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_8 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_fill_2 FILLER_2_70 ();
 sg13g2_fill_1 FILLER_2_72 ();
 sg13g2_fill_2 FILLER_2_83 ();
 sg13g2_fill_1 FILLER_2_85 ();
 sg13g2_fill_1 FILLER_2_112 ();
 sg13g2_decap_4 FILLER_2_139 ();
 sg13g2_fill_1 FILLER_2_143 ();
 sg13g2_decap_8 FILLER_2_170 ();
 sg13g2_decap_8 FILLER_2_177 ();
 sg13g2_decap_8 FILLER_2_184 ();
 sg13g2_decap_8 FILLER_2_191 ();
 sg13g2_decap_8 FILLER_2_198 ();
 sg13g2_decap_8 FILLER_2_205 ();
 sg13g2_decap_8 FILLER_2_212 ();
 sg13g2_decap_8 FILLER_2_219 ();
 sg13g2_decap_8 FILLER_2_226 ();
 sg13g2_decap_8 FILLER_2_233 ();
 sg13g2_decap_8 FILLER_2_240 ();
 sg13g2_decap_8 FILLER_2_247 ();
 sg13g2_decap_8 FILLER_2_254 ();
 sg13g2_decap_8 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_268 ();
 sg13g2_decap_8 FILLER_2_275 ();
 sg13g2_decap_8 FILLER_2_282 ();
 sg13g2_decap_8 FILLER_2_289 ();
 sg13g2_decap_8 FILLER_2_296 ();
 sg13g2_decap_8 FILLER_2_303 ();
 sg13g2_decap_8 FILLER_2_310 ();
 sg13g2_decap_8 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_331 ();
 sg13g2_decap_8 FILLER_2_338 ();
 sg13g2_decap_8 FILLER_2_345 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_4 FILLER_3_63 ();
 sg13g2_fill_1 FILLER_3_67 ();
 sg13g2_fill_1 FILLER_3_94 ();
 sg13g2_fill_2 FILLER_3_105 ();
 sg13g2_fill_1 FILLER_3_143 ();
 sg13g2_fill_2 FILLER_3_159 ();
 sg13g2_decap_8 FILLER_3_187 ();
 sg13g2_decap_8 FILLER_3_194 ();
 sg13g2_decap_8 FILLER_3_201 ();
 sg13g2_decap_8 FILLER_3_208 ();
 sg13g2_decap_8 FILLER_3_215 ();
 sg13g2_decap_8 FILLER_3_222 ();
 sg13g2_decap_8 FILLER_3_229 ();
 sg13g2_decap_8 FILLER_3_236 ();
 sg13g2_decap_8 FILLER_3_243 ();
 sg13g2_decap_8 FILLER_3_250 ();
 sg13g2_decap_8 FILLER_3_257 ();
 sg13g2_decap_8 FILLER_3_264 ();
 sg13g2_decap_8 FILLER_3_271 ();
 sg13g2_decap_8 FILLER_3_278 ();
 sg13g2_decap_8 FILLER_3_285 ();
 sg13g2_decap_8 FILLER_3_292 ();
 sg13g2_decap_8 FILLER_3_299 ();
 sg13g2_decap_8 FILLER_3_306 ();
 sg13g2_decap_8 FILLER_3_313 ();
 sg13g2_decap_8 FILLER_3_320 ();
 sg13g2_decap_8 FILLER_3_327 ();
 sg13g2_decap_8 FILLER_3_334 ();
 sg13g2_decap_8 FILLER_3_341 ();
 sg13g2_decap_8 FILLER_3_348 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_decap_8 FILLER_3_362 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_fill_1 FILLER_4_77 ();
 sg13g2_fill_2 FILLER_4_95 ();
 sg13g2_decap_4 FILLER_4_101 ();
 sg13g2_fill_1 FILLER_4_105 ();
 sg13g2_fill_1 FILLER_4_115 ();
 sg13g2_decap_4 FILLER_4_138 ();
 sg13g2_fill_1 FILLER_4_150 ();
 sg13g2_fill_1 FILLER_4_176 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_fill_2 FILLER_5_70 ();
 sg13g2_fill_1 FILLER_5_72 ();
 sg13g2_fill_2 FILLER_5_83 ();
 sg13g2_fill_1 FILLER_5_85 ();
 sg13g2_decap_8 FILLER_5_100 ();
 sg13g2_decap_8 FILLER_5_107 ();
 sg13g2_fill_2 FILLER_5_114 ();
 sg13g2_fill_1 FILLER_5_126 ();
 sg13g2_decap_4 FILLER_5_131 ();
 sg13g2_decap_8 FILLER_5_145 ();
 sg13g2_decap_8 FILLER_5_152 ();
 sg13g2_decap_4 FILLER_5_166 ();
 sg13g2_fill_2 FILLER_5_170 ();
 sg13g2_decap_8 FILLER_5_176 ();
 sg13g2_decap_8 FILLER_5_183 ();
 sg13g2_decap_8 FILLER_5_190 ();
 sg13g2_decap_8 FILLER_5_197 ();
 sg13g2_decap_8 FILLER_5_204 ();
 sg13g2_decap_8 FILLER_5_211 ();
 sg13g2_decap_8 FILLER_5_218 ();
 sg13g2_decap_8 FILLER_5_225 ();
 sg13g2_decap_8 FILLER_5_232 ();
 sg13g2_decap_8 FILLER_5_239 ();
 sg13g2_decap_8 FILLER_5_246 ();
 sg13g2_decap_8 FILLER_5_253 ();
 sg13g2_decap_8 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_267 ();
 sg13g2_decap_8 FILLER_5_274 ();
 sg13g2_decap_8 FILLER_5_281 ();
 sg13g2_decap_8 FILLER_5_288 ();
 sg13g2_decap_8 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_4 FILLER_6_63 ();
 sg13g2_fill_2 FILLER_6_67 ();
 sg13g2_decap_4 FILLER_6_105 ();
 sg13g2_fill_2 FILLER_6_109 ();
 sg13g2_decap_8 FILLER_6_142 ();
 sg13g2_fill_2 FILLER_6_159 ();
 sg13g2_fill_1 FILLER_6_161 ();
 sg13g2_fill_2 FILLER_6_171 ();
 sg13g2_fill_1 FILLER_6_173 ();
 sg13g2_decap_8 FILLER_6_179 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_4 FILLER_7_63 ();
 sg13g2_decap_4 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_205 ();
 sg13g2_decap_8 FILLER_7_212 ();
 sg13g2_decap_8 FILLER_7_219 ();
 sg13g2_decap_8 FILLER_7_226 ();
 sg13g2_decap_8 FILLER_7_233 ();
 sg13g2_decap_8 FILLER_7_240 ();
 sg13g2_decap_8 FILLER_7_247 ();
 sg13g2_decap_8 FILLER_7_254 ();
 sg13g2_decap_8 FILLER_7_277 ();
 sg13g2_decap_8 FILLER_7_284 ();
 sg13g2_decap_8 FILLER_7_291 ();
 sg13g2_decap_8 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_decap_8 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_326 ();
 sg13g2_decap_8 FILLER_7_333 ();
 sg13g2_decap_8 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_347 ();
 sg13g2_decap_8 FILLER_7_354 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_4 FILLER_8_56 ();
 sg13g2_fill_1 FILLER_8_60 ();
 sg13g2_decap_4 FILLER_8_87 ();
 sg13g2_fill_2 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_149 ();
 sg13g2_fill_1 FILLER_8_156 ();
 sg13g2_decap_4 FILLER_8_167 ();
 sg13g2_fill_2 FILLER_8_171 ();
 sg13g2_fill_2 FILLER_8_177 ();
 sg13g2_decap_8 FILLER_8_209 ();
 sg13g2_decap_8 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_fill_2 FILLER_8_285 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_4 FILLER_9_42 ();
 sg13g2_fill_2 FILLER_9_46 ();
 sg13g2_fill_1 FILLER_9_78 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_fill_2 FILLER_9_95 ();
 sg13g2_fill_2 FILLER_9_114 ();
 sg13g2_fill_1 FILLER_9_116 ();
 sg13g2_fill_2 FILLER_9_127 ();
 sg13g2_fill_2 FILLER_9_152 ();
 sg13g2_fill_2 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_181 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_215 ();
 sg13g2_decap_8 FILLER_9_222 ();
 sg13g2_decap_8 FILLER_9_229 ();
 sg13g2_decap_4 FILLER_9_236 ();
 sg13g2_fill_2 FILLER_9_243 ();
 sg13g2_fill_1 FILLER_9_245 ();
 sg13g2_fill_2 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_307 ();
 sg13g2_decap_8 FILLER_9_314 ();
 sg13g2_decap_8 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_328 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_4 FILLER_10_49 ();
 sg13g2_fill_2 FILLER_10_53 ();
 sg13g2_fill_1 FILLER_10_78 ();
 sg13g2_fill_2 FILLER_10_89 ();
 sg13g2_fill_2 FILLER_10_100 ();
 sg13g2_fill_1 FILLER_10_102 ();
 sg13g2_fill_1 FILLER_10_113 ();
 sg13g2_fill_2 FILLER_10_131 ();
 sg13g2_fill_1 FILLER_10_133 ();
 sg13g2_fill_2 FILLER_10_153 ();
 sg13g2_fill_1 FILLER_10_155 ();
 sg13g2_fill_2 FILLER_10_176 ();
 sg13g2_fill_1 FILLER_10_178 ();
 sg13g2_decap_4 FILLER_10_188 ();
 sg13g2_decap_8 FILLER_10_211 ();
 sg13g2_decap_8 FILLER_10_218 ();
 sg13g2_decap_8 FILLER_10_225 ();
 sg13g2_fill_2 FILLER_10_232 ();
 sg13g2_fill_2 FILLER_10_249 ();
 sg13g2_fill_2 FILLER_10_263 ();
 sg13g2_fill_1 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_decap_8 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_334 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_decap_8 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_4 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_53 ();
 sg13g2_decap_4 FILLER_11_69 ();
 sg13g2_fill_2 FILLER_11_109 ();
 sg13g2_fill_2 FILLER_11_116 ();
 sg13g2_fill_1 FILLER_11_161 ();
 sg13g2_fill_1 FILLER_11_188 ();
 sg13g2_decap_8 FILLER_11_215 ();
 sg13g2_decap_8 FILLER_11_222 ();
 sg13g2_fill_2 FILLER_11_229 ();
 sg13g2_fill_1 FILLER_11_231 ();
 sg13g2_fill_2 FILLER_11_280 ();
 sg13g2_fill_1 FILLER_11_282 ();
 sg13g2_fill_2 FILLER_11_288 ();
 sg13g2_fill_1 FILLER_11_290 ();
 sg13g2_decap_8 FILLER_11_300 ();
 sg13g2_decap_8 FILLER_11_307 ();
 sg13g2_decap_8 FILLER_11_314 ();
 sg13g2_decap_8 FILLER_11_321 ();
 sg13g2_decap_8 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_335 ();
 sg13g2_decap_8 FILLER_11_342 ();
 sg13g2_decap_8 FILLER_11_349 ();
 sg13g2_decap_8 FILLER_11_356 ();
 sg13g2_decap_8 FILLER_11_363 ();
 sg13g2_decap_8 FILLER_11_370 ();
 sg13g2_decap_8 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_4 FILLER_12_42 ();
 sg13g2_fill_2 FILLER_12_46 ();
 sg13g2_fill_1 FILLER_12_83 ();
 sg13g2_decap_8 FILLER_12_88 ();
 sg13g2_fill_2 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_152 ();
 sg13g2_fill_2 FILLER_12_158 ();
 sg13g2_decap_8 FILLER_12_177 ();
 sg13g2_decap_8 FILLER_12_184 ();
 sg13g2_fill_2 FILLER_12_191 ();
 sg13g2_fill_2 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_222 ();
 sg13g2_decap_4 FILLER_12_229 ();
 sg13g2_fill_2 FILLER_12_233 ();
 sg13g2_decap_4 FILLER_12_245 ();
 sg13g2_fill_2 FILLER_12_249 ();
 sg13g2_fill_1 FILLER_12_260 ();
 sg13g2_decap_4 FILLER_12_269 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_fill_2 FILLER_12_298 ();
 sg13g2_fill_1 FILLER_12_300 ();
 sg13g2_decap_8 FILLER_12_306 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_348 ();
 sg13g2_decap_8 FILLER_12_355 ();
 sg13g2_decap_8 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_369 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_fill_2 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_58 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_decap_4 FILLER_13_98 ();
 sg13g2_fill_1 FILLER_13_102 ();
 sg13g2_decap_4 FILLER_13_114 ();
 sg13g2_fill_2 FILLER_13_122 ();
 sg13g2_fill_1 FILLER_13_124 ();
 sg13g2_decap_8 FILLER_13_138 ();
 sg13g2_decap_4 FILLER_13_145 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_decap_8 FILLER_13_160 ();
 sg13g2_decap_8 FILLER_13_167 ();
 sg13g2_decap_8 FILLER_13_174 ();
 sg13g2_fill_2 FILLER_13_191 ();
 sg13g2_fill_1 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_220 ();
 sg13g2_decap_8 FILLER_13_227 ();
 sg13g2_decap_8 FILLER_13_234 ();
 sg13g2_fill_2 FILLER_13_241 ();
 sg13g2_fill_1 FILLER_13_243 ();
 sg13g2_fill_2 FILLER_13_256 ();
 sg13g2_fill_1 FILLER_13_258 ();
 sg13g2_decap_4 FILLER_13_270 ();
 sg13g2_fill_2 FILLER_13_274 ();
 sg13g2_fill_2 FILLER_13_281 ();
 sg13g2_fill_1 FILLER_13_283 ();
 sg13g2_decap_4 FILLER_13_288 ();
 sg13g2_fill_2 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_320 ();
 sg13g2_decap_8 FILLER_13_327 ();
 sg13g2_decap_8 FILLER_13_334 ();
 sg13g2_decap_8 FILLER_13_341 ();
 sg13g2_decap_8 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_fill_2 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_87 ();
 sg13g2_decap_8 FILLER_14_97 ();
 sg13g2_fill_2 FILLER_14_104 ();
 sg13g2_fill_1 FILLER_14_106 ();
 sg13g2_decap_8 FILLER_14_117 ();
 sg13g2_decap_8 FILLER_14_124 ();
 sg13g2_fill_1 FILLER_14_131 ();
 sg13g2_decap_4 FILLER_14_137 ();
 sg13g2_decap_4 FILLER_14_146 ();
 sg13g2_fill_2 FILLER_14_150 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_fill_2 FILLER_14_168 ();
 sg13g2_decap_4 FILLER_14_204 ();
 sg13g2_fill_2 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_218 ();
 sg13g2_decap_8 FILLER_14_225 ();
 sg13g2_decap_8 FILLER_14_232 ();
 sg13g2_decap_8 FILLER_14_239 ();
 sg13g2_fill_2 FILLER_14_246 ();
 sg13g2_fill_1 FILLER_14_248 ();
 sg13g2_decap_8 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_265 ();
 sg13g2_fill_1 FILLER_14_272 ();
 sg13g2_fill_2 FILLER_14_282 ();
 sg13g2_fill_2 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_328 ();
 sg13g2_decap_8 FILLER_14_335 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_356 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_4 FILLER_15_56 ();
 sg13g2_fill_2 FILLER_15_60 ();
 sg13g2_fill_2 FILLER_15_66 ();
 sg13g2_fill_1 FILLER_15_68 ();
 sg13g2_fill_1 FILLER_15_95 ();
 sg13g2_decap_4 FILLER_15_117 ();
 sg13g2_fill_2 FILLER_15_121 ();
 sg13g2_decap_8 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_135 ();
 sg13g2_decap_8 FILLER_15_141 ();
 sg13g2_decap_8 FILLER_15_148 ();
 sg13g2_fill_1 FILLER_15_155 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_172 ();
 sg13g2_decap_4 FILLER_15_195 ();
 sg13g2_fill_1 FILLER_15_199 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_fill_2 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_233 ();
 sg13g2_fill_2 FILLER_15_245 ();
 sg13g2_fill_1 FILLER_15_247 ();
 sg13g2_fill_1 FILLER_15_273 ();
 sg13g2_fill_2 FILLER_15_295 ();
 sg13g2_fill_1 FILLER_15_297 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_64 ();
 sg13g2_decap_8 FILLER_16_71 ();
 sg13g2_fill_2 FILLER_16_78 ();
 sg13g2_fill_1 FILLER_16_118 ();
 sg13g2_fill_2 FILLER_16_124 ();
 sg13g2_fill_1 FILLER_16_126 ();
 sg13g2_fill_2 FILLER_16_148 ();
 sg13g2_fill_1 FILLER_16_160 ();
 sg13g2_fill_1 FILLER_16_171 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_4 FILLER_16_196 ();
 sg13g2_fill_2 FILLER_16_226 ();
 sg13g2_fill_1 FILLER_16_228 ();
 sg13g2_decap_4 FILLER_16_247 ();
 sg13g2_fill_2 FILLER_16_251 ();
 sg13g2_fill_2 FILLER_16_278 ();
 sg13g2_fill_1 FILLER_16_280 ();
 sg13g2_fill_2 FILLER_16_289 ();
 sg13g2_fill_1 FILLER_16_291 ();
 sg13g2_fill_2 FILLER_16_302 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_4 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_74 ();
 sg13g2_fill_1 FILLER_17_81 ();
 sg13g2_decap_8 FILLER_17_184 ();
 sg13g2_decap_8 FILLER_17_191 ();
 sg13g2_decap_4 FILLER_17_225 ();
 sg13g2_fill_2 FILLER_17_229 ();
 sg13g2_decap_8 FILLER_17_235 ();
 sg13g2_decap_8 FILLER_17_242 ();
 sg13g2_decap_4 FILLER_17_249 ();
 sg13g2_fill_1 FILLER_17_253 ();
 sg13g2_fill_2 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_decap_8 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_340 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_35 ();
 sg13g2_fill_1 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_75 ();
 sg13g2_decap_8 FILLER_18_82 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_fill_1 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_100 ();
 sg13g2_fill_1 FILLER_18_107 ();
 sg13g2_fill_2 FILLER_18_116 ();
 sg13g2_fill_2 FILLER_18_128 ();
 sg13g2_fill_1 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_239 ();
 sg13g2_fill_1 FILLER_18_246 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_4 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_decap_8 FILLER_18_282 ();
 sg13g2_decap_4 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_320 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_fill_1 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_64 ();
 sg13g2_decap_8 FILLER_19_94 ();
 sg13g2_decap_8 FILLER_19_101 ();
 sg13g2_decap_8 FILLER_19_108 ();
 sg13g2_decap_8 FILLER_19_115 ();
 sg13g2_decap_8 FILLER_19_122 ();
 sg13g2_fill_1 FILLER_19_129 ();
 sg13g2_decap_4 FILLER_19_144 ();
 sg13g2_fill_1 FILLER_19_148 ();
 sg13g2_decap_8 FILLER_19_162 ();
 sg13g2_decap_8 FILLER_19_219 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_decap_8 FILLER_19_253 ();
 sg13g2_fill_2 FILLER_19_260 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_337 ();
 sg13g2_decap_8 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_8 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_4 FILLER_20_49 ();
 sg13g2_fill_1 FILLER_20_53 ();
 sg13g2_fill_2 FILLER_20_80 ();
 sg13g2_fill_1 FILLER_20_82 ();
 sg13g2_decap_8 FILLER_20_128 ();
 sg13g2_decap_8 FILLER_20_135 ();
 sg13g2_decap_8 FILLER_20_142 ();
 sg13g2_decap_8 FILLER_20_149 ();
 sg13g2_decap_4 FILLER_20_156 ();
 sg13g2_fill_1 FILLER_20_160 ();
 sg13g2_decap_4 FILLER_20_166 ();
 sg13g2_fill_1 FILLER_20_170 ();
 sg13g2_decap_8 FILLER_20_191 ();
 sg13g2_fill_2 FILLER_20_198 ();
 sg13g2_decap_8 FILLER_20_209 ();
 sg13g2_decap_4 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_220 ();
 sg13g2_decap_8 FILLER_20_261 ();
 sg13g2_decap_8 FILLER_20_268 ();
 sg13g2_decap_8 FILLER_20_279 ();
 sg13g2_decap_4 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_324 ();
 sg13g2_decap_8 FILLER_20_331 ();
 sg13g2_decap_8 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_345 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_66 ();
 sg13g2_fill_1 FILLER_21_68 ();
 sg13g2_fill_1 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_124 ();
 sg13g2_fill_2 FILLER_21_131 ();
 sg13g2_decap_8 FILLER_21_138 ();
 sg13g2_decap_4 FILLER_21_145 ();
 sg13g2_fill_2 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_164 ();
 sg13g2_decap_8 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_181 ();
 sg13g2_decap_8 FILLER_21_218 ();
 sg13g2_decap_4 FILLER_21_225 ();
 sg13g2_fill_2 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_242 ();
 sg13g2_fill_2 FILLER_21_249 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_fill_2 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_265 ();
 sg13g2_fill_2 FILLER_21_271 ();
 sg13g2_fill_2 FILLER_21_289 ();
 sg13g2_fill_1 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_296 ();
 sg13g2_decap_4 FILLER_21_303 ();
 sg13g2_fill_2 FILLER_21_307 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_fill_2 FILLER_22_49 ();
 sg13g2_fill_1 FILLER_22_51 ();
 sg13g2_fill_2 FILLER_22_71 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_fill_2 FILLER_22_123 ();
 sg13g2_fill_2 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_188 ();
 sg13g2_decap_4 FILLER_22_199 ();
 sg13g2_decap_8 FILLER_22_211 ();
 sg13g2_decap_8 FILLER_22_218 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_fill_2 FILLER_22_241 ();
 sg13g2_fill_2 FILLER_22_263 ();
 sg13g2_decap_4 FILLER_22_305 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_decap_8 FILLER_22_316 ();
 sg13g2_decap_8 FILLER_22_323 ();
 sg13g2_decap_8 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_90 ();
 sg13g2_fill_1 FILLER_23_92 ();
 sg13g2_fill_1 FILLER_23_114 ();
 sg13g2_fill_2 FILLER_23_151 ();
 sg13g2_fill_1 FILLER_23_153 ();
 sg13g2_fill_1 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_219 ();
 sg13g2_decap_4 FILLER_23_226 ();
 sg13g2_fill_1 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_241 ();
 sg13g2_fill_2 FILLER_23_256 ();
 sg13g2_fill_1 FILLER_23_258 ();
 sg13g2_fill_2 FILLER_23_283 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_61 ();
 sg13g2_fill_1 FILLER_24_93 ();
 sg13g2_fill_2 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_143 ();
 sg13g2_fill_1 FILLER_24_160 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_204 ();
 sg13g2_decap_4 FILLER_24_216 ();
 sg13g2_decap_8 FILLER_24_223 ();
 sg13g2_decap_8 FILLER_24_230 ();
 sg13g2_decap_4 FILLER_24_237 ();
 sg13g2_decap_8 FILLER_24_246 ();
 sg13g2_fill_2 FILLER_24_253 ();
 sg13g2_fill_1 FILLER_24_255 ();
 sg13g2_fill_2 FILLER_24_302 ();
 sg13g2_fill_1 FILLER_24_304 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_4 FILLER_25_28 ();
 sg13g2_fill_2 FILLER_25_32 ();
 sg13g2_fill_2 FILLER_25_83 ();
 sg13g2_decap_8 FILLER_25_159 ();
 sg13g2_decap_4 FILLER_25_166 ();
 sg13g2_fill_2 FILLER_25_175 ();
 sg13g2_fill_1 FILLER_25_177 ();
 sg13g2_fill_2 FILLER_25_191 ();
 sg13g2_fill_1 FILLER_25_193 ();
 sg13g2_fill_2 FILLER_25_229 ();
 sg13g2_decap_4 FILLER_25_236 ();
 sg13g2_fill_2 FILLER_25_240 ();
 sg13g2_decap_8 FILLER_25_255 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_decap_4 FILLER_25_271 ();
 sg13g2_fill_2 FILLER_25_275 ();
 sg13g2_fill_2 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_85 ();
 sg13g2_decap_4 FILLER_26_92 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_fill_2 FILLER_26_116 ();
 sg13g2_fill_2 FILLER_26_156 ();
 sg13g2_fill_1 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_164 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_decap_8 FILLER_26_187 ();
 sg13g2_fill_2 FILLER_26_194 ();
 sg13g2_fill_2 FILLER_26_232 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_fill_2 FILLER_26_241 ();
 sg13g2_fill_1 FILLER_26_243 ();
 sg13g2_decap_8 FILLER_26_264 ();
 sg13g2_decap_8 FILLER_26_271 ();
 sg13g2_decap_8 FILLER_26_278 ();
 sg13g2_decap_8 FILLER_26_285 ();
 sg13g2_decap_8 FILLER_26_292 ();
 sg13g2_decap_8 FILLER_26_299 ();
 sg13g2_decap_4 FILLER_26_306 ();
 sg13g2_fill_2 FILLER_26_310 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_8 FILLER_26_323 ();
 sg13g2_decap_4 FILLER_26_330 ();
 sg13g2_fill_1 FILLER_26_334 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_37 ();
 sg13g2_decap_4 FILLER_27_48 ();
 sg13g2_fill_2 FILLER_27_52 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_4 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_84 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_fill_1 FILLER_27_176 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_decap_4 FILLER_27_212 ();
 sg13g2_fill_1 FILLER_27_229 ();
 sg13g2_decap_4 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_decap_4 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_decap_8 FILLER_27_276 ();
 sg13g2_decap_8 FILLER_27_283 ();
 sg13g2_decap_8 FILLER_27_290 ();
 sg13g2_decap_8 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_66 ();
 sg13g2_fill_2 FILLER_28_94 ();
 sg13g2_fill_2 FILLER_28_100 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_fill_2 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_decap_4 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_219 ();
 sg13g2_decap_8 FILLER_28_226 ();
 sg13g2_fill_2 FILLER_28_233 ();
 sg13g2_fill_1 FILLER_28_246 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_fill_2 FILLER_28_297 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_decap_4 FILLER_28_342 ();
 sg13g2_fill_2 FILLER_28_350 ();
 sg13g2_fill_1 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_14 ();
 sg13g2_fill_2 FILLER_29_41 ();
 sg13g2_decap_4 FILLER_29_69 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_decap_8 FILLER_29_87 ();
 sg13g2_decap_8 FILLER_29_94 ();
 sg13g2_decap_8 FILLER_29_101 ();
 sg13g2_decap_4 FILLER_29_108 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_fill_2 FILLER_29_122 ();
 sg13g2_decap_8 FILLER_29_132 ();
 sg13g2_decap_4 FILLER_29_139 ();
 sg13g2_fill_1 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_168 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_fill_2 FILLER_29_189 ();
 sg13g2_fill_2 FILLER_29_199 ();
 sg13g2_fill_1 FILLER_29_201 ();
 sg13g2_decap_4 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_253 ();
 sg13g2_decap_8 FILLER_29_260 ();
 sg13g2_fill_2 FILLER_29_267 ();
 sg13g2_decap_4 FILLER_29_274 ();
 sg13g2_fill_2 FILLER_29_278 ();
 sg13g2_fill_2 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_318 ();
 sg13g2_fill_2 FILLER_29_325 ();
 sg13g2_fill_1 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_335 ();
 sg13g2_decap_8 FILLER_29_342 ();
 sg13g2_decap_8 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_363 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_36 ();
 sg13g2_fill_2 FILLER_30_50 ();
 sg13g2_fill_1 FILLER_30_66 ();
 sg13g2_decap_8 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_89 ();
 sg13g2_decap_8 FILLER_30_103 ();
 sg13g2_decap_8 FILLER_30_110 ();
 sg13g2_decap_4 FILLER_30_117 ();
 sg13g2_decap_8 FILLER_30_135 ();
 sg13g2_fill_2 FILLER_30_142 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_fill_1 FILLER_30_155 ();
 sg13g2_decap_8 FILLER_30_164 ();
 sg13g2_fill_1 FILLER_30_171 ();
 sg13g2_decap_8 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_201 ();
 sg13g2_fill_1 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_decap_8 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_decap_8 FILLER_30_276 ();
 sg13g2_fill_1 FILLER_30_283 ();
 sg13g2_decap_8 FILLER_30_304 ();
 sg13g2_decap_4 FILLER_30_311 ();
 sg13g2_fill_2 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_320 ();
 sg13g2_fill_2 FILLER_30_324 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_11 ();
 sg13g2_decap_4 FILLER_31_112 ();
 sg13g2_fill_2 FILLER_31_116 ();
 sg13g2_fill_2 FILLER_31_158 ();
 sg13g2_fill_1 FILLER_31_165 ();
 sg13g2_decap_4 FILLER_31_197 ();
 sg13g2_fill_2 FILLER_31_211 ();
 sg13g2_fill_2 FILLER_31_230 ();
 sg13g2_decap_8 FILLER_31_265 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_decap_8 FILLER_31_279 ();
 sg13g2_decap_4 FILLER_31_286 ();
 sg13g2_fill_2 FILLER_31_290 ();
 sg13g2_fill_2 FILLER_31_303 ();
 sg13g2_fill_1 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_311 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_decap_8 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_379 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_393 ();
 sg13g2_decap_8 FILLER_31_400 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_28 ();
 sg13g2_fill_2 FILLER_32_32 ();
 sg13g2_decap_8 FILLER_32_43 ();
 sg13g2_decap_8 FILLER_32_59 ();
 sg13g2_fill_2 FILLER_32_66 ();
 sg13g2_decap_8 FILLER_32_86 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_112 ();
 sg13g2_fill_1 FILLER_32_141 ();
 sg13g2_fill_1 FILLER_32_149 ();
 sg13g2_decap_4 FILLER_32_158 ();
 sg13g2_decap_4 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_fill_2 FILLER_32_186 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_decap_4 FILLER_32_194 ();
 sg13g2_fill_2 FILLER_32_198 ();
 sg13g2_fill_2 FILLER_32_226 ();
 sg13g2_decap_4 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_fill_2 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_281 ();
 sg13g2_fill_2 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_383 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_4 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_39 ();
 sg13g2_decap_4 FILLER_33_80 ();
 sg13g2_decap_8 FILLER_33_99 ();
 sg13g2_fill_1 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_121 ();
 sg13g2_fill_2 FILLER_33_167 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_214 ();
 sg13g2_decap_4 FILLER_33_221 ();
 sg13g2_decap_8 FILLER_33_230 ();
 sg13g2_decap_8 FILLER_33_237 ();
 sg13g2_decap_4 FILLER_33_244 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_decap_8 FILLER_33_254 ();
 sg13g2_decap_4 FILLER_33_283 ();
 sg13g2_fill_2 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_347 ();
 sg13g2_fill_2 FILLER_33_353 ();
 sg13g2_fill_1 FILLER_33_355 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_21 ();
 sg13g2_fill_1 FILLER_34_48 ();
 sg13g2_fill_1 FILLER_34_75 ();
 sg13g2_fill_2 FILLER_34_86 ();
 sg13g2_decap_8 FILLER_34_93 ();
 sg13g2_decap_8 FILLER_34_100 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_decap_4 FILLER_34_120 ();
 sg13g2_fill_1 FILLER_34_124 ();
 sg13g2_fill_2 FILLER_34_129 ();
 sg13g2_fill_1 FILLER_34_131 ();
 sg13g2_decap_8 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_143 ();
 sg13g2_decap_8 FILLER_34_155 ();
 sg13g2_fill_2 FILLER_34_162 ();
 sg13g2_fill_2 FILLER_34_178 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_4 FILLER_34_222 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_fill_1 FILLER_34_238 ();
 sg13g2_fill_1 FILLER_34_313 ();
 sg13g2_decap_8 FILLER_34_341 ();
 sg13g2_decap_8 FILLER_34_348 ();
 sg13g2_decap_4 FILLER_34_355 ();
 sg13g2_fill_2 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_370 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_34 ();
 sg13g2_fill_2 FILLER_35_61 ();
 sg13g2_decap_4 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_81 ();
 sg13g2_decap_8 FILLER_35_87 ();
 sg13g2_decap_8 FILLER_35_94 ();
 sg13g2_decap_4 FILLER_35_101 ();
 sg13g2_fill_2 FILLER_35_113 ();
 sg13g2_decap_4 FILLER_35_125 ();
 sg13g2_fill_1 FILLER_35_129 ();
 sg13g2_fill_1 FILLER_35_139 ();
 sg13g2_decap_4 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_fill_2 FILLER_35_165 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_fill_1 FILLER_35_180 ();
 sg13g2_decap_4 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_255 ();
 sg13g2_fill_1 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_269 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_2 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_318 ();
 sg13g2_fill_2 FILLER_35_329 ();
 sg13g2_decap_4 FILLER_35_334 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_fill_2 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_43 ();
 sg13g2_fill_2 FILLER_36_58 ();
 sg13g2_fill_1 FILLER_36_60 ();
 sg13g2_decap_4 FILLER_36_69 ();
 sg13g2_fill_1 FILLER_36_73 ();
 sg13g2_fill_1 FILLER_36_115 ();
 sg13g2_fill_2 FILLER_36_153 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_decap_4 FILLER_36_179 ();
 sg13g2_decap_4 FILLER_36_188 ();
 sg13g2_fill_1 FILLER_36_204 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_246 ();
 sg13g2_decap_8 FILLER_36_253 ();
 sg13g2_decap_8 FILLER_36_260 ();
 sg13g2_decap_8 FILLER_36_267 ();
 sg13g2_fill_2 FILLER_36_274 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_decap_4 FILLER_36_283 ();
 sg13g2_decap_8 FILLER_36_291 ();
 sg13g2_decap_4 FILLER_36_298 ();
 sg13g2_fill_1 FILLER_36_302 ();
 sg13g2_fill_2 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_350 ();
 sg13g2_fill_1 FILLER_36_356 ();
 sg13g2_fill_2 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_393 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_decap_8 FILLER_37_66 ();
 sg13g2_fill_1 FILLER_37_73 ();
 sg13g2_fill_2 FILLER_37_82 ();
 sg13g2_fill_1 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_146 ();
 sg13g2_fill_2 FILLER_37_161 ();
 sg13g2_fill_1 FILLER_37_163 ();
 sg13g2_decap_4 FILLER_37_225 ();
 sg13g2_decap_8 FILLER_37_233 ();
 sg13g2_decap_8 FILLER_37_240 ();
 sg13g2_decap_8 FILLER_37_247 ();
 sg13g2_decap_8 FILLER_37_254 ();
 sg13g2_decap_8 FILLER_37_261 ();
 sg13g2_decap_8 FILLER_37_302 ();
 sg13g2_decap_8 FILLER_37_309 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_fill_2 FILLER_37_323 ();
 sg13g2_fill_1 FILLER_37_325 ();
 sg13g2_decap_8 FILLER_37_330 ();
 sg13g2_decap_4 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_11 ();
 sg13g2_decap_8 FILLER_38_17 ();
 sg13g2_decap_4 FILLER_38_24 ();
 sg13g2_decap_4 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_67 ();
 sg13g2_decap_4 FILLER_38_74 ();
 sg13g2_fill_2 FILLER_38_83 ();
 sg13g2_fill_2 FILLER_38_94 ();
 sg13g2_fill_2 FILLER_38_121 ();
 sg13g2_fill_1 FILLER_38_131 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_153 ();
 sg13g2_fill_2 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_decap_4 FILLER_38_234 ();
 sg13g2_fill_2 FILLER_38_238 ();
 sg13g2_fill_1 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_268 ();
 sg13g2_fill_2 FILLER_38_275 ();
 sg13g2_decap_8 FILLER_38_293 ();
 sg13g2_decap_4 FILLER_38_300 ();
 sg13g2_fill_2 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_309 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_324 ();
 sg13g2_fill_2 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_fill_1 FILLER_39_35 ();
 sg13g2_fill_1 FILLER_39_96 ();
 sg13g2_decap_4 FILLER_39_107 ();
 sg13g2_fill_2 FILLER_39_131 ();
 sg13g2_decap_8 FILLER_39_162 ();
 sg13g2_fill_2 FILLER_39_169 ();
 sg13g2_fill_1 FILLER_39_171 ();
 sg13g2_decap_8 FILLER_39_195 ();
 sg13g2_decap_8 FILLER_39_202 ();
 sg13g2_decap_8 FILLER_39_209 ();
 sg13g2_decap_4 FILLER_39_216 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_fill_2 FILLER_39_231 ();
 sg13g2_fill_1 FILLER_39_233 ();
 sg13g2_fill_2 FILLER_39_270 ();
 sg13g2_fill_1 FILLER_39_272 ();
 sg13g2_decap_4 FILLER_39_284 ();
 sg13g2_fill_2 FILLER_39_288 ();
 sg13g2_fill_1 FILLER_39_294 ();
 sg13g2_fill_2 FILLER_39_316 ();
 sg13g2_fill_1 FILLER_39_328 ();
 sg13g2_fill_2 FILLER_39_362 ();
 sg13g2_fill_2 FILLER_39_369 ();
 sg13g2_fill_1 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_384 ();
 sg13g2_decap_8 FILLER_39_391 ();
 sg13g2_decap_8 FILLER_39_398 ();
 sg13g2_decap_4 FILLER_39_405 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_9 ();
 sg13g2_decap_8 FILLER_40_36 ();
 sg13g2_fill_1 FILLER_40_43 ();
 sg13g2_fill_2 FILLER_40_54 ();
 sg13g2_fill_2 FILLER_40_69 ();
 sg13g2_fill_1 FILLER_40_71 ();
 sg13g2_decap_4 FILLER_40_90 ();
 sg13g2_fill_1 FILLER_40_94 ();
 sg13g2_decap_8 FILLER_40_121 ();
 sg13g2_decap_4 FILLER_40_128 ();
 sg13g2_fill_2 FILLER_40_132 ();
 sg13g2_fill_2 FILLER_40_196 ();
 sg13g2_fill_1 FILLER_40_198 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_fill_2 FILLER_40_231 ();
 sg13g2_decap_4 FILLER_40_237 ();
 sg13g2_fill_2 FILLER_40_250 ();
 sg13g2_fill_2 FILLER_40_262 ();
 sg13g2_decap_4 FILLER_40_281 ();
 sg13g2_fill_2 FILLER_40_346 ();
 sg13g2_decap_8 FILLER_40_356 ();
 sg13g2_decap_8 FILLER_40_363 ();
 sg13g2_decap_8 FILLER_40_374 ();
 sg13g2_decap_8 FILLER_40_381 ();
 sg13g2_decap_8 FILLER_40_388 ();
 sg13g2_decap_8 FILLER_40_395 ();
 sg13g2_decap_8 FILLER_40_402 ();
 sg13g2_decap_4 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_4 ();
 sg13g2_fill_2 FILLER_41_41 ();
 sg13g2_fill_1 FILLER_41_43 ();
 sg13g2_fill_1 FILLER_41_53 ();
 sg13g2_fill_2 FILLER_41_63 ();
 sg13g2_fill_1 FILLER_41_65 ();
 sg13g2_fill_2 FILLER_41_74 ();
 sg13g2_decap_8 FILLER_41_80 ();
 sg13g2_decap_8 FILLER_41_87 ();
 sg13g2_decap_8 FILLER_41_94 ();
 sg13g2_decap_4 FILLER_41_101 ();
 sg13g2_fill_1 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_110 ();
 sg13g2_decap_8 FILLER_41_117 ();
 sg13g2_decap_8 FILLER_41_124 ();
 sg13g2_fill_2 FILLER_41_131 ();
 sg13g2_decap_8 FILLER_41_146 ();
 sg13g2_fill_2 FILLER_41_153 ();
 sg13g2_decap_8 FILLER_41_159 ();
 sg13g2_decap_8 FILLER_41_166 ();
 sg13g2_fill_1 FILLER_41_173 ();
 sg13g2_fill_1 FILLER_41_188 ();
 sg13g2_fill_1 FILLER_41_227 ();
 sg13g2_fill_2 FILLER_41_242 ();
 sg13g2_fill_2 FILLER_41_258 ();
 sg13g2_fill_1 FILLER_41_265 ();
 sg13g2_decap_8 FILLER_41_274 ();
 sg13g2_decap_8 FILLER_41_281 ();
 sg13g2_decap_4 FILLER_41_288 ();
 sg13g2_fill_1 FILLER_41_292 ();
 sg13g2_fill_1 FILLER_41_297 ();
 sg13g2_decap_4 FILLER_41_315 ();
 sg13g2_fill_1 FILLER_41_319 ();
 sg13g2_fill_1 FILLER_41_330 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_fill_2 FILLER_41_356 ();
 sg13g2_fill_1 FILLER_41_358 ();
 sg13g2_decap_4 FILLER_41_367 ();
 sg13g2_fill_2 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_fill_2 FILLER_42_14 ();
 sg13g2_fill_1 FILLER_42_16 ();
 sg13g2_fill_1 FILLER_42_21 ();
 sg13g2_fill_2 FILLER_42_68 ();
 sg13g2_fill_1 FILLER_42_74 ();
 sg13g2_decap_8 FILLER_42_83 ();
 sg13g2_decap_8 FILLER_42_90 ();
 sg13g2_fill_2 FILLER_42_97 ();
 sg13g2_decap_8 FILLER_42_107 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_fill_1 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_170 ();
 sg13g2_decap_4 FILLER_42_177 ();
 sg13g2_decap_4 FILLER_42_189 ();
 sg13g2_decap_4 FILLER_42_253 ();
 sg13g2_decap_8 FILLER_42_277 ();
 sg13g2_fill_1 FILLER_42_284 ();
 sg13g2_decap_8 FILLER_42_289 ();
 sg13g2_fill_2 FILLER_42_296 ();
 sg13g2_fill_1 FILLER_42_298 ();
 sg13g2_decap_8 FILLER_42_302 ();
 sg13g2_fill_2 FILLER_42_309 ();
 sg13g2_decap_4 FILLER_42_322 ();
 sg13g2_fill_1 FILLER_42_326 ();
 sg13g2_decap_4 FILLER_42_352 ();
 sg13g2_fill_1 FILLER_42_364 ();
 sg13g2_fill_2 FILLER_42_370 ();
 sg13g2_decap_8 FILLER_42_384 ();
 sg13g2_decap_8 FILLER_42_391 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_decap_4 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_4 FILLER_43_21 ();
 sg13g2_fill_1 FILLER_43_25 ();
 sg13g2_decap_4 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_177 ();
 sg13g2_decap_8 FILLER_43_184 ();
 sg13g2_decap_8 FILLER_43_191 ();
 sg13g2_fill_2 FILLER_43_198 ();
 sg13g2_fill_2 FILLER_43_207 ();
 sg13g2_decap_4 FILLER_43_268 ();
 sg13g2_decap_4 FILLER_43_303 ();
 sg13g2_fill_1 FILLER_43_307 ();
 sg13g2_decap_8 FILLER_43_311 ();
 sg13g2_decap_8 FILLER_43_318 ();
 sg13g2_decap_8 FILLER_43_325 ();
 sg13g2_fill_1 FILLER_43_340 ();
 sg13g2_fill_1 FILLER_43_347 ();
 sg13g2_fill_2 FILLER_43_363 ();
 sg13g2_fill_1 FILLER_43_370 ();
 sg13g2_decap_8 FILLER_43_382 ();
 sg13g2_decap_8 FILLER_43_389 ();
 sg13g2_decap_8 FILLER_43_396 ();
 sg13g2_decap_4 FILLER_43_403 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_fill_1 FILLER_44_35 ();
 sg13g2_fill_1 FILLER_44_56 ();
 sg13g2_fill_2 FILLER_44_82 ();
 sg13g2_fill_2 FILLER_44_97 ();
 sg13g2_decap_8 FILLER_44_107 ();
 sg13g2_fill_1 FILLER_44_124 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_fill_2 FILLER_44_161 ();
 sg13g2_fill_2 FILLER_44_174 ();
 sg13g2_decap_4 FILLER_44_182 ();
 sg13g2_fill_1 FILLER_44_192 ();
 sg13g2_decap_8 FILLER_44_206 ();
 sg13g2_decap_4 FILLER_44_213 ();
 sg13g2_fill_1 FILLER_44_217 ();
 sg13g2_fill_2 FILLER_44_228 ();
 sg13g2_decap_8 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_fill_2 FILLER_44_273 ();
 sg13g2_fill_2 FILLER_44_279 ();
 sg13g2_fill_1 FILLER_44_281 ();
 sg13g2_decap_4 FILLER_44_286 ();
 sg13g2_fill_1 FILLER_44_290 ();
 sg13g2_decap_8 FILLER_44_319 ();
 sg13g2_decap_8 FILLER_44_326 ();
 sg13g2_decap_4 FILLER_44_333 ();
 sg13g2_fill_2 FILLER_44_349 ();
 sg13g2_fill_1 FILLER_44_351 ();
 sg13g2_fill_2 FILLER_44_359 ();
 sg13g2_fill_1 FILLER_44_361 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_4 FILLER_45_28 ();
 sg13g2_decap_4 FILLER_45_48 ();
 sg13g2_fill_1 FILLER_45_52 ();
 sg13g2_decap_8 FILLER_45_57 ();
 sg13g2_decap_4 FILLER_45_73 ();
 sg13g2_decap_8 FILLER_45_87 ();
 sg13g2_fill_2 FILLER_45_94 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_fill_2 FILLER_45_119 ();
 sg13g2_fill_1 FILLER_45_121 ();
 sg13g2_fill_2 FILLER_45_147 ();
 sg13g2_fill_1 FILLER_45_149 ();
 sg13g2_decap_4 FILLER_45_155 ();
 sg13g2_fill_1 FILLER_45_171 ();
 sg13g2_decap_8 FILLER_45_214 ();
 sg13g2_fill_2 FILLER_45_221 ();
 sg13g2_decap_8 FILLER_45_247 ();
 sg13g2_fill_2 FILLER_45_254 ();
 sg13g2_decap_8 FILLER_45_333 ();
 sg13g2_fill_2 FILLER_45_340 ();
 sg13g2_fill_1 FILLER_45_342 ();
 sg13g2_decap_8 FILLER_45_352 ();
 sg13g2_fill_1 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_fill_2 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_46 ();
 sg13g2_fill_1 FILLER_46_50 ();
 sg13g2_decap_8 FILLER_46_65 ();
 sg13g2_decap_8 FILLER_46_72 ();
 sg13g2_decap_8 FILLER_46_79 ();
 sg13g2_decap_4 FILLER_46_86 ();
 sg13g2_fill_2 FILLER_46_90 ();
 sg13g2_decap_8 FILLER_46_110 ();
 sg13g2_decap_8 FILLER_46_122 ();
 sg13g2_decap_4 FILLER_46_129 ();
 sg13g2_fill_1 FILLER_46_133 ();
 sg13g2_decap_4 FILLER_46_144 ();
 sg13g2_fill_2 FILLER_46_148 ();
 sg13g2_fill_2 FILLER_46_156 ();
 sg13g2_fill_1 FILLER_46_170 ();
 sg13g2_fill_2 FILLER_46_175 ();
 sg13g2_fill_1 FILLER_46_177 ();
 sg13g2_fill_1 FILLER_46_188 ();
 sg13g2_decap_8 FILLER_46_220 ();
 sg13g2_decap_8 FILLER_46_227 ();
 sg13g2_fill_2 FILLER_46_234 ();
 sg13g2_decap_8 FILLER_46_239 ();
 sg13g2_decap_4 FILLER_46_246 ();
 sg13g2_fill_2 FILLER_46_250 ();
 sg13g2_decap_8 FILLER_46_257 ();
 sg13g2_decap_8 FILLER_46_264 ();
 sg13g2_decap_8 FILLER_46_271 ();
 sg13g2_fill_2 FILLER_46_278 ();
 sg13g2_fill_1 FILLER_46_280 ();
 sg13g2_fill_2 FILLER_46_296 ();
 sg13g2_fill_1 FILLER_46_298 ();
 sg13g2_fill_2 FILLER_46_314 ();
 sg13g2_fill_2 FILLER_46_326 ();
 sg13g2_fill_2 FILLER_46_362 ();
 sg13g2_fill_2 FILLER_46_370 ();
 sg13g2_decap_8 FILLER_46_387 ();
 sg13g2_decap_8 FILLER_46_394 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_9 ();
 sg13g2_decap_8 FILLER_47_62 ();
 sg13g2_fill_2 FILLER_47_69 ();
 sg13g2_fill_1 FILLER_47_80 ();
 sg13g2_decap_8 FILLER_47_93 ();
 sg13g2_fill_2 FILLER_47_100 ();
 sg13g2_fill_1 FILLER_47_102 ();
 sg13g2_fill_1 FILLER_47_113 ();
 sg13g2_decap_4 FILLER_47_157 ();
 sg13g2_fill_2 FILLER_47_161 ();
 sg13g2_decap_4 FILLER_47_176 ();
 sg13g2_fill_1 FILLER_47_180 ();
 sg13g2_fill_2 FILLER_47_194 ();
 sg13g2_decap_8 FILLER_47_222 ();
 sg13g2_decap_8 FILLER_47_229 ();
 sg13g2_fill_2 FILLER_47_236 ();
 sg13g2_fill_1 FILLER_47_242 ();
 sg13g2_decap_4 FILLER_47_248 ();
 sg13g2_fill_2 FILLER_47_282 ();
 sg13g2_decap_8 FILLER_47_300 ();
 sg13g2_decap_8 FILLER_47_307 ();
 sg13g2_fill_1 FILLER_47_324 ();
 sg13g2_decap_4 FILLER_47_336 ();
 sg13g2_fill_1 FILLER_47_340 ();
 sg13g2_fill_1 FILLER_47_346 ();
 sg13g2_decap_8 FILLER_47_353 ();
 sg13g2_fill_2 FILLER_47_360 ();
 sg13g2_decap_8 FILLER_47_376 ();
 sg13g2_decap_8 FILLER_47_383 ();
 sg13g2_decap_8 FILLER_47_390 ();
 sg13g2_decap_8 FILLER_47_397 ();
 sg13g2_decap_4 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_4 FILLER_48_14 ();
 sg13g2_decap_4 FILLER_48_104 ();
 sg13g2_fill_1 FILLER_48_108 ();
 sg13g2_fill_2 FILLER_48_113 ();
 sg13g2_decap_4 FILLER_48_119 ();
 sg13g2_fill_2 FILLER_48_123 ();
 sg13g2_fill_2 FILLER_48_146 ();
 sg13g2_fill_2 FILLER_48_153 ();
 sg13g2_decap_8 FILLER_48_163 ();
 sg13g2_decap_8 FILLER_48_170 ();
 sg13g2_fill_2 FILLER_48_177 ();
 sg13g2_decap_8 FILLER_48_213 ();
 sg13g2_decap_8 FILLER_48_220 ();
 sg13g2_decap_4 FILLER_48_227 ();
 sg13g2_fill_1 FILLER_48_235 ();
 sg13g2_fill_2 FILLER_48_263 ();
 sg13g2_fill_1 FILLER_48_265 ();
 sg13g2_decap_8 FILLER_48_293 ();
 sg13g2_decap_8 FILLER_48_300 ();
 sg13g2_decap_8 FILLER_48_307 ();
 sg13g2_decap_4 FILLER_48_321 ();
 sg13g2_fill_1 FILLER_48_325 ();
 sg13g2_decap_4 FILLER_48_331 ();
 sg13g2_fill_1 FILLER_48_335 ();
 sg13g2_decap_4 FILLER_48_346 ();
 sg13g2_fill_1 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_380 ();
 sg13g2_decap_8 FILLER_48_387 ();
 sg13g2_decap_8 FILLER_48_394 ();
 sg13g2_decap_8 FILLER_48_401 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_4 FILLER_49_28 ();
 sg13g2_fill_1 FILLER_49_32 ();
 sg13g2_fill_2 FILLER_49_42 ();
 sg13g2_fill_1 FILLER_49_44 ();
 sg13g2_decap_4 FILLER_49_97 ();
 sg13g2_fill_2 FILLER_49_106 ();
 sg13g2_fill_1 FILLER_49_108 ();
 sg13g2_fill_2 FILLER_49_144 ();
 sg13g2_fill_2 FILLER_49_153 ();
 sg13g2_fill_1 FILLER_49_155 ();
 sg13g2_decap_4 FILLER_49_161 ();
 sg13g2_decap_4 FILLER_49_171 ();
 sg13g2_fill_2 FILLER_49_175 ();
 sg13g2_decap_4 FILLER_49_182 ();
 sg13g2_fill_1 FILLER_49_186 ();
 sg13g2_decap_8 FILLER_49_201 ();
 sg13g2_decap_8 FILLER_49_208 ();
 sg13g2_decap_8 FILLER_49_215 ();
 sg13g2_decap_4 FILLER_49_222 ();
 sg13g2_fill_2 FILLER_49_226 ();
 sg13g2_fill_2 FILLER_49_236 ();
 sg13g2_fill_1 FILLER_49_238 ();
 sg13g2_fill_2 FILLER_49_247 ();
 sg13g2_fill_1 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_49_270 ();
 sg13g2_fill_1 FILLER_49_277 ();
 sg13g2_decap_4 FILLER_49_286 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_fill_1 FILLER_49_301 ();
 sg13g2_fill_2 FILLER_49_307 ();
 sg13g2_fill_1 FILLER_49_309 ();
 sg13g2_decap_8 FILLER_49_326 ();
 sg13g2_decap_8 FILLER_49_333 ();
 sg13g2_decap_8 FILLER_49_383 ();
 sg13g2_decap_8 FILLER_49_390 ();
 sg13g2_decap_8 FILLER_49_397 ();
 sg13g2_decap_4 FILLER_49_404 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_fill_1 FILLER_50_28 ();
 sg13g2_decap_4 FILLER_50_52 ();
 sg13g2_fill_1 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_64 ();
 sg13g2_fill_1 FILLER_50_71 ();
 sg13g2_decap_4 FILLER_50_75 ();
 sg13g2_fill_2 FILLER_50_79 ();
 sg13g2_fill_2 FILLER_50_89 ();
 sg13g2_fill_1 FILLER_50_91 ();
 sg13g2_decap_4 FILLER_50_125 ();
 sg13g2_decap_4 FILLER_50_133 ();
 sg13g2_fill_1 FILLER_50_137 ();
 sg13g2_fill_1 FILLER_50_141 ();
 sg13g2_fill_2 FILLER_50_151 ();
 sg13g2_fill_1 FILLER_50_153 ();
 sg13g2_fill_2 FILLER_50_175 ();
 sg13g2_fill_1 FILLER_50_177 ();
 sg13g2_decap_8 FILLER_50_197 ();
 sg13g2_fill_2 FILLER_50_209 ();
 sg13g2_decap_4 FILLER_50_216 ();
 sg13g2_fill_1 FILLER_50_220 ();
 sg13g2_decap_4 FILLER_50_226 ();
 sg13g2_fill_2 FILLER_50_288 ();
 sg13g2_decap_4 FILLER_50_305 ();
 sg13g2_decap_8 FILLER_50_335 ();
 sg13g2_decap_4 FILLER_50_342 ();
 sg13g2_fill_2 FILLER_50_346 ();
 sg13g2_fill_2 FILLER_50_362 ();
 sg13g2_fill_1 FILLER_50_364 ();
 sg13g2_decap_8 FILLER_50_374 ();
 sg13g2_decap_8 FILLER_50_381 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_decap_8 FILLER_50_402 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_7 ();
 sg13g2_fill_2 FILLER_51_11 ();
 sg13g2_fill_1 FILLER_51_44 ();
 sg13g2_decap_8 FILLER_51_55 ();
 sg13g2_decap_8 FILLER_51_71 ();
 sg13g2_decap_4 FILLER_51_78 ();
 sg13g2_decap_8 FILLER_51_92 ();
 sg13g2_decap_8 FILLER_51_99 ();
 sg13g2_decap_4 FILLER_51_106 ();
 sg13g2_decap_8 FILLER_51_115 ();
 sg13g2_decap_8 FILLER_51_122 ();
 sg13g2_decap_8 FILLER_51_129 ();
 sg13g2_fill_2 FILLER_51_136 ();
 sg13g2_fill_1 FILLER_51_138 ();
 sg13g2_decap_8 FILLER_51_144 ();
 sg13g2_fill_2 FILLER_51_156 ();
 sg13g2_fill_1 FILLER_51_158 ();
 sg13g2_decap_4 FILLER_51_171 ();
 sg13g2_fill_1 FILLER_51_175 ();
 sg13g2_decap_4 FILLER_51_210 ();
 sg13g2_fill_2 FILLER_51_214 ();
 sg13g2_decap_8 FILLER_51_232 ();
 sg13g2_decap_4 FILLER_51_239 ();
 sg13g2_decap_8 FILLER_51_258 ();
 sg13g2_fill_1 FILLER_51_265 ();
 sg13g2_fill_2 FILLER_51_276 ();
 sg13g2_fill_1 FILLER_51_278 ();
 sg13g2_fill_2 FILLER_51_305 ();
 sg13g2_fill_1 FILLER_51_307 ();
 sg13g2_decap_4 FILLER_51_347 ();
 sg13g2_fill_2 FILLER_51_357 ();
 sg13g2_fill_1 FILLER_51_359 ();
 sg13g2_decap_8 FILLER_51_365 ();
 sg13g2_decap_4 FILLER_51_372 ();
 sg13g2_decap_8 FILLER_51_383 ();
 sg13g2_decap_8 FILLER_51_390 ();
 sg13g2_decap_8 FILLER_51_397 ();
 sg13g2_decap_4 FILLER_51_404 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_14 ();
 sg13g2_fill_1 FILLER_52_16 ();
 sg13g2_fill_1 FILLER_52_47 ();
 sg13g2_fill_1 FILLER_52_74 ();
 sg13g2_fill_1 FILLER_52_78 ();
 sg13g2_fill_1 FILLER_52_92 ();
 sg13g2_decap_8 FILLER_52_109 ();
 sg13g2_fill_1 FILLER_52_116 ();
 sg13g2_decap_8 FILLER_52_128 ();
 sg13g2_fill_2 FILLER_52_151 ();
 sg13g2_fill_1 FILLER_52_153 ();
 sg13g2_decap_4 FILLER_52_159 ();
 sg13g2_decap_8 FILLER_52_170 ();
 sg13g2_decap_4 FILLER_52_177 ();
 sg13g2_fill_1 FILLER_52_186 ();
 sg13g2_fill_2 FILLER_52_191 ();
 sg13g2_fill_2 FILLER_52_206 ();
 sg13g2_fill_1 FILLER_52_208 ();
 sg13g2_fill_2 FILLER_52_220 ();
 sg13g2_fill_1 FILLER_52_222 ();
 sg13g2_fill_2 FILLER_52_229 ();
 sg13g2_fill_1 FILLER_52_239 ();
 sg13g2_decap_8 FILLER_52_266 ();
 sg13g2_decap_8 FILLER_52_273 ();
 sg13g2_fill_2 FILLER_52_285 ();
 sg13g2_fill_2 FILLER_52_297 ();
 sg13g2_fill_1 FILLER_52_304 ();
 sg13g2_decap_8 FILLER_52_308 ();
 sg13g2_fill_1 FILLER_52_315 ();
 sg13g2_decap_4 FILLER_52_324 ();
 sg13g2_fill_1 FILLER_52_328 ();
 sg13g2_fill_2 FILLER_52_335 ();
 sg13g2_fill_1 FILLER_52_337 ();
 sg13g2_fill_2 FILLER_52_344 ();
 sg13g2_fill_1 FILLER_52_346 ();
 sg13g2_fill_2 FILLER_52_375 ();
 sg13g2_fill_1 FILLER_52_377 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_decap_8 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_fill_2 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_72 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_decap_4 FILLER_53_106 ();
 sg13g2_fill_1 FILLER_53_110 ();
 sg13g2_decap_8 FILLER_53_116 ();
 sg13g2_fill_1 FILLER_53_123 ();
 sg13g2_fill_1 FILLER_53_167 ();
 sg13g2_fill_1 FILLER_53_175 ();
 sg13g2_fill_2 FILLER_53_212 ();
 sg13g2_decap_8 FILLER_53_227 ();
 sg13g2_decap_4 FILLER_53_234 ();
 sg13g2_fill_2 FILLER_53_238 ();
 sg13g2_decap_8 FILLER_53_255 ();
 sg13g2_fill_2 FILLER_53_262 ();
 sg13g2_fill_1 FILLER_53_264 ();
 sg13g2_decap_8 FILLER_53_273 ();
 sg13g2_fill_1 FILLER_53_280 ();
 sg13g2_decap_4 FILLER_53_287 ();
 sg13g2_fill_2 FILLER_53_291 ();
 sg13g2_decap_8 FILLER_53_303 ();
 sg13g2_fill_2 FILLER_53_310 ();
 sg13g2_fill_1 FILLER_53_312 ();
 sg13g2_fill_2 FILLER_53_322 ();
 sg13g2_fill_1 FILLER_53_324 ();
 sg13g2_decap_8 FILLER_53_354 ();
 sg13g2_decap_8 FILLER_53_361 ();
 sg13g2_fill_2 FILLER_53_368 ();
 sg13g2_fill_1 FILLER_53_375 ();
 sg13g2_decap_8 FILLER_53_390 ();
 sg13g2_decap_8 FILLER_53_397 ();
 sg13g2_decap_4 FILLER_53_404 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_fill_2 FILLER_54_42 ();
 sg13g2_fill_1 FILLER_54_44 ();
 sg13g2_fill_2 FILLER_54_72 ();
 sg13g2_decap_4 FILLER_54_79 ();
 sg13g2_fill_1 FILLER_54_83 ();
 sg13g2_decap_4 FILLER_54_124 ();
 sg13g2_fill_2 FILLER_54_161 ();
 sg13g2_fill_1 FILLER_54_163 ();
 sg13g2_fill_2 FILLER_54_169 ();
 sg13g2_fill_1 FILLER_54_171 ();
 sg13g2_fill_2 FILLER_54_183 ();
 sg13g2_decap_8 FILLER_54_237 ();
 sg13g2_decap_8 FILLER_54_244 ();
 sg13g2_decap_8 FILLER_54_251 ();
 sg13g2_decap_8 FILLER_54_258 ();
 sg13g2_decap_4 FILLER_54_265 ();
 sg13g2_fill_1 FILLER_54_269 ();
 sg13g2_decap_8 FILLER_54_275 ();
 sg13g2_decap_8 FILLER_54_282 ();
 sg13g2_decap_4 FILLER_54_289 ();
 sg13g2_decap_8 FILLER_54_343 ();
 sg13g2_decap_4 FILLER_54_350 ();
 sg13g2_fill_2 FILLER_54_359 ();
 sg13g2_fill_2 FILLER_54_372 ();
 sg13g2_fill_1 FILLER_54_374 ();
 sg13g2_fill_2 FILLER_54_380 ();
 sg13g2_decap_8 FILLER_54_400 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_4 FILLER_55_28 ();
 sg13g2_fill_2 FILLER_55_32 ();
 sg13g2_decap_8 FILLER_55_47 ();
 sg13g2_decap_8 FILLER_55_54 ();
 sg13g2_fill_1 FILLER_55_61 ();
 sg13g2_decap_8 FILLER_55_79 ();
 sg13g2_fill_1 FILLER_55_137 ();
 sg13g2_decap_4 FILLER_55_145 ();
 sg13g2_fill_1 FILLER_55_149 ();
 sg13g2_decap_8 FILLER_55_176 ();
 sg13g2_fill_1 FILLER_55_183 ();
 sg13g2_decap_8 FILLER_55_205 ();
 sg13g2_decap_4 FILLER_55_212 ();
 sg13g2_fill_1 FILLER_55_216 ();
 sg13g2_decap_8 FILLER_55_226 ();
 sg13g2_decap_8 FILLER_55_245 ();
 sg13g2_fill_1 FILLER_55_252 ();
 sg13g2_decap_8 FILLER_55_288 ();
 sg13g2_decap_4 FILLER_55_299 ();
 sg13g2_fill_1 FILLER_55_303 ();
 sg13g2_decap_8 FILLER_55_320 ();
 sg13g2_decap_8 FILLER_55_327 ();
 sg13g2_fill_1 FILLER_55_334 ();
 sg13g2_fill_2 FILLER_55_345 ();
 sg13g2_fill_2 FILLER_55_371 ();
 sg13g2_fill_1 FILLER_55_373 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_65 ();
 sg13g2_fill_1 FILLER_56_67 ();
 sg13g2_decap_8 FILLER_56_108 ();
 sg13g2_fill_1 FILLER_56_115 ();
 sg13g2_fill_1 FILLER_56_121 ();
 sg13g2_fill_2 FILLER_56_126 ();
 sg13g2_fill_1 FILLER_56_136 ();
 sg13g2_fill_1 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_175 ();
 sg13g2_decap_8 FILLER_56_182 ();
 sg13g2_decap_8 FILLER_56_189 ();
 sg13g2_decap_4 FILLER_56_196 ();
 sg13g2_fill_1 FILLER_56_200 ();
 sg13g2_fill_1 FILLER_56_230 ();
 sg13g2_decap_8 FILLER_56_246 ();
 sg13g2_decap_8 FILLER_56_253 ();
 sg13g2_fill_2 FILLER_56_260 ();
 sg13g2_fill_1 FILLER_56_262 ();
 sg13g2_decap_4 FILLER_56_293 ();
 sg13g2_decap_4 FILLER_56_323 ();
 sg13g2_fill_1 FILLER_56_327 ();
 sg13g2_fill_2 FILLER_56_351 ();
 sg13g2_fill_1 FILLER_56_353 ();
 sg13g2_fill_2 FILLER_56_376 ();
 sg13g2_fill_1 FILLER_56_378 ();
 sg13g2_decap_4 FILLER_56_382 ();
 sg13g2_decap_8 FILLER_56_395 ();
 sg13g2_decap_8 FILLER_56_402 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_fill_2 FILLER_57_21 ();
 sg13g2_fill_1 FILLER_57_23 ();
 sg13g2_decap_4 FILLER_57_51 ();
 sg13g2_decap_8 FILLER_57_101 ();
 sg13g2_decap_8 FILLER_57_108 ();
 sg13g2_decap_8 FILLER_57_115 ();
 sg13g2_decap_8 FILLER_57_122 ();
 sg13g2_fill_2 FILLER_57_129 ();
 sg13g2_fill_1 FILLER_57_131 ();
 sg13g2_fill_1 FILLER_57_139 ();
 sg13g2_decap_4 FILLER_57_150 ();
 sg13g2_fill_1 FILLER_57_154 ();
 sg13g2_decap_4 FILLER_57_160 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_decap_4 FILLER_57_175 ();
 sg13g2_decap_4 FILLER_57_193 ();
 sg13g2_fill_2 FILLER_57_197 ();
 sg13g2_fill_1 FILLER_57_225 ();
 sg13g2_fill_2 FILLER_57_240 ();
 sg13g2_fill_1 FILLER_57_242 ();
 sg13g2_decap_4 FILLER_57_265 ();
 sg13g2_fill_1 FILLER_57_269 ();
 sg13g2_decap_4 FILLER_57_275 ();
 sg13g2_decap_8 FILLER_57_302 ();
 sg13g2_decap_8 FILLER_57_309 ();
 sg13g2_fill_2 FILLER_57_316 ();
 sg13g2_decap_8 FILLER_57_322 ();
 sg13g2_decap_4 FILLER_57_329 ();
 sg13g2_fill_1 FILLER_57_358 ();
 sg13g2_decap_8 FILLER_57_364 ();
 sg13g2_fill_2 FILLER_57_371 ();
 sg13g2_decap_8 FILLER_57_397 ();
 sg13g2_decap_4 FILLER_57_404 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_4 FILLER_58_42 ();
 sg13g2_fill_1 FILLER_58_46 ();
 sg13g2_fill_1 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_99 ();
 sg13g2_fill_2 FILLER_58_106 ();
 sg13g2_fill_2 FILLER_58_118 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_4 FILLER_58_140 ();
 sg13g2_fill_2 FILLER_58_144 ();
 sg13g2_decap_8 FILLER_58_164 ();
 sg13g2_decap_8 FILLER_58_171 ();
 sg13g2_fill_2 FILLER_58_178 ();
 sg13g2_decap_8 FILLER_58_193 ();
 sg13g2_decap_8 FILLER_58_200 ();
 sg13g2_decap_4 FILLER_58_207 ();
 sg13g2_fill_1 FILLER_58_211 ();
 sg13g2_fill_2 FILLER_58_233 ();
 sg13g2_fill_1 FILLER_58_235 ();
 sg13g2_fill_1 FILLER_58_262 ();
 sg13g2_fill_2 FILLER_58_272 ();
 sg13g2_fill_1 FILLER_58_274 ();
 sg13g2_fill_2 FILLER_58_280 ();
 sg13g2_decap_8 FILLER_58_332 ();
 sg13g2_decap_4 FILLER_58_339 ();
 sg13g2_fill_2 FILLER_58_360 ();
 sg13g2_decap_4 FILLER_58_404 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_38 ();
 sg13g2_fill_1 FILLER_59_45 ();
 sg13g2_fill_2 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_100 ();
 sg13g2_fill_2 FILLER_59_107 ();
 sg13g2_fill_1 FILLER_59_109 ();
 sg13g2_fill_1 FILLER_59_141 ();
 sg13g2_fill_1 FILLER_59_157 ();
 sg13g2_decap_4 FILLER_59_162 ();
 sg13g2_fill_2 FILLER_59_166 ();
 sg13g2_decap_4 FILLER_59_211 ();
 sg13g2_fill_1 FILLER_59_215 ();
 sg13g2_decap_8 FILLER_59_220 ();
 sg13g2_decap_4 FILLER_59_227 ();
 sg13g2_fill_2 FILLER_59_236 ();
 sg13g2_decap_8 FILLER_59_262 ();
 sg13g2_fill_2 FILLER_59_311 ();
 sg13g2_fill_1 FILLER_59_313 ();
 sg13g2_fill_2 FILLER_59_340 ();
 sg13g2_fill_1 FILLER_59_342 ();
 sg13g2_decap_8 FILLER_59_347 ();
 sg13g2_fill_2 FILLER_59_354 ();
 sg13g2_fill_2 FILLER_59_361 ();
 sg13g2_fill_2 FILLER_59_375 ();
 sg13g2_fill_2 FILLER_59_391 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_fill_2 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_55 ();
 sg13g2_decap_8 FILLER_60_62 ();
 sg13g2_decap_8 FILLER_60_69 ();
 sg13g2_decap_4 FILLER_60_76 ();
 sg13g2_fill_2 FILLER_60_83 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_4 FILLER_60_98 ();
 sg13g2_fill_1 FILLER_60_128 ();
 sg13g2_fill_2 FILLER_60_136 ();
 sg13g2_fill_1 FILLER_60_138 ();
 sg13g2_decap_8 FILLER_60_173 ();
 sg13g2_decap_8 FILLER_60_180 ();
 sg13g2_decap_8 FILLER_60_191 ();
 sg13g2_decap_8 FILLER_60_198 ();
 sg13g2_decap_8 FILLER_60_205 ();
 sg13g2_decap_4 FILLER_60_212 ();
 sg13g2_fill_1 FILLER_60_216 ();
 sg13g2_decap_4 FILLER_60_220 ();
 sg13g2_fill_2 FILLER_60_224 ();
 sg13g2_fill_2 FILLER_60_230 ();
 sg13g2_decap_4 FILLER_60_236 ();
 sg13g2_decap_4 FILLER_60_245 ();
 sg13g2_fill_1 FILLER_60_249 ();
 sg13g2_fill_2 FILLER_60_286 ();
 sg13g2_fill_1 FILLER_60_288 ();
 sg13g2_fill_1 FILLER_60_311 ();
 sg13g2_fill_2 FILLER_60_322 ();
 sg13g2_fill_1 FILLER_60_324 ();
 sg13g2_decap_8 FILLER_60_329 ();
 sg13g2_decap_8 FILLER_60_336 ();
 sg13g2_decap_8 FILLER_60_343 ();
 sg13g2_decap_8 FILLER_60_350 ();
 sg13g2_fill_2 FILLER_60_357 ();
 sg13g2_fill_1 FILLER_60_375 ();
 sg13g2_decap_8 FILLER_60_402 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_14 ();
 sg13g2_fill_1 FILLER_61_16 ();
 sg13g2_fill_2 FILLER_61_69 ();
 sg13g2_fill_1 FILLER_61_71 ();
 sg13g2_decap_8 FILLER_61_85 ();
 sg13g2_fill_1 FILLER_61_92 ();
 sg13g2_decap_4 FILLER_61_106 ();
 sg13g2_fill_1 FILLER_61_133 ();
 sg13g2_fill_1 FILLER_61_149 ();
 sg13g2_decap_8 FILLER_61_163 ();
 sg13g2_fill_2 FILLER_61_170 ();
 sg13g2_fill_1 FILLER_61_172 ();
 sg13g2_decap_8 FILLER_61_181 ();
 sg13g2_decap_8 FILLER_61_188 ();
 sg13g2_decap_4 FILLER_61_245 ();
 sg13g2_fill_2 FILLER_61_260 ();
 sg13g2_fill_1 FILLER_61_262 ();
 sg13g2_fill_2 FILLER_61_288 ();
 sg13g2_fill_1 FILLER_61_290 ();
 sg13g2_fill_1 FILLER_61_296 ();
 sg13g2_fill_2 FILLER_61_311 ();
 sg13g2_decap_8 FILLER_61_317 ();
 sg13g2_decap_4 FILLER_61_324 ();
 sg13g2_decap_4 FILLER_61_333 ();
 sg13g2_fill_1 FILLER_61_337 ();
 sg13g2_decap_4 FILLER_61_343 ();
 sg13g2_fill_1 FILLER_61_347 ();
 sg13g2_fill_2 FILLER_61_352 ();
 sg13g2_decap_4 FILLER_61_358 ();
 sg13g2_fill_2 FILLER_61_362 ();
 sg13g2_fill_2 FILLER_61_373 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_4 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_103 ();
 sg13g2_decap_8 FILLER_62_110 ();
 sg13g2_fill_2 FILLER_62_127 ();
 sg13g2_fill_1 FILLER_62_134 ();
 sg13g2_decap_4 FILLER_62_174 ();
 sg13g2_fill_2 FILLER_62_178 ();
 sg13g2_fill_2 FILLER_62_190 ();
 sg13g2_fill_1 FILLER_62_192 ();
 sg13g2_decap_4 FILLER_62_260 ();
 sg13g2_fill_2 FILLER_62_264 ();
 sg13g2_decap_8 FILLER_62_271 ();
 sg13g2_decap_8 FILLER_62_278 ();
 sg13g2_decap_4 FILLER_62_285 ();
 sg13g2_fill_2 FILLER_62_289 ();
 sg13g2_fill_2 FILLER_62_305 ();
 sg13g2_fill_1 FILLER_62_316 ();
 sg13g2_fill_1 FILLER_62_382 ();
 sg13g2_decap_4 FILLER_62_405 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_4 FILLER_63_28 ();
 sg13g2_fill_2 FILLER_63_45 ();
 sg13g2_fill_1 FILLER_63_47 ();
 sg13g2_fill_1 FILLER_63_76 ();
 sg13g2_decap_8 FILLER_63_96 ();
 sg13g2_decap_4 FILLER_63_103 ();
 sg13g2_fill_2 FILLER_63_107 ();
 sg13g2_decap_8 FILLER_63_138 ();
 sg13g2_decap_8 FILLER_63_145 ();
 sg13g2_decap_4 FILLER_63_152 ();
 sg13g2_fill_2 FILLER_63_156 ();
 sg13g2_fill_2 FILLER_63_167 ();
 sg13g2_fill_1 FILLER_63_204 ();
 sg13g2_decap_8 FILLER_63_262 ();
 sg13g2_decap_4 FILLER_63_269 ();
 sg13g2_fill_2 FILLER_63_273 ();
 sg13g2_decap_4 FILLER_63_327 ();
 sg13g2_fill_1 FILLER_63_331 ();
 sg13g2_decap_4 FILLER_63_336 ();
 sg13g2_decap_8 FILLER_63_345 ();
 sg13g2_fill_1 FILLER_63_352 ();
 sg13g2_decap_8 FILLER_63_394 ();
 sg13g2_decap_8 FILLER_63_401 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_4 FILLER_64_79 ();
 sg13g2_fill_2 FILLER_64_83 ();
 sg13g2_fill_2 FILLER_64_114 ();
 sg13g2_decap_4 FILLER_64_129 ();
 sg13g2_fill_1 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_155 ();
 sg13g2_decap_8 FILLER_64_162 ();
 sg13g2_fill_1 FILLER_64_177 ();
 sg13g2_fill_2 FILLER_64_188 ();
 sg13g2_decap_4 FILLER_64_226 ();
 sg13g2_fill_2 FILLER_64_230 ();
 sg13g2_decap_8 FILLER_64_236 ();
 sg13g2_decap_8 FILLER_64_243 ();
 sg13g2_decap_8 FILLER_64_250 ();
 sg13g2_fill_2 FILLER_64_257 ();
 sg13g2_fill_1 FILLER_64_259 ();
 sg13g2_fill_1 FILLER_64_335 ();
 sg13g2_decap_8 FILLER_64_392 ();
 sg13g2_decap_8 FILLER_64_399 ();
 sg13g2_fill_2 FILLER_64_406 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_4 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_65 ();
 sg13g2_fill_1 FILLER_65_82 ();
 sg13g2_decap_8 FILLER_65_107 ();
 sg13g2_decap_4 FILLER_65_114 ();
 sg13g2_fill_1 FILLER_65_118 ();
 sg13g2_decap_4 FILLER_65_127 ();
 sg13g2_fill_1 FILLER_65_152 ();
 sg13g2_decap_8 FILLER_65_192 ();
 sg13g2_fill_2 FILLER_65_199 ();
 sg13g2_decap_8 FILLER_65_214 ();
 sg13g2_decap_8 FILLER_65_224 ();
 sg13g2_decap_4 FILLER_65_231 ();
 sg13g2_fill_2 FILLER_65_235 ();
 sg13g2_fill_2 FILLER_65_242 ();
 sg13g2_decap_8 FILLER_65_275 ();
 sg13g2_fill_1 FILLER_65_282 ();
 sg13g2_decap_8 FILLER_65_327 ();
 sg13g2_decap_8 FILLER_65_334 ();
 sg13g2_decap_8 FILLER_65_341 ();
 sg13g2_decap_8 FILLER_65_348 ();
 sg13g2_fill_2 FILLER_65_355 ();
 sg13g2_decap_8 FILLER_65_361 ();
 sg13g2_decap_8 FILLER_65_368 ();
 sg13g2_decap_8 FILLER_65_375 ();
 sg13g2_decap_8 FILLER_65_382 ();
 sg13g2_decap_8 FILLER_65_389 ();
 sg13g2_decap_8 FILLER_65_396 ();
 sg13g2_decap_4 FILLER_65_403 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_fill_1 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_54 ();
 sg13g2_decap_8 FILLER_66_61 ();
 sg13g2_fill_1 FILLER_66_68 ();
 sg13g2_fill_1 FILLER_66_107 ();
 sg13g2_decap_8 FILLER_66_138 ();
 sg13g2_fill_1 FILLER_66_145 ();
 sg13g2_fill_2 FILLER_66_172 ();
 sg13g2_fill_1 FILLER_66_174 ();
 sg13g2_decap_8 FILLER_66_188 ();
 sg13g2_fill_2 FILLER_66_195 ();
 sg13g2_decap_8 FILLER_66_256 ();
 sg13g2_decap_8 FILLER_66_263 ();
 sg13g2_decap_8 FILLER_66_270 ();
 sg13g2_decap_8 FILLER_66_277 ();
 sg13g2_decap_8 FILLER_66_284 ();
 sg13g2_fill_2 FILLER_66_291 ();
 sg13g2_fill_1 FILLER_66_293 ();
 sg13g2_decap_8 FILLER_66_298 ();
 sg13g2_decap_8 FILLER_66_305 ();
 sg13g2_decap_8 FILLER_66_312 ();
 sg13g2_fill_2 FILLER_66_324 ();
 sg13g2_fill_1 FILLER_66_326 ();
 sg13g2_decap_8 FILLER_66_348 ();
 sg13g2_fill_1 FILLER_66_355 ();
 sg13g2_decap_8 FILLER_66_365 ();
 sg13g2_decap_8 FILLER_66_372 ();
 sg13g2_decap_8 FILLER_66_379 ();
 sg13g2_decap_8 FILLER_66_386 ();
 sg13g2_decap_8 FILLER_66_393 ();
 sg13g2_decap_8 FILLER_66_400 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_fill_2 FILLER_67_49 ();
 sg13g2_fill_2 FILLER_67_77 ();
 sg13g2_decap_4 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_fill_2 FILLER_67_119 ();
 sg13g2_fill_1 FILLER_67_121 ();
 sg13g2_decap_8 FILLER_67_141 ();
 sg13g2_fill_1 FILLER_67_161 ();
 sg13g2_fill_2 FILLER_67_165 ();
 sg13g2_fill_1 FILLER_67_167 ();
 sg13g2_decap_8 FILLER_67_177 ();
 sg13g2_decap_8 FILLER_67_184 ();
 sg13g2_decap_8 FILLER_67_191 ();
 sg13g2_decap_8 FILLER_67_198 ();
 sg13g2_fill_1 FILLER_67_205 ();
 sg13g2_fill_2 FILLER_67_219 ();
 sg13g2_fill_1 FILLER_67_221 ();
 sg13g2_fill_2 FILLER_67_254 ();
 sg13g2_decap_8 FILLER_67_264 ();
 sg13g2_decap_8 FILLER_67_302 ();
 sg13g2_fill_2 FILLER_67_309 ();
 sg13g2_fill_1 FILLER_67_311 ();
 sg13g2_decap_8 FILLER_67_378 ();
 sg13g2_decap_8 FILLER_67_385 ();
 sg13g2_decap_8 FILLER_67_392 ();
 sg13g2_decap_8 FILLER_67_399 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_fill_2 FILLER_68_49 ();
 sg13g2_fill_1 FILLER_68_51 ();
 sg13g2_fill_1 FILLER_68_66 ();
 sg13g2_decap_8 FILLER_68_76 ();
 sg13g2_decap_8 FILLER_68_83 ();
 sg13g2_decap_8 FILLER_68_90 ();
 sg13g2_decap_4 FILLER_68_97 ();
 sg13g2_fill_2 FILLER_68_111 ();
 sg13g2_fill_1 FILLER_68_113 ();
 sg13g2_decap_4 FILLER_68_135 ();
 sg13g2_decap_4 FILLER_68_160 ();
 sg13g2_fill_2 FILLER_68_164 ();
 sg13g2_decap_8 FILLER_68_169 ();
 sg13g2_fill_1 FILLER_68_176 ();
 sg13g2_decap_8 FILLER_68_187 ();
 sg13g2_decap_4 FILLER_68_194 ();
 sg13g2_fill_1 FILLER_68_269 ();
 sg13g2_fill_1 FILLER_68_291 ();
 sg13g2_fill_2 FILLER_68_318 ();
 sg13g2_fill_1 FILLER_68_320 ();
 sg13g2_fill_2 FILLER_68_326 ();
 sg13g2_decap_4 FILLER_68_332 ();
 sg13g2_fill_1 FILLER_68_336 ();
 sg13g2_decap_8 FILLER_68_368 ();
 sg13g2_decap_8 FILLER_68_375 ();
 sg13g2_decap_8 FILLER_68_382 ();
 sg13g2_decap_8 FILLER_68_389 ();
 sg13g2_decap_8 FILLER_68_396 ();
 sg13g2_decap_4 FILLER_68_403 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_fill_2 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_61 ();
 sg13g2_decap_8 FILLER_69_68 ();
 sg13g2_fill_2 FILLER_69_78 ();
 sg13g2_fill_1 FILLER_69_80 ();
 sg13g2_decap_8 FILLER_69_193 ();
 sg13g2_decap_8 FILLER_69_200 ();
 sg13g2_fill_2 FILLER_69_207 ();
 sg13g2_decap_8 FILLER_69_213 ();
 sg13g2_decap_8 FILLER_69_220 ();
 sg13g2_fill_2 FILLER_69_227 ();
 sg13g2_decap_8 FILLER_69_232 ();
 sg13g2_fill_2 FILLER_69_239 ();
 sg13g2_fill_1 FILLER_69_241 ();
 sg13g2_fill_1 FILLER_69_245 ();
 sg13g2_fill_2 FILLER_69_255 ();
 sg13g2_fill_1 FILLER_69_261 ();
 sg13g2_fill_1 FILLER_69_272 ();
 sg13g2_decap_8 FILLER_69_277 ();
 sg13g2_fill_1 FILLER_69_284 ();
 sg13g2_decap_8 FILLER_69_362 ();
 sg13g2_decap_8 FILLER_69_369 ();
 sg13g2_decap_8 FILLER_69_376 ();
 sg13g2_decap_8 FILLER_69_383 ();
 sg13g2_decap_8 FILLER_69_390 ();
 sg13g2_decap_8 FILLER_69_397 ();
 sg13g2_decap_4 FILLER_69_404 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_fill_1 FILLER_70_42 ();
 sg13g2_fill_1 FILLER_70_142 ();
 sg13g2_fill_2 FILLER_70_159 ();
 sg13g2_fill_2 FILLER_70_173 ();
 sg13g2_decap_8 FILLER_70_188 ();
 sg13g2_decap_8 FILLER_70_195 ();
 sg13g2_decap_8 FILLER_70_202 ();
 sg13g2_decap_8 FILLER_70_209 ();
 sg13g2_fill_2 FILLER_70_216 ();
 sg13g2_fill_2 FILLER_70_228 ();
 sg13g2_decap_4 FILLER_70_234 ();
 sg13g2_fill_1 FILLER_70_243 ();
 sg13g2_fill_2 FILLER_70_249 ();
 sg13g2_fill_1 FILLER_70_282 ();
 sg13g2_fill_2 FILLER_70_288 ();
 sg13g2_fill_1 FILLER_70_311 ();
 sg13g2_fill_2 FILLER_70_329 ();
 sg13g2_decap_8 FILLER_70_335 ();
 sg13g2_decap_8 FILLER_70_342 ();
 sg13g2_decap_8 FILLER_70_349 ();
 sg13g2_decap_8 FILLER_70_356 ();
 sg13g2_decap_8 FILLER_70_363 ();
 sg13g2_decap_8 FILLER_70_370 ();
 sg13g2_decap_8 FILLER_70_377 ();
 sg13g2_decap_8 FILLER_70_384 ();
 sg13g2_decap_8 FILLER_70_391 ();
 sg13g2_decap_8 FILLER_70_398 ();
 sg13g2_decap_4 FILLER_70_405 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_fill_1 FILLER_71_49 ();
 sg13g2_decap_4 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_fill_2 FILLER_71_84 ();
 sg13g2_fill_1 FILLER_71_86 ();
 sg13g2_fill_2 FILLER_71_97 ();
 sg13g2_fill_1 FILLER_71_99 ();
 sg13g2_fill_1 FILLER_71_118 ();
 sg13g2_decap_8 FILLER_71_122 ();
 sg13g2_decap_4 FILLER_71_132 ();
 sg13g2_fill_1 FILLER_71_145 ();
 sg13g2_decap_8 FILLER_71_186 ();
 sg13g2_decap_4 FILLER_71_193 ();
 sg13g2_fill_1 FILLER_71_197 ();
 sg13g2_fill_1 FILLER_71_238 ();
 sg13g2_fill_1 FILLER_71_244 ();
 sg13g2_fill_1 FILLER_71_256 ();
 sg13g2_decap_8 FILLER_71_278 ();
 sg13g2_decap_4 FILLER_71_285 ();
 sg13g2_decap_4 FILLER_71_295 ();
 sg13g2_decap_8 FILLER_71_317 ();
 sg13g2_decap_8 FILLER_71_324 ();
 sg13g2_decap_8 FILLER_71_331 ();
 sg13g2_decap_8 FILLER_71_338 ();
 sg13g2_decap_8 FILLER_71_345 ();
 sg13g2_decap_8 FILLER_71_352 ();
 sg13g2_decap_8 FILLER_71_359 ();
 sg13g2_decap_8 FILLER_71_366 ();
 sg13g2_decap_8 FILLER_71_373 ();
 sg13g2_decap_8 FILLER_71_380 ();
 sg13g2_decap_8 FILLER_71_387 ();
 sg13g2_decap_8 FILLER_71_394 ();
 sg13g2_decap_8 FILLER_71_401 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_4 FILLER_72_63 ();
 sg13g2_fill_2 FILLER_72_67 ();
 sg13g2_decap_8 FILLER_72_104 ();
 sg13g2_fill_2 FILLER_72_121 ();
 sg13g2_fill_1 FILLER_72_123 ();
 sg13g2_fill_2 FILLER_72_160 ();
 sg13g2_decap_8 FILLER_72_169 ();
 sg13g2_decap_8 FILLER_72_176 ();
 sg13g2_decap_8 FILLER_72_183 ();
 sg13g2_decap_8 FILLER_72_190 ();
 sg13g2_decap_8 FILLER_72_197 ();
 sg13g2_decap_4 FILLER_72_204 ();
 sg13g2_fill_1 FILLER_72_208 ();
 sg13g2_decap_8 FILLER_72_213 ();
 sg13g2_fill_2 FILLER_72_220 ();
 sg13g2_fill_1 FILLER_72_242 ();
 sg13g2_fill_2 FILLER_72_256 ();
 sg13g2_decap_8 FILLER_72_266 ();
 sg13g2_decap_4 FILLER_72_273 ();
 sg13g2_fill_1 FILLER_72_277 ();
 sg13g2_decap_4 FILLER_72_282 ();
 sg13g2_fill_2 FILLER_72_286 ();
 sg13g2_decap_8 FILLER_72_292 ();
 sg13g2_fill_2 FILLER_72_299 ();
 sg13g2_fill_1 FILLER_72_315 ();
 sg13g2_decap_8 FILLER_72_337 ();
 sg13g2_decap_8 FILLER_72_344 ();
 sg13g2_decap_8 FILLER_72_351 ();
 sg13g2_decap_8 FILLER_72_358 ();
 sg13g2_decap_8 FILLER_72_365 ();
 sg13g2_decap_8 FILLER_72_372 ();
 sg13g2_decap_8 FILLER_72_379 ();
 sg13g2_decap_8 FILLER_72_386 ();
 sg13g2_decap_8 FILLER_72_393 ();
 sg13g2_decap_8 FILLER_72_400 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_fill_1 FILLER_73_70 ();
 sg13g2_fill_2 FILLER_73_81 ();
 sg13g2_decap_4 FILLER_73_96 ();
 sg13g2_decap_4 FILLER_73_136 ();
 sg13g2_fill_2 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_177 ();
 sg13g2_decap_8 FILLER_73_184 ();
 sg13g2_decap_8 FILLER_73_191 ();
 sg13g2_fill_2 FILLER_73_198 ();
 sg13g2_fill_1 FILLER_73_200 ();
 sg13g2_decap_4 FILLER_73_260 ();
 sg13g2_fill_2 FILLER_73_264 ();
 sg13g2_fill_2 FILLER_73_269 ();
 sg13g2_fill_1 FILLER_73_271 ();
 sg13g2_fill_2 FILLER_73_278 ();
 sg13g2_fill_1 FILLER_73_294 ();
 sg13g2_fill_1 FILLER_73_310 ();
 sg13g2_decap_8 FILLER_73_337 ();
 sg13g2_decap_8 FILLER_73_344 ();
 sg13g2_decap_8 FILLER_73_351 ();
 sg13g2_decap_8 FILLER_73_358 ();
 sg13g2_decap_8 FILLER_73_365 ();
 sg13g2_decap_8 FILLER_73_372 ();
 sg13g2_decap_8 FILLER_73_379 ();
 sg13g2_decap_8 FILLER_73_386 ();
 sg13g2_decap_8 FILLER_73_393 ();
 sg13g2_decap_8 FILLER_73_400 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_fill_2 FILLER_74_96 ();
 sg13g2_fill_1 FILLER_74_98 ();
 sg13g2_fill_1 FILLER_74_125 ();
 sg13g2_fill_1 FILLER_74_135 ();
 sg13g2_decap_8 FILLER_74_159 ();
 sg13g2_decap_8 FILLER_74_166 ();
 sg13g2_decap_8 FILLER_74_173 ();
 sg13g2_decap_8 FILLER_74_180 ();
 sg13g2_decap_8 FILLER_74_187 ();
 sg13g2_decap_8 FILLER_74_194 ();
 sg13g2_decap_8 FILLER_74_201 ();
 sg13g2_fill_2 FILLER_74_208 ();
 sg13g2_fill_1 FILLER_74_265 ();
 sg13g2_fill_2 FILLER_74_300 ();
 sg13g2_fill_1 FILLER_74_302 ();
 sg13g2_decap_8 FILLER_74_329 ();
 sg13g2_decap_8 FILLER_74_336 ();
 sg13g2_decap_8 FILLER_74_343 ();
 sg13g2_decap_8 FILLER_74_350 ();
 sg13g2_decap_8 FILLER_74_357 ();
 sg13g2_decap_8 FILLER_74_364 ();
 sg13g2_decap_8 FILLER_74_371 ();
 sg13g2_decap_8 FILLER_74_378 ();
 sg13g2_decap_8 FILLER_74_385 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_fill_2 FILLER_75_77 ();
 sg13g2_fill_1 FILLER_75_79 ();
 sg13g2_fill_1 FILLER_75_85 ();
 sg13g2_decap_8 FILLER_75_95 ();
 sg13g2_decap_8 FILLER_75_102 ();
 sg13g2_fill_1 FILLER_75_109 ();
 sg13g2_fill_1 FILLER_75_114 ();
 sg13g2_fill_1 FILLER_75_124 ();
 sg13g2_decap_8 FILLER_75_136 ();
 sg13g2_decap_4 FILLER_75_143 ();
 sg13g2_decap_8 FILLER_75_150 ();
 sg13g2_decap_8 FILLER_75_157 ();
 sg13g2_decap_8 FILLER_75_164 ();
 sg13g2_decap_8 FILLER_75_171 ();
 sg13g2_decap_8 FILLER_75_178 ();
 sg13g2_decap_8 FILLER_75_185 ();
 sg13g2_decap_8 FILLER_75_192 ();
 sg13g2_decap_8 FILLER_75_199 ();
 sg13g2_decap_4 FILLER_75_206 ();
 sg13g2_fill_2 FILLER_75_210 ();
 sg13g2_fill_2 FILLER_75_216 ();
 sg13g2_decap_8 FILLER_75_239 ();
 sg13g2_decap_4 FILLER_75_246 ();
 sg13g2_fill_1 FILLER_75_250 ();
 sg13g2_fill_2 FILLER_75_287 ();
 sg13g2_fill_1 FILLER_75_289 ();
 sg13g2_decap_8 FILLER_75_328 ();
 sg13g2_decap_8 FILLER_75_335 ();
 sg13g2_decap_8 FILLER_75_342 ();
 sg13g2_decap_8 FILLER_75_349 ();
 sg13g2_decap_8 FILLER_75_356 ();
 sg13g2_decap_8 FILLER_75_363 ();
 sg13g2_decap_8 FILLER_75_370 ();
 sg13g2_decap_8 FILLER_75_377 ();
 sg13g2_decap_8 FILLER_75_384 ();
 sg13g2_decap_8 FILLER_75_391 ();
 sg13g2_decap_8 FILLER_75_398 ();
 sg13g2_decap_4 FILLER_75_405 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_fill_1 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_89 ();
 sg13g2_decap_8 FILLER_76_96 ();
 sg13g2_decap_8 FILLER_76_103 ();
 sg13g2_decap_8 FILLER_76_110 ();
 sg13g2_decap_8 FILLER_76_117 ();
 sg13g2_decap_8 FILLER_76_124 ();
 sg13g2_decap_8 FILLER_76_131 ();
 sg13g2_decap_8 FILLER_76_138 ();
 sg13g2_decap_8 FILLER_76_145 ();
 sg13g2_decap_8 FILLER_76_152 ();
 sg13g2_decap_8 FILLER_76_159 ();
 sg13g2_decap_8 FILLER_76_166 ();
 sg13g2_decap_8 FILLER_76_173 ();
 sg13g2_decap_8 FILLER_76_180 ();
 sg13g2_decap_8 FILLER_76_187 ();
 sg13g2_decap_8 FILLER_76_194 ();
 sg13g2_decap_8 FILLER_76_201 ();
 sg13g2_decap_8 FILLER_76_208 ();
 sg13g2_decap_8 FILLER_76_215 ();
 sg13g2_decap_8 FILLER_76_222 ();
 sg13g2_decap_8 FILLER_76_229 ();
 sg13g2_fill_1 FILLER_76_244 ();
 sg13g2_fill_1 FILLER_76_262 ();
 sg13g2_fill_2 FILLER_76_279 ();
 sg13g2_decap_4 FILLER_76_288 ();
 sg13g2_fill_2 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_323 ();
 sg13g2_decap_8 FILLER_76_330 ();
 sg13g2_decap_8 FILLER_76_337 ();
 sg13g2_decap_8 FILLER_76_344 ();
 sg13g2_decap_8 FILLER_76_351 ();
 sg13g2_decap_8 FILLER_76_358 ();
 sg13g2_decap_8 FILLER_76_365 ();
 sg13g2_decap_8 FILLER_76_372 ();
 sg13g2_decap_8 FILLER_76_379 ();
 sg13g2_decap_8 FILLER_76_386 ();
 sg13g2_decap_8 FILLER_76_393 ();
 sg13g2_decap_8 FILLER_76_400 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_4 FILLER_77_217 ();
 sg13g2_fill_1 FILLER_77_221 ();
 sg13g2_fill_1 FILLER_77_283 ();
 sg13g2_decap_8 FILLER_77_328 ();
 sg13g2_decap_8 FILLER_77_335 ();
 sg13g2_decap_8 FILLER_77_342 ();
 sg13g2_decap_8 FILLER_77_349 ();
 sg13g2_decap_8 FILLER_77_356 ();
 sg13g2_decap_8 FILLER_77_363 ();
 sg13g2_decap_8 FILLER_77_370 ();
 sg13g2_decap_8 FILLER_77_377 ();
 sg13g2_decap_8 FILLER_77_384 ();
 sg13g2_decap_8 FILLER_77_391 ();
 sg13g2_decap_8 FILLER_77_398 ();
 sg13g2_decap_4 FILLER_77_405 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_fill_2 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_240 ();
 sg13g2_decap_8 FILLER_78_247 ();
 sg13g2_decap_8 FILLER_78_258 ();
 sg13g2_decap_4 FILLER_78_265 ();
 sg13g2_fill_2 FILLER_78_269 ();
 sg13g2_decap_8 FILLER_78_323 ();
 sg13g2_decap_8 FILLER_78_330 ();
 sg13g2_decap_8 FILLER_78_337 ();
 sg13g2_decap_8 FILLER_78_344 ();
 sg13g2_decap_8 FILLER_78_351 ();
 sg13g2_decap_8 FILLER_78_358 ();
 sg13g2_decap_8 FILLER_78_365 ();
 sg13g2_decap_8 FILLER_78_372 ();
 sg13g2_decap_8 FILLER_78_379 ();
 sg13g2_decap_8 FILLER_78_386 ();
 sg13g2_decap_8 FILLER_78_393 ();
 sg13g2_decap_8 FILLER_78_400 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_4 FILLER_79_238 ();
 sg13g2_fill_2 FILLER_79_268 ();
 sg13g2_fill_2 FILLER_79_296 ();
 sg13g2_fill_1 FILLER_79_298 ();
 sg13g2_decap_8 FILLER_79_303 ();
 sg13g2_decap_8 FILLER_79_310 ();
 sg13g2_decap_8 FILLER_79_317 ();
 sg13g2_decap_8 FILLER_79_324 ();
 sg13g2_decap_8 FILLER_79_331 ();
 sg13g2_decap_8 FILLER_79_338 ();
 sg13g2_decap_8 FILLER_79_345 ();
 sg13g2_decap_8 FILLER_79_352 ();
 sg13g2_decap_8 FILLER_79_359 ();
 sg13g2_decap_8 FILLER_79_366 ();
 sg13g2_decap_8 FILLER_79_373 ();
 sg13g2_decap_8 FILLER_79_380 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_8 FILLER_80_123 ();
 sg13g2_decap_8 FILLER_80_130 ();
 sg13g2_decap_8 FILLER_80_137 ();
 sg13g2_decap_8 FILLER_80_144 ();
 sg13g2_decap_8 FILLER_80_151 ();
 sg13g2_decap_8 FILLER_80_158 ();
 sg13g2_decap_8 FILLER_80_165 ();
 sg13g2_decap_8 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_179 ();
 sg13g2_decap_8 FILLER_80_186 ();
 sg13g2_decap_8 FILLER_80_193 ();
 sg13g2_decap_8 FILLER_80_200 ();
 sg13g2_decap_8 FILLER_80_207 ();
 sg13g2_decap_8 FILLER_80_214 ();
 sg13g2_decap_8 FILLER_80_221 ();
 sg13g2_decap_8 FILLER_80_228 ();
 sg13g2_decap_8 FILLER_80_235 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_decap_4 FILLER_80_249 ();
 sg13g2_decap_8 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_fill_2 FILLER_80_278 ();
 sg13g2_fill_1 FILLER_80_280 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_4 FILLER_80_306 ();
 sg13g2_fill_2 FILLER_80_310 ();
 sg13g2_fill_2 FILLER_80_317 ();
 sg13g2_fill_1 FILLER_80_319 ();
 sg13g2_fill_2 FILLER_80_325 ();
 sg13g2_fill_1 FILLER_80_327 ();
 sg13g2_fill_2 FILLER_80_333 ();
 sg13g2_fill_1 FILLER_80_335 ();
 sg13g2_fill_2 FILLER_80_341 ();
 sg13g2_fill_1 FILLER_80_343 ();
 sg13g2_decap_8 FILLER_80_376 ();
 sg13g2_decap_8 FILLER_80_383 ();
 sg13g2_decap_8 FILLER_80_390 ();
 sg13g2_decap_8 FILLER_80_397 ();
 sg13g2_decap_4 FILLER_80_404 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net198;
 assign uio_oe[1] = net199;
 assign uio_oe[2] = net200;
 assign uio_oe[3] = net201;
 assign uio_oe[4] = net202;
 assign uio_oe[5] = net203;
 assign uio_oe[6] = net204;
 assign uio_oe[7] = net205;
endmodule
