module tt_um_Xelef2000 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire clknet_0_clk;
 wire \byte_counter_r[0] ;
 wire \byte_counter_r[1] ;
 wire fsm_state_next;
 wire fsm_state_r;
 wire \i_random.bit_count[0] ;
 wire \i_random.bit_count[1] ;
 wire \i_random.bit_count[2] ;
 wire \i_random.bit_count[3] ;
 wire \i_random.bit_count[4] ;
 wire \i_random.combined_ring_bit ;
 wire \i_random.debiased_bit ;
 wire \i_random.debiased_bit_valid ;
 wire \i_random.first_bit ;
 wire \i_random.ready ;
 wire \i_random.ring_bit_12 ;
 wire \i_random.ring_bit_24 ;
 wire \i_random.ring_bit_6 ;
 wire \i_random.rnd_out[0] ;
 wire \i_random.rnd_out[10] ;
 wire \i_random.rnd_out[11] ;
 wire \i_random.rnd_out[12] ;
 wire \i_random.rnd_out[13] ;
 wire \i_random.rnd_out[14] ;
 wire \i_random.rnd_out[15] ;
 wire \i_random.rnd_out[16] ;
 wire \i_random.rnd_out[17] ;
 wire \i_random.rnd_out[18] ;
 wire \i_random.rnd_out[19] ;
 wire \i_random.rnd_out[1] ;
 wire \i_random.rnd_out[20] ;
 wire \i_random.rnd_out[21] ;
 wire \i_random.rnd_out[22] ;
 wire \i_random.rnd_out[23] ;
 wire \i_random.rnd_out[24] ;
 wire \i_random.rnd_out[25] ;
 wire \i_random.rnd_out[26] ;
 wire \i_random.rnd_out[27] ;
 wire \i_random.rnd_out[28] ;
 wire \i_random.rnd_out[29] ;
 wire \i_random.rnd_out[2] ;
 wire \i_random.rnd_out[30] ;
 wire \i_random.rnd_out[31] ;
 wire \i_random.rnd_out[3] ;
 wire \i_random.rnd_out[4] ;
 wire \i_random.rnd_out[5] ;
 wire \i_random.rnd_out[6] ;
 wire \i_random.rnd_out[7] ;
 wire \i_random.rnd_out[8] ;
 wire \i_random.rnd_out[9] ;
 wire \i_random.rnd_sync ;
 wire \i_random.state ;
 wire \i_random.sync1 ;
 wire \i_random.u_ring12.gated ;
 wire \i_random.u_ring12.n1 ;
 wire \i_random.u_ring12.n10 ;
 wire \i_random.u_ring12.n2 ;
 wire \i_random.u_ring12.n3 ;
 wire \i_random.u_ring12.n4 ;
 wire \i_random.u_ring12.n5 ;
 wire \i_random.u_ring12.n6 ;
 wire \i_random.u_ring12.n7 ;
 wire \i_random.u_ring12.n8 ;
 wire \i_random.u_ring12.n9 ;
 wire \i_random.u_ring24.gated ;
 wire \i_random.u_ring24.n1 ;
 wire \i_random.u_ring24.n10 ;
 wire \i_random.u_ring24.n11 ;
 wire \i_random.u_ring24.n12 ;
 wire \i_random.u_ring24.n13 ;
 wire \i_random.u_ring24.n14 ;
 wire \i_random.u_ring24.n15 ;
 wire \i_random.u_ring24.n16 ;
 wire \i_random.u_ring24.n17 ;
 wire \i_random.u_ring24.n18 ;
 wire \i_random.u_ring24.n19 ;
 wire \i_random.u_ring24.n2 ;
 wire \i_random.u_ring24.n20 ;
 wire \i_random.u_ring24.n21 ;
 wire \i_random.u_ring24.n22 ;
 wire \i_random.u_ring24.n3 ;
 wire \i_random.u_ring24.n4 ;
 wire \i_random.u_ring24.n5 ;
 wire \i_random.u_ring24.n6 ;
 wire \i_random.u_ring24.n7 ;
 wire \i_random.u_ring24.n8 ;
 wire \i_random.u_ring24.n9 ;
 wire \i_random.u_ring6.gated ;
 wire \i_random.u_ring6.n1 ;
 wire \i_random.u_ring6.n2 ;
 wire \i_random.u_ring6.n3 ;
 wire \i_random.u_ring6.n4 ;
 wire \i_uart_tx.bit_counter[0] ;
 wire \i_uart_tx.bit_counter[1] ;
 wire \i_uart_tx.bit_counter[2] ;
 wire \i_uart_tx.bit_counter[3] ;
 wire \i_uart_tx.cycle_counter[0] ;
 wire \i_uart_tx.cycle_counter[1] ;
 wire \i_uart_tx.cycle_counter[2] ;
 wire \i_uart_tx.cycle_counter[3] ;
 wire \i_uart_tx.cycle_counter[4] ;
 wire \i_uart_tx.cycle_counter[5] ;
 wire \i_uart_tx.cycle_counter[6] ;
 wire \i_uart_tx.data_to_send[0] ;
 wire \i_uart_tx.data_to_send[1] ;
 wire \i_uart_tx.data_to_send[2] ;
 wire \i_uart_tx.data_to_send[3] ;
 wire \i_uart_tx.data_to_send[4] ;
 wire \i_uart_tx.data_to_send[5] ;
 wire \i_uart_tx.data_to_send[6] ;
 wire \i_uart_tx.data_to_send[7] ;
 wire \i_uart_tx.fsm_state[0] ;
 wire \i_uart_tx.fsm_state[1] ;
 wire \i_uart_tx.txd_reg ;
 wire \i_uart_tx.uart_tx_data[0] ;
 wire \i_uart_tx.uart_tx_data[1] ;
 wire \i_uart_tx.uart_tx_data[2] ;
 wire \i_uart_tx.uart_tx_data[3] ;
 wire \i_uart_tx.uart_tx_data[4] ;
 wire \i_uart_tx.uart_tx_data[5] ;
 wire \i_uart_tx.uart_tx_data[6] ;
 wire \i_uart_tx.uart_tx_data[7] ;
 wire \i_uart_tx.uart_tx_en ;
 wire \random_buffer_r[0] ;
 wire \random_buffer_r[10] ;
 wire \random_buffer_r[11] ;
 wire \random_buffer_r[12] ;
 wire \random_buffer_r[13] ;
 wire \random_buffer_r[14] ;
 wire \random_buffer_r[15] ;
 wire \random_buffer_r[16] ;
 wire \random_buffer_r[17] ;
 wire \random_buffer_r[18] ;
 wire \random_buffer_r[19] ;
 wire \random_buffer_r[1] ;
 wire \random_buffer_r[20] ;
 wire \random_buffer_r[21] ;
 wire \random_buffer_r[22] ;
 wire \random_buffer_r[23] ;
 wire \random_buffer_r[24] ;
 wire \random_buffer_r[25] ;
 wire \random_buffer_r[26] ;
 wire \random_buffer_r[27] ;
 wire \random_buffer_r[28] ;
 wire \random_buffer_r[29] ;
 wire \random_buffer_r[2] ;
 wire \random_buffer_r[30] ;
 wire \random_buffer_r[31] ;
 wire \random_buffer_r[3] ;
 wire \random_buffer_r[4] ;
 wire \random_buffer_r[5] ;
 wire \random_buffer_r[6] ;
 wire \random_buffer_r[7] ;
 wire \random_buffer_r[8] ;
 wire \random_buffer_r[9] ;
 wire uart_tx_en_next;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net1;
 wire net2;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;

 sg13g2_inv_1 _377_ (.Y(_110_),
    .A(\i_uart_tx.bit_counter[3] ));
 sg13g2_inv_1 _378_ (.Y(_111_),
    .A(net84));
 sg13g2_inv_1 _379_ (.Y(_112_),
    .A(\i_uart_tx.fsm_state[0] ));
 sg13g2_inv_2 _380_ (.Y(_113_),
    .A(net142));
 sg13g2_inv_1 _381_ (.Y(_114_),
    .A(net153));
 sg13g2_inv_1 _382_ (.Y(_115_),
    .A(net67));
 sg13g2_inv_1 _383_ (.Y(_116_),
    .A(\random_buffer_r[0] ));
 sg13g2_inv_1 _384_ (.Y(_117_),
    .A(\random_buffer_r[1] ));
 sg13g2_inv_1 _385_ (.Y(_118_),
    .A(\random_buffer_r[3] ));
 sg13g2_inv_1 _386_ (.Y(_119_),
    .A(\random_buffer_r[5] ));
 sg13g2_inv_1 _387_ (.Y(_120_),
    .A(\random_buffer_r[6] ));
 sg13g2_inv_1 _388_ (.Y(_121_),
    .A(net51));
 sg13g2_inv_1 _389_ (.Y(_122_),
    .A(net234));
 sg13g2_inv_1 _390_ (.Y(_123_),
    .A(net208));
 sg13g2_inv_1 _391_ (.Y(_124_),
    .A(net75));
 sg13g2_nor2_2 _392_ (.A(net127),
    .B(\i_uart_tx.fsm_state[0] ),
    .Y(_125_));
 sg13g2_or2_1 _393_ (.X(_126_),
    .B(\i_uart_tx.fsm_state[0] ),
    .A(net127));
 sg13g2_nand2b_2 _394_ (.Y(_127_),
    .B(_125_),
    .A_N(net210));
 sg13g2_inv_2 _395_ (.Y(uart_tx_en_next),
    .A(_127_));
 sg13g2_nor2b_1 _396_ (.A(fsm_state_r),
    .B_N(\i_random.ready ),
    .Y(_128_));
 sg13g2_and2_1 _397_ (.A(\byte_counter_r[0] ),
    .B(\byte_counter_r[1] ),
    .X(_129_));
 sg13g2_nand2_1 _398_ (.Y(_130_),
    .A(_125_),
    .B(_129_));
 sg13g2_nand2_1 _399_ (.Y(_131_),
    .A(fsm_state_r),
    .B(_125_));
 sg13g2_a21o_1 _400_ (.A2(_130_),
    .A1(net250),
    .B1(net126),
    .X(fsm_state_next));
 sg13g2_xnor2_1 _401_ (.Y(_132_),
    .A(\i_random.ring_bit_6 ),
    .B(\i_random.ring_bit_24 ));
 sg13g2_xnor2_1 _402_ (.Y(\i_random.combined_ring_bit ),
    .A(\i_random.ring_bit_12 ),
    .B(_132_));
 sg13g2_nor3_1 _403_ (.A(\i_uart_tx.bit_counter[3] ),
    .B(\i_uart_tx.bit_counter[2] ),
    .C(\i_uart_tx.bit_counter[1] ),
    .Y(_133_));
 sg13g2_nand2_1 _404_ (.Y(_134_),
    .A(\i_uart_tx.bit_counter[0] ),
    .B(_133_));
 sg13g2_and2_1 _405_ (.A(\i_uart_tx.cycle_counter[5] ),
    .B(\i_uart_tx.cycle_counter[4] ),
    .X(_135_));
 sg13g2_nor3_2 _406_ (.A(\i_uart_tx.cycle_counter[6] ),
    .B(\i_uart_tx.cycle_counter[3] ),
    .C(\i_uart_tx.cycle_counter[1] ),
    .Y(_136_));
 sg13g2_nor2b_2 _407_ (.A(\i_uart_tx.cycle_counter[0] ),
    .B_N(\i_uart_tx.cycle_counter[2] ),
    .Y(_137_));
 sg13g2_and3_1 _408_ (.X(_138_),
    .A(_135_),
    .B(_136_),
    .C(_137_));
 sg13g2_nand3_1 _409_ (.B(_136_),
    .C(_137_),
    .A(_135_),
    .Y(_139_));
 sg13g2_and2_2 _410_ (.A(net241),
    .B(_125_),
    .X(_140_));
 sg13g2_nand2_1 _411_ (.Y(_141_),
    .A(net241),
    .B(_125_));
 sg13g2_nor4_1 _412_ (.A(_110_),
    .B(\i_uart_tx.bit_counter[2] ),
    .C(\i_uart_tx.bit_counter[1] ),
    .D(\i_uart_tx.bit_counter[0] ),
    .Y(_142_));
 sg13g2_a21o_1 _413_ (.A2(_134_),
    .A1(\i_uart_tx.fsm_state[0] ),
    .B1(_142_),
    .X(_143_));
 sg13g2_nor2_1 _414_ (.A(net127),
    .B(_112_),
    .Y(_144_));
 sg13g2_a221oi_1 _415_ (.B2(_139_),
    .C1(_140_),
    .B1(_144_),
    .A1(net127),
    .Y(_145_),
    .A2(_143_));
 sg13g2_nor2_1 _416_ (.A(_113_),
    .B(_145_),
    .Y(_004_));
 sg13g2_nor2b_1 _417_ (.A(\i_uart_tx.fsm_state[0] ),
    .B_N(net127),
    .Y(_146_));
 sg13g2_a221oi_1 _418_ (.B2(_144_),
    .C1(_146_),
    .B1(_138_),
    .A1(net256),
    .Y(_147_),
    .A2(_134_));
 sg13g2_nor2_1 _419_ (.A(_113_),
    .B(net257),
    .Y(_005_));
 sg13g2_nand4_1 _420_ (.B(_135_),
    .C(_136_),
    .A(\i_uart_tx.fsm_state[1] ),
    .Y(_148_),
    .D(_137_));
 sg13g2_nor2_2 _421_ (.A(net204),
    .B(_148_),
    .Y(_149_));
 sg13g2_nand4_1 _422_ (.B(_136_),
    .C(_137_),
    .A(_135_),
    .Y(_150_),
    .D(_146_));
 sg13g2_nand2_2 _423_ (.Y(_151_),
    .A(_141_),
    .B(_150_));
 sg13g2_nor2_1 _424_ (.A(net186),
    .B(_151_),
    .Y(_152_));
 sg13g2_o21ai_1 _425_ (.B1(net143),
    .Y(_153_),
    .A1(net171),
    .A2(net111));
 sg13g2_nor2_1 _426_ (.A(net181),
    .B(_150_),
    .Y(_154_));
 sg13g2_nor3_1 _427_ (.A(_152_),
    .B(_153_),
    .C(_154_),
    .Y(_006_));
 sg13g2_nor2_1 _428_ (.A(net181),
    .B(_151_),
    .Y(_155_));
 sg13g2_o21ai_1 _429_ (.B1(net143),
    .Y(_156_),
    .A1(net155),
    .A2(net111));
 sg13g2_nor2_1 _430_ (.A(\i_uart_tx.data_to_send[2] ),
    .B(_150_),
    .Y(_157_));
 sg13g2_nor3_1 _431_ (.A(net182),
    .B(_156_),
    .C(_157_),
    .Y(_007_));
 sg13g2_nor2_1 _432_ (.A(\i_uart_tx.data_to_send[2] ),
    .B(_151_),
    .Y(_158_));
 sg13g2_o21ai_1 _433_ (.B1(net140),
    .Y(_159_),
    .A1(\i_uart_tx.uart_tx_data[2] ),
    .A2(net111));
 sg13g2_nor2_1 _434_ (.A(net105),
    .B(_150_),
    .Y(_160_));
 sg13g2_nor3_1 _435_ (.A(_158_),
    .B(_159_),
    .C(_160_),
    .Y(_008_));
 sg13g2_nand2b_1 _436_ (.Y(_161_),
    .B(_140_),
    .A_N(net73));
 sg13g2_o21ai_1 _437_ (.B1(_161_),
    .Y(_162_),
    .A1(net239),
    .A2(_140_));
 sg13g2_o21ai_1 _438_ (.B1(net142),
    .Y(_163_),
    .A1(net105),
    .A2(_151_));
 sg13g2_a21oi_1 _439_ (.A1(_151_),
    .A2(_162_),
    .Y(_009_),
    .B1(_163_));
 sg13g2_nor2_1 _440_ (.A(_122_),
    .B(net111),
    .Y(_164_));
 sg13g2_a21oi_1 _441_ (.A1(net80),
    .A2(net111),
    .Y(_165_),
    .B1(_164_));
 sg13g2_o21ai_1 _442_ (.B1(net140),
    .Y(_166_),
    .A1(net239),
    .A2(_151_));
 sg13g2_a21oi_1 _443_ (.A1(_151_),
    .A2(_165_),
    .Y(_010_),
    .B1(_166_));
 sg13g2_nand3_1 _444_ (.B(net111),
    .C(_150_),
    .A(net80),
    .Y(_167_));
 sg13g2_and2_1 _445_ (.A(net235),
    .B(net111),
    .X(_168_));
 sg13g2_a22oi_1 _446_ (.Y(_169_),
    .B1(_149_),
    .B2(_168_),
    .A2(_140_),
    .A1(net78));
 sg13g2_a21oi_1 _447_ (.A1(_167_),
    .A2(_169_),
    .Y(_011_),
    .B1(_113_));
 sg13g2_nand2_1 _448_ (.Y(_170_),
    .A(_150_),
    .B(_168_));
 sg13g2_and2_1 _449_ (.A(\i_uart_tx.data_to_send[7] ),
    .B(net111),
    .X(_171_));
 sg13g2_a22oi_1 _450_ (.Y(_172_),
    .B1(_149_),
    .B2(_171_),
    .A2(_140_),
    .A1(net57));
 sg13g2_a21oi_1 _451_ (.A1(_170_),
    .A2(_172_),
    .Y(_012_),
    .B1(_113_));
 sg13g2_nor2_1 _452_ (.A(\byte_counter_r[0] ),
    .B(\byte_counter_r[1] ),
    .Y(_173_));
 sg13g2_nor2b_2 _453_ (.A(\byte_counter_r[1] ),
    .B_N(\byte_counter_r[0] ),
    .Y(_174_));
 sg13g2_nor2b_2 _454_ (.A(\byte_counter_r[0] ),
    .B_N(\byte_counter_r[1] ),
    .Y(_175_));
 sg13g2_a22oi_1 _455_ (.Y(_176_),
    .B1(_175_),
    .B2(net103),
    .A2(_174_),
    .A1(\random_buffer_r[8] ));
 sg13g2_a21oi_1 _456_ (.A1(net96),
    .A2(net120),
    .Y(_177_),
    .B1(net118));
 sg13g2_a22oi_1 _457_ (.Y(_178_),
    .B1(_176_),
    .B2(_177_),
    .A2(net119),
    .A1(_116_));
 sg13g2_mux2_1 _458_ (.A0(net171),
    .A1(_178_),
    .S(uart_tx_en_next),
    .X(_013_));
 sg13g2_a22oi_1 _459_ (.Y(_179_),
    .B1(_175_),
    .B2(net94),
    .A2(_174_),
    .A1(\random_buffer_r[9] ));
 sg13g2_a21oi_1 _460_ (.A1(\random_buffer_r[25] ),
    .A2(net120),
    .Y(_180_),
    .B1(net118));
 sg13g2_a22oi_1 _461_ (.Y(_181_),
    .B1(_179_),
    .B2(_180_),
    .A2(net119),
    .A1(_117_));
 sg13g2_mux2_1 _462_ (.A0(net155),
    .A1(_181_),
    .S(uart_tx_en_next),
    .X(_014_));
 sg13g2_and2_1 _463_ (.A(net163),
    .B(_175_),
    .X(_182_));
 sg13g2_a221oi_1 _464_ (.B2(net151),
    .C1(_182_),
    .B1(_174_),
    .A1(net192),
    .Y(_183_),
    .A2(net120));
 sg13g2_a21oi_1 _465_ (.A1(net159),
    .A2(net119),
    .Y(_184_),
    .B1(_127_));
 sg13g2_a22oi_1 _466_ (.Y(_015_),
    .B1(_183_),
    .B2(_184_),
    .A2(_127_),
    .A1(_123_));
 sg13g2_a22oi_1 _467_ (.Y(_185_),
    .B1(_175_),
    .B2(\random_buffer_r[19] ),
    .A2(_174_),
    .A1(\random_buffer_r[11] ));
 sg13g2_a21oi_1 _468_ (.A1(\random_buffer_r[27] ),
    .A2(net120),
    .Y(_186_),
    .B1(net118));
 sg13g2_a22oi_1 _469_ (.Y(_187_),
    .B1(_185_),
    .B2(_186_),
    .A2(net118),
    .A1(_118_));
 sg13g2_mux2_1 _470_ (.A0(net73),
    .A1(_187_),
    .S(uart_tx_en_next),
    .X(_016_));
 sg13g2_and2_1 _471_ (.A(net167),
    .B(_175_),
    .X(_188_));
 sg13g2_a221oi_1 _472_ (.B2(net90),
    .C1(_188_),
    .B1(_174_),
    .A1(net109),
    .Y(_189_),
    .A2(net120));
 sg13g2_a21oi_1 _473_ (.A1(net146),
    .A2(net119),
    .Y(_190_),
    .B1(_127_));
 sg13g2_a22oi_1 _474_ (.Y(_017_),
    .B1(_189_),
    .B2(_190_),
    .A2(_127_),
    .A1(_122_));
 sg13g2_a22oi_1 _475_ (.Y(_191_),
    .B1(_175_),
    .B2(\random_buffer_r[21] ),
    .A2(_174_),
    .A1(\random_buffer_r[13] ));
 sg13g2_a21oi_1 _476_ (.A1(\random_buffer_r[29] ),
    .A2(net120),
    .Y(_192_),
    .B1(net118));
 sg13g2_a22oi_1 _477_ (.Y(_193_),
    .B1(_191_),
    .B2(_192_),
    .A2(net118),
    .A1(_119_));
 sg13g2_mux2_1 _478_ (.A0(net78),
    .A1(_193_),
    .S(uart_tx_en_next),
    .X(_018_));
 sg13g2_a22oi_1 _479_ (.Y(_194_),
    .B1(_175_),
    .B2(\random_buffer_r[22] ),
    .A2(_174_),
    .A1(\random_buffer_r[14] ));
 sg13g2_a21oi_1 _480_ (.A1(\random_buffer_r[30] ),
    .A2(net120),
    .Y(_195_),
    .B1(net118));
 sg13g2_a22oi_1 _481_ (.Y(_196_),
    .B1(_194_),
    .B2(_195_),
    .A2(net118),
    .A1(_120_));
 sg13g2_mux2_1 _482_ (.A0(net57),
    .A1(_196_),
    .S(uart_tx_en_next),
    .X(_019_));
 sg13g2_and2_1 _483_ (.A(net157),
    .B(_175_),
    .X(_197_));
 sg13g2_a221oi_1 _484_ (.B2(net175),
    .C1(_197_),
    .B1(_174_),
    .A1(net161),
    .Y(_198_),
    .A2(net120));
 sg13g2_a21oi_1 _485_ (.A1(net179),
    .A2(net119),
    .Y(_199_),
    .B1(_127_));
 sg13g2_a22oi_1 _486_ (.Y(_020_),
    .B1(_198_),
    .B2(_199_),
    .A2(_127_),
    .A1(_111_));
 sg13g2_nand2_1 _487_ (.Y(_200_),
    .A(net53),
    .B(net126));
 sg13g2_o21ai_1 _488_ (.B1(_200_),
    .Y(_021_),
    .A1(_116_),
    .A2(net126));
 sg13g2_nand2_1 _489_ (.Y(_201_),
    .A(net62),
    .B(_128_));
 sg13g2_o21ai_1 _490_ (.B1(net63),
    .Y(_022_),
    .A1(_117_),
    .A2(net126));
 sg13g2_mux2_1 _491_ (.A0(net159),
    .A1(\i_random.rnd_out[2] ),
    .S(net126),
    .X(_023_));
 sg13g2_nand2_1 _492_ (.Y(_202_),
    .A(net55),
    .B(net124));
 sg13g2_o21ai_1 _493_ (.B1(_202_),
    .Y(_024_),
    .A1(_118_),
    .A2(net123));
 sg13g2_mux2_1 _494_ (.A0(net146),
    .A1(\i_random.rnd_out[4] ),
    .S(net124),
    .X(_025_));
 sg13g2_nand2_1 _495_ (.Y(_203_),
    .A(net92),
    .B(net124));
 sg13g2_o21ai_1 _496_ (.B1(_203_),
    .Y(_026_),
    .A1(_119_),
    .A2(net123));
 sg13g2_nand2_1 _497_ (.Y(_204_),
    .A(net69),
    .B(net123));
 sg13g2_o21ai_1 _498_ (.B1(_204_),
    .Y(_027_),
    .A1(_120_),
    .A2(net123));
 sg13g2_mux2_1 _499_ (.A0(net179),
    .A1(\i_random.rnd_out[7] ),
    .S(net123),
    .X(_028_));
 sg13g2_mux2_1 _500_ (.A0(net86),
    .A1(\i_random.rnd_out[8] ),
    .S(net123),
    .X(_029_));
 sg13g2_mux2_1 _501_ (.A0(net65),
    .A1(\i_random.rnd_out[9] ),
    .S(net123),
    .X(_030_));
 sg13g2_mux2_1 _502_ (.A0(net151),
    .A1(\i_random.rnd_out[10] ),
    .S(net123),
    .X(_031_));
 sg13g2_mux2_1 _503_ (.A0(net71),
    .A1(\i_random.rnd_out[11] ),
    .S(net121),
    .X(_032_));
 sg13g2_mux2_1 _504_ (.A0(net90),
    .A1(\i_random.rnd_out[12] ),
    .S(net122),
    .X(_033_));
 sg13g2_mux2_1 _505_ (.A0(net76),
    .A1(\i_random.rnd_out[13] ),
    .S(net121),
    .X(_034_));
 sg13g2_mux2_1 _506_ (.A0(net101),
    .A1(\i_random.rnd_out[14] ),
    .S(net121),
    .X(_035_));
 sg13g2_mux2_1 _507_ (.A0(net175),
    .A1(\i_random.rnd_out[15] ),
    .S(net122),
    .X(_036_));
 sg13g2_mux2_1 _508_ (.A0(net103),
    .A1(\i_random.rnd_out[16] ),
    .S(net121),
    .X(_037_));
 sg13g2_mux2_1 _509_ (.A0(net94),
    .A1(\i_random.rnd_out[17] ),
    .S(net121),
    .X(_038_));
 sg13g2_mux2_1 _510_ (.A0(net163),
    .A1(\i_random.rnd_out[18] ),
    .S(net121),
    .X(_039_));
 sg13g2_mux2_1 _511_ (.A0(net88),
    .A1(\i_random.rnd_out[19] ),
    .S(net121),
    .X(_040_));
 sg13g2_mux2_1 _512_ (.A0(net167),
    .A1(\i_random.rnd_out[20] ),
    .S(net121),
    .X(_041_));
 sg13g2_mux2_1 _513_ (.A0(net173),
    .A1(\i_random.rnd_out[21] ),
    .S(net122),
    .X(_042_));
 sg13g2_mux2_1 _514_ (.A0(net169),
    .A1(\i_random.rnd_out[22] ),
    .S(net122),
    .X(_043_));
 sg13g2_mux2_1 _515_ (.A0(net157),
    .A1(\i_random.rnd_out[23] ),
    .S(net125),
    .X(_044_));
 sg13g2_mux2_1 _516_ (.A0(net96),
    .A1(\i_random.rnd_out[24] ),
    .S(net125),
    .X(_045_));
 sg13g2_mux2_1 _517_ (.A0(net165),
    .A1(\i_random.rnd_out[25] ),
    .S(net125),
    .X(_046_));
 sg13g2_mux2_1 _518_ (.A0(net192),
    .A1(\i_random.rnd_out[26] ),
    .S(net125),
    .X(_047_));
 sg13g2_mux2_1 _519_ (.A0(net219),
    .A1(net198),
    .S(net125),
    .X(_048_));
 sg13g2_mux2_1 _520_ (.A0(net109),
    .A1(\i_random.rnd_out[28] ),
    .S(net126),
    .X(_049_));
 sg13g2_mux2_1 _521_ (.A0(net107),
    .A1(\i_random.rnd_out[29] ),
    .S(net125),
    .X(_050_));
 sg13g2_mux2_1 _522_ (.A0(net177),
    .A1(\i_random.rnd_out[30] ),
    .S(net125),
    .X(_051_));
 sg13g2_mux2_1 _523_ (.A0(net161),
    .A1(\i_random.rnd_out[31] ),
    .S(net125),
    .X(_052_));
 sg13g2_nand2b_1 _524_ (.Y(_205_),
    .B(net1),
    .A_N(\i_random.state ));
 sg13g2_mux2_1 _525_ (.A0(net98),
    .A1(net229),
    .S(_205_),
    .X(_053_));
 sg13g2_mux2_1 _526_ (.A0(\i_random.state ),
    .A1(net47),
    .S(net1),
    .X(_054_));
 sg13g2_nand2_1 _527_ (.Y(_206_),
    .A(\i_random.state ),
    .B(net145));
 sg13g2_a21oi_1 _528_ (.A1(net98),
    .A2(\i_random.first_bit ),
    .Y(_207_),
    .B1(_206_));
 sg13g2_o21ai_1 _529_ (.B1(_207_),
    .Y(_208_),
    .A1(net98),
    .A2(\i_random.first_bit ));
 sg13g2_a22oi_1 _530_ (.Y(_055_),
    .B1(_208_),
    .B2(_124_),
    .A2(_207_),
    .A1(net98));
 sg13g2_and2_1 _531_ (.A(net145),
    .B(\i_random.debiased_bit_valid ),
    .X(_209_));
 sg13g2_nand2_1 _532_ (.Y(_210_),
    .A(net145),
    .B(\i_random.debiased_bit_valid ));
 sg13g2_xnor2_1 _533_ (.Y(_056_),
    .A(net100),
    .B(net115));
 sg13g2_nand3_1 _534_ (.B(net100),
    .C(_209_),
    .A(net254),
    .Y(_211_));
 sg13g2_a21o_1 _535_ (.A2(_209_),
    .A1(net100),
    .B1(net254),
    .X(_212_));
 sg13g2_and2_1 _536_ (.A(_211_),
    .B(_212_),
    .X(_057_));
 sg13g2_nor2_1 _537_ (.A(_121_),
    .B(_211_),
    .Y(_213_));
 sg13g2_xnor2_1 _538_ (.Y(_058_),
    .A(net51),
    .B(_211_));
 sg13g2_xor2_1 _539_ (.B(_213_),
    .A(net82),
    .X(_059_));
 sg13g2_nand3_1 _540_ (.B(net255),
    .C(_213_),
    .A(net82),
    .Y(_214_));
 sg13g2_a21o_1 _541_ (.A2(_213_),
    .A1(net82),
    .B1(net255),
    .X(_215_));
 sg13g2_and2_1 _542_ (.A(_214_),
    .B(_215_),
    .X(_060_));
 sg13g2_o21ai_1 _543_ (.B1(_214_),
    .Y(_061_),
    .A1(net145),
    .A2(_115_));
 sg13g2_nand2_1 _544_ (.Y(_216_),
    .A(net53),
    .B(net116));
 sg13g2_o21ai_1 _545_ (.B1(_216_),
    .Y(_062_),
    .A1(_124_),
    .A2(net116));
 sg13g2_mux2_1 _546_ (.A0(net53),
    .A1(net62),
    .S(net116),
    .X(_063_));
 sg13g2_mux2_1 _547_ (.A0(net62),
    .A1(net196),
    .S(net116),
    .X(_064_));
 sg13g2_mux2_1 _548_ (.A0(net196),
    .A1(net55),
    .S(net115),
    .X(_065_));
 sg13g2_mux2_1 _549_ (.A0(net55),
    .A1(net222),
    .S(net116),
    .X(_066_));
 sg13g2_mux2_1 _550_ (.A0(net222),
    .A1(net92),
    .S(net115),
    .X(_067_));
 sg13g2_mux2_1 _551_ (.A0(net92),
    .A1(net69),
    .S(net115),
    .X(_068_));
 sg13g2_mux2_1 _552_ (.A0(net69),
    .A1(net231),
    .S(net115),
    .X(_069_));
 sg13g2_mux2_1 _553_ (.A0(net231),
    .A1(net218),
    .S(net115),
    .X(_070_));
 sg13g2_mux2_1 _554_ (.A0(net218),
    .A1(net214),
    .S(net115),
    .X(_071_));
 sg13g2_mux2_1 _555_ (.A0(net214),
    .A1(\i_random.rnd_out[10] ),
    .S(net115),
    .X(_072_));
 sg13g2_mux2_1 _556_ (.A0(\i_random.rnd_out[10] ),
    .A1(net206),
    .S(net113),
    .X(_073_));
 sg13g2_mux2_1 _557_ (.A0(net206),
    .A1(net216),
    .S(net113),
    .X(_074_));
 sg13g2_mux2_1 _558_ (.A0(net216),
    .A1(net226),
    .S(net112),
    .X(_075_));
 sg13g2_mux2_1 _559_ (.A0(net226),
    .A1(net237),
    .S(net112),
    .X(_076_));
 sg13g2_mux2_1 _560_ (.A0(net237),
    .A1(net238),
    .S(net112),
    .X(_077_));
 sg13g2_mux2_1 _561_ (.A0(net238),
    .A1(net217),
    .S(net113),
    .X(_078_));
 sg13g2_mux2_1 _562_ (.A0(net217),
    .A1(net197),
    .S(net113),
    .X(_079_));
 sg13g2_mux2_1 _563_ (.A0(net197),
    .A1(net194),
    .S(net113),
    .X(_080_));
 sg13g2_mux2_1 _564_ (.A0(net194),
    .A1(\i_random.rnd_out[19] ),
    .S(net112),
    .X(_081_));
 sg13g2_mux2_1 _565_ (.A0(net202),
    .A1(\i_random.rnd_out[20] ),
    .S(net112),
    .X(_082_));
 sg13g2_mux2_1 _566_ (.A0(net223),
    .A1(net200),
    .S(net112),
    .X(_083_));
 sg13g2_mux2_1 _567_ (.A0(net200),
    .A1(\i_random.rnd_out[22] ),
    .S(net112),
    .X(_084_));
 sg13g2_mux2_1 _568_ (.A0(net211),
    .A1(net184),
    .S(net112),
    .X(_085_));
 sg13g2_mux2_1 _569_ (.A0(net184),
    .A1(\i_random.rnd_out[24] ),
    .S(net114),
    .X(_086_));
 sg13g2_mux2_1 _570_ (.A0(net212),
    .A1(\i_random.rnd_out[25] ),
    .S(net117),
    .X(_087_));
 sg13g2_mux2_1 _571_ (.A0(net232),
    .A1(net205),
    .S(net117),
    .X(_088_));
 sg13g2_mux2_1 _572_ (.A0(net205),
    .A1(net198),
    .S(net114),
    .X(_089_));
 sg13g2_mux2_1 _573_ (.A0(net198),
    .A1(\i_random.rnd_out[28] ),
    .S(net114),
    .X(_090_));
 sg13g2_mux2_1 _574_ (.A0(net233),
    .A1(net220),
    .S(net114),
    .X(_091_));
 sg13g2_mux2_1 _575_ (.A0(net220),
    .A1(\i_random.rnd_out[30] ),
    .S(net114),
    .X(_092_));
 sg13g2_mux2_1 _576_ (.A0(\i_random.rnd_out[30] ),
    .A1(net227),
    .S(net114),
    .X(_093_));
 sg13g2_a21oi_1 _577_ (.A1(fsm_state_r),
    .A2(_125_),
    .Y(_217_),
    .B1(net126));
 sg13g2_a21oi_1 _578_ (.A1(uart_tx_en_next),
    .A2(_129_),
    .Y(_218_),
    .B1(_217_));
 sg13g2_a21oi_1 _579_ (.A1(fsm_state_r),
    .A2(_125_),
    .Y(_219_),
    .B1(net242));
 sg13g2_a21oi_1 _580_ (.A1(net242),
    .A2(_218_),
    .Y(_094_),
    .B1(_219_));
 sg13g2_nand2b_1 _581_ (.Y(_220_),
    .B(net244),
    .A_N(_218_));
 sg13g2_or2_1 _582_ (.X(_221_),
    .B(net119),
    .A(_129_));
 sg13g2_o21ai_1 _583_ (.B1(_220_),
    .Y(_095_),
    .A1(_131_),
    .A2(_221_));
 sg13g2_a21oi_1 _584_ (.A1(net84),
    .A2(_140_),
    .Y(_222_),
    .B1(_171_));
 sg13g2_nor2_1 _585_ (.A(_113_),
    .B(net85),
    .Y(_096_));
 sg13g2_nor2_1 _586_ (.A(net49),
    .B(_148_),
    .Y(_223_));
 sg13g2_nand2_1 _587_ (.Y(_224_),
    .A(net127),
    .B(net143));
 sg13g2_a21o_1 _588_ (.A2(_142_),
    .A1(_112_),
    .B1(_224_),
    .X(_225_));
 sg13g2_nor2b_1 _589_ (.A(\i_uart_tx.bit_counter[0] ),
    .B_N(_148_),
    .Y(_226_));
 sg13g2_nor3_1 _590_ (.A(_223_),
    .B(_225_),
    .C(_226_),
    .Y(_097_));
 sg13g2_nand3_1 _591_ (.B(net127),
    .C(_138_),
    .A(\i_uart_tx.bit_counter[0] ),
    .Y(_227_));
 sg13g2_nor2b_1 _592_ (.A(net190),
    .B_N(_227_),
    .Y(_228_));
 sg13g2_and4_1 _593_ (.A(net190),
    .B(\i_uart_tx.bit_counter[0] ),
    .C(net127),
    .D(_138_),
    .X(_229_));
 sg13g2_nor3_1 _594_ (.A(_225_),
    .B(net191),
    .C(_229_),
    .Y(_098_));
 sg13g2_nor2_1 _595_ (.A(net252),
    .B(_229_),
    .Y(_230_));
 sg13g2_a21oi_1 _596_ (.A1(net252),
    .A2(_229_),
    .Y(_231_),
    .B1(_225_));
 sg13g2_nor2b_1 _597_ (.A(net253),
    .B_N(_231_),
    .Y(_099_));
 sg13g2_a21oi_1 _598_ (.A1(\i_uart_tx.bit_counter[2] ),
    .A2(_229_),
    .Y(_232_),
    .B1(net187));
 sg13g2_and3_1 _599_ (.X(_233_),
    .A(net187),
    .B(\i_uart_tx.bit_counter[2] ),
    .C(_229_));
 sg13g2_nor3_1 _600_ (.A(_225_),
    .B(net188),
    .C(_233_),
    .Y(_100_));
 sg13g2_nand2_2 _601_ (.Y(_234_),
    .A(net142),
    .B(_139_));
 sg13g2_nand2_1 _602_ (.Y(_235_),
    .A(net45),
    .B(_126_));
 sg13g2_nand2_1 _603_ (.Y(_236_),
    .A(\i_uart_tx.cycle_counter[0] ),
    .B(_125_));
 sg13g2_a21oi_1 _604_ (.A1(_235_),
    .A2(_236_),
    .Y(_101_),
    .B1(_234_));
 sg13g2_and3_1 _605_ (.X(_237_),
    .A(net148),
    .B(\i_uart_tx.cycle_counter[0] ),
    .C(_126_));
 sg13g2_a21oi_1 _606_ (.A1(\i_uart_tx.cycle_counter[0] ),
    .A2(_126_),
    .Y(_238_),
    .B1(net148));
 sg13g2_nor3_1 _607_ (.A(_234_),
    .B(_237_),
    .C(net149),
    .Y(_102_));
 sg13g2_nor2_1 _608_ (.A(net246),
    .B(_237_),
    .Y(_239_));
 sg13g2_and2_1 _609_ (.A(net246),
    .B(_237_),
    .X(_240_));
 sg13g2_nor3_1 _610_ (.A(_234_),
    .B(net247),
    .C(_240_),
    .Y(_103_));
 sg13g2_nor2_1 _611_ (.A(net251),
    .B(_240_),
    .Y(_241_));
 sg13g2_and3_1 _612_ (.X(_242_),
    .A(net251),
    .B(net246),
    .C(_237_));
 sg13g2_nor3_1 _613_ (.A(_234_),
    .B(_241_),
    .C(_242_),
    .Y(_104_));
 sg13g2_xnor2_1 _614_ (.Y(_243_),
    .A(net224),
    .B(_242_));
 sg13g2_nor2_1 _615_ (.A(_234_),
    .B(net225),
    .Y(_105_));
 sg13g2_a21oi_1 _616_ (.A1(\i_uart_tx.cycle_counter[4] ),
    .A2(_242_),
    .Y(_244_),
    .B1(net59));
 sg13g2_nand4_1 _617_ (.B(net246),
    .C(_135_),
    .A(\i_uart_tx.cycle_counter[3] ),
    .Y(_245_),
    .D(_237_));
 sg13g2_inv_1 _618_ (.Y(_246_),
    .A(_245_));
 sg13g2_nor3_1 _619_ (.A(_234_),
    .B(net60),
    .C(_246_),
    .Y(_106_));
 sg13g2_xor2_1 _620_ (.B(_245_),
    .A(net248),
    .X(_247_));
 sg13g2_nor2_1 _621_ (.A(_234_),
    .B(net249),
    .Y(_107_));
 sg13g2_o21ai_1 _622_ (.B1(_208_),
    .Y(_108_),
    .A1(net145),
    .A2(_114_));
 sg13g2_nor2b_1 _623_ (.A(net186),
    .B_N(_146_),
    .Y(_248_));
 sg13g2_o21ai_1 _624_ (.B1(net142),
    .Y(_109_),
    .A1(_144_),
    .A2(_248_));
 sg13g2_dfrbp_1 _625_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net22),
    .D(_004_),
    .Q_N(_350_),
    .Q(\i_uart_tx.fsm_state[0] ));
 sg13g2_dfrbp_1 _626_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net36),
    .D(_005_),
    .Q_N(_349_),
    .Q(\i_uart_tx.fsm_state[1] ));
 sg13g2_dfrbp_1 _627_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net35),
    .D(_006_),
    .Q_N(_348_),
    .Q(\i_uart_tx.data_to_send[0] ));
 sg13g2_dfrbp_1 _628_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net33),
    .D(net183),
    .Q_N(_347_),
    .Q(\i_uart_tx.data_to_send[1] ));
 sg13g2_dfrbp_1 _629_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net32),
    .D(net106),
    .Q_N(_346_),
    .Q(\i_uart_tx.data_to_send[2] ));
 sg13g2_dfrbp_1 _630_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net30),
    .D(_009_),
    .Q_N(_345_),
    .Q(\i_uart_tx.data_to_send[3] ));
 sg13g2_dfrbp_1 _631_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net28),
    .D(net240),
    .Q_N(_344_),
    .Q(\i_uart_tx.data_to_send[4] ));
 sg13g2_dfrbp_1 _632_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net26),
    .D(net81),
    .Q_N(_343_),
    .Q(\i_uart_tx.data_to_send[5] ));
 sg13g2_dfrbp_1 _633_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net23),
    .D(net236),
    .Q_N(_351_),
    .Q(\i_uart_tx.data_to_send[6] ));
 sg13g2_dfrbp_1 _634_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net143),
    .D(uart_tx_en_next),
    .Q_N(_342_),
    .Q(\i_uart_tx.uart_tx_en ));
 sg13g2_dfrbp_1 _635_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net141),
    .D(net172),
    .Q_N(_341_),
    .Q(\i_uart_tx.uart_tx_data[0] ));
 sg13g2_dfrbp_1 _636_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net141),
    .D(net156),
    .Q_N(_340_),
    .Q(\i_uart_tx.uart_tx_data[1] ));
 sg13g2_dfrbp_1 _637_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net139),
    .D(net209),
    .Q_N(_339_),
    .Q(\i_uart_tx.uart_tx_data[2] ));
 sg13g2_dfrbp_1 _638_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net140),
    .D(net74),
    .Q_N(_338_),
    .Q(\i_uart_tx.uart_tx_data[3] ));
 sg13g2_dfrbp_1 _639_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net139),
    .D(_017_),
    .Q_N(_337_),
    .Q(\i_uart_tx.uart_tx_data[4] ));
 sg13g2_dfrbp_1 _640_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net140),
    .D(net79),
    .Q_N(_336_),
    .Q(\i_uart_tx.uart_tx_data[5] ));
 sg13g2_dfrbp_1 _641_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net140),
    .D(net58),
    .Q_N(_335_),
    .Q(\i_uart_tx.uart_tx_data[6] ));
 sg13g2_dfrbp_1 _642_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net139),
    .D(_020_),
    .Q_N(_352_),
    .Q(\i_uart_tx.uart_tx_data[7] ));
 sg13g2_dfrbp_1 _643_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net141),
    .D(fsm_state_next),
    .Q_N(_001_),
    .Q(fsm_state_r));
 sg13g2_dfrbp_1 _644_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net141),
    .D(net54),
    .Q_N(_334_),
    .Q(\random_buffer_r[0] ));
 sg13g2_dfrbp_1 _645_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net135),
    .D(net64),
    .Q_N(_333_),
    .Q(\random_buffer_r[1] ));
 sg13g2_dfrbp_1 _646_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net135),
    .D(net160),
    .Q_N(_332_),
    .Q(\random_buffer_r[2] ));
 sg13g2_dfrbp_1 _647_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net135),
    .D(net56),
    .Q_N(_331_),
    .Q(\random_buffer_r[3] ));
 sg13g2_dfrbp_1 _648_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net135),
    .D(net147),
    .Q_N(_330_),
    .Q(\random_buffer_r[4] ));
 sg13g2_dfrbp_1 _649_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net131),
    .D(net93),
    .Q_N(_329_),
    .Q(\random_buffer_r[5] ));
 sg13g2_dfrbp_1 _650_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net131),
    .D(net70),
    .Q_N(_328_),
    .Q(\random_buffer_r[6] ));
 sg13g2_dfrbp_1 _651_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net135),
    .D(net180),
    .Q_N(_327_),
    .Q(\random_buffer_r[7] ));
 sg13g2_dfrbp_1 _652_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net133),
    .D(net87),
    .Q_N(_326_),
    .Q(\random_buffer_r[8] ));
 sg13g2_dfrbp_1 _653_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net132),
    .D(net66),
    .Q_N(_325_),
    .Q(\random_buffer_r[9] ));
 sg13g2_dfrbp_1 _654_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net131),
    .D(net152),
    .Q_N(_324_),
    .Q(\random_buffer_r[10] ));
 sg13g2_dfrbp_1 _655_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net128),
    .D(net72),
    .Q_N(_323_),
    .Q(\random_buffer_r[11] ));
 sg13g2_dfrbp_1 _656_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net131),
    .D(net91),
    .Q_N(_322_),
    .Q(\random_buffer_r[12] ));
 sg13g2_dfrbp_1 _657_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net130),
    .D(net77),
    .Q_N(_321_),
    .Q(\random_buffer_r[13] ));
 sg13g2_dfrbp_1 _658_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net130),
    .D(net102),
    .Q_N(_320_),
    .Q(\random_buffer_r[14] ));
 sg13g2_dfrbp_1 _659_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net131),
    .D(net176),
    .Q_N(_319_),
    .Q(\random_buffer_r[15] ));
 sg13g2_dfrbp_1 _660_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net132),
    .D(net104),
    .Q_N(_318_),
    .Q(\random_buffer_r[16] ));
 sg13g2_dfrbp_1 _661_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net128),
    .D(net95),
    .Q_N(_317_),
    .Q(\random_buffer_r[17] ));
 sg13g2_dfrbp_1 _662_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net128),
    .D(net164),
    .Q_N(_316_),
    .Q(\random_buffer_r[18] ));
 sg13g2_dfrbp_1 _663_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net129),
    .D(net89),
    .Q_N(_315_),
    .Q(\random_buffer_r[19] ));
 sg13g2_dfrbp_1 _664_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net130),
    .D(net168),
    .Q_N(_314_),
    .Q(\random_buffer_r[20] ));
 sg13g2_dfrbp_1 _665_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net130),
    .D(net174),
    .Q_N(_313_),
    .Q(\random_buffer_r[21] ));
 sg13g2_dfrbp_1 _666_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net130),
    .D(net170),
    .Q_N(_312_),
    .Q(\random_buffer_r[22] ));
 sg13g2_dfrbp_1 _667_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net130),
    .D(net158),
    .Q_N(_311_),
    .Q(\random_buffer_r[23] ));
 sg13g2_dfrbp_1 _668_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net137),
    .D(net97),
    .Q_N(_310_),
    .Q(\random_buffer_r[24] ));
 sg13g2_dfrbp_1 _669_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net137),
    .D(net166),
    .Q_N(_309_),
    .Q(\random_buffer_r[25] ));
 sg13g2_dfrbp_1 _670_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net137),
    .D(net193),
    .Q_N(_308_),
    .Q(\random_buffer_r[26] ));
 sg13g2_dfrbp_1 _671_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net137),
    .D(_048_),
    .Q_N(_307_),
    .Q(\random_buffer_r[27] ));
 sg13g2_dfrbp_1 _672_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net138),
    .D(net110),
    .Q_N(_306_),
    .Q(\random_buffer_r[28] ));
 sg13g2_dfrbp_1 _673_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net138),
    .D(net108),
    .Q_N(_305_),
    .Q(\random_buffer_r[29] ));
 sg13g2_dfrbp_1 _674_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net137),
    .D(net178),
    .Q_N(_304_),
    .Q(\random_buffer_r[30] ));
 sg13g2_dfrbp_1 _675_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net137),
    .D(net162),
    .Q_N(_303_),
    .Q(\random_buffer_r[31] ));
 sg13g2_dfrbp_1 _676_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net141),
    .D(net230),
    .Q_N(_302_),
    .Q(\i_random.first_bit ));
 sg13g2_dfrbp_1 _677_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net141),
    .D(net48),
    .Q_N(_000_),
    .Q(\i_random.state ));
 sg13g2_dfrbp_1 _678_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net142),
    .D(net99),
    .Q_N(_301_),
    .Q(\i_random.debiased_bit ));
 sg13g2_dfrbp_1 _679_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(_056_),
    .Q_N(_300_),
    .Q(\i_random.bit_count[0] ));
 sg13g2_dfrbp_1 _680_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net133),
    .D(_057_),
    .Q_N(_299_),
    .Q(\i_random.bit_count[1] ));
 sg13g2_dfrbp_1 _681_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(net52),
    .Q_N(_298_),
    .Q(\i_random.bit_count[2] ));
 sg13g2_dfrbp_1 _682_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net134),
    .D(net83),
    .Q_N(_297_),
    .Q(\i_random.bit_count[3] ));
 sg13g2_dfrbp_1 _683_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net134),
    .D(_060_),
    .Q_N(_353_),
    .Q(\i_random.bit_count[4] ));
 sg13g2_dfrbp_1 _684_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net135),
    .D(\i_random.combined_ring_bit ),
    .Q_N(_296_),
    .Q(\i_random.sync1 ));
 sg13g2_dfrbp_1 _685_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net136),
    .D(net68),
    .Q_N(_295_),
    .Q(\i_random.ready ));
 sg13g2_dfrbp_1 _686_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net142),
    .D(_062_),
    .Q_N(_294_),
    .Q(\i_random.rnd_out[0] ));
 sg13g2_dfrbp_1 _687_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net136),
    .D(_063_),
    .Q_N(_293_),
    .Q(\i_random.rnd_out[1] ));
 sg13g2_dfrbp_1 _688_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net135),
    .D(_064_),
    .Q_N(_292_),
    .Q(\i_random.rnd_out[2] ));
 sg13g2_dfrbp_1 _689_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net135),
    .D(_065_),
    .Q_N(_291_),
    .Q(\i_random.rnd_out[3] ));
 sg13g2_dfrbp_1 _690_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net133),
    .D(_066_),
    .Q_N(_290_),
    .Q(\i_random.rnd_out[4] ));
 sg13g2_dfrbp_1 _691_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net133),
    .D(_067_),
    .Q_N(_289_),
    .Q(\i_random.rnd_out[5] ));
 sg13g2_dfrbp_1 _692_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net133),
    .D(_068_),
    .Q_N(_288_),
    .Q(\i_random.rnd_out[6] ));
 sg13g2_dfrbp_1 _693_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net133),
    .D(_069_),
    .Q_N(_287_),
    .Q(\i_random.rnd_out[7] ));
 sg13g2_dfrbp_1 _694_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net133),
    .D(_070_),
    .Q_N(_286_),
    .Q(\i_random.rnd_out[8] ));
 sg13g2_dfrbp_1 _695_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net133),
    .D(_071_),
    .Q_N(_285_),
    .Q(\i_random.rnd_out[9] ));
 sg13g2_dfrbp_1 _696_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net128),
    .D(net215),
    .Q_N(_284_),
    .Q(\i_random.rnd_out[10] ));
 sg13g2_dfrbp_1 _697_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net128),
    .D(net207),
    .Q_N(_283_),
    .Q(\i_random.rnd_out[11] ));
 sg13g2_dfrbp_1 _698_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net128),
    .D(_074_),
    .Q_N(_282_),
    .Q(\i_random.rnd_out[12] ));
 sg13g2_dfrbp_1 _699_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net129),
    .D(_075_),
    .Q_N(_281_),
    .Q(\i_random.rnd_out[13] ));
 sg13g2_dfrbp_1 _700_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net129),
    .D(_076_),
    .Q_N(_280_),
    .Q(\i_random.rnd_out[14] ));
 sg13g2_dfrbp_1 _701_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net129),
    .D(_077_),
    .Q_N(_279_),
    .Q(\i_random.rnd_out[15] ));
 sg13g2_dfrbp_1 _702_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net128),
    .D(_078_),
    .Q_N(_278_),
    .Q(\i_random.rnd_out[16] ));
 sg13g2_dfrbp_1 _703_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net128),
    .D(_079_),
    .Q_N(_277_),
    .Q(\i_random.rnd_out[17] ));
 sg13g2_dfrbp_1 _704_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net129),
    .D(_080_),
    .Q_N(_276_),
    .Q(\i_random.rnd_out[18] ));
 sg13g2_dfrbp_1 _705_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net129),
    .D(net195),
    .Q_N(_275_),
    .Q(\i_random.rnd_out[19] ));
 sg13g2_dfrbp_1 _706_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net129),
    .D(net203),
    .Q_N(_274_),
    .Q(\i_random.rnd_out[20] ));
 sg13g2_dfrbp_1 _707_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net129),
    .D(_083_),
    .Q_N(_273_),
    .Q(\i_random.rnd_out[21] ));
 sg13g2_dfrbp_1 _708_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net130),
    .D(net201),
    .Q_N(_272_),
    .Q(\i_random.rnd_out[22] ));
 sg13g2_dfrbp_1 _709_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net130),
    .D(_085_),
    .Q_N(_271_),
    .Q(\i_random.rnd_out[23] ));
 sg13g2_dfrbp_1 _710_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net131),
    .D(net185),
    .Q_N(_270_),
    .Q(\i_random.rnd_out[24] ));
 sg13g2_dfrbp_1 _711_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net137),
    .D(net213),
    .Q_N(_269_),
    .Q(\i_random.rnd_out[25] ));
 sg13g2_dfrbp_1 _712_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net137),
    .D(_088_),
    .Q_N(_268_),
    .Q(\i_random.rnd_out[26] ));
 sg13g2_dfrbp_1 _713_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net138),
    .D(_089_),
    .Q_N(_267_),
    .Q(\i_random.rnd_out[27] ));
 sg13g2_dfrbp_1 _714_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net138),
    .D(net199),
    .Q_N(_266_),
    .Q(\i_random.rnd_out[28] ));
 sg13g2_dfrbp_1 _715_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net140),
    .D(_091_),
    .Q_N(_265_),
    .Q(\i_random.rnd_out[29] ));
 sg13g2_dfrbp_1 _716_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net144),
    .D(net221),
    .Q_N(_264_),
    .Q(\i_random.rnd_out[30] ));
 sg13g2_dfrbp_1 _717_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net140),
    .D(net228),
    .Q_N(_354_),
    .Q(\i_random.rnd_out[31] ));
 sg13g2_dfrbp_1 _718_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net142),
    .D(net44),
    .Q_N(_263_),
    .Q(\i_random.rnd_sync ));
 sg13g2_dfrbp_1 _719_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net141),
    .D(net243),
    .Q_N(_262_),
    .Q(\byte_counter_r[0] ));
 sg13g2_dfrbp_1 _720_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net141),
    .D(net245),
    .Q_N(_261_),
    .Q(\byte_counter_r[1] ));
 sg13g2_dfrbp_1 _721_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net43),
    .D(_096_),
    .Q_N(_260_),
    .Q(\i_uart_tx.data_to_send[7] ));
 sg13g2_dfrbp_1 _722_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net41),
    .D(net50),
    .Q_N(_003_),
    .Q(\i_uart_tx.bit_counter[0] ));
 sg13g2_dfrbp_1 _723_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net39),
    .D(_098_),
    .Q_N(_259_),
    .Q(\i_uart_tx.bit_counter[1] ));
 sg13g2_dfrbp_1 _724_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net38),
    .D(_099_),
    .Q_N(_258_),
    .Q(\i_uart_tx.bit_counter[2] ));
 sg13g2_dfrbp_1 _725_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net34),
    .D(net189),
    .Q_N(_257_),
    .Q(\i_uart_tx.bit_counter[3] ));
 sg13g2_dfrbp_1 _726_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net31),
    .D(net46),
    .Q_N(_002_),
    .Q(\i_uart_tx.cycle_counter[0] ));
 sg13g2_dfrbp_1 _727_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net27),
    .D(net150),
    .Q_N(_256_),
    .Q(\i_uart_tx.cycle_counter[1] ));
 sg13g2_dfrbp_1 _728_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net24),
    .D(_103_),
    .Q_N(_255_),
    .Q(\i_uart_tx.cycle_counter[2] ));
 sg13g2_dfrbp_1 _729_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net40),
    .D(_104_),
    .Q_N(_254_),
    .Q(\i_uart_tx.cycle_counter[3] ));
 sg13g2_dfrbp_1 _730_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net37),
    .D(_105_),
    .Q_N(_253_),
    .Q(\i_uart_tx.cycle_counter[4] ));
 sg13g2_dfrbp_1 _731_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net29),
    .D(net61),
    .Q_N(_252_),
    .Q(\i_uart_tx.cycle_counter[5] ));
 sg13g2_dfrbp_1 _732_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net42),
    .D(_107_),
    .Q_N(_251_),
    .Q(\i_uart_tx.cycle_counter[6] ));
 sg13g2_dfrbp_1 _733_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net136),
    .D(net154),
    .Q_N(_250_),
    .Q(\i_random.debiased_bit_valid ));
 sg13g2_dfrbp_1 _734_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net25),
    .D(_109_),
    .Q_N(_249_),
    .Q(\i_uart_tx.txd_reg ));
 sg13g2_tiehi _633__23 (.L_HI(net23));
 sg13g2_tiehi _728__24 (.L_HI(net24));
 sg13g2_tiehi _734__25 (.L_HI(net25));
 sg13g2_tiehi _632__26 (.L_HI(net26));
 sg13g2_tiehi _727__27 (.L_HI(net27));
 sg13g2_tiehi _631__28 (.L_HI(net28));
 sg13g2_tiehi _731__29 (.L_HI(net29));
 sg13g2_tiehi _630__30 (.L_HI(net30));
 sg13g2_tiehi _726__31 (.L_HI(net31));
 sg13g2_tiehi _629__32 (.L_HI(net32));
 sg13g2_tiehi _628__33 (.L_HI(net33));
 sg13g2_tiehi _725__34 (.L_HI(net34));
 sg13g2_tiehi _627__35 (.L_HI(net35));
 sg13g2_tiehi _626__36 (.L_HI(net36));
 sg13g2_tiehi _730__37 (.L_HI(net37));
 sg13g2_tiehi _724__38 (.L_HI(net38));
 sg13g2_tiehi _723__39 (.L_HI(net39));
 sg13g2_tiehi _729__40 (.L_HI(net40));
 sg13g2_tiehi _722__41 (.L_HI(net41));
 sg13g2_tiehi _732__42 (.L_HI(net42));
 sg13g2_tiehi _721__43 (.L_HI(net43));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_Xelef2000_3 (.L_LO(net3));
 sg13g2_tielo tt_um_Xelef2000_4 (.L_LO(net4));
 sg13g2_tielo tt_um_Xelef2000_5 (.L_LO(net5));
 sg13g2_tielo tt_um_Xelef2000_6 (.L_LO(net6));
 sg13g2_tielo tt_um_Xelef2000_7 (.L_LO(net7));
 sg13g2_tielo tt_um_Xelef2000_8 (.L_LO(net8));
 sg13g2_tielo tt_um_Xelef2000_9 (.L_LO(net9));
 sg13g2_tielo tt_um_Xelef2000_10 (.L_LO(net10));
 sg13g2_tielo tt_um_Xelef2000_11 (.L_LO(net11));
 sg13g2_tielo tt_um_Xelef2000_12 (.L_LO(net12));
 sg13g2_tielo tt_um_Xelef2000_13 (.L_LO(net13));
 sg13g2_tielo tt_um_Xelef2000_14 (.L_LO(net14));
 sg13g2_tielo tt_um_Xelef2000_15 (.L_LO(net15));
 sg13g2_tielo tt_um_Xelef2000_16 (.L_LO(net16));
 sg13g2_tielo tt_um_Xelef2000_17 (.L_LO(net17));
 sg13g2_tielo tt_um_Xelef2000_18 (.L_LO(net18));
 sg13g2_tielo tt_um_Xelef2000_19 (.L_LO(net19));
 sg13g2_tielo tt_um_Xelef2000_20 (.L_LO(net20));
 sg13g2_tielo tt_um_Xelef2000_21 (.L_LO(net21));
 sg13g2_tiehi _625__22 (.L_HI(net22));
 sg13g2_buf_1 _777_ (.A(\i_uart_tx.txd_reg ),
    .X(uo_out[0]));
 sg13g2_buf_1 _778_ (.A(\i_random.ring_bit_6 ),
    .X(uo_out[1]));
 sg13g2_buf_1 _779_ (.A(\i_random.ring_bit_12 ),
    .X(uo_out[2]));
 sg13g2_buf_1 _780_ (.A(\i_random.ring_bit_24 ),
    .X(uo_out[3]));
 sg13g2_nand2_1 \i_random.u_ring12.u0  (.Y(\i_random.u_ring12.gated ),
    .A(\i_random.ring_bit_12 ),
    .B(net145));
 sg13g2_inv_2 \i_random.u_ring12.u1  (.Y(\i_random.u_ring12.n1 ),
    .A(\i_random.u_ring12.gated ));
 sg13g2_inv_2 \i_random.u_ring12.u10  (.Y(\i_random.u_ring12.n10 ),
    .A(\i_random.u_ring12.n9 ));
 sg13g2_inv_2 \i_random.u_ring12.u11  (.Y(\i_random.ring_bit_12 ),
    .A(\i_random.u_ring12.n10 ));
 sg13g2_inv_2 \i_random.u_ring12.u2  (.Y(\i_random.u_ring12.n2 ),
    .A(\i_random.u_ring12.n1 ));
 sg13g2_inv_2 \i_random.u_ring12.u3  (.Y(\i_random.u_ring12.n3 ),
    .A(\i_random.u_ring12.n2 ));
 sg13g2_inv_2 \i_random.u_ring12.u4  (.Y(\i_random.u_ring12.n4 ),
    .A(\i_random.u_ring12.n3 ));
 sg13g2_inv_2 \i_random.u_ring12.u5  (.Y(\i_random.u_ring12.n5 ),
    .A(\i_random.u_ring12.n4 ));
 sg13g2_inv_2 \i_random.u_ring12.u6  (.Y(\i_random.u_ring12.n6 ),
    .A(\i_random.u_ring12.n5 ));
 sg13g2_inv_2 \i_random.u_ring12.u7  (.Y(\i_random.u_ring12.n7 ),
    .A(\i_random.u_ring12.n6 ));
 sg13g2_inv_2 \i_random.u_ring12.u8  (.Y(\i_random.u_ring12.n8 ),
    .A(\i_random.u_ring12.n7 ));
 sg13g2_inv_2 \i_random.u_ring12.u9  (.Y(\i_random.u_ring12.n9 ),
    .A(\i_random.u_ring12.n8 ));
 sg13g2_nand2_1 \i_random.u_ring24.u0  (.Y(\i_random.u_ring24.gated ),
    .A(\i_random.ring_bit_24 ),
    .B(net145));
 sg13g2_inv_2 \i_random.u_ring24.u1  (.Y(\i_random.u_ring24.n1 ),
    .A(\i_random.u_ring24.gated ));
 sg13g2_inv_2 \i_random.u_ring24.u10  (.Y(\i_random.u_ring24.n10 ),
    .A(\i_random.u_ring24.n9 ));
 sg13g2_inv_2 \i_random.u_ring24.u11  (.Y(\i_random.u_ring24.n11 ),
    .A(\i_random.u_ring24.n10 ));
 sg13g2_inv_2 \i_random.u_ring24.u12  (.Y(\i_random.u_ring24.n12 ),
    .A(\i_random.u_ring24.n11 ));
 sg13g2_inv_2 \i_random.u_ring24.u13  (.Y(\i_random.u_ring24.n13 ),
    .A(\i_random.u_ring24.n12 ));
 sg13g2_inv_2 \i_random.u_ring24.u14  (.Y(\i_random.u_ring24.n14 ),
    .A(\i_random.u_ring24.n13 ));
 sg13g2_inv_2 \i_random.u_ring24.u15  (.Y(\i_random.u_ring24.n15 ),
    .A(\i_random.u_ring24.n14 ));
 sg13g2_inv_2 \i_random.u_ring24.u16  (.Y(\i_random.u_ring24.n16 ),
    .A(\i_random.u_ring24.n15 ));
 sg13g2_inv_2 \i_random.u_ring24.u17  (.Y(\i_random.u_ring24.n17 ),
    .A(\i_random.u_ring24.n16 ));
 sg13g2_inv_2 \i_random.u_ring24.u18  (.Y(\i_random.u_ring24.n18 ),
    .A(\i_random.u_ring24.n17 ));
 sg13g2_inv_2 \i_random.u_ring24.u19  (.Y(\i_random.u_ring24.n19 ),
    .A(\i_random.u_ring24.n18 ));
 sg13g2_inv_2 \i_random.u_ring24.u2  (.Y(\i_random.u_ring24.n2 ),
    .A(\i_random.u_ring24.n1 ));
 sg13g2_inv_2 \i_random.u_ring24.u20  (.Y(\i_random.u_ring24.n20 ),
    .A(\i_random.u_ring24.n19 ));
 sg13g2_inv_2 \i_random.u_ring24.u21  (.Y(\i_random.u_ring24.n21 ),
    .A(\i_random.u_ring24.n20 ));
 sg13g2_inv_2 \i_random.u_ring24.u22  (.Y(\i_random.u_ring24.n22 ),
    .A(\i_random.u_ring24.n21 ));
 sg13g2_inv_2 \i_random.u_ring24.u23  (.Y(\i_random.ring_bit_24 ),
    .A(\i_random.u_ring24.n22 ));
 sg13g2_inv_2 \i_random.u_ring24.u3  (.Y(\i_random.u_ring24.n3 ),
    .A(\i_random.u_ring24.n2 ));
 sg13g2_inv_2 \i_random.u_ring24.u4  (.Y(\i_random.u_ring24.n4 ),
    .A(\i_random.u_ring24.n3 ));
 sg13g2_inv_2 \i_random.u_ring24.u5  (.Y(\i_random.u_ring24.n5 ),
    .A(\i_random.u_ring24.n4 ));
 sg13g2_inv_2 \i_random.u_ring24.u6  (.Y(\i_random.u_ring24.n6 ),
    .A(\i_random.u_ring24.n5 ));
 sg13g2_inv_2 \i_random.u_ring24.u7  (.Y(\i_random.u_ring24.n7 ),
    .A(\i_random.u_ring24.n6 ));
 sg13g2_inv_2 \i_random.u_ring24.u8  (.Y(\i_random.u_ring24.n8 ),
    .A(\i_random.u_ring24.n7 ));
 sg13g2_inv_2 \i_random.u_ring24.u9  (.Y(\i_random.u_ring24.n9 ),
    .A(\i_random.u_ring24.n8 ));
 sg13g2_nand2_1 \i_random.u_ring6.u0  (.Y(\i_random.u_ring6.gated ),
    .A(\i_random.ring_bit_6 ),
    .B(net145));
 sg13g2_inv_2 \i_random.u_ring6.u1  (.Y(\i_random.u_ring6.n1 ),
    .A(\i_random.u_ring6.gated ));
 sg13g2_inv_2 \i_random.u_ring6.u2  (.Y(\i_random.u_ring6.n2 ),
    .A(\i_random.u_ring6.n1 ));
 sg13g2_inv_2 \i_random.u_ring6.u3  (.Y(\i_random.u_ring6.n3 ),
    .A(\i_random.u_ring6.n2 ));
 sg13g2_inv_2 \i_random.u_ring6.u4  (.Y(\i_random.u_ring6.n4 ),
    .A(\i_random.u_ring6.n3 ));
 sg13g2_inv_2 \i_random.u_ring6.u5  (.Y(\i_random.ring_bit_6 ),
    .A(\i_random.u_ring6.n4 ));
 sg13g2_buf_2 fanout111 (.A(_141_),
    .X(net111));
 sg13g2_buf_4 fanout112 (.X(net112),
    .A(net114));
 sg13g2_buf_2 fanout113 (.A(net114),
    .X(net113));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(net117));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(net116));
 sg13g2_buf_2 fanout116 (.A(net117),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_210_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_173_),
    .X(net118));
 sg13g2_buf_1 fanout119 (.A(_173_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_129_),
    .X(net120));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(net124));
 sg13g2_buf_2 fanout122 (.A(net124),
    .X(net122));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(net124));
 sg13g2_buf_2 fanout124 (.A(_128_),
    .X(net124));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(net126));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(_128_));
 sg13g2_buf_2 fanout127 (.A(\i_uart_tx.fsm_state[1] ),
    .X(net127));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(net132));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(net132));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(net131));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(net132));
 sg13g2_buf_2 fanout132 (.A(rst_n),
    .X(net132));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(net136));
 sg13g2_buf_2 fanout134 (.A(net136),
    .X(net134));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net136));
 sg13g2_buf_2 fanout136 (.A(rst_n),
    .X(net136));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net139));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(net144));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(net142));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net144));
 sg13g2_buf_2 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(rst_n),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(net1),
    .X(net145));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_tielo tt_um_Xelef2000_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\i_random.sync1 ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold2 (.A(_002_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold3 (.A(_101_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold4 (.A(_000_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold5 (.A(_054_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold6 (.A(_003_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold7 (.A(_097_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold8 (.A(\i_random.bit_count[2] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold9 (.A(_058_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_random.rnd_out[0] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold11 (.A(_021_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_random.rnd_out[3] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold13 (.A(_024_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_uart_tx.uart_tx_data[6] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold15 (.A(_019_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_uart_tx.cycle_counter[5] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold17 (.A(_244_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold18 (.A(_106_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i_random.rnd_out[1] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold20 (.A(_201_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold21 (.A(_022_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold22 (.A(\random_buffer_r[9] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold23 (.A(_030_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i_random.ready ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold25 (.A(_061_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i_random.rnd_out[6] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold27 (.A(_027_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold28 (.A(\random_buffer_r[11] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold29 (.A(_032_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_uart_tx.uart_tx_data[3] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold31 (.A(_016_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_random.debiased_bit ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold33 (.A(\random_buffer_r[13] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold34 (.A(_034_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold35 (.A(\i_uart_tx.uart_tx_data[5] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold36 (.A(_018_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold37 (.A(\i_uart_tx.data_to_send[5] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold38 (.A(_011_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold39 (.A(\i_random.bit_count[3] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold40 (.A(_059_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold41 (.A(\i_uart_tx.uart_tx_data[7] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold42 (.A(_222_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold43 (.A(\random_buffer_r[8] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold44 (.A(_029_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold45 (.A(\random_buffer_r[19] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold46 (.A(_040_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold47 (.A(\random_buffer_r[12] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold48 (.A(_033_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold49 (.A(\i_random.rnd_out[5] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold50 (.A(_026_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold51 (.A(\random_buffer_r[17] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold52 (.A(_038_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold53 (.A(\random_buffer_r[24] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold54 (.A(_045_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold55 (.A(\i_random.rnd_sync ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold56 (.A(_055_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold57 (.A(\i_random.bit_count[0] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold58 (.A(\random_buffer_r[14] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold59 (.A(_035_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold60 (.A(\random_buffer_r[16] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold61 (.A(_037_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold62 (.A(\i_uart_tx.data_to_send[3] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold63 (.A(_008_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold64 (.A(\random_buffer_r[29] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold65 (.A(_050_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold66 (.A(\random_buffer_r[28] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold67 (.A(_049_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold68 (.A(\random_buffer_r[4] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold69 (.A(_025_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_uart_tx.cycle_counter[1] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold71 (.A(_238_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold72 (.A(_102_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold73 (.A(\random_buffer_r[10] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold74 (.A(_031_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold75 (.A(\i_random.debiased_bit_valid ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold76 (.A(_108_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold77 (.A(\i_uart_tx.uart_tx_data[1] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold78 (.A(_014_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold79 (.A(\random_buffer_r[23] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold80 (.A(_044_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold81 (.A(\random_buffer_r[2] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold82 (.A(_023_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold83 (.A(\random_buffer_r[31] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold84 (.A(_052_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold85 (.A(\random_buffer_r[18] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold86 (.A(_039_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold87 (.A(\random_buffer_r[25] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold88 (.A(_046_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold89 (.A(\random_buffer_r[20] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold90 (.A(_041_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold91 (.A(\random_buffer_r[22] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold92 (.A(_043_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_uart_tx.uart_tx_data[0] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold94 (.A(_013_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold95 (.A(\random_buffer_r[21] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold96 (.A(_042_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold97 (.A(\random_buffer_r[15] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold98 (.A(_036_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold99 (.A(\random_buffer_r[30] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold100 (.A(_051_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold101 (.A(\random_buffer_r[7] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold102 (.A(_028_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_uart_tx.data_to_send[1] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold104 (.A(_155_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold105 (.A(_007_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_random.rnd_out[23] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold107 (.A(_086_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold108 (.A(\i_uart_tx.data_to_send[0] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_uart_tx.bit_counter[3] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold110 (.A(_232_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold111 (.A(_100_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold112 (.A(\i_uart_tx.bit_counter[1] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold113 (.A(_228_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold114 (.A(\random_buffer_r[26] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold115 (.A(_047_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_random.rnd_out[18] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold117 (.A(_081_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_random.rnd_out[2] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold119 (.A(\i_random.rnd_out[17] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_random.rnd_out[27] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold121 (.A(_090_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_random.rnd_out[21] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold123 (.A(_084_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold124 (.A(\i_random.rnd_out[19] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold125 (.A(_082_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold126 (.A(\i_uart_tx.fsm_state[0] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_random.rnd_out[26] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold128 (.A(\i_random.rnd_out[11] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold129 (.A(_073_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_uart_tx.uart_tx_data[2] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold131 (.A(_015_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold132 (.A(_001_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_random.rnd_out[22] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_random.rnd_out[24] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold135 (.A(_087_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold136 (.A(\i_random.rnd_out[9] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold137 (.A(_072_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_random.rnd_out[12] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold139 (.A(\i_random.rnd_out[16] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_random.rnd_out[8] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold141 (.A(\random_buffer_r[27] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold142 (.A(\i_random.rnd_out[29] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold143 (.A(_092_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold144 (.A(\i_random.rnd_out[4] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold145 (.A(\i_random.rnd_out[20] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold146 (.A(\i_uart_tx.cycle_counter[4] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold147 (.A(_243_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold148 (.A(\i_random.rnd_out[13] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_random.rnd_out[31] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold150 (.A(_093_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_random.first_bit ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold152 (.A(_053_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_random.rnd_out[7] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold154 (.A(\i_random.rnd_out[25] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_random.rnd_out[28] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold156 (.A(\i_uart_tx.uart_tx_data[4] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_uart_tx.data_to_send[6] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold158 (.A(_012_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold159 (.A(\i_random.rnd_out[14] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_random.rnd_out[15] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_uart_tx.data_to_send[4] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold162 (.A(_010_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold163 (.A(\i_uart_tx.uart_tx_en ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold164 (.A(\byte_counter_r[0] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold165 (.A(_094_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold166 (.A(\byte_counter_r[1] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold167 (.A(_095_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold168 (.A(\i_uart_tx.cycle_counter[2] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold169 (.A(_239_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_uart_tx.cycle_counter[6] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold171 (.A(_247_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold172 (.A(fsm_state_r),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_uart_tx.cycle_counter[3] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_uart_tx.bit_counter[2] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold175 (.A(_230_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_random.bit_count[1] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold177 (.A(\i_random.bit_count[4] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold178 (.A(\i_uart_tx.fsm_state[1] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold179 (.A(_147_),
    .X(net257));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_4 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_209 ();
 sg13g2_decap_8 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_251 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_265 ();
 sg13g2_decap_8 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_4 FILLER_9_168 ();
 sg13g2_fill_1 FILLER_9_172 ();
 sg13g2_fill_1 FILLER_9_182 ();
 sg13g2_fill_2 FILLER_9_192 ();
 sg13g2_decap_4 FILLER_9_204 ();
 sg13g2_fill_1 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_218 ();
 sg13g2_decap_8 FILLER_9_225 ();
 sg13g2_decap_8 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_239 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_decap_8 FILLER_9_253 ();
 sg13g2_decap_8 FILLER_9_260 ();
 sg13g2_decap_8 FILLER_9_267 ();
 sg13g2_decap_8 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_281 ();
 sg13g2_decap_8 FILLER_9_288 ();
 sg13g2_decap_8 FILLER_9_295 ();
 sg13g2_decap_8 FILLER_9_302 ();
 sg13g2_decap_8 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_316 ();
 sg13g2_decap_8 FILLER_9_323 ();
 sg13g2_decap_8 FILLER_9_330 ();
 sg13g2_decap_8 FILLER_9_337 ();
 sg13g2_decap_8 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_351 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_decap_8 FILLER_9_365 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_4 FILLER_10_105 ();
 sg13g2_fill_1 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_fill_2 FILLER_10_147 ();
 sg13g2_decap_4 FILLER_10_168 ();
 sg13g2_decap_4 FILLER_10_191 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_fill_2 FILLER_10_249 ();
 sg13g2_fill_1 FILLER_10_251 ();
 sg13g2_decap_4 FILLER_10_260 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_289 ();
 sg13g2_decap_8 FILLER_10_296 ();
 sg13g2_decap_8 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_4 FILLER_11_131 ();
 sg13g2_fill_2 FILLER_11_170 ();
 sg13g2_fill_1 FILLER_11_172 ();
 sg13g2_fill_2 FILLER_11_209 ();
 sg13g2_fill_1 FILLER_11_211 ();
 sg13g2_decap_4 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_fill_2 FILLER_12_98 ();
 sg13g2_fill_1 FILLER_12_100 ();
 sg13g2_fill_1 FILLER_12_127 ();
 sg13g2_decap_4 FILLER_12_164 ();
 sg13g2_fill_1 FILLER_12_168 ();
 sg13g2_fill_2 FILLER_12_178 ();
 sg13g2_decap_4 FILLER_12_216 ();
 sg13g2_fill_2 FILLER_12_220 ();
 sg13g2_decap_4 FILLER_12_284 ();
 sg13g2_fill_1 FILLER_12_288 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_4 FILLER_13_84 ();
 sg13g2_fill_1 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_151 ();
 sg13g2_fill_1 FILLER_13_158 ();
 sg13g2_fill_1 FILLER_13_195 ();
 sg13g2_decap_4 FILLER_13_205 ();
 sg13g2_fill_2 FILLER_13_218 ();
 sg13g2_fill_1 FILLER_13_220 ();
 sg13g2_fill_1 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_297 ();
 sg13g2_decap_8 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_decap_4 FILLER_14_120 ();
 sg13g2_decap_4 FILLER_14_134 ();
 sg13g2_fill_2 FILLER_14_138 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_1 FILLER_14_216 ();
 sg13g2_decap_8 FILLER_14_243 ();
 sg13g2_decap_4 FILLER_14_278 ();
 sg13g2_fill_2 FILLER_14_282 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_4 FILLER_15_84 ();
 sg13g2_fill_1 FILLER_15_88 ();
 sg13g2_fill_2 FILLER_15_99 ();
 sg13g2_fill_1 FILLER_15_101 ();
 sg13g2_fill_2 FILLER_15_137 ();
 sg13g2_fill_1 FILLER_15_139 ();
 sg13g2_decap_4 FILLER_15_169 ();
 sg13g2_decap_4 FILLER_15_208 ();
 sg13g2_fill_2 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_decap_8 FILLER_15_317 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_fill_1 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_4 FILLER_15_403 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_fill_2 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_72 ();
 sg13g2_fill_2 FILLER_16_108 ();
 sg13g2_decap_8 FILLER_16_164 ();
 sg13g2_fill_2 FILLER_16_189 ();
 sg13g2_fill_1 FILLER_16_191 ();
 sg13g2_decap_4 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_233 ();
 sg13g2_fill_2 FILLER_16_240 ();
 sg13g2_decap_4 FILLER_16_252 ();
 sg13g2_fill_2 FILLER_16_256 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_283 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_decap_4 FILLER_16_317 ();
 sg13g2_fill_2 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_fill_2 FILLER_17_63 ();
 sg13g2_fill_2 FILLER_17_167 ();
 sg13g2_fill_1 FILLER_17_178 ();
 sg13g2_fill_1 FILLER_17_188 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_fill_2 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_4 FILLER_18_56 ();
 sg13g2_fill_2 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_117 ();
 sg13g2_fill_1 FILLER_18_119 ();
 sg13g2_fill_2 FILLER_18_181 ();
 sg13g2_fill_1 FILLER_18_183 ();
 sg13g2_fill_1 FILLER_18_208 ();
 sg13g2_decap_8 FILLER_18_218 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_8 FILLER_18_232 ();
 sg13g2_decap_4 FILLER_18_239 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_4 FILLER_19_70 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_fill_1 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_130 ();
 sg13g2_fill_1 FILLER_19_137 ();
 sg13g2_fill_2 FILLER_19_147 ();
 sg13g2_fill_1 FILLER_19_149 ();
 sg13g2_decap_4 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_179 ();
 sg13g2_decap_4 FILLER_19_186 ();
 sg13g2_decap_4 FILLER_19_224 ();
 sg13g2_fill_2 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_265 ();
 sg13g2_fill_1 FILLER_19_272 ();
 sg13g2_fill_2 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_fill_2 FILLER_19_322 ();
 sg13g2_fill_1 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_330 ();
 sg13g2_fill_2 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_4 FILLER_20_84 ();
 sg13g2_fill_1 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_108 ();
 sg13g2_fill_1 FILLER_20_115 ();
 sg13g2_decap_8 FILLER_20_152 ();
 sg13g2_decap_8 FILLER_20_159 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_decap_8 FILLER_20_177 ();
 sg13g2_fill_2 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_226 ();
 sg13g2_decap_8 FILLER_20_233 ();
 sg13g2_fill_2 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_242 ();
 sg13g2_decap_4 FILLER_20_249 ();
 sg13g2_fill_2 FILLER_20_253 ();
 sg13g2_decap_8 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_267 ();
 sg13g2_fill_1 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_323 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_113 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_decap_8 FILLER_21_226 ();
 sg13g2_decap_8 FILLER_21_233 ();
 sg13g2_decap_8 FILLER_21_240 ();
 sg13g2_decap_8 FILLER_21_247 ();
 sg13g2_fill_1 FILLER_21_259 ();
 sg13g2_fill_2 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_376 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_4 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_81 ();
 sg13g2_decap_4 FILLER_22_108 ();
 sg13g2_fill_1 FILLER_22_112 ();
 sg13g2_fill_2 FILLER_22_173 ();
 sg13g2_decap_4 FILLER_22_212 ();
 sg13g2_fill_1 FILLER_22_216 ();
 sg13g2_decap_8 FILLER_22_220 ();
 sg13g2_decap_8 FILLER_22_227 ();
 sg13g2_fill_2 FILLER_22_234 ();
 sg13g2_fill_1 FILLER_22_236 ();
 sg13g2_decap_8 FILLER_22_240 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_249 ();
 sg13g2_fill_1 FILLER_22_311 ();
 sg13g2_fill_1 FILLER_22_325 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_4 FILLER_23_77 ();
 sg13g2_fill_1 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_127 ();
 sg13g2_fill_2 FILLER_23_142 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_2 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_fill_1 FILLER_23_254 ();
 sg13g2_fill_2 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_316 ();
 sg13g2_fill_1 FILLER_23_386 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_140 ();
 sg13g2_fill_2 FILLER_24_163 ();
 sg13g2_fill_1 FILLER_24_174 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_decap_4 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_314 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_fill_2 FILLER_24_380 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_fill_2 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_114 ();
 sg13g2_decap_4 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_decap_4 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_265 ();
 sg13g2_decap_4 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_335 ();
 sg13g2_fill_2 FILLER_25_361 ();
 sg13g2_fill_1 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_4 FILLER_26_91 ();
 sg13g2_fill_2 FILLER_26_95 ();
 sg13g2_decap_4 FILLER_26_123 ();
 sg13g2_fill_2 FILLER_26_127 ();
 sg13g2_fill_2 FILLER_26_181 ();
 sg13g2_fill_1 FILLER_26_183 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_fill_2 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_290 ();
 sg13g2_fill_1 FILLER_26_292 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_fill_2 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_fill_2 FILLER_26_366 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_4 FILLER_27_105 ();
 sg13g2_fill_1 FILLER_27_109 ();
 sg13g2_decap_4 FILLER_27_134 ();
 sg13g2_fill_1 FILLER_27_138 ();
 sg13g2_fill_2 FILLER_27_149 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_decap_4 FILLER_27_299 ();
 sg13g2_fill_2 FILLER_27_361 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_fill_2 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_121 ();
 sg13g2_decap_4 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_134 ();
 sg13g2_decap_8 FILLER_28_144 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_decap_8 FILLER_28_170 ();
 sg13g2_decap_8 FILLER_28_177 ();
 sg13g2_decap_8 FILLER_28_184 ();
 sg13g2_decap_4 FILLER_28_191 ();
 sg13g2_fill_2 FILLER_28_195 ();
 sg13g2_fill_2 FILLER_28_223 ();
 sg13g2_fill_2 FILLER_28_229 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_291 ();
 sg13g2_decap_4 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_312 ();
 sg13g2_fill_2 FILLER_28_322 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_decap_8 FILLER_28_333 ();
 sg13g2_decap_4 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_344 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_152 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_decap_8 FILLER_29_177 ();
 sg13g2_decap_4 FILLER_29_184 ();
 sg13g2_fill_2 FILLER_29_188 ();
 sg13g2_fill_2 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_219 ();
 sg13g2_fill_2 FILLER_29_226 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_234 ();
 sg13g2_decap_8 FILLER_29_239 ();
 sg13g2_decap_8 FILLER_29_246 ();
 sg13g2_decap_4 FILLER_29_253 ();
 sg13g2_decap_8 FILLER_29_282 ();
 sg13g2_decap_8 FILLER_29_289 ();
 sg13g2_decap_8 FILLER_29_296 ();
 sg13g2_decap_8 FILLER_29_303 ();
 sg13g2_fill_2 FILLER_29_310 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_8 FILLER_29_331 ();
 sg13g2_decap_8 FILLER_29_338 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_144 ();
 sg13g2_decap_8 FILLER_30_159 ();
 sg13g2_fill_2 FILLER_30_166 ();
 sg13g2_fill_1 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_decap_8 FILLER_30_229 ();
 sg13g2_decap_8 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_249 ();
 sg13g2_decap_8 FILLER_30_290 ();
 sg13g2_decap_8 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_304 ();
 sg13g2_fill_2 FILLER_30_324 ();
 sg13g2_fill_1 FILLER_30_326 ();
 sg13g2_fill_1 FILLER_30_332 ();
 sg13g2_fill_2 FILLER_30_338 ();
 sg13g2_decap_4 FILLER_30_344 ();
 sg13g2_fill_2 FILLER_30_365 ();
 sg13g2_fill_2 FILLER_30_376 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_4 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_decap_4 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_158 ();
 sg13g2_fill_2 FILLER_31_185 ();
 sg13g2_fill_1 FILLER_31_187 ();
 sg13g2_decap_4 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_299 ();
 sg13g2_fill_2 FILLER_31_341 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_fill_2 FILLER_32_126 ();
 sg13g2_fill_1 FILLER_32_128 ();
 sg13g2_decap_4 FILLER_32_138 ();
 sg13g2_decap_4 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_336 ();
 sg13g2_fill_2 FILLER_32_362 ();
 sg13g2_fill_2 FILLER_32_372 ();
 sg13g2_fill_1 FILLER_32_374 ();
 sg13g2_fill_2 FILLER_32_384 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_4 FILLER_33_126 ();
 sg13g2_fill_2 FILLER_33_130 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_fill_1 FILLER_33_161 ();
 sg13g2_decap_4 FILLER_33_171 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_195 ();
 sg13g2_decap_8 FILLER_33_202 ();
 sg13g2_fill_1 FILLER_33_209 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_decap_8 FILLER_33_227 ();
 sg13g2_decap_8 FILLER_33_234 ();
 sg13g2_decap_8 FILLER_33_241 ();
 sg13g2_fill_2 FILLER_33_271 ();
 sg13g2_fill_1 FILLER_33_282 ();
 sg13g2_fill_2 FILLER_33_292 ();
 sg13g2_fill_2 FILLER_33_303 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_178 ();
 sg13g2_decap_8 FILLER_34_185 ();
 sg13g2_decap_8 FILLER_34_192 ();
 sg13g2_decap_4 FILLER_34_199 ();
 sg13g2_decap_8 FILLER_34_207 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_4 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_fill_2 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_289 ();
 sg13g2_fill_2 FILLER_34_356 ();
 sg13g2_decap_4 FILLER_34_392 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_4 FILLER_35_189 ();
 sg13g2_decap_4 FILLER_35_249 ();
 sg13g2_decap_8 FILLER_35_261 ();
 sg13g2_decap_8 FILLER_35_268 ();
 sg13g2_decap_4 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_365 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_fill_1 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_208 ();
 sg13g2_decap_4 FILLER_36_215 ();
 sg13g2_fill_2 FILLER_36_271 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_4 FILLER_37_224 ();
 sg13g2_fill_1 FILLER_37_228 ();
 sg13g2_decap_8 FILLER_37_265 ();
 sg13g2_decap_4 FILLER_37_272 ();
 sg13g2_fill_2 FILLER_37_276 ();
 sg13g2_fill_2 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_219 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_decap_8 FILLER_38_233 ();
 sg13g2_fill_2 FILLER_38_240 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_255 ();
 sg13g2_decap_8 FILLER_38_262 ();
 sg13g2_decap_4 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_273 ();
 sg13g2_fill_2 FILLER_38_300 ();
 sg13g2_fill_1 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_347 ();
 sg13g2_fill_2 FILLER_38_354 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[4] = net18;
 assign uo_out[5] = net19;
 assign uo_out[6] = net20;
 assign uo_out[7] = net21;
endmodule
