module tt_um_wokwi_434917200607612929 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire params_ready;
 wire spike_out;
 wire \system_inst.leak_cycles_1[0] ;
 wire \system_inst.leak_cycles_1[1] ;
 wire \system_inst.leak_cycles_1[2] ;
 wire \system_inst.leak_cycles_1[3] ;
 wire \system_inst.leak_cycles_2[0] ;
 wire \system_inst.leak_cycles_2[1] ;
 wire \system_inst.leak_cycles_2[2] ;
 wire \system_inst.leak_cycles_2[3] ;
 wire \system_inst.leak_rate_1[0] ;
 wire \system_inst.leak_rate_1[1] ;
 wire \system_inst.leak_rate_1[2] ;
 wire \system_inst.leak_rate_1[3] ;
 wire \system_inst.leak_rate_1[4] ;
 wire \system_inst.leak_rate_1[5] ;
 wire \system_inst.leak_rate_1[6] ;
 wire \system_inst.leak_rate_1[7] ;
 wire \system_inst.leak_rate_2[0] ;
 wire \system_inst.leak_rate_2[1] ;
 wire \system_inst.leak_rate_2[2] ;
 wire \system_inst.leak_rate_2[3] ;
 wire \system_inst.leak_rate_2[4] ;
 wire \system_inst.leak_rate_2[5] ;
 wire \system_inst.leak_rate_2[6] ;
 wire \system_inst.leak_rate_2[7] ;
 wire \system_inst.loader.bit_count[0] ;
 wire \system_inst.loader.bit_count[1] ;
 wire \system_inst.loader.bit_count[2] ;
 wire \system_inst.loader.current_state[0] ;
 wire \system_inst.loader.current_state[1] ;
 wire \system_inst.loader.current_state[2] ;
 wire \system_inst.loader.current_state[3] ;
 wire \system_inst.loader.current_state[4] ;
 wire \system_inst.loader.current_state[5] ;
 wire \system_inst.loader.current_state[6] ;
 wire \system_inst.loader.shift_reg[0] ;
 wire \system_inst.loader.shift_reg[1] ;
 wire \system_inst.loader.shift_reg[2] ;
 wire \system_inst.loader.shift_reg[3] ;
 wire \system_inst.loader.shift_reg[4] ;
 wire \system_inst.loader.shift_reg[5] ;
 wire \system_inst.loader.shift_reg[6] ;
 wire \system_inst.loader.threshold[0] ;
 wire \system_inst.loader.threshold[1] ;
 wire \system_inst.loader.threshold[2] ;
 wire \system_inst.loader.threshold[3] ;
 wire \system_inst.loader.threshold[4] ;
 wire \system_inst.loader.threshold[5] ;
 wire \system_inst.loader.threshold[6] ;
 wire \system_inst.loader.threshold[7] ;
 wire \system_inst.loader.weight_a[0] ;
 wire \system_inst.loader.weight_a[1] ;
 wire \system_inst.loader.weight_a[2] ;
 wire \system_inst.neuron.leak_counter_1[0] ;
 wire \system_inst.neuron.leak_counter_1[1] ;
 wire \system_inst.neuron.leak_counter_1[2] ;
 wire \system_inst.neuron.leak_counter_1[3] ;
 wire \system_inst.neuron.leak_counter_2[0] ;
 wire \system_inst.neuron.leak_counter_2[1] ;
 wire \system_inst.neuron.leak_counter_2[2] ;
 wire \system_inst.neuron.leak_counter_2[3] ;
 wire \system_inst.neuron.refr_cnt[0] ;
 wire \system_inst.neuron.refr_cnt[1] ;
 wire \system_inst.neuron.refr_cnt[2] ;
 wire \system_inst.neuron.refr_cnt[3] ;
 wire \system_inst.neuron.v_mem[0] ;
 wire \system_inst.neuron.v_mem[1] ;
 wire \system_inst.neuron.v_mem[2] ;
 wire \system_inst.neuron.v_mem[3] ;
 wire \system_inst.neuron.v_mem[4] ;
 wire \system_inst.neuron.v_mem[5] ;
 wire \system_inst.neuron.v_mem[6] ;
 wire \system_inst.neuron.v_mem[7] ;
 wire \system_inst.neuron.v_mem[8] ;
 wire clknet_0_clk;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;

 sg13g2_inv_1 _0786_ (.Y(_0099_),
    .A(net167));
 sg13g2_inv_2 _0787_ (.Y(_0100_),
    .A(net180));
 sg13g2_inv_2 _0788_ (.Y(_0101_),
    .A(net182));
 sg13g2_inv_1 _0789_ (.Y(_0102_),
    .A(net217));
 sg13g2_inv_2 _0790_ (.Y(_0103_),
    .A(net165));
 sg13g2_inv_2 _0791_ (.Y(_0104_),
    .A(net223));
 sg13g2_inv_2 _0792_ (.Y(_0105_),
    .A(net221));
 sg13g2_inv_1 _0793_ (.Y(_0106_),
    .A(\system_inst.leak_cycles_2[3] ));
 sg13g2_inv_1 _0794_ (.Y(_0107_),
    .A(net160));
 sg13g2_inv_2 _0795_ (.Y(_0108_),
    .A(net4));
 sg13g2_inv_1 _0796_ (.Y(_0109_),
    .A(net158));
 sg13g2_inv_1 _0797_ (.Y(_0110_),
    .A(\system_inst.loader.threshold[7] ));
 sg13g2_inv_1 _0798_ (.Y(_0111_),
    .A(net237));
 sg13g2_inv_1 _0799_ (.Y(_0112_),
    .A(net227));
 sg13g2_inv_1 _0800_ (.Y(_0113_),
    .A(net240));
 sg13g2_inv_1 _0801_ (.Y(_0114_),
    .A(net170));
 sg13g2_inv_1 _0802_ (.Y(_0115_),
    .A(net235));
 sg13g2_inv_1 _0803_ (.Y(_0116_),
    .A(\system_inst.neuron.leak_counter_2[2] ));
 sg13g2_inv_1 _0804_ (.Y(_0117_),
    .A(\system_inst.neuron.leak_counter_2[1] ));
 sg13g2_inv_1 _0805_ (.Y(_0118_),
    .A(net5));
 sg13g2_inv_1 _0806_ (.Y(_0119_),
    .A(_0026_));
 sg13g2_inv_1 _0807_ (.Y(_0120_),
    .A(_0027_));
 sg13g2_inv_1 _0808_ (.Y(_0121_),
    .A(_0028_));
 sg13g2_inv_2 _0809_ (.Y(_0122_),
    .A(net140));
 sg13g2_inv_1 _0810_ (.Y(_0123_),
    .A(\system_inst.loader.current_state[0] ));
 sg13g2_inv_1 _0811_ (.Y(_0124_),
    .A(net148));
 sg13g2_and2_1 _0812_ (.A(net1),
    .B(net3),
    .X(_0125_));
 sg13g2_nand2_1 _0813_ (.Y(_0126_),
    .A(net140),
    .B(net130));
 sg13g2_nand2b_1 _0814_ (.Y(_0127_),
    .B(net140),
    .A_N(net1));
 sg13g2_nor2_1 _0815_ (.A(net153),
    .B(_0127_),
    .Y(_0128_));
 sg13g2_a21oi_1 _0816_ (.A1(net138),
    .A2(net130),
    .Y(_0000_),
    .B1(_0128_));
 sg13g2_nand2_2 _0817_ (.Y(_0129_),
    .A(net174),
    .B(net154));
 sg13g2_nor2_2 _0818_ (.A(_0029_),
    .B(_0129_),
    .Y(_0130_));
 sg13g2_o21ai_1 _0819_ (.B1(_0127_),
    .Y(_0131_),
    .A1(_0126_),
    .A2(net125));
 sg13g2_nand3_1 _0820_ (.B(net130),
    .C(net125),
    .A(net103),
    .Y(_0132_));
 sg13g2_inv_1 _0821_ (.Y(_0133_),
    .A(_0132_));
 sg13g2_a22oi_1 _0822_ (.Y(_0134_),
    .B1(_0133_),
    .B2(net140),
    .A2(_0131_),
    .A1(net147));
 sg13g2_inv_1 _0823_ (.Y(_0002_),
    .A(_0134_));
 sg13g2_and3_1 _0824_ (.X(_0135_),
    .A(\system_inst.loader.current_state[5] ),
    .B(net130),
    .C(net125));
 sg13g2_a22oi_1 _0825_ (.Y(_0136_),
    .B1(_0135_),
    .B2(net138),
    .A2(_0131_),
    .A1(net148));
 sg13g2_inv_1 _0826_ (.Y(_0003_),
    .A(net149));
 sg13g2_nand2_1 _0827_ (.Y(_0137_),
    .A(net103),
    .B(_0131_));
 sg13g2_o21ai_1 _0828_ (.B1(_0137_),
    .Y(_0004_),
    .A1(_0123_),
    .A2(_0126_));
 sg13g2_and3_1 _0829_ (.X(_0138_),
    .A(\system_inst.loader.current_state[1] ),
    .B(_0125_),
    .C(_0130_));
 sg13g2_nand3_1 _0830_ (.B(net130),
    .C(_0130_),
    .A(net198),
    .Y(_0139_));
 sg13g2_a22oi_1 _0831_ (.Y(_0140_),
    .B1(net123),
    .B2(net138),
    .A2(_0131_),
    .A1(net177));
 sg13g2_inv_1 _0832_ (.Y(_0005_),
    .A(_0140_));
 sg13g2_and3_1 _0833_ (.X(_0141_),
    .A(net147),
    .B(net130),
    .C(net125));
 sg13g2_a22oi_1 _0834_ (.Y(_0142_),
    .B1(net121),
    .B2(net137),
    .A2(_0131_),
    .A1(net157));
 sg13g2_inv_1 _0835_ (.Y(_0006_),
    .A(_0142_));
 sg13g2_and3_1 _0836_ (.X(_0143_),
    .A(\system_inst.loader.current_state[6] ),
    .B(net130),
    .C(net125));
 sg13g2_a22oi_1 _0837_ (.Y(_0144_),
    .B1(net118),
    .B2(net137),
    .A2(_0131_),
    .A1(net198));
 sg13g2_inv_1 _0838_ (.Y(_0001_),
    .A(_0144_));
 sg13g2_nor2b_1 _0839_ (.A(net129),
    .B_N(\system_inst.neuron.v_mem[0] ),
    .Y(uo_out[1]));
 sg13g2_nor2b_1 _0840_ (.A(net129),
    .B_N(\system_inst.neuron.v_mem[1] ),
    .Y(uo_out[2]));
 sg13g2_nor2b_1 _0841_ (.A(net129),
    .B_N(\system_inst.neuron.v_mem[2] ),
    .Y(uo_out[3]));
 sg13g2_nor2b_1 _0842_ (.A(net129),
    .B_N(\system_inst.neuron.v_mem[3] ),
    .Y(uo_out[4]));
 sg13g2_nor2b_1 _0843_ (.A(net129),
    .B_N(\system_inst.neuron.v_mem[4] ),
    .Y(uo_out[5]));
 sg13g2_nor2b_1 _0844_ (.A(net129),
    .B_N(\system_inst.neuron.v_mem[5] ),
    .Y(uo_out[6]));
 sg13g2_nor2b_1 _0845_ (.A(net129),
    .B_N(\system_inst.neuron.v_mem[6] ),
    .Y(uo_out[7]));
 sg13g2_and3_1 _0846_ (.X(_0145_),
    .A(net127),
    .B(\system_inst.neuron.v_mem[4] ),
    .C(net7));
 sg13g2_nand3_1 _0847_ (.B(\system_inst.neuron.v_mem[4] ),
    .C(net7),
    .A(net128),
    .Y(_0146_));
 sg13g2_nand2_1 _0848_ (.Y(_0147_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net8));
 sg13g2_a21oi_1 _0849_ (.A1(net128),
    .A2(net7),
    .Y(_0148_),
    .B1(\system_inst.neuron.v_mem[4] ));
 sg13g2_nor2_1 _0850_ (.A(_0145_),
    .B(_0148_),
    .Y(_0149_));
 sg13g2_o21ai_1 _0851_ (.B1(_0146_),
    .Y(_0150_),
    .A1(_0147_),
    .A2(_0148_));
 sg13g2_nand2_1 _0852_ (.Y(_0151_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net9));
 sg13g2_nand3_1 _0853_ (.B(\system_inst.neuron.v_mem[5] ),
    .C(net8),
    .A(net127),
    .Y(_0152_));
 sg13g2_a21o_1 _0854_ (.A2(net8),
    .A1(net127),
    .B1(\system_inst.neuron.v_mem[5] ),
    .X(_0153_));
 sg13g2_nand2_1 _0855_ (.Y(_0154_),
    .A(_0152_),
    .B(_0153_));
 sg13g2_xor2_1 _0856_ (.B(_0154_),
    .A(_0151_),
    .X(_0155_));
 sg13g2_nand2_1 _0857_ (.Y(_0156_),
    .A(_0150_),
    .B(_0155_));
 sg13g2_nand2_1 _0858_ (.Y(_0157_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net10));
 sg13g2_xnor2_1 _0859_ (.Y(_0158_),
    .A(_0150_),
    .B(_0155_));
 sg13g2_or2_1 _0860_ (.X(_0159_),
    .B(_0158_),
    .A(_0157_));
 sg13g2_o21ai_1 _0861_ (.B1(_0152_),
    .Y(_0160_),
    .A1(_0151_),
    .A2(_0154_));
 sg13g2_nand2_1 _0862_ (.Y(_0161_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net10));
 sg13g2_nand3_1 _0863_ (.B(\system_inst.neuron.v_mem[6] ),
    .C(net9),
    .A(net127),
    .Y(_0162_));
 sg13g2_a21o_1 _0864_ (.A2(net9),
    .A1(net127),
    .B1(\system_inst.neuron.v_mem[6] ),
    .X(_0163_));
 sg13g2_nand2_1 _0865_ (.Y(_0164_),
    .A(_0162_),
    .B(_0163_));
 sg13g2_xor2_1 _0866_ (.B(_0164_),
    .A(_0161_),
    .X(_0165_));
 sg13g2_nand2_1 _0867_ (.Y(_0166_),
    .A(_0160_),
    .B(_0165_));
 sg13g2_xnor2_1 _0868_ (.Y(_0167_),
    .A(_0160_),
    .B(_0165_));
 sg13g2_a21oi_1 _0869_ (.A1(_0156_),
    .A2(_0159_),
    .Y(_0168_),
    .B1(_0167_));
 sg13g2_nand3_1 _0870_ (.B(_0159_),
    .C(_0167_),
    .A(_0156_),
    .Y(_0169_));
 sg13g2_nand2b_1 _0871_ (.Y(_0170_),
    .B(_0169_),
    .A_N(_0168_));
 sg13g2_and3_1 _0872_ (.X(_0171_),
    .A(net128),
    .B(\system_inst.neuron.v_mem[3] ),
    .C(net6));
 sg13g2_nand3_1 _0873_ (.B(\system_inst.neuron.v_mem[3] ),
    .C(net6),
    .A(net127),
    .Y(_0172_));
 sg13g2_nand2_1 _0874_ (.Y(_0173_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net7));
 sg13g2_a21oi_1 _0875_ (.A1(net127),
    .A2(net6),
    .Y(_0174_),
    .B1(\system_inst.neuron.v_mem[3] ));
 sg13g2_nor2_1 _0876_ (.A(_0171_),
    .B(_0174_),
    .Y(_0175_));
 sg13g2_o21ai_1 _0877_ (.B1(_0172_),
    .Y(_0176_),
    .A1(_0173_),
    .A2(_0174_));
 sg13g2_xnor2_1 _0878_ (.Y(_0177_),
    .A(_0147_),
    .B(_0149_));
 sg13g2_nand2_1 _0879_ (.Y(_0178_),
    .A(_0176_),
    .B(_0177_));
 sg13g2_nand2_1 _0880_ (.Y(_0179_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net9));
 sg13g2_xnor2_1 _0881_ (.Y(_0180_),
    .A(_0176_),
    .B(_0177_));
 sg13g2_o21ai_1 _0882_ (.B1(_0178_),
    .Y(_0181_),
    .A1(_0179_),
    .A2(_0180_));
 sg13g2_xor2_1 _0883_ (.B(_0158_),
    .A(_0157_),
    .X(_0182_));
 sg13g2_nor2_1 _0884_ (.A(_0181_),
    .B(_0182_),
    .Y(_0183_));
 sg13g2_and3_1 _0885_ (.X(_0184_),
    .A(net128),
    .B(\system_inst.neuron.v_mem[2] ),
    .C(net5));
 sg13g2_nand2_1 _0886_ (.Y(_0185_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net6));
 sg13g2_a21oi_1 _0887_ (.A1(net128),
    .A2(net5),
    .Y(_0186_),
    .B1(\system_inst.neuron.v_mem[2] ));
 sg13g2_or3_1 _0888_ (.A(_0184_),
    .B(_0185_),
    .C(_0186_),
    .X(_0187_));
 sg13g2_nand2b_1 _0889_ (.Y(_0188_),
    .B(_0187_),
    .A_N(_0184_));
 sg13g2_xnor2_1 _0890_ (.Y(_0189_),
    .A(_0173_),
    .B(_0175_));
 sg13g2_nand2_1 _0891_ (.Y(_0190_),
    .A(_0188_),
    .B(_0189_));
 sg13g2_nand2_1 _0892_ (.Y(_0191_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net8));
 sg13g2_xnor2_1 _0893_ (.Y(_0192_),
    .A(_0188_),
    .B(_0189_));
 sg13g2_o21ai_1 _0894_ (.B1(_0190_),
    .Y(_0193_),
    .A1(_0191_),
    .A2(_0192_));
 sg13g2_xor2_1 _0895_ (.B(_0180_),
    .A(_0179_),
    .X(_0194_));
 sg13g2_nand2_1 _0896_ (.Y(_0195_),
    .A(_0193_),
    .B(_0194_));
 sg13g2_xor2_1 _0897_ (.B(_0194_),
    .A(_0193_),
    .X(_0196_));
 sg13g2_and3_1 _0898_ (.X(_0197_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(\system_inst.neuron.v_mem[1] ),
    .C(net5));
 sg13g2_o21ai_1 _0899_ (.B1(_0185_),
    .Y(_0198_),
    .A1(_0184_),
    .A2(_0186_));
 sg13g2_and3_1 _0900_ (.X(_0199_),
    .A(_0187_),
    .B(_0197_),
    .C(_0198_));
 sg13g2_nand2_1 _0901_ (.Y(_0200_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net7));
 sg13g2_a21oi_1 _0902_ (.A1(_0187_),
    .A2(_0198_),
    .Y(_0201_),
    .B1(_0197_));
 sg13g2_or3_1 _0903_ (.A(_0199_),
    .B(_0200_),
    .C(_0201_),
    .X(_0202_));
 sg13g2_nand2b_2 _0904_ (.Y(_0203_),
    .B(_0202_),
    .A_N(_0199_));
 sg13g2_xor2_1 _0905_ (.B(_0192_),
    .A(_0191_),
    .X(_0204_));
 sg13g2_nor2_1 _0906_ (.A(_0203_),
    .B(_0204_),
    .Y(_0205_));
 sg13g2_or2_1 _0907_ (.X(_0206_),
    .B(_0204_),
    .A(_0203_));
 sg13g2_a21oi_1 _0908_ (.A1(\system_inst.loader.weight_a[1] ),
    .A2(net5),
    .Y(_0207_),
    .B1(\system_inst.neuron.v_mem[1] ));
 sg13g2_nand2_1 _0909_ (.Y(_0208_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net6));
 sg13g2_nor3_1 _0910_ (.A(_0197_),
    .B(_0207_),
    .C(_0208_),
    .Y(_0209_));
 sg13g2_o21ai_1 _0911_ (.B1(_0200_),
    .Y(_0210_),
    .A1(_0199_),
    .A2(_0201_));
 sg13g2_and3_1 _0912_ (.X(_0211_),
    .A(_0202_),
    .B(_0209_),
    .C(_0210_));
 sg13g2_nand3b_1 _0913_ (.B(net5),
    .C(\system_inst.loader.weight_a[0] ),
    .Y(_0212_),
    .A_N(_0008_));
 sg13g2_o21ai_1 _0914_ (.B1(_0208_),
    .Y(_0213_),
    .A1(_0197_),
    .A2(_0207_));
 sg13g2_nor2b_1 _0915_ (.A(_0209_),
    .B_N(_0213_),
    .Y(_0214_));
 sg13g2_nor2b_1 _0916_ (.A(_0212_),
    .B_N(_0214_),
    .Y(_0215_));
 sg13g2_a21o_1 _0917_ (.A2(_0210_),
    .A1(_0202_),
    .B1(_0209_),
    .X(_0216_));
 sg13g2_nand2b_1 _0918_ (.Y(_0217_),
    .B(_0216_),
    .A_N(_0211_));
 sg13g2_a221oi_1 _0919_ (.B2(_0216_),
    .C1(_0211_),
    .B1(_0215_),
    .A1(_0203_),
    .Y(_0218_),
    .A2(_0204_));
 sg13g2_xnor2_1 _0920_ (.Y(_0219_),
    .A(_0203_),
    .B(_0204_));
 sg13g2_nor2_1 _0921_ (.A(_0205_),
    .B(_0218_),
    .Y(_0220_));
 sg13g2_nand3b_1 _0922_ (.B(_0196_),
    .C(_0206_),
    .Y(_0221_),
    .A_N(_0218_));
 sg13g2_nand2_1 _0923_ (.Y(_0222_),
    .A(_0181_),
    .B(_0182_));
 sg13g2_and2_1 _0924_ (.A(_0195_),
    .B(_0222_),
    .X(_0223_));
 sg13g2_a21oi_1 _0925_ (.A1(_0221_),
    .A2(_0223_),
    .Y(_0224_),
    .B1(_0183_));
 sg13g2_a21oi_1 _0926_ (.A1(_0169_),
    .A2(_0224_),
    .Y(_0225_),
    .B1(_0168_));
 sg13g2_o21ai_1 _0927_ (.B1(_0162_),
    .Y(_0226_),
    .A1(_0161_),
    .A2(_0164_));
 sg13g2_nand2_1 _0928_ (.Y(_0227_),
    .A(net127),
    .B(net10));
 sg13g2_nor2_1 _0929_ (.A(_0007_),
    .B(_0227_),
    .Y(_0228_));
 sg13g2_nand2_1 _0930_ (.Y(_0229_),
    .A(_0007_),
    .B(_0227_));
 sg13g2_nor2b_1 _0931_ (.A(_0228_),
    .B_N(_0229_),
    .Y(_0230_));
 sg13g2_xnor2_1 _0932_ (.Y(_0231_),
    .A(_0226_),
    .B(_0230_));
 sg13g2_or2_1 _0933_ (.X(_0232_),
    .B(_0231_),
    .A(_0166_));
 sg13g2_xnor2_1 _0934_ (.Y(_0233_),
    .A(_0166_),
    .B(_0231_));
 sg13g2_xor2_1 _0935_ (.B(_0233_),
    .A(_0225_),
    .X(_0234_));
 sg13g2_or3_2 _0936_ (.A(\system_inst.leak_rate_1[2] ),
    .B(\system_inst.leak_rate_1[1] ),
    .C(\system_inst.leak_rate_1[0] ),
    .X(_0235_));
 sg13g2_nor2_1 _0937_ (.A(\system_inst.leak_rate_1[3] ),
    .B(_0235_),
    .Y(_0236_));
 sg13g2_nor3_1 _0938_ (.A(\system_inst.leak_rate_1[4] ),
    .B(\system_inst.leak_rate_1[3] ),
    .C(_0235_),
    .Y(_0237_));
 sg13g2_nor2b_1 _0939_ (.A(\system_inst.leak_rate_1[5] ),
    .B_N(_0237_),
    .Y(_0238_));
 sg13g2_nand2b_1 _0940_ (.Y(_0239_),
    .B(_0238_),
    .A_N(\system_inst.leak_rate_1[6] ));
 sg13g2_nand2_1 _0941_ (.Y(_0240_),
    .A(\system_inst.leak_rate_1[7] ),
    .B(_0239_));
 sg13g2_xnor2_1 _0942_ (.Y(_0241_),
    .A(_0170_),
    .B(_0224_));
 sg13g2_xnor2_1 _0943_ (.Y(_0242_),
    .A(_0009_),
    .B(_0241_));
 sg13g2_nand2b_1 _0944_ (.Y(_0243_),
    .B(_0222_),
    .A_N(_0183_));
 sg13g2_nand3_1 _0945_ (.B(_0221_),
    .C(_0243_),
    .A(_0195_),
    .Y(_0244_));
 sg13g2_a21o_1 _0946_ (.A2(_0221_),
    .A1(_0195_),
    .B1(_0243_),
    .X(_0245_));
 sg13g2_and2_2 _0947_ (.A(_0244_),
    .B(_0245_),
    .X(_0246_));
 sg13g2_a21oi_1 _0948_ (.A1(_0244_),
    .A2(_0245_),
    .Y(_0247_),
    .B1(_0010_));
 sg13g2_xor2_1 _0949_ (.B(_0220_),
    .A(_0196_),
    .X(_0248_));
 sg13g2_nor2_1 _0950_ (.A(_0011_),
    .B(_0248_),
    .Y(_0249_));
 sg13g2_nand3_1 _0951_ (.B(_0244_),
    .C(_0245_),
    .A(_0010_),
    .Y(_0250_));
 sg13g2_xor2_1 _0952_ (.B(_0248_),
    .A(_0011_),
    .X(_0251_));
 sg13g2_nand3b_1 _0953_ (.B(_0250_),
    .C(_0251_),
    .Y(_0252_),
    .A_N(_0247_));
 sg13g2_nor3_1 _0954_ (.A(_0234_),
    .B(_0242_),
    .C(_0252_),
    .Y(_0253_));
 sg13g2_a21oi_1 _0955_ (.A1(_0215_),
    .A2(_0216_),
    .Y(_0254_),
    .B1(_0211_));
 sg13g2_xnor2_1 _0956_ (.Y(_0255_),
    .A(_0219_),
    .B(_0254_));
 sg13g2_inv_1 _0957_ (.Y(_0256_),
    .A(_0255_));
 sg13g2_xor2_1 _0958_ (.B(_0217_),
    .A(_0215_),
    .X(_0257_));
 sg13g2_inv_1 _0959_ (.Y(_0258_),
    .A(_0257_));
 sg13g2_xor2_1 _0960_ (.B(_0257_),
    .A(_0012_),
    .X(_0259_));
 sg13g2_xnor2_1 _0961_ (.Y(_0260_),
    .A(\system_inst.loader.threshold[4] ),
    .B(_0255_));
 sg13g2_nor2_1 _0962_ (.A(_0259_),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_xnor2_1 _0963_ (.Y(_0262_),
    .A(_0212_),
    .B(_0214_));
 sg13g2_inv_1 _0964_ (.Y(_0263_),
    .A(_0262_));
 sg13g2_nand2_1 _0965_ (.Y(_0264_),
    .A(\system_inst.loader.threshold[2] ),
    .B(_0263_));
 sg13g2_o21ai_1 _0966_ (.B1(_0008_),
    .Y(_0265_),
    .A1(_0115_),
    .A2(_0118_));
 sg13g2_nand2_2 _0967_ (.Y(_0266_),
    .A(_0212_),
    .B(_0265_));
 sg13g2_nor2_1 _0968_ (.A(\system_inst.loader.threshold[1] ),
    .B(_0266_),
    .Y(_0267_));
 sg13g2_xnor2_1 _0969_ (.Y(_0268_),
    .A(_0013_),
    .B(_0262_));
 sg13g2_o21ai_1 _0970_ (.B1(_0264_),
    .Y(_0269_),
    .A1(_0267_),
    .A2(_0268_));
 sg13g2_a22oi_1 _0971_ (.Y(_0270_),
    .B1(_0257_),
    .B2(\system_inst.loader.threshold[3] ),
    .A2(_0255_),
    .A1(\system_inst.loader.threshold[4] ));
 sg13g2_a21oi_1 _0972_ (.A1(_0111_),
    .A2(_0256_),
    .Y(_0271_),
    .B1(_0270_));
 sg13g2_a21oi_1 _0973_ (.A1(_0261_),
    .A2(_0269_),
    .Y(_0272_),
    .B1(_0271_));
 sg13g2_nor4_2 _0974_ (.A(_0234_),
    .B(_0242_),
    .C(_0252_),
    .Y(_0273_),
    .D(_0272_));
 sg13g2_a21oi_1 _0975_ (.A1(_0249_),
    .A2(_0250_),
    .Y(_0274_),
    .B1(_0247_));
 sg13g2_nor3_1 _0976_ (.A(_0234_),
    .B(_0242_),
    .C(_0274_),
    .Y(_0275_));
 sg13g2_nor3_1 _0977_ (.A(_0110_),
    .B(_0234_),
    .C(_0241_),
    .Y(_0276_));
 sg13g2_nor3_2 _0978_ (.A(_0273_),
    .B(_0275_),
    .C(_0276_),
    .Y(_0277_));
 sg13g2_or3_2 _0979_ (.A(_0273_),
    .B(_0275_),
    .C(_0276_),
    .X(_0278_));
 sg13g2_xor2_1 _0980_ (.B(_0266_),
    .A(_0014_),
    .X(_0279_));
 sg13g2_nor4_2 _0981_ (.A(_0259_),
    .B(_0260_),
    .C(_0268_),
    .Y(_0280_),
    .D(_0279_));
 sg13g2_o21ai_1 _0982_ (.B1(_0232_),
    .Y(_0281_),
    .A1(_0225_),
    .A2(_0233_));
 sg13g2_o21ai_1 _0983_ (.B1(_0229_),
    .Y(_0282_),
    .A1(_0226_),
    .A2(_0228_));
 sg13g2_xor2_1 _0984_ (.B(_0282_),
    .A(\system_inst.neuron.v_mem[8] ),
    .X(_0283_));
 sg13g2_xnor2_1 _0985_ (.Y(_0284_),
    .A(_0281_),
    .B(_0283_));
 sg13g2_a21oi_2 _0986_ (.B1(_0284_),
    .Y(_0285_),
    .A2(_0280_),
    .A1(_0253_));
 sg13g2_a21o_2 _0987_ (.A2(_0280_),
    .A1(_0253_),
    .B1(_0284_),
    .X(_0286_));
 sg13g2_nor2_2 _0988_ (.A(_0277_),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_nor2_1 _0989_ (.A(\system_inst.leak_rate_1[7] ),
    .B(_0239_),
    .Y(_0288_));
 sg13g2_nor3_2 _0990_ (.A(_0277_),
    .B(_0286_),
    .C(_0288_),
    .Y(_0289_));
 sg13g2_nor2_1 _0991_ (.A(_0015_),
    .B(_0287_),
    .Y(_0290_));
 sg13g2_a21oi_2 _0992_ (.B1(_0290_),
    .Y(_0291_),
    .A2(_0289_),
    .A1(_0240_));
 sg13g2_nand2_1 _0993_ (.Y(_0292_),
    .A(_0234_),
    .B(_0291_));
 sg13g2_xnor2_1 _0994_ (.Y(_0293_),
    .A(_0234_),
    .B(_0291_));
 sg13g2_inv_1 _0995_ (.Y(_0294_),
    .A(_0293_));
 sg13g2_xnor2_1 _0996_ (.Y(_0295_),
    .A(\system_inst.leak_rate_1[6] ),
    .B(_0238_));
 sg13g2_nor2_1 _0997_ (.A(_0016_),
    .B(_0287_),
    .Y(_0296_));
 sg13g2_a21oi_1 _0998_ (.A1(_0287_),
    .A2(_0295_),
    .Y(_0297_),
    .B1(_0296_));
 sg13g2_nand2_1 _0999_ (.Y(_0298_),
    .A(_0241_),
    .B(_0297_));
 sg13g2_xnor2_1 _1000_ (.Y(_0299_),
    .A(_0241_),
    .B(_0297_));
 sg13g2_xnor2_1 _1001_ (.Y(_0300_),
    .A(\system_inst.leak_rate_1[1] ),
    .B(\system_inst.leak_rate_1[0] ));
 sg13g2_a21oi_1 _1002_ (.A1(_0278_),
    .A2(_0285_),
    .Y(_0301_),
    .B1(_0021_));
 sg13g2_nor3_1 _1003_ (.A(_0277_),
    .B(_0286_),
    .C(_0300_),
    .Y(_0302_));
 sg13g2_nor3_1 _1004_ (.A(_0263_),
    .B(_0301_),
    .C(_0302_),
    .Y(_0303_));
 sg13g2_nand2_1 _1005_ (.Y(_0304_),
    .A(\system_inst.leak_rate_1[0] ),
    .B(_0266_));
 sg13g2_o21ai_1 _1006_ (.B1(_0263_),
    .Y(_0305_),
    .A1(_0301_),
    .A2(_0302_));
 sg13g2_nor2b_1 _1007_ (.A(_0303_),
    .B_N(_0305_),
    .Y(_0306_));
 sg13g2_a21oi_2 _1008_ (.B1(_0303_),
    .Y(_0307_),
    .A2(_0305_),
    .A1(_0304_));
 sg13g2_o21ai_1 _1009_ (.B1(_0019_),
    .Y(_0308_),
    .A1(_0277_),
    .A2(_0286_));
 sg13g2_xnor2_1 _1010_ (.Y(_0309_),
    .A(\system_inst.leak_rate_1[3] ),
    .B(_0235_));
 sg13g2_nand3_1 _1011_ (.B(_0285_),
    .C(_0309_),
    .A(_0278_),
    .Y(_0310_));
 sg13g2_a21oi_1 _1012_ (.A1(_0278_),
    .A2(_0285_),
    .Y(_0311_),
    .B1(_0019_));
 sg13g2_nor3_1 _1013_ (.A(_0277_),
    .B(_0286_),
    .C(_0309_),
    .Y(_0312_));
 sg13g2_and3_1 _1014_ (.X(_0313_),
    .A(_0255_),
    .B(_0308_),
    .C(_0310_));
 sg13g2_o21ai_1 _1015_ (.B1(_0255_),
    .Y(_0314_),
    .A1(_0311_),
    .A2(_0312_));
 sg13g2_nor3_1 _1016_ (.A(_0255_),
    .B(_0311_),
    .C(_0312_),
    .Y(_0315_));
 sg13g2_nor2_1 _1017_ (.A(_0313_),
    .B(_0315_),
    .Y(_0316_));
 sg13g2_o21ai_1 _1018_ (.B1(\system_inst.leak_rate_1[2] ),
    .Y(_0317_),
    .A1(\system_inst.leak_rate_1[1] ),
    .A2(\system_inst.leak_rate_1[0] ));
 sg13g2_a21o_1 _1019_ (.A2(_0285_),
    .A1(_0278_),
    .B1(_0020_),
    .X(_0318_));
 sg13g2_nand4_1 _1020_ (.B(_0278_),
    .C(_0285_),
    .A(_0235_),
    .Y(_0319_),
    .D(_0317_));
 sg13g2_and3_1 _1021_ (.X(_0320_),
    .A(_0258_),
    .B(_0318_),
    .C(_0319_));
 sg13g2_nand3_1 _1022_ (.B(_0318_),
    .C(_0319_),
    .A(_0258_),
    .Y(_0321_));
 sg13g2_a21oi_1 _1023_ (.A1(_0318_),
    .A2(_0319_),
    .Y(_0322_),
    .B1(_0258_));
 sg13g2_or2_1 _1024_ (.X(_0323_),
    .B(_0322_),
    .A(_0320_));
 sg13g2_or4_1 _1025_ (.A(_0313_),
    .B(_0315_),
    .C(_0320_),
    .D(_0322_),
    .X(_0324_));
 sg13g2_a21oi_1 _1026_ (.A1(_0314_),
    .A2(_0320_),
    .Y(_0325_),
    .B1(_0315_));
 sg13g2_o21ai_1 _1027_ (.B1(_0325_),
    .Y(_0326_),
    .A1(_0307_),
    .A2(_0324_));
 sg13g2_xor2_1 _1028_ (.B(_0236_),
    .A(\system_inst.leak_rate_1[4] ),
    .X(_0327_));
 sg13g2_mux2_1 _1029_ (.A0(_0018_),
    .A1(_0327_),
    .S(_0287_),
    .X(_0328_));
 sg13g2_and2_1 _1030_ (.A(_0248_),
    .B(_0328_),
    .X(_0329_));
 sg13g2_xor2_1 _1031_ (.B(_0328_),
    .A(_0248_),
    .X(_0330_));
 sg13g2_xor2_1 _1032_ (.B(_0237_),
    .A(\system_inst.leak_rate_1[5] ),
    .X(_0331_));
 sg13g2_mux2_1 _1033_ (.A0(_0017_),
    .A1(_0331_),
    .S(_0287_),
    .X(_0332_));
 sg13g2_and2_1 _1034_ (.A(_0246_),
    .B(_0332_),
    .X(_0333_));
 sg13g2_or2_1 _1035_ (.X(_0334_),
    .B(_0332_),
    .A(_0246_));
 sg13g2_xor2_1 _1036_ (.B(_0332_),
    .A(_0246_),
    .X(_0335_));
 sg13g2_and2_1 _1037_ (.A(_0330_),
    .B(_0335_),
    .X(_0336_));
 sg13g2_a221oi_1 _1038_ (.B2(_0326_),
    .C1(_0333_),
    .B1(_0336_),
    .A1(_0329_),
    .Y(_0337_),
    .A2(_0334_));
 sg13g2_o21ai_1 _1039_ (.B1(_0298_),
    .Y(_0338_),
    .A1(_0299_),
    .A2(_0337_));
 sg13g2_nand2b_1 _1040_ (.Y(_0339_),
    .B(_0293_),
    .A_N(_0338_));
 sg13g2_nand2b_1 _1041_ (.Y(_0340_),
    .B(\system_inst.leak_cycles_1[3] ),
    .A_N(\system_inst.neuron.leak_counter_1[3] ));
 sg13g2_nor2b_1 _1042_ (.A(\system_inst.leak_cycles_1[3] ),
    .B_N(\system_inst.neuron.leak_counter_1[3] ),
    .Y(_0341_));
 sg13g2_nor2b_1 _1043_ (.A(\system_inst.neuron.leak_counter_1[2] ),
    .B_N(\system_inst.leak_cycles_1[2] ),
    .Y(_0342_));
 sg13g2_nand2b_1 _1044_ (.Y(_0343_),
    .B(\system_inst.neuron.leak_counter_1[2] ),
    .A_N(\system_inst.leak_cycles_1[2] ));
 sg13g2_nand2_1 _1045_ (.Y(_0344_),
    .A(_0109_),
    .B(\system_inst.neuron.leak_counter_1[1] ));
 sg13g2_nand3b_1 _1046_ (.B(_0344_),
    .C(\system_inst.leak_cycles_1[0] ),
    .Y(_0345_),
    .A_N(\system_inst.neuron.leak_counter_1[0] ));
 sg13g2_o21ai_1 _1047_ (.B1(_0345_),
    .Y(_0346_),
    .A1(_0109_),
    .A2(\system_inst.neuron.leak_counter_1[1] ));
 sg13g2_a21oi_1 _1048_ (.A1(_0343_),
    .A2(_0346_),
    .Y(_0347_),
    .B1(_0342_));
 sg13g2_a21o_1 _1049_ (.A2(_0347_),
    .A1(_0340_),
    .B1(_0341_),
    .X(_0348_));
 sg13g2_a21oi_2 _1050_ (.B1(_0341_),
    .Y(_0349_),
    .A2(_0347_),
    .A1(_0340_));
 sg13g2_a21oi_1 _1051_ (.A1(_0294_),
    .A2(_0338_),
    .Y(_0350_),
    .B1(_0349_));
 sg13g2_a22oi_1 _1052_ (.Y(_0351_),
    .B1(_0350_),
    .B2(_0339_),
    .A2(_0349_),
    .A1(_0234_));
 sg13g2_nor3_1 _1053_ (.A(\system_inst.leak_rate_2[2] ),
    .B(\system_inst.leak_rate_2[1] ),
    .C(\system_inst.leak_rate_2[0] ),
    .Y(_0352_));
 sg13g2_nor2b_1 _1054_ (.A(\system_inst.leak_rate_2[3] ),
    .B_N(_0352_),
    .Y(_0353_));
 sg13g2_nor2b_1 _1055_ (.A(\system_inst.leak_rate_2[4] ),
    .B_N(_0353_),
    .Y(_0354_));
 sg13g2_nor2b_1 _1056_ (.A(\system_inst.leak_rate_2[5] ),
    .B_N(_0354_),
    .Y(_0355_));
 sg13g2_nor2b_1 _1057_ (.A(\system_inst.leak_rate_2[6] ),
    .B_N(_0355_),
    .Y(_0356_));
 sg13g2_nand2b_1 _1058_ (.Y(_0357_),
    .B(\system_inst.leak_rate_2[7] ),
    .A_N(_0356_));
 sg13g2_xnor2_1 _1059_ (.Y(_0358_),
    .A(_0299_),
    .B(_0337_));
 sg13g2_nor2_1 _1060_ (.A(_0241_),
    .B(net111),
    .Y(_0359_));
 sg13g2_a21oi_2 _1061_ (.B1(_0359_),
    .Y(_0360_),
    .A2(_0358_),
    .A1(net111));
 sg13g2_xor2_1 _1062_ (.B(_0360_),
    .A(_0009_),
    .X(_0361_));
 sg13g2_a21oi_1 _1063_ (.A1(_0326_),
    .A2(_0330_),
    .Y(_0362_),
    .B1(_0329_));
 sg13g2_nor2_1 _1064_ (.A(_0246_),
    .B(net111),
    .Y(_0363_));
 sg13g2_xor2_1 _1065_ (.B(_0362_),
    .A(_0335_),
    .X(_0364_));
 sg13g2_a21oi_2 _1066_ (.B1(_0363_),
    .Y(_0365_),
    .A2(_0364_),
    .A1(net111));
 sg13g2_or2_1 _1067_ (.X(_0366_),
    .B(_0365_),
    .A(_0010_));
 sg13g2_nand2_1 _1068_ (.Y(_0367_),
    .A(_0010_),
    .B(_0365_));
 sg13g2_xnor2_1 _1069_ (.Y(_0368_),
    .A(_0326_),
    .B(_0330_));
 sg13g2_nor2_1 _1070_ (.A(_0248_),
    .B(net111),
    .Y(_0369_));
 sg13g2_a21oi_2 _1071_ (.B1(_0369_),
    .Y(_0370_),
    .A2(_0368_),
    .A1(net111));
 sg13g2_or2_1 _1072_ (.X(_0371_),
    .B(_0370_),
    .A(_0011_));
 sg13g2_xnor2_1 _1073_ (.Y(_0372_),
    .A(_0011_),
    .B(_0370_));
 sg13g2_a21oi_1 _1074_ (.A1(_0010_),
    .A2(_0365_),
    .Y(_0373_),
    .B1(_0372_));
 sg13g2_and4_1 _1075_ (.A(_0351_),
    .B(_0361_),
    .C(_0366_),
    .D(_0373_),
    .X(_0374_));
 sg13g2_o21ai_1 _1076_ (.B1(_0321_),
    .Y(_0375_),
    .A1(_0307_),
    .A2(_0323_));
 sg13g2_xor2_1 _1077_ (.B(_0375_),
    .A(_0316_),
    .X(_0376_));
 sg13g2_nand2_1 _1078_ (.Y(_0377_),
    .A(_0255_),
    .B(_0349_));
 sg13g2_o21ai_1 _1079_ (.B1(_0377_),
    .Y(_0378_),
    .A1(_0349_),
    .A2(_0376_));
 sg13g2_inv_1 _1080_ (.Y(_0379_),
    .A(_0378_));
 sg13g2_and2_1 _1081_ (.A(\system_inst.loader.threshold[4] ),
    .B(_0378_),
    .X(_0380_));
 sg13g2_nand2_1 _1082_ (.Y(_0381_),
    .A(\system_inst.loader.threshold[4] ),
    .B(_0378_));
 sg13g2_nor2_1 _1083_ (.A(\system_inst.loader.threshold[4] ),
    .B(_0378_),
    .Y(_0382_));
 sg13g2_nor2_1 _1084_ (.A(_0258_),
    .B(net112),
    .Y(_0383_));
 sg13g2_xnor2_1 _1085_ (.Y(_0384_),
    .A(_0307_),
    .B(_0323_));
 sg13g2_a21oi_2 _1086_ (.B1(_0383_),
    .Y(_0385_),
    .A2(_0384_),
    .A1(net111));
 sg13g2_xnor2_1 _1087_ (.Y(_0386_),
    .A(_0012_),
    .B(_0385_));
 sg13g2_nor3_1 _1088_ (.A(_0380_),
    .B(_0382_),
    .C(_0386_),
    .Y(_0387_));
 sg13g2_nand2_1 _1089_ (.Y(_0388_),
    .A(\system_inst.leak_rate_1[0] ),
    .B(net112));
 sg13g2_xnor2_1 _1090_ (.Y(_0389_),
    .A(_0266_),
    .B(_0388_));
 sg13g2_xnor2_1 _1091_ (.Y(_0390_),
    .A(_0304_),
    .B(_0306_));
 sg13g2_nor2_1 _1092_ (.A(_0262_),
    .B(net112),
    .Y(_0391_));
 sg13g2_a21oi_2 _1093_ (.B1(_0391_),
    .Y(_0392_),
    .A2(_0390_),
    .A1(net112));
 sg13g2_xor2_1 _1094_ (.B(_0392_),
    .A(_0013_),
    .X(_0393_));
 sg13g2_o21ai_1 _1095_ (.B1(_0393_),
    .Y(_0394_),
    .A1(\system_inst.loader.threshold[1] ),
    .A2(_0389_));
 sg13g2_o21ai_1 _1096_ (.B1(_0394_),
    .Y(_0395_),
    .A1(_0112_),
    .A2(_0392_));
 sg13g2_nand2b_1 _1097_ (.Y(_0396_),
    .B(\system_inst.loader.threshold[3] ),
    .A_N(_0385_));
 sg13g2_a21oi_1 _1098_ (.A1(_0381_),
    .A2(_0396_),
    .Y(_0397_),
    .B1(_0382_));
 sg13g2_a21o_1 _1099_ (.A2(_0395_),
    .A1(_0387_),
    .B1(_0397_),
    .X(_0398_));
 sg13g2_o21ai_1 _1100_ (.B1(_0371_),
    .Y(_0399_),
    .A1(_0010_),
    .A2(_0365_));
 sg13g2_and4_1 _1101_ (.A(_0351_),
    .B(_0361_),
    .C(_0367_),
    .D(_0399_),
    .X(_0400_));
 sg13g2_nor2_1 _1102_ (.A(_0110_),
    .B(_0360_),
    .Y(_0401_));
 sg13g2_a221oi_1 _1103_ (.B2(_0351_),
    .C1(_0400_),
    .B1(_0401_),
    .A1(_0374_),
    .Y(_0402_),
    .A2(_0398_));
 sg13g2_xor2_1 _1104_ (.B(_0388_),
    .A(_0279_),
    .X(_0403_));
 sg13g2_and3_1 _1105_ (.X(_0404_),
    .A(_0387_),
    .B(_0393_),
    .C(_0403_));
 sg13g2_nand2_1 _1106_ (.Y(_0405_),
    .A(_0292_),
    .B(_0350_));
 sg13g2_a21oi_1 _1107_ (.A1(_0289_),
    .A2(net111),
    .Y(_0406_),
    .B1(_0284_));
 sg13g2_xor2_1 _1108_ (.B(_0406_),
    .A(_0405_),
    .X(_0407_));
 sg13g2_a21oi_1 _1109_ (.A1(_0374_),
    .A2(_0404_),
    .Y(_0408_),
    .B1(_0407_));
 sg13g2_a21o_2 _1110_ (.A2(_0404_),
    .A1(_0374_),
    .B1(_0407_),
    .X(_0409_));
 sg13g2_nor2_2 _1111_ (.A(_0402_),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_nand2b_1 _1112_ (.Y(_0411_),
    .B(_0356_),
    .A_N(\system_inst.leak_rate_2[7] ));
 sg13g2_and2_1 _1113_ (.A(_0410_),
    .B(_0411_),
    .X(_0412_));
 sg13g2_nand3_1 _1114_ (.B(_0410_),
    .C(_0411_),
    .A(_0357_),
    .Y(_0413_));
 sg13g2_o21ai_1 _1115_ (.B1(_0413_),
    .Y(_0414_),
    .A1(_0022_),
    .A2(_0410_));
 sg13g2_xor2_1 _1116_ (.B(_0414_),
    .A(_0351_),
    .X(_0415_));
 sg13g2_xor2_1 _1117_ (.B(\system_inst.leak_rate_2[0] ),
    .A(\system_inst.leak_rate_2[1] ),
    .X(_0416_));
 sg13g2_o21ai_1 _1118_ (.B1(_0121_),
    .Y(_0417_),
    .A1(_0402_),
    .A2(_0409_));
 sg13g2_nand3b_1 _1119_ (.B(_0408_),
    .C(_0416_),
    .Y(_0418_),
    .A_N(_0402_));
 sg13g2_nand3_1 _1120_ (.B(_0417_),
    .C(_0418_),
    .A(_0392_),
    .Y(_0419_));
 sg13g2_nand2_1 _1121_ (.Y(_0420_),
    .A(\system_inst.leak_rate_2[0] ),
    .B(_0389_));
 sg13g2_inv_1 _1122_ (.Y(_0421_),
    .A(_0420_));
 sg13g2_a21oi_1 _1123_ (.A1(_0417_),
    .A2(_0418_),
    .Y(_0422_),
    .B1(_0392_));
 sg13g2_a21o_1 _1124_ (.A2(_0418_),
    .A1(_0417_),
    .B1(_0392_),
    .X(_0423_));
 sg13g2_and3_1 _1125_ (.X(_0424_),
    .A(_0419_),
    .B(_0420_),
    .C(_0423_));
 sg13g2_o21ai_1 _1126_ (.B1(_0419_),
    .Y(_0425_),
    .A1(_0421_),
    .A2(_0422_));
 sg13g2_o21ai_1 _1127_ (.B1(\system_inst.leak_rate_2[2] ),
    .Y(_0426_),
    .A1(\system_inst.leak_rate_2[1] ),
    .A2(\system_inst.leak_rate_2[0] ));
 sg13g2_nor2b_1 _1128_ (.A(_0352_),
    .B_N(_0426_),
    .Y(_0427_));
 sg13g2_o21ai_1 _1129_ (.B1(_0120_),
    .Y(_0428_),
    .A1(_0402_),
    .A2(_0409_));
 sg13g2_nand3b_1 _1130_ (.B(_0408_),
    .C(_0427_),
    .Y(_0429_),
    .A_N(_0402_));
 sg13g2_and3_1 _1131_ (.X(_0430_),
    .A(_0385_),
    .B(_0428_),
    .C(_0429_));
 sg13g2_a21oi_1 _1132_ (.A1(_0428_),
    .A2(_0429_),
    .Y(_0431_),
    .B1(_0385_));
 sg13g2_nor2_1 _1133_ (.A(_0430_),
    .B(_0431_),
    .Y(_0432_));
 sg13g2_nor2b_1 _1134_ (.A(_0352_),
    .B_N(\system_inst.leak_rate_2[3] ),
    .Y(_0433_));
 sg13g2_o21ai_1 _1135_ (.B1(_0119_),
    .Y(_0434_),
    .A1(_0402_),
    .A2(_0409_));
 sg13g2_or4_1 _1136_ (.A(_0353_),
    .B(_0402_),
    .C(_0409_),
    .D(_0433_),
    .X(_0435_));
 sg13g2_a21oi_1 _1137_ (.A1(_0434_),
    .A2(_0435_),
    .Y(_0436_),
    .B1(_0379_));
 sg13g2_a21o_1 _1138_ (.A2(_0435_),
    .A1(_0434_),
    .B1(_0379_),
    .X(_0437_));
 sg13g2_and3_1 _1139_ (.X(_0438_),
    .A(_0379_),
    .B(_0434_),
    .C(_0435_));
 sg13g2_or2_1 _1140_ (.X(_0439_),
    .B(_0438_),
    .A(_0436_));
 sg13g2_nor4_1 _1141_ (.A(_0430_),
    .B(_0431_),
    .C(_0436_),
    .D(_0438_),
    .Y(_0440_));
 sg13g2_a221oi_1 _1142_ (.B2(_0425_),
    .C1(_0438_),
    .B1(_0440_),
    .A1(_0430_),
    .Y(_0441_),
    .A2(_0437_));
 sg13g2_xor2_1 _1143_ (.B(_0353_),
    .A(\system_inst.leak_rate_2[4] ),
    .X(_0442_));
 sg13g2_mux2_1 _1144_ (.A0(_0025_),
    .A1(_0442_),
    .S(_0410_),
    .X(_0443_));
 sg13g2_and2_1 _1145_ (.A(_0370_),
    .B(_0443_),
    .X(_0444_));
 sg13g2_nand2_1 _1146_ (.Y(_0445_),
    .A(_0370_),
    .B(_0443_));
 sg13g2_xnor2_1 _1147_ (.Y(_0446_),
    .A(_0370_),
    .B(_0443_));
 sg13g2_xor2_1 _1148_ (.B(_0354_),
    .A(\system_inst.leak_rate_2[5] ),
    .X(_0447_));
 sg13g2_mux2_1 _1149_ (.A0(_0024_),
    .A1(_0447_),
    .S(_0410_),
    .X(_0448_));
 sg13g2_or2_1 _1150_ (.X(_0449_),
    .B(_0448_),
    .A(_0365_));
 sg13g2_and2_1 _1151_ (.A(_0365_),
    .B(_0448_),
    .X(_0450_));
 sg13g2_xor2_1 _1152_ (.B(_0448_),
    .A(_0365_),
    .X(_0451_));
 sg13g2_nand2b_1 _1153_ (.Y(_0452_),
    .B(_0451_),
    .A_N(_0446_));
 sg13g2_a21oi_1 _1154_ (.A1(_0444_),
    .A2(_0449_),
    .Y(_0453_),
    .B1(_0450_));
 sg13g2_o21ai_1 _1155_ (.B1(_0453_),
    .Y(_0454_),
    .A1(_0441_),
    .A2(_0452_));
 sg13g2_xor2_1 _1156_ (.B(_0355_),
    .A(\system_inst.leak_rate_2[6] ),
    .X(_0455_));
 sg13g2_mux2_1 _1157_ (.A0(_0023_),
    .A1(_0455_),
    .S(_0410_),
    .X(_0456_));
 sg13g2_nand2_1 _1158_ (.Y(_0457_),
    .A(_0360_),
    .B(_0456_));
 sg13g2_inv_1 _1159_ (.Y(_0458_),
    .A(_0457_));
 sg13g2_xor2_1 _1160_ (.B(_0456_),
    .A(_0360_),
    .X(_0459_));
 sg13g2_and2_1 _1161_ (.A(_0415_),
    .B(_0459_),
    .X(_0460_));
 sg13g2_a21oi_1 _1162_ (.A1(_0351_),
    .A2(_0414_),
    .Y(_0461_),
    .B1(_0457_));
 sg13g2_nor2_1 _1163_ (.A(\system_inst.leak_cycles_2[1] ),
    .B(_0117_),
    .Y(_0462_));
 sg13g2_nand2b_1 _1164_ (.Y(_0463_),
    .B(\system_inst.leak_cycles_2[0] ),
    .A_N(\system_inst.neuron.leak_counter_2[0] ));
 sg13g2_a22oi_1 _1165_ (.Y(_0464_),
    .B1(_0117_),
    .B2(\system_inst.leak_cycles_2[1] ),
    .A2(_0116_),
    .A1(\system_inst.leak_cycles_2[2] ));
 sg13g2_o21ai_1 _1166_ (.B1(_0464_),
    .Y(_0465_),
    .A1(_0462_),
    .A2(_0463_));
 sg13g2_a22oi_1 _1167_ (.Y(_0466_),
    .B1(\system_inst.neuron.leak_counter_2[2] ),
    .B2(_0107_),
    .A2(\system_inst.neuron.leak_counter_2[3] ),
    .A1(_0106_));
 sg13g2_nand2_1 _1168_ (.Y(_0467_),
    .A(_0465_),
    .B(_0466_));
 sg13g2_o21ai_1 _1169_ (.B1(_0467_),
    .Y(_0468_),
    .A1(_0106_),
    .A2(\system_inst.neuron.leak_counter_2[3] ));
 sg13g2_inv_1 _1170_ (.Y(_0469_),
    .A(_0468_));
 sg13g2_o21ai_1 _1171_ (.B1(net110),
    .Y(_0470_),
    .A1(_0351_),
    .A2(_0414_));
 sg13g2_or2_1 _1172_ (.X(_0471_),
    .B(_0470_),
    .A(_0461_));
 sg13g2_a21o_1 _1173_ (.A2(_0460_),
    .A1(_0454_),
    .B1(_0471_),
    .X(_0472_));
 sg13g2_a21oi_1 _1174_ (.A1(_0412_),
    .A2(net110),
    .Y(_0473_),
    .B1(_0407_));
 sg13g2_xor2_1 _1175_ (.B(_0473_),
    .A(_0472_),
    .X(_0474_));
 sg13g2_xnor2_1 _1176_ (.Y(_0475_),
    .A(_0472_),
    .B(_0473_));
 sg13g2_xnor2_1 _1177_ (.Y(_0476_),
    .A(_0454_),
    .B(_0459_));
 sg13g2_nand2_1 _1178_ (.Y(_0477_),
    .A(_0360_),
    .B(_0468_));
 sg13g2_o21ai_1 _1179_ (.B1(_0477_),
    .Y(_0478_),
    .A1(_0468_),
    .A2(_0476_));
 sg13g2_nand2_1 _1180_ (.Y(_0479_),
    .A(net108),
    .B(_0478_));
 sg13g2_xnor2_1 _1181_ (.Y(_0480_),
    .A(\system_inst.loader.threshold[6] ),
    .B(_0479_));
 sg13g2_a21oi_1 _1182_ (.A1(_0454_),
    .A2(_0459_),
    .Y(_0481_),
    .B1(_0458_));
 sg13g2_or2_1 _1183_ (.X(_0482_),
    .B(_0481_),
    .A(_0415_));
 sg13g2_a21oi_1 _1184_ (.A1(_0415_),
    .A2(_0481_),
    .Y(_0483_),
    .B1(_0468_));
 sg13g2_a221oi_1 _1185_ (.B2(_0483_),
    .C1(_0474_),
    .B1(_0482_),
    .A1(_0351_),
    .Y(_0484_),
    .A2(_0468_));
 sg13g2_nand2_1 _1186_ (.Y(_0485_),
    .A(_0009_),
    .B(_0484_));
 sg13g2_nor2_1 _1187_ (.A(_0009_),
    .B(_0484_),
    .Y(_0486_));
 sg13g2_xnor2_1 _1188_ (.Y(_0487_),
    .A(_0009_),
    .B(_0484_));
 sg13g2_nor2_1 _1189_ (.A(_0480_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_nor2_1 _1190_ (.A(_0365_),
    .B(net110),
    .Y(_0489_));
 sg13g2_o21ai_1 _1191_ (.B1(_0445_),
    .Y(_0490_),
    .A1(_0441_),
    .A2(_0446_));
 sg13g2_xnor2_1 _1192_ (.Y(_0491_),
    .A(_0451_),
    .B(_0490_));
 sg13g2_a21oi_1 _1193_ (.A1(net110),
    .A2(_0491_),
    .Y(_0492_),
    .B1(_0489_));
 sg13g2_nand2_1 _1194_ (.Y(_0493_),
    .A(net108),
    .B(_0492_));
 sg13g2_xor2_1 _1195_ (.B(_0493_),
    .A(_0011_),
    .X(_0494_));
 sg13g2_xor2_1 _1196_ (.B(_0446_),
    .A(_0441_),
    .X(_0495_));
 sg13g2_mux2_1 _1197_ (.A0(_0370_),
    .A1(_0495_),
    .S(net110),
    .X(_0496_));
 sg13g2_nand2_1 _1198_ (.Y(_0497_),
    .A(net108),
    .B(_0496_));
 sg13g2_nand2_1 _1199_ (.Y(_0498_),
    .A(\system_inst.loader.threshold[4] ),
    .B(_0497_));
 sg13g2_xnor2_1 _1200_ (.Y(_0499_),
    .A(\system_inst.loader.threshold[4] ),
    .B(_0497_));
 sg13g2_nor4_2 _1201_ (.A(_0480_),
    .B(_0487_),
    .C(_0494_),
    .Y(_0500_),
    .D(_0499_));
 sg13g2_a21oi_1 _1202_ (.A1(_0425_),
    .A2(_0432_),
    .Y(_0501_),
    .B1(_0430_));
 sg13g2_nand2_1 _1203_ (.Y(_0502_),
    .A(_0439_),
    .B(_0501_));
 sg13g2_nor2_1 _1204_ (.A(_0439_),
    .B(_0501_),
    .Y(_0503_));
 sg13g2_nand3b_1 _1205_ (.B(_0469_),
    .C(_0502_),
    .Y(_0504_),
    .A_N(_0503_));
 sg13g2_o21ai_1 _1206_ (.B1(_0504_),
    .Y(_0505_),
    .A1(_0378_),
    .A2(net110));
 sg13g2_and2_1 _1207_ (.A(net108),
    .B(_0505_),
    .X(_0506_));
 sg13g2_a21o_1 _1208_ (.A2(_0505_),
    .A1(net107),
    .B1(_0012_),
    .X(_0507_));
 sg13g2_nand3_1 _1209_ (.B(net107),
    .C(_0505_),
    .A(_0012_),
    .Y(_0508_));
 sg13g2_xor2_1 _1210_ (.B(_0432_),
    .A(_0425_),
    .X(_0509_));
 sg13g2_mux2_1 _1211_ (.A0(_0385_),
    .A1(_0509_),
    .S(net110),
    .X(_0510_));
 sg13g2_and2_1 _1212_ (.A(net107),
    .B(_0510_),
    .X(_0511_));
 sg13g2_nand2_1 _1213_ (.Y(_0512_),
    .A(net107),
    .B(_0510_));
 sg13g2_nand3_1 _1214_ (.B(net107),
    .C(_0510_),
    .A(_0112_),
    .Y(_0513_));
 sg13g2_a21o_1 _1215_ (.A2(_0510_),
    .A1(net107),
    .B1(_0112_),
    .X(_0514_));
 sg13g2_nand4_1 _1216_ (.B(_0508_),
    .C(_0513_),
    .A(_0507_),
    .Y(_0515_),
    .D(_0514_));
 sg13g2_nor2_1 _1217_ (.A(_0113_),
    .B(_0468_),
    .Y(_0516_));
 sg13g2_xnor2_1 _1218_ (.Y(_0517_),
    .A(_0389_),
    .B(_0516_));
 sg13g2_nand2_1 _1219_ (.Y(_0518_),
    .A(net108),
    .B(_0517_));
 sg13g2_nand3b_1 _1220_ (.B(_0475_),
    .C(_0517_),
    .Y(_0519_),
    .A_N(\system_inst.loader.threshold[0] ));
 sg13g2_nand2b_1 _1221_ (.Y(_0520_),
    .B(_0468_),
    .A_N(_0392_));
 sg13g2_a21oi_1 _1222_ (.A1(_0419_),
    .A2(_0423_),
    .Y(_0521_),
    .B1(_0420_));
 sg13g2_o21ai_1 _1223_ (.B1(net110),
    .Y(_0522_),
    .A1(_0424_),
    .A2(_0521_));
 sg13g2_and2_1 _1224_ (.A(_0520_),
    .B(_0522_),
    .X(_0523_));
 sg13g2_and2_1 _1225_ (.A(net107),
    .B(_0523_),
    .X(_0524_));
 sg13g2_and3_1 _1226_ (.X(_0525_),
    .A(\system_inst.loader.threshold[1] ),
    .B(net108),
    .C(_0523_));
 sg13g2_a21oi_1 _1227_ (.A1(net107),
    .A2(_0523_),
    .Y(_0526_),
    .B1(\system_inst.loader.threshold[1] ));
 sg13g2_o21ai_1 _1228_ (.B1(_0519_),
    .Y(_0527_),
    .A1(_0525_),
    .A2(_0526_));
 sg13g2_or2_1 _1229_ (.X(_0528_),
    .B(_0524_),
    .A(_0014_));
 sg13g2_a21oi_1 _1230_ (.A1(_0527_),
    .A2(_0528_),
    .Y(_0529_),
    .B1(_0515_));
 sg13g2_o21ai_1 _1231_ (.B1(_0507_),
    .Y(_0530_),
    .A1(_0013_),
    .A2(_0511_));
 sg13g2_and2_1 _1232_ (.A(_0508_),
    .B(_0530_),
    .X(_0531_));
 sg13g2_o21ai_1 _1233_ (.B1(_0500_),
    .Y(_0532_),
    .A1(_0529_),
    .A2(_0531_));
 sg13g2_nand2_1 _1234_ (.Y(_0533_),
    .A(\system_inst.loader.threshold[5] ),
    .B(_0493_));
 sg13g2_o21ai_1 _1235_ (.B1(_0533_),
    .Y(_0534_),
    .A1(_0494_),
    .A2(_0498_));
 sg13g2_a21oi_1 _1236_ (.A1(net108),
    .A2(_0478_),
    .Y(_0535_),
    .B1(_0010_));
 sg13g2_a221oi_1 _1237_ (.B2(_0485_),
    .C1(_0486_),
    .B1(_0535_),
    .A1(_0488_),
    .Y(_0536_),
    .A2(_0534_));
 sg13g2_and2_1 _1238_ (.A(\system_inst.loader.threshold[0] ),
    .B(_0518_),
    .X(_0537_));
 sg13g2_nor3_1 _1239_ (.A(_0515_),
    .B(_0527_),
    .C(_0537_),
    .Y(_0538_));
 sg13g2_a22oi_1 _1240_ (.Y(_0539_),
    .B1(_0538_),
    .B2(_0500_),
    .A2(_0536_),
    .A1(_0532_));
 sg13g2_or3_2 _1241_ (.A(\system_inst.neuron.refr_cnt[2] ),
    .B(\system_inst.neuron.refr_cnt[1] ),
    .C(\system_inst.neuron.refr_cnt[0] ),
    .X(_0540_));
 sg13g2_nor2_1 _1242_ (.A(\system_inst.neuron.refr_cnt[3] ),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_and2_1 _1243_ (.A(params_ready),
    .B(net1),
    .X(_0542_));
 sg13g2_nand2_2 _1244_ (.Y(_0543_),
    .A(params_ready),
    .B(net1));
 sg13g2_nand2_1 _1245_ (.Y(_0544_),
    .A(net2),
    .B(_0542_));
 sg13g2_nor3_2 _1246_ (.A(net155),
    .B(_0540_),
    .C(_0544_),
    .Y(_0545_));
 sg13g2_nand3_1 _1247_ (.B(_0541_),
    .C(_0542_),
    .A(net2),
    .Y(_0546_));
 sg13g2_nor3_1 _1248_ (.A(net132),
    .B(net106),
    .C(net114),
    .Y(_0031_));
 sg13g2_o21ai_1 _1249_ (.B1(net137),
    .Y(_0547_),
    .A1(_0468_),
    .A2(_0543_));
 sg13g2_xnor2_1 _1250_ (.Y(_0548_),
    .A(net197),
    .B(net126));
 sg13g2_nor2_1 _1251_ (.A(_0547_),
    .B(_0548_),
    .Y(_0032_));
 sg13g2_and3_1 _1252_ (.X(_0549_),
    .A(net105),
    .B(net197),
    .C(net126));
 sg13g2_a21oi_1 _1253_ (.A1(\system_inst.neuron.leak_counter_2[0] ),
    .A2(net126),
    .Y(_0550_),
    .B1(net105));
 sg13g2_nor3_1 _1254_ (.A(_0547_),
    .B(_0549_),
    .C(net142),
    .Y(_0033_));
 sg13g2_nand2_1 _1255_ (.Y(_0551_),
    .A(\system_inst.neuron.leak_counter_2[2] ),
    .B(_0549_));
 sg13g2_xnor2_1 _1256_ (.Y(_0552_),
    .A(net204),
    .B(_0549_));
 sg13g2_nor2_1 _1257_ (.A(_0547_),
    .B(_0552_),
    .Y(_0034_));
 sg13g2_xor2_1 _1258_ (.B(_0551_),
    .A(net190),
    .X(_0553_));
 sg13g2_nor2_1 _1259_ (.A(_0547_),
    .B(net191),
    .Y(_0035_));
 sg13g2_nor2_1 _1260_ (.A(_0518_),
    .B(net114),
    .Y(_0554_));
 sg13g2_a22oi_1 _1261_ (.Y(_0555_),
    .B1(_0554_),
    .B2(_0539_),
    .A2(net114),
    .A1(net146));
 sg13g2_nor2_1 _1262_ (.A(net131),
    .B(_0555_),
    .Y(_0036_));
 sg13g2_nand2_1 _1263_ (.Y(_0556_),
    .A(net169),
    .B(net114));
 sg13g2_nand3_1 _1264_ (.B(net106),
    .C(_0545_),
    .A(_0524_),
    .Y(_0557_));
 sg13g2_a21oi_1 _1265_ (.A1(_0556_),
    .A2(_0557_),
    .Y(_0037_),
    .B1(net131));
 sg13g2_nor2_1 _1266_ (.A(_0512_),
    .B(net114),
    .Y(_0558_));
 sg13g2_a22oi_1 _1267_ (.Y(_0559_),
    .B1(_0558_),
    .B2(net106),
    .A2(net113),
    .A1(net192));
 sg13g2_nor2_1 _1268_ (.A(net131),
    .B(_0559_),
    .Y(_0038_));
 sg13g2_nand2_1 _1269_ (.Y(_0560_),
    .A(net208),
    .B(net114));
 sg13g2_nand3_1 _1270_ (.B(net106),
    .C(_0545_),
    .A(_0506_),
    .Y(_0561_));
 sg13g2_a21oi_1 _1271_ (.A1(_0560_),
    .A2(_0561_),
    .Y(_0039_),
    .B1(net131));
 sg13g2_nor2_1 _1272_ (.A(_0497_),
    .B(net113),
    .Y(_0562_));
 sg13g2_a22oi_1 _1273_ (.Y(_0563_),
    .B1(_0562_),
    .B2(net106),
    .A2(net113),
    .A1(net216));
 sg13g2_nor2_1 _1274_ (.A(net131),
    .B(_0563_),
    .Y(_0040_));
 sg13g2_nor2_1 _1275_ (.A(_0493_),
    .B(net113),
    .Y(_0564_));
 sg13g2_a22oi_1 _1276_ (.Y(_0565_),
    .B1(_0564_),
    .B2(net106),
    .A2(net113),
    .A1(net193));
 sg13g2_nor2_1 _1277_ (.A(net131),
    .B(_0565_),
    .Y(_0041_));
 sg13g2_nor2_1 _1278_ (.A(_0479_),
    .B(net113),
    .Y(_0566_));
 sg13g2_a22oi_1 _1279_ (.Y(_0567_),
    .B1(_0566_),
    .B2(net106),
    .A2(net113),
    .A1(net183));
 sg13g2_nor2_1 _1280_ (.A(net131),
    .B(_0567_),
    .Y(_0042_));
 sg13g2_nand2_1 _1281_ (.Y(_0568_),
    .A(net101),
    .B(net114));
 sg13g2_nand3_1 _1282_ (.B(net106),
    .C(_0545_),
    .A(_0484_),
    .Y(_0569_));
 sg13g2_a21oi_1 _1283_ (.A1(_0568_),
    .A2(_0569_),
    .Y(_0043_),
    .B1(net131));
 sg13g2_and3_1 _1284_ (.X(_0044_),
    .A(net129),
    .B(net136),
    .C(net113));
 sg13g2_o21ai_1 _1285_ (.B1(net126),
    .Y(_0570_),
    .A1(\system_inst.neuron.refr_cnt[3] ),
    .A2(_0540_));
 sg13g2_o21ai_1 _1286_ (.B1(_0570_),
    .Y(_0571_),
    .A1(_0539_),
    .A2(_0544_));
 sg13g2_o21ai_1 _1287_ (.B1(_0571_),
    .Y(_0572_),
    .A1(net236),
    .A2(_0541_));
 sg13g2_o21ai_1 _1288_ (.B1(net141),
    .Y(_0573_),
    .A1(net236),
    .A2(_0571_));
 sg13g2_nor2b_1 _1289_ (.A(_0573_),
    .B_N(_0572_),
    .Y(_0045_));
 sg13g2_xor2_1 _1290_ (.B(\system_inst.neuron.refr_cnt[0] ),
    .A(net231),
    .X(_0574_));
 sg13g2_o21ai_1 _1291_ (.B1(_0571_),
    .Y(_0575_),
    .A1(_0541_),
    .A2(_0574_));
 sg13g2_o21ai_1 _1292_ (.B1(net140),
    .Y(_0576_),
    .A1(net231),
    .A2(_0571_));
 sg13g2_nor2b_1 _1293_ (.A(_0576_),
    .B_N(_0575_),
    .Y(_0046_));
 sg13g2_o21ai_1 _1294_ (.B1(net185),
    .Y(_0577_),
    .A1(\system_inst.neuron.refr_cnt[1] ),
    .A2(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_nand3_1 _1295_ (.B(net126),
    .C(_0577_),
    .A(_0540_),
    .Y(_0578_));
 sg13g2_o21ai_1 _1296_ (.B1(net140),
    .Y(_0579_),
    .A1(net185),
    .A2(_0571_));
 sg13g2_nor2b_1 _1297_ (.A(_0579_),
    .B_N(_0578_),
    .Y(_0047_));
 sg13g2_o21ai_1 _1298_ (.B1(net155),
    .Y(_0580_),
    .A1(_0540_),
    .A2(_0543_));
 sg13g2_nor2_1 _1299_ (.A(net133),
    .B(net156),
    .Y(_0048_));
 sg13g2_o21ai_1 _1300_ (.B1(net138),
    .Y(_0581_),
    .A1(_0349_),
    .A2(_0543_));
 sg13g2_xnor2_1 _1301_ (.Y(_0582_),
    .A(net196),
    .B(net126));
 sg13g2_nor2_1 _1302_ (.A(_0581_),
    .B(_0582_),
    .Y(_0049_));
 sg13g2_and3_1 _1303_ (.X(_0583_),
    .A(net150),
    .B(net196),
    .C(net126));
 sg13g2_a21oi_1 _1304_ (.A1(\system_inst.neuron.leak_counter_1[0] ),
    .A2(net126),
    .Y(_0584_),
    .B1(net150));
 sg13g2_nor3_1 _1305_ (.A(_0581_),
    .B(_0583_),
    .C(net151),
    .Y(_0050_));
 sg13g2_nand2_1 _1306_ (.Y(_0585_),
    .A(\system_inst.neuron.leak_counter_1[2] ),
    .B(_0583_));
 sg13g2_xnor2_1 _1307_ (.Y(_0586_),
    .A(net206),
    .B(_0583_));
 sg13g2_nor2_1 _1308_ (.A(_0581_),
    .B(_0586_),
    .Y(_0051_));
 sg13g2_xor2_1 _1309_ (.B(_0585_),
    .A(net194),
    .X(_0587_));
 sg13g2_nor2_1 _1310_ (.A(_0581_),
    .B(net195),
    .Y(_0052_));
 sg13g2_or2_1 _1311_ (.X(_0588_),
    .B(\system_inst.loader.current_state[4] ),
    .A(\system_inst.loader.current_state[2] ));
 sg13g2_nor4_2 _1312_ (.A(\system_inst.loader.current_state[1] ),
    .B(\system_inst.loader.current_state[6] ),
    .C(\system_inst.loader.current_state[5] ),
    .Y(_0589_),
    .D(_0588_));
 sg13g2_nand2_1 _1313_ (.Y(_0590_),
    .A(_0030_),
    .B(_0589_));
 sg13g2_nor2_1 _1314_ (.A(net153),
    .B(_0590_),
    .Y(_0591_));
 sg13g2_o21ai_1 _1315_ (.B1(net1),
    .Y(_0592_),
    .A1(_0123_),
    .A2(net3));
 sg13g2_nor2_1 _1316_ (.A(_0591_),
    .B(_0592_),
    .Y(_0593_));
 sg13g2_o21ai_1 _1317_ (.B1(_0589_),
    .Y(_0594_),
    .A1(_0124_),
    .A2(net125));
 sg13g2_nand2_1 _1318_ (.Y(_0595_),
    .A(net3),
    .B(_0594_));
 sg13g2_nand2_1 _1319_ (.Y(_0596_),
    .A(_0593_),
    .B(_0595_));
 sg13g2_and2_1 _1320_ (.A(_0124_),
    .B(_0589_),
    .X(_0597_));
 sg13g2_a21oi_1 _1321_ (.A1(net210),
    .A2(_0596_),
    .Y(_0598_),
    .B1(net133));
 sg13g2_o21ai_1 _1322_ (.B1(_0598_),
    .Y(_0053_),
    .A1(_0596_),
    .A2(_0597_));
 sg13g2_o21ai_1 _1323_ (.B1(net140),
    .Y(_0599_),
    .A1(net4),
    .A2(_0132_));
 sg13g2_a21oi_1 _1324_ (.A1(_0115_),
    .A2(_0132_),
    .Y(_0054_),
    .B1(_0599_));
 sg13g2_a21oi_1 _1325_ (.A1(net234),
    .A2(_0132_),
    .Y(_0600_),
    .B1(net133));
 sg13g2_o21ai_1 _1326_ (.B1(_0600_),
    .Y(_0055_),
    .A1(_0105_),
    .A2(_0132_));
 sg13g2_o21ai_1 _1327_ (.B1(net140),
    .Y(_0601_),
    .A1(net228),
    .A2(_0133_));
 sg13g2_a21oi_1 _1328_ (.A1(_0104_),
    .A2(_0133_),
    .Y(_0056_),
    .B1(_0601_));
 sg13g2_o21ai_1 _1329_ (.B1(net139),
    .Y(_0602_),
    .A1(net239),
    .A2(net121));
 sg13g2_a21oi_1 _1330_ (.A1(_0108_),
    .A2(net121),
    .Y(_0057_),
    .B1(_0602_));
 sg13g2_a21oi_1 _1331_ (.A1(\system_inst.loader.shift_reg[0] ),
    .A2(net121),
    .Y(_0603_),
    .B1(net132));
 sg13g2_o21ai_1 _1332_ (.B1(_0603_),
    .Y(_0058_),
    .A1(_0114_),
    .A2(net121));
 sg13g2_o21ai_1 _1333_ (.B1(net135),
    .Y(_0604_),
    .A1(net202),
    .A2(net120));
 sg13g2_a21oi_1 _1334_ (.A1(_0104_),
    .A2(net120),
    .Y(_0059_),
    .B1(_0604_));
 sg13g2_o21ai_1 _1335_ (.B1(net135),
    .Y(_0605_),
    .A1(net233),
    .A2(net120));
 sg13g2_a21oi_1 _1336_ (.A1(_0103_),
    .A2(net120),
    .Y(_0060_),
    .B1(_0605_));
 sg13g2_o21ai_1 _1337_ (.B1(net136),
    .Y(_0606_),
    .A1(net212),
    .A2(net119));
 sg13g2_a21oi_1 _1338_ (.A1(_0102_),
    .A2(net119),
    .Y(_0061_),
    .B1(_0606_));
 sg13g2_o21ai_1 _1339_ (.B1(net136),
    .Y(_0607_),
    .A1(net207),
    .A2(net119));
 sg13g2_a21oi_1 _1340_ (.A1(_0101_),
    .A2(net119),
    .Y(_0062_),
    .B1(_0607_));
 sg13g2_o21ai_1 _1341_ (.B1(net134),
    .Y(_0608_),
    .A1(net189),
    .A2(net119));
 sg13g2_a21oi_1 _1342_ (.A1(_0100_),
    .A2(net119),
    .Y(_0063_),
    .B1(_0608_));
 sg13g2_o21ai_1 _1343_ (.B1(net134),
    .Y(_0609_),
    .A1(net209),
    .A2(net119));
 sg13g2_a21oi_1 _1344_ (.A1(_0099_),
    .A2(net119),
    .Y(_0064_),
    .B1(_0609_));
 sg13g2_a21oi_1 _1345_ (.A1(net4),
    .A2(net118),
    .Y(_0610_),
    .B1(net133));
 sg13g2_o21ai_1 _1346_ (.B1(_0610_),
    .Y(_0065_),
    .A1(_0113_),
    .A2(net118));
 sg13g2_o21ai_1 _1347_ (.B1(net135),
    .Y(_0611_),
    .A1(net225),
    .A2(net117));
 sg13g2_a21oi_1 _1348_ (.A1(_0105_),
    .A2(net117),
    .Y(_0066_),
    .B1(_0611_));
 sg13g2_o21ai_1 _1349_ (.B1(net134),
    .Y(_0612_),
    .A1(net200),
    .A2(net116));
 sg13g2_a21oi_1 _1350_ (.A1(_0104_),
    .A2(net116),
    .Y(_0067_),
    .B1(_0612_));
 sg13g2_o21ai_1 _1351_ (.B1(net135),
    .Y(_0613_),
    .A1(net184),
    .A2(net116));
 sg13g2_a21oi_1 _1352_ (.A1(_0103_),
    .A2(net116),
    .Y(_0068_),
    .B1(_0613_));
 sg13g2_o21ai_1 _1353_ (.B1(net134),
    .Y(_0614_),
    .A1(net226),
    .A2(net115));
 sg13g2_a21oi_1 _1354_ (.A1(_0102_),
    .A2(net115),
    .Y(_0069_),
    .B1(_0614_));
 sg13g2_o21ai_1 _1355_ (.B1(net135),
    .Y(_0615_),
    .A1(net220),
    .A2(net115));
 sg13g2_a21oi_1 _1356_ (.A1(_0101_),
    .A2(net115),
    .Y(_0070_),
    .B1(_0615_));
 sg13g2_o21ai_1 _1357_ (.B1(net136),
    .Y(_0616_),
    .A1(net188),
    .A2(net115));
 sg13g2_a21oi_1 _1358_ (.A1(_0100_),
    .A2(net115),
    .Y(_0071_),
    .B1(_0616_));
 sg13g2_o21ai_1 _1359_ (.B1(net136),
    .Y(_0617_),
    .A1(net199),
    .A2(net115));
 sg13g2_a21oi_1 _1360_ (.A1(_0099_),
    .A2(net115),
    .Y(_0072_),
    .B1(_0617_));
 sg13g2_o21ai_1 _1361_ (.B1(net141),
    .Y(_0618_),
    .A1(net224),
    .A2(net123));
 sg13g2_a21oi_1 _1362_ (.A1(_0108_),
    .A2(net123),
    .Y(_0073_),
    .B1(_0618_));
 sg13g2_a21oi_1 _1363_ (.A1(net229),
    .A2(_0139_),
    .Y(_0619_),
    .B1(_0122_));
 sg13g2_o21ai_1 _1364_ (.B1(_0619_),
    .Y(_0074_),
    .A1(_0105_),
    .A2(_0139_));
 sg13g2_a21oi_1 _1365_ (.A1(net223),
    .A2(net123),
    .Y(_0620_),
    .B1(net132));
 sg13g2_o21ai_1 _1366_ (.B1(_0620_),
    .Y(_0075_),
    .A1(_0112_),
    .A2(net123));
 sg13g2_a21oi_1 _1367_ (.A1(net218),
    .A2(_0139_),
    .Y(_0621_),
    .B1(net133));
 sg13g2_o21ai_1 _1368_ (.B1(_0621_),
    .Y(_0076_),
    .A1(_0103_),
    .A2(_0139_));
 sg13g2_a21oi_1 _1369_ (.A1(net217),
    .A2(net122),
    .Y(_0622_),
    .B1(net132));
 sg13g2_o21ai_1 _1370_ (.B1(_0622_),
    .Y(_0077_),
    .A1(_0111_),
    .A2(net122));
 sg13g2_o21ai_1 _1371_ (.B1(net136),
    .Y(_0623_),
    .A1(net172),
    .A2(net122));
 sg13g2_a21oi_1 _1372_ (.A1(_0101_),
    .A2(net122),
    .Y(_0078_),
    .B1(_0623_));
 sg13g2_o21ai_1 _1373_ (.B1(net136),
    .Y(_0624_),
    .A1(\system_inst.loader.threshold[6] ),
    .A2(net122));
 sg13g2_a21oi_1 _1374_ (.A1(_0100_),
    .A2(net122),
    .Y(_0079_),
    .B1(_0624_));
 sg13g2_o21ai_1 _1375_ (.B1(net134),
    .Y(_0625_),
    .A1(net187),
    .A2(net122));
 sg13g2_a21oi_1 _1376_ (.A1(_0099_),
    .A2(net122),
    .Y(_0080_),
    .B1(_0625_));
 sg13g2_o21ai_1 _1377_ (.B1(net137),
    .Y(_0626_),
    .A1(net164),
    .A2(net124));
 sg13g2_a21oi_1 _1378_ (.A1(_0108_),
    .A2(net124),
    .Y(_0081_),
    .B1(_0626_));
 sg13g2_a21oi_1 _1379_ (.A1(\system_inst.loader.shift_reg[0] ),
    .A2(net124),
    .Y(_0627_),
    .B1(net133));
 sg13g2_o21ai_1 _1380_ (.B1(_0627_),
    .Y(_0082_),
    .A1(_0109_),
    .A2(net124));
 sg13g2_o21ai_1 _1381_ (.B1(net137),
    .Y(_0628_),
    .A1(net178),
    .A2(net124));
 sg13g2_a21oi_1 _1382_ (.A1(_0104_),
    .A2(net124),
    .Y(_0083_),
    .B1(_0628_));
 sg13g2_o21ai_1 _1383_ (.B1(net139),
    .Y(_0629_),
    .A1(net205),
    .A2(net124));
 sg13g2_a21oi_1 _1384_ (.A1(_0103_),
    .A2(net124),
    .Y(_0084_),
    .B1(_0629_));
 sg13g2_and3_2 _1385_ (.X(_0630_),
    .A(net148),
    .B(net130),
    .C(net125));
 sg13g2_o21ai_1 _1386_ (.B1(net137),
    .Y(_0631_),
    .A1(net176),
    .A2(_0630_));
 sg13g2_a21oi_1 _1387_ (.A1(_0108_),
    .A2(_0630_),
    .Y(_0085_),
    .B1(_0631_));
 sg13g2_o21ai_1 _1388_ (.B1(net139),
    .Y(_0632_),
    .A1(net214),
    .A2(_0630_));
 sg13g2_a21oi_1 _1389_ (.A1(_0105_),
    .A2(_0630_),
    .Y(_0086_),
    .B1(_0632_));
 sg13g2_a21oi_1 _1390_ (.A1(\system_inst.loader.shift_reg[1] ),
    .A2(_0630_),
    .Y(_0633_),
    .B1(net133));
 sg13g2_o21ai_1 _1391_ (.B1(_0633_),
    .Y(_0087_),
    .A1(_0107_),
    .A2(_0630_));
 sg13g2_o21ai_1 _1392_ (.B1(net139),
    .Y(_0634_),
    .A1(net162),
    .A2(_0630_));
 sg13g2_a21oi_1 _1393_ (.A1(_0103_),
    .A2(_0630_),
    .Y(_0088_),
    .B1(_0634_));
 sg13g2_nor2_1 _1394_ (.A(net3),
    .B(_0597_),
    .Y(_0635_));
 sg13g2_nor2b_2 _1395_ (.A(_0635_),
    .B_N(_0593_),
    .Y(_0636_));
 sg13g2_nand2b_1 _1396_ (.Y(_0637_),
    .B(_0593_),
    .A_N(_0635_));
 sg13g2_o21ai_1 _1397_ (.B1(_0124_),
    .Y(_0638_),
    .A1(net125),
    .A2(_0589_));
 sg13g2_a21oi_1 _1398_ (.A1(net4),
    .A2(_0638_),
    .Y(_0639_),
    .B1(net109));
 sg13g2_o21ai_1 _1399_ (.B1(net139),
    .Y(_0640_),
    .A1(net221),
    .A2(_0636_));
 sg13g2_nor2_1 _1400_ (.A(_0639_),
    .B(_0640_),
    .Y(_0089_));
 sg13g2_a21oi_1 _1401_ (.A1(net221),
    .A2(_0638_),
    .Y(_0641_),
    .B1(net109));
 sg13g2_o21ai_1 _1402_ (.B1(net139),
    .Y(_0642_),
    .A1(\system_inst.loader.shift_reg[1] ),
    .A2(_0636_));
 sg13g2_nor2_1 _1403_ (.A(_0641_),
    .B(_0642_),
    .Y(_0090_));
 sg13g2_a21oi_1 _1404_ (.A1(net223),
    .A2(_0638_),
    .Y(_0643_),
    .B1(net109));
 sg13g2_o21ai_1 _1405_ (.B1(net135),
    .Y(_0644_),
    .A1(net165),
    .A2(_0636_));
 sg13g2_nor2_1 _1406_ (.A(_0643_),
    .B(_0644_),
    .Y(_0091_));
 sg13g2_a21oi_1 _1407_ (.A1(net165),
    .A2(_0638_),
    .Y(_0645_),
    .B1(net109));
 sg13g2_o21ai_1 _1408_ (.B1(net135),
    .Y(_0646_),
    .A1(\system_inst.loader.shift_reg[3] ),
    .A2(_0636_));
 sg13g2_nor2_1 _1409_ (.A(_0645_),
    .B(_0646_),
    .Y(_0092_));
 sg13g2_a21oi_1 _1410_ (.A1(net217),
    .A2(_0638_),
    .Y(_0647_),
    .B1(net109));
 sg13g2_o21ai_1 _1411_ (.B1(net134),
    .Y(_0648_),
    .A1(net182),
    .A2(_0636_));
 sg13g2_nor2_1 _1412_ (.A(_0647_),
    .B(_0648_),
    .Y(_0093_));
 sg13g2_a21oi_1 _1413_ (.A1(net182),
    .A2(_0638_),
    .Y(_0649_),
    .B1(net109));
 sg13g2_o21ai_1 _1414_ (.B1(net134),
    .Y(_0650_),
    .A1(net180),
    .A2(_0636_));
 sg13g2_nor2_1 _1415_ (.A(_0649_),
    .B(_0650_),
    .Y(_0094_));
 sg13g2_a21oi_1 _1416_ (.A1(\system_inst.loader.shift_reg[5] ),
    .A2(_0638_),
    .Y(_0651_),
    .B1(net109));
 sg13g2_o21ai_1 _1417_ (.B1(net134),
    .Y(_0652_),
    .A1(net167),
    .A2(_0636_));
 sg13g2_nor2_1 _1418_ (.A(_0651_),
    .B(_0652_),
    .Y(_0095_));
 sg13g2_nor2_1 _1419_ (.A(_0597_),
    .B(_0637_),
    .Y(_0653_));
 sg13g2_o21ai_1 _1420_ (.B1(net137),
    .Y(_0654_),
    .A1(net154),
    .A2(_0653_));
 sg13g2_a21oi_1 _1421_ (.A1(net154),
    .A2(_0636_),
    .Y(_0096_),
    .B1(_0654_));
 sg13g2_and2_1 _1422_ (.A(_0590_),
    .B(_0653_),
    .X(_0655_));
 sg13g2_a22oi_1 _1423_ (.Y(_0656_),
    .B1(_0655_),
    .B2(_0129_),
    .A2(net109),
    .A1(net174));
 sg13g2_o21ai_1 _1424_ (.B1(net137),
    .Y(_0657_),
    .A1(net174),
    .A2(net154));
 sg13g2_nor2_1 _1425_ (.A(net175),
    .B(_0657_),
    .Y(_0097_));
 sg13g2_xor2_1 _1426_ (.B(_0129_),
    .A(_0029_),
    .X(_0658_));
 sg13g2_a22oi_1 _1427_ (.Y(_0659_),
    .B1(_0655_),
    .B2(_0658_),
    .A2(_0637_),
    .A1(net144));
 sg13g2_nor2_1 _1428_ (.A(net133),
    .B(net145),
    .Y(_0098_));
 sg13g2_dfrbp_1 _1429_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net27),
    .D(_0031_),
    .Q_N(_0705_),
    .Q(spike_out));
 sg13g2_dfrbp_1 _1430_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net28),
    .D(_0000_),
    .Q_N(_0706_),
    .Q(\system_inst.loader.current_state[0] ));
 sg13g2_dfrbp_1 _1431_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net29),
    .D(_0001_),
    .Q_N(_0707_),
    .Q(\system_inst.loader.current_state[1] ));
 sg13g2_dfrbp_1 _1432_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net30),
    .D(_0002_),
    .Q_N(_0708_),
    .Q(\system_inst.loader.current_state[2] ));
 sg13g2_dfrbp_1 _1433_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net31),
    .D(_0003_),
    .Q_N(_0030_),
    .Q(\system_inst.loader.current_state[3] ));
 sg13g2_dfrbp_1 _1434_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net32),
    .D(net104),
    .Q_N(_0709_),
    .Q(\system_inst.loader.current_state[4] ));
 sg13g2_dfrbp_1 _1435_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net68),
    .D(_0005_),
    .Q_N(_0710_),
    .Q(\system_inst.loader.current_state[5] ));
 sg13g2_dfrbp_1 _1436_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net26),
    .D(_0006_),
    .Q_N(_0704_),
    .Q(\system_inst.loader.current_state[6] ));
 sg13g2_dfrbp_1 _1437_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net75),
    .D(_0032_),
    .Q_N(_0703_),
    .Q(\system_inst.neuron.leak_counter_2[0] ));
 sg13g2_dfrbp_1 _1438_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net73),
    .D(net143),
    .Q_N(_0702_),
    .Q(\system_inst.neuron.leak_counter_2[1] ));
 sg13g2_dfrbp_1 _1439_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net71),
    .D(_0034_),
    .Q_N(_0701_),
    .Q(\system_inst.neuron.leak_counter_2[2] ));
 sg13g2_dfrbp_1 _1440_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net69),
    .D(_0035_),
    .Q_N(_0700_),
    .Q(\system_inst.neuron.leak_counter_2[3] ));
 sg13g2_dfrbp_1 _1441_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net67),
    .D(_0036_),
    .Q_N(_0008_),
    .Q(\system_inst.neuron.v_mem[0] ));
 sg13g2_dfrbp_1 _1442_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net65),
    .D(_0037_),
    .Q_N(_0699_),
    .Q(\system_inst.neuron.v_mem[1] ));
 sg13g2_dfrbp_1 _1443_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net63),
    .D(_0038_),
    .Q_N(_0698_),
    .Q(\system_inst.neuron.v_mem[2] ));
 sg13g2_dfrbp_1 _1444_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net61),
    .D(_0039_),
    .Q_N(_0697_),
    .Q(\system_inst.neuron.v_mem[3] ));
 sg13g2_dfrbp_1 _1445_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net59),
    .D(_0040_),
    .Q_N(_0696_),
    .Q(\system_inst.neuron.v_mem[4] ));
 sg13g2_dfrbp_1 _1446_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net57),
    .D(_0041_),
    .Q_N(_0695_),
    .Q(\system_inst.neuron.v_mem[5] ));
 sg13g2_dfrbp_1 _1447_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net55),
    .D(_0042_),
    .Q_N(_0694_),
    .Q(\system_inst.neuron.v_mem[6] ));
 sg13g2_dfrbp_1 _1448_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net53),
    .D(net102),
    .Q_N(_0007_),
    .Q(\system_inst.neuron.v_mem[7] ));
 sg13g2_dfrbp_1 _1449_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net51),
    .D(_0044_),
    .Q_N(_0693_),
    .Q(\system_inst.neuron.v_mem[8] ));
 sg13g2_dfrbp_1 _1450_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net49),
    .D(_0045_),
    .Q_N(_0692_),
    .Q(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_dfrbp_1 _1451_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net47),
    .D(net232),
    .Q_N(_0691_),
    .Q(\system_inst.neuron.refr_cnt[1] ));
 sg13g2_dfrbp_1 _1452_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net45),
    .D(net186),
    .Q_N(_0690_),
    .Q(\system_inst.neuron.refr_cnt[2] ));
 sg13g2_dfrbp_1 _1453_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net43),
    .D(_0048_),
    .Q_N(_0689_),
    .Q(\system_inst.neuron.refr_cnt[3] ));
 sg13g2_dfrbp_1 _1454_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net41),
    .D(_0049_),
    .Q_N(_0688_),
    .Q(\system_inst.neuron.leak_counter_1[0] ));
 sg13g2_dfrbp_1 _1455_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net39),
    .D(net152),
    .Q_N(_0687_),
    .Q(\system_inst.neuron.leak_counter_1[1] ));
 sg13g2_dfrbp_1 _1456_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net37),
    .D(_0051_),
    .Q_N(_0686_),
    .Q(\system_inst.neuron.leak_counter_1[2] ));
 sg13g2_dfrbp_1 _1457_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net35),
    .D(_0052_),
    .Q_N(_0685_),
    .Q(\system_inst.neuron.leak_counter_1[3] ));
 sg13g2_dfrbp_1 _1458_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net33),
    .D(net211),
    .Q_N(_0684_),
    .Q(params_ready));
 sg13g2_dfrbp_1 _1459_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net99),
    .D(_0054_),
    .Q_N(_0683_),
    .Q(\system_inst.loader.weight_a[0] ));
 sg13g2_dfrbp_1 _1460_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net97),
    .D(_0055_),
    .Q_N(_0682_),
    .Q(\system_inst.loader.weight_a[1] ));
 sg13g2_dfrbp_1 _1461_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net95),
    .D(_0056_),
    .Q_N(_0681_),
    .Q(\system_inst.loader.weight_a[2] ));
 sg13g2_dfrbp_1 _1462_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net93),
    .D(_0057_),
    .Q_N(_0680_),
    .Q(\system_inst.leak_rate_1[0] ));
 sg13g2_dfrbp_1 _1463_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net91),
    .D(net171),
    .Q_N(_0021_),
    .Q(\system_inst.leak_rate_1[1] ));
 sg13g2_dfrbp_1 _1464_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net89),
    .D(net203),
    .Q_N(_0020_),
    .Q(\system_inst.leak_rate_1[2] ));
 sg13g2_dfrbp_1 _1465_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net87),
    .D(_0060_),
    .Q_N(_0019_),
    .Q(\system_inst.leak_rate_1[3] ));
 sg13g2_dfrbp_1 _1466_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net85),
    .D(net213),
    .Q_N(_0018_),
    .Q(\system_inst.leak_rate_1[4] ));
 sg13g2_dfrbp_1 _1467_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net83),
    .D(_0062_),
    .Q_N(_0017_),
    .Q(\system_inst.leak_rate_1[5] ));
 sg13g2_dfrbp_1 _1468_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net81),
    .D(_0063_),
    .Q_N(_0016_),
    .Q(\system_inst.leak_rate_1[6] ));
 sg13g2_dfrbp_1 _1469_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net79),
    .D(_0064_),
    .Q_N(_0015_),
    .Q(\system_inst.leak_rate_1[7] ));
 sg13g2_dfrbp_1 _1470_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net77),
    .D(_0065_),
    .Q_N(_0679_),
    .Q(\system_inst.leak_rate_2[0] ));
 sg13g2_dfrbp_1 _1471_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net74),
    .D(_0066_),
    .Q_N(_0028_),
    .Q(\system_inst.leak_rate_2[1] ));
 sg13g2_dfrbp_1 _1472_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net70),
    .D(net201),
    .Q_N(_0027_),
    .Q(\system_inst.leak_rate_2[2] ));
 sg13g2_dfrbp_1 _1473_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net66),
    .D(_0068_),
    .Q_N(_0026_),
    .Q(\system_inst.leak_rate_2[3] ));
 sg13g2_dfrbp_1 _1474_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net62),
    .D(_0069_),
    .Q_N(_0025_),
    .Q(\system_inst.leak_rate_2[4] ));
 sg13g2_dfrbp_1 _1475_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net58),
    .D(_0070_),
    .Q_N(_0024_),
    .Q(\system_inst.leak_rate_2[5] ));
 sg13g2_dfrbp_1 _1476_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net54),
    .D(_0071_),
    .Q_N(_0023_),
    .Q(\system_inst.leak_rate_2[6] ));
 sg13g2_dfrbp_1 _1477_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net50),
    .D(_0072_),
    .Q_N(_0022_),
    .Q(\system_inst.leak_rate_2[7] ));
 sg13g2_dfrbp_1 _1478_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net46),
    .D(_0073_),
    .Q_N(_0678_),
    .Q(\system_inst.loader.threshold[0] ));
 sg13g2_dfrbp_1 _1479_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net42),
    .D(net230),
    .Q_N(_0014_),
    .Q(\system_inst.loader.threshold[1] ));
 sg13g2_dfrbp_1 _1480_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net38),
    .D(_0075_),
    .Q_N(_0013_),
    .Q(\system_inst.loader.threshold[2] ));
 sg13g2_dfrbp_1 _1481_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net34),
    .D(net219),
    .Q_N(_0012_),
    .Q(\system_inst.loader.threshold[3] ));
 sg13g2_dfrbp_1 _1482_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net98),
    .D(_0077_),
    .Q_N(_0677_),
    .Q(\system_inst.loader.threshold[4] ));
 sg13g2_dfrbp_1 _1483_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net94),
    .D(net173),
    .Q_N(_0011_),
    .Q(\system_inst.loader.threshold[5] ));
 sg13g2_dfrbp_1 _1484_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net90),
    .D(net181),
    .Q_N(_0010_),
    .Q(\system_inst.loader.threshold[6] ));
 sg13g2_dfrbp_1 _1485_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net86),
    .D(_0080_),
    .Q_N(_0009_),
    .Q(\system_inst.loader.threshold[7] ));
 sg13g2_dfrbp_1 _1486_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net82),
    .D(_0081_),
    .Q_N(_0676_),
    .Q(\system_inst.leak_cycles_1[0] ));
 sg13g2_dfrbp_1 _1487_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net78),
    .D(net159),
    .Q_N(_0675_),
    .Q(\system_inst.leak_cycles_1[1] ));
 sg13g2_dfrbp_1 _1488_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net72),
    .D(net179),
    .Q_N(_0674_),
    .Q(\system_inst.leak_cycles_1[2] ));
 sg13g2_dfrbp_1 _1489_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net64),
    .D(_0084_),
    .Q_N(_0673_),
    .Q(\system_inst.leak_cycles_1[3] ));
 sg13g2_dfrbp_1 _1490_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net56),
    .D(_0085_),
    .Q_N(_0672_),
    .Q(\system_inst.leak_cycles_2[0] ));
 sg13g2_dfrbp_1 _1491_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net48),
    .D(net215),
    .Q_N(_0671_),
    .Q(\system_inst.leak_cycles_2[1] ));
 sg13g2_dfrbp_1 _1492_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net40),
    .D(net161),
    .Q_N(_0670_),
    .Q(\system_inst.leak_cycles_2[2] ));
 sg13g2_dfrbp_1 _1493_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net25),
    .D(net163),
    .Q_N(_0669_),
    .Q(\system_inst.leak_cycles_2[3] ));
 sg13g2_dfrbp_1 _1494_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net92),
    .D(_0089_),
    .Q_N(_0668_),
    .Q(\system_inst.loader.shift_reg[0] ));
 sg13g2_dfrbp_1 _1495_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net84),
    .D(net222),
    .Q_N(_0667_),
    .Q(\system_inst.loader.shift_reg[1] ));
 sg13g2_dfrbp_1 _1496_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net76),
    .D(_0091_),
    .Q_N(_0666_),
    .Q(\system_inst.loader.shift_reg[2] ));
 sg13g2_dfrbp_1 _1497_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net60),
    .D(net166),
    .Q_N(_0665_),
    .Q(\system_inst.loader.shift_reg[3] ));
 sg13g2_dfrbp_1 _1498_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net44),
    .D(_0093_),
    .Q_N(_0664_),
    .Q(\system_inst.loader.shift_reg[4] ));
 sg13g2_dfrbp_1 _1499_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net96),
    .D(_0094_),
    .Q_N(_0663_),
    .Q(\system_inst.loader.shift_reg[5] ));
 sg13g2_dfrbp_1 _1500_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net80),
    .D(net168),
    .Q_N(_0662_),
    .Q(\system_inst.loader.shift_reg[6] ));
 sg13g2_dfrbp_1 _1501_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net52),
    .D(_0096_),
    .Q_N(_0661_),
    .Q(\system_inst.loader.bit_count[0] ));
 sg13g2_dfrbp_1 _1502_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net88),
    .D(_0097_),
    .Q_N(_0660_),
    .Q(\system_inst.loader.bit_count[1] ));
 sg13g2_dfrbp_1 _1503_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net36),
    .D(_0098_),
    .Q_N(_0029_),
    .Q(\system_inst.loader.bit_count[2] ));
 sg13g2_tiehi _1436__26 (.L_HI(net26));
 sg13g2_tiehi _1429__27 (.L_HI(net27));
 sg13g2_tiehi _1430__28 (.L_HI(net28));
 sg13g2_tiehi _1431__29 (.L_HI(net29));
 sg13g2_tiehi _1432__30 (.L_HI(net30));
 sg13g2_tiehi _1433__31 (.L_HI(net31));
 sg13g2_tiehi _1434__32 (.L_HI(net32));
 sg13g2_tiehi _1458__33 (.L_HI(net33));
 sg13g2_tiehi _1481__34 (.L_HI(net34));
 sg13g2_tiehi _1457__35 (.L_HI(net35));
 sg13g2_tiehi _1503__36 (.L_HI(net36));
 sg13g2_tiehi _1456__37 (.L_HI(net37));
 sg13g2_tiehi _1480__38 (.L_HI(net38));
 sg13g2_tiehi _1455__39 (.L_HI(net39));
 sg13g2_tiehi _1492__40 (.L_HI(net40));
 sg13g2_tiehi _1454__41 (.L_HI(net41));
 sg13g2_tiehi _1479__42 (.L_HI(net42));
 sg13g2_tiehi _1453__43 (.L_HI(net43));
 sg13g2_tiehi _1498__44 (.L_HI(net44));
 sg13g2_tiehi _1452__45 (.L_HI(net45));
 sg13g2_tiehi _1478__46 (.L_HI(net46));
 sg13g2_tiehi _1451__47 (.L_HI(net47));
 sg13g2_tiehi _1491__48 (.L_HI(net48));
 sg13g2_tiehi _1450__49 (.L_HI(net49));
 sg13g2_tiehi _1477__50 (.L_HI(net50));
 sg13g2_tiehi _1449__51 (.L_HI(net51));
 sg13g2_tiehi _1501__52 (.L_HI(net52));
 sg13g2_tiehi _1448__53 (.L_HI(net53));
 sg13g2_tiehi _1476__54 (.L_HI(net54));
 sg13g2_tiehi _1447__55 (.L_HI(net55));
 sg13g2_tiehi _1490__56 (.L_HI(net56));
 sg13g2_tiehi _1446__57 (.L_HI(net57));
 sg13g2_tiehi _1475__58 (.L_HI(net58));
 sg13g2_tiehi _1445__59 (.L_HI(net59));
 sg13g2_tiehi _1497__60 (.L_HI(net60));
 sg13g2_tiehi _1444__61 (.L_HI(net61));
 sg13g2_tiehi _1474__62 (.L_HI(net62));
 sg13g2_tiehi _1443__63 (.L_HI(net63));
 sg13g2_tiehi _1489__64 (.L_HI(net64));
 sg13g2_tiehi _1442__65 (.L_HI(net65));
 sg13g2_tiehi _1473__66 (.L_HI(net66));
 sg13g2_tiehi _1441__67 (.L_HI(net67));
 sg13g2_tiehi _1435__68 (.L_HI(net68));
 sg13g2_tiehi _1440__69 (.L_HI(net69));
 sg13g2_tiehi _1472__70 (.L_HI(net70));
 sg13g2_tiehi _1439__71 (.L_HI(net71));
 sg13g2_tiehi _1488__72 (.L_HI(net72));
 sg13g2_tiehi _1438__73 (.L_HI(net73));
 sg13g2_tiehi _1471__74 (.L_HI(net74));
 sg13g2_tiehi _1437__75 (.L_HI(net75));
 sg13g2_tiehi _1496__76 (.L_HI(net76));
 sg13g2_tiehi _1470__77 (.L_HI(net77));
 sg13g2_tiehi _1487__78 (.L_HI(net78));
 sg13g2_tiehi _1469__79 (.L_HI(net79));
 sg13g2_tiehi _1500__80 (.L_HI(net80));
 sg13g2_tiehi _1468__81 (.L_HI(net81));
 sg13g2_tiehi _1486__82 (.L_HI(net82));
 sg13g2_tiehi _1467__83 (.L_HI(net83));
 sg13g2_tiehi _1495__84 (.L_HI(net84));
 sg13g2_tiehi _1466__85 (.L_HI(net85));
 sg13g2_tiehi _1485__86 (.L_HI(net86));
 sg13g2_tiehi _1465__87 (.L_HI(net87));
 sg13g2_tiehi _1502__88 (.L_HI(net88));
 sg13g2_tiehi _1464__89 (.L_HI(net89));
 sg13g2_tiehi _1484__90 (.L_HI(net90));
 sg13g2_tiehi _1463__91 (.L_HI(net91));
 sg13g2_tiehi _1494__92 (.L_HI(net92));
 sg13g2_tiehi _1462__93 (.L_HI(net93));
 sg13g2_tiehi _1483__94 (.L_HI(net94));
 sg13g2_tiehi _1461__95 (.L_HI(net95));
 sg13g2_tiehi _1499__96 (.L_HI(net96));
 sg13g2_tiehi _1460__97 (.L_HI(net97));
 sg13g2_tiehi _1482__98 (.L_HI(net98));
 sg13g2_tiehi _1459__99 (.L_HI(net99));
 sg13g2_tiehi tt_um_wokwi_434917200607612929_100 (.L_HI(net100));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_wokwi_434917200607612929_12 (.L_LO(net12));
 sg13g2_tielo tt_um_wokwi_434917200607612929_13 (.L_LO(net13));
 sg13g2_tielo tt_um_wokwi_434917200607612929_14 (.L_LO(net14));
 sg13g2_tielo tt_um_wokwi_434917200607612929_15 (.L_LO(net15));
 sg13g2_tielo tt_um_wokwi_434917200607612929_16 (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_434917200607612929_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_434917200607612929_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_434917200607612929_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_434917200607612929_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_434917200607612929_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_434917200607612929_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_434917200607612929_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_434917200607612929_24 (.L_LO(net24));
 sg13g2_tiehi _1493__25 (.L_HI(net25));
 sg13g2_buf_2 _1594_ (.A(params_ready),
    .X(uio_out[0]));
 sg13g2_buf_1 _1595_ (.A(spike_out),
    .X(uo_out[0]));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(_0539_));
 sg13g2_buf_2 fanout107 (.A(net108),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_0475_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_0637_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_0469_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_0348_),
    .X(net111));
 sg13g2_buf_1 fanout112 (.A(_0348_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(net114),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0546_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(net117),
    .X(net115));
 sg13g2_buf_1 fanout116 (.A(net117),
    .X(net116));
 sg13g2_buf_1 fanout117 (.A(net118),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_0143_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(net121),
    .X(net119));
 sg13g2_buf_1 fanout120 (.A(net121),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_0141_),
    .X(net121));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(_0138_));
 sg13g2_buf_2 fanout123 (.A(_0138_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_0135_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_0130_),
    .X(net125));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(_0542_));
 sg13g2_buf_2 fanout127 (.A(\system_inst.loader.weight_a[2] ),
    .X(net127));
 sg13g2_buf_1 fanout128 (.A(\system_inst.loader.weight_a[2] ),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(net238),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_0125_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_0122_),
    .X(net132));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(_0122_));
 sg13g2_buf_2 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net136));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(rst_n));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net139));
 sg13g2_buf_1 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(net141),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(net141),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(rst_n),
    .X(net141));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_tielo tt_um_wokwi_434917200607612929_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\system_inst.neuron.v_mem[7] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0043_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold3 (.A(\system_inst.loader.current_state[4] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0004_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold5 (.A(\system_inst.neuron.leak_counter_2[1] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0550_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0033_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold8 (.A(\system_inst.loader.bit_count[2] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0659_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold10 (.A(\system_inst.neuron.v_mem[0] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold11 (.A(\system_inst.loader.current_state[2] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold12 (.A(\system_inst.loader.current_state[3] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0136_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold14 (.A(\system_inst.neuron.leak_counter_1[1] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0584_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0050_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold17 (.A(\system_inst.loader.current_state[0] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold18 (.A(\system_inst.loader.bit_count[0] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold19 (.A(\system_inst.neuron.refr_cnt[3] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0580_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold21 (.A(\system_inst.loader.current_state[6] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold22 (.A(\system_inst.leak_cycles_1[1] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0082_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold24 (.A(\system_inst.leak_cycles_2[2] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0087_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold26 (.A(\system_inst.leak_cycles_2[3] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0088_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold28 (.A(\system_inst.leak_cycles_1[0] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold29 (.A(\system_inst.loader.shift_reg[2] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0092_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold31 (.A(\system_inst.loader.shift_reg[6] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0095_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold33 (.A(\system_inst.neuron.v_mem[1] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold34 (.A(\system_inst.leak_rate_1[1] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0058_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold36 (.A(\system_inst.loader.threshold[5] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0078_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold38 (.A(\system_inst.loader.bit_count[1] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0656_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold40 (.A(\system_inst.leak_cycles_2[0] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold41 (.A(\system_inst.loader.current_state[5] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold42 (.A(\system_inst.leak_cycles_1[2] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0083_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold44 (.A(\system_inst.loader.shift_reg[5] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0079_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold46 (.A(\system_inst.loader.shift_reg[4] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold47 (.A(\system_inst.neuron.v_mem[6] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold48 (.A(\system_inst.leak_rate_2[3] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold49 (.A(\system_inst.neuron.refr_cnt[2] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0047_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold51 (.A(\system_inst.loader.threshold[7] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold52 (.A(\system_inst.leak_rate_2[6] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold53 (.A(\system_inst.leak_rate_1[6] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold54 (.A(\system_inst.neuron.leak_counter_2[3] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0553_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold56 (.A(\system_inst.neuron.v_mem[2] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold57 (.A(\system_inst.neuron.v_mem[5] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold58 (.A(\system_inst.neuron.leak_counter_1[3] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0587_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold60 (.A(\system_inst.neuron.leak_counter_1[0] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold61 (.A(\system_inst.neuron.leak_counter_2[0] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold62 (.A(\system_inst.loader.current_state[1] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold63 (.A(\system_inst.leak_rate_2[7] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold64 (.A(\system_inst.leak_rate_2[2] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0067_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold66 (.A(\system_inst.leak_rate_1[2] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0059_),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold68 (.A(\system_inst.neuron.leak_counter_2[2] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold69 (.A(\system_inst.leak_cycles_1[3] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold70 (.A(\system_inst.neuron.leak_counter_1[2] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold71 (.A(\system_inst.leak_rate_1[5] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold72 (.A(\system_inst.neuron.v_mem[3] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold73 (.A(\system_inst.leak_rate_1[7] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold74 (.A(params_ready),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0053_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold76 (.A(\system_inst.leak_rate_1[4] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0061_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold78 (.A(\system_inst.leak_cycles_2[1] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0086_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold80 (.A(\system_inst.neuron.v_mem[4] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold81 (.A(\system_inst.loader.shift_reg[3] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold82 (.A(\system_inst.loader.threshold[3] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0076_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold84 (.A(\system_inst.leak_rate_2[5] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold85 (.A(\system_inst.loader.shift_reg[0] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0090_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold87 (.A(\system_inst.loader.shift_reg[1] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold88 (.A(\system_inst.loader.threshold[0] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold89 (.A(\system_inst.leak_rate_2[1] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold90 (.A(\system_inst.leak_rate_2[4] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold91 (.A(\system_inst.loader.threshold[2] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold92 (.A(\system_inst.loader.weight_a[2] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold93 (.A(\system_inst.loader.threshold[1] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0074_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold95 (.A(\system_inst.neuron.refr_cnt[1] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0046_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold97 (.A(\system_inst.leak_rate_1[3] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold98 (.A(\system_inst.loader.weight_a[1] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold99 (.A(\system_inst.loader.weight_a[0] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold100 (.A(\system_inst.neuron.refr_cnt[0] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold101 (.A(\system_inst.loader.threshold[4] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold102 (.A(\system_inst.neuron.v_mem[8] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold103 (.A(\system_inst.leak_rate_1[0] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold104 (.A(\system_inst.leak_rate_2[0] ),
    .X(net240));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_fill_2 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_230 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_251 ();
 sg13g2_decap_8 FILLER_8_258 ();
 sg13g2_decap_8 FILLER_8_265 ();
 sg13g2_decap_8 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_4 FILLER_9_203 ();
 sg13g2_fill_1 FILLER_9_207 ();
 sg13g2_fill_1 FILLER_9_242 ();
 sg13g2_fill_1 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_319 ();
 sg13g2_decap_4 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_334 ();
 sg13g2_fill_2 FILLER_9_341 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_fill_2 FILLER_9_363 ();
 sg13g2_decap_4 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_4 FILLER_10_203 ();
 sg13g2_fill_1 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_212 ();
 sg13g2_fill_2 FILLER_10_219 ();
 sg13g2_fill_1 FILLER_10_221 ();
 sg13g2_fill_1 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_fill_2 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_fill_1 FILLER_10_324 ();
 sg13g2_decap_4 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_fill_2 FILLER_11_244 ();
 sg13g2_decap_8 FILLER_11_278 ();
 sg13g2_decap_8 FILLER_11_285 ();
 sg13g2_decap_4 FILLER_11_292 ();
 sg13g2_fill_1 FILLER_11_296 ();
 sg13g2_fill_2 FILLER_11_323 ();
 sg13g2_decap_8 FILLER_11_346 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_fill_2 FILLER_12_196 ();
 sg13g2_decap_4 FILLER_12_288 ();
 sg13g2_fill_1 FILLER_12_292 ();
 sg13g2_fill_1 FILLER_12_316 ();
 sg13g2_decap_8 FILLER_12_346 ();
 sg13g2_fill_1 FILLER_12_353 ();
 sg13g2_fill_2 FILLER_12_379 ();
 sg13g2_fill_1 FILLER_12_381 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_4 FILLER_13_203 ();
 sg13g2_fill_2 FILLER_13_207 ();
 sg13g2_fill_1 FILLER_13_222 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_266 ();
 sg13g2_decap_4 FILLER_13_285 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_decap_4 FILLER_13_325 ();
 sg13g2_fill_2 FILLER_13_360 ();
 sg13g2_fill_1 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_4 FILLER_14_105 ();
 sg13g2_fill_2 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_115 ();
 sg13g2_decap_8 FILLER_14_122 ();
 sg13g2_decap_8 FILLER_14_129 ();
 sg13g2_decap_8 FILLER_14_136 ();
 sg13g2_decap_8 FILLER_14_143 ();
 sg13g2_decap_8 FILLER_14_150 ();
 sg13g2_fill_1 FILLER_14_157 ();
 sg13g2_decap_8 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_169 ();
 sg13g2_fill_1 FILLER_14_171 ();
 sg13g2_decap_4 FILLER_14_177 ();
 sg13g2_decap_8 FILLER_14_185 ();
 sg13g2_decap_8 FILLER_14_192 ();
 sg13g2_decap_8 FILLER_14_199 ();
 sg13g2_fill_2 FILLER_14_206 ();
 sg13g2_fill_2 FILLER_14_234 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_decap_4 FILLER_14_280 ();
 sg13g2_fill_2 FILLER_14_310 ();
 sg13g2_fill_1 FILLER_14_312 ();
 sg13g2_fill_1 FILLER_14_330 ();
 sg13g2_decap_4 FILLER_14_340 ();
 sg13g2_fill_1 FILLER_14_344 ();
 sg13g2_fill_2 FILLER_14_362 ();
 sg13g2_fill_1 FILLER_14_364 ();
 sg13g2_fill_1 FILLER_14_370 ();
 sg13g2_fill_2 FILLER_14_380 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_fill_1 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_82 ();
 sg13g2_fill_2 FILLER_15_89 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_fill_2 FILLER_15_173 ();
 sg13g2_fill_1 FILLER_15_175 ();
 sg13g2_decap_4 FILLER_15_215 ();
 sg13g2_decap_8 FILLER_15_223 ();
 sg13g2_fill_1 FILLER_15_230 ();
 sg13g2_decap_4 FILLER_15_244 ();
 sg13g2_fill_2 FILLER_15_253 ();
 sg13g2_fill_1 FILLER_15_255 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_fill_2 FILLER_15_287 ();
 sg13g2_fill_1 FILLER_15_294 ();
 sg13g2_fill_1 FILLER_15_299 ();
 sg13g2_fill_2 FILLER_15_305 ();
 sg13g2_decap_4 FILLER_15_316 ();
 sg13g2_decap_4 FILLER_15_333 ();
 sg13g2_fill_2 FILLER_15_337 ();
 sg13g2_fill_2 FILLER_15_365 ();
 sg13g2_fill_1 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_4 FILLER_16_56 ();
 sg13g2_fill_2 FILLER_16_60 ();
 sg13g2_fill_2 FILLER_16_98 ();
 sg13g2_decap_4 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_114 ();
 sg13g2_decap_8 FILLER_16_130 ();
 sg13g2_decap_4 FILLER_16_142 ();
 sg13g2_decap_8 FILLER_16_150 ();
 sg13g2_fill_1 FILLER_16_194 ();
 sg13g2_fill_1 FILLER_16_214 ();
 sg13g2_fill_1 FILLER_16_224 ();
 sg13g2_fill_1 FILLER_16_234 ();
 sg13g2_decap_8 FILLER_16_258 ();
 sg13g2_fill_1 FILLER_16_269 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_decap_4 FILLER_16_290 ();
 sg13g2_fill_1 FILLER_16_294 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_309 ();
 sg13g2_fill_1 FILLER_16_316 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_4 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_67 ();
 sg13g2_fill_1 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_103 ();
 sg13g2_fill_1 FILLER_17_105 ();
 sg13g2_decap_4 FILLER_17_162 ();
 sg13g2_fill_2 FILLER_17_192 ();
 sg13g2_fill_1 FILLER_17_194 ();
 sg13g2_decap_8 FILLER_17_226 ();
 sg13g2_fill_2 FILLER_17_263 ();
 sg13g2_fill_1 FILLER_17_265 ();
 sg13g2_fill_2 FILLER_17_301 ();
 sg13g2_fill_1 FILLER_17_303 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_56 ();
 sg13g2_fill_1 FILLER_18_83 ();
 sg13g2_fill_1 FILLER_18_93 ();
 sg13g2_fill_2 FILLER_18_108 ();
 sg13g2_fill_1 FILLER_18_110 ();
 sg13g2_fill_2 FILLER_18_148 ();
 sg13g2_fill_2 FILLER_18_169 ();
 sg13g2_fill_1 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_198 ();
 sg13g2_fill_2 FILLER_18_209 ();
 sg13g2_fill_1 FILLER_18_211 ();
 sg13g2_decap_8 FILLER_18_218 ();
 sg13g2_decap_4 FILLER_18_225 ();
 sg13g2_fill_2 FILLER_18_229 ();
 sg13g2_fill_2 FILLER_18_258 ();
 sg13g2_fill_2 FILLER_18_265 ();
 sg13g2_fill_1 FILLER_18_267 ();
 sg13g2_fill_1 FILLER_18_285 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_317 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_decap_4 FILLER_18_335 ();
 sg13g2_fill_1 FILLER_18_339 ();
 sg13g2_fill_1 FILLER_18_348 ();
 sg13g2_fill_2 FILLER_18_359 ();
 sg13g2_fill_2 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_63 ();
 sg13g2_fill_1 FILLER_19_65 ();
 sg13g2_fill_2 FILLER_19_74 ();
 sg13g2_fill_2 FILLER_19_86 ();
 sg13g2_fill_1 FILLER_19_88 ();
 sg13g2_fill_2 FILLER_19_115 ();
 sg13g2_fill_1 FILLER_19_117 ();
 sg13g2_fill_2 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_128 ();
 sg13g2_fill_2 FILLER_19_152 ();
 sg13g2_decap_8 FILLER_19_172 ();
 sg13g2_decap_4 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_4 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_223 ();
 sg13g2_fill_2 FILLER_19_320 ();
 sg13g2_fill_2 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_330 ();
 sg13g2_fill_1 FILLER_19_353 ();
 sg13g2_fill_1 FILLER_19_377 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_4 FILLER_20_49 ();
 sg13g2_fill_2 FILLER_20_53 ();
 sg13g2_fill_2 FILLER_20_81 ();
 sg13g2_decap_4 FILLER_20_92 ();
 sg13g2_fill_1 FILLER_20_96 ();
 sg13g2_decap_4 FILLER_20_115 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_146 ();
 sg13g2_decap_8 FILLER_20_153 ();
 sg13g2_fill_2 FILLER_20_160 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_decap_8 FILLER_20_173 ();
 sg13g2_fill_2 FILLER_20_180 ();
 sg13g2_fill_2 FILLER_20_199 ();
 sg13g2_fill_1 FILLER_20_206 ();
 sg13g2_fill_1 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_225 ();
 sg13g2_fill_2 FILLER_20_237 ();
 sg13g2_fill_1 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_decap_8 FILLER_20_255 ();
 sg13g2_fill_1 FILLER_20_262 ();
 sg13g2_fill_2 FILLER_20_268 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_decap_8 FILLER_20_282 ();
 sg13g2_decap_4 FILLER_20_289 ();
 sg13g2_decap_8 FILLER_20_296 ();
 sg13g2_decap_4 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_324 ();
 sg13g2_decap_8 FILLER_20_331 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_344 ();
 sg13g2_decap_4 FILLER_20_351 ();
 sg13g2_fill_2 FILLER_20_363 ();
 sg13g2_fill_1 FILLER_20_365 ();
 sg13g2_fill_2 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_fill_1 FILLER_21_87 ();
 sg13g2_decap_8 FILLER_21_92 ();
 sg13g2_fill_1 FILLER_21_99 ();
 sg13g2_decap_8 FILLER_21_113 ();
 sg13g2_fill_1 FILLER_21_120 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_4 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_144 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_decap_8 FILLER_21_174 ();
 sg13g2_decap_4 FILLER_21_181 ();
 sg13g2_fill_2 FILLER_21_205 ();
 sg13g2_fill_1 FILLER_21_207 ();
 sg13g2_decap_8 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_250 ();
 sg13g2_fill_2 FILLER_21_288 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_fill_2 FILLER_21_368 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_65 ();
 sg13g2_decap_4 FILLER_22_81 ();
 sg13g2_decap_4 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_145 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_4 FILLER_22_182 ();
 sg13g2_decap_4 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_226 ();
 sg13g2_decap_8 FILLER_22_233 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_fill_2 FILLER_22_271 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_fill_2 FILLER_22_304 ();
 sg13g2_fill_1 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_338 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_decap_4 FILLER_22_350 ();
 sg13g2_fill_2 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_decap_4 FILLER_22_387 ();
 sg13g2_fill_1 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_49 ();
 sg13g2_decap_4 FILLER_23_54 ();
 sg13g2_decap_8 FILLER_23_85 ();
 sg13g2_decap_4 FILLER_23_92 ();
 sg13g2_fill_2 FILLER_23_96 ();
 sg13g2_decap_8 FILLER_23_103 ();
 sg13g2_decap_4 FILLER_23_110 ();
 sg13g2_fill_2 FILLER_23_114 ();
 sg13g2_decap_8 FILLER_23_120 ();
 sg13g2_decap_8 FILLER_23_127 ();
 sg13g2_decap_8 FILLER_23_134 ();
 sg13g2_decap_8 FILLER_23_141 ();
 sg13g2_decap_4 FILLER_23_148 ();
 sg13g2_fill_2 FILLER_23_160 ();
 sg13g2_decap_8 FILLER_23_172 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_decap_4 FILLER_23_186 ();
 sg13g2_decap_4 FILLER_23_207 ();
 sg13g2_fill_1 FILLER_23_211 ();
 sg13g2_fill_2 FILLER_23_221 ();
 sg13g2_fill_2 FILLER_23_231 ();
 sg13g2_decap_4 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_250 ();
 sg13g2_fill_1 FILLER_23_256 ();
 sg13g2_decap_4 FILLER_23_283 ();
 sg13g2_fill_2 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_294 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_fill_1 FILLER_23_301 ();
 sg13g2_fill_1 FILLER_23_311 ();
 sg13g2_fill_1 FILLER_23_317 ();
 sg13g2_fill_2 FILLER_23_331 ();
 sg13g2_fill_2 FILLER_23_350 ();
 sg13g2_decap_4 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_368 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_32 ();
 sg13g2_fill_2 FILLER_24_59 ();
 sg13g2_decap_4 FILLER_24_75 ();
 sg13g2_fill_2 FILLER_24_102 ();
 sg13g2_fill_1 FILLER_24_104 ();
 sg13g2_fill_2 FILLER_24_169 ();
 sg13g2_fill_2 FILLER_24_179 ();
 sg13g2_fill_1 FILLER_24_181 ();
 sg13g2_decap_8 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_238 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_245 ();
 sg13g2_fill_1 FILLER_24_247 ();
 sg13g2_decap_4 FILLER_24_251 ();
 sg13g2_fill_1 FILLER_24_255 ();
 sg13g2_decap_4 FILLER_24_259 ();
 sg13g2_fill_2 FILLER_24_263 ();
 sg13g2_fill_2 FILLER_24_283 ();
 sg13g2_fill_1 FILLER_24_285 ();
 sg13g2_decap_4 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_4 FILLER_24_343 ();
 sg13g2_fill_2 FILLER_24_347 ();
 sg13g2_fill_1 FILLER_24_357 ();
 sg13g2_decap_4 FILLER_24_364 ();
 sg13g2_decap_4 FILLER_24_375 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_48 ();
 sg13g2_fill_1 FILLER_25_55 ();
 sg13g2_fill_1 FILLER_25_68 ();
 sg13g2_decap_4 FILLER_25_94 ();
 sg13g2_decap_8 FILLER_25_103 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_fill_2 FILLER_25_130 ();
 sg13g2_fill_2 FILLER_25_135 ();
 sg13g2_decap_4 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_149 ();
 sg13g2_decap_8 FILLER_25_158 ();
 sg13g2_fill_1 FILLER_25_170 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_4 FILLER_25_182 ();
 sg13g2_fill_2 FILLER_25_186 ();
 sg13g2_decap_8 FILLER_25_205 ();
 sg13g2_decap_4 FILLER_25_212 ();
 sg13g2_decap_4 FILLER_25_236 ();
 sg13g2_decap_4 FILLER_25_252 ();
 sg13g2_decap_4 FILLER_25_273 ();
 sg13g2_fill_2 FILLER_25_277 ();
 sg13g2_decap_4 FILLER_25_284 ();
 sg13g2_fill_2 FILLER_25_288 ();
 sg13g2_decap_4 FILLER_25_304 ();
 sg13g2_fill_1 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_fill_2 FILLER_25_347 ();
 sg13g2_fill_2 FILLER_25_375 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_83 ();
 sg13g2_fill_1 FILLER_26_108 ();
 sg13g2_decap_4 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_179 ();
 sg13g2_decap_4 FILLER_26_185 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_decap_4 FILLER_26_199 ();
 sg13g2_fill_2 FILLER_26_208 ();
 sg13g2_fill_2 FILLER_26_221 ();
 sg13g2_fill_1 FILLER_26_223 ();
 sg13g2_decap_4 FILLER_26_236 ();
 sg13g2_fill_2 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_264 ();
 sg13g2_fill_2 FILLER_26_281 ();
 sg13g2_fill_1 FILLER_26_283 ();
 sg13g2_decap_8 FILLER_26_310 ();
 sg13g2_decap_8 FILLER_26_317 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_fill_2 FILLER_26_336 ();
 sg13g2_fill_2 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_40 ();
 sg13g2_fill_2 FILLER_27_47 ();
 sg13g2_fill_1 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_65 ();
 sg13g2_decap_8 FILLER_27_72 ();
 sg13g2_fill_2 FILLER_27_87 ();
 sg13g2_fill_1 FILLER_27_89 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_decap_8 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_107 ();
 sg13g2_decap_8 FILLER_27_131 ();
 sg13g2_decap_8 FILLER_27_142 ();
 sg13g2_decap_8 FILLER_27_149 ();
 sg13g2_decap_8 FILLER_27_156 ();
 sg13g2_fill_2 FILLER_27_163 ();
 sg13g2_decap_8 FILLER_27_170 ();
 sg13g2_decap_4 FILLER_27_177 ();
 sg13g2_fill_2 FILLER_27_181 ();
 sg13g2_fill_2 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_218 ();
 sg13g2_decap_4 FILLER_27_225 ();
 sg13g2_decap_8 FILLER_27_237 ();
 sg13g2_decap_8 FILLER_27_244 ();
 sg13g2_decap_4 FILLER_27_251 ();
 sg13g2_decap_4 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_decap_8 FILLER_27_331 ();
 sg13g2_decap_4 FILLER_27_338 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_fill_2 FILLER_27_388 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_39 ();
 sg13g2_decap_4 FILLER_28_46 ();
 sg13g2_fill_1 FILLER_28_50 ();
 sg13g2_fill_2 FILLER_28_69 ();
 sg13g2_decap_4 FILLER_28_85 ();
 sg13g2_decap_8 FILLER_28_124 ();
 sg13g2_decap_4 FILLER_28_152 ();
 sg13g2_decap_8 FILLER_28_176 ();
 sg13g2_decap_4 FILLER_28_183 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_fill_2 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_202 ();
 sg13g2_decap_8 FILLER_28_211 ();
 sg13g2_decap_8 FILLER_28_218 ();
 sg13g2_fill_2 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_237 ();
 sg13g2_decap_8 FILLER_28_244 ();
 sg13g2_fill_2 FILLER_28_251 ();
 sg13g2_decap_8 FILLER_28_269 ();
 sg13g2_decap_4 FILLER_28_276 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_decap_4 FILLER_28_316 ();
 sg13g2_fill_1 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_346 ();
 sg13g2_fill_2 FILLER_28_378 ();
 sg13g2_fill_1 FILLER_28_380 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_fill_2 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_23 ();
 sg13g2_fill_2 FILLER_29_50 ();
 sg13g2_decap_4 FILLER_29_76 ();
 sg13g2_fill_1 FILLER_29_80 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_decap_4 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_4 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_177 ();
 sg13g2_decap_8 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_209 ();
 sg13g2_fill_1 FILLER_29_211 ();
 sg13g2_fill_2 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_248 ();
 sg13g2_fill_2 FILLER_29_255 ();
 sg13g2_fill_1 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_4 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_decap_8 FILLER_29_283 ();
 sg13g2_fill_1 FILLER_29_290 ();
 sg13g2_decap_4 FILLER_29_317 ();
 sg13g2_fill_2 FILLER_29_321 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_fill_2 FILLER_29_374 ();
 sg13g2_fill_2 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_37 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_4 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_101 ();
 sg13g2_decap_8 FILLER_30_107 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_116 ();
 sg13g2_decap_4 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_130 ();
 sg13g2_decap_8 FILLER_30_141 ();
 sg13g2_fill_2 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_150 ();
 sg13g2_decap_4 FILLER_30_156 ();
 sg13g2_decap_8 FILLER_30_165 ();
 sg13g2_decap_8 FILLER_30_172 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_decap_8 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_227 ();
 sg13g2_fill_1 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_254 ();
 sg13g2_decap_8 FILLER_30_260 ();
 sg13g2_fill_2 FILLER_30_267 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_fill_2 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_324 ();
 sg13g2_decap_8 FILLER_30_338 ();
 sg13g2_decap_8 FILLER_30_345 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_25 ();
 sg13g2_fill_2 FILLER_31_53 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_decap_4 FILLER_31_75 ();
 sg13g2_fill_2 FILLER_31_79 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_112 ();
 sg13g2_fill_1 FILLER_31_124 ();
 sg13g2_decap_4 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_183 ();
 sg13g2_decap_8 FILLER_31_190 ();
 sg13g2_decap_8 FILLER_31_202 ();
 sg13g2_fill_2 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_216 ();
 sg13g2_decap_8 FILLER_31_223 ();
 sg13g2_fill_2 FILLER_31_230 ();
 sg13g2_fill_1 FILLER_31_232 ();
 sg13g2_fill_2 FILLER_31_253 ();
 sg13g2_fill_1 FILLER_31_255 ();
 sg13g2_decap_8 FILLER_31_271 ();
 sg13g2_fill_1 FILLER_31_278 ();
 sg13g2_decap_8 FILLER_31_292 ();
 sg13g2_decap_8 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_decap_8 FILLER_31_319 ();
 sg13g2_fill_2 FILLER_31_326 ();
 sg13g2_decap_4 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_31_366 ();
 sg13g2_decap_4 FILLER_31_373 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_fill_2 FILLER_31_392 ();
 sg13g2_decap_4 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_53 ();
 sg13g2_fill_1 FILLER_32_60 ();
 sg13g2_decap_8 FILLER_32_74 ();
 sg13g2_decap_8 FILLER_32_81 ();
 sg13g2_decap_4 FILLER_32_88 ();
 sg13g2_fill_2 FILLER_32_92 ();
 sg13g2_decap_8 FILLER_32_109 ();
 sg13g2_decap_8 FILLER_32_116 ();
 sg13g2_decap_4 FILLER_32_123 ();
 sg13g2_fill_1 FILLER_32_127 ();
 sg13g2_fill_1 FILLER_32_141 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_4 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_164 ();
 sg13g2_decap_8 FILLER_32_171 ();
 sg13g2_fill_1 FILLER_32_178 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_fill_2 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_decap_8 FILLER_32_225 ();
 sg13g2_decap_4 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_256 ();
 sg13g2_decap_4 FILLER_32_296 ();
 sg13g2_fill_1 FILLER_32_300 ();
 sg13g2_decap_8 FILLER_32_317 ();
 sg13g2_decap_4 FILLER_32_324 ();
 sg13g2_fill_2 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_fill_2 FILLER_32_394 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_37 ();
 sg13g2_fill_2 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_117 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_decap_8 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_215 ();
 sg13g2_decap_4 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_4 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_279 ();
 sg13g2_decap_4 FILLER_33_286 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_decap_4 FILLER_33_299 ();
 sg13g2_decap_4 FILLER_33_330 ();
 sg13g2_fill_2 FILLER_33_339 ();
 sg13g2_decap_8 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_53 ();
 sg13g2_decap_4 FILLER_34_60 ();
 sg13g2_decap_8 FILLER_34_73 ();
 sg13g2_decap_8 FILLER_34_80 ();
 sg13g2_decap_4 FILLER_34_87 ();
 sg13g2_fill_2 FILLER_34_100 ();
 sg13g2_decap_8 FILLER_34_106 ();
 sg13g2_decap_8 FILLER_34_144 ();
 sg13g2_decap_8 FILLER_34_151 ();
 sg13g2_fill_2 FILLER_34_158 ();
 sg13g2_fill_1 FILLER_34_160 ();
 sg13g2_decap_8 FILLER_34_185 ();
 sg13g2_decap_4 FILLER_34_192 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_fill_2 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_214 ();
 sg13g2_fill_2 FILLER_34_221 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_decap_4 FILLER_34_263 ();
 sg13g2_fill_2 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_283 ();
 sg13g2_fill_1 FILLER_34_290 ();
 sg13g2_fill_2 FILLER_34_306 ();
 sg13g2_fill_1 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_313 ();
 sg13g2_decap_8 FILLER_34_320 ();
 sg13g2_decap_4 FILLER_34_327 ();
 sg13g2_decap_8 FILLER_34_344 ();
 sg13g2_fill_2 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_decap_4 FILLER_34_359 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_fill_2 FILLER_34_372 ();
 sg13g2_fill_1 FILLER_34_374 ();
 sg13g2_fill_1 FILLER_34_394 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_fill_1 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_127 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_fill_2 FILLER_35_166 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_184 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_fill_1 FILLER_35_196 ();
 sg13g2_fill_2 FILLER_35_237 ();
 sg13g2_fill_1 FILLER_35_239 ();
 sg13g2_decap_4 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_248 ();
 sg13g2_decap_4 FILLER_35_300 ();
 sg13g2_decap_8 FILLER_35_324 ();
 sg13g2_fill_2 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_337 ();
 sg13g2_fill_2 FILLER_35_344 ();
 sg13g2_fill_1 FILLER_35_346 ();
 sg13g2_fill_2 FILLER_35_351 ();
 sg13g2_fill_1 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_370 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_4 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_155 ();
 sg13g2_decap_4 FILLER_36_162 ();
 sg13g2_decap_8 FILLER_36_209 ();
 sg13g2_fill_2 FILLER_36_216 ();
 sg13g2_fill_1 FILLER_36_218 ();
 sg13g2_fill_1 FILLER_36_224 ();
 sg13g2_fill_2 FILLER_36_235 ();
 sg13g2_decap_8 FILLER_36_246 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_fill_2 FILLER_36_270 ();
 sg13g2_decap_8 FILLER_36_277 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_decap_8 FILLER_36_299 ();
 sg13g2_decap_8 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_342 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_fill_1 FILLER_36_355 ();
 sg13g2_decap_8 FILLER_36_360 ();
 sg13g2_fill_2 FILLER_36_367 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_fill_2 FILLER_36_386 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_fill_2 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_decap_4 FILLER_37_237 ();
 sg13g2_fill_2 FILLER_37_241 ();
 sg13g2_decap_4 FILLER_37_247 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_decap_4 FILLER_37_281 ();
 sg13g2_fill_1 FILLER_37_285 ();
 sg13g2_decap_4 FILLER_37_327 ();
 sg13g2_fill_1 FILLER_37_331 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_fill_1 FILLER_37_361 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_fill_2 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_174 ();
 sg13g2_decap_4 FILLER_38_184 ();
 sg13g2_decap_8 FILLER_38_192 ();
 sg13g2_decap_4 FILLER_38_217 ();
 sg13g2_fill_2 FILLER_38_221 ();
 sg13g2_decap_8 FILLER_38_258 ();
 sg13g2_fill_2 FILLER_38_265 ();
 sg13g2_fill_1 FILLER_38_267 ();
 sg13g2_decap_8 FILLER_38_281 ();
 sg13g2_fill_2 FILLER_38_288 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_decap_4 FILLER_38_300 ();
 sg13g2_fill_1 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_fill_2 FILLER_38_389 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net100;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net12;
 assign uio_oe[3] = net13;
 assign uio_oe[4] = net14;
 assign uio_oe[5] = net15;
 assign uio_oe[6] = net16;
 assign uio_oe[7] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule
