module tt_um_emmk_riscv (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire clknet_leaf_0_clk;
 wire \m_sys._GEN_11[3] ;
 wire \m_sys._GEN_11[4] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[0] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[10] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[11] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[1] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[2] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[3] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[4] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[5] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[6] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[7] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[8] ;
 wire \m_sys._m_bootloader_io_b_mem_addr[9] ;
 wire \m_sys._m_bootloader_io_b_mem_wdata[0] ;
 wire \m_sys._m_bootloader_io_b_mem_wdata[1] ;
 wire \m_sys._m_bootloader_io_b_mem_wdata[2] ;
 wire \m_sys._m_bootloader_io_b_mem_wdata[3] ;
 wire \m_sys._m_bootloader_io_b_mem_wdata[4] ;
 wire \m_sys._m_bootloader_io_b_mem_wdata[5] ;
 wire \m_sys._m_bootloader_io_b_mem_wdata[6] ;
 wire \m_sys._m_bootloader_io_b_mem_wdata[7] ;
 wire \m_sys._m_bootloader_io_b_mem_wen[0] ;
 wire \m_sys._m_bootloader_io_o_bl ;
 wire \m_sys._m_core_io_b_mem_wdata[0] ;
 wire \m_sys._m_core_io_b_mem_wdata[10] ;
 wire \m_sys._m_core_io_b_mem_wdata[11] ;
 wire \m_sys._m_core_io_b_mem_wdata[12] ;
 wire \m_sys._m_core_io_b_mem_wdata[13] ;
 wire \m_sys._m_core_io_b_mem_wdata[14] ;
 wire \m_sys._m_core_io_b_mem_wdata[15] ;
 wire \m_sys._m_core_io_b_mem_wdata[16] ;
 wire \m_sys._m_core_io_b_mem_wdata[17] ;
 wire \m_sys._m_core_io_b_mem_wdata[18] ;
 wire \m_sys._m_core_io_b_mem_wdata[19] ;
 wire \m_sys._m_core_io_b_mem_wdata[1] ;
 wire \m_sys._m_core_io_b_mem_wdata[20] ;
 wire \m_sys._m_core_io_b_mem_wdata[21] ;
 wire \m_sys._m_core_io_b_mem_wdata[22] ;
 wire \m_sys._m_core_io_b_mem_wdata[23] ;
 wire \m_sys._m_core_io_b_mem_wdata[24] ;
 wire \m_sys._m_core_io_b_mem_wdata[25] ;
 wire \m_sys._m_core_io_b_mem_wdata[26] ;
 wire \m_sys._m_core_io_b_mem_wdata[27] ;
 wire \m_sys._m_core_io_b_mem_wdata[28] ;
 wire \m_sys._m_core_io_b_mem_wdata[29] ;
 wire \m_sys._m_core_io_b_mem_wdata[2] ;
 wire \m_sys._m_core_io_b_mem_wdata[30] ;
 wire \m_sys._m_core_io_b_mem_wdata[31] ;
 wire \m_sys._m_core_io_b_mem_wdata[3] ;
 wire \m_sys._m_core_io_b_mem_wdata[4] ;
 wire \m_sys._m_core_io_b_mem_wdata[5] ;
 wire \m_sys._m_core_io_b_mem_wdata[6] ;
 wire \m_sys._m_core_io_b_mem_wdata[7] ;
 wire \m_sys._m_core_io_b_mem_wdata[8] ;
 wire \m_sys._m_core_io_b_mem_wdata[9] ;
 wire \m_sys._m_gpio8_io_b_mem_rdata[0] ;
 wire \m_sys._m_gpio8_io_b_mem_rdata[1] ;
 wire \m_sys._m_gpio8_io_b_mem_rdata[2] ;
 wire \m_sys._m_gpio8_io_b_mem_rdata[3] ;
 wire \m_sys._m_gpio8_io_b_mem_rdata[4] ;
 wire \m_sys._m_gpio8_io_b_mem_rdata[5] ;
 wire \m_sys._m_gpio8_io_b_mem_rdata[6] ;
 wire \m_sys._m_gpio8_io_b_mem_rdata[7] ;
 wire \m_sys._m_ram_io_b_port_rdata[0] ;
 wire \m_sys._m_ram_io_b_port_rdata[10] ;
 wire \m_sys._m_ram_io_b_port_rdata[11] ;
 wire \m_sys._m_ram_io_b_port_rdata[12] ;
 wire \m_sys._m_ram_io_b_port_rdata[13] ;
 wire \m_sys._m_ram_io_b_port_rdata[14] ;
 wire \m_sys._m_ram_io_b_port_rdata[15] ;
 wire \m_sys._m_ram_io_b_port_rdata[16] ;
 wire \m_sys._m_ram_io_b_port_rdata[17] ;
 wire \m_sys._m_ram_io_b_port_rdata[18] ;
 wire \m_sys._m_ram_io_b_port_rdata[19] ;
 wire \m_sys._m_ram_io_b_port_rdata[1] ;
 wire \m_sys._m_ram_io_b_port_rdata[20] ;
 wire \m_sys._m_ram_io_b_port_rdata[21] ;
 wire \m_sys._m_ram_io_b_port_rdata[22] ;
 wire \m_sys._m_ram_io_b_port_rdata[23] ;
 wire \m_sys._m_ram_io_b_port_rdata[24] ;
 wire \m_sys._m_ram_io_b_port_rdata[25] ;
 wire \m_sys._m_ram_io_b_port_rdata[26] ;
 wire \m_sys._m_ram_io_b_port_rdata[27] ;
 wire \m_sys._m_ram_io_b_port_rdata[28] ;
 wire \m_sys._m_ram_io_b_port_rdata[29] ;
 wire \m_sys._m_ram_io_b_port_rdata[2] ;
 wire \m_sys._m_ram_io_b_port_rdata[30] ;
 wire \m_sys._m_ram_io_b_port_rdata[31] ;
 wire \m_sys._m_ram_io_b_port_rdata[3] ;
 wire \m_sys._m_ram_io_b_port_rdata[4] ;
 wire \m_sys._m_ram_io_b_port_rdata[5] ;
 wire \m_sys._m_ram_io_b_port_rdata[6] ;
 wire \m_sys._m_ram_io_b_port_rdata[7] ;
 wire \m_sys._m_ram_io_b_port_rdata[8] ;
 wire \m_sys._m_ram_io_b_port_rdata[9] ;
 wire \m_sys._m_uart_io_b_mem_rdata[0] ;
 wire \m_sys._m_uart_io_b_mem_rdata[10] ;
 wire \m_sys._m_uart_io_b_mem_rdata[11] ;
 wire \m_sys._m_uart_io_b_mem_rdata[12] ;
 wire \m_sys._m_uart_io_b_mem_rdata[13] ;
 wire \m_sys._m_uart_io_b_mem_rdata[14] ;
 wire \m_sys._m_uart_io_b_mem_rdata[15] ;
 wire \m_sys._m_uart_io_b_mem_rdata[1] ;
 wire \m_sys._m_uart_io_b_mem_rdata[2] ;
 wire \m_sys._m_uart_io_b_mem_rdata[3] ;
 wire \m_sys._m_uart_io_b_mem_rdata[4] ;
 wire \m_sys._m_uart_io_b_mem_rdata[5] ;
 wire \m_sys._m_uart_io_b_mem_rdata[6] ;
 wire \m_sys._m_uart_io_b_mem_rdata[7] ;
 wire \m_sys._m_uart_io_b_mem_rdata[8] ;
 wire \m_sys._m_uart_io_b_mem_rdata[9] ;
 wire \m_sys._m_uart_io_o_bl_data[0] ;
 wire \m_sys._m_uart_io_o_bl_data[1] ;
 wire \m_sys._m_uart_io_o_bl_data[2] ;
 wire \m_sys._m_uart_io_o_bl_data[3] ;
 wire \m_sys._m_uart_io_o_bl_data[4] ;
 wire \m_sys._m_uart_io_o_bl_data[5] ;
 wire \m_sys._m_uart_io_o_bl_data[6] ;
 wire \m_sys._m_uart_io_o_bl_data[7] ;
 wire \m_sys.io_b_uart_tx ;
 wire \m_sys.m_bootloader._GEN_22[0] ;
 wire \m_sys.m_bootloader._GEN_22[10] ;
 wire \m_sys.m_bootloader._GEN_22[11] ;
 wire \m_sys.m_bootloader._GEN_22[1] ;
 wire \m_sys.m_bootloader._GEN_22[2] ;
 wire \m_sys.m_bootloader._GEN_22[3] ;
 wire \m_sys.m_bootloader._GEN_22[4] ;
 wire \m_sys.m_bootloader._GEN_22[5] ;
 wire \m_sys.m_bootloader._GEN_22[6] ;
 wire \m_sys.m_bootloader._GEN_22[7] ;
 wire \m_sys.m_bootloader._GEN_22[8] ;
 wire \m_sys.m_bootloader._GEN_22[9] ;
 wire \m_sys.m_bootloader.r_byte_cnt[0] ;
 wire \m_sys.m_bootloader.r_byte_cnt[10] ;
 wire \m_sys.m_bootloader.r_byte_cnt[11] ;
 wire \m_sys.m_bootloader.r_byte_cnt[12] ;
 wire \m_sys.m_bootloader.r_byte_cnt[13] ;
 wire \m_sys.m_bootloader.r_byte_cnt[14] ;
 wire \m_sys.m_bootloader.r_byte_cnt[15] ;
 wire \m_sys.m_bootloader.r_byte_cnt[1] ;
 wire \m_sys.m_bootloader.r_byte_cnt[2] ;
 wire \m_sys.m_bootloader.r_byte_cnt[3] ;
 wire \m_sys.m_bootloader.r_byte_cnt[4] ;
 wire \m_sys.m_bootloader.r_byte_cnt[5] ;
 wire \m_sys.m_bootloader.r_byte_cnt[6] ;
 wire \m_sys.m_bootloader.r_byte_cnt[7] ;
 wire \m_sys.m_bootloader.r_byte_cnt[8] ;
 wire \m_sys.m_bootloader.r_byte_cnt[9] ;
 wire \m_sys.m_bootloader.r_cstate[0] ;
 wire \m_sys.m_bootloader.r_cstate[1] ;
 wire \m_sys.m_bootloader.r_cstate[2] ;
 wire \m_sys.m_bootloader.r_cstate[3] ;
 wire \m_sys.m_bootloader.r_cstate[4] ;
 wire \m_sys.m_bootloader.r_num[0] ;
 wire \m_sys.m_bootloader.r_num[1] ;
 wire \m_sys.m_bootloader.r_num[2] ;
 wire \m_sys.m_bootloader.r_num[3] ;
 wire \m_sys.m_bootloader.r_num[4] ;
 wire \m_sys.m_bootloader.r_num[5] ;
 wire \m_sys.m_bootloader.r_num[6] ;
 wire \m_sys.m_bootloader.r_num[7] ;
 wire \m_sys.m_bootloader.r_num_cnt[0] ;
 wire \m_sys.m_bootloader.r_num_cnt[1] ;
 wire \m_sys.m_bootloader.r_num_cnt[2] ;
 wire \m_sys.m_bootloader.r_num_cnt[3] ;
 wire \m_sys.m_bootloader.r_num_cnt[4] ;
 wire \m_sys.m_bootloader.r_num_cnt[5] ;
 wire \m_sys.m_bootloader.r_num_cnt[6] ;
 wire \m_sys.m_bootloader.r_num_cnt[7] ;
 wire \m_sys.m_bootloader.r_offset_0[0] ;
 wire \m_sys.m_bootloader.r_offset_0[1] ;
 wire \m_sys.m_bootloader.r_offset_0[2] ;
 wire \m_sys.m_bootloader.r_offset_0[3] ;
 wire \m_sys.m_bootloader.r_offset_0[4] ;
 wire \m_sys.m_bootloader.r_offset_0[5] ;
 wire \m_sys.m_bootloader.r_offset_0[6] ;
 wire \m_sys.m_bootloader.r_offset_0[7] ;
 wire \m_sys.m_bootloader.r_offset_1[0] ;
 wire \m_sys.m_bootloader.r_offset_1[1] ;
 wire \m_sys.m_bootloader.r_offset_1[2] ;
 wire \m_sys.m_bootloader.r_offset_1[3] ;
 wire \m_sys.m_bootloader.r_offset_1[4] ;
 wire \m_sys.m_bootloader.r_offset_1[5] ;
 wire \m_sys.m_bootloader.r_offset_1[6] ;
 wire \m_sys.m_bootloader.r_offset_1[7] ;
 wire \m_sys.m_core._m_bru_io_o_res[0] ;
 wire \m_sys.m_core._m_bru_io_o_res[1] ;
 wire \m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[0] ;
 wire \m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[1] ;
 wire \m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[2] ;
 wire \m_sys.m_core._m_decoder_io_o_rs1[0] ;
 wire \m_sys.m_core._m_decoder_io_o_rs1[1] ;
 wire \m_sys.m_core._m_decoder_io_o_rs1[2] ;
 wire \m_sys.m_core._m_decoder_io_o_rs2[0] ;
 wire \m_sys.m_core._m_decoder_io_o_rs2[1] ;
 wire \m_sys.m_core._m_decoder_io_o_rs2[2] ;
 wire \m_sys.m_core.m_alu.io_i_signed ;
 wire \m_sys.m_core.m_alu.io_i_uop[0] ;
 wire \m_sys.m_core.m_alu.io_i_uop[1] ;
 wire \m_sys.m_core.m_alu.io_i_uop[2] ;
 wire \m_sys.m_core.m_bru.io_i_pc[10] ;
 wire \m_sys.m_core.m_bru.io_i_pc[11] ;
 wire \m_sys.m_core.m_bru.io_i_pc[2] ;
 wire \m_sys.m_core.m_bru.io_i_pc[3] ;
 wire \m_sys.m_core.m_bru.io_i_pc[4] ;
 wire \m_sys.m_core.m_bru.io_i_pc[5] ;
 wire \m_sys.m_core.m_bru.io_i_pc[6] ;
 wire \m_sys.m_core.m_bru.io_i_pc[7] ;
 wire \m_sys.m_core.m_bru.io_i_pc[8] ;
 wire \m_sys.m_core.m_bru.io_i_pc[9] ;
 wire \m_sys.m_core.m_bru.io_i_s1[0] ;
 wire \m_sys.m_core.m_bru.io_i_s1[10] ;
 wire \m_sys.m_core.m_bru.io_i_s1[11] ;
 wire \m_sys.m_core.m_bru.io_i_s1[12] ;
 wire \m_sys.m_core.m_bru.io_i_s1[13] ;
 wire \m_sys.m_core.m_bru.io_i_s1[14] ;
 wire \m_sys.m_core.m_bru.io_i_s1[18] ;
 wire \m_sys.m_core.m_bru.io_i_s1[19] ;
 wire \m_sys.m_core.m_bru.io_i_s1[1] ;
 wire \m_sys.m_core.m_bru.io_i_s1[23] ;
 wire \m_sys.m_core.m_bru.io_i_s1[24] ;
 wire \m_sys.m_core.m_bru.io_i_s1[25] ;
 wire \m_sys.m_core.m_bru.io_i_s1[26] ;
 wire \m_sys.m_core.m_bru.io_i_s1[27] ;
 wire \m_sys.m_core.m_bru.io_i_s1[28] ;
 wire \m_sys.m_core.m_bru.io_i_s1[29] ;
 wire \m_sys.m_core.m_bru.io_i_s1[2] ;
 wire \m_sys.m_core.m_bru.io_i_s1[30] ;
 wire \m_sys.m_core.m_bru.io_i_s1[31] ;
 wire \m_sys.m_core.m_bru.io_i_s1[3] ;
 wire \m_sys.m_core.m_bru.io_i_s1[4] ;
 wire \m_sys.m_core.m_bru.io_i_s1[5] ;
 wire \m_sys.m_core.m_bru.io_i_s1[6] ;
 wire \m_sys.m_core.m_bru.io_i_s2[0] ;
 wire \m_sys.m_core.m_bru.io_i_s2[10] ;
 wire \m_sys.m_core.m_bru.io_i_s2[11] ;
 wire \m_sys.m_core.m_bru.io_i_s2[12] ;
 wire \m_sys.m_core.m_bru.io_i_s2[13] ;
 wire \m_sys.m_core.m_bru.io_i_s2[14] ;
 wire \m_sys.m_core.m_bru.io_i_s2[15] ;
 wire \m_sys.m_core.m_bru.io_i_s2[16] ;
 wire \m_sys.m_core.m_bru.io_i_s2[17] ;
 wire \m_sys.m_core.m_bru.io_i_s2[18] ;
 wire \m_sys.m_core.m_bru.io_i_s2[19] ;
 wire \m_sys.m_core.m_bru.io_i_s2[1] ;
 wire \m_sys.m_core.m_bru.io_i_s2[20] ;
 wire \m_sys.m_core.m_bru.io_i_s2[21] ;
 wire \m_sys.m_core.m_bru.io_i_s2[22] ;
 wire \m_sys.m_core.m_bru.io_i_s2[23] ;
 wire \m_sys.m_core.m_bru.io_i_s2[24] ;
 wire \m_sys.m_core.m_bru.io_i_s2[25] ;
 wire \m_sys.m_core.m_bru.io_i_s2[26] ;
 wire \m_sys.m_core.m_bru.io_i_s2[27] ;
 wire \m_sys.m_core.m_bru.io_i_s2[28] ;
 wire \m_sys.m_core.m_bru.io_i_s2[29] ;
 wire \m_sys.m_core.m_bru.io_i_s2[2] ;
 wire \m_sys.m_core.m_bru.io_i_s2[30] ;
 wire \m_sys.m_core.m_bru.io_i_s2[31] ;
 wire \m_sys.m_core.m_bru.io_i_s2[3] ;
 wire \m_sys.m_core.m_bru.io_i_s2[4] ;
 wire \m_sys.m_core.m_bru.io_i_s2[5] ;
 wire \m_sys.m_core.m_bru.io_i_s2[6] ;
 wire \m_sys.m_core.m_bru.io_i_s2[7] ;
 wire \m_sys.m_core.m_bru.io_i_s2[8] ;
 wire \m_sys.m_core.m_bru.io_i_s2[9] ;
 wire \m_sys.m_core.m_bru.io_i_uop[0] ;
 wire \m_sys.m_core.m_bru.io_i_uop[1] ;
 wire \m_sys.m_core.m_bru.io_i_uop[2] ;
 wire \m_sys.m_core.m_fsm.r_cstate[0] ;
 wire \m_sys.m_core.m_fsm.r_cstate[1] ;
 wire \m_sys.m_core.m_fsm.r_cstate[2] ;
 wire \m_sys.m_core.m_fsm.r_cstate[3] ;
 wire \m_sys.m_core.m_gpr._GEN[100] ;
 wire \m_sys.m_core.m_gpr._GEN[101] ;
 wire \m_sys.m_core.m_gpr._GEN[102] ;
 wire \m_sys.m_core.m_gpr._GEN[103] ;
 wire \m_sys.m_core.m_gpr._GEN[104] ;
 wire \m_sys.m_core.m_gpr._GEN[105] ;
 wire \m_sys.m_core.m_gpr._GEN[106] ;
 wire \m_sys.m_core.m_gpr._GEN[107] ;
 wire \m_sys.m_core.m_gpr._GEN[108] ;
 wire \m_sys.m_core.m_gpr._GEN[109] ;
 wire \m_sys.m_core.m_gpr._GEN[110] ;
 wire \m_sys.m_core.m_gpr._GEN[111] ;
 wire \m_sys.m_core.m_gpr._GEN[112] ;
 wire \m_sys.m_core.m_gpr._GEN[113] ;
 wire \m_sys.m_core.m_gpr._GEN[114] ;
 wire \m_sys.m_core.m_gpr._GEN[115] ;
 wire \m_sys.m_core.m_gpr._GEN[116] ;
 wire \m_sys.m_core.m_gpr._GEN[117] ;
 wire \m_sys.m_core.m_gpr._GEN[118] ;
 wire \m_sys.m_core.m_gpr._GEN[119] ;
 wire \m_sys.m_core.m_gpr._GEN[120] ;
 wire \m_sys.m_core.m_gpr._GEN[121] ;
 wire \m_sys.m_core.m_gpr._GEN[122] ;
 wire \m_sys.m_core.m_gpr._GEN[123] ;
 wire \m_sys.m_core.m_gpr._GEN[124] ;
 wire \m_sys.m_core.m_gpr._GEN[125] ;
 wire \m_sys.m_core.m_gpr._GEN[126] ;
 wire \m_sys.m_core.m_gpr._GEN[127] ;
 wire \m_sys.m_core.m_gpr._GEN[128] ;
 wire \m_sys.m_core.m_gpr._GEN[129] ;
 wire \m_sys.m_core.m_gpr._GEN[130] ;
 wire \m_sys.m_core.m_gpr._GEN[131] ;
 wire \m_sys.m_core.m_gpr._GEN[132] ;
 wire \m_sys.m_core.m_gpr._GEN[133] ;
 wire \m_sys.m_core.m_gpr._GEN[134] ;
 wire \m_sys.m_core.m_gpr._GEN[135] ;
 wire \m_sys.m_core.m_gpr._GEN[136] ;
 wire \m_sys.m_core.m_gpr._GEN[137] ;
 wire \m_sys.m_core.m_gpr._GEN[138] ;
 wire \m_sys.m_core.m_gpr._GEN[139] ;
 wire \m_sys.m_core.m_gpr._GEN[140] ;
 wire \m_sys.m_core.m_gpr._GEN[141] ;
 wire \m_sys.m_core.m_gpr._GEN[142] ;
 wire \m_sys.m_core.m_gpr._GEN[143] ;
 wire \m_sys.m_core.m_gpr._GEN[144] ;
 wire \m_sys.m_core.m_gpr._GEN[145] ;
 wire \m_sys.m_core.m_gpr._GEN[146] ;
 wire \m_sys.m_core.m_gpr._GEN[147] ;
 wire \m_sys.m_core.m_gpr._GEN[148] ;
 wire \m_sys.m_core.m_gpr._GEN[149] ;
 wire \m_sys.m_core.m_gpr._GEN[150] ;
 wire \m_sys.m_core.m_gpr._GEN[151] ;
 wire \m_sys.m_core.m_gpr._GEN[152] ;
 wire \m_sys.m_core.m_gpr._GEN[153] ;
 wire \m_sys.m_core.m_gpr._GEN[154] ;
 wire \m_sys.m_core.m_gpr._GEN[155] ;
 wire \m_sys.m_core.m_gpr._GEN[156] ;
 wire \m_sys.m_core.m_gpr._GEN[157] ;
 wire \m_sys.m_core.m_gpr._GEN[158] ;
 wire \m_sys.m_core.m_gpr._GEN[159] ;
 wire \m_sys.m_core.m_gpr._GEN[160] ;
 wire \m_sys.m_core.m_gpr._GEN[161] ;
 wire \m_sys.m_core.m_gpr._GEN[162] ;
 wire \m_sys.m_core.m_gpr._GEN[163] ;
 wire \m_sys.m_core.m_gpr._GEN[164] ;
 wire \m_sys.m_core.m_gpr._GEN[165] ;
 wire \m_sys.m_core.m_gpr._GEN[166] ;
 wire \m_sys.m_core.m_gpr._GEN[167] ;
 wire \m_sys.m_core.m_gpr._GEN[168] ;
 wire \m_sys.m_core.m_gpr._GEN[169] ;
 wire \m_sys.m_core.m_gpr._GEN[170] ;
 wire \m_sys.m_core.m_gpr._GEN[171] ;
 wire \m_sys.m_core.m_gpr._GEN[172] ;
 wire \m_sys.m_core.m_gpr._GEN[173] ;
 wire \m_sys.m_core.m_gpr._GEN[174] ;
 wire \m_sys.m_core.m_gpr._GEN[175] ;
 wire \m_sys.m_core.m_gpr._GEN[176] ;
 wire \m_sys.m_core.m_gpr._GEN[177] ;
 wire \m_sys.m_core.m_gpr._GEN[178] ;
 wire \m_sys.m_core.m_gpr._GEN[179] ;
 wire \m_sys.m_core.m_gpr._GEN[180] ;
 wire \m_sys.m_core.m_gpr._GEN[181] ;
 wire \m_sys.m_core.m_gpr._GEN[182] ;
 wire \m_sys.m_core.m_gpr._GEN[183] ;
 wire \m_sys.m_core.m_gpr._GEN[184] ;
 wire \m_sys.m_core.m_gpr._GEN[185] ;
 wire \m_sys.m_core.m_gpr._GEN[186] ;
 wire \m_sys.m_core.m_gpr._GEN[187] ;
 wire \m_sys.m_core.m_gpr._GEN[188] ;
 wire \m_sys.m_core.m_gpr._GEN[189] ;
 wire \m_sys.m_core.m_gpr._GEN[190] ;
 wire \m_sys.m_core.m_gpr._GEN[191] ;
 wire \m_sys.m_core.m_gpr._GEN[192] ;
 wire \m_sys.m_core.m_gpr._GEN[193] ;
 wire \m_sys.m_core.m_gpr._GEN[194] ;
 wire \m_sys.m_core.m_gpr._GEN[195] ;
 wire \m_sys.m_core.m_gpr._GEN[196] ;
 wire \m_sys.m_core.m_gpr._GEN[197] ;
 wire \m_sys.m_core.m_gpr._GEN[198] ;
 wire \m_sys.m_core.m_gpr._GEN[199] ;
 wire \m_sys.m_core.m_gpr._GEN[200] ;
 wire \m_sys.m_core.m_gpr._GEN[201] ;
 wire \m_sys.m_core.m_gpr._GEN[202] ;
 wire \m_sys.m_core.m_gpr._GEN[203] ;
 wire \m_sys.m_core.m_gpr._GEN[204] ;
 wire \m_sys.m_core.m_gpr._GEN[205] ;
 wire \m_sys.m_core.m_gpr._GEN[206] ;
 wire \m_sys.m_core.m_gpr._GEN[207] ;
 wire \m_sys.m_core.m_gpr._GEN[208] ;
 wire \m_sys.m_core.m_gpr._GEN[209] ;
 wire \m_sys.m_core.m_gpr._GEN[210] ;
 wire \m_sys.m_core.m_gpr._GEN[211] ;
 wire \m_sys.m_core.m_gpr._GEN[212] ;
 wire \m_sys.m_core.m_gpr._GEN[213] ;
 wire \m_sys.m_core.m_gpr._GEN[214] ;
 wire \m_sys.m_core.m_gpr._GEN[215] ;
 wire \m_sys.m_core.m_gpr._GEN[216] ;
 wire \m_sys.m_core.m_gpr._GEN[217] ;
 wire \m_sys.m_core.m_gpr._GEN[218] ;
 wire \m_sys.m_core.m_gpr._GEN[219] ;
 wire \m_sys.m_core.m_gpr._GEN[220] ;
 wire \m_sys.m_core.m_gpr._GEN[221] ;
 wire \m_sys.m_core.m_gpr._GEN[222] ;
 wire \m_sys.m_core.m_gpr._GEN[223] ;
 wire \m_sys.m_core.m_gpr._GEN[224] ;
 wire \m_sys.m_core.m_gpr._GEN[225] ;
 wire \m_sys.m_core.m_gpr._GEN[226] ;
 wire \m_sys.m_core.m_gpr._GEN[227] ;
 wire \m_sys.m_core.m_gpr._GEN[228] ;
 wire \m_sys.m_core.m_gpr._GEN[229] ;
 wire \m_sys.m_core.m_gpr._GEN[230] ;
 wire \m_sys.m_core.m_gpr._GEN[231] ;
 wire \m_sys.m_core.m_gpr._GEN[232] ;
 wire \m_sys.m_core.m_gpr._GEN[233] ;
 wire \m_sys.m_core.m_gpr._GEN[234] ;
 wire \m_sys.m_core.m_gpr._GEN[235] ;
 wire \m_sys.m_core.m_gpr._GEN[236] ;
 wire \m_sys.m_core.m_gpr._GEN[237] ;
 wire \m_sys.m_core.m_gpr._GEN[238] ;
 wire \m_sys.m_core.m_gpr._GEN[239] ;
 wire \m_sys.m_core.m_gpr._GEN[240] ;
 wire \m_sys.m_core.m_gpr._GEN[241] ;
 wire \m_sys.m_core.m_gpr._GEN[242] ;
 wire \m_sys.m_core.m_gpr._GEN[243] ;
 wire \m_sys.m_core.m_gpr._GEN[244] ;
 wire \m_sys.m_core.m_gpr._GEN[245] ;
 wire \m_sys.m_core.m_gpr._GEN[246] ;
 wire \m_sys.m_core.m_gpr._GEN[247] ;
 wire \m_sys.m_core.m_gpr._GEN[248] ;
 wire \m_sys.m_core.m_gpr._GEN[249] ;
 wire \m_sys.m_core.m_gpr._GEN[250] ;
 wire \m_sys.m_core.m_gpr._GEN[251] ;
 wire \m_sys.m_core.m_gpr._GEN[252] ;
 wire \m_sys.m_core.m_gpr._GEN[253] ;
 wire \m_sys.m_core.m_gpr._GEN[254] ;
 wire \m_sys.m_core.m_gpr._GEN[255] ;
 wire \m_sys.m_core.m_gpr._GEN[32] ;
 wire \m_sys.m_core.m_gpr._GEN[33] ;
 wire \m_sys.m_core.m_gpr._GEN[34] ;
 wire \m_sys.m_core.m_gpr._GEN[35] ;
 wire \m_sys.m_core.m_gpr._GEN[36] ;
 wire \m_sys.m_core.m_gpr._GEN[37] ;
 wire \m_sys.m_core.m_gpr._GEN[38] ;
 wire \m_sys.m_core.m_gpr._GEN[39] ;
 wire \m_sys.m_core.m_gpr._GEN[40] ;
 wire \m_sys.m_core.m_gpr._GEN[41] ;
 wire \m_sys.m_core.m_gpr._GEN[42] ;
 wire \m_sys.m_core.m_gpr._GEN[43] ;
 wire \m_sys.m_core.m_gpr._GEN[44] ;
 wire \m_sys.m_core.m_gpr._GEN[45] ;
 wire \m_sys.m_core.m_gpr._GEN[46] ;
 wire \m_sys.m_core.m_gpr._GEN[47] ;
 wire \m_sys.m_core.m_gpr._GEN[48] ;
 wire \m_sys.m_core.m_gpr._GEN[49] ;
 wire \m_sys.m_core.m_gpr._GEN[50] ;
 wire \m_sys.m_core.m_gpr._GEN[51] ;
 wire \m_sys.m_core.m_gpr._GEN[52] ;
 wire \m_sys.m_core.m_gpr._GEN[53] ;
 wire \m_sys.m_core.m_gpr._GEN[54] ;
 wire \m_sys.m_core.m_gpr._GEN[55] ;
 wire \m_sys.m_core.m_gpr._GEN[56] ;
 wire \m_sys.m_core.m_gpr._GEN[57] ;
 wire \m_sys.m_core.m_gpr._GEN[58] ;
 wire \m_sys.m_core.m_gpr._GEN[59] ;
 wire \m_sys.m_core.m_gpr._GEN[60] ;
 wire \m_sys.m_core.m_gpr._GEN[61] ;
 wire \m_sys.m_core.m_gpr._GEN[62] ;
 wire \m_sys.m_core.m_gpr._GEN[63] ;
 wire \m_sys.m_core.m_gpr._GEN[64] ;
 wire \m_sys.m_core.m_gpr._GEN[65] ;
 wire \m_sys.m_core.m_gpr._GEN[66] ;
 wire \m_sys.m_core.m_gpr._GEN[67] ;
 wire \m_sys.m_core.m_gpr._GEN[68] ;
 wire \m_sys.m_core.m_gpr._GEN[69] ;
 wire \m_sys.m_core.m_gpr._GEN[70] ;
 wire \m_sys.m_core.m_gpr._GEN[71] ;
 wire \m_sys.m_core.m_gpr._GEN[72] ;
 wire \m_sys.m_core.m_gpr._GEN[73] ;
 wire \m_sys.m_core.m_gpr._GEN[74] ;
 wire \m_sys.m_core.m_gpr._GEN[75] ;
 wire \m_sys.m_core.m_gpr._GEN[76] ;
 wire \m_sys.m_core.m_gpr._GEN[77] ;
 wire \m_sys.m_core.m_gpr._GEN[78] ;
 wire \m_sys.m_core.m_gpr._GEN[79] ;
 wire \m_sys.m_core.m_gpr._GEN[80] ;
 wire \m_sys.m_core.m_gpr._GEN[81] ;
 wire \m_sys.m_core.m_gpr._GEN[82] ;
 wire \m_sys.m_core.m_gpr._GEN[83] ;
 wire \m_sys.m_core.m_gpr._GEN[84] ;
 wire \m_sys.m_core.m_gpr._GEN[85] ;
 wire \m_sys.m_core.m_gpr._GEN[86] ;
 wire \m_sys.m_core.m_gpr._GEN[87] ;
 wire \m_sys.m_core.m_gpr._GEN[88] ;
 wire \m_sys.m_core.m_gpr._GEN[89] ;
 wire \m_sys.m_core.m_gpr._GEN[90] ;
 wire \m_sys.m_core.m_gpr._GEN[91] ;
 wire \m_sys.m_core.m_gpr._GEN[92] ;
 wire \m_sys.m_core.m_gpr._GEN[93] ;
 wire \m_sys.m_core.m_gpr._GEN[94] ;
 wire \m_sys.m_core.m_gpr._GEN[95] ;
 wire \m_sys.m_core.m_gpr._GEN[96] ;
 wire \m_sys.m_core.m_gpr._GEN[97] ;
 wire \m_sys.m_core.m_gpr._GEN[98] ;
 wire \m_sys.m_core.m_gpr._GEN[99] ;
 wire \m_sys.m_core.m_gpr.io_b_write_addr[0] ;
 wire \m_sys.m_core.m_gpr.io_b_write_addr[1] ;
 wire \m_sys.m_core.m_gpr.io_b_write_addr[2] ;
 wire \m_sys.m_core.r_ctrl_bru_pc_rel ;
 wire \m_sys.m_core.r_ctrl_mem_rw ;
 wire \m_sys.m_core.r_ctrl_mem_signed ;
 wire \m_sys.m_core.r_ctrl_mem_size[0] ;
 wire \m_sys.m_core.r_ctrl_mem_size[1] ;
 wire \m_sys.m_core.r_ctrl_wb_en ;
 wire \m_sys.m_gpio8.r_in[0] ;
 wire \m_sys.m_gpio8.r_in[1] ;
 wire \m_sys.m_gpio8.r_in[2] ;
 wire \m_sys.m_gpio8.r_in[3] ;
 wire \m_sys.m_gpio8.r_in[4] ;
 wire \m_sys.m_gpio8.r_in[5] ;
 wire \m_sys.m_gpio8.r_in[6] ;
 wire \m_sys.m_gpio8.r_in[7] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[0][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[10][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[11][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[12][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[13][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[14][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[15][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[16][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[17][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[18][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[19][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[1][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[20][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[21][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[22][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[23][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[24][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[25][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[26][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[27][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[28][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[29][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[2][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[30][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[31][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[3][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[4][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[5][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[6][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[7][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[8][9] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][0] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][10] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][11] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][12] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][13] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][14] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][15] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][16] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][17] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][18] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][19] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][1] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][20] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][21] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][22] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][23] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][24] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][25] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][26] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][27] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][28] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][29] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][2] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][30] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][31] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][3] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][4] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][5] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][6] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][7] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][8] ;
 wire \m_sys.m_ram.m_ram.r_mem[9][9] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[0] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[10] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[11] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[12] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[13] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[14] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[15] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[1] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[2] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[3] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[4] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[5] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[6] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[7] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[8] ;
 wire \m_sys.m_uart.m_rx.io_i_ncycle[9] ;
 wire \m_sys.m_uart.m_rx.r_bit_cnt[0] ;
 wire \m_sys.m_uart.m_rx.r_bit_cnt[1] ;
 wire \m_sys.m_uart.m_rx.r_bit_cnt[2] ;
 wire \m_sys.m_uart.m_rx.r_cstate[0] ;
 wire \m_sys.m_uart.m_rx.r_cstate[1] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[0] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[10] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[11] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[12] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[13] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[14] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[15] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[1] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[2] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[3] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[4] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[5] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[6] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[7] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[8] ;
 wire \m_sys.m_uart.m_rx.r_cycle_cnt[9] ;
 wire \m_sys.m_uart.m_rx.r_rx ;
 wire \m_sys.m_uart.m_tx.r_bit_cnt[0] ;
 wire \m_sys.m_uart.m_tx.r_bit_cnt[1] ;
 wire \m_sys.m_uart.m_tx.r_bit_cnt[2] ;
 wire \m_sys.m_uart.m_tx.r_cstate[0] ;
 wire \m_sys.m_uart.m_tx.r_cstate[1] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[0] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[10] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[11] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[12] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[13] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[14] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[15] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[1] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[2] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[3] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[4] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[5] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[6] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[7] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[8] ;
 wire \m_sys.m_uart.m_tx.r_cycle_cnt[9] ;
 wire \m_sys.m_uart.m_tx.r_data[0] ;
 wire \m_sys.m_uart.m_tx.r_data[1] ;
 wire \m_sys.m_uart.m_tx.r_data[2] ;
 wire \m_sys.m_uart.m_tx.r_data[3] ;
 wire \m_sys.m_uart.m_tx.r_data[4] ;
 wire \m_sys.m_uart.m_tx.r_data[5] ;
 wire \m_sys.m_uart.m_tx.r_data[6] ;
 wire \m_sys.m_uart.m_tx.r_data[7] ;
 wire \m_sys.m_uart.r_rx_data[0] ;
 wire \m_sys.m_uart.r_rx_data[1] ;
 wire \m_sys.m_uart.r_rx_data[2] ;
 wire \m_sys.m_uart.r_rx_data[3] ;
 wire \m_sys.m_uart.r_rx_data[4] ;
 wire \m_sys.m_uart.r_rx_data[5] ;
 wire \m_sys.m_uart.r_rx_data[6] ;
 wire \m_sys.m_uart.r_rx_data[7] ;
 wire \m_sys.m_uart.r_rx_valid ;
 wire \m_sys.r_addr[10] ;
 wire \m_sys.r_addr[11] ;
 wire \m_sys.r_addr[6] ;
 wire \m_sys.r_addr[7] ;
 wire \m_sys.r_addr[8] ;
 wire \m_sys.r_addr[9] ;
 wire \m_sys.r_valid ;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;

 sg13g2_inv_1 _10778_ (.Y(_02323_),
    .A(\m_sys.m_core._m_bru_io_o_res[1] ));
 sg13g2_inv_1 _10779_ (.Y(_02324_),
    .A(\m_sys.m_core._m_bru_io_o_res[0] ));
 sg13g2_inv_1 _10780_ (.Y(_02325_),
    .A(net3306));
 sg13g2_inv_1 _10781_ (.Y(_02326_),
    .A(net3374));
 sg13g2_inv_1 _10782_ (.Y(_02327_),
    .A(net3390));
 sg13g2_inv_1 _10783_ (.Y(_02328_),
    .A(net3225));
 sg13g2_inv_1 _10784_ (.Y(_02329_),
    .A(net3391));
 sg13g2_inv_1 _10785_ (.Y(_02330_),
    .A(net3383));
 sg13g2_inv_1 _10786_ (.Y(_02331_),
    .A(net3409));
 sg13g2_inv_1 _10787_ (.Y(_02332_),
    .A(net3397));
 sg13g2_inv_1 _10788_ (.Y(_02333_),
    .A(net3386));
 sg13g2_inv_1 _10789_ (.Y(_02334_),
    .A(net3419));
 sg13g2_inv_1 _10790_ (.Y(_02335_),
    .A(net3426));
 sg13g2_inv_1 _10791_ (.Y(_02336_),
    .A(net3373));
 sg13g2_inv_1 _10792_ (.Y(_02337_),
    .A(net3439));
 sg13g2_inv_1 _10793_ (.Y(_02338_),
    .A(net3435));
 sg13g2_inv_1 _10794_ (.Y(_02339_),
    .A(net3438));
 sg13g2_inv_1 _10795_ (.Y(_02340_),
    .A(net3434));
 sg13g2_inv_4 _10796_ (.A(net2522),
    .Y(_02341_));
 sg13g2_inv_4 _10797_ (.A(net3443),
    .Y(_02342_));
 sg13g2_inv_1 _10798_ (.Y(_02343_),
    .A(net2828));
 sg13g2_inv_1 _10799_ (.Y(_02344_),
    .A(net3053));
 sg13g2_inv_1 _10800_ (.Y(_02345_),
    .A(net3216));
 sg13g2_inv_2 _10801_ (.Y(_02346_),
    .A(net3090));
 sg13g2_inv_1 _10802_ (.Y(_02347_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[12] ));
 sg13g2_inv_1 _10803_ (.Y(_02348_),
    .A(net3201));
 sg13g2_inv_1 _10804_ (.Y(_02349_),
    .A(net3109));
 sg13g2_inv_1 _10805_ (.Y(_02350_),
    .A(net2952));
 sg13g2_inv_1 _10806_ (.Y(_02351_),
    .A(net3368));
 sg13g2_inv_1 _10807_ (.Y(_02352_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[6] ));
 sg13g2_inv_1 _10808_ (.Y(_02353_),
    .A(net3358));
 sg13g2_inv_2 _10809_ (.Y(_02354_),
    .A(net3152));
 sg13g2_inv_1 _10810_ (.Y(_02355_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[3] ));
 sg13g2_inv_1 _10811_ (.Y(_02356_),
    .A(net3422));
 sg13g2_inv_1 _10812_ (.Y(_02357_),
    .A(net3356));
 sg13g2_inv_1 _10813_ (.Y(_02358_),
    .A(net3416));
 sg13g2_inv_1 _10814_ (.Y(_02359_),
    .A(net2985));
 sg13g2_inv_1 _10815_ (.Y(_02360_),
    .A(net5282));
 sg13g2_inv_2 _10816_ (.Y(_02361_),
    .A(net5286));
 sg13g2_inv_1 _10817_ (.Y(_02362_),
    .A(net3385));
 sg13g2_inv_1 _10818_ (.Y(_02363_),
    .A(net3366));
 sg13g2_inv_1 _10819_ (.Y(_02364_),
    .A(net2903));
 sg13g2_inv_2 _10820_ (.Y(_02365_),
    .A(net3125));
 sg13g2_inv_2 _10821_ (.Y(_02366_),
    .A(net5271));
 sg13g2_inv_1 _10822_ (.Y(_02367_),
    .A(net5267));
 sg13g2_inv_2 _10823_ (.Y(_02368_),
    .A(net5242));
 sg13g2_inv_1 _10824_ (.Y(_02369_),
    .A(net5309));
 sg13g2_inv_1 _10825_ (.Y(_02370_),
    .A(\m_sys._m_bootloader_io_b_mem_addr[4] ));
 sg13g2_inv_4 _10826_ (.A(\m_sys.m_core.m_bru.io_i_s1[2] ),
    .Y(_02371_));
 sg13g2_inv_2 _10827_ (.Y(_02372_),
    .A(net3415));
 sg13g2_inv_1 _10828_ (.Y(_02373_),
    .A(net3387));
 sg13g2_inv_1 _10829_ (.Y(_02374_),
    .A(_00013_));
 sg13g2_inv_1 _10830_ (.Y(_02375_),
    .A(\m_sys.m_uart.m_tx.r_cycle_cnt[2] ));
 sg13g2_inv_1 _10831_ (.Y(_02376_),
    .A(\m_sys.m_uart.m_tx.r_cycle_cnt[9] ));
 sg13g2_inv_1 _10832_ (.Y(_02377_),
    .A(\m_sys.m_uart.m_tx.r_cycle_cnt[10] ));
 sg13g2_inv_1 _10833_ (.Y(_02378_),
    .A(\m_sys.m_uart.m_tx.r_cycle_cnt[11] ));
 sg13g2_inv_1 _10834_ (.Y(_02379_),
    .A(\m_sys.m_uart.m_tx.r_cycle_cnt[12] ));
 sg13g2_inv_1 _10835_ (.Y(_02380_),
    .A(\m_sys.m_uart.m_tx.r_cycle_cnt[13] ));
 sg13g2_inv_4 _10836_ (.A(\m_sys.m_core.m_bru.io_i_s1[11] ),
    .Y(_02381_));
 sg13g2_inv_1 _10837_ (.Y(_02382_),
    .A(_00016_));
 sg13g2_inv_4 _10838_ (.A(\m_sys.m_core.m_bru.io_i_s1[10] ),
    .Y(_02383_));
 sg13g2_inv_1 _10839_ (.Y(_02384_),
    .A(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[2] ));
 sg13g2_inv_1 _10840_ (.Y(_02385_),
    .A(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[0] ));
 sg13g2_inv_1 _10841_ (.Y(_02386_),
    .A(\m_sys.m_core.m_bru.io_i_s1[6] ));
 sg13g2_inv_1 _10842_ (.Y(_02387_),
    .A(\m_sys._m_bootloader_io_b_mem_addr[11] ));
 sg13g2_inv_1 _10843_ (.Y(_02388_),
    .A(net3421));
 sg13g2_inv_1 _10844_ (.Y(_02389_),
    .A(net3037));
 sg13g2_inv_1 _10845_ (.Y(_02390_),
    .A(\m_sys.m_uart.m_rx.r_cycle_cnt[2] ));
 sg13g2_inv_1 _10846_ (.Y(_02391_),
    .A(\m_sys.m_uart.m_rx.r_cycle_cnt[3] ));
 sg13g2_inv_1 _10847_ (.Y(_02392_),
    .A(\m_sys.m_uart.m_rx.r_cycle_cnt[4] ));
 sg13g2_inv_1 _10848_ (.Y(_02393_),
    .A(\m_sys.m_uart.m_rx.r_cycle_cnt[8] ));
 sg13g2_inv_1 _10849_ (.Y(_02394_),
    .A(\m_sys.m_uart.m_rx.r_cycle_cnt[13] ));
 sg13g2_inv_1 _10850_ (.Y(_02395_),
    .A(\m_sys.m_uart.m_rx.r_cycle_cnt[14] ));
 sg13g2_inv_1 _10851_ (.Y(_02396_),
    .A(net5382));
 sg13g2_inv_4 _10852_ (.A(\m_sys.m_core.m_bru.io_i_s1[0] ),
    .Y(_02397_));
 sg13g2_inv_2 _10853_ (.Y(_02398_),
    .A(\m_sys.m_core.m_bru.io_i_s1[13] ));
 sg13g2_inv_4 _10854_ (.A(\m_sys.m_core.m_bru.io_i_s1[12] ),
    .Y(_02399_));
 sg13g2_inv_4 _10855_ (.A(\m_sys.m_core.m_bru.io_i_s1[14] ),
    .Y(_02400_));
 sg13g2_inv_1 _10856_ (.Y(_02401_),
    .A(\m_sys.m_bootloader.r_byte_cnt[0] ));
 sg13g2_inv_1 _10857_ (.Y(_02402_),
    .A(net5311));
 sg13g2_inv_1 _10858_ (.Y(_02403_),
    .A(_00033_));
 sg13g2_inv_1 _10859_ (.Y(_02404_),
    .A(net3315));
 sg13g2_inv_1 _10860_ (.Y(_02405_),
    .A(net3272));
 sg13g2_inv_1 _10861_ (.Y(_02406_),
    .A(net3323));
 sg13g2_inv_1 _10862_ (.Y(_02407_),
    .A(net3189));
 sg13g2_inv_1 _10863_ (.Y(_02408_),
    .A(\m_sys._m_core_io_b_mem_wdata[9] ));
 sg13g2_inv_1 _10864_ (.Y(_02409_),
    .A(\m_sys._m_core_io_b_mem_wdata[10] ));
 sg13g2_inv_1 _10865_ (.Y(_02410_),
    .A(\m_sys._m_core_io_b_mem_wdata[11] ));
 sg13g2_inv_2 _10866_ (.Y(_02411_),
    .A(net5278));
 sg13g2_inv_1 _10867_ (.Y(_02412_),
    .A(net3142));
 sg13g2_inv_1 _10868_ (.Y(_02413_),
    .A(net3164));
 sg13g2_inv_1 _10869_ (.Y(_02414_),
    .A(net3351));
 sg13g2_inv_1 _10870_ (.Y(_02415_),
    .A(net3234));
 sg13g2_inv_1 _10871_ (.Y(_02416_),
    .A(net3114));
 sg13g2_inv_1 _10872_ (.Y(_02417_),
    .A(\m_sys._m_uart_io_b_mem_rdata[7] ));
 sg13g2_inv_1 _10873_ (.Y(_02418_),
    .A(\m_sys._m_gpio8_io_b_mem_rdata[7] ));
 sg13g2_inv_1 _10874_ (.Y(_02419_),
    .A(_00062_));
 sg13g2_inv_1 _10875_ (.Y(_02420_),
    .A(_00063_));
 sg13g2_inv_1 _10876_ (.Y(_02421_),
    .A(net2590));
 sg13g2_inv_1 _10877_ (.Y(_02422_),
    .A(net5349));
 sg13g2_inv_1 _10878_ (.Y(_02423_),
    .A(net5351));
 sg13g2_inv_1 _10879_ (.Y(_02424_),
    .A(net5340));
 sg13g2_inv_1 _10880_ (.Y(_02425_),
    .A(net2511));
 sg13g2_inv_1 _10881_ (.Y(_02426_),
    .A(net3436));
 sg13g2_inv_2 _10882_ (.Y(_02427_),
    .A(\m_sys.m_core.m_bru.io_i_s1[23] ));
 sg13g2_inv_1 _10883_ (.Y(_02428_),
    .A(\m_sys.m_core.m_gpr._GEN[163] ));
 sg13g2_inv_1 _10884_ (.Y(_02429_),
    .A(net2986));
 sg13g2_inv_2 _10885_ (.Y(_02430_),
    .A(\m_sys.m_core.m_bru.io_i_s1[24] ));
 sg13g2_inv_1 _10886_ (.Y(_02431_),
    .A(net2510));
 sg13g2_inv_2 _10887_ (.Y(_02432_),
    .A(\m_sys.m_core.m_bru.io_i_s1[25] ));
 sg13g2_inv_1 _10888_ (.Y(_02433_),
    .A(net2802));
 sg13g2_inv_1 _10889_ (.Y(_02434_),
    .A(\m_sys.m_core.m_bru.io_i_s1[26] ));
 sg13g2_inv_1 _10890_ (.Y(_02435_),
    .A(\m_sys.m_core.m_gpr._GEN[102] ));
 sg13g2_inv_1 _10891_ (.Y(_02436_),
    .A(net2795));
 sg13g2_inv_1 _10892_ (.Y(_02437_),
    .A(\m_sys.m_core.m_bru.io_i_s1[27] ));
 sg13g2_inv_1 _10893_ (.Y(_02438_),
    .A(net2868));
 sg13g2_inv_4 _10894_ (.A(net3441),
    .Y(_02439_));
 sg13g2_inv_2 _10895_ (.Y(_02440_),
    .A(\m_sys.m_core.m_bru.io_i_s1[29] ));
 sg13g2_inv_1 _10896_ (.Y(_02441_),
    .A(net2918));
 sg13g2_inv_1 _10897_ (.Y(_02442_),
    .A(\m_sys.m_core.m_gpr._GEN[233] ));
 sg13g2_inv_4 _10898_ (.A(\m_sys.m_core.m_bru.io_i_s1[30] ),
    .Y(_02443_));
 sg13g2_inv_2 _10899_ (.Y(_02444_),
    .A(net3363));
 sg13g2_inv_2 _10900_ (.Y(_02445_),
    .A(\m_sys.m_core._m_decoder_io_o_rs1[0] ));
 sg13g2_inv_1 _10901_ (.Y(_02446_),
    .A(_00082_));
 sg13g2_inv_1 _10902_ (.Y(_02447_),
    .A(net5325));
 sg13g2_inv_2 _10903_ (.Y(_02448_),
    .A(net5330));
 sg13g2_inv_1 _10904_ (.Y(_02449_),
    .A(_00084_));
 sg13g2_inv_2 _10905_ (.Y(_02450_),
    .A(\m_sys.m_core.m_bru.io_i_s1[18] ));
 sg13g2_inv_1 _10906_ (.Y(_02451_),
    .A(_00085_));
 sg13g2_inv_2 _10907_ (.Y(_02452_),
    .A(\m_sys.m_core.m_bru.io_i_s1[19] ));
 sg13g2_inv_1 _10908_ (.Y(_02453_),
    .A(net2844));
 sg13g2_inv_1 _10909_ (.Y(_02454_),
    .A(net2827));
 sg13g2_inv_1 _10910_ (.Y(_02455_),
    .A(net2825));
 sg13g2_inv_1 _10911_ (.Y(_02456_),
    .A(net2749));
 sg13g2_inv_1 _10912_ (.Y(_02457_),
    .A(net2721));
 sg13g2_inv_1 _10913_ (.Y(_02458_),
    .A(net3179));
 sg13g2_inv_1 _10914_ (.Y(_02459_),
    .A(net3066));
 sg13g2_inv_1 _10915_ (.Y(_02460_),
    .A(net3243));
 sg13g2_inv_1 _10916_ (.Y(_02461_),
    .A(\m_sys.m_core.m_bru.io_i_s2[1] ));
 sg13g2_inv_1 _10917_ (.Y(_02462_),
    .A(net3382));
 sg13g2_inv_1 _10918_ (.Y(_02463_),
    .A(net3348));
 sg13g2_inv_1 _10919_ (.Y(_02464_),
    .A(net3233));
 sg13g2_inv_1 _10920_ (.Y(_02465_),
    .A(net3251));
 sg13g2_inv_1 _10921_ (.Y(_02466_),
    .A(net3298));
 sg13g2_inv_1 _10922_ (.Y(_02467_),
    .A(net3347));
 sg13g2_inv_1 _10923_ (.Y(_02468_),
    .A(\m_sys.m_core.m_bru.io_i_s2[14] ));
 sg13g2_inv_1 _10924_ (.Y(_02469_),
    .A(net3253));
 sg13g2_inv_1 _10925_ (.Y(_02470_),
    .A(net3388));
 sg13g2_inv_1 _10926_ (.Y(_02471_),
    .A(net3261));
 sg13g2_inv_1 _10927_ (.Y(_02472_),
    .A(net3019));
 sg13g2_inv_1 _10928_ (.Y(_02473_),
    .A(\m_sys.m_core.m_bru.io_i_s2[9] ));
 sg13g2_inv_1 _10929_ (.Y(_02474_),
    .A(net3296));
 sg13g2_inv_1 _10930_ (.Y(_02475_),
    .A(net3279));
 sg13g2_inv_1 _10931_ (.Y(_02476_),
    .A(net3231));
 sg13g2_inv_1 _10932_ (.Y(_02477_),
    .A(\m_sys.m_core.m_bru.io_i_s2[28] ));
 sg13g2_inv_1 _10933_ (.Y(_02478_),
    .A(net3372));
 sg13g2_inv_1 _10934_ (.Y(_02479_),
    .A(\m_sys.m_core.m_bru.io_i_s2[26] ));
 sg13g2_inv_2 _10935_ (.Y(_02480_),
    .A(net3393));
 sg13g2_inv_1 _10936_ (.Y(_02481_),
    .A(net3310));
 sg13g2_inv_1 _10937_ (.Y(_02482_),
    .A(\m_sys.m_core.m_bru.io_i_s2[22] ));
 sg13g2_inv_1 _10938_ (.Y(_02483_),
    .A(net3316));
 sg13g2_inv_1 _10939_ (.Y(_02484_),
    .A(net3328));
 sg13g2_inv_1 _10940_ (.Y(_02485_),
    .A(\m_sys.m_core.m_gpr._GEN[160] ));
 sg13g2_inv_1 _10941_ (.Y(_02486_),
    .A(net3131));
 sg13g2_inv_1 _10942_ (.Y(_02487_),
    .A(net5288));
 sg13g2_inv_1 _10943_ (.Y(_02488_),
    .A(net3080));
 sg13g2_inv_2 _10944_ (.Y(_02489_),
    .A(net5251));
 sg13g2_inv_1 _10945_ (.Y(_02490_),
    .A(net5302));
 sg13g2_inv_1 _10946_ (.Y(_02491_),
    .A(_00093_));
 sg13g2_inv_1 _10947_ (.Y(_02492_),
    .A(_00096_));
 sg13g2_inv_1 _10948_ (.Y(_02493_),
    .A(_00101_));
 sg13g2_inv_1 _10949_ (.Y(_02494_),
    .A(_00107_));
 sg13g2_inv_1 _10950_ (.Y(_02495_),
    .A(_00118_));
 sg13g2_inv_1 _10951_ (.Y(_02496_),
    .A(net5257));
 sg13g2_inv_1 _10952_ (.Y(_02497_),
    .A(_00124_));
 sg13g2_inv_1 _10953_ (.Y(_02498_),
    .A(_00126_));
 sg13g2_inv_1 _10954_ (.Y(_02499_),
    .A(_00128_));
 sg13g2_inv_1 _10955_ (.Y(_02500_),
    .A(_00132_));
 sg13g2_inv_1 _10956_ (.Y(_02501_),
    .A(net3071));
 sg13g2_inv_1 _10957_ (.Y(_02502_),
    .A(_00139_));
 sg13g2_inv_1 _10958_ (.Y(_02503_),
    .A(net2964));
 sg13g2_nand2b_1 _10959_ (.Y(_02504_),
    .B(\m_sys.m_uart.m_tx.r_cycle_cnt[10] ),
    .A_N(\m_sys.m_uart.m_rx.io_i_ncycle[10] ));
 sg13g2_nand2b_1 _10960_ (.Y(_02505_),
    .B(\m_sys.m_uart.m_rx.io_i_ncycle[0] ),
    .A_N(\m_sys.m_uart.m_tx.r_cycle_cnt[0] ));
 sg13g2_nand2b_1 _10961_ (.Y(_02506_),
    .B(\m_sys.m_uart.m_rx.io_i_ncycle[6] ),
    .A_N(\m_sys.m_uart.m_tx.r_cycle_cnt[6] ));
 sg13g2_xnor2_1 _10962_ (.Y(_02507_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[8] ),
    .B(\m_sys.m_uart.m_tx.r_cycle_cnt[8] ));
 sg13g2_xnor2_1 _10963_ (.Y(_02508_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[5] ),
    .B(\m_sys.m_uart.m_tx.r_cycle_cnt[5] ));
 sg13g2_xnor2_1 _10964_ (.Y(_02509_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[1] ),
    .B(\m_sys.m_uart.m_tx.r_cycle_cnt[1] ));
 sg13g2_a22oi_1 _10965_ (.Y(_02510_),
    .B1(_02380_),
    .B2(\m_sys.m_uart.m_rx.io_i_ncycle[13] ),
    .A2(_02376_),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[9] ));
 sg13g2_xnor2_1 _10966_ (.Y(_02511_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[14] ),
    .B(\m_sys.m_uart.m_tx.r_cycle_cnt[14] ));
 sg13g2_a22oi_1 _10967_ (.Y(_02512_),
    .B1(_02377_),
    .B2(\m_sys.m_uart.m_rx.io_i_ncycle[10] ),
    .A2(\m_sys.m_uart.m_tx.r_cycle_cnt[2] ),
    .A1(_02356_));
 sg13g2_o21ai_1 _10968_ (.B1(_02505_),
    .Y(_02513_),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[9] ),
    .A2(_02376_));
 sg13g2_a22oi_1 _10969_ (.Y(_02514_),
    .B1(\m_sys.m_uart.m_tx.r_cycle_cnt[13] ),
    .B2(_02346_),
    .A2(\m_sys.m_uart.m_tx.r_cycle_cnt[6] ),
    .A1(_02352_));
 sg13g2_nand4_1 _10970_ (.B(_02506_),
    .C(_02509_),
    .A(_02504_),
    .Y(_02515_),
    .D(_02514_));
 sg13g2_a22oi_1 _10971_ (.Y(_02516_),
    .B1(\m_sys.m_uart.m_tx.r_cycle_cnt[12] ),
    .B2(_02347_),
    .A2(\m_sys.m_uart.m_tx.r_cycle_cnt[0] ),
    .A1(_02358_));
 sg13g2_nand4_1 _10972_ (.B(_02511_),
    .C(_02512_),
    .A(_02510_),
    .Y(_02517_),
    .D(_02516_));
 sg13g2_xor2_1 _10973_ (.B(\m_sys.m_uart.m_tx.r_cycle_cnt[3] ),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[3] ),
    .X(_02518_));
 sg13g2_a221oi_1 _10974_ (.B2(\m_sys.m_uart.m_rx.io_i_ncycle[12] ),
    .C1(_02518_),
    .B1(_02379_),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[11] ),
    .Y(_02519_),
    .A2(_02378_));
 sg13g2_a22oi_1 _10975_ (.Y(_02520_),
    .B1(\m_sys.m_uart.m_tx.r_cycle_cnt[11] ),
    .B2(_02348_),
    .A2(_02375_),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[2] ));
 sg13g2_xnor2_1 _10976_ (.Y(_02521_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[15] ),
    .B(\m_sys.m_uart.m_tx.r_cycle_cnt[15] ));
 sg13g2_xnor2_1 _10977_ (.Y(_02522_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[7] ),
    .B(\m_sys.m_uart.m_tx.r_cycle_cnt[7] ));
 sg13g2_xnor2_1 _10978_ (.Y(_02523_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[4] ),
    .B(\m_sys.m_uart.m_tx.r_cycle_cnt[4] ));
 sg13g2_nand4_1 _10979_ (.B(_02521_),
    .C(_02522_),
    .A(_02508_),
    .Y(_02524_),
    .D(_02523_));
 sg13g2_nor4_1 _10980_ (.A(_02513_),
    .B(_02515_),
    .C(_02517_),
    .D(_02524_),
    .Y(_02525_));
 sg13g2_nand4_1 _10981_ (.B(_02519_),
    .C(_02520_),
    .A(_02507_),
    .Y(_02526_),
    .D(_02525_));
 sg13g2_nand2b_2 _10982_ (.Y(_02527_),
    .B(_00014_),
    .A_N(\m_sys.m_uart.m_tx.r_cstate[1] ));
 sg13g2_nand2_1 _10983_ (.Y(_02528_),
    .A(_02526_),
    .B(_02527_));
 sg13g2_nor2_1 _10984_ (.A(net3095),
    .B(net4692),
    .Y(_01760_));
 sg13g2_xnor2_1 _10985_ (.Y(_02529_),
    .A(net3095),
    .B(net3230));
 sg13g2_nor2_1 _10986_ (.A(net4692),
    .B(_02529_),
    .Y(_01767_));
 sg13g2_and3_1 _10987_ (.X(_02530_),
    .A(net3095),
    .B(\m_sys.m_uart.m_tx.r_cycle_cnt[1] ),
    .C(net2911));
 sg13g2_a21oi_1 _10988_ (.A1(\m_sys.m_uart.m_tx.r_cycle_cnt[0] ),
    .A2(\m_sys.m_uart.m_tx.r_cycle_cnt[1] ),
    .Y(_02531_),
    .B1(net2911));
 sg13g2_nor3_1 _10989_ (.A(net4692),
    .B(_02530_),
    .C(net2912),
    .Y(_01768_));
 sg13g2_nor2_1 _10990_ (.A(net3204),
    .B(_02530_),
    .Y(_02532_));
 sg13g2_and2_1 _10991_ (.A(net3204),
    .B(_02530_),
    .X(_02533_));
 sg13g2_nor3_1 _10992_ (.A(net4691),
    .B(net3205),
    .C(_02533_),
    .Y(_01769_));
 sg13g2_nor2_1 _10993_ (.A(net3168),
    .B(_02533_),
    .Y(_02534_));
 sg13g2_and2_1 _10994_ (.A(net3168),
    .B(_02533_),
    .X(_02535_));
 sg13g2_nor3_1 _10995_ (.A(net4691),
    .B(net3169),
    .C(_02535_),
    .Y(_01770_));
 sg13g2_xnor2_1 _10996_ (.Y(_02536_),
    .A(net3307),
    .B(_02535_));
 sg13g2_nor2_1 _10997_ (.A(net4691),
    .B(_02536_),
    .Y(_01771_));
 sg13g2_a21oi_1 _10998_ (.A1(\m_sys.m_uart.m_tx.r_cycle_cnt[5] ),
    .A2(_02535_),
    .Y(_02537_),
    .B1(net3098));
 sg13g2_and3_1 _10999_ (.X(_02538_),
    .A(\m_sys.m_uart.m_tx.r_cycle_cnt[5] ),
    .B(net3098),
    .C(_02535_));
 sg13g2_nor3_1 _11000_ (.A(net4691),
    .B(net3099),
    .C(_02538_),
    .Y(_01772_));
 sg13g2_and2_1 _11001_ (.A(net3213),
    .B(_02538_),
    .X(_02539_));
 sg13g2_nor2_1 _11002_ (.A(net3213),
    .B(_02538_),
    .Y(_02540_));
 sg13g2_nor3_1 _11003_ (.A(net4691),
    .B(_02539_),
    .C(net3214),
    .Y(_01773_));
 sg13g2_nor2_1 _11004_ (.A(net3221),
    .B(_02539_),
    .Y(_02541_));
 sg13g2_and2_1 _11005_ (.A(net3221),
    .B(_02539_),
    .X(_02542_));
 sg13g2_nor3_1 _11006_ (.A(net4691),
    .B(_02541_),
    .C(_02542_),
    .Y(_01774_));
 sg13g2_xnor2_1 _11007_ (.Y(_02543_),
    .A(net3140),
    .B(_02542_));
 sg13g2_nor2_1 _11008_ (.A(net4691),
    .B(net3141),
    .Y(_01775_));
 sg13g2_a21oi_1 _11009_ (.A1(\m_sys.m_uart.m_tx.r_cycle_cnt[9] ),
    .A2(_02542_),
    .Y(_02544_),
    .B1(net3031));
 sg13g2_and3_2 _11010_ (.X(_02545_),
    .A(net3140),
    .B(net3031),
    .C(_02542_));
 sg13g2_nor3_1 _11011_ (.A(net4691),
    .B(net3032),
    .C(_02545_),
    .Y(_01761_));
 sg13g2_xnor2_1 _11012_ (.Y(_02546_),
    .A(net3247),
    .B(_02545_));
 sg13g2_nor2_1 _11013_ (.A(net4692),
    .B(_02546_),
    .Y(_01762_));
 sg13g2_a21oi_1 _11014_ (.A1(\m_sys.m_uart.m_tx.r_cycle_cnt[11] ),
    .A2(_02545_),
    .Y(_02547_),
    .B1(net2936));
 sg13g2_and3_1 _11015_ (.X(_02548_),
    .A(\m_sys.m_uart.m_tx.r_cycle_cnt[11] ),
    .B(net2936),
    .C(_02545_));
 sg13g2_nor3_1 _11016_ (.A(net4692),
    .B(net2937),
    .C(_02548_),
    .Y(_01763_));
 sg13g2_nor2_1 _11017_ (.A(net3146),
    .B(_02548_),
    .Y(_02549_));
 sg13g2_and2_1 _11018_ (.A(net3146),
    .B(_02548_),
    .X(_02550_));
 sg13g2_nor3_1 _11019_ (.A(net4692),
    .B(net3147),
    .C(_02550_),
    .Y(_01764_));
 sg13g2_nor2_1 _11020_ (.A(net3163),
    .B(_02550_),
    .Y(_02551_));
 sg13g2_and2_1 _11021_ (.A(net3163),
    .B(_02550_),
    .X(_02552_));
 sg13g2_nor3_1 _11022_ (.A(net4692),
    .B(_02551_),
    .C(_02552_),
    .Y(_01765_));
 sg13g2_a21oi_1 _11023_ (.A1(net3278),
    .A2(_02552_),
    .Y(_02553_),
    .B1(net4692));
 sg13g2_o21ai_1 _11024_ (.B1(_02553_),
    .Y(_02554_),
    .A1(net3278),
    .A2(_02552_));
 sg13g2_inv_1 _11025_ (.Y(_01766_),
    .A(_02554_));
 sg13g2_nand2b_1 _11026_ (.Y(_02555_),
    .B(\m_sys.m_uart.m_rx.io_i_ncycle[8] ),
    .A_N(\m_sys.m_uart.m_rx.r_cycle_cnt[7] ));
 sg13g2_xnor2_1 _11027_ (.Y(_02556_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[7] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[6] ));
 sg13g2_xnor2_1 _11028_ (.Y(_02557_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[1] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[0] ));
 sg13g2_nand2b_1 _11029_ (.Y(_02558_),
    .B(\m_sys.m_uart.m_rx.io_i_ncycle[2] ),
    .A_N(\m_sys.m_uart.m_rx.r_cycle_cnt[1] ));
 sg13g2_a22oi_1 _11030_ (.Y(_02559_),
    .B1(_02395_),
    .B2(\m_sys.m_uart.m_rx.io_i_ncycle[15] ),
    .A2(\m_sys.m_uart.m_rx.r_cycle_cnt[8] ),
    .A1(_02349_));
 sg13g2_xnor2_1 _11031_ (.Y(_02560_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[12] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[11] ));
 sg13g2_xnor2_1 _11032_ (.Y(_02561_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[11] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[10] ));
 sg13g2_a22oi_1 _11033_ (.Y(_02562_),
    .B1(\m_sys.m_uart.m_rx.r_cycle_cnt[12] ),
    .B2(_02346_),
    .A2(_02390_),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[3] ));
 sg13g2_xnor2_1 _11034_ (.Y(_02563_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[5] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[4] ));
 sg13g2_a22oi_1 _11035_ (.Y(_02564_),
    .B1(\m_sys.m_uart.m_rx.r_cycle_cnt[7] ),
    .B2(_02350_),
    .A2(_02391_),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[4] ));
 sg13g2_a22oi_1 _11036_ (.Y(_02565_),
    .B1(\m_sys.m_uart.m_rx.r_cycle_cnt[14] ),
    .B2(_02344_),
    .A2(_02394_),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[14] ));
 sg13g2_xnor2_1 _11037_ (.Y(_02566_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[10] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[9] ));
 sg13g2_a22oi_1 _11038_ (.Y(_02567_),
    .B1(\m_sys.m_uart.m_rx.r_cycle_cnt[2] ),
    .B2(_02355_),
    .A2(\m_sys.m_uart.m_rx.r_cycle_cnt[1] ),
    .A1(_02356_));
 sg13g2_and4_1 _11039_ (.A(_02564_),
    .B(_02565_),
    .C(_02566_),
    .D(_02567_),
    .X(_02568_));
 sg13g2_o21ai_1 _11040_ (.B1(_02555_),
    .Y(_02569_),
    .A1(_02346_),
    .A2(\m_sys.m_uart.m_rx.r_cycle_cnt[12] ));
 sg13g2_a21oi_1 _11041_ (.A1(_02345_),
    .A2(\m_sys.m_uart.m_rx.r_cycle_cnt[13] ),
    .Y(_02570_),
    .B1(_02569_));
 sg13g2_o21ai_1 _11042_ (.B1(_02558_),
    .Y(_02571_),
    .A1(_02352_),
    .A2(\m_sys.m_uart.m_rx.r_cycle_cnt[5] ));
 sg13g2_a221oi_1 _11043_ (.B2(_02352_),
    .C1(_02571_),
    .B1(\m_sys.m_uart.m_rx.r_cycle_cnt[5] ),
    .A1(_02354_),
    .Y(_02572_),
    .A2(\m_sys.m_uart.m_rx.r_cycle_cnt[3] ));
 sg13g2_nand4_1 _11044_ (.B(_02557_),
    .C(_02559_),
    .A(_02556_),
    .Y(_02573_),
    .D(_02562_));
 sg13g2_a21oi_1 _11045_ (.A1(\m_sys.m_uart.m_rx.io_i_ncycle[9] ),
    .A2(_02393_),
    .Y(_02574_),
    .B1(\m_sys.m_uart.m_rx.r_cycle_cnt[15] ));
 sg13g2_nand4_1 _11046_ (.B(_02561_),
    .C(_02563_),
    .A(_02560_),
    .Y(_02575_),
    .D(_02574_));
 sg13g2_nor2_1 _11047_ (.A(_02573_),
    .B(_02575_),
    .Y(_02576_));
 sg13g2_nand4_1 _11048_ (.B(_02570_),
    .C(_02572_),
    .A(_02568_),
    .Y(_02577_),
    .D(_02576_));
 sg13g2_nand3_1 _11049_ (.B(_02365_),
    .C(_02577_),
    .A(net2903),
    .Y(_02578_));
 sg13g2_inv_1 _11050_ (.Y(_02579_),
    .A(_02578_));
 sg13g2_xor2_1 _11051_ (.B(\m_sys.m_uart.m_rx.r_cycle_cnt[7] ),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[7] ),
    .X(_02580_));
 sg13g2_a221oi_1 _11052_ (.B2(_02350_),
    .C1(_02580_),
    .B1(\m_sys.m_uart.m_rx.r_cycle_cnt[8] ),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[4] ),
    .Y(_02581_),
    .A2(_02392_));
 sg13g2_xnor2_1 _11053_ (.Y(_02582_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[6] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[6] ));
 sg13g2_a22oi_1 _11054_ (.Y(_02583_),
    .B1(\m_sys.m_uart.m_rx.r_cycle_cnt[13] ),
    .B2(_02346_),
    .A2(_02393_),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[8] ));
 sg13g2_xor2_1 _11055_ (.B(\m_sys.m_uart.m_rx.r_cycle_cnt[14] ),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[14] ),
    .X(_02584_));
 sg13g2_xor2_1 _11056_ (.B(\m_sys.m_uart.m_rx.r_cycle_cnt[0] ),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[0] ),
    .X(_02585_));
 sg13g2_xor2_1 _11057_ (.B(\m_sys.m_uart.m_rx.r_cycle_cnt[2] ),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[2] ),
    .X(_02586_));
 sg13g2_xor2_1 _11058_ (.B(\m_sys.m_uart.m_rx.r_cycle_cnt[3] ),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[3] ),
    .X(_02587_));
 sg13g2_nor4_1 _11059_ (.A(_02584_),
    .B(_02585_),
    .C(_02586_),
    .D(_02587_),
    .Y(_02588_));
 sg13g2_nand4_1 _11060_ (.B(_02582_),
    .C(_02583_),
    .A(_02581_),
    .Y(_02589_),
    .D(_02588_));
 sg13g2_xnor2_1 _11061_ (.Y(_02590_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[15] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[15] ));
 sg13g2_xnor2_1 _11062_ (.Y(_02591_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[9] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[9] ));
 sg13g2_xnor2_1 _11063_ (.Y(_02592_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[12] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[12] ));
 sg13g2_xnor2_1 _11064_ (.Y(_02593_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[11] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[11] ));
 sg13g2_nand4_1 _11065_ (.B(_02591_),
    .C(_02592_),
    .A(_02590_),
    .Y(_02594_),
    .D(_02593_));
 sg13g2_xnor2_1 _11066_ (.Y(_02595_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[1] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[1] ));
 sg13g2_a22oi_1 _11067_ (.Y(_02596_),
    .B1(_02394_),
    .B2(\m_sys.m_uart.m_rx.io_i_ncycle[13] ),
    .A2(\m_sys.m_uart.m_rx.r_cycle_cnt[4] ),
    .A1(_02354_));
 sg13g2_xnor2_1 _11068_ (.Y(_02597_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[5] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[5] ));
 sg13g2_xnor2_1 _11069_ (.Y(_02598_),
    .A(\m_sys.m_uart.m_rx.io_i_ncycle[10] ),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[10] ));
 sg13g2_nand4_1 _11070_ (.B(_02596_),
    .C(_02597_),
    .A(_02595_),
    .Y(_02599_),
    .D(_02598_));
 sg13g2_or3_1 _11071_ (.A(_02589_),
    .B(_02594_),
    .C(_02599_),
    .X(_02600_));
 sg13g2_a21oi_1 _11072_ (.A1(\m_sys.m_uart.m_rx.r_cstate[1] ),
    .A2(_02600_),
    .Y(_02601_),
    .B1(_02579_));
 sg13g2_inv_2 _11073_ (.Y(_02602_),
    .A(net4368));
 sg13g2_nor2_1 _11074_ (.A(net3236),
    .B(net4368),
    .Y(_01744_));
 sg13g2_o21ai_1 _11075_ (.B1(_02602_),
    .Y(_02603_),
    .A1(net3236),
    .A2(net3288));
 sg13g2_a21oi_1 _11076_ (.A1(net3236),
    .A2(net3288),
    .Y(_01751_),
    .B1(_02603_));
 sg13g2_a21oi_1 _11077_ (.A1(\m_sys.m_uart.m_rx.r_cycle_cnt[0] ),
    .A2(\m_sys.m_uart.m_rx.r_cycle_cnt[1] ),
    .Y(_02604_),
    .B1(net3182));
 sg13g2_and3_1 _11078_ (.X(_02605_),
    .A(net3451),
    .B(\m_sys.m_uart.m_rx.r_cycle_cnt[1] ),
    .C(net3182));
 sg13g2_nor3_1 _11079_ (.A(net4368),
    .B(net3183),
    .C(_02605_),
    .Y(_01752_));
 sg13g2_and2_1 _11080_ (.A(net3268),
    .B(_02605_),
    .X(_02606_));
 sg13g2_nor2_1 _11081_ (.A(net3268),
    .B(_02605_),
    .Y(_02607_));
 sg13g2_nor3_1 _11082_ (.A(net4368),
    .B(_02606_),
    .C(net3269),
    .Y(_01753_));
 sg13g2_and2_1 _11083_ (.A(net3317),
    .B(_02606_),
    .X(_02608_));
 sg13g2_nor2_1 _11084_ (.A(net3317),
    .B(_02606_),
    .Y(_02609_));
 sg13g2_nor3_1 _11085_ (.A(net4367),
    .B(_02608_),
    .C(_02609_),
    .Y(_01754_));
 sg13g2_and2_1 _11086_ (.A(net3273),
    .B(_02608_),
    .X(_02610_));
 sg13g2_nor2_1 _11087_ (.A(net3273),
    .B(_02608_),
    .Y(_02611_));
 sg13g2_nor3_1 _11088_ (.A(net4367),
    .B(_02610_),
    .C(net3274),
    .Y(_01755_));
 sg13g2_and2_1 _11089_ (.A(net3259),
    .B(_02610_),
    .X(_02612_));
 sg13g2_nor2_1 _11090_ (.A(net3259),
    .B(_02610_),
    .Y(_02613_));
 sg13g2_nor3_1 _11091_ (.A(net4367),
    .B(_02612_),
    .C(net3260),
    .Y(_01756_));
 sg13g2_and2_1 _11092_ (.A(net3277),
    .B(_02612_),
    .X(_02614_));
 sg13g2_nor2_1 _11093_ (.A(net3277),
    .B(_02612_),
    .Y(_02615_));
 sg13g2_nor3_1 _11094_ (.A(net4367),
    .B(_02614_),
    .C(_02615_),
    .Y(_01757_));
 sg13g2_and2_1 _11095_ (.A(net3266),
    .B(_02614_),
    .X(_02616_));
 sg13g2_nor2_1 _11096_ (.A(net3266),
    .B(_02614_),
    .Y(_02617_));
 sg13g2_nor3_1 _11097_ (.A(net4367),
    .B(_02616_),
    .C(net3267),
    .Y(_01758_));
 sg13g2_xnor2_1 _11098_ (.Y(_02618_),
    .A(net3379),
    .B(_02616_));
 sg13g2_nor2_1 _11099_ (.A(net4367),
    .B(_02618_),
    .Y(_01759_));
 sg13g2_a21oi_1 _11100_ (.A1(\m_sys.m_uart.m_rx.r_cycle_cnt[9] ),
    .A2(_02616_),
    .Y(_02619_),
    .B1(net3149));
 sg13g2_and3_1 _11101_ (.X(_02620_),
    .A(net3450),
    .B(net3149),
    .C(_02616_));
 sg13g2_nor3_1 _11102_ (.A(net4367),
    .B(net3150),
    .C(_02620_),
    .Y(_01745_));
 sg13g2_nor2_1 _11103_ (.A(net3193),
    .B(_02620_),
    .Y(_02621_));
 sg13g2_and2_1 _11104_ (.A(net3193),
    .B(_02620_),
    .X(_02622_));
 sg13g2_nor3_1 _11105_ (.A(net4367),
    .B(net3194),
    .C(_02622_),
    .Y(_01746_));
 sg13g2_and2_1 _11106_ (.A(net3341),
    .B(_02622_),
    .X(_02623_));
 sg13g2_o21ai_1 _11107_ (.B1(_02602_),
    .Y(_02624_),
    .A1(net3341),
    .A2(_02622_));
 sg13g2_nor2_1 _11108_ (.A(_02623_),
    .B(_02624_),
    .Y(_01747_));
 sg13g2_and2_1 _11109_ (.A(net3332),
    .B(_02623_),
    .X(_02625_));
 sg13g2_o21ai_1 _11110_ (.B1(_02602_),
    .Y(_02626_),
    .A1(net3332),
    .A2(_02623_));
 sg13g2_nor2_1 _11111_ (.A(_02625_),
    .B(net3333),
    .Y(_01748_));
 sg13g2_and2_1 _11112_ (.A(net3400),
    .B(_02625_),
    .X(_02627_));
 sg13g2_o21ai_1 _11113_ (.B1(_02602_),
    .Y(_02628_),
    .A1(net3400),
    .A2(_02625_));
 sg13g2_nor2_1 _11114_ (.A(_02627_),
    .B(_02628_),
    .Y(_01749_));
 sg13g2_a21oi_1 _11115_ (.A1(net3334),
    .A2(_02627_),
    .Y(_02629_),
    .B1(net4368));
 sg13g2_o21ai_1 _11116_ (.B1(_02629_),
    .Y(_02630_),
    .A1(net3334),
    .A2(_02627_));
 sg13g2_inv_1 _11117_ (.Y(_01750_),
    .A(net3335));
 sg13g2_and2_2 _11118_ (.A(\m_sys._m_bootloader_io_b_mem_addr[1] ),
    .B(net5268),
    .X(_02631_));
 sg13g2_nand2_1 _11119_ (.Y(_02632_),
    .A(net5270),
    .B(net5267));
 sg13g2_nand2b_2 _11120_ (.Y(_02633_),
    .B(_02632_),
    .A_N(net5159));
 sg13g2_nand2b_2 _11121_ (.Y(_02634_),
    .B(\m_sys.m_core.m_fsm.r_cstate[2] ),
    .A_N(\m_sys.m_core.m_fsm.r_cstate[3] ));
 sg13g2_nor2_2 _11122_ (.A(_02368_),
    .B(_02634_),
    .Y(_02635_));
 sg13g2_or2_1 _11123_ (.X(_02636_),
    .B(_02634_),
    .A(_02368_));
 sg13g2_a21oi_1 _11124_ (.A1(_02372_),
    .A2(net5142),
    .Y(_02637_),
    .B1(net5272));
 sg13g2_o21ai_1 _11125_ (.B1(_02637_),
    .Y(_02638_),
    .A1(_00010_),
    .A2(net5142));
 sg13g2_o21ai_1 _11126_ (.B1(_02638_),
    .Y(_02639_),
    .A1(net5234),
    .A2(\m_sys._m_bootloader_io_b_mem_addr[2] ));
 sg13g2_a21oi_1 _11127_ (.A1(_02374_),
    .A2(net5141),
    .Y(_02640_),
    .B1(net5272));
 sg13g2_o21ai_1 _11128_ (.B1(_02640_),
    .Y(_02641_),
    .A1(_00012_),
    .A2(net5141));
 sg13g2_o21ai_1 _11129_ (.B1(_02641_),
    .Y(_02642_),
    .A1(net5234),
    .A2(\m_sys._m_bootloader_io_b_mem_addr[3] ));
 sg13g2_nor2b_2 _11130_ (.A(_02639_),
    .B_N(_02642_),
    .Y(_02643_));
 sg13g2_nand2b_2 _11131_ (.Y(_02644_),
    .B(_02642_),
    .A_N(_02639_));
 sg13g2_nor2_2 _11132_ (.A(_02633_),
    .B(net4643),
    .Y(_02645_));
 sg13g2_and2_2 _11133_ (.A(_02639_),
    .B(_02642_),
    .X(_02646_));
 sg13g2_nand2_2 _11134_ (.Y(_02647_),
    .A(_02639_),
    .B(_02642_));
 sg13g2_nand2b_2 _11135_ (.Y(_02648_),
    .B(net4606),
    .A_N(_02633_));
 sg13g2_nor2b_1 _11136_ (.A(_02642_),
    .B_N(_02639_),
    .Y(_02649_));
 sg13g2_nand2b_1 _11137_ (.Y(_02650_),
    .B(_02639_),
    .A_N(_02642_));
 sg13g2_nor2_1 _11138_ (.A(_02633_),
    .B(net4551),
    .Y(_02651_));
 sg13g2_a22oi_1 _11139_ (.Y(_02652_),
    .B1(net4391),
    .B2(uio_out[0]),
    .A2(_02645_),
    .A1(net3293));
 sg13g2_nor2_1 _11140_ (.A(uio_oe[0]),
    .B(net4393),
    .Y(_02653_));
 sg13g2_a21oi_2 _11141_ (.B1(_02653_),
    .Y(_00000_),
    .A2(net3294),
    .A1(net4393));
 sg13g2_a22oi_1 _11142_ (.Y(_02654_),
    .B1(net4391),
    .B2(uio_out[1]),
    .A2(_02645_),
    .A1(net3227));
 sg13g2_nor2_1 _11143_ (.A(uio_oe[1]),
    .B(net4393),
    .Y(_02655_));
 sg13g2_a21oi_1 _11144_ (.A1(net4393),
    .A2(net3228),
    .Y(_00001_),
    .B1(_02655_));
 sg13g2_a22oi_1 _11145_ (.Y(_02656_),
    .B1(net4391),
    .B2(uio_out[2]),
    .A2(_02645_),
    .A1(net3254));
 sg13g2_nor2_1 _11146_ (.A(uio_oe[2]),
    .B(net4393),
    .Y(_02657_));
 sg13g2_a21oi_2 _11147_ (.B1(_02657_),
    .Y(_00002_),
    .A2(net3255),
    .A1(net4393));
 sg13g2_a22oi_1 _11148_ (.Y(_02658_),
    .B1(net4391),
    .B2(uio_out[3]),
    .A2(_02645_),
    .A1(net3217));
 sg13g2_nor2_1 _11149_ (.A(uio_oe[3]),
    .B(net4393),
    .Y(_02659_));
 sg13g2_a21oi_2 _11150_ (.B1(_02659_),
    .Y(_00003_),
    .A2(net3218),
    .A1(_02648_));
 sg13g2_a22oi_1 _11151_ (.Y(_02660_),
    .B1(net4391),
    .B2(net3225),
    .A2(_02645_),
    .A1(net3284));
 sg13g2_nor2_1 _11152_ (.A(uio_oe[4]),
    .B(net4394),
    .Y(_02661_));
 sg13g2_a21oi_2 _11153_ (.B1(_02661_),
    .Y(_00004_),
    .A2(_02660_),
    .A1(net4394));
 sg13g2_a22oi_1 _11154_ (.Y(_02662_),
    .B1(net4391),
    .B2(uio_out[5]),
    .A2(_02645_),
    .A1(net3198));
 sg13g2_nor2_1 _11155_ (.A(uio_oe[5]),
    .B(net4394),
    .Y(_02663_));
 sg13g2_a21oi_2 _11156_ (.B1(_02663_),
    .Y(_00005_),
    .A2(net3199),
    .A1(net4394));
 sg13g2_a22oi_1 _11157_ (.Y(_02664_),
    .B1(net4391),
    .B2(uio_out[6]),
    .A2(_02645_),
    .A1(net3281));
 sg13g2_nor2_1 _11158_ (.A(uio_oe[6]),
    .B(net4394),
    .Y(_02665_));
 sg13g2_a21oi_2 _11159_ (.B1(_02665_),
    .Y(_00006_),
    .A2(net3282),
    .A1(net4394));
 sg13g2_a22oi_1 _11160_ (.Y(_02666_),
    .B1(net4391),
    .B2(net3306),
    .A2(_02645_),
    .A1(net3345));
 sg13g2_nor2_1 _11161_ (.A(uio_oe[7]),
    .B(net4394),
    .Y(_02667_));
 sg13g2_a21oi_2 _11162_ (.B1(_02667_),
    .Y(_00007_),
    .A2(_02666_),
    .A1(net4394));
 sg13g2_nor2_2 _11163_ (.A(_02332_),
    .B(_02340_),
    .Y(uo_out[0]));
 sg13g2_nor2_2 _11164_ (.A(_02331_),
    .B(_02339_),
    .Y(uo_out[1]));
 sg13g2_nor2_2 _11165_ (.A(_02330_),
    .B(_02338_),
    .Y(uo_out[2]));
 sg13g2_nor2_2 _11166_ (.A(_02329_),
    .B(_02337_),
    .Y(uo_out[3]));
 sg13g2_nor2_2 _11167_ (.A(_02327_),
    .B(_02335_),
    .Y(uo_out[5]));
 sg13g2_nor2_2 _11168_ (.A(_02326_),
    .B(_02334_),
    .Y(uo_out[6]));
 sg13g2_nor2_1 _11169_ (.A(_02325_),
    .B(_02333_),
    .Y(uo_out[7]));
 sg13g2_a21o_1 _11170_ (.A2(_02635_),
    .A1(_00008_),
    .B1(net5272),
    .X(_02668_));
 sg13g2_a21oi_2 _11171_ (.B1(_02668_),
    .Y(_02669_),
    .A2(net5141),
    .A1(_00009_));
 sg13g2_a21oi_2 _11172_ (.B1(_02669_),
    .Y(_02670_),
    .A2(\m_sys._m_bootloader_io_b_mem_addr[4] ),
    .A1(net5268));
 sg13g2_a21o_2 _11173_ (.A2(\m_sys._m_bootloader_io_b_mem_addr[4] ),
    .A1(net5268),
    .B1(_02669_),
    .X(_02671_));
 sg13g2_nor3_1 _11174_ (.A(_02633_),
    .B(net4643),
    .C(_02671_),
    .Y(_02672_));
 sg13g2_and2_1 _11175_ (.A(net2952),
    .B(net4388),
    .X(_00147_));
 sg13g2_and2_1 _11176_ (.A(net3109),
    .B(net4388),
    .X(_00148_));
 sg13g2_and2_1 _11177_ (.A(net3076),
    .B(net4388),
    .X(_00149_));
 sg13g2_and2_1 _11178_ (.A(net3201),
    .B(net4388),
    .X(_00150_));
 sg13g2_and2_1 _11179_ (.A(net3319),
    .B(net4390),
    .X(_00151_));
 sg13g2_and2_1 _11180_ (.A(net3090),
    .B(net4388),
    .X(_00152_));
 sg13g2_and2_1 _11181_ (.A(net3216),
    .B(net4388),
    .X(_00153_));
 sg13g2_and2_1 _11182_ (.A(net3053),
    .B(net4388),
    .X(_00154_));
 sg13g2_nand2_1 _11183_ (.Y(_02673_),
    .A(net5274),
    .B(net2458));
 sg13g2_o21ai_1 _11184_ (.B1(_02673_),
    .Y(_00155_),
    .A1(net5274),
    .A2(_02632_));
 sg13g2_mux2_1 _11185_ (.A0(net5357),
    .A1(net5159),
    .S(_02411_),
    .X(_00156_));
 sg13g2_nor2_1 _11186_ (.A(_02639_),
    .B(_02642_),
    .Y(_02674_));
 sg13g2_or2_2 _11187_ (.X(_02675_),
    .B(_02642_),
    .A(_02639_));
 sg13g2_mux2_1 _11188_ (.A0(_00022_),
    .A1(_00023_),
    .S(net5141),
    .X(_02676_));
 sg13g2_mux2_2 _11189_ (.A0(_00045_),
    .A1(_02676_),
    .S(net5234),
    .X(_02677_));
 sg13g2_nand2_1 _11190_ (.Y(_02678_),
    .A(net5269),
    .B(_00044_));
 sg13g2_nor2_1 _11191_ (.A(_00020_),
    .B(net5141),
    .Y(_02679_));
 sg13g2_o21ai_1 _11192_ (.B1(net5234),
    .Y(_02680_),
    .A1(_00021_),
    .A2(_02635_));
 sg13g2_o21ai_1 _11193_ (.B1(_02678_),
    .Y(_02681_),
    .A1(_02679_),
    .A2(_02680_));
 sg13g2_nor2_1 _11194_ (.A(_02677_),
    .B(_02681_),
    .Y(_02682_));
 sg13g2_nand2_2 _11195_ (.Y(_02683_),
    .A(_02670_),
    .B(_02682_));
 sg13g2_nor2_2 _11196_ (.A(net4506),
    .B(_02683_),
    .Y(_02684_));
 sg13g2_a21oi_2 _11197_ (.B1(net5234),
    .Y(_02685_),
    .A2(\m_sys._m_bootloader_io_b_mem_wen[0] ),
    .A1(_02367_));
 sg13g2_nand2_1 _11198_ (.Y(_02686_),
    .A(\m_sys.m_core.m_bru.io_i_pc[10] ),
    .B(net5142));
 sg13g2_o21ai_1 _11199_ (.B1(_02686_),
    .Y(_02687_),
    .A1(net5229),
    .A2(net5142));
 sg13g2_mux2_1 _11200_ (.A0(net5320),
    .A1(\m_sys.m_core.m_bru.io_i_pc[8] ),
    .S(net5141),
    .X(_02688_));
 sg13g2_nand2_1 _11201_ (.Y(_02689_),
    .A(\m_sys.m_core.m_bru.io_i_pc[9] ),
    .B(net5142));
 sg13g2_o21ai_1 _11202_ (.B1(_02689_),
    .Y(_02690_),
    .A1(net5228),
    .A2(net5141));
 sg13g2_and2_1 _11203_ (.A(_00019_),
    .B(net5141),
    .X(_02691_));
 sg13g2_a21oi_1 _11204_ (.A1(_00018_),
    .A2(_02635_),
    .Y(_02692_),
    .B1(_02691_));
 sg13g2_nor4_2 _11205_ (.A(_02687_),
    .B(_02688_),
    .C(_02690_),
    .Y(_02693_),
    .D(_02692_));
 sg13g2_nand2_1 _11206_ (.Y(_02694_),
    .A(_00017_),
    .B(net5142));
 sg13g2_o21ai_1 _11207_ (.B1(_02694_),
    .Y(_02695_),
    .A1(_02382_),
    .A2(net5142));
 sg13g2_inv_1 _11208_ (.Y(_02696_),
    .A(_02695_));
 sg13g2_and2_1 _11209_ (.A(_02693_),
    .B(_02695_),
    .X(_02697_));
 sg13g2_inv_2 _11210_ (.Y(_02698_),
    .A(net4493));
 sg13g2_nand2_2 _11211_ (.Y(_02699_),
    .A(net5242),
    .B(net5232));
 sg13g2_nand2_1 _11212_ (.Y(_02700_),
    .A(net5232),
    .B(_02635_));
 sg13g2_nor2_1 _11213_ (.A(net3448),
    .B(_02699_),
    .Y(_02701_));
 sg13g2_nor2_1 _11214_ (.A(_02635_),
    .B(_02701_),
    .Y(_02702_));
 sg13g2_a21oi_1 _11215_ (.A1(net5232),
    .A2(_02635_),
    .Y(_02703_),
    .B1(_02702_));
 sg13g2_and2_1 _11216_ (.A(net5235),
    .B(_02703_),
    .X(_02704_));
 sg13g2_nand2_1 _11217_ (.Y(_02705_),
    .A(net4494),
    .B(_02704_));
 sg13g2_nand2_2 _11218_ (.Y(_02706_),
    .A(\m_sys.m_bootloader.r_cstate[1] ),
    .B(_00024_));
 sg13g2_nor2_1 _11219_ (.A(net5284),
    .B(_02706_),
    .Y(_02707_));
 sg13g2_nand3_1 _11220_ (.B(net5283),
    .C(_02707_),
    .A(\m_sys.m_bootloader.r_cstate[3] ),
    .Y(_02708_));
 sg13g2_nor2b_2 _11221_ (.A(\m_sys.m_bootloader.r_cstate[1] ),
    .B_N(_00024_),
    .Y(_02709_));
 sg13g2_nand2b_2 _11222_ (.Y(_02710_),
    .B(_00024_),
    .A_N(\m_sys.m_bootloader.r_cstate[1] ));
 sg13g2_nand2_2 _11223_ (.Y(_02711_),
    .A(net5284),
    .B(_02709_));
 sg13g2_nand2b_2 _11224_ (.Y(_02712_),
    .B(net5282),
    .A_N(\m_sys.m_bootloader.r_cstate[2] ));
 sg13g2_o21ai_1 _11225_ (.B1(_02708_),
    .Y(_02713_),
    .A1(_02711_),
    .A2(_02712_));
 sg13g2_nand2_1 _11226_ (.Y(_02714_),
    .A(net5268),
    .B(_02713_));
 sg13g2_nor4_2 _11227_ (.A(\m_sys._m_bootloader_io_b_mem_addr[10] ),
    .B(\m_sys._m_bootloader_io_b_mem_addr[8] ),
    .C(\m_sys._m_bootloader_io_b_mem_addr[9] ),
    .Y(_02715_),
    .D(\m_sys._m_bootloader_io_b_mem_addr[7] ));
 sg13g2_and2_1 _11228_ (.A(_02387_),
    .B(_02715_),
    .X(_02716_));
 sg13g2_nand2_2 _11229_ (.Y(_02717_),
    .A(_02387_),
    .B(_02715_));
 sg13g2_o21ai_1 _11230_ (.B1(_02705_),
    .Y(_02718_),
    .A1(_02714_),
    .A2(_02717_));
 sg13g2_nand2_1 _11231_ (.Y(_02719_),
    .A(net5384),
    .B(net4361));
 sg13g2_nor2b_1 _11232_ (.A(\m_sys.m_core.r_ctrl_mem_size[0] ),
    .B_N(\m_sys.m_core.r_ctrl_mem_size[1] ),
    .Y(_02720_));
 sg13g2_and2_1 _11233_ (.A(\m_sys.m_core.r_ctrl_mem_rw ),
    .B(_02635_),
    .X(_02721_));
 sg13g2_a21oi_1 _11234_ (.A1(_02720_),
    .A2(_02721_),
    .Y(_02722_),
    .B1(net5272));
 sg13g2_and2_2 _11235_ (.A(net5268),
    .B(_00043_),
    .X(_02723_));
 sg13g2_nor3_2 _11236_ (.A(_02719_),
    .B(_02722_),
    .C(_02723_),
    .Y(_02724_));
 sg13g2_nand2b_1 _11237_ (.Y(_02725_),
    .B(_02724_),
    .A_N(_02685_));
 sg13g2_nor3_1 _11238_ (.A(net4506),
    .B(net4501),
    .C(net4333),
    .Y(_02726_));
 sg13g2_nor2_1 _11239_ (.A(net2716),
    .B(net4308),
    .Y(_02727_));
 sg13g2_nor2b_1 _11240_ (.A(net5266),
    .B_N(\m_sys._m_bootloader_io_b_mem_wdata[0] ),
    .Y(_02728_));
 sg13g2_a22oi_1 _11241_ (.Y(_02729_),
    .B1(_02631_),
    .B2(_02728_),
    .A2(\m_sys._m_core_io_b_mem_wdata[16] ),
    .A1(net5241));
 sg13g2_a21oi_1 _11242_ (.A1(net4308),
    .A2(net5136),
    .Y(_00157_),
    .B1(_02727_));
 sg13g2_nor2_1 _11243_ (.A(net2697),
    .B(net4308),
    .Y(_02730_));
 sg13g2_nor2_1 _11244_ (.A(net5266),
    .B(_02404_),
    .Y(_02731_));
 sg13g2_a22oi_1 _11245_ (.Y(_02732_),
    .B1(_02631_),
    .B2(_02731_),
    .A2(\m_sys._m_core_io_b_mem_wdata[17] ),
    .A1(net5241));
 sg13g2_a21oi_1 _11246_ (.A1(net4308),
    .A2(net4997),
    .Y(_00158_),
    .B1(_02730_));
 sg13g2_nor2_1 _11247_ (.A(net2724),
    .B(net4309),
    .Y(_02733_));
 sg13g2_nor2b_1 _11248_ (.A(net5266),
    .B_N(\m_sys._m_bootloader_io_b_mem_wdata[2] ),
    .Y(_02734_));
 sg13g2_a22oi_1 _11249_ (.Y(_02735_),
    .B1(_02631_),
    .B2(_02734_),
    .A2(\m_sys._m_core_io_b_mem_wdata[18] ),
    .A1(net5240));
 sg13g2_a21oi_1 _11250_ (.A1(net4309),
    .A2(net5133),
    .Y(_00159_),
    .B1(_02733_));
 sg13g2_nor2_1 _11251_ (.A(net2711),
    .B(net4308),
    .Y(_02736_));
 sg13g2_nor2_1 _11252_ (.A(net5266),
    .B(_02405_),
    .Y(_02737_));
 sg13g2_a22oi_1 _11253_ (.Y(_02738_),
    .B1(net5159),
    .B2(_02737_),
    .A2(\m_sys._m_core_io_b_mem_wdata[19] ),
    .A1(net5240));
 sg13g2_a21oi_1 _11254_ (.A1(net4308),
    .A2(net4989),
    .Y(_00160_),
    .B1(_02736_));
 sg13g2_nor2_1 _11255_ (.A(net2645),
    .B(net4309),
    .Y(_02739_));
 sg13g2_nor2b_1 _11256_ (.A(net5266),
    .B_N(\m_sys._m_bootloader_io_b_mem_wdata[4] ),
    .Y(_02740_));
 sg13g2_a22oi_1 _11257_ (.Y(_02741_),
    .B1(net5159),
    .B2(_02740_),
    .A2(\m_sys._m_core_io_b_mem_wdata[20] ),
    .A1(net5239));
 sg13g2_a21oi_1 _11258_ (.A1(net4309),
    .A2(net5128),
    .Y(_00161_),
    .B1(_02739_));
 sg13g2_nor2_1 _11259_ (.A(net2696),
    .B(net4308),
    .Y(_02742_));
 sg13g2_nor2_1 _11260_ (.A(net5267),
    .B(_02406_),
    .Y(_02743_));
 sg13g2_a22oi_1 _11261_ (.Y(_02744_),
    .B1(net5159),
    .B2(_02743_),
    .A2(\m_sys._m_core_io_b_mem_wdata[21] ),
    .A1(net5239));
 sg13g2_a21oi_1 _11262_ (.A1(net4308),
    .A2(net4987),
    .Y(_00162_),
    .B1(_02742_));
 sg13g2_nor2_1 _11263_ (.A(net2707),
    .B(net4309),
    .Y(_02745_));
 sg13g2_nor2b_1 _11264_ (.A(net5266),
    .B_N(\m_sys._m_bootloader_io_b_mem_wdata[6] ),
    .Y(_02746_));
 sg13g2_a22oi_1 _11265_ (.Y(_02747_),
    .B1(net5159),
    .B2(_02746_),
    .A2(\m_sys._m_core_io_b_mem_wdata[22] ),
    .A1(net5239));
 sg13g2_a21oi_1 _11266_ (.A1(net4309),
    .A2(net5122),
    .Y(_00163_),
    .B1(_02745_));
 sg13g2_nor2_1 _11267_ (.A(net2406),
    .B(net4309),
    .Y(_02748_));
 sg13g2_nor2_1 _11268_ (.A(net5266),
    .B(_02407_),
    .Y(_02749_));
 sg13g2_a22oi_1 _11269_ (.Y(_02750_),
    .B1(net5159),
    .B2(_02749_),
    .A2(\m_sys._m_core_io_b_mem_wdata[23] ),
    .A1(net5239));
 sg13g2_a21oi_1 _11270_ (.A1(net4309),
    .A2(net4981),
    .Y(_00164_),
    .B1(_02748_));
 sg13g2_nor2_2 _11271_ (.A(net5242),
    .B(\m_sys.m_core.m_fsm.r_cstate[3] ),
    .Y(_02751_));
 sg13g2_nor2_1 _11272_ (.A(net5242),
    .B(net5309),
    .Y(_02752_));
 sg13g2_nand2b_2 _11273_ (.Y(_02753_),
    .B(\m_sys.m_core.m_fsm.r_cstate[3] ),
    .A_N(\m_sys.m_core.m_fsm.r_cstate[2] ));
 sg13g2_nand3b_1 _11274_ (.B(net5232),
    .C(_02368_),
    .Y(_02754_),
    .A_N(_02753_));
 sg13g2_nor3_2 _11275_ (.A(net5232),
    .B(\m_sys.m_core.m_fsm.r_cstate[3] ),
    .C(\m_sys.m_core.m_fsm.r_cstate[2] ),
    .Y(_02755_));
 sg13g2_and2_2 _11276_ (.A(net5242),
    .B(_02755_),
    .X(_02756_));
 sg13g2_nand2_1 _11277_ (.Y(_02757_),
    .A(net5242),
    .B(_02755_));
 sg13g2_nand2_1 _11278_ (.Y(_02758_),
    .A(_02754_),
    .B(net4958));
 sg13g2_a21oi_2 _11279_ (.B1(_02758_),
    .Y(_02759_),
    .A2(_02751_),
    .A1(\m_sys.m_core.m_fsm.r_cstate[2] ));
 sg13g2_mux2_1 _11280_ (.A0(\m_sys.m_core.m_gpr._GEN[193] ),
    .A1(\m_sys.m_core.m_gpr._GEN[225] ),
    .S(net5335),
    .X(_02760_));
 sg13g2_nor2_1 _11281_ (.A(net5347),
    .B(net5339),
    .Y(_02761_));
 sg13g2_nand2_1 _11282_ (.Y(_02762_),
    .A(\m_sys.m_core.m_gpr._GEN[129] ),
    .B(net5153));
 sg13g2_nor2_1 _11283_ (.A(net5347),
    .B(net5205),
    .Y(_02763_));
 sg13g2_a221oi_1 _11284_ (.B2(\m_sys.m_core.m_gpr._GEN[161] ),
    .C1(net5210),
    .B1(net5113),
    .A1(net5344),
    .Y(_02764_),
    .A2(_02760_));
 sg13g2_and2_1 _11285_ (.A(_00067_),
    .B(net5153),
    .X(_02765_));
 sg13g2_nand2_1 _11286_ (.Y(_02766_),
    .A(_00067_),
    .B(net5153));
 sg13g2_mux2_1 _11287_ (.A0(\m_sys.m_core.m_gpr._GEN[65] ),
    .A1(\m_sys.m_core.m_gpr._GEN[97] ),
    .S(net5334),
    .X(_02767_));
 sg13g2_a22oi_1 _11288_ (.Y(_02768_),
    .B1(_02767_),
    .B2(net5343),
    .A2(net5113),
    .A1(\m_sys.m_core.m_gpr._GEN[33] ));
 sg13g2_a221oi_1 _11289_ (.B2(net5210),
    .C1(net5108),
    .B1(_02768_),
    .A1(_02762_),
    .Y(_02769_),
    .A2(_02764_));
 sg13g2_nand2_1 _11290_ (.Y(_02770_),
    .A(net5312),
    .B(\m_sys.m_core.m_bru.io_i_s1[0] ));
 sg13g2_nor3_1 _11291_ (.A(\m_sys.m_core.m_bru.io_i_s1[2] ),
    .B(net5313),
    .C(_02770_),
    .Y(_02771_));
 sg13g2_and2_2 _11292_ (.A(net5226),
    .B(_02771_),
    .X(_02772_));
 sg13g2_nor2b_2 _11293_ (.A(net5315),
    .B_N(_02772_),
    .Y(_02773_));
 sg13g2_inv_1 _11294_ (.Y(_02774_),
    .A(_02773_));
 sg13g2_nand2b_2 _11295_ (.Y(_02775_),
    .B(net5317),
    .A_N(net5315));
 sg13g2_and4_2 _11296_ (.A(net5318),
    .B(_00022_),
    .C(net4972),
    .D(_02773_),
    .X(_02776_));
 sg13g2_nand4_1 _11297_ (.B(_00022_),
    .C(net4972),
    .A(net5317),
    .Y(_02777_),
    .D(_02773_));
 sg13g2_a22oi_1 _11298_ (.Y(_02778_),
    .B1(_02769_),
    .B2(net4733),
    .A2(net4735),
    .A1(\m_sys._m_core_io_b_mem_wdata[1] ));
 sg13g2_nor2_1 _11299_ (.A(_00022_),
    .B(_02775_),
    .Y(_02779_));
 sg13g2_nand2_1 _11300_ (.Y(_02780_),
    .A(\m_sys.m_core.m_bru.io_i_s1[2] ),
    .B(net5313));
 sg13g2_nor4_1 _11301_ (.A(_00022_),
    .B(_02770_),
    .C(_02775_),
    .D(_02780_),
    .Y(_02781_));
 sg13g2_and2_2 _11302_ (.A(_02771_),
    .B(_02779_),
    .X(_02782_));
 sg13g2_o21ai_1 _11303_ (.B1(net4973),
    .Y(_02783_),
    .A1(net5102),
    .A2(net4957));
 sg13g2_mux2_1 _11304_ (.A0(net3320),
    .A1(_00065_),
    .S(net5102),
    .X(_02784_));
 sg13g2_o21ai_1 _11305_ (.B1(_02778_),
    .Y(_00165_),
    .A1(net4786),
    .A2(_02784_));
 sg13g2_nor2_1 _11306_ (.A(net5205),
    .B(\m_sys.m_core.m_gpr._GEN[226] ),
    .Y(_02785_));
 sg13g2_o21ai_1 _11307_ (.B1(net5347),
    .Y(_02786_),
    .A1(net5339),
    .A2(\m_sys.m_core.m_gpr._GEN[194] ));
 sg13g2_a221oi_1 _11308_ (.B2(\m_sys.m_core.m_gpr._GEN[162] ),
    .C1(net5215),
    .B1(net5117),
    .A1(\m_sys.m_core.m_gpr._GEN[130] ),
    .Y(_02787_),
    .A2(net5156));
 sg13g2_o21ai_1 _11309_ (.B1(_02787_),
    .Y(_02788_),
    .A1(_02785_),
    .A2(_02786_));
 sg13g2_nor2_1 _11310_ (.A(net5339),
    .B(\m_sys.m_core.m_gpr._GEN[66] ),
    .Y(_02789_));
 sg13g2_o21ai_1 _11311_ (.B1(net5347),
    .Y(_02790_),
    .A1(net5205),
    .A2(\m_sys.m_core.m_gpr._GEN[98] ));
 sg13g2_a21oi_1 _11312_ (.A1(\m_sys.m_core.m_gpr._GEN[34] ),
    .A2(net5117),
    .Y(_02791_),
    .B1(net5351));
 sg13g2_o21ai_1 _11313_ (.B1(_02791_),
    .Y(_02792_),
    .A1(_02789_),
    .A2(_02790_));
 sg13g2_nand3_1 _11314_ (.B(_02788_),
    .C(_02792_),
    .A(net5106),
    .Y(_02793_));
 sg13g2_nor2_1 _11315_ (.A(net4732),
    .B(_02793_),
    .Y(_02794_));
 sg13g2_a21oi_1 _11316_ (.A1(\m_sys._m_core_io_b_mem_wdata[2] ),
    .A2(net4735),
    .Y(_02795_),
    .B1(_02794_));
 sg13g2_nand2_1 _11317_ (.Y(_02796_),
    .A(_00067_),
    .B(net5102));
 sg13g2_o21ai_1 _11318_ (.B1(_02796_),
    .Y(_02797_),
    .A1(_02426_),
    .A2(net5103));
 sg13g2_o21ai_1 _11319_ (.B1(_02795_),
    .Y(_00166_),
    .A1(net4787),
    .A2(_02797_));
 sg13g2_a21oi_1 _11320_ (.A1(net5205),
    .A2(_02429_),
    .Y(_02798_),
    .B1(net5220));
 sg13g2_o21ai_1 _11321_ (.B1(_02798_),
    .Y(_02799_),
    .A1(net5205),
    .A2(\m_sys.m_core.m_gpr._GEN[227] ));
 sg13g2_a221oi_1 _11322_ (.B2(\m_sys.m_core.m_gpr._GEN[163] ),
    .C1(net5215),
    .B1(net5117),
    .A1(\m_sys.m_core.m_gpr._GEN[131] ),
    .Y(_02800_),
    .A2(net5156));
 sg13g2_mux2_1 _11323_ (.A0(\m_sys.m_core.m_gpr._GEN[67] ),
    .A1(\m_sys.m_core.m_gpr._GEN[99] ),
    .S(net5339),
    .X(_02801_));
 sg13g2_a22oi_1 _11324_ (.Y(_02802_),
    .B1(_02801_),
    .B2(net5349),
    .A2(net5117),
    .A1(\m_sys.m_core.m_gpr._GEN[35] ));
 sg13g2_a221oi_1 _11325_ (.B2(net5215),
    .C1(net5109),
    .B1(_02802_),
    .A1(_02799_),
    .Y(_02803_),
    .A2(_02800_));
 sg13g2_mux2_1 _11326_ (.A0(net3299),
    .A1(_00069_),
    .S(net5103),
    .X(_02804_));
 sg13g2_a22oi_1 _11327_ (.Y(_02805_),
    .B1(net4733),
    .B2(_02803_),
    .A2(net4735),
    .A1(\m_sys._m_core_io_b_mem_wdata[3] ));
 sg13g2_o21ai_1 _11328_ (.B1(_02805_),
    .Y(_00167_),
    .A1(net4787),
    .A2(net3300));
 sg13g2_mux2_1 _11329_ (.A0(\m_sys.m_core.m_gpr._GEN[196] ),
    .A1(\m_sys.m_core.m_gpr._GEN[228] ),
    .S(net5334),
    .X(_02806_));
 sg13g2_nand2_1 _11330_ (.Y(_02807_),
    .A(\m_sys.m_core.m_gpr._GEN[132] ),
    .B(net5153));
 sg13g2_a221oi_1 _11331_ (.B2(net5344),
    .C1(net5211),
    .B1(_02806_),
    .A1(\m_sys.m_core.m_gpr._GEN[164] ),
    .Y(_02808_),
    .A2(net5112));
 sg13g2_mux2_1 _11332_ (.A0(\m_sys.m_core.m_gpr._GEN[68] ),
    .A1(\m_sys.m_core.m_gpr._GEN[100] ),
    .S(net5334),
    .X(_02809_));
 sg13g2_a22oi_1 _11333_ (.Y(_02810_),
    .B1(_02809_),
    .B2(net5343),
    .A2(net5112),
    .A1(\m_sys.m_core.m_gpr._GEN[36] ));
 sg13g2_a22oi_1 _11334_ (.Y(_02811_),
    .B1(_02810_),
    .B2(net5210),
    .A2(_02808_),
    .A1(_02807_));
 sg13g2_nand2_2 _11335_ (.Y(_02812_),
    .A(net5106),
    .B(_02811_));
 sg13g2_nor2_1 _11336_ (.A(net4732),
    .B(_02812_),
    .Y(_02813_));
 sg13g2_a21oi_1 _11337_ (.A1(net3402),
    .A2(net4735),
    .Y(_02814_),
    .B1(_02813_));
 sg13g2_nand2_1 _11338_ (.Y(_02815_),
    .A(net3423),
    .B(net5102));
 sg13g2_o21ai_1 _11339_ (.B1(_02815_),
    .Y(_02816_),
    .A1(_02382_),
    .A2(net5103));
 sg13g2_o21ai_1 _11340_ (.B1(_02814_),
    .Y(_00168_),
    .A1(net4787),
    .A2(net3424));
 sg13g2_a21oi_1 _11341_ (.A1(net5198),
    .A2(_02433_),
    .Y(_02817_),
    .B1(net5218));
 sg13g2_o21ai_1 _11342_ (.B1(_02817_),
    .Y(_02818_),
    .A1(net5199),
    .A2(\m_sys.m_core.m_gpr._GEN[229] ));
 sg13g2_a221oi_1 _11343_ (.B2(\m_sys.m_core.m_gpr._GEN[165] ),
    .C1(net5210),
    .B1(net5111),
    .A1(\m_sys.m_core.m_gpr._GEN[133] ),
    .Y(_02819_),
    .A2(net5154));
 sg13g2_mux2_1 _11344_ (.A0(\m_sys.m_core.m_gpr._GEN[69] ),
    .A1(\m_sys.m_core.m_gpr._GEN[101] ),
    .S(net5333),
    .X(_02820_));
 sg13g2_a22oi_1 _11345_ (.Y(_02821_),
    .B1(_02820_),
    .B2(net5342),
    .A2(net5111),
    .A1(\m_sys.m_core.m_gpr._GEN[37] ));
 sg13g2_a221oi_1 _11346_ (.B2(net5209),
    .C1(net5107),
    .B1(_02821_),
    .A1(_02818_),
    .Y(_02822_),
    .A2(_02819_));
 sg13g2_a22oi_1 _11347_ (.Y(_02823_),
    .B1(net4734),
    .B2(_02822_),
    .A2(net4735),
    .A1(\m_sys._m_core_io_b_mem_wdata[5] ));
 sg13g2_o21ai_1 _11348_ (.B1(_02823_),
    .Y(_00169_),
    .A1(net3128),
    .A2(net4787));
 sg13g2_a21oi_1 _11349_ (.A1(net5199),
    .A2(_02436_),
    .Y(_02824_),
    .B1(net5220));
 sg13g2_o21ai_1 _11350_ (.B1(_02824_),
    .Y(_02825_),
    .A1(net5199),
    .A2(\m_sys.m_core.m_gpr._GEN[230] ));
 sg13g2_a221oi_1 _11351_ (.B2(\m_sys.m_core.m_gpr._GEN[166] ),
    .C1(net5211),
    .B1(net5113),
    .A1(\m_sys.m_core.m_gpr._GEN[134] ),
    .Y(_02826_),
    .A2(net5153));
 sg13g2_nor2_1 _11352_ (.A(net5334),
    .B(\m_sys.m_core.m_gpr._GEN[70] ),
    .Y(_02827_));
 sg13g2_a21oi_1 _11353_ (.A1(net5334),
    .A2(_02435_),
    .Y(_02828_),
    .B1(_02827_));
 sg13g2_a22oi_1 _11354_ (.Y(_02829_),
    .B1(_02828_),
    .B2(net5343),
    .A2(net5113),
    .A1(\m_sys.m_core.m_gpr._GEN[38] ));
 sg13g2_a221oi_1 _11355_ (.B2(net5211),
    .C1(net5108),
    .B1(_02829_),
    .A1(_02825_),
    .Y(_02830_),
    .A2(_02826_));
 sg13g2_a22oi_1 _11356_ (.Y(_02831_),
    .B1(net4734),
    .B2(_02830_),
    .A2(net4736),
    .A1(\m_sys._m_core_io_b_mem_wdata[6] ));
 sg13g2_o21ai_1 _11357_ (.B1(_02831_),
    .Y(_00170_),
    .A1(net3232),
    .A2(net4786));
 sg13g2_a21oi_1 _11358_ (.A1(net5199),
    .A2(_02438_),
    .Y(_02832_),
    .B1(net5218));
 sg13g2_o21ai_1 _11359_ (.B1(_02832_),
    .Y(_02833_),
    .A1(net5199),
    .A2(\m_sys.m_core.m_gpr._GEN[231] ));
 sg13g2_a221oi_1 _11360_ (.B2(\m_sys.m_core.m_gpr._GEN[167] ),
    .C1(net5210),
    .B1(net5112),
    .A1(\m_sys.m_core.m_gpr._GEN[135] ),
    .Y(_02834_),
    .A2(net5153));
 sg13g2_mux2_1 _11361_ (.A0(\m_sys.m_core.m_gpr._GEN[71] ),
    .A1(\m_sys.m_core.m_gpr._GEN[103] ),
    .S(net5334),
    .X(_02835_));
 sg13g2_a22oi_1 _11362_ (.Y(_02836_),
    .B1(_02835_),
    .B2(net5343),
    .A2(net5112),
    .A1(\m_sys.m_core.m_gpr._GEN[39] ));
 sg13g2_a221oi_1 _11363_ (.B2(net5211),
    .C1(net5108),
    .B1(_02836_),
    .A1(_02833_),
    .Y(_02837_),
    .A2(_02834_));
 sg13g2_a22oi_1 _11364_ (.Y(_02838_),
    .B1(net4733),
    .B2(_02837_),
    .A2(net4735),
    .A1(\m_sys._m_core_io_b_mem_wdata[7] ));
 sg13g2_o21ai_1 _11365_ (.B1(_02838_),
    .Y(_00171_),
    .A1(net3360),
    .A2(net4786));
 sg13g2_mux2_1 _11366_ (.A0(\m_sys.m_core.m_gpr._GEN[200] ),
    .A1(\m_sys.m_core.m_gpr._GEN[232] ),
    .S(net5336),
    .X(_02839_));
 sg13g2_nand2_1 _11367_ (.Y(_02840_),
    .A(\m_sys.m_core.m_gpr._GEN[136] ),
    .B(net5157));
 sg13g2_a221oi_1 _11368_ (.B2(net5347),
    .C1(net5215),
    .B1(_02839_),
    .A1(\m_sys.m_core.m_gpr._GEN[168] ),
    .Y(_02841_),
    .A2(net5117));
 sg13g2_mux2_1 _11369_ (.A0(\m_sys.m_core.m_gpr._GEN[72] ),
    .A1(\m_sys.m_core.m_gpr._GEN[104] ),
    .S(net5339),
    .X(_02842_));
 sg13g2_a22oi_1 _11370_ (.Y(_02843_),
    .B1(_02842_),
    .B2(net5347),
    .A2(net5117),
    .A1(\m_sys.m_core.m_gpr._GEN[40] ));
 sg13g2_a221oi_1 _11371_ (.B2(net5215),
    .C1(net5109),
    .B1(_02843_),
    .A1(_02840_),
    .Y(_02844_),
    .A2(_02841_));
 sg13g2_a22oi_1 _11372_ (.Y(_02845_),
    .B1(net4733),
    .B2(_02844_),
    .A2(net4737),
    .A1(\m_sys._m_core_io_b_mem_wdata[8] ));
 sg13g2_o21ai_1 _11373_ (.B1(_02845_),
    .Y(_00172_),
    .A1(net1799),
    .A2(net4786));
 sg13g2_a21oi_1 _11374_ (.A1(net5200),
    .A2(_02441_),
    .Y(_02846_),
    .B1(net5218));
 sg13g2_o21ai_1 _11375_ (.B1(_02846_),
    .Y(_02847_),
    .A1(net5200),
    .A2(\m_sys.m_core.m_gpr._GEN[233] ));
 sg13g2_a221oi_1 _11376_ (.B2(\m_sys.m_core.m_gpr._GEN[169] ),
    .C1(net5210),
    .B1(net5112),
    .A1(\m_sys.m_core.m_gpr._GEN[137] ),
    .Y(_02848_),
    .A2(net5157));
 sg13g2_mux2_1 _11377_ (.A0(\m_sys.m_core.m_gpr._GEN[73] ),
    .A1(\m_sys.m_core.m_gpr._GEN[105] ),
    .S(net5335),
    .X(_02849_));
 sg13g2_a22oi_1 _11378_ (.Y(_02850_),
    .B1(_02849_),
    .B2(net5343),
    .A2(net5112),
    .A1(\m_sys.m_core.m_gpr._GEN[41] ));
 sg13g2_a221oi_1 _11379_ (.B2(net5211),
    .C1(net5108),
    .B1(_02850_),
    .A1(_02847_),
    .Y(_02851_),
    .A2(_02848_));
 sg13g2_a22oi_1 _11380_ (.Y(_02852_),
    .B1(net4733),
    .B2(_02851_),
    .A2(net4736),
    .A1(\m_sys._m_core_io_b_mem_wdata[9] ));
 sg13g2_o21ai_1 _11381_ (.B1(_02852_),
    .Y(_00173_),
    .A1(net2471),
    .A2(net4786));
 sg13g2_mux2_1 _11382_ (.A0(\m_sys.m_core.m_gpr._GEN[202] ),
    .A1(\m_sys.m_core.m_gpr._GEN[234] ),
    .S(net5334),
    .X(_02853_));
 sg13g2_nand2_1 _11383_ (.Y(_02854_),
    .A(\m_sys.m_core.m_gpr._GEN[138] ),
    .B(net5153));
 sg13g2_a221oi_1 _11384_ (.B2(net5343),
    .C1(net5210),
    .B1(_02853_),
    .A1(\m_sys.m_core.m_gpr._GEN[170] ),
    .Y(_02855_),
    .A2(net5112));
 sg13g2_mux2_1 _11385_ (.A0(\m_sys.m_core.m_gpr._GEN[74] ),
    .A1(\m_sys.m_core.m_gpr._GEN[106] ),
    .S(net5332),
    .X(_02856_));
 sg13g2_a22oi_1 _11386_ (.Y(_02857_),
    .B1(_02856_),
    .B2(net5343),
    .A2(net5112),
    .A1(\m_sys.m_core.m_gpr._GEN[42] ));
 sg13g2_a221oi_1 _11387_ (.B2(net5210),
    .C1(net5107),
    .B1(_02857_),
    .A1(_02854_),
    .Y(_02858_),
    .A2(_02855_));
 sg13g2_a22oi_1 _11388_ (.Y(_02859_),
    .B1(net4733),
    .B2(_02858_),
    .A2(net4736),
    .A1(\m_sys._m_core_io_b_mem_wdata[10] ));
 sg13g2_o21ai_1 _11389_ (.B1(_02859_),
    .Y(_00174_),
    .A1(net1655),
    .A2(net4786));
 sg13g2_nor2_1 _11390_ (.A(net5204),
    .B(\m_sys.m_core.m_gpr._GEN[235] ),
    .Y(_02860_));
 sg13g2_o21ai_1 _11391_ (.B1(net5346),
    .Y(_02861_),
    .A1(net5336),
    .A2(\m_sys.m_core.m_gpr._GEN[203] ));
 sg13g2_a221oi_1 _11392_ (.B2(\m_sys.m_core.m_gpr._GEN[171] ),
    .C1(net5214),
    .B1(net5115),
    .A1(\m_sys.m_core.m_gpr._GEN[139] ),
    .Y(_02862_),
    .A2(net5155));
 sg13g2_o21ai_1 _11393_ (.B1(_02862_),
    .Y(_02863_),
    .A1(_02860_),
    .A2(_02861_));
 sg13g2_nor2_1 _11394_ (.A(net5336),
    .B(\m_sys.m_core.m_gpr._GEN[75] ),
    .Y(_02864_));
 sg13g2_o21ai_1 _11395_ (.B1(net5346),
    .Y(_02865_),
    .A1(net5204),
    .A2(\m_sys.m_core.m_gpr._GEN[107] ));
 sg13g2_a21oi_1 _11396_ (.A1(\m_sys.m_core.m_gpr._GEN[43] ),
    .A2(net5115),
    .Y(_02866_),
    .B1(net5351));
 sg13g2_o21ai_1 _11397_ (.B1(_02866_),
    .Y(_02867_),
    .A1(_02864_),
    .A2(_02865_));
 sg13g2_nand3_1 _11398_ (.B(_02863_),
    .C(_02867_),
    .A(net5105),
    .Y(_02868_));
 sg13g2_nor2_1 _11399_ (.A(net4732),
    .B(_02868_),
    .Y(_02869_));
 sg13g2_a21oi_1 _11400_ (.A1(net3166),
    .A2(net4736),
    .Y(_02870_),
    .B1(_02869_));
 sg13g2_mux2_1 _11401_ (.A0(_00018_),
    .A1(_00078_),
    .S(net5102),
    .X(_02871_));
 sg13g2_o21ai_1 _11402_ (.B1(_02870_),
    .Y(_00175_),
    .A1(net4786),
    .A2(_02871_));
 sg13g2_nor2_1 _11403_ (.A(net5202),
    .B(\m_sys.m_core.m_gpr._GEN[236] ),
    .Y(_02872_));
 sg13g2_o21ai_1 _11404_ (.B1(net5345),
    .Y(_02873_),
    .A1(net5337),
    .A2(\m_sys.m_core.m_gpr._GEN[204] ));
 sg13g2_a221oi_1 _11405_ (.B2(\m_sys.m_core.m_gpr._GEN[172] ),
    .C1(net5213),
    .B1(net5114),
    .A1(\m_sys.m_core.m_gpr._GEN[140] ),
    .Y(_02874_),
    .A2(net5156));
 sg13g2_o21ai_1 _11406_ (.B1(_02874_),
    .Y(_02875_),
    .A1(_02872_),
    .A2(_02873_));
 sg13g2_nor2_1 _11407_ (.A(net5337),
    .B(\m_sys.m_core.m_gpr._GEN[76] ),
    .Y(_02876_));
 sg13g2_o21ai_1 _11408_ (.B1(net5345),
    .Y(_02877_),
    .A1(net5202),
    .A2(\m_sys.m_core.m_gpr._GEN[108] ));
 sg13g2_a21oi_1 _11409_ (.A1(\m_sys.m_core.m_gpr._GEN[44] ),
    .A2(net5114),
    .Y(_02878_),
    .B1(net5352));
 sg13g2_o21ai_1 _11410_ (.B1(_02878_),
    .Y(_02879_),
    .A1(_02876_),
    .A2(_02877_));
 sg13g2_nand3_1 _11411_ (.B(_02875_),
    .C(_02879_),
    .A(net5105),
    .Y(_02880_));
 sg13g2_nor2_1 _11412_ (.A(net4732),
    .B(_02880_),
    .Y(_02881_));
 sg13g2_a21oi_1 _11413_ (.A1(\m_sys._m_core_io_b_mem_wdata[12] ),
    .A2(net4737),
    .Y(_02882_),
    .B1(_02881_));
 sg13g2_or2_1 _11414_ (.X(_02883_),
    .B(net4788),
    .A(_00080_));
 sg13g2_nand2b_1 _11415_ (.Y(_02884_),
    .B(_00080_),
    .A_N(net5103));
 sg13g2_nand2b_2 _11416_ (.Y(_02885_),
    .B(_02884_),
    .A_N(net4788));
 sg13g2_a21oi_1 _11417_ (.A1(net3289),
    .A2(net5103),
    .Y(_02886_),
    .B1(_02885_));
 sg13g2_nand2b_1 _11418_ (.Y(_00176_),
    .B(_02882_),
    .A_N(_02886_));
 sg13g2_mux2_1 _11419_ (.A0(\m_sys.m_core.m_gpr._GEN[205] ),
    .A1(\m_sys.m_core.m_gpr._GEN[237] ),
    .S(net5336),
    .X(_02887_));
 sg13g2_nand2_1 _11420_ (.Y(_02888_),
    .A(\m_sys.m_core.m_gpr._GEN[141] ),
    .B(net5155));
 sg13g2_a221oi_1 _11421_ (.B2(net5346),
    .C1(net5214),
    .B1(_02887_),
    .A1(\m_sys.m_core.m_gpr._GEN[173] ),
    .Y(_02889_),
    .A2(net5115));
 sg13g2_mux2_1 _11422_ (.A0(\m_sys.m_core.m_gpr._GEN[77] ),
    .A1(\m_sys.m_core.m_gpr._GEN[109] ),
    .S(net5336),
    .X(_02890_));
 sg13g2_a22oi_1 _11423_ (.Y(_02891_),
    .B1(_02890_),
    .B2(net5346),
    .A2(net5115),
    .A1(\m_sys.m_core.m_gpr._GEN[45] ));
 sg13g2_a22oi_1 _11424_ (.Y(_02892_),
    .B1(_02891_),
    .B2(net5214),
    .A2(_02889_),
    .A1(_02888_));
 sg13g2_nand2_2 _11425_ (.Y(_02893_),
    .A(net5106),
    .B(_02892_));
 sg13g2_nor2_1 _11426_ (.A(net4732),
    .B(_02893_),
    .Y(_02894_));
 sg13g2_a21oi_1 _11427_ (.A1(net3093),
    .A2(net4737),
    .Y(_02895_),
    .B1(_02894_));
 sg13g2_a21oi_1 _11428_ (.A1(_00081_),
    .A2(net5103),
    .Y(_02896_),
    .B1(_02885_));
 sg13g2_nand2b_1 _11429_ (.Y(_00177_),
    .B(_02895_),
    .A_N(_02896_));
 sg13g2_mux2_1 _11430_ (.A0(\m_sys.m_core.m_gpr._GEN[206] ),
    .A1(\m_sys.m_core.m_gpr._GEN[238] ),
    .S(net5338),
    .X(_02897_));
 sg13g2_nand2_1 _11431_ (.Y(_02898_),
    .A(\m_sys.m_core.m_gpr._GEN[142] ),
    .B(net5155));
 sg13g2_a221oi_1 _11432_ (.B2(net5348),
    .C1(net5216),
    .B1(_02897_),
    .A1(\m_sys.m_core.m_gpr._GEN[174] ),
    .Y(_02899_),
    .A2(net5116));
 sg13g2_mux2_1 _11433_ (.A0(\m_sys.m_core.m_gpr._GEN[78] ),
    .A1(\m_sys.m_core.m_gpr._GEN[110] ),
    .S(net5338),
    .X(_02900_));
 sg13g2_a22oi_1 _11434_ (.Y(_02901_),
    .B1(_02900_),
    .B2(net5348),
    .A2(net5116),
    .A1(\m_sys.m_core.m_gpr._GEN[46] ));
 sg13g2_a22oi_1 _11435_ (.Y(_02902_),
    .B1(_02901_),
    .B2(net5216),
    .A2(_02899_),
    .A1(_02898_));
 sg13g2_nand2_2 _11436_ (.Y(_02903_),
    .A(net5105),
    .B(_02902_));
 sg13g2_nor2_1 _11437_ (.A(net4732),
    .B(_02903_),
    .Y(_02904_));
 sg13g2_a21oi_1 _11438_ (.A1(net3156),
    .A2(net4737),
    .Y(_02905_),
    .B1(_02904_));
 sg13g2_a21oi_1 _11439_ (.A1(_00026_),
    .A2(net5103),
    .Y(_02906_),
    .B1(_02885_));
 sg13g2_nand2b_1 _11440_ (.Y(_00178_),
    .B(_02905_),
    .A_N(_02906_));
 sg13g2_nor2_1 _11441_ (.A(net5206),
    .B(\m_sys.m_core.m_gpr._GEN[239] ),
    .Y(_02907_));
 sg13g2_o21ai_1 _11442_ (.B1(net5349),
    .Y(_02908_),
    .A1(net5338),
    .A2(\m_sys.m_core.m_gpr._GEN[207] ));
 sg13g2_a221oi_1 _11443_ (.B2(\m_sys.m_core.m_gpr._GEN[175] ),
    .C1(net5216),
    .B1(net5118),
    .A1(\m_sys.m_core.m_gpr._GEN[143] ),
    .Y(_02909_),
    .A2(net5156));
 sg13g2_o21ai_1 _11444_ (.B1(_02909_),
    .Y(_02910_),
    .A1(_02907_),
    .A2(_02908_));
 sg13g2_nor2_1 _11445_ (.A(net5338),
    .B(\m_sys.m_core.m_gpr._GEN[79] ),
    .Y(_02911_));
 sg13g2_o21ai_1 _11446_ (.B1(net5348),
    .Y(_02912_),
    .A1(net5206),
    .A2(\m_sys.m_core.m_gpr._GEN[111] ));
 sg13g2_a21oi_1 _11447_ (.A1(\m_sys.m_core.m_gpr._GEN[47] ),
    .A2(net5116),
    .Y(_02913_),
    .B1(net5352));
 sg13g2_o21ai_1 _11448_ (.B1(_02913_),
    .Y(_02914_),
    .A1(_02911_),
    .A2(_02912_));
 sg13g2_nand3_1 _11449_ (.B(_02910_),
    .C(_02914_),
    .A(net5106),
    .Y(_02915_));
 sg13g2_nor2_1 _11450_ (.A(net4731),
    .B(_02915_),
    .Y(_02916_));
 sg13g2_a21oi_1 _11451_ (.A1(net3226),
    .A2(net4739),
    .Y(_02917_),
    .B1(_02916_));
 sg13g2_a21oi_1 _11452_ (.A1(_00082_),
    .A2(net5104),
    .Y(_02918_),
    .B1(_02885_));
 sg13g2_nand2b_1 _11453_ (.Y(_00179_),
    .B(_02917_),
    .A_N(_02918_));
 sg13g2_nor2_1 _11454_ (.A(net5205),
    .B(\m_sys.m_core.m_gpr._GEN[240] ),
    .Y(_02919_));
 sg13g2_o21ai_1 _11455_ (.B1(net5348),
    .Y(_02920_),
    .A1(net5338),
    .A2(\m_sys.m_core.m_gpr._GEN[208] ));
 sg13g2_a221oi_1 _11456_ (.B2(\m_sys.m_core.m_gpr._GEN[176] ),
    .C1(net5216),
    .B1(net5116),
    .A1(\m_sys.m_core.m_gpr._GEN[144] ),
    .Y(_02921_),
    .A2(net5157));
 sg13g2_o21ai_1 _11457_ (.B1(_02921_),
    .Y(_02922_),
    .A1(_02919_),
    .A2(_02920_));
 sg13g2_nor2_1 _11458_ (.A(net5338),
    .B(\m_sys.m_core.m_gpr._GEN[80] ),
    .Y(_02923_));
 sg13g2_o21ai_1 _11459_ (.B1(net5348),
    .Y(_02924_),
    .A1(net5206),
    .A2(\m_sys.m_core.m_gpr._GEN[112] ));
 sg13g2_a21oi_1 _11460_ (.A1(\m_sys.m_core.m_gpr._GEN[48] ),
    .A2(net5116),
    .Y(_02925_),
    .B1(\m_sys.m_core._m_decoder_io_o_rs2[2] ));
 sg13g2_o21ai_1 _11461_ (.B1(_02925_),
    .Y(_02926_),
    .A1(_02923_),
    .A2(_02924_));
 sg13g2_nand3_1 _11462_ (.B(_02922_),
    .C(_02926_),
    .A(net5105),
    .Y(_02927_));
 sg13g2_nor2_1 _11463_ (.A(net4732),
    .B(_02927_),
    .Y(_02928_));
 sg13g2_a21oi_1 _11464_ (.A1(\m_sys._m_core_io_b_mem_wdata[16] ),
    .A2(net4738),
    .Y(_02929_),
    .B1(_02928_));
 sg13g2_a21oi_1 _11465_ (.A1(net2990),
    .A2(net5104),
    .Y(_02930_),
    .B1(_02885_));
 sg13g2_nand2b_1 _11466_ (.Y(_00180_),
    .B(_02929_),
    .A_N(_02930_));
 sg13g2_nor2_1 _11467_ (.A(net5206),
    .B(\m_sys.m_core.m_gpr._GEN[241] ),
    .Y(_02931_));
 sg13g2_o21ai_1 _11468_ (.B1(net5348),
    .Y(_02932_),
    .A1(net5338),
    .A2(\m_sys.m_core.m_gpr._GEN[209] ));
 sg13g2_a221oi_1 _11469_ (.B2(\m_sys.m_core.m_gpr._GEN[177] ),
    .C1(net5216),
    .B1(net5116),
    .A1(\m_sys.m_core.m_gpr._GEN[145] ),
    .Y(_02933_),
    .A2(net5156));
 sg13g2_o21ai_1 _11470_ (.B1(_02933_),
    .Y(_02934_),
    .A1(_02931_),
    .A2(_02932_));
 sg13g2_nor2_1 _11471_ (.A(net5338),
    .B(\m_sys.m_core.m_gpr._GEN[81] ),
    .Y(_02935_));
 sg13g2_o21ai_1 _11472_ (.B1(net5348),
    .Y(_02936_),
    .A1(net5206),
    .A2(\m_sys.m_core.m_gpr._GEN[113] ));
 sg13g2_a21oi_1 _11473_ (.A1(\m_sys.m_core.m_gpr._GEN[49] ),
    .A2(net5116),
    .Y(_02937_),
    .B1(net5351));
 sg13g2_o21ai_1 _11474_ (.B1(_02937_),
    .Y(_02938_),
    .A1(_02935_),
    .A2(_02936_));
 sg13g2_nand3_1 _11475_ (.B(_02934_),
    .C(_02938_),
    .A(net5105),
    .Y(_02939_));
 sg13g2_nor2_1 _11476_ (.A(net4731),
    .B(_02939_),
    .Y(_02940_));
 sg13g2_a21oi_1 _11477_ (.A1(\m_sys._m_core_io_b_mem_wdata[17] ),
    .A2(_02759_),
    .Y(_02941_),
    .B1(_02940_));
 sg13g2_a21oi_1 _11478_ (.A1(net3377),
    .A2(net5104),
    .Y(_02942_),
    .B1(_02885_));
 sg13g2_nand2b_1 _11479_ (.Y(_00181_),
    .B(_02941_),
    .A_N(_02942_));
 sg13g2_nor2_1 _11480_ (.A(net5205),
    .B(\m_sys.m_core.m_gpr._GEN[242] ),
    .Y(_02943_));
 sg13g2_o21ai_1 _11481_ (.B1(net5347),
    .Y(_02944_),
    .A1(net5339),
    .A2(\m_sys.m_core.m_gpr._GEN[210] ));
 sg13g2_a221oi_1 _11482_ (.B2(\m_sys.m_core.m_gpr._GEN[178] ),
    .C1(net5215),
    .B1(net5117),
    .A1(\m_sys.m_core.m_gpr._GEN[146] ),
    .Y(_02945_),
    .A2(net5156));
 sg13g2_o21ai_1 _11483_ (.B1(_02945_),
    .Y(_02946_),
    .A1(_02943_),
    .A2(_02944_));
 sg13g2_nor2_1 _11484_ (.A(net5339),
    .B(\m_sys.m_core.m_gpr._GEN[82] ),
    .Y(_02947_));
 sg13g2_o21ai_1 _11485_ (.B1(net5347),
    .Y(_02948_),
    .A1(net5205),
    .A2(\m_sys.m_core.m_gpr._GEN[114] ));
 sg13g2_a21oi_1 _11486_ (.A1(\m_sys.m_core.m_gpr._GEN[50] ),
    .A2(net5117),
    .Y(_02949_),
    .B1(net5351));
 sg13g2_o21ai_1 _11487_ (.B1(_02949_),
    .Y(_02950_),
    .A1(_02947_),
    .A2(_02948_));
 sg13g2_nand3_1 _11488_ (.B(_02946_),
    .C(_02950_),
    .A(net5106),
    .Y(_02951_));
 sg13g2_nor2_1 _11489_ (.A(net4731),
    .B(_02951_),
    .Y(_02952_));
 sg13g2_a21oi_1 _11490_ (.A1(\m_sys._m_core_io_b_mem_wdata[18] ),
    .A2(net4738),
    .Y(_02953_),
    .B1(_02952_));
 sg13g2_a21oi_1 _11491_ (.A1(net3240),
    .A2(net5104),
    .Y(_02954_),
    .B1(_02885_));
 sg13g2_nand2b_1 _11492_ (.Y(_00182_),
    .B(_02953_),
    .A_N(_02954_));
 sg13g2_mux2_1 _11493_ (.A0(\m_sys.m_core.m_gpr._GEN[211] ),
    .A1(\m_sys.m_core.m_gpr._GEN[243] ),
    .S(net5340),
    .X(_02955_));
 sg13g2_nand2_1 _11494_ (.Y(_02956_),
    .A(\m_sys.m_core.m_gpr._GEN[147] ),
    .B(net5156));
 sg13g2_a221oi_1 _11495_ (.B2(net5349),
    .C1(net5215),
    .B1(_02955_),
    .A1(\m_sys.m_core.m_gpr._GEN[179] ),
    .Y(_02957_),
    .A2(net5118));
 sg13g2_mux2_1 _11496_ (.A0(\m_sys.m_core.m_gpr._GEN[83] ),
    .A1(\m_sys.m_core.m_gpr._GEN[115] ),
    .S(net5340),
    .X(_02958_));
 sg13g2_a22oi_1 _11497_ (.Y(_02959_),
    .B1(_02958_),
    .B2(net5348),
    .A2(net5116),
    .A1(\m_sys.m_core.m_gpr._GEN[51] ));
 sg13g2_a22oi_1 _11498_ (.Y(_02960_),
    .B1(_02959_),
    .B2(net5215),
    .A2(_02957_),
    .A1(_02956_));
 sg13g2_nand2_2 _11499_ (.Y(_02961_),
    .A(net5105),
    .B(_02960_));
 sg13g2_nor2_1 _11500_ (.A(net4731),
    .B(_02961_),
    .Y(_02962_));
 sg13g2_a21oi_1 _11501_ (.A1(\m_sys._m_core_io_b_mem_wdata[19] ),
    .A2(net4738),
    .Y(_02963_),
    .B1(_02962_));
 sg13g2_a21oi_1 _11502_ (.A1(net3394),
    .A2(net5104),
    .Y(_02964_),
    .B1(_02885_));
 sg13g2_nand2b_1 _11503_ (.Y(_00183_),
    .B(_02963_),
    .A_N(_02964_));
 sg13g2_nand2_1 _11504_ (.Y(_02965_),
    .A(net3276),
    .B(net4739));
 sg13g2_mux2_1 _11505_ (.A0(\m_sys.m_core.m_gpr._GEN[212] ),
    .A1(\m_sys.m_core.m_gpr._GEN[244] ),
    .S(net5337),
    .X(_02966_));
 sg13g2_nand2_1 _11506_ (.Y(_02967_),
    .A(\m_sys.m_core.m_gpr._GEN[148] ),
    .B(net5155));
 sg13g2_a221oi_1 _11507_ (.B2(net5345),
    .C1(net5213),
    .B1(_02966_),
    .A1(\m_sys.m_core.m_gpr._GEN[180] ),
    .Y(_02968_),
    .A2(net5114));
 sg13g2_mux2_1 _11508_ (.A0(\m_sys.m_core.m_gpr._GEN[84] ),
    .A1(\m_sys.m_core.m_gpr._GEN[116] ),
    .S(net5337),
    .X(_02969_));
 sg13g2_a22oi_1 _11509_ (.Y(_02970_),
    .B1(_02969_),
    .B2(net5345),
    .A2(net5114),
    .A1(\m_sys.m_core.m_gpr._GEN[52] ));
 sg13g2_a221oi_1 _11510_ (.B2(net5213),
    .C1(net5109),
    .B1(_02970_),
    .A1(_02967_),
    .Y(_02971_),
    .A2(_02968_));
 sg13g2_nand2_1 _11511_ (.Y(_02972_),
    .A(_02776_),
    .B(_02971_));
 sg13g2_nand3_1 _11512_ (.B(_02965_),
    .C(_02972_),
    .A(net4730),
    .Y(_00184_));
 sg13g2_a21oi_1 _11513_ (.A1(net5203),
    .A2(_02453_),
    .Y(_02973_),
    .B1(net5219));
 sg13g2_o21ai_1 _11514_ (.B1(_02973_),
    .Y(_02974_),
    .A1(net5203),
    .A2(\m_sys.m_core.m_gpr._GEN[245] ));
 sg13g2_a221oi_1 _11515_ (.B2(\m_sys.m_core.m_gpr._GEN[181] ),
    .C1(net5212),
    .B1(net5118),
    .A1(\m_sys.m_core.m_gpr._GEN[149] ),
    .Y(_02975_),
    .A2(net5155));
 sg13g2_mux2_1 _11516_ (.A0(\m_sys.m_core.m_gpr._GEN[85] ),
    .A1(\m_sys.m_core.m_gpr._GEN[117] ),
    .S(net5337),
    .X(_02976_));
 sg13g2_a22oi_1 _11517_ (.Y(_02977_),
    .B1(_02976_),
    .B2(net5345),
    .A2(net5118),
    .A1(\m_sys.m_core.m_gpr._GEN[53] ));
 sg13g2_a221oi_1 _11518_ (.B2(net5212),
    .C1(net5109),
    .B1(_02977_),
    .A1(_02974_),
    .Y(_02978_),
    .A2(_02975_));
 sg13g2_a22oi_1 _11519_ (.Y(_02979_),
    .B1(net4734),
    .B2(_02978_),
    .A2(net4738),
    .A1(net3322));
 sg13g2_nand2_1 _11520_ (.Y(_00185_),
    .A(net4730),
    .B(_02979_));
 sg13g2_nand2_1 _11521_ (.Y(_02980_),
    .A(net3399),
    .B(net4738));
 sg13g2_a21oi_1 _11522_ (.A1(net5203),
    .A2(_02454_),
    .Y(_02981_),
    .B1(net5219));
 sg13g2_o21ai_1 _11523_ (.B1(_02981_),
    .Y(_02982_),
    .A1(net5203),
    .A2(\m_sys.m_core.m_gpr._GEN[246] ));
 sg13g2_a221oi_1 _11524_ (.B2(\m_sys.m_core.m_gpr._GEN[182] ),
    .C1(net5212),
    .B1(net5114),
    .A1(\m_sys.m_core.m_gpr._GEN[150] ),
    .Y(_02983_),
    .A2(net5155));
 sg13g2_mux2_1 _11525_ (.A0(\m_sys.m_core.m_gpr._GEN[86] ),
    .A1(\m_sys.m_core.m_gpr._GEN[118] ),
    .S(net5337),
    .X(_02984_));
 sg13g2_a22oi_1 _11526_ (.Y(_02985_),
    .B1(_02984_),
    .B2(net5345),
    .A2(net5114),
    .A1(\m_sys.m_core.m_gpr._GEN[54] ));
 sg13g2_a221oi_1 _11527_ (.B2(net5213),
    .C1(net5109),
    .B1(_02985_),
    .A1(_02982_),
    .Y(_02986_),
    .A2(_02983_));
 sg13g2_nand2_1 _11528_ (.Y(_02987_),
    .A(_02776_),
    .B(_02986_));
 sg13g2_nand3_1 _11529_ (.B(_02980_),
    .C(_02987_),
    .A(net4730),
    .Y(_00186_));
 sg13g2_nor2_1 _11530_ (.A(net5201),
    .B(\m_sys.m_core.m_gpr._GEN[247] ),
    .Y(_02988_));
 sg13g2_o21ai_1 _11531_ (.B1(net5345),
    .Y(_02989_),
    .A1(net5337),
    .A2(\m_sys.m_core.m_gpr._GEN[215] ));
 sg13g2_a221oi_1 _11532_ (.B2(\m_sys.m_core.m_gpr._GEN[183] ),
    .C1(net5213),
    .B1(net5114),
    .A1(\m_sys.m_core.m_gpr._GEN[151] ),
    .Y(_02990_),
    .A2(net5155));
 sg13g2_o21ai_1 _11533_ (.B1(_02990_),
    .Y(_02991_),
    .A1(_02988_),
    .A2(_02989_));
 sg13g2_nor2_1 _11534_ (.A(net5337),
    .B(\m_sys.m_core.m_gpr._GEN[87] ),
    .Y(_02992_));
 sg13g2_o21ai_1 _11535_ (.B1(net5345),
    .Y(_02993_),
    .A1(net5201),
    .A2(\m_sys.m_core.m_gpr._GEN[119] ));
 sg13g2_a21oi_1 _11536_ (.A1(\m_sys.m_core.m_gpr._GEN[55] ),
    .A2(net5114),
    .Y(_02994_),
    .B1(net5351));
 sg13g2_o21ai_1 _11537_ (.B1(_02994_),
    .Y(_02995_),
    .A1(_02992_),
    .A2(_02993_));
 sg13g2_nand3_1 _11538_ (.B(_02991_),
    .C(_02995_),
    .A(net5105),
    .Y(_02996_));
 sg13g2_o21ai_1 _11539_ (.B1(net4729),
    .Y(_02997_),
    .A1(net4731),
    .A2(_02996_));
 sg13g2_a21o_1 _11540_ (.A2(net4738),
    .A1(net3384),
    .B1(_02997_),
    .X(_00187_));
 sg13g2_mux2_1 _11541_ (.A0(\m_sys.m_core.m_gpr._GEN[216] ),
    .A1(\m_sys.m_core.m_gpr._GEN[248] ),
    .S(net5333),
    .X(_02998_));
 sg13g2_nand2_1 _11542_ (.Y(_02999_),
    .A(\m_sys.m_core.m_gpr._GEN[152] ),
    .B(net5154));
 sg13g2_a221oi_1 _11543_ (.B2(net5341),
    .C1(net5209),
    .B1(_02998_),
    .A1(\m_sys.m_core.m_gpr._GEN[184] ),
    .Y(_03000_),
    .A2(net5111));
 sg13g2_mux2_1 _11544_ (.A0(\m_sys.m_core.m_gpr._GEN[88] ),
    .A1(\m_sys.m_core.m_gpr._GEN[120] ),
    .S(net5332),
    .X(_03001_));
 sg13g2_a22oi_1 _11545_ (.Y(_03002_),
    .B1(_03001_),
    .B2(net5341),
    .A2(net5111),
    .A1(\m_sys.m_core.m_gpr._GEN[56] ));
 sg13g2_a221oi_1 _11546_ (.B2(net5209),
    .C1(net5107),
    .B1(_03002_),
    .A1(_02999_),
    .Y(_03003_),
    .A2(_03000_));
 sg13g2_a22oi_1 _11547_ (.Y(_03004_),
    .B1(_02776_),
    .B2(_03003_),
    .A2(net4738),
    .A1(net3442));
 sg13g2_nand2_1 _11548_ (.Y(_00188_),
    .A(net4730),
    .B(_03004_));
 sg13g2_nor2_1 _11549_ (.A(net5204),
    .B(\m_sys.m_core.m_gpr._GEN[249] ),
    .Y(_03005_));
 sg13g2_o21ai_1 _11550_ (.B1(net5342),
    .Y(_03006_),
    .A1(net5333),
    .A2(\m_sys.m_core.m_gpr._GEN[217] ));
 sg13g2_a221oi_1 _11551_ (.B2(\m_sys.m_core.m_gpr._GEN[185] ),
    .C1(net5209),
    .B1(net5111),
    .A1(\m_sys.m_core.m_gpr._GEN[153] ),
    .Y(_03007_),
    .A2(net5154));
 sg13g2_o21ai_1 _11552_ (.B1(_03007_),
    .Y(_03008_),
    .A1(_03005_),
    .A2(_03006_));
 sg13g2_nor2_1 _11553_ (.A(net5336),
    .B(\m_sys.m_core.m_gpr._GEN[89] ),
    .Y(_03009_));
 sg13g2_o21ai_1 _11554_ (.B1(net5346),
    .Y(_03010_),
    .A1(net5204),
    .A2(\m_sys.m_core.m_gpr._GEN[121] ));
 sg13g2_a21oi_1 _11555_ (.A1(\m_sys.m_core.m_gpr._GEN[57] ),
    .A2(net5115),
    .Y(_03011_),
    .B1(net5351));
 sg13g2_o21ai_1 _11556_ (.B1(_03011_),
    .Y(_03012_),
    .A1(_03009_),
    .A2(_03010_));
 sg13g2_nand3_1 _11557_ (.B(_03008_),
    .C(_03012_),
    .A(net5106),
    .Y(_03013_));
 sg13g2_o21ai_1 _11558_ (.B1(net4729),
    .Y(_03014_),
    .A1(net4731),
    .A2(_03013_));
 sg13g2_a21o_1 _11559_ (.A2(net4739),
    .A1(net3371),
    .B1(_03014_),
    .X(_00189_));
 sg13g2_nand2_1 _11560_ (.Y(_03015_),
    .A(net3440),
    .B(net4739));
 sg13g2_mux2_1 _11561_ (.A0(\m_sys.m_core.m_gpr._GEN[218] ),
    .A1(\m_sys.m_core.m_gpr._GEN[250] ),
    .S(net5332),
    .X(_03016_));
 sg13g2_nand2_1 _11562_ (.Y(_03017_),
    .A(\m_sys.m_core.m_gpr._GEN[154] ),
    .B(net5154));
 sg13g2_a221oi_1 _11563_ (.B2(net5341),
    .C1(net5208),
    .B1(_03016_),
    .A1(\m_sys.m_core.m_gpr._GEN[186] ),
    .Y(_03018_),
    .A2(net5110));
 sg13g2_mux2_1 _11564_ (.A0(\m_sys.m_core.m_gpr._GEN[90] ),
    .A1(\m_sys.m_core.m_gpr._GEN[122] ),
    .S(net5332),
    .X(_03019_));
 sg13g2_a22oi_1 _11565_ (.Y(_03020_),
    .B1(_03019_),
    .B2(net5341),
    .A2(net5110),
    .A1(\m_sys.m_core.m_gpr._GEN[58] ));
 sg13g2_a221oi_1 _11566_ (.B2(net5208),
    .C1(net5107),
    .B1(_03020_),
    .A1(_03017_),
    .Y(_03021_),
    .A2(_03018_));
 sg13g2_nand2_1 _11567_ (.Y(_03022_),
    .A(net4734),
    .B(_03021_));
 sg13g2_nand3_1 _11568_ (.B(_03015_),
    .C(_03022_),
    .A(net4729),
    .Y(_00190_));
 sg13g2_nor2_1 _11569_ (.A(net5200),
    .B(\m_sys.m_core.m_gpr._GEN[251] ),
    .Y(_03023_));
 sg13g2_o21ai_1 _11570_ (.B1(net5342),
    .Y(_03024_),
    .A1(net5333),
    .A2(\m_sys.m_core.m_gpr._GEN[219] ));
 sg13g2_a221oi_1 _11571_ (.B2(\m_sys.m_core.m_gpr._GEN[187] ),
    .C1(net5209),
    .B1(net5110),
    .A1(\m_sys.m_core.m_gpr._GEN[155] ),
    .Y(_03025_),
    .A2(net5154));
 sg13g2_o21ai_1 _11572_ (.B1(_03025_),
    .Y(_03026_),
    .A1(_03023_),
    .A2(_03024_));
 sg13g2_a21oi_1 _11573_ (.A1(net5198),
    .A2(_02455_),
    .Y(_03027_),
    .B1(net5218));
 sg13g2_o21ai_1 _11574_ (.B1(_03027_),
    .Y(_03028_),
    .A1(net5198),
    .A2(\m_sys.m_core.m_gpr._GEN[123] ));
 sg13g2_a21oi_1 _11575_ (.A1(\m_sys.m_core.m_gpr._GEN[59] ),
    .A2(net5110),
    .Y(_03029_),
    .B1(net5352));
 sg13g2_a21oi_1 _11576_ (.A1(_03028_),
    .A2(_03029_),
    .Y(_03030_),
    .B1(net5107));
 sg13g2_nand2_2 _11577_ (.Y(_03031_),
    .A(_03026_),
    .B(_03030_));
 sg13g2_o21ai_1 _11578_ (.B1(net4729),
    .Y(_03032_),
    .A1(net4731),
    .A2(_03031_));
 sg13g2_a21o_1 _11579_ (.A2(net4738),
    .A1(net3389),
    .B1(_03032_),
    .X(_00191_));
 sg13g2_nand2_1 _11580_ (.Y(_03033_),
    .A(net3429),
    .B(net4739));
 sg13g2_mux2_1 _11581_ (.A0(\m_sys.m_core.m_gpr._GEN[220] ),
    .A1(\m_sys.m_core.m_gpr._GEN[252] ),
    .S(net5333),
    .X(_03034_));
 sg13g2_nand2_1 _11582_ (.Y(_03035_),
    .A(\m_sys.m_core.m_gpr._GEN[156] ),
    .B(net5154));
 sg13g2_a221oi_1 _11583_ (.B2(net5342),
    .C1(net5209),
    .B1(_03034_),
    .A1(\m_sys.m_core.m_gpr._GEN[188] ),
    .Y(_03036_),
    .A2(net5111));
 sg13g2_mux2_1 _11584_ (.A0(\m_sys.m_core.m_gpr._GEN[92] ),
    .A1(\m_sys.m_core.m_gpr._GEN[124] ),
    .S(net5333),
    .X(_03037_));
 sg13g2_a22oi_1 _11585_ (.Y(_03038_),
    .B1(_03037_),
    .B2(net5342),
    .A2(net5111),
    .A1(\m_sys.m_core.m_gpr._GEN[60] ));
 sg13g2_a221oi_1 _11586_ (.B2(net5209),
    .C1(net5107),
    .B1(_03038_),
    .A1(_03035_),
    .Y(_03039_),
    .A2(_03036_));
 sg13g2_nand2_1 _11587_ (.Y(_03040_),
    .A(net4734),
    .B(_03039_));
 sg13g2_nand3_1 _11588_ (.B(_03033_),
    .C(_03040_),
    .A(net4729),
    .Y(_00192_));
 sg13g2_mux2_1 _11589_ (.A0(\m_sys.m_core.m_gpr._GEN[221] ),
    .A1(\m_sys.m_core.m_gpr._GEN[253] ),
    .S(net5336),
    .X(_03041_));
 sg13g2_nand2_1 _11590_ (.Y(_03042_),
    .A(\m_sys.m_core.m_gpr._GEN[157] ),
    .B(net5155));
 sg13g2_a221oi_1 _11591_ (.B2(net5346),
    .C1(net5214),
    .B1(_03041_),
    .A1(\m_sys.m_core.m_gpr._GEN[189] ),
    .Y(_03043_),
    .A2(net5115));
 sg13g2_mux2_1 _11592_ (.A0(\m_sys.m_core.m_gpr._GEN[93] ),
    .A1(\m_sys.m_core.m_gpr._GEN[125] ),
    .S(net5336),
    .X(_03044_));
 sg13g2_a22oi_1 _11593_ (.Y(_03045_),
    .B1(_03044_),
    .B2(net5346),
    .A2(net5115),
    .A1(\m_sys.m_core.m_gpr._GEN[61] ));
 sg13g2_a22oi_1 _11594_ (.Y(_03046_),
    .B1(_03045_),
    .B2(net5214),
    .A2(_03043_),
    .A1(_03042_));
 sg13g2_nand2_2 _11595_ (.Y(_03047_),
    .A(net5105),
    .B(_03046_));
 sg13g2_o21ai_1 _11596_ (.B1(net4729),
    .Y(_03048_),
    .A1(net4731),
    .A2(_03047_));
 sg13g2_a21o_1 _11597_ (.A2(net4739),
    .A1(net3331),
    .B1(_03048_),
    .X(_00193_));
 sg13g2_nand2_1 _11598_ (.Y(_03049_),
    .A(net3411),
    .B(net4737));
 sg13g2_a21oi_1 _11599_ (.A1(net5198),
    .A2(_02456_),
    .Y(_03050_),
    .B1(net5218));
 sg13g2_o21ai_1 _11600_ (.B1(_03050_),
    .Y(_03051_),
    .A1(net5198),
    .A2(\m_sys.m_core.m_gpr._GEN[254] ));
 sg13g2_a221oi_1 _11601_ (.B2(\m_sys.m_core.m_gpr._GEN[190] ),
    .C1(net5208),
    .B1(net5110),
    .A1(\m_sys.m_core.m_gpr._GEN[158] ),
    .Y(_03052_),
    .A2(net5154));
 sg13g2_mux2_1 _11602_ (.A0(\m_sys.m_core.m_gpr._GEN[94] ),
    .A1(\m_sys.m_core.m_gpr._GEN[126] ),
    .S(net5332),
    .X(_03053_));
 sg13g2_a22oi_1 _11603_ (.Y(_03054_),
    .B1(_03053_),
    .B2(net5341),
    .A2(net5110),
    .A1(\m_sys.m_core.m_gpr._GEN[62] ));
 sg13g2_a221oi_1 _11604_ (.B2(net5208),
    .C1(net5107),
    .B1(_03054_),
    .A1(_03051_),
    .Y(_03055_),
    .A2(_03052_));
 sg13g2_nand2_1 _11605_ (.Y(_03056_),
    .A(net4734),
    .B(_03055_));
 sg13g2_nand3_1 _11606_ (.B(_03049_),
    .C(_03056_),
    .A(net4729),
    .Y(_00194_));
 sg13g2_a21oi_1 _11607_ (.A1(net5198),
    .A2(_02457_),
    .Y(_03057_),
    .B1(net5218));
 sg13g2_o21ai_1 _11608_ (.B1(_03057_),
    .Y(_03058_),
    .A1(net5198),
    .A2(\m_sys.m_core.m_gpr._GEN[255] ));
 sg13g2_a221oi_1 _11609_ (.B2(\m_sys.m_core.m_gpr._GEN[191] ),
    .C1(net5208),
    .B1(net5110),
    .A1(\m_sys.m_core.m_gpr._GEN[159] ),
    .Y(_03059_),
    .A2(net5154));
 sg13g2_mux2_1 _11610_ (.A0(\m_sys.m_core.m_gpr._GEN[95] ),
    .A1(\m_sys.m_core.m_gpr._GEN[127] ),
    .S(net5332),
    .X(_03060_));
 sg13g2_a22oi_1 _11611_ (.Y(_03061_),
    .B1(_03060_),
    .B2(net5341),
    .A2(net5110),
    .A1(\m_sys.m_core.m_gpr._GEN[63] ));
 sg13g2_a221oi_1 _11612_ (.B2(net5208),
    .C1(net5107),
    .B1(_03061_),
    .A1(_03058_),
    .Y(_03062_),
    .A2(_03059_));
 sg13g2_a22oi_1 _11613_ (.Y(_03063_),
    .B1(net4734),
    .B2(_03062_),
    .A2(net4739),
    .A1(net3330));
 sg13g2_nand2_1 _11614_ (.Y(_00195_),
    .A(net4729),
    .B(_03063_));
 sg13g2_a21oi_2 _11615_ (.B1(_02634_),
    .Y(_03064_),
    .A2(net5309),
    .A1(\m_sys.m_core.m_fsm.r_cstate[0] ));
 sg13g2_a21o_2 _11616_ (.A2(net5309),
    .A1(net5242),
    .B1(_02634_),
    .X(_03065_));
 sg13g2_nor3_1 _11617_ (.A(net5242),
    .B(net5232),
    .C(_02634_),
    .Y(_03066_));
 sg13g2_nand3_1 _11618_ (.B(\m_sys.m_core.m_fsm.r_cstate[2] ),
    .C(_02751_),
    .A(net5309),
    .Y(_03067_));
 sg13g2_nor2_2 _11619_ (.A(_02488_),
    .B(net5093),
    .Y(_03068_));
 sg13g2_nand4_1 _11620_ (.B(\m_sys.m_core.m_fsm.r_cstate[2] ),
    .C(\m_sys.m_core.r_ctrl_bru_pc_rel ),
    .A(net5309),
    .Y(_03069_),
    .D(_02751_));
 sg13g2_mux2_2 _11621_ (.A0(\m_sys._m_core_io_b_mem_wdata[30] ),
    .A1(\m_sys.m_core.m_bru.io_i_s1[30] ),
    .S(net5082),
    .X(_03070_));
 sg13g2_nand2_1 _11622_ (.Y(_03071_),
    .A(\m_sys.m_core.m_bru.io_i_s2[30] ),
    .B(net5083));
 sg13g2_nor2b_1 _11623_ (.A(_03070_),
    .B_N(_03071_),
    .Y(_03072_));
 sg13g2_nand2_2 _11624_ (.Y(_03073_),
    .A(\m_sys.m_core.m_bru.io_i_s2[15] ),
    .B(net5084));
 sg13g2_nor2_1 _11625_ (.A(_00082_),
    .B(_03073_),
    .Y(_03074_));
 sg13g2_mux2_2 _11626_ (.A0(_00096_),
    .A1(_00082_),
    .S(net5084),
    .X(_03075_));
 sg13g2_mux2_1 _11627_ (.A0(_02492_),
    .A1(_02446_),
    .S(net5082),
    .X(_03076_));
 sg13g2_and2_1 _11628_ (.A(_03073_),
    .B(_03075_),
    .X(_03077_));
 sg13g2_mux2_2 _11629_ (.A0(_00082_),
    .A1(_03076_),
    .S(_03073_),
    .X(_03078_));
 sg13g2_nor2b_1 _11630_ (.A(_00026_),
    .B_N(net5082),
    .Y(_03079_));
 sg13g2_nand2_2 _11631_ (.Y(_03080_),
    .A(\m_sys.m_core.m_bru.io_i_s2[14] ),
    .B(net5092));
 sg13g2_nand2_2 _11632_ (.Y(_03081_),
    .A(\m_sys.m_core.m_bru.io_i_s2[14] ),
    .B(_03079_));
 sg13g2_mux2_2 _11633_ (.A0(_00097_),
    .A1(_00026_),
    .S(net5082),
    .X(_03082_));
 sg13g2_nand2_1 _11634_ (.Y(_03083_),
    .A(_03080_),
    .B(_03082_));
 sg13g2_a22oi_1 _11635_ (.Y(_03084_),
    .B1(_03080_),
    .B2(_03082_),
    .A2(_03079_),
    .A1(\m_sys.m_core.m_bru.io_i_s2[14] ));
 sg13g2_nand2_1 _11636_ (.Y(_03085_),
    .A(_03081_),
    .B(_03083_));
 sg13g2_nand2_1 _11637_ (.Y(_03086_),
    .A(_03078_),
    .B(_03084_));
 sg13g2_nor2b_1 _11638_ (.A(_00081_),
    .B_N(net5077),
    .Y(_03087_));
 sg13g2_mux2_2 _11639_ (.A0(_00098_),
    .A1(_00081_),
    .S(net5078),
    .X(_03088_));
 sg13g2_nand2_1 _11640_ (.Y(_03089_),
    .A(\m_sys.m_core.m_bru.io_i_s2[13] ),
    .B(net5082));
 sg13g2_nand2_1 _11641_ (.Y(_03090_),
    .A(_03088_),
    .B(_03089_));
 sg13g2_a22oi_1 _11642_ (.Y(_03091_),
    .B1(_03088_),
    .B2(_03089_),
    .A2(_03087_),
    .A1(\m_sys.m_core.m_bru.io_i_s2[13] ));
 sg13g2_nor2b_1 _11643_ (.A(_00079_),
    .B_N(net5077),
    .Y(_03092_));
 sg13g2_nand2_1 _11644_ (.Y(_03093_),
    .A(\m_sys.m_core.m_bru.io_i_s2[12] ),
    .B(net5077));
 sg13g2_nor2_1 _11645_ (.A(_00079_),
    .B(_03093_),
    .Y(_03094_));
 sg13g2_mux2_2 _11646_ (.A0(_00099_),
    .A1(_00079_),
    .S(net5078),
    .X(_03095_));
 sg13g2_nand2_1 _11647_ (.Y(_03096_),
    .A(_03093_),
    .B(_03095_));
 sg13g2_a22oi_1 _11648_ (.Y(_03097_),
    .B1(_03093_),
    .B2(_03095_),
    .A2(_03092_),
    .A1(\m_sys.m_core.m_bru.io_i_s2[12] ));
 sg13g2_and2_1 _11649_ (.A(_03091_),
    .B(_03097_),
    .X(_03098_));
 sg13g2_nor2b_1 _11650_ (.A(_03086_),
    .B_N(_03098_),
    .Y(_03099_));
 sg13g2_mux2_2 _11651_ (.A0(_02409_),
    .A1(net5229),
    .S(net5078),
    .X(_03100_));
 sg13g2_mux2_2 _11652_ (.A0(_00103_),
    .A1(_00102_),
    .S(net5078),
    .X(_03101_));
 sg13g2_nand2b_1 _11653_ (.Y(_03102_),
    .B(_03101_),
    .A_N(_03100_));
 sg13g2_or2_2 _11654_ (.X(_03103_),
    .B(_03101_),
    .A(_03100_));
 sg13g2_xnor2_1 _11655_ (.Y(_03104_),
    .A(_03100_),
    .B(_03101_));
 sg13g2_mux2_2 _11656_ (.A0(_00017_),
    .A1(_00100_),
    .S(net5081),
    .X(_03105_));
 sg13g2_mux2_2 _11657_ (.A0(\m_sys._m_core_io_b_mem_wdata[11] ),
    .A1(\m_sys.m_core.m_bru.io_i_s1[11] ),
    .S(net5077),
    .X(_03106_));
 sg13g2_nand2b_1 _11658_ (.Y(_03107_),
    .B(_03106_),
    .A_N(_03105_));
 sg13g2_nand2_1 _11659_ (.Y(_03108_),
    .A(_03105_),
    .B(_03106_));
 sg13g2_xor2_1 _11660_ (.B(_03106_),
    .A(_03105_),
    .X(_03109_));
 sg13g2_nor2_1 _11661_ (.A(_03104_),
    .B(_03109_),
    .Y(_03110_));
 sg13g2_mux2_2 _11662_ (.A0(\m_sys._m_core_io_b_mem_wdata[7] ),
    .A1(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[0] ),
    .S(net5079),
    .X(_03111_));
 sg13g2_mux2_2 _11663_ (.A0(_00019_),
    .A1(_00110_),
    .S(net5075),
    .X(_03112_));
 sg13g2_nand2b_2 _11664_ (.Y(_03113_),
    .B(_03111_),
    .A_N(_03112_));
 sg13g2_nor2b_1 _11665_ (.A(_03111_),
    .B_N(_03112_),
    .Y(_03114_));
 sg13g2_nand2b_2 _11666_ (.Y(_03115_),
    .B(_03112_),
    .A_N(_03111_));
 sg13g2_mux2_1 _11667_ (.A0(_00023_),
    .A1(_00111_),
    .S(net5076),
    .X(_03116_));
 sg13g2_mux2_2 _11668_ (.A0(\m_sys._m_core_io_b_mem_wdata[6] ),
    .A1(\m_sys.m_core.m_bru.io_i_s1[6] ),
    .S(net5079),
    .X(_03117_));
 sg13g2_inv_1 _11669_ (.Y(_03118_),
    .A(_03117_));
 sg13g2_nand2b_2 _11670_ (.Y(_03119_),
    .B(_03117_),
    .A_N(_03116_));
 sg13g2_o21ai_1 _11671_ (.B1(_03113_),
    .Y(_03120_),
    .A1(_03114_),
    .A2(_03119_));
 sg13g2_nand2_1 _11672_ (.Y(_03121_),
    .A(_02462_),
    .B(net5074));
 sg13g2_mux2_2 _11673_ (.A0(\m_sys.m_core.m_bru.io_i_pc[3] ),
    .A1(\m_sys.m_core.m_bru.io_i_s2[3] ),
    .S(net5074),
    .X(_03122_));
 sg13g2_o21ai_1 _11674_ (.B1(_03121_),
    .Y(_03123_),
    .A1(\m_sys.m_core.m_bru.io_i_pc[3] ),
    .A2(net5074));
 sg13g2_mux2_2 _11675_ (.A0(_00116_),
    .A1(_00012_),
    .S(net5075),
    .X(_03124_));
 sg13g2_nor2b_1 _11676_ (.A(net4948),
    .B_N(_03124_),
    .Y(_03125_));
 sg13g2_nor2_1 _11677_ (.A(net4785),
    .B(_03124_),
    .Y(_03126_));
 sg13g2_mux2_2 _11678_ (.A0(\m_sys.m_core.m_bru.io_i_pc[2] ),
    .A1(\m_sys.m_core.m_bru.io_i_s2[2] ),
    .S(net5074),
    .X(_03127_));
 sg13g2_mux2_1 _11679_ (.A0(_02363_),
    .A1(_02463_),
    .S(net5074),
    .X(_03128_));
 sg13g2_mux2_2 _11680_ (.A0(_00117_),
    .A1(_00010_),
    .S(net5076),
    .X(_03129_));
 sg13g2_nor2_1 _11681_ (.A(net4936),
    .B(_03129_),
    .Y(_03130_));
 sg13g2_mux2_1 _11682_ (.A0(_02323_),
    .A1(_02461_),
    .S(net5076),
    .X(_03131_));
 sg13g2_mux2_1 _11683_ (.A0(\m_sys.m_core._m_bru_io_o_res[1] ),
    .A1(\m_sys.m_core.m_bru.io_i_s2[1] ),
    .S(net5076),
    .X(_03132_));
 sg13g2_mux2_2 _11684_ (.A0(_00120_),
    .A1(_00119_),
    .S(net5080),
    .X(_03133_));
 sg13g2_nor2_1 _11685_ (.A(net4927),
    .B(_03133_),
    .Y(_03134_));
 sg13g2_nand2b_1 _11686_ (.Y(_03135_),
    .B(net4913),
    .A_N(_03133_));
 sg13g2_mux2_1 _11687_ (.A0(_02324_),
    .A1(_02460_),
    .S(net5076),
    .X(_03136_));
 sg13g2_mux2_1 _11688_ (.A0(\m_sys.m_core._m_bru_io_o_res[0] ),
    .A1(\m_sys.m_core.m_bru.io_i_s2[0] ),
    .S(net5076),
    .X(_03137_));
 sg13g2_mux2_2 _11689_ (.A0(_00027_),
    .A1(_00089_),
    .S(net5080),
    .X(_03138_));
 sg13g2_nor2_1 _11690_ (.A(net4904),
    .B(_03138_),
    .Y(_03139_));
 sg13g2_nand2b_1 _11691_ (.Y(_03140_),
    .B(net4897),
    .A_N(_03138_));
 sg13g2_and2_1 _11692_ (.A(net4927),
    .B(_03133_),
    .X(_03141_));
 sg13g2_a21oi_1 _11693_ (.A1(_03135_),
    .A2(_03140_),
    .Y(_03142_),
    .B1(_03141_));
 sg13g2_nor2_1 _11694_ (.A(net4945),
    .B(_03129_),
    .Y(_03143_));
 sg13g2_nand2b_1 _11695_ (.Y(_03144_),
    .B(net4936),
    .A_N(_03129_));
 sg13g2_nand2_1 _11696_ (.Y(_03145_),
    .A(net4945),
    .B(_03129_));
 sg13g2_nand2_1 _11697_ (.Y(_03146_),
    .A(_03144_),
    .B(_03145_));
 sg13g2_a221oi_1 _11698_ (.B2(_03145_),
    .C1(_03141_),
    .B1(_03144_),
    .A1(_03135_),
    .Y(_03147_),
    .A2(_03140_));
 sg13g2_nor2_1 _11699_ (.A(_03130_),
    .B(_03147_),
    .Y(_03148_));
 sg13g2_nor3_1 _11700_ (.A(_03126_),
    .B(_03130_),
    .C(_03147_),
    .Y(_03149_));
 sg13g2_nor2_1 _11701_ (.A(_03125_),
    .B(_03149_),
    .Y(_03150_));
 sg13g2_mux2_2 _11702_ (.A0(\m_sys.m_core.m_bru.io_i_pc[4] ),
    .A1(\m_sys.m_core.m_bru.io_i_s2[4] ),
    .S(net5074),
    .X(_03151_));
 sg13g2_mux2_1 _11703_ (.A0(_02362_),
    .A1(_02466_),
    .S(net5074),
    .X(_03152_));
 sg13g2_mux2_2 _11704_ (.A0(_00115_),
    .A1(_00008_),
    .S(net5079),
    .X(_03153_));
 sg13g2_nor2_1 _11705_ (.A(net4894),
    .B(_03153_),
    .Y(_03154_));
 sg13g2_or2_1 _11706_ (.X(_03155_),
    .B(_03153_),
    .A(net4894));
 sg13g2_nand2_1 _11707_ (.Y(_03156_),
    .A(net4894),
    .B(_03153_));
 sg13g2_nand2_2 _11708_ (.Y(_03157_),
    .A(_03155_),
    .B(_03156_));
 sg13g2_mux2_2 _11709_ (.A0(_00021_),
    .A1(_00113_),
    .S(net5075),
    .X(_03158_));
 sg13g2_mux2_2 _11710_ (.A0(\m_sys._m_core_io_b_mem_wdata[5] ),
    .A1(net5319),
    .S(net5079),
    .X(_03159_));
 sg13g2_nand2b_1 _11711_ (.Y(_03160_),
    .B(_03159_),
    .A_N(_03158_));
 sg13g2_nand2b_1 _11712_ (.Y(_03161_),
    .B(_03158_),
    .A_N(_03159_));
 sg13g2_inv_1 _11713_ (.Y(_03162_),
    .A(_03161_));
 sg13g2_nand2_2 _11714_ (.Y(_03163_),
    .A(_03160_),
    .B(_03161_));
 sg13g2_nor2_1 _11715_ (.A(_03157_),
    .B(_03163_),
    .Y(_03164_));
 sg13g2_or4_1 _11716_ (.A(_03125_),
    .B(_03149_),
    .C(_03157_),
    .D(_03163_),
    .X(_03165_));
 sg13g2_a21oi_1 _11717_ (.A1(_03155_),
    .A2(_03160_),
    .Y(_03166_),
    .B1(_03162_));
 sg13g2_a21oi_1 _11718_ (.A1(_03150_),
    .A2(_03164_),
    .Y(_03167_),
    .B1(_03166_));
 sg13g2_nor2_1 _11719_ (.A(_03120_),
    .B(_03166_),
    .Y(_03168_));
 sg13g2_nor2b_1 _11720_ (.A(_03117_),
    .B_N(_03116_),
    .Y(_03169_));
 sg13g2_inv_1 _11721_ (.Y(_03170_),
    .A(_03169_));
 sg13g2_a221oi_1 _11722_ (.B2(_03113_),
    .C1(_03114_),
    .B1(_03169_),
    .A1(_03165_),
    .Y(_03171_),
    .A2(_03168_));
 sg13g2_mux2_2 _11723_ (.A0(\m_sys._m_core_io_b_mem_wdata[8] ),
    .A1(net5320),
    .S(net5077),
    .X(_03172_));
 sg13g2_mux2_2 _11724_ (.A0(_00109_),
    .A1(_00108_),
    .S(net5076),
    .X(_03173_));
 sg13g2_nand2b_2 _11725_ (.Y(_03174_),
    .B(_03172_),
    .A_N(_03173_));
 sg13g2_nand2b_1 _11726_ (.Y(_03175_),
    .B(_03173_),
    .A_N(_03172_));
 sg13g2_nand2_2 _11727_ (.Y(_03176_),
    .A(_03174_),
    .B(_03175_));
 sg13g2_mux2_2 _11728_ (.A0(\m_sys._m_core_io_b_mem_wdata[9] ),
    .A1(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[2] ),
    .S(net5077),
    .X(_03177_));
 sg13g2_mux2_2 _11729_ (.A0(_00106_),
    .A1(_00105_),
    .S(net5079),
    .X(_03178_));
 sg13g2_nand2_1 _11730_ (.Y(_03179_),
    .A(_03177_),
    .B(_03178_));
 sg13g2_nand2b_1 _11731_ (.Y(_03180_),
    .B(_03177_),
    .A_N(_03178_));
 sg13g2_xor2_1 _11732_ (.B(_03178_),
    .A(_03177_),
    .X(_03181_));
 sg13g2_nor2_2 _11733_ (.A(_03176_),
    .B(_03181_),
    .Y(_03182_));
 sg13g2_o21ai_1 _11734_ (.B1(_03180_),
    .Y(_03183_),
    .A1(_03174_),
    .A2(_03181_));
 sg13g2_a21oi_2 _11735_ (.B1(_03183_),
    .Y(_03184_),
    .A2(_03182_),
    .A1(_03171_));
 sg13g2_a22oi_1 _11736_ (.Y(_03185_),
    .B1(_03090_),
    .B2(_03094_),
    .A2(_03087_),
    .A1(\m_sys.m_core.m_bru.io_i_s2[13] ));
 sg13g2_nor2_1 _11737_ (.A(_03077_),
    .B(_03081_),
    .Y(_03186_));
 sg13g2_nor2_1 _11738_ (.A(_03074_),
    .B(_03186_),
    .Y(_03187_));
 sg13g2_o21ai_1 _11739_ (.B1(_03187_),
    .Y(_03188_),
    .A1(_03086_),
    .A2(_03185_));
 sg13g2_o21ai_1 _11740_ (.B1(_03107_),
    .Y(_03189_),
    .A1(_03103_),
    .A2(_03109_));
 sg13g2_and3_1 _11741_ (.X(_03190_),
    .A(_03099_),
    .B(_03110_),
    .C(_03182_));
 sg13g2_a21o_1 _11742_ (.A2(_03183_),
    .A1(_03110_),
    .B1(_03189_),
    .X(_03191_));
 sg13g2_a21o_1 _11743_ (.A2(_03191_),
    .A1(_03099_),
    .B1(_03188_),
    .X(_03192_));
 sg13g2_a21oi_2 _11744_ (.B1(_03192_),
    .Y(_03193_),
    .A2(_03190_),
    .A1(_03171_));
 sg13g2_a21o_2 _11745_ (.A2(_03190_),
    .A1(_03171_),
    .B1(_03192_),
    .X(_03194_));
 sg13g2_nand2_1 _11746_ (.Y(_03195_),
    .A(\m_sys.m_core.m_bru.io_i_s2[23] ),
    .B(net5088));
 sg13g2_nand3_1 _11747_ (.B(\m_sys.m_core.m_bru.io_i_s2[23] ),
    .C(net5087),
    .A(\m_sys.m_core.m_bru.io_i_s1[23] ),
    .Y(_03196_));
 sg13g2_mux2_2 _11748_ (.A0(\m_sys._m_core_io_b_mem_wdata[23] ),
    .A1(\m_sys.m_core.m_bru.io_i_s1[23] ),
    .S(net5088),
    .X(_03197_));
 sg13g2_nand2b_1 _11749_ (.Y(_03198_),
    .B(_03195_),
    .A_N(_03197_));
 sg13g2_inv_1 _11750_ (.Y(_03199_),
    .A(_03198_));
 sg13g2_nand2_2 _11751_ (.Y(_03200_),
    .A(_03196_),
    .B(_03198_));
 sg13g2_mux2_2 _11752_ (.A0(\m_sys._m_core_io_b_mem_wdata[22] ),
    .A1(net5352),
    .S(net5088),
    .X(_03201_));
 sg13g2_nand2_1 _11753_ (.Y(_03202_),
    .A(\m_sys.m_core.m_bru.io_i_s2[22] ),
    .B(net5087));
 sg13g2_nand2b_2 _11754_ (.Y(_03203_),
    .B(_03202_),
    .A_N(_03201_));
 sg13g2_inv_1 _11755_ (.Y(_03204_),
    .A(_03203_));
 sg13g2_nand3_1 _11756_ (.B(\m_sys.m_core.m_bru.io_i_s2[22] ),
    .C(net5087),
    .A(net5352),
    .Y(_03205_));
 sg13g2_and2_1 _11757_ (.A(_03203_),
    .B(_03205_),
    .X(_03206_));
 sg13g2_nand2_2 _11758_ (.Y(_03207_),
    .A(_03203_),
    .B(_03205_));
 sg13g2_nand2_1 _11759_ (.Y(_03208_),
    .A(\m_sys.m_core.m_bru.io_i_s2[20] ),
    .B(net5087));
 sg13g2_nor2_2 _11760_ (.A(_00078_),
    .B(_03208_),
    .Y(_03209_));
 sg13g2_mux2_2 _11761_ (.A0(_00091_),
    .A1(_00078_),
    .S(net5086),
    .X(_03210_));
 sg13g2_and2_1 _11762_ (.A(_03208_),
    .B(_03210_),
    .X(_03211_));
 sg13g2_nor2_2 _11763_ (.A(_03209_),
    .B(_03211_),
    .Y(_03212_));
 sg13g2_nand2_2 _11764_ (.Y(_03213_),
    .A(\m_sys.m_core.m_bru.io_i_s2[21] ),
    .B(net5087));
 sg13g2_nor2_2 _11765_ (.A(_00065_),
    .B(_03213_),
    .Y(_03214_));
 sg13g2_mux2_2 _11766_ (.A0(_00090_),
    .A1(_00065_),
    .S(net5087),
    .X(_03215_));
 sg13g2_inv_1 _11767_ (.Y(_03216_),
    .A(_03215_));
 sg13g2_nand2_1 _11768_ (.Y(_03217_),
    .A(_03213_),
    .B(_03215_));
 sg13g2_nor2b_2 _11769_ (.A(_03214_),
    .B_N(_03217_),
    .Y(_03218_));
 sg13g2_nand2b_1 _11770_ (.Y(_03219_),
    .B(_03217_),
    .A_N(_03214_));
 sg13g2_and2_1 _11771_ (.A(_03212_),
    .B(_03218_),
    .X(_03220_));
 sg13g2_nand4_1 _11772_ (.B(_03198_),
    .C(_03206_),
    .A(_03196_),
    .Y(_03221_),
    .D(_03220_));
 sg13g2_nor2b_1 _11773_ (.A(_00086_),
    .B_N(net5090),
    .Y(_03222_));
 sg13g2_mux2_2 _11774_ (.A0(_00092_),
    .A1(_00086_),
    .S(net5090),
    .X(_03223_));
 sg13g2_nand2_2 _11775_ (.Y(_03224_),
    .A(\m_sys.m_core.m_bru.io_i_s2[19] ),
    .B(net5090));
 sg13g2_a22oi_1 _11776_ (.Y(_03225_),
    .B1(_03223_),
    .B2(_03224_),
    .A2(_03222_),
    .A1(\m_sys.m_core.m_bru.io_i_s2[19] ));
 sg13g2_inv_1 _11777_ (.Y(_03226_),
    .A(_03225_));
 sg13g2_nand2_1 _11778_ (.Y(_03227_),
    .A(\m_sys.m_core.m_bru.io_i_s2[18] ),
    .B(net5090));
 sg13g2_nand3_1 _11779_ (.B(\m_sys.m_core.m_bru.io_i_s2[18] ),
    .C(net5089),
    .A(_02451_),
    .Y(_03228_));
 sg13g2_nor2_1 _11780_ (.A(_00093_),
    .B(net5090),
    .Y(_03229_));
 sg13g2_a21oi_2 _11781_ (.B1(_03229_),
    .Y(_03230_),
    .A2(net5089),
    .A1(_02451_));
 sg13g2_mux2_1 _11782_ (.A0(_02491_),
    .A1(_02451_),
    .S(net5090),
    .X(_03231_));
 sg13g2_nor2b_1 _11783_ (.A(_03231_),
    .B_N(_03227_),
    .Y(_03232_));
 sg13g2_mux2_2 _11784_ (.A0(_00085_),
    .A1(_03231_),
    .S(_03227_),
    .X(_03233_));
 sg13g2_and2_1 _11785_ (.A(_03225_),
    .B(_03233_),
    .X(_03234_));
 sg13g2_nand2_1 _11786_ (.Y(_03235_),
    .A(\m_sys.m_core.m_bru.io_i_s2[16] ),
    .B(net5089));
 sg13g2_or2_1 _11787_ (.X(_03236_),
    .B(_03235_),
    .A(_00083_));
 sg13g2_mux2_2 _11788_ (.A0(_00095_),
    .A1(_00083_),
    .S(net5089),
    .X(_03237_));
 sg13g2_nand2_1 _11789_ (.Y(_03238_),
    .A(_03235_),
    .B(_03237_));
 sg13g2_nand2_2 _11790_ (.Y(_03239_),
    .A(_03236_),
    .B(_03238_));
 sg13g2_nand2_1 _11791_ (.Y(_03240_),
    .A(\m_sys.m_core.m_bru.io_i_s2[17] ),
    .B(net5089));
 sg13g2_nor2_1 _11792_ (.A(_00084_),
    .B(_03240_),
    .Y(_03241_));
 sg13g2_inv_1 _11793_ (.Y(_03242_),
    .A(_03241_));
 sg13g2_mux2_2 _11794_ (.A0(_00094_),
    .A1(_00084_),
    .S(net5089),
    .X(_03243_));
 sg13g2_and2_1 _11795_ (.A(_03240_),
    .B(_03243_),
    .X(_03244_));
 sg13g2_mux2_2 _11796_ (.A0(_02449_),
    .A1(_03243_),
    .S(_03240_),
    .X(_03245_));
 sg13g2_nor2_1 _11797_ (.A(_03239_),
    .B(_03245_),
    .Y(_03246_));
 sg13g2_nand2_1 _11798_ (.Y(_03247_),
    .A(_03234_),
    .B(_03246_));
 sg13g2_nor2_1 _11799_ (.A(_03221_),
    .B(_03247_),
    .Y(_03248_));
 sg13g2_o21ai_1 _11800_ (.B1(_03242_),
    .Y(_03249_),
    .A1(_03236_),
    .A2(_03244_));
 sg13g2_a21oi_1 _11801_ (.A1(_03223_),
    .A2(_03224_),
    .Y(_03250_),
    .B1(_03228_));
 sg13g2_a221oi_1 _11802_ (.B2(_03249_),
    .C1(_03250_),
    .B1(_03234_),
    .A1(\m_sys.m_core.m_bru.io_i_s2[19] ),
    .Y(_03251_),
    .A2(_03222_));
 sg13g2_a21oi_1 _11803_ (.A1(_03196_),
    .A2(_03205_),
    .Y(_03252_),
    .B1(_03199_));
 sg13g2_a21oi_1 _11804_ (.A1(_03209_),
    .A2(_03217_),
    .Y(_03253_),
    .B1(_03214_));
 sg13g2_nor3_1 _11805_ (.A(_03200_),
    .B(_03207_),
    .C(_03253_),
    .Y(_03254_));
 sg13g2_nor2_1 _11806_ (.A(_03252_),
    .B(_03254_),
    .Y(_03255_));
 sg13g2_o21ai_1 _11807_ (.B1(_03255_),
    .Y(_03256_),
    .A1(_03221_),
    .A2(_03251_));
 sg13g2_a21oi_1 _11808_ (.A1(_03194_),
    .A2(_03248_),
    .Y(_03257_),
    .B1(_03256_));
 sg13g2_a21o_1 _11809_ (.A2(_03248_),
    .A1(_03194_),
    .B1(_03256_),
    .X(_03258_));
 sg13g2_nand2_1 _11810_ (.Y(_03259_),
    .A(\m_sys.m_core.m_bru.io_i_s2[27] ),
    .B(net5086));
 sg13g2_nand3_1 _11811_ (.B(\m_sys.m_core.m_bru.io_i_s2[27] ),
    .C(net5085),
    .A(\m_sys.m_core.m_bru.io_i_s1[27] ),
    .Y(_03260_));
 sg13g2_mux2_2 _11812_ (.A0(\m_sys._m_core_io_b_mem_wdata[27] ),
    .A1(\m_sys.m_core.m_bru.io_i_s1[27] ),
    .S(net5085),
    .X(_03261_));
 sg13g2_a21o_1 _11813_ (.A2(net5085),
    .A1(\m_sys.m_core.m_bru.io_i_s2[27] ),
    .B1(_03261_),
    .X(_03262_));
 sg13g2_and2_1 _11814_ (.A(_03260_),
    .B(_03262_),
    .X(_03263_));
 sg13g2_nand2_1 _11815_ (.Y(_03264_),
    .A(_03260_),
    .B(_03262_));
 sg13g2_nor2_2 _11816_ (.A(_02479_),
    .B(_03068_),
    .Y(_03265_));
 sg13g2_nand2_1 _11817_ (.Y(_03266_),
    .A(\m_sys.m_core.m_bru.io_i_s1[26] ),
    .B(_03265_));
 sg13g2_mux2_2 _11818_ (.A0(\m_sys._m_core_io_b_mem_wdata[26] ),
    .A1(\m_sys.m_core.m_bru.io_i_s1[26] ),
    .S(net5085),
    .X(_03267_));
 sg13g2_inv_2 _11819_ (.Y(_03268_),
    .A(_03267_));
 sg13g2_nor2_1 _11820_ (.A(_03265_),
    .B(_03267_),
    .Y(_03269_));
 sg13g2_o21ai_1 _11821_ (.B1(_03266_),
    .Y(_03270_),
    .A1(_03265_),
    .A2(_03267_));
 sg13g2_nor2_1 _11822_ (.A(_03264_),
    .B(_03270_),
    .Y(_03271_));
 sg13g2_nand2_1 _11823_ (.Y(_03272_),
    .A(\m_sys.m_core.m_bru.io_i_s2[25] ),
    .B(net5085));
 sg13g2_nand3_1 _11824_ (.B(\m_sys.m_core.m_bru.io_i_s2[25] ),
    .C(net5086),
    .A(\m_sys.m_core.m_bru.io_i_s1[25] ),
    .Y(_03273_));
 sg13g2_mux2_2 _11825_ (.A0(\m_sys._m_core_io_b_mem_wdata[25] ),
    .A1(\m_sys.m_core.m_bru.io_i_s1[25] ),
    .S(net5085),
    .X(_03274_));
 sg13g2_a21oi_1 _11826_ (.A1(\m_sys.m_core.m_bru.io_i_s2[25] ),
    .A2(net5085),
    .Y(_03275_),
    .B1(_03274_));
 sg13g2_inv_1 _11827_ (.Y(_03276_),
    .A(_03275_));
 sg13g2_nand2_2 _11828_ (.Y(_03277_),
    .A(_03273_),
    .B(_03276_));
 sg13g2_nand3_1 _11829_ (.B(\m_sys.m_core.m_bru.io_i_s2[24] ),
    .C(net5088),
    .A(\m_sys.m_core.m_bru.io_i_s1[24] ),
    .Y(_03278_));
 sg13g2_mux2_2 _11830_ (.A0(\m_sys._m_core_io_b_mem_wdata[24] ),
    .A1(\m_sys.m_core.m_bru.io_i_s1[24] ),
    .S(net5086),
    .X(_03279_));
 sg13g2_inv_2 _11831_ (.Y(_03280_),
    .A(_03279_));
 sg13g2_o21ai_1 _11832_ (.B1(_03280_),
    .Y(_03281_),
    .A1(_02480_),
    .A2(_03068_));
 sg13g2_nand2_2 _11833_ (.Y(_03282_),
    .A(_03278_),
    .B(_03281_));
 sg13g2_nor2_1 _11834_ (.A(_03277_),
    .B(_03282_),
    .Y(_03283_));
 sg13g2_nand2_1 _11835_ (.Y(_03284_),
    .A(_03271_),
    .B(_03283_));
 sg13g2_a21oi_1 _11836_ (.A1(_03273_),
    .A2(_03278_),
    .Y(_03285_),
    .B1(_03275_));
 sg13g2_nand2_1 _11837_ (.Y(_03286_),
    .A(_03260_),
    .B(_03266_));
 sg13g2_a22oi_1 _11838_ (.Y(_03287_),
    .B1(_03286_),
    .B2(_03262_),
    .A2(_03285_),
    .A1(_03271_));
 sg13g2_o21ai_1 _11839_ (.B1(_03287_),
    .Y(_03288_),
    .A1(_03257_),
    .A2(_03284_));
 sg13g2_nand2_1 _11840_ (.Y(_03289_),
    .A(\m_sys.m_core.m_bru.io_i_s2[29] ),
    .B(net5084));
 sg13g2_nand3_1 _11841_ (.B(\m_sys.m_core.m_bru.io_i_s2[29] ),
    .C(net5084),
    .A(\m_sys.m_core.m_bru.io_i_s1[29] ),
    .Y(_03290_));
 sg13g2_mux2_2 _11842_ (.A0(\m_sys._m_core_io_b_mem_wdata[29] ),
    .A1(\m_sys.m_core.m_bru.io_i_s1[29] ),
    .S(net5083),
    .X(_03291_));
 sg13g2_a21o_1 _11843_ (.A2(net5083),
    .A1(\m_sys.m_core.m_bru.io_i_s2[29] ),
    .B1(_03291_),
    .X(_03292_));
 sg13g2_nand2_2 _11844_ (.Y(_03293_),
    .A(_03290_),
    .B(_03292_));
 sg13g2_nand3_1 _11845_ (.B(\m_sys.m_core.m_bru.io_i_s2[28] ),
    .C(net5084),
    .A(\m_sys.m_core.m_bru.io_i_s1[28] ),
    .Y(_03294_));
 sg13g2_mux2_2 _11846_ (.A0(\m_sys._m_core_io_b_mem_wdata[28] ),
    .A1(\m_sys.m_core.m_bru.io_i_s1[28] ),
    .S(net5083),
    .X(_03295_));
 sg13g2_inv_2 _11847_ (.Y(_03296_),
    .A(_03295_));
 sg13g2_o21ai_1 _11848_ (.B1(_03296_),
    .Y(_03297_),
    .A1(_02477_),
    .A2(_03068_));
 sg13g2_nand2_2 _11849_ (.Y(_03298_),
    .A(_03294_),
    .B(_03297_));
 sg13g2_nor2_1 _11850_ (.A(_03293_),
    .B(_03298_),
    .Y(_03299_));
 sg13g2_nand2_1 _11851_ (.Y(_03300_),
    .A(_03290_),
    .B(_03294_));
 sg13g2_a22oi_1 _11852_ (.Y(_03301_),
    .B1(_03300_),
    .B2(_03292_),
    .A2(_03299_),
    .A1(_03288_));
 sg13g2_nand3_1 _11853_ (.B(\m_sys.m_core.m_bru.io_i_s2[30] ),
    .C(net5083),
    .A(\m_sys.m_core.m_bru.io_i_s1[30] ),
    .Y(_03302_));
 sg13g2_o21ai_1 _11854_ (.B1(_03302_),
    .Y(_03303_),
    .A1(_03072_),
    .A2(_03301_));
 sg13g2_nor2b_2 _11855_ (.A(_03072_),
    .B_N(_03302_),
    .Y(_03304_));
 sg13g2_nand2_1 _11856_ (.Y(_03305_),
    .A(_03113_),
    .B(_03115_));
 sg13g2_mux2_2 _11857_ (.A0(_00112_),
    .A1(_00022_),
    .S(net5079),
    .X(_03306_));
 sg13g2_nand2_2 _11858_ (.Y(_03307_),
    .A(_03116_),
    .B(_03306_));
 sg13g2_nand2_1 _11859_ (.Y(_03308_),
    .A(_03119_),
    .B(_03307_));
 sg13g2_a22oi_1 _11860_ (.Y(_03309_),
    .B1(_03119_),
    .B2(_03307_),
    .A2(_03115_),
    .A1(_03113_));
 sg13g2_mux2_2 _11861_ (.A0(_00114_),
    .A1(_00020_),
    .S(net5079),
    .X(_03310_));
 sg13g2_mux2_1 _11862_ (.A0(_03159_),
    .A1(_03310_),
    .S(_03158_),
    .X(_03311_));
 sg13g2_xnor2_1 _11863_ (.Y(_03312_),
    .A(net4927),
    .B(_03133_));
 sg13g2_nand2_2 _11864_ (.Y(_03313_),
    .A(net4897),
    .B(_03138_));
 sg13g2_nor2_1 _11865_ (.A(net4913),
    .B(_03133_),
    .Y(_03314_));
 sg13g2_a21oi_1 _11866_ (.A1(_03312_),
    .A2(_03313_),
    .Y(_03315_),
    .B1(_03314_));
 sg13g2_a21o_1 _11867_ (.A2(_03313_),
    .A1(_03312_),
    .B1(_03314_),
    .X(_03316_));
 sg13g2_nand2_1 _11868_ (.Y(_03317_),
    .A(_00118_),
    .B(net5075));
 sg13g2_mux2_1 _11869_ (.A0(_02372_),
    .A1(_02495_),
    .S(net5075),
    .X(_03318_));
 sg13g2_o21ai_1 _11870_ (.B1(_03317_),
    .Y(_03319_),
    .A1(_02372_),
    .A2(net5074));
 sg13g2_mux2_1 _11871_ (.A0(net4936),
    .A1(net4887),
    .S(_03129_),
    .X(_03320_));
 sg13g2_nor2_1 _11872_ (.A(net4948),
    .B(_03124_),
    .Y(_03321_));
 sg13g2_xor2_1 _11873_ (.B(_03124_),
    .A(net4948),
    .X(_03322_));
 sg13g2_nor2b_1 _11874_ (.A(_03320_),
    .B_N(_03322_),
    .Y(_03323_));
 sg13g2_a221oi_1 _11875_ (.B2(_03316_),
    .C1(_03321_),
    .B1(_03323_),
    .A1(_03143_),
    .Y(_03324_),
    .A2(_03322_));
 sg13g2_nor2b_1 _11876_ (.A(_03324_),
    .B_N(_03157_),
    .Y(_03325_));
 sg13g2_nand3_1 _11877_ (.B(_03309_),
    .C(_03311_),
    .A(_03157_),
    .Y(_03326_));
 sg13g2_nor2_1 _11878_ (.A(_03151_),
    .B(_03153_),
    .Y(_03327_));
 sg13g2_and2_1 _11879_ (.A(_03158_),
    .B(_03159_),
    .X(_03328_));
 sg13g2_a21o_1 _11880_ (.A2(_03327_),
    .A1(_03311_),
    .B1(_03328_),
    .X(_03329_));
 sg13g2_nand2_1 _11881_ (.Y(_03330_),
    .A(_03116_),
    .B(_03117_));
 sg13g2_a21oi_1 _11882_ (.A1(_03113_),
    .A2(_03115_),
    .Y(_03331_),
    .B1(_03330_));
 sg13g2_a221oi_1 _11883_ (.B2(_03329_),
    .C1(_03331_),
    .B1(_03309_),
    .A1(_03111_),
    .Y(_03332_),
    .A2(_03112_));
 sg13g2_o21ai_1 _11884_ (.B1(_03332_),
    .Y(_03333_),
    .A1(_03324_),
    .A2(_03326_));
 sg13g2_or2_1 _11885_ (.X(_03334_),
    .B(_03097_),
    .A(_03091_));
 sg13g2_nor2_1 _11886_ (.A(_03078_),
    .B(_03084_),
    .Y(_03335_));
 sg13g2_nand2b_1 _11887_ (.Y(_03336_),
    .B(_03335_),
    .A_N(_03334_));
 sg13g2_nand2_1 _11888_ (.Y(_03337_),
    .A(_00016_),
    .B(net5081));
 sg13g2_o21ai_1 _11889_ (.B1(_03337_),
    .Y(_03338_),
    .A1(_02493_),
    .A2(net5077));
 sg13g2_mux4_1 _11890_ (.S0(_03105_),
    .A0(net5230),
    .A1(_02382_),
    .A2(_02410_),
    .A3(_02493_),
    .S1(_03068_),
    .X(_03339_));
 sg13g2_mux2_2 _11891_ (.A0(_00104_),
    .A1(_00070_),
    .S(net5077),
    .X(_03340_));
 sg13g2_nand2_1 _11892_ (.Y(_03341_),
    .A(_03101_),
    .B(_03340_));
 sg13g2_and2_1 _11893_ (.A(_03103_),
    .B(_03341_),
    .X(_03342_));
 sg13g2_a21oi_1 _11894_ (.A1(_03103_),
    .A2(_03341_),
    .Y(_03343_),
    .B1(_03339_));
 sg13g2_inv_1 _11895_ (.Y(_03344_),
    .A(_03343_));
 sg13g2_mux2_2 _11896_ (.A0(_00107_),
    .A1(_00068_),
    .S(net5079),
    .X(_03345_));
 sg13g2_nand2_1 _11897_ (.Y(_03346_),
    .A(_03178_),
    .B(_03345_));
 sg13g2_mux4_1 _11898_ (.S0(_03068_),
    .A0(net5228),
    .A1(_02408_),
    .A2(_02426_),
    .A3(_02494_),
    .S1(_03178_),
    .X(_03347_));
 sg13g2_nand2_1 _11899_ (.Y(_03348_),
    .A(_03180_),
    .B(_03346_));
 sg13g2_nand3_1 _11900_ (.B(_03343_),
    .C(_03348_),
    .A(_03176_),
    .Y(_03349_));
 sg13g2_nor2_1 _11901_ (.A(_03336_),
    .B(_03349_),
    .Y(_03350_));
 sg13g2_o21ai_1 _11902_ (.B1(_03108_),
    .Y(_03351_),
    .A1(_03102_),
    .A2(_03339_));
 sg13g2_nand2_1 _11903_ (.Y(_03352_),
    .A(_03172_),
    .B(_03173_));
 sg13g2_or2_1 _11904_ (.X(_03353_),
    .B(_03352_),
    .A(_03347_));
 sg13g2_o21ai_1 _11905_ (.B1(_03179_),
    .Y(_03354_),
    .A1(_03347_),
    .A2(_03352_));
 sg13g2_inv_1 _11906_ (.Y(_03355_),
    .A(_03354_));
 sg13g2_a21oi_1 _11907_ (.A1(_03343_),
    .A2(_03354_),
    .Y(_03356_),
    .B1(_03351_));
 sg13g2_a21o_1 _11908_ (.A2(net5082),
    .A1(\m_sys.m_core.m_bru.io_i_s2[12] ),
    .B1(_03095_),
    .X(_03357_));
 sg13g2_nand2b_1 _11909_ (.Y(_03358_),
    .B(_03089_),
    .A_N(_03088_));
 sg13g2_o21ai_1 _11910_ (.B1(_03358_),
    .Y(_03359_),
    .A1(_03091_),
    .A2(_03357_));
 sg13g2_a21oi_1 _11911_ (.A1(\m_sys.m_core.m_bru.io_i_s2[14] ),
    .A2(net5082),
    .Y(_03360_),
    .B1(_03082_));
 sg13g2_nor2b_1 _11912_ (.A(_03078_),
    .B_N(_03360_),
    .Y(_03361_));
 sg13g2_a221oi_1 _11913_ (.B2(_03359_),
    .C1(_03361_),
    .B1(_03335_),
    .A1(_03073_),
    .Y(_03362_),
    .A2(_03076_));
 sg13g2_o21ai_1 _11914_ (.B1(_03362_),
    .Y(_03363_),
    .A1(_03336_),
    .A2(_03356_));
 sg13g2_a21oi_2 _11915_ (.B1(_03363_),
    .Y(_03364_),
    .A2(_03350_),
    .A1(_03333_));
 sg13g2_nand2_1 _11916_ (.Y(_03365_),
    .A(_03200_),
    .B(_03207_));
 sg13g2_nor2_1 _11917_ (.A(_03225_),
    .B(_03233_),
    .Y(_03366_));
 sg13g2_nand2_1 _11918_ (.Y(_03367_),
    .A(_03239_),
    .B(_03245_));
 sg13g2_nand3_1 _11919_ (.B(_03245_),
    .C(_03366_),
    .A(_03239_),
    .Y(_03368_));
 sg13g2_or4_1 _11920_ (.A(_03212_),
    .B(_03218_),
    .C(_03365_),
    .D(_03368_),
    .X(_03369_));
 sg13g2_a21oi_1 _11921_ (.A1(\m_sys.m_core.m_bru.io_i_s2[16] ),
    .A2(net5089),
    .Y(_03370_),
    .B1(_03237_));
 sg13g2_a21oi_1 _11922_ (.A1(\m_sys.m_core.m_bru.io_i_s2[17] ),
    .A2(net5089),
    .Y(_03371_),
    .B1(_03243_));
 sg13g2_a21o_1 _11923_ (.A2(_03370_),
    .A1(_03245_),
    .B1(_03371_),
    .X(_03372_));
 sg13g2_nor2b_1 _11924_ (.A(_03223_),
    .B_N(_03224_),
    .Y(_03373_));
 sg13g2_and2_1 _11925_ (.A(_03227_),
    .B(_03231_),
    .X(_03374_));
 sg13g2_a221oi_1 _11926_ (.B2(_03226_),
    .C1(_03373_),
    .B1(_03374_),
    .A1(_03366_),
    .Y(_03375_),
    .A2(_03372_));
 sg13g2_nor4_1 _11927_ (.A(_03212_),
    .B(_03218_),
    .C(_03365_),
    .D(_03375_),
    .Y(_03376_));
 sg13g2_a21oi_2 _11928_ (.B1(_03210_),
    .Y(_03377_),
    .A2(net5087),
    .A1(\m_sys.m_core.m_bru.io_i_s2[20] ));
 sg13g2_a22oi_1 _11929_ (.Y(_03378_),
    .B1(_03219_),
    .B2(_03377_),
    .A2(_03216_),
    .A1(_03213_));
 sg13g2_and2_1 _11930_ (.A(_03201_),
    .B(_03202_),
    .X(_03379_));
 sg13g2_a22oi_1 _11931_ (.Y(_03380_),
    .B1(_03200_),
    .B2(_03379_),
    .A2(_03197_),
    .A1(_03195_));
 sg13g2_o21ai_1 _11932_ (.B1(_03380_),
    .Y(_03381_),
    .A1(_03365_),
    .A2(_03378_));
 sg13g2_nor2_1 _11933_ (.A(_03376_),
    .B(_03381_),
    .Y(_03382_));
 sg13g2_o21ai_1 _11934_ (.B1(_03382_),
    .Y(_03383_),
    .A1(_03364_),
    .A2(_03369_));
 sg13g2_nand2_1 _11935_ (.Y(_03384_),
    .A(_03277_),
    .B(_03282_));
 sg13g2_and4_1 _11936_ (.A(_03264_),
    .B(_03270_),
    .C(_03277_),
    .D(_03282_),
    .X(_03385_));
 sg13g2_a21oi_1 _11937_ (.A1(\m_sys.m_core.m_bru.io_i_s2[24] ),
    .A2(net5087),
    .Y(_03386_),
    .B1(_03280_));
 sg13g2_and2_1 _11938_ (.A(_03272_),
    .B(_03274_),
    .X(_03387_));
 sg13g2_a21o_1 _11939_ (.A2(_03386_),
    .A1(_03277_),
    .B1(_03387_),
    .X(_03388_));
 sg13g2_nand3_1 _11940_ (.B(_03270_),
    .C(_03388_),
    .A(_03264_),
    .Y(_03389_));
 sg13g2_nor2_1 _11941_ (.A(_03265_),
    .B(_03268_),
    .Y(_03390_));
 sg13g2_a22oi_1 _11942_ (.Y(_03391_),
    .B1(_03264_),
    .B2(_03390_),
    .A2(_03261_),
    .A1(_03259_));
 sg13g2_nand2_1 _11943_ (.Y(_03392_),
    .A(_03389_),
    .B(_03391_));
 sg13g2_a21oi_2 _11944_ (.B1(_03392_),
    .Y(_03393_),
    .A2(_03385_),
    .A1(_03383_));
 sg13g2_nand2_1 _11945_ (.Y(_03394_),
    .A(_03293_),
    .B(_03298_));
 sg13g2_a21oi_1 _11946_ (.A1(\m_sys.m_core.m_bru.io_i_s2[28] ),
    .A2(net5085),
    .Y(_03395_),
    .B1(_03296_));
 sg13g2_a22oi_1 _11947_ (.Y(_03396_),
    .B1(_03293_),
    .B2(_03395_),
    .A2(_03291_),
    .A1(_03289_));
 sg13g2_o21ai_1 _11948_ (.B1(_03396_),
    .Y(_03397_),
    .A1(_03393_),
    .A2(_03394_));
 sg13g2_nand2b_1 _11949_ (.Y(_03398_),
    .B(_03397_),
    .A_N(_03304_));
 sg13g2_nand2_1 _11950_ (.Y(_03399_),
    .A(_03070_),
    .B(_03071_));
 sg13g2_a21o_1 _11951_ (.A2(_03399_),
    .A1(_03398_),
    .B1(net5169),
    .X(_03400_));
 sg13g2_o21ai_1 _11952_ (.B1(_03400_),
    .Y(_03401_),
    .A1(net5247),
    .A2(_03303_));
 sg13g2_mux2_2 _11953_ (.A0(\m_sys._m_core_io_b_mem_wdata[31] ),
    .A1(net5353),
    .S(net5082),
    .X(_03402_));
 sg13g2_nand2_1 _11954_ (.Y(_03403_),
    .A(\m_sys.m_core.m_bru.io_i_s2[31] ),
    .B(net5083));
 sg13g2_nor2_2 _11955_ (.A(net5353),
    .B(_02475_),
    .Y(_03404_));
 sg13g2_nand2b_1 _11956_ (.Y(_03405_),
    .B(_03403_),
    .A_N(net4884));
 sg13g2_nand3_1 _11957_ (.B(\m_sys.m_core.m_bru.io_i_s2[31] ),
    .C(net5083),
    .A(net5353),
    .Y(_03406_));
 sg13g2_nand2_1 _11958_ (.Y(_03407_),
    .A(_03405_),
    .B(_03406_));
 sg13g2_a21oi_1 _11959_ (.A1(_03405_),
    .A2(_03406_),
    .Y(_03408_),
    .B1(net5303));
 sg13g2_nor2_1 _11960_ (.A(net5162),
    .B(net4893),
    .Y(_03409_));
 sg13g2_nand2_2 _11961_ (.Y(_03410_),
    .A(net5300),
    .B(net4895));
 sg13g2_nand2_1 _11962_ (.Y(_03411_),
    .A(_03082_),
    .B(net4903));
 sg13g2_nand2_1 _11963_ (.Y(_03412_),
    .A(_03075_),
    .B(net4910));
 sg13g2_nand2_1 _11964_ (.Y(_03413_),
    .A(_03411_),
    .B(_03412_));
 sg13g2_nand2_1 _11965_ (.Y(_03414_),
    .A(_03095_),
    .B(net4899));
 sg13g2_nand2_1 _11966_ (.Y(_03415_),
    .A(_03088_),
    .B(net4911));
 sg13g2_nand2_1 _11967_ (.Y(_03416_),
    .A(_03414_),
    .B(_03415_));
 sg13g2_mux2_1 _11968_ (.A0(_03413_),
    .A1(_03416_),
    .S(net4916),
    .X(_03417_));
 sg13g2_mux2_1 _11969_ (.A0(_03338_),
    .A1(_03340_),
    .S(net4899),
    .X(_03418_));
 sg13g2_nand2_1 _11970_ (.Y(_03419_),
    .A(net4898),
    .B(_03172_));
 sg13g2_o21ai_1 _11971_ (.B1(_03419_),
    .Y(_03420_),
    .A1(net4899),
    .A2(_03345_));
 sg13g2_nor2_1 _11972_ (.A(net4934),
    .B(_03420_),
    .Y(_03421_));
 sg13g2_a21oi_1 _11973_ (.A1(net4934),
    .A2(_03418_),
    .Y(_03422_),
    .B1(_03421_));
 sg13g2_nand2_1 _11974_ (.Y(_03423_),
    .A(net4940),
    .B(_03422_));
 sg13g2_o21ai_1 _11975_ (.B1(_03423_),
    .Y(_03424_),
    .A1(net4944),
    .A2(_03417_));
 sg13g2_nand2b_1 _11976_ (.Y(_03425_),
    .B(net4897),
    .A_N(_03129_));
 sg13g2_nor2_1 _11977_ (.A(_03124_),
    .B(net4896),
    .Y(_03426_));
 sg13g2_o21ai_1 _11978_ (.B1(_03425_),
    .Y(_03427_),
    .A1(_03124_),
    .A2(net4896));
 sg13g2_nor2_1 _11979_ (.A(_03133_),
    .B(net4896),
    .Y(_03428_));
 sg13g2_or3_1 _11980_ (.A(net4924),
    .B(_03139_),
    .C(_03428_),
    .X(_03429_));
 sg13g2_o21ai_1 _11981_ (.B1(_03429_),
    .Y(_03430_),
    .A1(net4915),
    .A2(_03427_));
 sg13g2_nor2_1 _11982_ (.A(net4898),
    .B(_03310_),
    .Y(_03431_));
 sg13g2_nor2_1 _11983_ (.A(net4904),
    .B(_03153_),
    .Y(_03432_));
 sg13g2_nor2_1 _11984_ (.A(_03431_),
    .B(_03432_),
    .Y(_03433_));
 sg13g2_nand2_1 _11985_ (.Y(_03434_),
    .A(net4914),
    .B(_03433_));
 sg13g2_nand2_1 _11986_ (.Y(_03435_),
    .A(_03111_),
    .B(net4905));
 sg13g2_o21ai_1 _11987_ (.B1(_03435_),
    .Y(_03436_),
    .A1(net4905),
    .A2(_03306_));
 sg13g2_o21ai_1 _11988_ (.B1(_03434_),
    .Y(_03437_),
    .A1(net4914),
    .A2(_03436_));
 sg13g2_mux2_1 _11989_ (.A0(_03430_),
    .A1(_03437_),
    .S(net4935),
    .X(_03438_));
 sg13g2_nor2_1 _11990_ (.A(net4780),
    .B(_03438_),
    .Y(_03439_));
 sg13g2_a21oi_1 _11991_ (.A1(net4780),
    .A2(_03424_),
    .Y(_03440_),
    .B1(_03439_));
 sg13g2_nand2_1 _11992_ (.Y(_03441_),
    .A(net4770),
    .B(_03440_));
 sg13g2_nor2_1 _11993_ (.A(net5291),
    .B(net5258),
    .Y(_03442_));
 sg13g2_nand2_2 _11994_ (.Y(_03443_),
    .A(net5175),
    .B(net5160));
 sg13g2_nand2_1 _11995_ (.Y(_03444_),
    .A(net4906),
    .B(_03261_));
 sg13g2_o21ai_1 _11996_ (.B1(_03444_),
    .Y(_03445_),
    .A1(net4907),
    .A2(_03268_));
 sg13g2_and2_1 _11997_ (.A(net4906),
    .B(_03274_),
    .X(_03446_));
 sg13g2_a21oi_1 _11998_ (.A1(net4901),
    .A2(_03279_),
    .Y(_03447_),
    .B1(_03446_));
 sg13g2_nor2_1 _11999_ (.A(net4919),
    .B(_03445_),
    .Y(_03448_));
 sg13g2_a21oi_1 _12000_ (.A1(net4919),
    .A2(_03447_),
    .Y(_03449_),
    .B1(_03448_));
 sg13g2_nand2_1 _12001_ (.Y(_03450_),
    .A(_03070_),
    .B(net4901));
 sg13g2_and2_1 _12002_ (.A(net4910),
    .B(_03402_),
    .X(_03451_));
 sg13g2_nor2_1 _12003_ (.A(net4918),
    .B(_03451_),
    .Y(_03452_));
 sg13g2_nand2_1 _12004_ (.Y(_03453_),
    .A(net4901),
    .B(_03295_));
 sg13g2_nand2_1 _12005_ (.Y(_03454_),
    .A(net4907),
    .B(_03291_));
 sg13g2_and2_1 _12006_ (.A(_03453_),
    .B(_03454_),
    .X(_03455_));
 sg13g2_a221oi_1 _12007_ (.B2(net4918),
    .C1(net4943),
    .B1(_03455_),
    .A1(_03450_),
    .Y(_03456_),
    .A2(_03452_));
 sg13g2_a21oi_1 _12008_ (.A1(net4944),
    .A2(_03449_),
    .Y(_03457_),
    .B1(_03456_));
 sg13g2_nand2_1 _12009_ (.Y(_03458_),
    .A(net4928),
    .B(_03451_));
 sg13g2_nor2_1 _12010_ (.A(net5163),
    .B(net4895),
    .Y(_03459_));
 sg13g2_nand2_1 _12011_ (.Y(_03460_),
    .A(net5298),
    .B(net4894));
 sg13g2_nand2_1 _12012_ (.Y(_03461_),
    .A(net4902),
    .B(_03230_));
 sg13g2_nand2_1 _12013_ (.Y(_03462_),
    .A(net4908),
    .B(_03223_));
 sg13g2_nand2_1 _12014_ (.Y(_03463_),
    .A(_03461_),
    .B(_03462_));
 sg13g2_nand2_1 _12015_ (.Y(_03464_),
    .A(net4901),
    .B(_03237_));
 sg13g2_nand2_1 _12016_ (.Y(_03465_),
    .A(net4909),
    .B(_03243_));
 sg13g2_nand2_1 _12017_ (.Y(_03466_),
    .A(_03464_),
    .B(_03465_));
 sg13g2_mux2_1 _12018_ (.A0(_03463_),
    .A1(_03466_),
    .S(net4921),
    .X(_03467_));
 sg13g2_nand2_1 _12019_ (.Y(_03468_),
    .A(net4908),
    .B(_03197_));
 sg13g2_nand2_1 _12020_ (.Y(_03469_),
    .A(net4902),
    .B(_03201_));
 sg13g2_nand2_1 _12021_ (.Y(_03470_),
    .A(_03468_),
    .B(_03469_));
 sg13g2_nand2_1 _12022_ (.Y(_03471_),
    .A(net4931),
    .B(_03470_));
 sg13g2_nand2_1 _12023_ (.Y(_03472_),
    .A(net4902),
    .B(_03210_));
 sg13g2_nand2_1 _12024_ (.Y(_03473_),
    .A(net4909),
    .B(_03215_));
 sg13g2_nand2_1 _12025_ (.Y(_03474_),
    .A(_03472_),
    .B(_03473_));
 sg13g2_o21ai_1 _12026_ (.B1(_03471_),
    .Y(_03475_),
    .A1(net4930),
    .A2(_03474_));
 sg13g2_inv_1 _12027_ (.Y(_03476_),
    .A(_03475_));
 sg13g2_nor2_1 _12028_ (.A(net4944),
    .B(_03475_),
    .Y(_03477_));
 sg13g2_a21oi_1 _12029_ (.A1(net4941),
    .A2(_03467_),
    .Y(_03478_),
    .B1(_03477_));
 sg13g2_a21oi_1 _12030_ (.A1(net4954),
    .A2(_03478_),
    .Y(_03479_),
    .B1(net4763));
 sg13g2_o21ai_1 _12031_ (.B1(_03479_),
    .Y(_03480_),
    .A1(net4954),
    .A2(_03457_));
 sg13g2_nand3_1 _12032_ (.B(_03442_),
    .C(_03480_),
    .A(_03441_),
    .Y(_03481_));
 sg13g2_nor2_1 _12033_ (.A(net5303),
    .B(_03407_),
    .Y(_03482_));
 sg13g2_mux2_1 _12034_ (.A0(_03482_),
    .A1(_03408_),
    .S(_03401_),
    .X(_03483_));
 sg13g2_nand3_1 _12035_ (.B(net5303),
    .C(_03402_),
    .A(net5247),
    .Y(_03484_));
 sg13g2_and2_2 _12036_ (.A(net4761),
    .B(_03484_),
    .X(_03485_));
 sg13g2_nand2_1 _12037_ (.Y(_03486_),
    .A(net4761),
    .B(_03484_));
 sg13g2_nor2_1 _12038_ (.A(net5253),
    .B(net4953),
    .Y(_03487_));
 sg13g2_inv_1 _12039_ (.Y(_03488_),
    .A(_03487_));
 sg13g2_nand4_1 _12040_ (.B(net4929),
    .C(_03451_),
    .A(net4937),
    .Y(_03489_),
    .D(_03487_));
 sg13g2_o21ai_1 _12041_ (.B1(_03484_),
    .Y(_03490_),
    .A1(net4761),
    .A2(_03489_));
 sg13g2_or3_1 _12042_ (.A(net5289),
    .B(_03482_),
    .C(_03490_),
    .X(_03491_));
 sg13g2_nand2_1 _12043_ (.Y(_03492_),
    .A(net5163),
    .B(_03405_));
 sg13g2_nand3_1 _12044_ (.B(_03406_),
    .C(_03492_),
    .A(net5289),
    .Y(_03493_));
 sg13g2_nand3_1 _12045_ (.B(_03491_),
    .C(_03493_),
    .A(net5257),
    .Y(_03494_));
 sg13g2_o21ai_1 _12046_ (.B1(_03494_),
    .Y(_03495_),
    .A1(_03481_),
    .A2(_03483_));
 sg13g2_nor2_1 _12047_ (.A(net4975),
    .B(net5096),
    .Y(_03496_));
 sg13g2_nand2_1 _12048_ (.Y(_03497_),
    .A(net4958),
    .B(net5093));
 sg13g2_and3_2 _12049_ (.X(_03498_),
    .A(_02676_),
    .B(_02693_),
    .C(_02696_));
 sg13g2_mux2_1 _12050_ (.A0(_00136_),
    .A1(_00135_),
    .S(_03498_),
    .X(_03499_));
 sg13g2_nor4_2 _12051_ (.A(\m_sys.r_addr[8] ),
    .B(\m_sys.r_addr[9] ),
    .C(\m_sys.r_addr[10] ),
    .Y(_03500_),
    .D(\m_sys.r_addr[7] ));
 sg13g2_nand4_1 _12052_ (.B(_02413_),
    .C(_02415_),
    .A(_02412_),
    .Y(_03501_),
    .D(_02416_));
 sg13g2_mux2_1 _12053_ (.A0(\m_sys._m_ram_io_b_port_rdata[23] ),
    .A1(\m_sys._m_ram_io_b_port_rdata[31] ),
    .S(net5363),
    .X(_03502_));
 sg13g2_nand2_1 _12054_ (.Y(_03503_),
    .A(net5360),
    .B(_00063_));
 sg13g2_o21ai_1 _12055_ (.B1(_03503_),
    .Y(_03504_),
    .A1(net5360),
    .A2(_02419_));
 sg13g2_nor2_1 _12056_ (.A(net5354),
    .B(_03504_),
    .Y(_03505_));
 sg13g2_nor2_1 _12057_ (.A(\m_sys.r_addr[11] ),
    .B(_03501_),
    .Y(_03506_));
 sg13g2_nand2_1 _12058_ (.Y(_03507_),
    .A(_02414_),
    .B(_03500_));
 sg13g2_a21o_1 _12059_ (.A2(_03502_),
    .A1(net5354),
    .B1(net5072),
    .X(_03508_));
 sg13g2_o21ai_1 _12060_ (.B1(net5277),
    .Y(_03509_),
    .A1(_03505_),
    .A2(_03508_));
 sg13g2_nand2_1 _12061_ (.Y(_03510_),
    .A(\m_sys.r_addr[11] ),
    .B(_03500_));
 sg13g2_nor2_2 _12062_ (.A(\m_sys.r_addr[6] ),
    .B(_03510_),
    .Y(_03511_));
 sg13g2_or2_2 _12063_ (.X(_03512_),
    .B(_03510_),
    .A(\m_sys.r_addr[6] ));
 sg13g2_nand2_2 _12064_ (.Y(_03513_),
    .A(\m_sys.r_addr[11] ),
    .B(\m_sys.r_addr[6] ));
 sg13g2_nor2_2 _12065_ (.A(_03501_),
    .B(_03513_),
    .Y(_03514_));
 sg13g2_or2_1 _12066_ (.X(_03515_),
    .B(_03513_),
    .A(_03501_));
 sg13g2_a221oi_1 _12067_ (.B2(_00136_),
    .C1(_03509_),
    .B1(net4882),
    .A1(_00135_),
    .Y(_03516_),
    .A2(_03511_));
 sg13g2_a22oi_1 _12068_ (.Y(_03517_),
    .B1(_03500_),
    .B2(_03516_),
    .A2(net4493),
    .A1(_02419_));
 sg13g2_o21ai_1 _12069_ (.B1(_03517_),
    .Y(_03518_),
    .A1(net4493),
    .A2(_03499_));
 sg13g2_o21ai_1 _12070_ (.B1(_03518_),
    .Y(_03519_),
    .A1(_02411_),
    .A2(_03516_));
 sg13g2_nor2_1 _12071_ (.A(_02501_),
    .B(_03519_),
    .Y(_03520_));
 sg13g2_nor2_1 _12072_ (.A(\m_sys.m_core.r_ctrl_mem_size[0] ),
    .B(_03520_),
    .Y(_03521_));
 sg13g2_nor2_1 _12073_ (.A(\m_sys.m_core.r_ctrl_mem_size[1] ),
    .B(_03521_),
    .Y(_03522_));
 sg13g2_nor2_2 _12074_ (.A(net4493),
    .B(_03498_),
    .Y(_03523_));
 sg13g2_nand2b_1 _12075_ (.Y(_03524_),
    .B(_03523_),
    .A_N(_00143_));
 sg13g2_nor2_1 _12076_ (.A(net5364),
    .B(_02420_),
    .Y(_03525_));
 sg13g2_a21oi_1 _12077_ (.A1(net5363),
    .A2(_00144_),
    .Y(_03526_),
    .B1(_03525_));
 sg13g2_nand2b_1 _12078_ (.Y(_03527_),
    .B(\m_sys._m_ram_io_b_port_rdata[31] ),
    .A_N(net5363));
 sg13g2_o21ai_1 _12079_ (.B1(_03506_),
    .Y(_03528_),
    .A1(net5358),
    .A2(_03526_));
 sg13g2_a21oi_1 _12080_ (.A1(net5358),
    .A2(_03527_),
    .Y(_03529_),
    .B1(_03528_));
 sg13g2_or2_1 _12081_ (.X(_03530_),
    .B(_03529_),
    .A(_03514_));
 sg13g2_a22oi_1 _12082_ (.Y(_03531_),
    .B1(_03530_),
    .B2(net5278),
    .A2(net4497),
    .A1(_02420_));
 sg13g2_nor2_1 _12083_ (.A(_02411_),
    .B(_03501_),
    .Y(_03532_));
 sg13g2_nand2_1 _12084_ (.Y(_03533_),
    .A(net5274),
    .B(_03500_));
 sg13g2_o21ai_1 _12085_ (.B1(net4879),
    .Y(_03534_),
    .A1(_00143_),
    .A2(_03513_));
 sg13g2_nor2_1 _12086_ (.A(_03529_),
    .B(_03534_),
    .Y(_03535_));
 sg13g2_a21oi_1 _12087_ (.A1(_03524_),
    .A2(_03531_),
    .Y(_03536_),
    .B1(_03535_));
 sg13g2_nand2_1 _12088_ (.Y(_03537_),
    .A(\m_sys.m_core.r_ctrl_mem_signed ),
    .B(_03536_));
 sg13g2_or2_2 _12089_ (.X(_03538_),
    .B(_02754_),
    .A(\m_sys.m_core.r_ctrl_mem_rw ));
 sg13g2_a21oi_1 _12090_ (.A1(\m_sys.m_core.r_ctrl_mem_size[0] ),
    .A2(_03537_),
    .Y(_03539_),
    .B1(_03538_));
 sg13g2_a21oi_1 _12091_ (.A1(_03522_),
    .A2(_03539_),
    .Y(_03540_),
    .B1(net5101));
 sg13g2_nor2_1 _12092_ (.A(_02720_),
    .B(_03538_),
    .Y(_03541_));
 sg13g2_nor3_2 _12093_ (.A(_02411_),
    .B(net5356),
    .C(net5073),
    .Y(_03542_));
 sg13g2_nand2b_1 _12094_ (.Y(_03543_),
    .B(_03542_),
    .A_N(_03527_));
 sg13g2_nand3_1 _12095_ (.B(net4496),
    .C(net5070),
    .A(\m_sys._m_ram_io_b_port_rdata[31] ),
    .Y(_03544_));
 sg13g2_a21o_1 _12096_ (.A2(_03544_),
    .A1(_03543_),
    .B1(net4745),
    .X(_03545_));
 sg13g2_a21oi_2 _12097_ (.B1(net4748),
    .Y(_03546_),
    .A2(_03545_),
    .A1(net4040));
 sg13g2_o21ai_1 _12098_ (.B1(_03546_),
    .Y(_03547_),
    .A1(net5098),
    .A2(_03495_));
 sg13g2_nand2_2 _12099_ (.Y(_03548_),
    .A(\m_sys.m_core.r_ctrl_mem_size[1] ),
    .B(\m_sys.m_core.r_ctrl_mem_size[0] ));
 sg13g2_nand3b_1 _12100_ (.B(net5097),
    .C(_03538_),
    .Y(_03549_),
    .A_N(_02755_));
 sg13g2_o21ai_1 _12101_ (.B1(_03549_),
    .Y(_03550_),
    .A1(_03538_),
    .A2(_03548_));
 sg13g2_nor3_1 _12102_ (.A(net5231),
    .B(net5313),
    .C(_02770_),
    .Y(_03551_));
 sg13g2_nand3_1 _12103_ (.B(net5226),
    .C(_03551_),
    .A(net5316),
    .Y(_03552_));
 sg13g2_nand2b_1 _12104_ (.Y(_03553_),
    .B(_03552_),
    .A_N(net5102));
 sg13g2_nor2_1 _12105_ (.A(\m_sys.m_core._m_decoder_io_o_rs1[0] ),
    .B(net5325),
    .Y(_03554_));
 sg13g2_nor2_2 _12106_ (.A(_02772_),
    .B(_02782_),
    .Y(_03555_));
 sg13g2_and2_2 _12107_ (.A(_02779_),
    .B(_03551_),
    .X(_03556_));
 sg13g2_nor2_2 _12108_ (.A(net4744),
    .B(_03556_),
    .Y(_03557_));
 sg13g2_a221oi_1 _12109_ (.B2(_03557_),
    .C1(net4743),
    .B1(_03555_),
    .A1(net5179),
    .Y(_03558_),
    .A2(net5148));
 sg13g2_and2_2 _12110_ (.A(net4975),
    .B(net4492),
    .X(_03559_));
 sg13g2_nand2_2 _12111_ (.Y(_03560_),
    .A(net4976),
    .B(_03558_));
 sg13g2_nor2_1 _12112_ (.A(_02445_),
    .B(net5189),
    .Y(_03561_));
 sg13g2_nand2_1 _12113_ (.Y(_03562_),
    .A(\m_sys.m_core.m_gpr._GEN[127] ),
    .B(net5060));
 sg13g2_nor2_2 _12114_ (.A(net5324),
    .B(net5185),
    .Y(_03563_));
 sg13g2_a221oi_1 _12115_ (.B2(net5051),
    .C1(net5328),
    .B1(\m_sys.m_core.m_gpr._GEN[95] ),
    .A1(net5184),
    .Y(_03564_),
    .A2(\m_sys.m_core.m_gpr._GEN[63] ));
 sg13g2_nor2_1 _12116_ (.A(net5191),
    .B(net5325),
    .Y(_03565_));
 sg13g2_a22oi_1 _12117_ (.Y(_03566_),
    .B1(net5046),
    .B2(\m_sys.m_core.m_gpr._GEN[191] ),
    .A2(net5060),
    .A1(\m_sys.m_core.m_gpr._GEN[255] ));
 sg13g2_a221oi_1 _12118_ (.B2(\m_sys.m_core.m_gpr._GEN[223] ),
    .C1(net5178),
    .B1(net5051),
    .A1(\m_sys.m_core.m_gpr._GEN[159] ),
    .Y(_03567_),
    .A2(net5148));
 sg13g2_a22oi_1 _12119_ (.Y(_03568_),
    .B1(_03566_),
    .B2(_03567_),
    .A2(_03564_),
    .A1(_03562_));
 sg13g2_a21oi_1 _12120_ (.A1(_03559_),
    .A2(_03568_),
    .Y(_03569_),
    .B1(net4724));
 sg13g2_a22oi_1 _12121_ (.Y(_00196_),
    .B1(_03569_),
    .B2(_03547_),
    .A2(net4724),
    .A1(_02444_));
 sg13g2_a221oi_1 _12122_ (.B2(_03292_),
    .C1(net5247),
    .B1(_03300_),
    .A1(_03288_),
    .Y(_03570_),
    .A2(_03299_));
 sg13g2_and2_1 _12123_ (.A(net5247),
    .B(_03397_),
    .X(_03571_));
 sg13g2_o21ai_1 _12124_ (.B1(_03304_),
    .Y(_03572_),
    .A1(_03570_),
    .A2(_03571_));
 sg13g2_or3_1 _12125_ (.A(_03304_),
    .B(_03570_),
    .C(_03571_),
    .X(_03573_));
 sg13g2_nand3_1 _12126_ (.B(_03572_),
    .C(_03573_),
    .A(net5163),
    .Y(_03574_));
 sg13g2_mux2_1 _12127_ (.A0(_03306_),
    .A1(_03310_),
    .S(net4898),
    .X(_03575_));
 sg13g2_nand2_1 _12128_ (.Y(_03576_),
    .A(net4924),
    .B(_03575_));
 sg13g2_nor2_1 _12129_ (.A(_03124_),
    .B(net4904),
    .Y(_03577_));
 sg13g2_nor2_1 _12130_ (.A(net4896),
    .B(_03153_),
    .Y(_03578_));
 sg13g2_or2_1 _12131_ (.X(_03579_),
    .B(_03578_),
    .A(_03577_));
 sg13g2_o21ai_1 _12132_ (.B1(_03576_),
    .Y(_03580_),
    .A1(net4924),
    .A2(_03579_));
 sg13g2_nor2_1 _12133_ (.A(net4945),
    .B(_03580_),
    .Y(_03581_));
 sg13g2_nor2_1 _12134_ (.A(_03133_),
    .B(net4904),
    .Y(_03582_));
 sg13g2_nor2_2 _12135_ (.A(_03129_),
    .B(net4897),
    .Y(_03583_));
 sg13g2_o21ai_1 _12136_ (.B1(net4924),
    .Y(_03584_),
    .A1(_03582_),
    .A2(_03583_));
 sg13g2_or2_2 _12137_ (.X(_03585_),
    .B(_03138_),
    .A(net4899));
 sg13g2_o21ai_1 _12138_ (.B1(_03584_),
    .Y(_03586_),
    .A1(net4925),
    .A2(_03585_));
 sg13g2_a21oi_1 _12139_ (.A1(net4945),
    .A2(_03586_),
    .Y(_03587_),
    .B1(_03581_));
 sg13g2_nand2_1 _12140_ (.Y(_03588_),
    .A(net4949),
    .B(_03587_));
 sg13g2_mux2_1 _12141_ (.A0(_03340_),
    .A1(_03345_),
    .S(net4899),
    .X(_03589_));
 sg13g2_nand2_1 _12142_ (.Y(_03590_),
    .A(_03111_),
    .B(net4896));
 sg13g2_and2_1 _12143_ (.A(net4905),
    .B(_03172_),
    .X(_03591_));
 sg13g2_a21o_1 _12144_ (.A2(net4898),
    .A1(_03111_),
    .B1(_03591_),
    .X(_03592_));
 sg13g2_nand2_1 _12145_ (.Y(_03593_),
    .A(net4915),
    .B(_03592_));
 sg13g2_o21ai_1 _12146_ (.B1(_03593_),
    .Y(_03594_),
    .A1(net4915),
    .A2(_03589_));
 sg13g2_nand2_1 _12147_ (.Y(_03595_),
    .A(net4940),
    .B(_03594_));
 sg13g2_nand2_1 _12148_ (.Y(_03596_),
    .A(_03088_),
    .B(net4899));
 sg13g2_nand2_1 _12149_ (.Y(_03597_),
    .A(_03082_),
    .B(net4910));
 sg13g2_and2_1 _12150_ (.A(_03596_),
    .B(_03597_),
    .X(_03598_));
 sg13g2_nand2_1 _12151_ (.Y(_03599_),
    .A(net4899),
    .B(_03338_));
 sg13g2_nand2_1 _12152_ (.Y(_03600_),
    .A(_03095_),
    .B(net4911));
 sg13g2_nand2_1 _12153_ (.Y(_03601_),
    .A(_03599_),
    .B(_03600_));
 sg13g2_nand2_1 _12154_ (.Y(_03602_),
    .A(net4916),
    .B(_03601_));
 sg13g2_o21ai_1 _12155_ (.B1(_03602_),
    .Y(_03603_),
    .A1(net4916),
    .A2(_03598_));
 sg13g2_o21ai_1 _12156_ (.B1(_03595_),
    .Y(_03604_),
    .A1(net4940),
    .A2(_03603_));
 sg13g2_o21ai_1 _12157_ (.B1(_03588_),
    .Y(_03605_),
    .A1(net4949),
    .A2(_03604_));
 sg13g2_nor2b_1 _12158_ (.A(net5259),
    .B_N(_00088_),
    .Y(_03606_));
 sg13g2_nand2_2 _12159_ (.Y(_03607_),
    .A(net5160),
    .B(_00088_));
 sg13g2_nor2_1 _12160_ (.A(net4906),
    .B(_03274_),
    .Y(_03608_));
 sg13g2_a21oi_1 _12161_ (.A1(net4906),
    .A2(_03268_),
    .Y(_03609_),
    .B1(_03608_));
 sg13g2_inv_1 _12162_ (.Y(_03610_),
    .A(_03609_));
 sg13g2_nand2_1 _12163_ (.Y(_03611_),
    .A(net4932),
    .B(_03609_));
 sg13g2_nor2_1 _12164_ (.A(net4908),
    .B(_03197_),
    .Y(_03612_));
 sg13g2_a21o_1 _12165_ (.A2(_03280_),
    .A1(net4908),
    .B1(_03612_),
    .X(_03613_));
 sg13g2_o21ai_1 _12166_ (.B1(_03611_),
    .Y(_03614_),
    .A1(net4932),
    .A2(_03613_));
 sg13g2_nor2_1 _12167_ (.A(_03070_),
    .B(net4901),
    .Y(_03615_));
 sg13g2_nor2_1 _12168_ (.A(net4907),
    .B(_03291_),
    .Y(_03616_));
 sg13g2_or3_1 _12169_ (.A(net4918),
    .B(_03615_),
    .C(_03616_),
    .X(_03617_));
 sg13g2_nor2_1 _12170_ (.A(net4906),
    .B(_03261_),
    .Y(_03618_));
 sg13g2_a21oi_1 _12171_ (.A1(net4907),
    .A2(_03296_),
    .Y(_03619_),
    .B1(_03618_));
 sg13g2_a21oi_1 _12172_ (.A1(net4919),
    .A2(_03619_),
    .Y(_03620_),
    .B1(net4942));
 sg13g2_a21oi_1 _12173_ (.A1(_03617_),
    .A2(_03620_),
    .Y(_03621_),
    .B1(net4954));
 sg13g2_o21ai_1 _12174_ (.B1(_03621_),
    .Y(_03622_),
    .A1(net4937),
    .A2(_03614_));
 sg13g2_nor2_1 _12175_ (.A(net4902),
    .B(_03201_),
    .Y(_03623_));
 sg13g2_a21oi_1 _12176_ (.A1(net4901),
    .A2(_03215_),
    .Y(_03624_),
    .B1(_03623_));
 sg13g2_nand2_1 _12177_ (.Y(_03625_),
    .A(net4901),
    .B(_03223_));
 sg13g2_nand2_1 _12178_ (.Y(_03626_),
    .A(net4909),
    .B(_03210_));
 sg13g2_nand2_1 _12179_ (.Y(_03627_),
    .A(_03625_),
    .B(_03626_));
 sg13g2_nor2_1 _12180_ (.A(net4931),
    .B(_03627_),
    .Y(_03628_));
 sg13g2_a21oi_1 _12181_ (.A1(net4930),
    .A2(_03624_),
    .Y(_03629_),
    .B1(_03628_));
 sg13g2_or2_1 _12182_ (.X(_03630_),
    .B(_03629_),
    .A(net4941));
 sg13g2_nand2_1 _12183_ (.Y(_03631_),
    .A(net4901),
    .B(_03243_));
 sg13g2_nand2_2 _12184_ (.Y(_03632_),
    .A(net4908),
    .B(_03230_));
 sg13g2_nand2_1 _12185_ (.Y(_03633_),
    .A(_03075_),
    .B(net4903));
 sg13g2_nand2_1 _12186_ (.Y(_03634_),
    .A(net4910),
    .B(_03237_));
 sg13g2_nand2_1 _12187_ (.Y(_03635_),
    .A(_03633_),
    .B(_03634_));
 sg13g2_a21oi_1 _12188_ (.A1(_03631_),
    .A2(_03632_),
    .Y(_03636_),
    .B1(net4921));
 sg13g2_a21o_1 _12189_ (.A2(_03635_),
    .A1(net4921),
    .B1(_03636_),
    .X(_03637_));
 sg13g2_o21ai_1 _12190_ (.B1(_03630_),
    .Y(_03638_),
    .A1(net4939),
    .A2(_03637_));
 sg13g2_a21oi_1 _12191_ (.A1(net4949),
    .A2(_03638_),
    .Y(_03639_),
    .B1(net4762));
 sg13g2_a221oi_1 _12192_ (.B2(_03639_),
    .C1(_03607_),
    .B1(_03622_),
    .A1(net4769),
    .Y(_03640_),
    .A2(_03605_));
 sg13g2_nor2_1 _12193_ (.A(net5167),
    .B(_03485_),
    .Y(_03641_));
 sg13g2_nand2_2 _12194_ (.Y(_03642_),
    .A(net4953),
    .B(net4884));
 sg13g2_nor2_2 _12195_ (.A(net4937),
    .B(net4884),
    .Y(_03643_));
 sg13g2_nor2_1 _12196_ (.A(net4907),
    .B(net4884),
    .Y(_03644_));
 sg13g2_nor2_1 _12197_ (.A(_03615_),
    .B(_03644_),
    .Y(_03645_));
 sg13g2_nand2_2 _12198_ (.Y(_03646_),
    .A(net4928),
    .B(_03645_));
 sg13g2_nand2_1 _12199_ (.Y(_03647_),
    .A(net4918),
    .B(net4884));
 sg13g2_nand3_1 _12200_ (.B(_03646_),
    .C(_03647_),
    .A(net4937),
    .Y(_03648_));
 sg13g2_nand2b_1 _12201_ (.Y(_03649_),
    .B(_03648_),
    .A_N(_03643_));
 sg13g2_o21ai_1 _12202_ (.B1(_03642_),
    .Y(_03650_),
    .A1(net4953),
    .A2(_03649_));
 sg13g2_o21ai_1 _12203_ (.B1(_03641_),
    .Y(_03651_),
    .A1(net4895),
    .A2(_03650_));
 sg13g2_nor3_1 _12204_ (.A(net4943),
    .B(_03488_),
    .C(_03646_),
    .Y(_03652_));
 sg13g2_nand2_1 _12205_ (.Y(_03653_),
    .A(net5174),
    .B(net5307));
 sg13g2_a221oi_1 _12206_ (.B2(_03652_),
    .C1(net5289),
    .B1(net4766),
    .A1(net5163),
    .Y(_03654_),
    .A2(_03304_));
 sg13g2_o21ai_1 _12207_ (.B1(_03302_),
    .Y(_03655_),
    .A1(net5303),
    .A2(_03072_));
 sg13g2_o21ai_1 _12208_ (.B1(net5257),
    .Y(_03656_),
    .A1(net5174),
    .A2(_03655_));
 sg13g2_a21oi_1 _12209_ (.A1(_03651_),
    .A2(_03654_),
    .Y(_03657_),
    .B1(_03656_));
 sg13g2_a21oi_2 _12210_ (.B1(_03657_),
    .Y(_03658_),
    .A2(_03640_),
    .A1(_03574_));
 sg13g2_nand2_1 _12211_ (.Y(_03659_),
    .A(net5099),
    .B(_03658_));
 sg13g2_nor2b_1 _12212_ (.A(net5361),
    .B_N(\m_sys._m_ram_io_b_port_rdata[30] ),
    .Y(_03660_));
 sg13g2_and2_1 _12213_ (.A(\m_sys._m_ram_io_b_port_rdata[30] ),
    .B(net5069),
    .X(_03661_));
 sg13g2_a22oi_1 _12214_ (.Y(_03662_),
    .B1(_03661_),
    .B2(net4493),
    .A2(_03660_),
    .A1(_03542_));
 sg13g2_o21ai_1 _12215_ (.B1(net4040),
    .Y(_03663_),
    .A1(net4747),
    .A2(_03662_));
 sg13g2_nand3_1 _12216_ (.B(_03659_),
    .C(_03663_),
    .A(net4757),
    .Y(_03664_));
 sg13g2_nand2_1 _12217_ (.Y(_03665_),
    .A(\m_sys.m_core.m_gpr._GEN[126] ),
    .B(net5060));
 sg13g2_a221oi_1 _12218_ (.B2(net5051),
    .C1(net5328),
    .B1(\m_sys.m_core.m_gpr._GEN[94] ),
    .A1(net5184),
    .Y(_03666_),
    .A2(\m_sys.m_core.m_gpr._GEN[62] ));
 sg13g2_a22oi_1 _12219_ (.Y(_03667_),
    .B1(net5046),
    .B2(\m_sys.m_core.m_gpr._GEN[190] ),
    .A2(net5060),
    .A1(\m_sys.m_core.m_gpr._GEN[254] ));
 sg13g2_a221oi_1 _12220_ (.B2(\m_sys.m_core.m_gpr._GEN[222] ),
    .C1(net5178),
    .B1(net5051),
    .A1(\m_sys.m_core.m_gpr._GEN[158] ),
    .Y(_03668_),
    .A2(net5148));
 sg13g2_a22oi_1 _12221_ (.Y(_03669_),
    .B1(_03667_),
    .B2(_03668_),
    .A2(_03666_),
    .A1(_03665_));
 sg13g2_a21oi_2 _12222_ (.B1(net4724),
    .Y(_03670_),
    .A2(_03669_),
    .A1(_03559_));
 sg13g2_a22oi_1 _12223_ (.Y(_00197_),
    .B1(_03664_),
    .B2(_03670_),
    .A2(net4723),
    .A1(_02443_));
 sg13g2_nor2_1 _12224_ (.A(net5167),
    .B(_03393_),
    .Y(_03671_));
 sg13g2_a22oi_1 _12225_ (.Y(_03672_),
    .B1(_03671_),
    .B2(_03298_),
    .A2(_03395_),
    .A1(net5247));
 sg13g2_nand2_1 _12226_ (.Y(_03673_),
    .A(net5167),
    .B(_03294_));
 sg13g2_a21o_1 _12227_ (.A2(_03297_),
    .A1(_03288_),
    .B1(_03673_),
    .X(_03674_));
 sg13g2_a21o_1 _12228_ (.A2(_03674_),
    .A1(_03672_),
    .B1(_03293_),
    .X(_03675_));
 sg13g2_nand3_1 _12229_ (.B(_03672_),
    .C(_03674_),
    .A(_03293_),
    .Y(_03676_));
 sg13g2_nand3_1 _12230_ (.B(_03675_),
    .C(_03676_),
    .A(net5163),
    .Y(_03677_));
 sg13g2_nor2_1 _12231_ (.A(net4914),
    .B(_03433_),
    .Y(_03678_));
 sg13g2_a21oi_1 _12232_ (.A1(net4914),
    .A2(_03427_),
    .Y(_03679_),
    .B1(_03678_));
 sg13g2_nand2b_1 _12233_ (.Y(_03680_),
    .B(net4935),
    .A_N(_03679_));
 sg13g2_o21ai_1 _12234_ (.B1(net4924),
    .Y(_03681_),
    .A1(_03139_),
    .A2(_03428_));
 sg13g2_o21ai_1 _12235_ (.B1(_03680_),
    .Y(_03682_),
    .A1(net4935),
    .A2(_03681_));
 sg13g2_mux2_1 _12236_ (.A0(_03420_),
    .A1(_03436_),
    .S(net4914),
    .X(_03683_));
 sg13g2_mux2_1 _12237_ (.A0(_03416_),
    .A1(_03418_),
    .S(net4916),
    .X(_03684_));
 sg13g2_nor2_1 _12238_ (.A(net4940),
    .B(_03684_),
    .Y(_03685_));
 sg13g2_a21oi_1 _12239_ (.A1(net4940),
    .A2(_03683_),
    .Y(_03686_),
    .B1(_03685_));
 sg13g2_nand2_1 _12240_ (.Y(_03687_),
    .A(net4778),
    .B(_03686_));
 sg13g2_o21ai_1 _12241_ (.B1(_03687_),
    .Y(_03688_),
    .A1(net4778),
    .A2(_03682_));
 sg13g2_nor2_1 _12242_ (.A(net4920),
    .B(_03447_),
    .Y(_03689_));
 sg13g2_a21oi_2 _12243_ (.B1(_03689_),
    .Y(_03690_),
    .A2(_03470_),
    .A1(net4920));
 sg13g2_a21oi_1 _12244_ (.A1(net4928),
    .A2(_03455_),
    .Y(_03691_),
    .B1(net4942));
 sg13g2_o21ai_1 _12245_ (.B1(_03691_),
    .Y(_03692_),
    .A1(net4928),
    .A2(_03445_));
 sg13g2_o21ai_1 _12246_ (.B1(_03692_),
    .Y(_03693_),
    .A1(net4937),
    .A2(_03690_));
 sg13g2_mux2_1 _12247_ (.A0(_03463_),
    .A1(_03474_),
    .S(net4930),
    .X(_03694_));
 sg13g2_mux2_1 _12248_ (.A0(_03413_),
    .A1(_03466_),
    .S(net4933),
    .X(_03695_));
 sg13g2_mux2_1 _12249_ (.A0(_03694_),
    .A1(_03695_),
    .S(net4941),
    .X(_03696_));
 sg13g2_nand2b_1 _12250_ (.Y(_03697_),
    .B(net4951),
    .A_N(_03696_));
 sg13g2_a21oi_1 _12251_ (.A1(net4783),
    .A2(_03693_),
    .Y(_03698_),
    .B1(net4763));
 sg13g2_a221oi_1 _12252_ (.B2(_03698_),
    .C1(_03443_),
    .B1(_03697_),
    .A1(net4770),
    .Y(_03699_),
    .A2(_03688_));
 sg13g2_a21oi_1 _12253_ (.A1(_03450_),
    .A2(_03454_),
    .Y(_03700_),
    .B1(net4918));
 sg13g2_a21oi_1 _12254_ (.A1(net4918),
    .A2(net4884),
    .Y(_03701_),
    .B1(_03700_));
 sg13g2_a21oi_1 _12255_ (.A1(net4937),
    .A2(_03701_),
    .Y(_03702_),
    .B1(_03643_));
 sg13g2_nand2_1 _12256_ (.Y(_03703_),
    .A(net4783),
    .B(_03702_));
 sg13g2_nand2_1 _12257_ (.Y(_03704_),
    .A(_03642_),
    .B(_03703_));
 sg13g2_o21ai_1 _12258_ (.B1(_03641_),
    .Y(_03705_),
    .A1(net4895),
    .A2(_03704_));
 sg13g2_a21oi_1 _12259_ (.A1(net4918),
    .A2(_03451_),
    .Y(_03706_),
    .B1(_03700_));
 sg13g2_or2_1 _12260_ (.X(_03707_),
    .B(_03706_),
    .A(net4889));
 sg13g2_or2_1 _12261_ (.X(_03708_),
    .B(_03707_),
    .A(_03488_));
 sg13g2_nor2_1 _12262_ (.A(net4761),
    .B(_03708_),
    .Y(_03709_));
 sg13g2_o21ai_1 _12263_ (.B1(net5174),
    .Y(_03710_),
    .A1(net5303),
    .A2(_03293_));
 sg13g2_nor2_1 _12264_ (.A(_03709_),
    .B(_03710_),
    .Y(_03711_));
 sg13g2_nand2_1 _12265_ (.Y(_03712_),
    .A(net5163),
    .B(_03292_));
 sg13g2_nand3_1 _12266_ (.B(_03290_),
    .C(_03712_),
    .A(net5289),
    .Y(_03713_));
 sg13g2_a21oi_1 _12267_ (.A1(_03705_),
    .A2(_03711_),
    .Y(_03714_),
    .B1(net5160));
 sg13g2_a22oi_1 _12268_ (.Y(_03715_),
    .B1(_03713_),
    .B2(_03714_),
    .A2(_03699_),
    .A1(_03677_));
 sg13g2_nand2b_1 _12269_ (.Y(_03716_),
    .B(\m_sys._m_ram_io_b_port_rdata[29] ),
    .A_N(net5362));
 sg13g2_nand3b_1 _12270_ (.B(_03542_),
    .C(\m_sys._m_ram_io_b_port_rdata[29] ),
    .Y(_03717_),
    .A_N(net5365));
 sg13g2_nand3_1 _12271_ (.B(net4495),
    .C(net5070),
    .A(\m_sys._m_ram_io_b_port_rdata[29] ),
    .Y(_03718_));
 sg13g2_a21o_2 _12272_ (.A2(_03718_),
    .A1(_03717_),
    .B1(net4745),
    .X(_03719_));
 sg13g2_a221oi_1 _12273_ (.B2(net4039),
    .C1(net4753),
    .B1(_03719_),
    .A1(net5099),
    .Y(_03720_),
    .A2(_03715_));
 sg13g2_nand2_1 _12274_ (.Y(_03721_),
    .A(\m_sys.m_core.m_gpr._GEN[125] ),
    .B(net5065));
 sg13g2_a221oi_1 _12275_ (.B2(net5055),
    .C1(net5329),
    .B1(\m_sys.m_core.m_gpr._GEN[93] ),
    .A1(net5186),
    .Y(_03722_),
    .A2(\m_sys.m_core.m_gpr._GEN[61] ));
 sg13g2_a22oi_1 _12276_ (.Y(_03723_),
    .B1(net5048),
    .B2(\m_sys.m_core.m_gpr._GEN[189] ),
    .A2(net5065),
    .A1(\m_sys.m_core.m_gpr._GEN[253] ));
 sg13g2_a221oi_1 _12277_ (.B2(\m_sys.m_core.m_gpr._GEN[221] ),
    .C1(net5181),
    .B1(net5055),
    .A1(\m_sys.m_core.m_gpr._GEN[157] ),
    .Y(_03724_),
    .A2(net5151));
 sg13g2_a221oi_1 _12278_ (.B2(_03724_),
    .C1(_03560_),
    .B1(_03723_),
    .A1(_03721_),
    .Y(_03725_),
    .A2(_03722_));
 sg13g2_nor3_1 _12279_ (.A(net4723),
    .B(_03720_),
    .C(_03725_),
    .Y(_03726_));
 sg13g2_a21oi_1 _12280_ (.A1(net5192),
    .A2(net4723),
    .Y(_00198_),
    .B1(_03726_));
 sg13g2_mux2_1 _12281_ (.A0(_03288_),
    .A1(_03393_),
    .S(net5247),
    .X(_03727_));
 sg13g2_a21oi_1 _12282_ (.A1(_03298_),
    .A2(_03727_),
    .Y(_03728_),
    .B1(net5303));
 sg13g2_o21ai_1 _12283_ (.B1(_03728_),
    .Y(_03729_),
    .A1(_03298_),
    .A2(_03727_));
 sg13g2_nor2_1 _12284_ (.A(net4914),
    .B(_03592_),
    .Y(_03730_));
 sg13g2_a21oi_2 _12285_ (.B1(_03730_),
    .Y(_03731_),
    .A2(_03575_),
    .A1(net4914));
 sg13g2_mux2_1 _12286_ (.A0(_03589_),
    .A1(_03601_),
    .S(net4926),
    .X(_03732_));
 sg13g2_nand2_1 _12287_ (.Y(_03733_),
    .A(net4938),
    .B(_03732_));
 sg13g2_o21ai_1 _12288_ (.B1(_03733_),
    .Y(_03734_),
    .A1(net4938),
    .A2(_03731_));
 sg13g2_nor2_1 _12289_ (.A(net4947),
    .B(_03734_),
    .Y(_03735_));
 sg13g2_or3_1 _12290_ (.A(net4935),
    .B(net4915),
    .C(_03585_),
    .X(_03736_));
 sg13g2_nor3_1 _12291_ (.A(net4927),
    .B(_03582_),
    .C(_03583_),
    .Y(_03737_));
 sg13g2_nor2_1 _12292_ (.A(net4915),
    .B(_03579_),
    .Y(_03738_));
 sg13g2_or2_1 _12293_ (.X(_03739_),
    .B(_03738_),
    .A(_03737_));
 sg13g2_o21ai_1 _12294_ (.B1(_03736_),
    .Y(_03740_),
    .A1(net4945),
    .A2(_03739_));
 sg13g2_a21oi_2 _12295_ (.B1(_03735_),
    .Y(_03741_),
    .A2(_03740_),
    .A1(net4947));
 sg13g2_a21oi_1 _12296_ (.A1(net4920),
    .A2(_03610_),
    .Y(_03742_),
    .B1(net4942));
 sg13g2_o21ai_1 _12297_ (.B1(_03742_),
    .Y(_03743_),
    .A1(net4919),
    .A2(_03619_));
 sg13g2_nand2_1 _12298_ (.Y(_03744_),
    .A(net4920),
    .B(_03624_));
 sg13g2_o21ai_1 _12299_ (.B1(_03744_),
    .Y(_03745_),
    .A1(net4920),
    .A2(_03613_));
 sg13g2_nand2_1 _12300_ (.Y(_03746_),
    .A(net4942),
    .B(_03745_));
 sg13g2_a21oi_2 _12301_ (.B1(net4954),
    .Y(_03747_),
    .A2(_03746_),
    .A1(_03743_));
 sg13g2_nor2_1 _12302_ (.A(net4917),
    .B(_03635_),
    .Y(_03748_));
 sg13g2_a21oi_1 _12303_ (.A1(net4917),
    .A2(_03598_),
    .Y(_03749_),
    .B1(_03748_));
 sg13g2_a21oi_1 _12304_ (.A1(_03631_),
    .A2(_03632_),
    .Y(_03750_),
    .B1(net4930));
 sg13g2_a21o_1 _12305_ (.A2(_03627_),
    .A1(net4930),
    .B1(_03750_),
    .X(_03751_));
 sg13g2_mux2_1 _12306_ (.A0(_03749_),
    .A1(_03751_),
    .S(net4939),
    .X(_03752_));
 sg13g2_o21ai_1 _12307_ (.B1(net4765),
    .Y(_03753_),
    .A1(net4779),
    .A2(_03752_));
 sg13g2_o21ai_1 _12308_ (.B1(_03442_),
    .Y(_03754_),
    .A1(_03747_),
    .A2(_03753_));
 sg13g2_a21oi_1 _12309_ (.A1(net4770),
    .A2(_03741_),
    .Y(_03755_),
    .B1(_03754_));
 sg13g2_a21oi_1 _12310_ (.A1(net4907),
    .A2(_03296_),
    .Y(_03756_),
    .B1(_03616_));
 sg13g2_mux2_1 _12311_ (.A0(_03645_),
    .A1(_03756_),
    .S(net4928),
    .X(_03757_));
 sg13g2_nor2_1 _12312_ (.A(net4943),
    .B(_03757_),
    .Y(_03758_));
 sg13g2_or3_1 _12313_ (.A(net4952),
    .B(_03643_),
    .C(_03758_),
    .X(_03759_));
 sg13g2_nand2_1 _12314_ (.Y(_03760_),
    .A(_03642_),
    .B(_03759_));
 sg13g2_o21ai_1 _12315_ (.B1(_03641_),
    .Y(_03761_),
    .A1(net4895),
    .A2(_03760_));
 sg13g2_nand2_2 _12316_ (.Y(_03762_),
    .A(net4771),
    .B(_03757_));
 sg13g2_nor3_1 _12317_ (.A(net4761),
    .B(_03488_),
    .C(_03762_),
    .Y(_03763_));
 sg13g2_o21ai_1 _12318_ (.B1(net5174),
    .Y(_03764_),
    .A1(net5303),
    .A2(_03298_));
 sg13g2_nor2_1 _12319_ (.A(_03763_),
    .B(_03764_),
    .Y(_03765_));
 sg13g2_nand2_1 _12320_ (.Y(_03766_),
    .A(net5163),
    .B(_03297_));
 sg13g2_nand3_1 _12321_ (.B(_03294_),
    .C(_03766_),
    .A(net5289),
    .Y(_03767_));
 sg13g2_a21oi_1 _12322_ (.A1(_03761_),
    .A2(_03765_),
    .Y(_03768_),
    .B1(net5160));
 sg13g2_a22oi_1 _12323_ (.Y(_03769_),
    .B1(_03767_),
    .B2(_03768_),
    .A2(_03755_),
    .A1(_03729_));
 sg13g2_nand2b_1 _12324_ (.Y(_03770_),
    .B(\m_sys._m_ram_io_b_port_rdata[28] ),
    .A_N(net5362));
 sg13g2_nand3b_1 _12325_ (.B(_03542_),
    .C(\m_sys._m_ram_io_b_port_rdata[28] ),
    .Y(_03771_),
    .A_N(net5365));
 sg13g2_nand3_1 _12326_ (.B(net4495),
    .C(net5070),
    .A(\m_sys._m_ram_io_b_port_rdata[28] ),
    .Y(_03772_));
 sg13g2_a21o_2 _12327_ (.A2(_03772_),
    .A1(_03771_),
    .B1(net4745),
    .X(_03773_));
 sg13g2_a22oi_1 _12328_ (.Y(_03774_),
    .B1(_03773_),
    .B2(net4039),
    .A2(_03769_),
    .A1(net5099));
 sg13g2_nand2_1 _12329_ (.Y(_03775_),
    .A(\m_sys.m_core.m_gpr._GEN[124] ),
    .B(net5059));
 sg13g2_a221oi_1 _12330_ (.B2(net5050),
    .C1(net5328),
    .B1(\m_sys.m_core.m_gpr._GEN[92] ),
    .A1(net5185),
    .Y(_03776_),
    .A2(\m_sys.m_core.m_gpr._GEN[60] ));
 sg13g2_a22oi_1 _12331_ (.Y(_03777_),
    .B1(net5046),
    .B2(\m_sys.m_core.m_gpr._GEN[188] ),
    .A2(net5059),
    .A1(\m_sys.m_core.m_gpr._GEN[252] ));
 sg13g2_a221oi_1 _12332_ (.B2(\m_sys.m_core.m_gpr._GEN[220] ),
    .C1(net5179),
    .B1(net5050),
    .A1(\m_sys.m_core.m_gpr._GEN[156] ),
    .Y(_03778_),
    .A2(net5149));
 sg13g2_a22oi_1 _12333_ (.Y(_03779_),
    .B1(_03777_),
    .B2(_03778_),
    .A2(_03776_),
    .A1(_03775_));
 sg13g2_a221oi_1 _12334_ (.B2(net4385),
    .C1(net4728),
    .B1(_03779_),
    .A1(net4757),
    .Y(_03780_),
    .A2(_03774_));
 sg13g2_a21oi_1 _12335_ (.A1(_02439_),
    .A2(net4728),
    .Y(_00199_),
    .B1(_03780_));
 sg13g2_a21oi_1 _12336_ (.A1(_03258_),
    .A2(_03283_),
    .Y(_03781_),
    .B1(_03285_));
 sg13g2_a21oi_1 _12337_ (.A1(\m_sys.m_core.m_bru.io_i_s1[26] ),
    .A2(_03265_),
    .Y(_03782_),
    .B1(net5248));
 sg13g2_o21ai_1 _12338_ (.B1(_03782_),
    .Y(_03783_),
    .A1(_03269_),
    .A2(_03781_));
 sg13g2_nand2_1 _12339_ (.Y(_03784_),
    .A(net5248),
    .B(_03388_));
 sg13g2_nand2_1 _12340_ (.Y(_03785_),
    .A(net5248),
    .B(_03383_));
 sg13g2_inv_1 _12341_ (.Y(_03786_),
    .A(_03785_));
 sg13g2_o21ai_1 _12342_ (.B1(_03784_),
    .Y(_03787_),
    .A1(_03384_),
    .A2(_03785_));
 sg13g2_a22oi_1 _12343_ (.Y(_03788_),
    .B1(_03787_),
    .B2(_03270_),
    .A2(_03390_),
    .A1(net5248));
 sg13g2_nand2_1 _12344_ (.Y(_03789_),
    .A(_03783_),
    .B(_03788_));
 sg13g2_xnor2_1 _12345_ (.Y(_03790_),
    .A(_03263_),
    .B(_03789_));
 sg13g2_nor2_1 _12346_ (.A(net4938),
    .B(_03437_),
    .Y(_03791_));
 sg13g2_a21oi_1 _12347_ (.A1(net4938),
    .A2(_03422_),
    .Y(_03792_),
    .B1(_03791_));
 sg13g2_nand2_1 _12348_ (.Y(_03793_),
    .A(net4775),
    .B(_03792_));
 sg13g2_nor2_1 _12349_ (.A(net4945),
    .B(_03430_),
    .Y(_03794_));
 sg13g2_o21ai_1 _12350_ (.B1(_03793_),
    .Y(_03795_),
    .A1(net4775),
    .A2(_03794_));
 sg13g2_a21oi_1 _12351_ (.A1(net4942),
    .A2(_03476_),
    .Y(_03796_),
    .B1(net4954));
 sg13g2_o21ai_1 _12352_ (.B1(_03796_),
    .Y(_03797_),
    .A1(net4942),
    .A2(_03449_));
 sg13g2_nand2b_1 _12353_ (.Y(_03798_),
    .B(net4940),
    .A_N(_03417_));
 sg13g2_o21ai_1 _12354_ (.B1(_03798_),
    .Y(_03799_),
    .A1(net4941),
    .A2(_03467_));
 sg13g2_a21oi_1 _12355_ (.A1(net4950),
    .A2(_03799_),
    .Y(_03800_),
    .B1(net4763));
 sg13g2_a221oi_1 _12356_ (.B2(_03800_),
    .C1(_03607_),
    .B1(_03797_),
    .A1(net4769),
    .Y(_03801_),
    .A2(_03795_));
 sg13g2_o21ai_1 _12357_ (.B1(_03801_),
    .Y(_03802_),
    .A1(net5304),
    .A2(_03790_));
 sg13g2_nand2_2 _12358_ (.Y(_03803_),
    .A(net5247),
    .B(_03642_));
 sg13g2_and2_1 _12359_ (.A(_03444_),
    .B(_03453_),
    .X(_03804_));
 sg13g2_a21o_1 _12360_ (.A2(_03454_),
    .A1(_03450_),
    .B1(net4928),
    .X(_03805_));
 sg13g2_o21ai_1 _12361_ (.B1(_03805_),
    .Y(_03806_),
    .A1(net4918),
    .A2(_03804_));
 sg13g2_nor2_1 _12362_ (.A(net4943),
    .B(_03806_),
    .Y(_03807_));
 sg13g2_nor2_1 _12363_ (.A(_03643_),
    .B(_03807_),
    .Y(_03808_));
 sg13g2_a21oi_1 _12364_ (.A1(net4781),
    .A2(_03808_),
    .Y(_03809_),
    .B1(_03803_));
 sg13g2_nand2_1 _12365_ (.Y(_03810_),
    .A(net4771),
    .B(_03806_));
 sg13g2_o21ai_1 _12366_ (.B1(_03810_),
    .Y(_03811_),
    .A1(net4771),
    .A2(_03458_));
 sg13g2_a21oi_1 _12367_ (.A1(net4781),
    .A2(_03811_),
    .Y(_03812_),
    .B1(net5250));
 sg13g2_a21oi_1 _12368_ (.A1(net4892),
    .A2(_03809_),
    .Y(_03813_),
    .B1(_03812_));
 sg13g2_a221oi_1 _12369_ (.B2(_03813_),
    .C1(net5289),
    .B1(_03486_),
    .A1(net5164),
    .Y(_03814_),
    .A2(_03263_));
 sg13g2_nand2_1 _12370_ (.Y(_03815_),
    .A(net5164),
    .B(_03262_));
 sg13g2_nand3_1 _12371_ (.B(_03260_),
    .C(_03815_),
    .A(net5290),
    .Y(_03816_));
 sg13g2_nand2_1 _12372_ (.Y(_03817_),
    .A(net5257),
    .B(_03816_));
 sg13g2_o21ai_1 _12373_ (.B1(_03802_),
    .Y(_03818_),
    .A1(_03814_),
    .A2(_03817_));
 sg13g2_and3_1 _12374_ (.X(_03819_),
    .A(net5278),
    .B(_00047_),
    .C(net4883));
 sg13g2_nand3_1 _12375_ (.B(_00047_),
    .C(net4883),
    .A(net5278),
    .Y(_03820_));
 sg13g2_nand2b_1 _12376_ (.Y(_03821_),
    .B(\m_sys._m_ram_io_b_port_rdata[27] ),
    .A_N(net5364));
 sg13g2_nand3_1 _12377_ (.B(net4495),
    .C(net5071),
    .A(\m_sys._m_ram_io_b_port_rdata[27] ),
    .Y(_03822_));
 sg13g2_o21ai_1 _12378_ (.B1(_03822_),
    .Y(_03823_),
    .A1(_03820_),
    .A2(_03821_));
 sg13g2_nand2b_2 _12379_ (.Y(_03824_),
    .B(_03823_),
    .A_N(net4746));
 sg13g2_a21oi_1 _12380_ (.A1(net4039),
    .A2(_03824_),
    .Y(_03825_),
    .B1(net4751));
 sg13g2_o21ai_1 _12381_ (.B1(_03825_),
    .Y(_03826_),
    .A1(net5098),
    .A2(_03818_));
 sg13g2_nand2_1 _12382_ (.Y(_03827_),
    .A(net3016),
    .B(net5060));
 sg13g2_a221oi_1 _12383_ (.B2(net5051),
    .C1(net5328),
    .B1(\m_sys.m_core.m_gpr._GEN[91] ),
    .A1(net5184),
    .Y(_03828_),
    .A2(\m_sys.m_core.m_gpr._GEN[59] ));
 sg13g2_a22oi_1 _12384_ (.Y(_03829_),
    .B1(net5046),
    .B2(net3449),
    .A2(net5062),
    .A1(\m_sys.m_core.m_gpr._GEN[251] ));
 sg13g2_a221oi_1 _12385_ (.B2(\m_sys.m_core.m_gpr._GEN[219] ),
    .C1(net5178),
    .B1(net5053),
    .A1(\m_sys.m_core.m_gpr._GEN[155] ),
    .Y(_03830_),
    .A2(net5149));
 sg13g2_a22oi_1 _12386_ (.Y(_03831_),
    .B1(_03829_),
    .B2(_03830_),
    .A2(_03828_),
    .A1(_03827_));
 sg13g2_a21oi_1 _12387_ (.A1(_03559_),
    .A2(_03831_),
    .Y(_03832_),
    .B1(net4724));
 sg13g2_a22oi_1 _12388_ (.Y(_00200_),
    .B1(_03826_),
    .B2(_03832_),
    .A2(net4724),
    .A1(net5193));
 sg13g2_a21oi_1 _12389_ (.A1(net5167),
    .A2(_03781_),
    .Y(_03833_),
    .B1(_03787_));
 sg13g2_a21oi_1 _12390_ (.A1(_03270_),
    .A2(_03833_),
    .Y(_03834_),
    .B1(net5304));
 sg13g2_o21ai_1 _12391_ (.B1(_03834_),
    .Y(_03835_),
    .A1(_03270_),
    .A2(_03833_));
 sg13g2_nor2_1 _12392_ (.A(net4935),
    .B(_03580_),
    .Y(_03836_));
 sg13g2_a21oi_1 _12393_ (.A1(net4938),
    .A2(_03594_),
    .Y(_03837_),
    .B1(_03836_));
 sg13g2_a21oi_1 _12394_ (.A1(net4938),
    .A2(_03586_),
    .Y(_03838_),
    .B1(net4776));
 sg13g2_a21o_1 _12395_ (.A2(_03837_),
    .A1(net4776),
    .B1(_03838_),
    .X(_03839_));
 sg13g2_o21ai_1 _12396_ (.B1(net4784),
    .Y(_03840_),
    .A1(net4943),
    .A2(_03614_));
 sg13g2_a21o_1 _12397_ (.A2(_03629_),
    .A1(net4942),
    .B1(_03840_),
    .X(_03841_));
 sg13g2_or2_1 _12398_ (.X(_03842_),
    .B(_03637_),
    .A(net4941));
 sg13g2_o21ai_1 _12399_ (.B1(_03842_),
    .Y(_03843_),
    .A1(net4938),
    .A2(_03603_));
 sg13g2_a21oi_1 _12400_ (.A1(net4950),
    .A2(_03843_),
    .Y(_03844_),
    .B1(net4762));
 sg13g2_a221oi_1 _12401_ (.B2(_03844_),
    .C1(_03443_),
    .B1(_03841_),
    .A1(net4770),
    .Y(_03845_),
    .A2(_03839_));
 sg13g2_a21oi_1 _12402_ (.A1(net4906),
    .A2(_03268_),
    .Y(_03846_),
    .B1(_03618_));
 sg13g2_mux2_1 _12403_ (.A0(_03756_),
    .A1(_03846_),
    .S(net4929),
    .X(_03847_));
 sg13g2_nor2_1 _12404_ (.A(net4888),
    .B(_03847_),
    .Y(_03848_));
 sg13g2_nand3_1 _12405_ (.B(_03646_),
    .C(_03647_),
    .A(net4888),
    .Y(_03849_));
 sg13g2_nor2b_1 _12406_ (.A(_03848_),
    .B_N(_03849_),
    .Y(_03850_));
 sg13g2_a21oi_2 _12407_ (.B1(_03803_),
    .Y(_03851_),
    .A2(_03850_),
    .A1(net4781));
 sg13g2_a21oi_1 _12408_ (.A1(net4888),
    .A2(_03646_),
    .Y(_03852_),
    .B1(_03848_));
 sg13g2_a21o_1 _12409_ (.A2(_03852_),
    .A1(net4781),
    .B1(net5249),
    .X(_03853_));
 sg13g2_a21oi_1 _12410_ (.A1(net4892),
    .A2(_03851_),
    .Y(_03854_),
    .B1(_03485_));
 sg13g2_o21ai_1 _12411_ (.B1(net5173),
    .Y(_03855_),
    .A1(net5305),
    .A2(_03270_));
 sg13g2_a21oi_1 _12412_ (.A1(_03853_),
    .A2(_03854_),
    .Y(_03856_),
    .B1(_03855_));
 sg13g2_a21oi_1 _12413_ (.A1(\m_sys.m_core.m_bru.io_i_s1[26] ),
    .A2(_03265_),
    .Y(_03857_),
    .B1(net5173));
 sg13g2_o21ai_1 _12414_ (.B1(_03857_),
    .Y(_03858_),
    .A1(net5304),
    .A2(_03269_));
 sg13g2_nor2b_1 _12415_ (.A(_03856_),
    .B_N(_03858_),
    .Y(_03859_));
 sg13g2_a22oi_1 _12416_ (.Y(_03860_),
    .B1(_03859_),
    .B2(net5257),
    .A2(_03845_),
    .A1(_03835_));
 sg13g2_nand3b_1 _12417_ (.B(net4740),
    .C(\m_sys._m_ram_io_b_port_rdata[26] ),
    .Y(_03861_),
    .A_N(net5365));
 sg13g2_nand3_1 _12418_ (.B(net4496),
    .C(net5070),
    .A(\m_sys._m_ram_io_b_port_rdata[26] ),
    .Y(_03862_));
 sg13g2_a21o_2 _12419_ (.A2(_03862_),
    .A1(_03861_),
    .B1(net4745),
    .X(_03863_));
 sg13g2_a22oi_1 _12420_ (.Y(_03864_),
    .B1(_03863_),
    .B2(net4038),
    .A2(_03860_),
    .A1(net5100));
 sg13g2_nand2_1 _12421_ (.Y(_03865_),
    .A(\m_sys.m_core.m_gpr._GEN[122] ),
    .B(net5060));
 sg13g2_a221oi_1 _12422_ (.B2(net5051),
    .C1(net5328),
    .B1(\m_sys.m_core.m_gpr._GEN[90] ),
    .A1(net5184),
    .Y(_03866_),
    .A2(\m_sys.m_core.m_gpr._GEN[58] ));
 sg13g2_a22oi_1 _12423_ (.Y(_03867_),
    .B1(net5046),
    .B2(\m_sys.m_core.m_gpr._GEN[186] ),
    .A2(net5060),
    .A1(\m_sys.m_core.m_gpr._GEN[250] ));
 sg13g2_a221oi_1 _12424_ (.B2(\m_sys.m_core.m_gpr._GEN[218] ),
    .C1(net5178),
    .B1(net5051),
    .A1(\m_sys.m_core.m_gpr._GEN[154] ),
    .Y(_03868_),
    .A2(net5148));
 sg13g2_a22oi_1 _12425_ (.Y(_03869_),
    .B1(_03867_),
    .B2(_03868_),
    .A2(_03866_),
    .A1(_03865_));
 sg13g2_a221oi_1 _12426_ (.B2(net4385),
    .C1(net4723),
    .B1(_03869_),
    .A1(net4758),
    .Y(_03870_),
    .A2(_03864_));
 sg13g2_a21oi_1 _12427_ (.A1(net5194),
    .A2(net4723),
    .Y(_00201_),
    .B1(_03870_));
 sg13g2_nand2_1 _12428_ (.Y(_03871_),
    .A(net5167),
    .B(_03278_));
 sg13g2_a21oi_1 _12429_ (.A1(_03258_),
    .A2(_03281_),
    .Y(_03872_),
    .B1(_03871_));
 sg13g2_a221oi_1 _12430_ (.B2(_03282_),
    .C1(_03872_),
    .B1(_03786_),
    .A1(net5248),
    .Y(_03873_),
    .A2(_03386_));
 sg13g2_xnor2_1 _12431_ (.Y(_03874_),
    .A(_03277_),
    .B(_03873_));
 sg13g2_nor2_1 _12432_ (.A(net4945),
    .B(_03681_),
    .Y(_03875_));
 sg13g2_nor2_1 _12433_ (.A(net4935),
    .B(_03679_),
    .Y(_03876_));
 sg13g2_a21oi_1 _12434_ (.A1(net4935),
    .A2(_03683_),
    .Y(_03877_),
    .B1(_03876_));
 sg13g2_nor2_1 _12435_ (.A(net4947),
    .B(_03877_),
    .Y(_03878_));
 sg13g2_a21oi_2 _12436_ (.B1(_03878_),
    .Y(_03879_),
    .A2(_03875_),
    .A1(net4947));
 sg13g2_nand2_1 _12437_ (.Y(_03880_),
    .A(net4941),
    .B(_03694_));
 sg13g2_a21oi_1 _12438_ (.A1(net4937),
    .A2(_03690_),
    .Y(_03881_),
    .B1(net4954));
 sg13g2_nand2_1 _12439_ (.Y(_03882_),
    .A(_03880_),
    .B(_03881_));
 sg13g2_or2_1 _12440_ (.X(_03883_),
    .B(_03684_),
    .A(net4938));
 sg13g2_o21ai_1 _12441_ (.B1(_03883_),
    .Y(_03884_),
    .A1(net4940),
    .A2(_03695_));
 sg13g2_a21oi_1 _12442_ (.A1(net4950),
    .A2(_03884_),
    .Y(_03885_),
    .B1(net4762));
 sg13g2_a221oi_1 _12443_ (.B2(_03885_),
    .C1(_03443_),
    .B1(_03882_),
    .A1(_03409_),
    .Y(_03886_),
    .A2(_03879_));
 sg13g2_o21ai_1 _12444_ (.B1(_03886_),
    .Y(_03887_),
    .A1(net5304),
    .A2(_03874_));
 sg13g2_mux2_1 _12445_ (.A0(_03267_),
    .A1(_03274_),
    .S(net4906),
    .X(_03888_));
 sg13g2_nand2_1 _12446_ (.Y(_03889_),
    .A(net4928),
    .B(_03888_));
 sg13g2_o21ai_1 _12447_ (.B1(_03889_),
    .Y(_03890_),
    .A1(net4929),
    .A2(_03804_));
 sg13g2_nor2_1 _12448_ (.A(net4888),
    .B(_03890_),
    .Y(_03891_));
 sg13g2_a21oi_1 _12449_ (.A1(net4888),
    .A2(_03701_),
    .Y(_03892_),
    .B1(_03891_));
 sg13g2_a21o_1 _12450_ (.A2(_03892_),
    .A1(net4781),
    .B1(_03803_),
    .X(_03893_));
 sg13g2_a21oi_1 _12451_ (.A1(net4888),
    .A2(_03706_),
    .Y(_03894_),
    .B1(_03891_));
 sg13g2_a21oi_1 _12452_ (.A1(net4781),
    .A2(_03894_),
    .Y(_03895_),
    .B1(net5253));
 sg13g2_o21ai_1 _12453_ (.B1(_03486_),
    .Y(_03896_),
    .A1(net4895),
    .A2(_03893_));
 sg13g2_nor2_1 _12454_ (.A(_03895_),
    .B(_03896_),
    .Y(_03897_));
 sg13g2_o21ai_1 _12455_ (.B1(net5173),
    .Y(_03898_),
    .A1(net5304),
    .A2(_03277_));
 sg13g2_nor2_1 _12456_ (.A(_03897_),
    .B(_03898_),
    .Y(_03899_));
 sg13g2_nor2_1 _12457_ (.A(net5304),
    .B(_03275_),
    .Y(_03900_));
 sg13g2_nand2_1 _12458_ (.Y(_03901_),
    .A(net5290),
    .B(_03273_));
 sg13g2_o21ai_1 _12459_ (.B1(net5257),
    .Y(_03902_),
    .A1(_03900_),
    .A2(_03901_));
 sg13g2_o21ai_1 _12460_ (.B1(_03887_),
    .Y(_03903_),
    .A1(_03899_),
    .A2(_03902_));
 sg13g2_nand2b_1 _12461_ (.Y(_03904_),
    .B(\m_sys._m_ram_io_b_port_rdata[25] ),
    .A_N(net5364));
 sg13g2_nand3_1 _12462_ (.B(net4495),
    .C(net5071),
    .A(\m_sys._m_ram_io_b_port_rdata[25] ),
    .Y(_03905_));
 sg13g2_o21ai_1 _12463_ (.B1(_03905_),
    .Y(_03906_),
    .A1(_03820_),
    .A2(_03904_));
 sg13g2_nand2b_2 _12464_ (.Y(_03907_),
    .B(_03906_),
    .A_N(net4745));
 sg13g2_a21oi_1 _12465_ (.A1(net4038),
    .A2(_03907_),
    .Y(_03908_),
    .B1(net4753));
 sg13g2_o21ai_1 _12466_ (.B1(_03908_),
    .Y(_03909_),
    .A1(_03065_),
    .A2(_03903_));
 sg13g2_nand2_1 _12467_ (.Y(_03910_),
    .A(\m_sys.m_core.m_gpr._GEN[121] ),
    .B(net5059));
 sg13g2_a221oi_1 _12468_ (.B2(net5055),
    .C1(net5329),
    .B1(\m_sys.m_core.m_gpr._GEN[89] ),
    .A1(net5186),
    .Y(_03911_),
    .A2(\m_sys.m_core.m_gpr._GEN[57] ));
 sg13g2_a22oi_1 _12469_ (.Y(_03912_),
    .B1(net5046),
    .B2(\m_sys.m_core.m_gpr._GEN[185] ),
    .A2(net5059),
    .A1(\m_sys.m_core.m_gpr._GEN[249] ));
 sg13g2_a221oi_1 _12470_ (.B2(\m_sys.m_core.m_gpr._GEN[217] ),
    .C1(net5178),
    .B1(net5050),
    .A1(\m_sys.m_core.m_gpr._GEN[153] ),
    .Y(_03913_),
    .A2(net5148));
 sg13g2_a22oi_1 _12471_ (.Y(_03914_),
    .B1(_03912_),
    .B2(_03913_),
    .A2(_03911_),
    .A1(_03910_));
 sg13g2_a21oi_1 _12472_ (.A1(net4385),
    .A2(_03914_),
    .Y(_03915_),
    .B1(net4723));
 sg13g2_a22oi_1 _12473_ (.Y(_00202_),
    .B1(_03909_),
    .B2(_03915_),
    .A2(net4723),
    .A1(net5195));
 sg13g2_o21ai_1 _12474_ (.B1(_03785_),
    .Y(_03916_),
    .A1(net5248),
    .A2(_03258_));
 sg13g2_xnor2_1 _12475_ (.Y(_03917_),
    .A(_03282_),
    .B(_03916_));
 sg13g2_nand2_1 _12476_ (.Y(_03918_),
    .A(net5164),
    .B(_03917_));
 sg13g2_nor2_1 _12477_ (.A(net4935),
    .B(_03739_),
    .Y(_03919_));
 sg13g2_a21oi_2 _12478_ (.B1(_03919_),
    .Y(_03920_),
    .A2(_03731_),
    .A1(net4936));
 sg13g2_nand2_1 _12479_ (.Y(_03921_),
    .A(net4775),
    .B(_03920_));
 sg13g2_nor3_1 _12480_ (.A(net4945),
    .B(net4914),
    .C(_03585_),
    .Y(_03922_));
 sg13g2_o21ai_1 _12481_ (.B1(_03921_),
    .Y(_03923_),
    .A1(net4775),
    .A2(_03922_));
 sg13g2_a21oi_1 _12482_ (.A1(net4941),
    .A2(_03751_),
    .Y(_03924_),
    .B1(net4955));
 sg13g2_o21ai_1 _12483_ (.B1(_03924_),
    .Y(_03925_),
    .A1(net4941),
    .A2(_03745_));
 sg13g2_and2_1 _12484_ (.A(net4940),
    .B(_03732_),
    .X(_03926_));
 sg13g2_a21oi_1 _12485_ (.A1(net4937),
    .A2(_03749_),
    .Y(_03927_),
    .B1(_03926_));
 sg13g2_a21oi_1 _12486_ (.A1(net4949),
    .A2(_03927_),
    .Y(_03928_),
    .B1(net4762));
 sg13g2_a221oi_1 _12487_ (.B2(_03928_),
    .C1(_03607_),
    .B1(_03925_),
    .A1(net4769),
    .Y(_03929_),
    .A2(_03923_));
 sg13g2_and2_1 _12488_ (.A(net4888),
    .B(_03757_),
    .X(_03930_));
 sg13g2_a21oi_1 _12489_ (.A1(net4906),
    .A2(_03280_),
    .Y(_03931_),
    .B1(_03608_));
 sg13g2_mux2_1 _12490_ (.A0(_03846_),
    .A1(_03931_),
    .S(net4928),
    .X(_03932_));
 sg13g2_a21oi_1 _12491_ (.A1(net4771),
    .A2(_03932_),
    .Y(_03933_),
    .B1(_03930_));
 sg13g2_nor2_1 _12492_ (.A(net4952),
    .B(_03933_),
    .Y(_03934_));
 sg13g2_nor2_1 _12493_ (.A(_03803_),
    .B(_03934_),
    .Y(_03935_));
 sg13g2_nor2_1 _12494_ (.A(net5253),
    .B(_03934_),
    .Y(_03936_));
 sg13g2_a221oi_1 _12495_ (.B2(net4892),
    .C1(_03936_),
    .B1(_03935_),
    .A1(net4761),
    .Y(_03937_),
    .A2(_03484_));
 sg13g2_o21ai_1 _12496_ (.B1(net5173),
    .Y(_03938_),
    .A1(net5305),
    .A2(_03282_));
 sg13g2_nor2_1 _12497_ (.A(_03937_),
    .B(_03938_),
    .Y(_03939_));
 sg13g2_nand2_1 _12498_ (.Y(_03940_),
    .A(net5164),
    .B(_03281_));
 sg13g2_nand3_1 _12499_ (.B(_03278_),
    .C(_03940_),
    .A(net5290),
    .Y(_03941_));
 sg13g2_nor2b_1 _12500_ (.A(_03939_),
    .B_N(_03941_),
    .Y(_03942_));
 sg13g2_a22oi_1 _12501_ (.Y(_03943_),
    .B1(_03942_),
    .B2(net5257),
    .A2(_03929_),
    .A1(_03918_));
 sg13g2_nand2b_1 _12502_ (.Y(_03944_),
    .B(\m_sys._m_ram_io_b_port_rdata[24] ),
    .A_N(net5362));
 sg13g2_nand3_1 _12503_ (.B(net4497),
    .C(net5071),
    .A(\m_sys._m_ram_io_b_port_rdata[24] ),
    .Y(_03945_));
 sg13g2_o21ai_1 _12504_ (.B1(_03945_),
    .Y(_03946_),
    .A1(_03820_),
    .A2(_03944_));
 sg13g2_nand2b_2 _12505_ (.Y(_03947_),
    .B(_03946_),
    .A_N(net4745));
 sg13g2_a221oi_1 _12506_ (.B2(net4038),
    .C1(net4751),
    .B1(_03947_),
    .A1(net5100),
    .Y(_03948_),
    .A2(_03943_));
 sg13g2_nand2_1 _12507_ (.Y(_03949_),
    .A(\m_sys.m_core.m_gpr._GEN[120] ),
    .B(net5059));
 sg13g2_a221oi_1 _12508_ (.B2(net5050),
    .C1(net5328),
    .B1(\m_sys.m_core.m_gpr._GEN[88] ),
    .A1(net5184),
    .Y(_03950_),
    .A2(\m_sys.m_core.m_gpr._GEN[56] ));
 sg13g2_a22oi_1 _12509_ (.Y(_03951_),
    .B1(net5046),
    .B2(\m_sys.m_core.m_gpr._GEN[184] ),
    .A2(net5059),
    .A1(\m_sys.m_core.m_gpr._GEN[248] ));
 sg13g2_a221oi_1 _12510_ (.B2(\m_sys.m_core.m_gpr._GEN[216] ),
    .C1(net5178),
    .B1(net5050),
    .A1(\m_sys.m_core.m_gpr._GEN[152] ),
    .Y(_03952_),
    .A2(net5148));
 sg13g2_a221oi_1 _12511_ (.B2(_03952_),
    .C1(_03560_),
    .B1(_03951_),
    .A1(_03949_),
    .Y(_03953_),
    .A2(_03950_));
 sg13g2_nor3_1 _12512_ (.A(net4726),
    .B(_03948_),
    .C(_03953_),
    .Y(_03954_));
 sg13g2_a21oi_1 _12513_ (.A1(net5196),
    .A2(net4726),
    .Y(_00203_),
    .B1(_03954_));
 sg13g2_o21ai_1 _12514_ (.B1(_03251_),
    .Y(_03955_),
    .A1(_03193_),
    .A2(_03247_));
 sg13g2_a221oi_1 _12515_ (.B2(_03955_),
    .C1(_03214_),
    .B1(_03220_),
    .A1(_03209_),
    .Y(_03956_),
    .A2(_03217_));
 sg13g2_o21ai_1 _12516_ (.B1(_03205_),
    .Y(_03957_),
    .A1(_03204_),
    .A2(_03956_));
 sg13g2_o21ai_1 _12517_ (.B1(_03375_),
    .Y(_03958_),
    .A1(_03364_),
    .A2(_03368_));
 sg13g2_nand3b_1 _12518_ (.B(_03219_),
    .C(_03958_),
    .Y(_03959_),
    .A_N(_03212_));
 sg13g2_nand2b_1 _12519_ (.Y(_03960_),
    .B(net5251),
    .A_N(_03364_));
 sg13g2_inv_1 _12520_ (.Y(_03961_),
    .A(_03960_));
 sg13g2_nand2_1 _12521_ (.Y(_03962_),
    .A(net5251),
    .B(_03958_));
 sg13g2_a21oi_1 _12522_ (.A1(_03378_),
    .A2(_03959_),
    .Y(_03963_),
    .B1(net5167));
 sg13g2_a22oi_1 _12523_ (.Y(_03964_),
    .B1(_03963_),
    .B2(_03207_),
    .A2(_03379_),
    .A1(net5249));
 sg13g2_o21ai_1 _12524_ (.B1(_03964_),
    .Y(_03965_),
    .A1(net5249),
    .A2(_03957_));
 sg13g2_xor2_1 _12525_ (.B(_03965_),
    .A(_03200_),
    .X(_03966_));
 sg13g2_nand2_1 _12526_ (.Y(_03967_),
    .A(net4951),
    .B(_03424_));
 sg13g2_a21oi_1 _12527_ (.A1(net4779),
    .A2(_03478_),
    .Y(_03968_),
    .B1(net4762));
 sg13g2_nand2_1 _12528_ (.Y(_03969_),
    .A(net4768),
    .B(_03606_));
 sg13g2_or2_1 _12529_ (.X(_03970_),
    .B(_03438_),
    .A(net4951));
 sg13g2_a221oi_1 _12530_ (.B2(net4770),
    .C1(_03607_),
    .B1(_03970_),
    .A1(_03967_),
    .Y(_03971_),
    .A2(_03968_));
 sg13g2_o21ai_1 _12531_ (.B1(_03971_),
    .Y(_03972_),
    .A1(net5304),
    .A2(_03966_));
 sg13g2_o21ai_1 _12532_ (.B1(_03468_),
    .Y(_03973_),
    .A1(net4908),
    .A2(_03280_));
 sg13g2_mux2_1 _12533_ (.A0(_03888_),
    .A1(_03973_),
    .S(net4932),
    .X(_03974_));
 sg13g2_mux2_1 _12534_ (.A0(_03806_),
    .A1(_03974_),
    .S(net4771),
    .X(_03975_));
 sg13g2_and2_1 _12535_ (.A(net4781),
    .B(_03975_),
    .X(_03976_));
 sg13g2_nor2_1 _12536_ (.A(_03803_),
    .B(_03976_),
    .Y(_03977_));
 sg13g2_nor3_1 _12537_ (.A(net4781),
    .B(net4943),
    .C(_03458_),
    .Y(_03978_));
 sg13g2_nor3_1 _12538_ (.A(net5253),
    .B(_03976_),
    .C(_03978_),
    .Y(_03979_));
 sg13g2_a221oi_1 _12539_ (.B2(net4892),
    .C1(_03979_),
    .B1(_03977_),
    .A1(net4764),
    .Y(_03980_),
    .A2(_03484_));
 sg13g2_o21ai_1 _12540_ (.B1(net5173),
    .Y(_03981_),
    .A1(net5305),
    .A2(_03200_));
 sg13g2_nor2_1 _12541_ (.A(_03980_),
    .B(_03981_),
    .Y(_03982_));
 sg13g2_nor2_1 _12542_ (.A(net5305),
    .B(_03199_),
    .Y(_03983_));
 sg13g2_nand2_1 _12543_ (.Y(_03984_),
    .A(net5290),
    .B(_03196_));
 sg13g2_o21ai_1 _12544_ (.B1(net5257),
    .Y(_03985_),
    .A1(_03983_),
    .A2(_03984_));
 sg13g2_o21ai_1 _12545_ (.B1(_03972_),
    .Y(_03986_),
    .A1(_03982_),
    .A2(_03985_));
 sg13g2_and2_1 _12546_ (.A(\m_sys._m_ram_io_b_port_rdata[23] ),
    .B(net5070),
    .X(_03987_));
 sg13g2_a22oi_1 _12547_ (.Y(_03988_),
    .B1(_03987_),
    .B2(net4496),
    .A2(net4740),
    .A1(_03502_));
 sg13g2_or2_2 _12548_ (.X(_03989_),
    .B(_03988_),
    .A(net4746));
 sg13g2_a21oi_1 _12549_ (.A1(net4038),
    .A2(_03989_),
    .Y(_03990_),
    .B1(net4752));
 sg13g2_o21ai_1 _12550_ (.B1(_03990_),
    .Y(_03991_),
    .A1(net5098),
    .A2(_03986_));
 sg13g2_nand2_1 _12551_ (.Y(_03992_),
    .A(\m_sys.m_core.m_gpr._GEN[119] ),
    .B(net5063));
 sg13g2_a221oi_1 _12552_ (.B2(net5054),
    .C1(net5331),
    .B1(\m_sys.m_core.m_gpr._GEN[87] ),
    .A1(net5190),
    .Y(_03993_),
    .A2(\m_sys.m_core.m_gpr._GEN[55] ));
 sg13g2_a22oi_1 _12553_ (.Y(_03994_),
    .B1(net5048),
    .B2(\m_sys.m_core.m_gpr._GEN[183] ),
    .A2(net5063),
    .A1(\m_sys.m_core.m_gpr._GEN[247] ));
 sg13g2_a221oi_1 _12554_ (.B2(\m_sys.m_core.m_gpr._GEN[215] ),
    .C1(net5180),
    .B1(net5054),
    .A1(\m_sys.m_core.m_gpr._GEN[151] ),
    .Y(_03995_),
    .A2(net5150));
 sg13g2_a22oi_1 _12555_ (.Y(_03996_),
    .B1(_03994_),
    .B2(_03995_),
    .A2(_03993_),
    .A1(_03992_));
 sg13g2_a21oi_1 _12556_ (.A1(net4385),
    .A2(_03996_),
    .Y(_03997_),
    .B1(net4724));
 sg13g2_a22oi_1 _12557_ (.Y(_00204_),
    .B1(_03991_),
    .B2(_03997_),
    .A2(net4726),
    .A1(net5197));
 sg13g2_a21oi_1 _12558_ (.A1(net5167),
    .A2(_03956_),
    .Y(_03998_),
    .B1(_03963_));
 sg13g2_a21oi_1 _12559_ (.A1(_03207_),
    .A2(_03998_),
    .Y(_03999_),
    .B1(net5304));
 sg13g2_o21ai_1 _12560_ (.B1(_03999_),
    .Y(_04000_),
    .A1(_03207_),
    .A2(_03998_));
 sg13g2_nand2_1 _12561_ (.Y(_04001_),
    .A(net4949),
    .B(_03604_));
 sg13g2_a21oi_1 _12562_ (.A1(net4779),
    .A2(_03638_),
    .Y(_04002_),
    .B1(net4762));
 sg13g2_nand2_1 _12563_ (.Y(_04003_),
    .A(net4767),
    .B(_03442_));
 sg13g2_or2_1 _12564_ (.X(_04004_),
    .B(_03587_),
    .A(net4946));
 sg13g2_a221oi_1 _12565_ (.B2(net4769),
    .C1(_03443_),
    .B1(_04004_),
    .A1(_04001_),
    .Y(_04005_),
    .A2(_04002_));
 sg13g2_nor2_1 _12566_ (.A(_03612_),
    .B(_03623_),
    .Y(_04006_));
 sg13g2_mux2_1 _12567_ (.A0(_03931_),
    .A1(_04006_),
    .S(net4932),
    .X(_04007_));
 sg13g2_mux2_1 _12568_ (.A0(_03847_),
    .A1(_04007_),
    .S(net4771),
    .X(_04008_));
 sg13g2_nor2_1 _12569_ (.A(net4952),
    .B(_04008_),
    .Y(_04009_));
 sg13g2_a21oi_1 _12570_ (.A1(net4952),
    .A2(_03649_),
    .Y(_04010_),
    .B1(_04009_));
 sg13g2_nor2_1 _12571_ (.A(net5168),
    .B(_04010_),
    .Y(_04011_));
 sg13g2_o21ai_1 _12572_ (.B1(net4952),
    .Y(_04012_),
    .A1(net4943),
    .A2(_03646_));
 sg13g2_o21ai_1 _12573_ (.B1(_04012_),
    .Y(_04013_),
    .A1(net4952),
    .A2(_04008_));
 sg13g2_and2_1 _12574_ (.A(net5168),
    .B(_04013_),
    .X(_04014_));
 sg13g2_a21o_1 _12575_ (.A2(_04011_),
    .A1(net4892),
    .B1(_03485_),
    .X(_04015_));
 sg13g2_a21oi_1 _12576_ (.A1(net5164),
    .A2(_03206_),
    .Y(_04016_),
    .B1(net5289));
 sg13g2_o21ai_1 _12577_ (.B1(_04016_),
    .Y(_04017_),
    .A1(_04014_),
    .A2(_04015_));
 sg13g2_nand2_1 _12578_ (.Y(_04018_),
    .A(net5164),
    .B(_03203_));
 sg13g2_and2_1 _12579_ (.A(net5289),
    .B(_03205_),
    .X(_04019_));
 sg13g2_a21oi_1 _12580_ (.A1(_04018_),
    .A2(_04019_),
    .Y(_04020_),
    .B1(_02496_));
 sg13g2_a22oi_1 _12581_ (.Y(_04021_),
    .B1(_04017_),
    .B2(_04020_),
    .A2(_04005_),
    .A1(_04000_));
 sg13g2_mux2_1 _12582_ (.A0(\m_sys._m_ram_io_b_port_rdata[22] ),
    .A1(\m_sys._m_ram_io_b_port_rdata[30] ),
    .S(net5360),
    .X(_04022_));
 sg13g2_and2_1 _12583_ (.A(\m_sys._m_ram_io_b_port_rdata[22] ),
    .B(net5069),
    .X(_04023_));
 sg13g2_a22oi_1 _12584_ (.Y(_04024_),
    .B1(_04023_),
    .B2(net4497),
    .A2(_04022_),
    .A1(net4740));
 sg13g2_or2_2 _12585_ (.X(_04025_),
    .B(_04024_),
    .A(net4747));
 sg13g2_a221oi_1 _12586_ (.B2(net4038),
    .C1(net4752),
    .B1(_04025_),
    .A1(net5099),
    .Y(_04026_),
    .A2(_04021_));
 sg13g2_nand2_1 _12587_ (.Y(_04027_),
    .A(\m_sys.m_core.m_gpr._GEN[118] ),
    .B(net5064));
 sg13g2_a221oi_1 _12588_ (.B2(net5058),
    .C1(net5329),
    .B1(\m_sys.m_core.m_gpr._GEN[86] ),
    .A1(net5186),
    .Y(_04028_),
    .A2(\m_sys.m_core.m_gpr._GEN[54] ));
 sg13g2_a22oi_1 _12589_ (.Y(_04029_),
    .B1(net5048),
    .B2(\m_sys.m_core.m_gpr._GEN[182] ),
    .A2(net5064),
    .A1(\m_sys.m_core.m_gpr._GEN[246] ));
 sg13g2_a221oi_1 _12590_ (.B2(\m_sys.m_core.m_gpr._GEN[214] ),
    .C1(net5180),
    .B1(net5054),
    .A1(\m_sys.m_core.m_gpr._GEN[150] ),
    .Y(_04030_),
    .A2(net5150));
 sg13g2_a221oi_1 _12591_ (.B2(_04030_),
    .C1(_03560_),
    .B1(_04029_),
    .A1(_04027_),
    .Y(_04031_),
    .A2(_04028_));
 sg13g2_nor3_1 _12592_ (.A(net4725),
    .B(_04026_),
    .C(_04031_),
    .Y(_04032_));
 sg13g2_a21oi_1 _12593_ (.A1(net5208),
    .A2(net4725),
    .Y(_00205_),
    .B1(_04032_));
 sg13g2_nand2b_1 _12594_ (.Y(_04033_),
    .B(_03955_),
    .A_N(_03211_));
 sg13g2_nor2_1 _12595_ (.A(net5249),
    .B(_03209_),
    .Y(_04034_));
 sg13g2_nor2_1 _12596_ (.A(_03212_),
    .B(_03962_),
    .Y(_04035_));
 sg13g2_a221oi_1 _12597_ (.B2(_04034_),
    .C1(_04035_),
    .B1(_04033_),
    .A1(net5248),
    .Y(_04036_),
    .A2(_03377_));
 sg13g2_xnor2_1 _12598_ (.Y(_04037_),
    .A(_03218_),
    .B(_04036_));
 sg13g2_nor2_1 _12599_ (.A(net4780),
    .B(_03686_),
    .Y(_04038_));
 sg13g2_o21ai_1 _12600_ (.B1(net4765),
    .Y(_04039_),
    .A1(net4951),
    .A2(_03696_));
 sg13g2_nand2_1 _12601_ (.Y(_04040_),
    .A(net4778),
    .B(_03682_));
 sg13g2_a21oi_1 _12602_ (.A1(net4770),
    .A2(_04040_),
    .Y(_04041_),
    .B1(_03443_));
 sg13g2_o21ai_1 _12603_ (.B1(_04041_),
    .Y(_04042_),
    .A1(_04038_),
    .A2(_04039_));
 sg13g2_a21oi_1 _12604_ (.A1(net5165),
    .A2(_04037_),
    .Y(_04043_),
    .B1(_04042_));
 sg13g2_o21ai_1 _12605_ (.B1(_03473_),
    .Y(_04044_),
    .A1(net4908),
    .A2(_03201_));
 sg13g2_nor2_1 _12606_ (.A(net4921),
    .B(_04044_),
    .Y(_04045_));
 sg13g2_and2_1 _12607_ (.A(net4920),
    .B(_03973_),
    .X(_04046_));
 sg13g2_nor2_1 _12608_ (.A(_04045_),
    .B(_04046_),
    .Y(_04047_));
 sg13g2_nand2_1 _12609_ (.Y(_04048_),
    .A(net4889),
    .B(_03890_));
 sg13g2_o21ai_1 _12610_ (.B1(_04048_),
    .Y(_04049_),
    .A1(net4888),
    .A2(_04047_));
 sg13g2_nand2b_1 _12611_ (.Y(_04050_),
    .B(net4783),
    .A_N(_04049_));
 sg13g2_o21ai_1 _12612_ (.B1(_04050_),
    .Y(_04051_),
    .A1(net4783),
    .A2(_03702_));
 sg13g2_nand3_1 _12613_ (.B(net4892),
    .C(_04051_),
    .A(net5250),
    .Y(_04052_));
 sg13g2_nand2_1 _12614_ (.Y(_04053_),
    .A(net4953),
    .B(_03707_));
 sg13g2_a21o_1 _12615_ (.A2(_04053_),
    .A1(_04050_),
    .B1(net5253),
    .X(_04054_));
 sg13g2_and2_1 _12616_ (.A(_03486_),
    .B(_04054_),
    .X(_04055_));
 sg13g2_a221oi_1 _12617_ (.B2(_04055_),
    .C1(net5291),
    .B1(_04052_),
    .A1(net5165),
    .Y(_04056_),
    .A2(_03218_));
 sg13g2_a21oi_1 _12618_ (.A1(_03213_),
    .A2(_03215_),
    .Y(_04057_),
    .B1(net5305));
 sg13g2_nor3_1 _12619_ (.A(net5173),
    .B(_03214_),
    .C(_04057_),
    .Y(_04058_));
 sg13g2_nor3_1 _12620_ (.A(_02496_),
    .B(_04056_),
    .C(_04058_),
    .Y(_04059_));
 sg13g2_nor2_2 _12621_ (.A(_04043_),
    .B(_04059_),
    .Y(_04060_));
 sg13g2_mux2_1 _12622_ (.A0(\m_sys._m_ram_io_b_port_rdata[21] ),
    .A1(\m_sys._m_ram_io_b_port_rdata[29] ),
    .S(net5364),
    .X(_04061_));
 sg13g2_and2_1 _12623_ (.A(\m_sys._m_ram_io_b_port_rdata[21] ),
    .B(net5070),
    .X(_04062_));
 sg13g2_a22oi_1 _12624_ (.Y(_04063_),
    .B1(_04062_),
    .B2(net4495),
    .A2(_04061_),
    .A1(_03819_));
 sg13g2_or2_2 _12625_ (.X(_04064_),
    .B(_04063_),
    .A(net4746));
 sg13g2_a221oi_1 _12626_ (.B2(net4038),
    .C1(net4751),
    .B1(_04064_),
    .A1(net5099),
    .Y(_04065_),
    .A2(_04060_));
 sg13g2_nand2_1 _12627_ (.Y(_04066_),
    .A(\m_sys.m_core.m_gpr._GEN[117] ),
    .B(net5064));
 sg13g2_a221oi_1 _12628_ (.B2(net5058),
    .C1(net5329),
    .B1(\m_sys.m_core.m_gpr._GEN[85] ),
    .A1(net5186),
    .Y(_04067_),
    .A2(\m_sys.m_core.m_gpr._GEN[53] ));
 sg13g2_a22oi_1 _12629_ (.Y(_04068_),
    .B1(net5048),
    .B2(\m_sys.m_core.m_gpr._GEN[181] ),
    .A2(net5064),
    .A1(\m_sys.m_core.m_gpr._GEN[245] ));
 sg13g2_a221oi_1 _12630_ (.B2(\m_sys.m_core.m_gpr._GEN[213] ),
    .C1(net5180),
    .B1(net5058),
    .A1(\m_sys.m_core.m_gpr._GEN[149] ),
    .Y(_04069_),
    .A2(net5150));
 sg13g2_a221oi_1 _12631_ (.B2(_04069_),
    .C1(_03560_),
    .B1(_04068_),
    .A1(_04066_),
    .Y(_04070_),
    .A2(_04067_));
 sg13g2_nor3_1 _12632_ (.A(net4725),
    .B(_04065_),
    .C(_04070_),
    .Y(_04071_));
 sg13g2_a21oi_1 _12633_ (.A1(net5218),
    .A2(net4725),
    .Y(_00206_),
    .B1(_04071_));
 sg13g2_o21ai_1 _12634_ (.B1(_03962_),
    .Y(_04072_),
    .A1(net5248),
    .A2(_03955_));
 sg13g2_xnor2_1 _12635_ (.Y(_04073_),
    .A(_03212_),
    .B(_04072_));
 sg13g2_nor2_1 _12636_ (.A(net4780),
    .B(_03734_),
    .Y(_04074_));
 sg13g2_o21ai_1 _12637_ (.B1(net4765),
    .Y(_04075_),
    .A1(net4950),
    .A2(_03752_));
 sg13g2_nor2_1 _12638_ (.A(_04074_),
    .B(_04075_),
    .Y(_04076_));
 sg13g2_and2_1 _12639_ (.A(net4778),
    .B(_03740_),
    .X(_04077_));
 sg13g2_o21ai_1 _12640_ (.B1(_03606_),
    .Y(_04078_),
    .A1(net4768),
    .A2(_04077_));
 sg13g2_nor2_2 _12641_ (.A(_04076_),
    .B(_04078_),
    .Y(_04079_));
 sg13g2_o21ai_1 _12642_ (.B1(_04079_),
    .Y(_04080_),
    .A1(net5307),
    .A2(_04073_));
 sg13g2_o21ai_1 _12643_ (.B1(_03626_),
    .Y(_04081_),
    .A1(net4908),
    .A2(_03216_));
 sg13g2_nor2_1 _12644_ (.A(net4921),
    .B(_04081_),
    .Y(_04082_));
 sg13g2_a21oi_1 _12645_ (.A1(net4920),
    .A2(_04006_),
    .Y(_04083_),
    .B1(_04082_));
 sg13g2_nor2_1 _12646_ (.A(net4890),
    .B(_04083_),
    .Y(_04084_));
 sg13g2_a21oi_2 _12647_ (.B1(_04084_),
    .Y(_04085_),
    .A2(_03932_),
    .A1(net4890));
 sg13g2_nand2_1 _12648_ (.Y(_04086_),
    .A(net4782),
    .B(_04085_));
 sg13g2_o21ai_1 _12649_ (.B1(net4952),
    .Y(_04087_),
    .A1(_03643_),
    .A2(_03758_));
 sg13g2_a21oi_1 _12650_ (.A1(_04086_),
    .A2(_04087_),
    .Y(_04088_),
    .B1(net5168));
 sg13g2_nand2_1 _12651_ (.Y(_04089_),
    .A(net4952),
    .B(_03762_));
 sg13g2_a21oi_1 _12652_ (.A1(_04086_),
    .A2(_04089_),
    .Y(_04090_),
    .B1(net5250));
 sg13g2_a21o_1 _12653_ (.A2(_04088_),
    .A1(net4892),
    .B1(_03485_),
    .X(_04091_));
 sg13g2_a21oi_1 _12654_ (.A1(net5165),
    .A2(_03212_),
    .Y(_04092_),
    .B1(net5291));
 sg13g2_o21ai_1 _12655_ (.B1(_04092_),
    .Y(_04093_),
    .A1(_04090_),
    .A2(_04091_));
 sg13g2_nor2_1 _12656_ (.A(net5173),
    .B(_03209_),
    .Y(_04094_));
 sg13g2_o21ai_1 _12657_ (.B1(_04094_),
    .Y(_04095_),
    .A1(net5308),
    .A2(_03211_));
 sg13g2_nand3_1 _12658_ (.B(_04093_),
    .C(_04095_),
    .A(net5258),
    .Y(_04096_));
 sg13g2_and2_1 _12659_ (.A(_04080_),
    .B(_04096_),
    .X(_04097_));
 sg13g2_mux2_1 _12660_ (.A0(\m_sys._m_ram_io_b_port_rdata[20] ),
    .A1(\m_sys._m_ram_io_b_port_rdata[28] ),
    .S(net5363),
    .X(_04098_));
 sg13g2_and2_1 _12661_ (.A(\m_sys._m_ram_io_b_port_rdata[20] ),
    .B(net5071),
    .X(_04099_));
 sg13g2_a22oi_1 _12662_ (.Y(_04100_),
    .B1(_04099_),
    .B2(net4496),
    .A2(_04098_),
    .A1(net4740));
 sg13g2_or2_2 _12663_ (.X(_04101_),
    .B(_04100_),
    .A(net4745));
 sg13g2_a221oi_1 _12664_ (.B2(net4038),
    .C1(net4751),
    .B1(_04101_),
    .A1(net5100),
    .Y(_04102_),
    .A2(_04097_));
 sg13g2_nand2_1 _12665_ (.Y(_04103_),
    .A(\m_sys.m_core.m_gpr._GEN[116] ),
    .B(net5063));
 sg13g2_a221oi_1 _12666_ (.B2(net5054),
    .C1(net5329),
    .B1(\m_sys.m_core.m_gpr._GEN[84] ),
    .A1(net5186),
    .Y(_04104_),
    .A2(\m_sys.m_core.m_gpr._GEN[52] ));
 sg13g2_a22oi_1 _12667_ (.Y(_04105_),
    .B1(net5048),
    .B2(\m_sys.m_core.m_gpr._GEN[180] ),
    .A2(net5063),
    .A1(\m_sys.m_core.m_gpr._GEN[244] ));
 sg13g2_a221oi_1 _12668_ (.B2(\m_sys.m_core.m_gpr._GEN[212] ),
    .C1(net5180),
    .B1(net5054),
    .A1(\m_sys.m_core.m_gpr._GEN[148] ),
    .Y(_04106_),
    .A2(net5150));
 sg13g2_a221oi_1 _12669_ (.B2(_04106_),
    .C1(_03560_),
    .B1(_04105_),
    .A1(_04103_),
    .Y(_04107_),
    .A2(_04104_));
 sg13g2_nor3_1 _12670_ (.A(net4724),
    .B(_04102_),
    .C(_04107_),
    .Y(_04108_));
 sg13g2_a21oi_1 _12671_ (.A1(net5198),
    .A2(net4724),
    .Y(_00207_),
    .B1(_04108_));
 sg13g2_a21oi_1 _12672_ (.A1(_03194_),
    .A2(_03246_),
    .Y(_04109_),
    .B1(_03249_));
 sg13g2_o21ai_1 _12673_ (.B1(_03228_),
    .Y(_04110_),
    .A1(_03232_),
    .A2(_04109_));
 sg13g2_nand2_1 _12674_ (.Y(_04111_),
    .A(net5252),
    .B(_03372_));
 sg13g2_o21ai_1 _12675_ (.B1(_04111_),
    .Y(_04112_),
    .A1(_03367_),
    .A2(_03960_));
 sg13g2_nor2b_1 _12676_ (.A(_03233_),
    .B_N(_04112_),
    .Y(_04113_));
 sg13g2_a21oi_1 _12677_ (.A1(net5252),
    .A2(_03374_),
    .Y(_04114_),
    .B1(_04113_));
 sg13g2_o21ai_1 _12678_ (.B1(_04114_),
    .Y(_04115_),
    .A1(net5252),
    .A2(_04110_));
 sg13g2_xnor2_1 _12679_ (.Y(_04116_),
    .A(_03225_),
    .B(_04115_));
 sg13g2_nand2b_1 _12680_ (.Y(_04117_),
    .B(net4949),
    .A_N(_03792_));
 sg13g2_a21oi_1 _12681_ (.A1(net4785),
    .A2(_03799_),
    .Y(_04118_),
    .B1(net4763));
 sg13g2_nand2_1 _12682_ (.Y(_04119_),
    .A(net4775),
    .B(_03794_));
 sg13g2_a221oi_1 _12683_ (.B2(net4769),
    .C1(_03443_),
    .B1(_04119_),
    .A1(_04117_),
    .Y(_04120_),
    .A2(_04118_));
 sg13g2_o21ai_1 _12684_ (.B1(_04120_),
    .Y(_04121_),
    .A1(net5308),
    .A2(_04116_));
 sg13g2_nand2_1 _12685_ (.Y(_04122_),
    .A(_03462_),
    .B(_03472_));
 sg13g2_mux2_1 _12686_ (.A0(_04044_),
    .A1(_04122_),
    .S(net4931),
    .X(_04123_));
 sg13g2_nand2_1 _12687_ (.Y(_04124_),
    .A(net4772),
    .B(_04123_));
 sg13g2_o21ai_1 _12688_ (.B1(_04124_),
    .Y(_04125_),
    .A1(net4772),
    .A2(_03974_));
 sg13g2_nand2_1 _12689_ (.Y(_04126_),
    .A(net4784),
    .B(_04125_));
 sg13g2_o21ai_1 _12690_ (.B1(_04126_),
    .Y(_04127_),
    .A1(net4782),
    .A2(_03808_));
 sg13g2_and2_1 _12691_ (.A(net5252),
    .B(_04127_),
    .X(_04128_));
 sg13g2_nand2_1 _12692_ (.Y(_04129_),
    .A(net4893),
    .B(_04128_));
 sg13g2_o21ai_1 _12693_ (.B1(_04126_),
    .Y(_04130_),
    .A1(net4782),
    .A2(_03811_));
 sg13g2_and2_1 _12694_ (.A(net5167),
    .B(_04130_),
    .X(_04131_));
 sg13g2_nor2_1 _12695_ (.A(_03485_),
    .B(_04131_),
    .Y(_04132_));
 sg13g2_a221oi_1 _12696_ (.B2(_04132_),
    .C1(net5291),
    .B1(_04129_),
    .A1(net5165),
    .Y(_04133_),
    .A2(_03225_));
 sg13g2_a21oi_1 _12697_ (.A1(_03223_),
    .A2(_03224_),
    .Y(_04134_),
    .B1(net5307));
 sg13g2_o21ai_1 _12698_ (.B1(net5291),
    .Y(_04135_),
    .A1(_00086_),
    .A2(_03224_));
 sg13g2_o21ai_1 _12699_ (.B1(net5258),
    .Y(_04136_),
    .A1(_04134_),
    .A2(_04135_));
 sg13g2_o21ai_1 _12700_ (.B1(_04121_),
    .Y(_04137_),
    .A1(_04133_),
    .A2(_04136_));
 sg13g2_mux2_1 _12701_ (.A0(\m_sys._m_ram_io_b_port_rdata[19] ),
    .A1(\m_sys._m_ram_io_b_port_rdata[27] ),
    .S(net5364),
    .X(_04138_));
 sg13g2_and2_1 _12702_ (.A(\m_sys._m_ram_io_b_port_rdata[19] ),
    .B(net5070),
    .X(_04139_));
 sg13g2_a22oi_1 _12703_ (.Y(_04140_),
    .B1(_04139_),
    .B2(net4495),
    .A2(_04138_),
    .A1(net4740));
 sg13g2_or2_1 _12704_ (.X(_04141_),
    .B(_04140_),
    .A(net4746));
 sg13g2_a21oi_2 _12705_ (.B1(net4748),
    .Y(_04142_),
    .A2(_04141_),
    .A1(net4040));
 sg13g2_o21ai_1 _12706_ (.B1(_04142_),
    .Y(_04143_),
    .A1(net5098),
    .A2(_04137_));
 sg13g2_nand2_1 _12707_ (.Y(_04144_),
    .A(\m_sys.m_core.m_gpr._GEN[115] ),
    .B(net5067));
 sg13g2_a221oi_1 _12708_ (.B2(net5056),
    .C1(net5330),
    .B1(\m_sys.m_core.m_gpr._GEN[83] ),
    .A1(net5187),
    .Y(_04145_),
    .A2(\m_sys.m_core.m_gpr._GEN[51] ));
 sg13g2_a22oi_1 _12709_ (.Y(_04146_),
    .B1(net5047),
    .B2(\m_sys.m_core.m_gpr._GEN[179] ),
    .A2(net5067),
    .A1(\m_sys.m_core.m_gpr._GEN[243] ));
 sg13g2_a221oi_1 _12710_ (.B2(\m_sys.m_core.m_gpr._GEN[211] ),
    .C1(net5182),
    .B1(net5056),
    .A1(\m_sys.m_core.m_gpr._GEN[147] ),
    .Y(_04147_),
    .A2(net5150));
 sg13g2_a22oi_1 _12711_ (.Y(_04148_),
    .B1(_04146_),
    .B2(_04147_),
    .A2(_04145_),
    .A1(_04144_));
 sg13g2_a21oi_1 _12712_ (.A1(net4385),
    .A2(_04148_),
    .Y(_04149_),
    .B1(net4727));
 sg13g2_a22oi_1 _12713_ (.Y(_00208_),
    .B1(_04143_),
    .B2(_04149_),
    .A2(net4728),
    .A1(net5176));
 sg13g2_a21oi_1 _12714_ (.A1(net5168),
    .A2(_04109_),
    .Y(_04150_),
    .B1(_04112_));
 sg13g2_xnor2_1 _12715_ (.Y(_04151_),
    .A(_03233_),
    .B(_04150_));
 sg13g2_nand2_1 _12716_ (.Y(_04152_),
    .A(net5165),
    .B(_04151_));
 sg13g2_nand2b_1 _12717_ (.Y(_04153_),
    .B(net4949),
    .A_N(_03837_));
 sg13g2_a21oi_1 _12718_ (.A1(net4780),
    .A2(_03843_),
    .Y(_04154_),
    .B1(net4762));
 sg13g2_nand3_1 _12719_ (.B(net4936),
    .C(_03586_),
    .A(net4777),
    .Y(_04155_));
 sg13g2_a221oi_1 _12720_ (.B2(net4769),
    .C1(_03607_),
    .B1(_04155_),
    .A1(_04153_),
    .Y(_04156_),
    .A2(_04154_));
 sg13g2_a21oi_1 _12721_ (.A1(_03625_),
    .A2(_03632_),
    .Y(_04157_),
    .B1(net4920));
 sg13g2_a21o_1 _12722_ (.A2(_04081_),
    .A1(net4921),
    .B1(_04157_),
    .X(_04158_));
 sg13g2_nor2_1 _12723_ (.A(net4890),
    .B(_04158_),
    .Y(_04159_));
 sg13g2_a21oi_2 _12724_ (.B1(_04159_),
    .Y(_04160_),
    .A2(_04007_),
    .A1(net4889));
 sg13g2_nand2_1 _12725_ (.Y(_04161_),
    .A(net4782),
    .B(_04160_));
 sg13g2_o21ai_1 _12726_ (.B1(_04161_),
    .Y(_04162_),
    .A1(net4782),
    .A2(_03850_));
 sg13g2_nand3_1 _12727_ (.B(net4893),
    .C(_04162_),
    .A(net5250),
    .Y(_04163_));
 sg13g2_nand2b_1 _12728_ (.Y(_04164_),
    .B(net4956),
    .A_N(_03852_));
 sg13g2_a21oi_1 _12729_ (.A1(_04161_),
    .A2(_04164_),
    .Y(_04165_),
    .B1(net5250));
 sg13g2_nor2_1 _12730_ (.A(_03485_),
    .B(_04165_),
    .Y(_04166_));
 sg13g2_nand2_1 _12731_ (.Y(_04167_),
    .A(_04163_),
    .B(_04166_));
 sg13g2_a21oi_1 _12732_ (.A1(net5165),
    .A2(_03233_),
    .Y(_04168_),
    .B1(net5291));
 sg13g2_o21ai_1 _12733_ (.B1(_03228_),
    .Y(_04169_),
    .A1(net5307),
    .A2(_03232_));
 sg13g2_o21ai_1 _12734_ (.B1(net5258),
    .Y(_04170_),
    .A1(net5174),
    .A2(_04169_));
 sg13g2_a21oi_1 _12735_ (.A1(_04167_),
    .A2(_04168_),
    .Y(_04171_),
    .B1(_04170_));
 sg13g2_a21oi_2 _12736_ (.B1(_04171_),
    .Y(_04172_),
    .A2(_04156_),
    .A1(_04152_));
 sg13g2_nand2_1 _12737_ (.Y(_04173_),
    .A(net5099),
    .B(_04172_));
 sg13g2_mux2_1 _12738_ (.A0(\m_sys._m_ram_io_b_port_rdata[18] ),
    .A1(\m_sys._m_ram_io_b_port_rdata[26] ),
    .S(net5363),
    .X(_04174_));
 sg13g2_and2_1 _12739_ (.A(\m_sys._m_ram_io_b_port_rdata[18] ),
    .B(net5071),
    .X(_04175_));
 sg13g2_a22oi_1 _12740_ (.Y(_04176_),
    .B1(_04175_),
    .B2(net4495),
    .A2(_04174_),
    .A1(net4740));
 sg13g2_o21ai_1 _12741_ (.B1(net4040),
    .Y(_04177_),
    .A1(net4745),
    .A2(_04176_));
 sg13g2_nand3_1 _12742_ (.B(_04173_),
    .C(_04177_),
    .A(net4759),
    .Y(_04178_));
 sg13g2_nand2_1 _12743_ (.Y(_04179_),
    .A(\m_sys.m_core.m_gpr._GEN[114] ),
    .B(net5066));
 sg13g2_a221oi_1 _12744_ (.B2(net5057),
    .C1(net5330),
    .B1(\m_sys.m_core.m_gpr._GEN[82] ),
    .A1(net5189),
    .Y(_04180_),
    .A2(\m_sys.m_core.m_gpr._GEN[50] ));
 sg13g2_a22oi_1 _12745_ (.Y(_04181_),
    .B1(net5047),
    .B2(\m_sys.m_core.m_gpr._GEN[178] ),
    .A2(net5066),
    .A1(\m_sys.m_core.m_gpr._GEN[242] ));
 sg13g2_a221oi_1 _12746_ (.B2(\m_sys.m_core.m_gpr._GEN[210] ),
    .C1(net5182),
    .B1(net5057),
    .A1(\m_sys.m_core.m_gpr._GEN[146] ),
    .Y(_04182_),
    .A2(net5151));
 sg13g2_a22oi_1 _12747_ (.Y(_04183_),
    .B1(_04181_),
    .B2(_04182_),
    .A2(_04180_),
    .A1(_04179_));
 sg13g2_a21oi_1 _12748_ (.A1(net4385),
    .A2(_04183_),
    .Y(_04184_),
    .B1(net4727));
 sg13g2_a22oi_1 _12749_ (.Y(_00209_),
    .B1(_04178_),
    .B2(_04184_),
    .A2(net4727),
    .A1(net5177));
 sg13g2_nand2_1 _12750_ (.Y(_04185_),
    .A(net5168),
    .B(_03236_));
 sg13g2_a21oi_1 _12751_ (.A1(_03194_),
    .A2(_03238_),
    .Y(_04186_),
    .B1(_04185_));
 sg13g2_a221oi_1 _12752_ (.B2(_03239_),
    .C1(_04186_),
    .B1(_03961_),
    .A1(net5251),
    .Y(_04187_),
    .A2(_03370_));
 sg13g2_xnor2_1 _12753_ (.Y(_04188_),
    .A(_03245_),
    .B(_04187_));
 sg13g2_nor2_1 _12754_ (.A(net4775),
    .B(_03877_),
    .Y(_04189_));
 sg13g2_a21oi_1 _12755_ (.A1(net4779),
    .A2(_03884_),
    .Y(_04190_),
    .B1(_04189_));
 sg13g2_nand2_1 _12756_ (.Y(_04191_),
    .A(net4775),
    .B(_03875_));
 sg13g2_a221oi_1 _12757_ (.B2(net4769),
    .C1(_03607_),
    .B1(_04191_),
    .A1(net4765),
    .Y(_04192_),
    .A2(_04190_));
 sg13g2_o21ai_1 _12758_ (.B1(_04192_),
    .Y(_04193_),
    .A1(net5307),
    .A2(_04188_));
 sg13g2_and2_1 _12759_ (.A(_03461_),
    .B(_03465_),
    .X(_04194_));
 sg13g2_nor2_1 _12760_ (.A(net4930),
    .B(_04122_),
    .Y(_04195_));
 sg13g2_a21oi_2 _12761_ (.B1(_04195_),
    .Y(_04196_),
    .A2(_04194_),
    .A1(net4930));
 sg13g2_nor3_1 _12762_ (.A(net4771),
    .B(_04045_),
    .C(_04046_),
    .Y(_04197_));
 sg13g2_a21oi_2 _12763_ (.B1(_04197_),
    .Y(_04198_),
    .A2(_04196_),
    .A1(net4772));
 sg13g2_nand2b_1 _12764_ (.Y(_04199_),
    .B(net4784),
    .A_N(_04198_));
 sg13g2_o21ai_1 _12765_ (.B1(_04199_),
    .Y(_04200_),
    .A1(net4782),
    .A2(_03892_));
 sg13g2_and3_1 _12766_ (.X(_04201_),
    .A(net5250),
    .B(net4893),
    .C(_04200_));
 sg13g2_nand2b_1 _12767_ (.Y(_04202_),
    .B(net4956),
    .A_N(_03894_));
 sg13g2_a21oi_1 _12768_ (.A1(_04199_),
    .A2(_04202_),
    .Y(_04203_),
    .B1(net5253));
 sg13g2_nor3_1 _12769_ (.A(_03485_),
    .B(_04201_),
    .C(_04203_),
    .Y(_04204_));
 sg13g2_o21ai_1 _12770_ (.B1(net5174),
    .Y(_04205_),
    .A1(net5307),
    .A2(_03245_));
 sg13g2_nor2_1 _12771_ (.A(net5307),
    .B(_03244_),
    .Y(_04206_));
 sg13g2_nor3_1 _12772_ (.A(net5173),
    .B(_03241_),
    .C(_04206_),
    .Y(_04207_));
 sg13g2_nor2_1 _12773_ (.A(net5160),
    .B(_04207_),
    .Y(_04208_));
 sg13g2_o21ai_1 _12774_ (.B1(_04208_),
    .Y(_04209_),
    .A1(_04204_),
    .A2(_04205_));
 sg13g2_and2_1 _12775_ (.A(_04193_),
    .B(_04209_),
    .X(_04210_));
 sg13g2_mux2_1 _12776_ (.A0(\m_sys._m_ram_io_b_port_rdata[17] ),
    .A1(\m_sys._m_ram_io_b_port_rdata[25] ),
    .S(net5364),
    .X(_04211_));
 sg13g2_and2_1 _12777_ (.A(\m_sys._m_ram_io_b_port_rdata[17] ),
    .B(net5070),
    .X(_04212_));
 sg13g2_a22oi_1 _12778_ (.Y(_04213_),
    .B1(_04212_),
    .B2(net4495),
    .A2(_04211_),
    .A1(net4740));
 sg13g2_or2_2 _12779_ (.X(_04214_),
    .B(_04213_),
    .A(net4746));
 sg13g2_a221oi_1 _12780_ (.B2(net4038),
    .C1(net4751),
    .B1(_04214_),
    .A1(net5099),
    .Y(_04215_),
    .A2(_04210_));
 sg13g2_nand2_1 _12781_ (.Y(_04216_),
    .A(\m_sys.m_core.m_gpr._GEN[113] ),
    .B(net5063));
 sg13g2_a221oi_1 _12782_ (.B2(net5056),
    .C1(net5331),
    .B1(\m_sys.m_core.m_gpr._GEN[81] ),
    .A1(net5188),
    .Y(_04217_),
    .A2(\m_sys.m_core.m_gpr._GEN[49] ));
 sg13g2_a22oi_1 _12783_ (.Y(_04218_),
    .B1(net5049),
    .B2(\m_sys.m_core.m_gpr._GEN[177] ),
    .A2(net5063),
    .A1(\m_sys.m_core.m_gpr._GEN[241] ));
 sg13g2_a221oi_1 _12784_ (.B2(\m_sys.m_core.m_gpr._GEN[209] ),
    .C1(net5182),
    .B1(net5056),
    .A1(\m_sys.m_core.m_gpr._GEN[145] ),
    .Y(_04219_),
    .A2(net5152));
 sg13g2_a221oi_1 _12785_ (.B2(_04219_),
    .C1(_03560_),
    .B1(_04218_),
    .A1(_04216_),
    .Y(_04220_),
    .A2(_04217_));
 sg13g2_nor3_1 _12786_ (.A(net4725),
    .B(_04215_),
    .C(_04220_),
    .Y(_04221_));
 sg13g2_a21oi_1 _12787_ (.A1(net5178),
    .A2(net4725),
    .Y(_00210_),
    .B1(_04221_));
 sg13g2_o21ai_1 _12788_ (.B1(_03960_),
    .Y(_04222_),
    .A1(net5250),
    .A2(_03194_));
 sg13g2_xnor2_1 _12789_ (.Y(_04223_),
    .A(_03239_),
    .B(_04222_));
 sg13g2_a21oi_1 _12790_ (.A1(net4779),
    .A2(_03927_),
    .Y(_04224_),
    .B1(net4762));
 sg13g2_o21ai_1 _12791_ (.B1(_04224_),
    .Y(_04225_),
    .A1(net4779),
    .A2(_03920_));
 sg13g2_and2_1 _12792_ (.A(net4775),
    .B(_03922_),
    .X(_04226_));
 sg13g2_o21ai_1 _12793_ (.B1(_03606_),
    .Y(_04227_),
    .A1(net4767),
    .A2(_04226_));
 sg13g2_a21oi_1 _12794_ (.A1(net5166),
    .A2(_04223_),
    .Y(_04228_),
    .B1(_04227_));
 sg13g2_and2_1 _12795_ (.A(net4890),
    .B(_04083_),
    .X(_04229_));
 sg13g2_nand2_1 _12796_ (.Y(_04230_),
    .A(_03631_),
    .B(_03634_));
 sg13g2_a21oi_1 _12797_ (.A1(_03625_),
    .A2(_03632_),
    .Y(_04231_),
    .B1(net4930));
 sg13g2_a21o_1 _12798_ (.A2(_04230_),
    .A1(net4933),
    .B1(_04231_),
    .X(_04232_));
 sg13g2_a21oi_2 _12799_ (.B1(_04229_),
    .Y(_04233_),
    .A2(_04232_),
    .A1(net4772));
 sg13g2_nor2_1 _12800_ (.A(net4784),
    .B(_03933_),
    .Y(_04234_));
 sg13g2_a21oi_2 _12801_ (.B1(_04234_),
    .Y(_04235_),
    .A2(_04233_),
    .A1(net4784));
 sg13g2_a21oi_2 _12802_ (.B1(net4767),
    .Y(_04236_),
    .A2(net4884),
    .A1(net5253));
 sg13g2_a221oi_1 _12803_ (.B2(_04235_),
    .C1(_04236_),
    .B1(net4765),
    .A1(net5165),
    .Y(_04237_),
    .A2(_03239_));
 sg13g2_nand2_1 _12804_ (.Y(_04238_),
    .A(net5165),
    .B(_03238_));
 sg13g2_nand3_1 _12805_ (.B(_03236_),
    .C(_04238_),
    .A(net5291),
    .Y(_04239_));
 sg13g2_o21ai_1 _12806_ (.B1(_04239_),
    .Y(_04240_),
    .A1(net5291),
    .A2(_04237_));
 sg13g2_inv_1 _12807_ (.Y(_04241_),
    .A(_04240_));
 sg13g2_a22oi_1 _12808_ (.Y(_04242_),
    .B1(_04241_),
    .B2(net5258),
    .A2(_04228_),
    .A1(_04225_));
 sg13g2_nand2_1 _12809_ (.Y(_04243_),
    .A(net5100),
    .B(_04242_));
 sg13g2_mux2_1 _12810_ (.A0(\m_sys._m_ram_io_b_port_rdata[16] ),
    .A1(\m_sys._m_ram_io_b_port_rdata[24] ),
    .S(net5366),
    .X(_04244_));
 sg13g2_and2_1 _12811_ (.A(\m_sys._m_ram_io_b_port_rdata[16] ),
    .B(net5071),
    .X(_04245_));
 sg13g2_a22oi_1 _12812_ (.Y(_04246_),
    .B1(_04245_),
    .B2(net4497),
    .A2(_04244_),
    .A1(net4740));
 sg13g2_o21ai_1 _12813_ (.B1(net4040),
    .Y(_04247_),
    .A1(net4747),
    .A2(_04246_));
 sg13g2_nand3_1 _12814_ (.B(_04243_),
    .C(_04247_),
    .A(net4759),
    .Y(_04248_));
 sg13g2_nand2_1 _12815_ (.Y(_04249_),
    .A(\m_sys.m_core.m_gpr._GEN[112] ),
    .B(net5067));
 sg13g2_a221oi_1 _12816_ (.B2(net5056),
    .C1(net5331),
    .B1(\m_sys.m_core.m_gpr._GEN[80] ),
    .A1(net5187),
    .Y(_04250_),
    .A2(\m_sys.m_core.m_gpr._GEN[48] ));
 sg13g2_a22oi_1 _12817_ (.Y(_04251_),
    .B1(net5047),
    .B2(\m_sys.m_core.m_gpr._GEN[176] ),
    .A2(net5067),
    .A1(\m_sys.m_core.m_gpr._GEN[240] ));
 sg13g2_a221oi_1 _12818_ (.B2(\m_sys.m_core.m_gpr._GEN[208] ),
    .C1(net5182),
    .B1(net5056),
    .A1(\m_sys.m_core.m_gpr._GEN[144] ),
    .Y(_04252_),
    .A2(net5152));
 sg13g2_a22oi_1 _12819_ (.Y(_04253_),
    .B1(_04251_),
    .B2(_04252_),
    .A2(_04250_),
    .A1(_04249_));
 sg13g2_a21oi_1 _12820_ (.A1(net4385),
    .A2(_04253_),
    .Y(_04254_),
    .B1(net4727));
 sg13g2_a22oi_1 _12821_ (.Y(_00211_),
    .B1(_04248_),
    .B2(_04254_),
    .A2(net4727),
    .A1(net5185));
 sg13g2_o21ai_1 _12822_ (.B1(_03103_),
    .Y(_04255_),
    .A1(_03104_),
    .A2(_03184_));
 sg13g2_nor3_2 _12823_ (.A(_03104_),
    .B(_03109_),
    .C(_03184_),
    .Y(_04256_));
 sg13g2_o21ai_1 _12824_ (.B1(_03098_),
    .Y(_04257_),
    .A1(_03189_),
    .A2(_04256_));
 sg13g2_a22oi_1 _12825_ (.Y(_04258_),
    .B1(_03185_),
    .B2(_04257_),
    .A2(_03082_),
    .A1(_03080_));
 sg13g2_nand2_1 _12826_ (.Y(_04259_),
    .A(net5169),
    .B(_03081_));
 sg13g2_nand2_1 _12827_ (.Y(_04260_),
    .A(net5243),
    .B(_03359_));
 sg13g2_nand2_1 _12828_ (.Y(_04261_),
    .A(_03176_),
    .B(_03333_));
 sg13g2_nand3_1 _12829_ (.B(_03333_),
    .C(_03348_),
    .A(_03176_),
    .Y(_04262_));
 sg13g2_and2_1 _12830_ (.A(_03355_),
    .B(_04262_),
    .X(_04263_));
 sg13g2_a21oi_1 _12831_ (.A1(_03355_),
    .A2(_04262_),
    .Y(_04264_),
    .B1(_03344_));
 sg13g2_nor2_1 _12832_ (.A(_03351_),
    .B(_04264_),
    .Y(_04265_));
 sg13g2_nor2_1 _12833_ (.A(net5169),
    .B(_04265_),
    .Y(_04266_));
 sg13g2_o21ai_1 _12834_ (.B1(net5243),
    .Y(_04267_),
    .A1(_03351_),
    .A2(_04264_));
 sg13g2_o21ai_1 _12835_ (.B1(_04260_),
    .Y(_04268_),
    .A1(_03334_),
    .A2(_04267_));
 sg13g2_a22oi_1 _12836_ (.Y(_04269_),
    .B1(_04268_),
    .B2(_03085_),
    .A2(_03360_),
    .A1(net5243));
 sg13g2_o21ai_1 _12837_ (.B1(_04269_),
    .Y(_04270_),
    .A1(_04258_),
    .A2(_04259_));
 sg13g2_xnor2_1 _12838_ (.Y(_04271_),
    .A(_03078_),
    .B(_04270_));
 sg13g2_a21oi_1 _12839_ (.A1(net5307),
    .A2(_03440_),
    .Y(_04272_),
    .B1(_04003_));
 sg13g2_o21ai_1 _12840_ (.B1(_04272_),
    .Y(_04273_),
    .A1(net5306),
    .A2(_04271_));
 sg13g2_nand2_1 _12841_ (.Y(_04274_),
    .A(_03412_),
    .B(_03464_));
 sg13g2_nor2_1 _12842_ (.A(net4917),
    .B(_04274_),
    .Y(_04275_));
 sg13g2_a21oi_2 _12843_ (.B1(_04275_),
    .Y(_04276_),
    .A2(_04194_),
    .A1(net4921));
 sg13g2_mux2_1 _12844_ (.A0(_04123_),
    .A1(_04276_),
    .S(net4771),
    .X(_04277_));
 sg13g2_nor2_1 _12845_ (.A(net4955),
    .B(_04277_),
    .Y(_04278_));
 sg13g2_a21oi_1 _12846_ (.A1(net4953),
    .A2(_03975_),
    .Y(_04279_),
    .B1(_04278_));
 sg13g2_nor2_1 _12847_ (.A(net5306),
    .B(_03078_),
    .Y(_04280_));
 sg13g2_a221oi_1 _12848_ (.B2(net4766),
    .C1(_04280_),
    .B1(_04279_),
    .A1(_03489_),
    .Y(_04281_),
    .A2(_04236_));
 sg13g2_nor2_1 _12849_ (.A(net5172),
    .B(_03074_),
    .Y(_04282_));
 sg13g2_o21ai_1 _12850_ (.B1(_04282_),
    .Y(_04283_),
    .A1(net5306),
    .A2(_03077_));
 sg13g2_o21ai_1 _12851_ (.B1(_04283_),
    .Y(_04284_),
    .A1(net5287),
    .A2(_04281_));
 sg13g2_o21ai_1 _12852_ (.B1(_04273_),
    .Y(_04285_),
    .A1(net5160),
    .A2(_04284_));
 sg13g2_or2_1 _12853_ (.X(_04286_),
    .B(\m_sys.m_core.r_ctrl_mem_size[0] ),
    .A(\m_sys.m_core.r_ctrl_mem_size[1] ));
 sg13g2_nor2_1 _12854_ (.A(_03538_),
    .B(_04286_),
    .Y(_04287_));
 sg13g2_a21oi_2 _12855_ (.B1(net5101),
    .Y(_04288_),
    .A2(_04287_),
    .A1(_03520_));
 sg13g2_a21oi_2 _12856_ (.B1(_03538_),
    .Y(_04289_),
    .A2(_04286_),
    .A1(_03548_));
 sg13g2_nor2b_1 _12857_ (.A(_03522_),
    .B_N(net4747),
    .Y(_04290_));
 sg13g2_nand2b_1 _12858_ (.Y(_04291_),
    .B(_03536_),
    .A_N(_04290_));
 sg13g2_a21oi_2 _12859_ (.B1(net4748),
    .Y(_04292_),
    .A2(_04291_),
    .A1(_04288_));
 sg13g2_o21ai_1 _12860_ (.B1(_04292_),
    .Y(_04293_),
    .A1(net5098),
    .A2(_04285_));
 sg13g2_nand2_1 _12861_ (.Y(_04294_),
    .A(\m_sys.m_core.m_gpr._GEN[111] ),
    .B(net5067));
 sg13g2_a221oi_1 _12862_ (.B2(\m_sys.m_core.m_gpr._GEN[79] ),
    .C1(net5330),
    .B1(net5056),
    .A1(\m_sys.m_core.m_gpr._GEN[47] ),
    .Y(_04295_),
    .A2(net5188));
 sg13g2_a22oi_1 _12863_ (.Y(_04296_),
    .B1(net5047),
    .B2(\m_sys.m_core.m_gpr._GEN[175] ),
    .A2(net5067),
    .A1(\m_sys.m_core.m_gpr._GEN[239] ));
 sg13g2_a221oi_1 _12864_ (.B2(\m_sys.m_core.m_gpr._GEN[207] ),
    .C1(net5182),
    .B1(net5058),
    .A1(\m_sys.m_core.m_gpr._GEN[143] ),
    .Y(_04297_),
    .A2(net5150));
 sg13g2_a22oi_1 _12865_ (.Y(_04298_),
    .B1(_04296_),
    .B2(_04297_),
    .A2(_04295_),
    .A1(_04294_));
 sg13g2_a21oi_1 _12866_ (.A1(net4385),
    .A2(_04298_),
    .Y(_04299_),
    .B1(net4727));
 sg13g2_a22oi_1 _12867_ (.Y(_00212_),
    .B1(_04293_),
    .B2(_04299_),
    .A2(net4727),
    .A1(net5191));
 sg13g2_nand3_1 _12868_ (.B(_03185_),
    .C(_04257_),
    .A(net5169),
    .Y(_04300_));
 sg13g2_nand2b_1 _12869_ (.Y(_04301_),
    .B(_04300_),
    .A_N(_04268_));
 sg13g2_xnor2_1 _12870_ (.Y(_04302_),
    .A(_03084_),
    .B(_04301_));
 sg13g2_a21oi_1 _12871_ (.A1(net5300),
    .A2(_03605_),
    .Y(_04303_),
    .B1(net4717));
 sg13g2_o21ai_1 _12872_ (.B1(_04303_),
    .Y(_04304_),
    .A1(net5293),
    .A2(_04302_));
 sg13g2_nand2_1 _12873_ (.Y(_04305_),
    .A(net5247),
    .B(_03650_));
 sg13g2_nor2_1 _12874_ (.A(net4767),
    .B(_03652_),
    .Y(_04306_));
 sg13g2_a21oi_1 _12875_ (.A1(_03597_),
    .A2(_03633_),
    .Y(_04307_),
    .B1(net4917));
 sg13g2_a21o_1 _12876_ (.A2(_04230_),
    .A1(net4916),
    .B1(_04307_),
    .X(_04308_));
 sg13g2_mux2_2 _12877_ (.A0(_04158_),
    .A1(_04308_),
    .S(net4773),
    .X(_04309_));
 sg13g2_o21ai_1 _12878_ (.B1(net4766),
    .Y(_04310_),
    .A1(net4950),
    .A2(_04309_));
 sg13g2_a21oi_1 _12879_ (.A1(net4953),
    .A2(_04008_),
    .Y(_04311_),
    .B1(_04310_));
 sg13g2_a221oi_1 _12880_ (.B2(_04306_),
    .C1(_04311_),
    .B1(_04305_),
    .A1(net5163),
    .Y(_04312_),
    .A2(_03085_));
 sg13g2_nor2_1 _12881_ (.A(net5287),
    .B(_04312_),
    .Y(_04313_));
 sg13g2_a21oi_1 _12882_ (.A1(_03080_),
    .A2(_03082_),
    .Y(_04314_),
    .B1(net5294));
 sg13g2_nand2_1 _12883_ (.Y(_04315_),
    .A(net5287),
    .B(_03081_));
 sg13g2_o21ai_1 _12884_ (.B1(net5256),
    .Y(_04316_),
    .A1(_04314_),
    .A2(_04315_));
 sg13g2_o21ai_1 _12885_ (.B1(_04304_),
    .Y(_04317_),
    .A1(_04313_),
    .A2(_04316_));
 sg13g2_nand2b_1 _12886_ (.Y(_04318_),
    .B(net4387),
    .A_N(_00141_));
 sg13g2_o21ai_1 _12887_ (.B1(_04318_),
    .Y(_04319_),
    .A1(_00061_),
    .A2(_02698_));
 sg13g2_mux2_1 _12888_ (.A0(_00061_),
    .A1(_00142_),
    .S(net5360),
    .X(_04320_));
 sg13g2_a21oi_1 _12889_ (.A1(net5356),
    .A2(_03660_),
    .Y(_04321_),
    .B1(net5072));
 sg13g2_o21ai_1 _12890_ (.B1(_04321_),
    .Y(_04322_),
    .A1(net5356),
    .A2(_04320_));
 sg13g2_nand2_1 _12891_ (.Y(_04323_),
    .A(net5073),
    .B(net4881));
 sg13g2_nand2_1 _12892_ (.Y(_04324_),
    .A(net5277),
    .B(_04323_));
 sg13g2_a21oi_1 _12893_ (.A1(_00141_),
    .A2(net5073),
    .Y(_04325_),
    .B1(_04324_));
 sg13g2_a22oi_1 _12894_ (.Y(_04326_),
    .B1(_04322_),
    .B2(_04325_),
    .A2(_04319_),
    .A1(net5069));
 sg13g2_o21ai_1 _12895_ (.B1(_04288_),
    .Y(_04327_),
    .A1(_04290_),
    .A2(_04326_));
 sg13g2_and2_1 _12896_ (.A(net4755),
    .B(_04327_),
    .X(_04328_));
 sg13g2_o21ai_1 _12897_ (.B1(_04328_),
    .Y(_04329_),
    .A1(net5098),
    .A2(_04317_));
 sg13g2_nand2_1 _12898_ (.Y(_04330_),
    .A(\m_sys.m_core.m_gpr._GEN[110] ),
    .B(net5067));
 sg13g2_a221oi_1 _12899_ (.B2(\m_sys.m_core.m_gpr._GEN[78] ),
    .C1(net5331),
    .B1(net5056),
    .A1(\m_sys.m_core.m_gpr._GEN[46] ),
    .Y(_04331_),
    .A2(net5188));
 sg13g2_a22oi_1 _12900_ (.Y(_04332_),
    .B1(net5047),
    .B2(\m_sys.m_core.m_gpr._GEN[174] ),
    .A2(net5067),
    .A1(\m_sys.m_core.m_gpr._GEN[238] ));
 sg13g2_a221oi_1 _12901_ (.B2(\m_sys.m_core.m_gpr._GEN[206] ),
    .C1(net5181),
    .B1(net5054),
    .A1(\m_sys.m_core.m_gpr._GEN[142] ),
    .Y(_04333_),
    .A2(net5150));
 sg13g2_a22oi_1 _12902_ (.Y(_04334_),
    .B1(_04332_),
    .B2(_04333_),
    .A2(_04331_),
    .A1(_04330_));
 sg13g2_a21oi_1 _12903_ (.A1(net4386),
    .A2(_04334_),
    .Y(_04335_),
    .B1(net4723));
 sg13g2_a22oi_1 _12904_ (.Y(_00213_),
    .B1(_04329_),
    .B2(_04335_),
    .A2(net4722),
    .A1(net5222));
 sg13g2_o21ai_1 _12905_ (.B1(_03096_),
    .Y(_04336_),
    .A1(_03189_),
    .A2(_04256_));
 sg13g2_nor2_1 _12906_ (.A(net5243),
    .B(_03094_),
    .Y(_04337_));
 sg13g2_o21ai_1 _12907_ (.B1(_03357_),
    .Y(_04338_),
    .A1(_03097_),
    .A2(_04265_));
 sg13g2_a22oi_1 _12908_ (.Y(_04339_),
    .B1(_04338_),
    .B2(net5243),
    .A2(_04337_),
    .A1(_04336_));
 sg13g2_xor2_1 _12909_ (.B(_04339_),
    .A(_03091_),
    .X(_04340_));
 sg13g2_or2_1 _12910_ (.X(_04341_),
    .B(_04340_),
    .A(net5294));
 sg13g2_a21oi_1 _12911_ (.A1(net5300),
    .A2(_03688_),
    .Y(_04342_),
    .B1(net4717));
 sg13g2_a21oi_1 _12912_ (.A1(net5249),
    .A2(_03704_),
    .Y(_04343_),
    .B1(net4767));
 sg13g2_nor2_1 _12913_ (.A(net5294),
    .B(_03091_),
    .Y(_04344_));
 sg13g2_nand2_1 _12914_ (.Y(_04345_),
    .A(net4953),
    .B(_04049_));
 sg13g2_a21oi_1 _12915_ (.A1(_03411_),
    .A2(_03415_),
    .Y(_04346_),
    .B1(net4916));
 sg13g2_a21o_1 _12916_ (.A2(_04274_),
    .A1(net4916),
    .B1(_04346_),
    .X(_04347_));
 sg13g2_or2_1 _12917_ (.X(_04348_),
    .B(_04347_),
    .A(net4891));
 sg13g2_o21ai_1 _12918_ (.B1(_04348_),
    .Y(_04349_),
    .A1(net4773),
    .A2(_04196_));
 sg13g2_a21oi_1 _12919_ (.A1(net4780),
    .A2(_04349_),
    .Y(_04350_),
    .B1(net4761));
 sg13g2_a221oi_1 _12920_ (.B2(_04350_),
    .C1(_04344_),
    .B1(_04345_),
    .A1(_03708_),
    .Y(_04351_),
    .A2(_04343_));
 sg13g2_nor2_1 _12921_ (.A(net5287),
    .B(_04351_),
    .Y(_04352_));
 sg13g2_a221oi_1 _12922_ (.B2(net5162),
    .C1(net5172),
    .B1(_03090_),
    .A1(\m_sys.m_core.m_bru.io_i_s2[13] ),
    .Y(_04353_),
    .A2(_03087_));
 sg13g2_nor2_1 _12923_ (.A(_04352_),
    .B(_04353_),
    .Y(_04354_));
 sg13g2_a22oi_1 _12924_ (.Y(_04355_),
    .B1(_04354_),
    .B2(net5256),
    .A2(_04342_),
    .A1(_04341_));
 sg13g2_nor2b_1 _12925_ (.A(net5364),
    .B_N(_00059_),
    .Y(_04356_));
 sg13g2_a21oi_1 _12926_ (.A1(net5364),
    .A2(_00140_),
    .Y(_04357_),
    .B1(_04356_));
 sg13g2_o21ai_1 _12927_ (.B1(net4883),
    .Y(_04358_),
    .A1(net5358),
    .A2(_04357_));
 sg13g2_a21oi_1 _12928_ (.A1(net5357),
    .A2(_03716_),
    .Y(_04359_),
    .B1(_04358_));
 sg13g2_o21ai_1 _12929_ (.B1(net5279),
    .Y(_04360_),
    .A1(_03514_),
    .A2(_04359_));
 sg13g2_o21ai_1 _12930_ (.B1(_04360_),
    .Y(_04361_),
    .A1(_00059_),
    .A2(_02698_));
 sg13g2_a21oi_1 _12931_ (.A1(_02502_),
    .A2(net4387),
    .Y(_04362_),
    .B1(_04361_));
 sg13g2_o21ai_1 _12932_ (.B1(_03532_),
    .Y(_04363_),
    .A1(_00139_),
    .A2(_03513_));
 sg13g2_nor2_1 _12933_ (.A(_04359_),
    .B(_04363_),
    .Y(_04364_));
 sg13g2_or3_1 _12934_ (.A(_04290_),
    .B(_04362_),
    .C(_04364_),
    .X(_04365_));
 sg13g2_a221oi_1 _12935_ (.B2(_04288_),
    .C1(net4748),
    .B1(_04365_),
    .A1(net5101),
    .Y(_04366_),
    .A2(_04355_));
 sg13g2_nand2_1 _12936_ (.Y(_04367_),
    .A(\m_sys.m_core.m_gpr._GEN[109] ),
    .B(net5065));
 sg13g2_a221oi_1 _12937_ (.B2(\m_sys.m_core.m_gpr._GEN[77] ),
    .C1(net5329),
    .B1(net5055),
    .A1(\m_sys.m_core.m_gpr._GEN[45] ),
    .Y(_04368_),
    .A2(net5186));
 sg13g2_a22oi_1 _12938_ (.Y(_04369_),
    .B1(net5048),
    .B2(\m_sys.m_core.m_gpr._GEN[173] ),
    .A2(net5065),
    .A1(\m_sys.m_core.m_gpr._GEN[237] ));
 sg13g2_a221oi_1 _12939_ (.B2(\m_sys.m_core.m_gpr._GEN[205] ),
    .C1(net5181),
    .B1(net5055),
    .A1(\m_sys.m_core.m_gpr._GEN[141] ),
    .Y(_04370_),
    .A2(net5151));
 sg13g2_a221oi_1 _12940_ (.B2(_04370_),
    .C1(_03560_),
    .B1(_04369_),
    .A1(_04367_),
    .Y(_04371_),
    .A2(_04368_));
 sg13g2_nor3_1 _12941_ (.A(net4722),
    .B(_04366_),
    .C(_04371_),
    .Y(_04372_));
 sg13g2_a21oi_1 _12942_ (.A1(net5224),
    .A2(net4722),
    .Y(_00214_),
    .B1(_04372_));
 sg13g2_nor3_1 _12943_ (.A(net5243),
    .B(_03189_),
    .C(_04256_),
    .Y(_04373_));
 sg13g2_nor2_1 _12944_ (.A(_04266_),
    .B(_04373_),
    .Y(_04374_));
 sg13g2_xnor2_1 _12945_ (.Y(_04375_),
    .A(_03097_),
    .B(_04374_));
 sg13g2_nand2_1 _12946_ (.Y(_04376_),
    .A(net5162),
    .B(_04375_));
 sg13g2_a21oi_1 _12947_ (.A1(net5298),
    .A2(_03741_),
    .Y(_04377_),
    .B1(net4717));
 sg13g2_o21ai_1 _12948_ (.B1(net5303),
    .Y(_04378_),
    .A1(_03488_),
    .A2(_03762_));
 sg13g2_a21oi_1 _12949_ (.A1(net5249),
    .A2(_03760_),
    .Y(_04379_),
    .B1(_04378_));
 sg13g2_nand2_1 _12950_ (.Y(_04380_),
    .A(_03596_),
    .B(_03600_));
 sg13g2_a21oi_1 _12951_ (.A1(_03597_),
    .A2(_03633_),
    .Y(_04381_),
    .B1(net4933));
 sg13g2_a21o_1 _12952_ (.A2(_04380_),
    .A1(net4933),
    .B1(_04381_),
    .X(_04382_));
 sg13g2_and2_1 _12953_ (.A(net4773),
    .B(_04382_),
    .X(_04383_));
 sg13g2_a21oi_2 _12954_ (.B1(_04383_),
    .Y(_04384_),
    .A2(_04232_),
    .A1(net4890));
 sg13g2_a21oi_1 _12955_ (.A1(net4954),
    .A2(_04085_),
    .Y(_04385_),
    .B1(_03151_));
 sg13g2_o21ai_1 _12956_ (.B1(_04385_),
    .Y(_04386_),
    .A1(net4954),
    .A2(_04384_));
 sg13g2_o21ai_1 _12957_ (.B1(_04386_),
    .Y(_04387_),
    .A1(net4766),
    .A2(_04379_));
 sg13g2_o21ai_1 _12958_ (.B1(_04387_),
    .Y(_04388_),
    .A1(net5293),
    .A2(_03097_));
 sg13g2_a221oi_1 _12959_ (.B2(net5162),
    .C1(net5172),
    .B1(_03096_),
    .A1(\m_sys.m_core.m_bru.io_i_s2[12] ),
    .Y(_04389_),
    .A2(_03092_));
 sg13g2_a21oi_1 _12960_ (.A1(net5172),
    .A2(_04388_),
    .Y(_04390_),
    .B1(_04389_));
 sg13g2_a22oi_1 _12961_ (.Y(_04391_),
    .B1(_04390_),
    .B2(net5256),
    .A2(_04377_),
    .A1(_04376_));
 sg13g2_nand2_1 _12962_ (.Y(_04392_),
    .A(net5099),
    .B(_04391_));
 sg13g2_nor2b_1 _12963_ (.A(net5363),
    .B_N(_00057_),
    .Y(_04393_));
 sg13g2_a21oi_1 _12964_ (.A1(net5363),
    .A2(_00138_),
    .Y(_04394_),
    .B1(_04393_));
 sg13g2_o21ai_1 _12965_ (.B1(net4883),
    .Y(_04395_),
    .A1(net5358),
    .A2(_04394_));
 sg13g2_a21oi_1 _12966_ (.A1(net5357),
    .A2(_03770_),
    .Y(_04396_),
    .B1(_04395_));
 sg13g2_o21ai_1 _12967_ (.B1(net4879),
    .Y(_04397_),
    .A1(_00137_),
    .A2(_03513_));
 sg13g2_or2_1 _12968_ (.X(_04398_),
    .B(_04397_),
    .A(_04396_));
 sg13g2_nor3_1 _12969_ (.A(_00137_),
    .B(net4493),
    .C(_03498_),
    .Y(_04399_));
 sg13g2_o21ai_1 _12970_ (.B1(net5278),
    .Y(_04400_),
    .A1(_03514_),
    .A2(_04396_));
 sg13g2_o21ai_1 _12971_ (.B1(_04400_),
    .Y(_04401_),
    .A1(_00057_),
    .A2(_02698_));
 sg13g2_o21ai_1 _12972_ (.B1(_04398_),
    .Y(_04402_),
    .A1(_04399_),
    .A2(_04401_));
 sg13g2_o21ai_1 _12973_ (.B1(_04288_),
    .Y(_04403_),
    .A1(_04290_),
    .A2(_04402_));
 sg13g2_nand3_1 _12974_ (.B(_04392_),
    .C(_04403_),
    .A(net4756),
    .Y(_04404_));
 sg13g2_nand2_1 _12975_ (.Y(_04405_),
    .A(\m_sys.m_core.m_gpr._GEN[108] ),
    .B(net5063));
 sg13g2_a221oi_1 _12976_ (.B2(\m_sys.m_core.m_gpr._GEN[76] ),
    .C1(net5329),
    .B1(net5054),
    .A1(\m_sys.m_core.m_gpr._GEN[44] ),
    .Y(_04406_),
    .A2(net5186));
 sg13g2_a22oi_1 _12977_ (.Y(_04407_),
    .B1(net5048),
    .B2(\m_sys.m_core.m_gpr._GEN[172] ),
    .A2(net5063),
    .A1(\m_sys.m_core.m_gpr._GEN[236] ));
 sg13g2_a221oi_1 _12978_ (.B2(\m_sys.m_core.m_gpr._GEN[204] ),
    .C1(net5180),
    .B1(net5054),
    .A1(\m_sys.m_core.m_gpr._GEN[140] ),
    .Y(_04408_),
    .A2(net5150));
 sg13g2_a22oi_1 _12979_ (.Y(_04409_),
    .B1(_04407_),
    .B2(_04408_),
    .A2(_04406_),
    .A1(_04405_));
 sg13g2_a21oi_1 _12980_ (.A1(net4386),
    .A2(_04409_),
    .Y(_04410_),
    .B1(net4722));
 sg13g2_a22oi_1 _12981_ (.Y(_00215_),
    .B1(_04404_),
    .B2(_04410_),
    .A2(net4722),
    .A1(net5223));
 sg13g2_nand2_1 _12982_ (.Y(_04411_),
    .A(\m_sys.m_core.m_bru.io_i_pc[3] ),
    .B(\m_sys.m_core.m_bru.io_i_pc[2] ));
 sg13g2_nand4_1 _12983_ (.B(\m_sys.m_core.m_bru.io_i_pc[4] ),
    .C(\m_sys.m_core.m_bru.io_i_pc[3] ),
    .A(\m_sys.m_core.m_bru.io_i_pc[5] ),
    .Y(_04412_),
    .D(\m_sys.m_core.m_bru.io_i_pc[2] ));
 sg13g2_nand2_1 _12984_ (.Y(_04413_),
    .A(\m_sys.m_core.m_bru.io_i_pc[7] ),
    .B(\m_sys.m_core.m_bru.io_i_pc[6] ));
 sg13g2_nor2_1 _12985_ (.A(_04412_),
    .B(_04413_),
    .Y(_04414_));
 sg13g2_nand3_1 _12986_ (.B(\m_sys.m_core.m_bru.io_i_pc[8] ),
    .C(_04414_),
    .A(\m_sys.m_core.m_bru.io_i_pc[9] ),
    .Y(_04415_));
 sg13g2_nor2_1 _12987_ (.A(_00103_),
    .B(_04415_),
    .Y(_04416_));
 sg13g2_xnor2_1 _12988_ (.Y(_04417_),
    .A(net3083),
    .B(_04416_));
 sg13g2_nor2_1 _12989_ (.A(net5093),
    .B(_04417_),
    .Y(_04418_));
 sg13g2_nor3_2 _12990_ (.A(net4768),
    .B(_03809_),
    .C(_03812_),
    .Y(_04419_));
 sg13g2_nand2_1 _12991_ (.Y(_04420_),
    .A(net4891),
    .B(_04276_));
 sg13g2_o21ai_1 _12992_ (.B1(_03414_),
    .Y(_04421_),
    .A1(_03106_),
    .A2(net4899));
 sg13g2_nand3_1 _12993_ (.B(_03411_),
    .C(_03415_),
    .A(net4916),
    .Y(_04422_));
 sg13g2_o21ai_1 _12994_ (.B1(_04422_),
    .Y(_04423_),
    .A1(net4915),
    .A2(_04421_));
 sg13g2_o21ai_1 _12995_ (.B1(_04420_),
    .Y(_04424_),
    .A1(net4891),
    .A2(_04423_));
 sg13g2_a21o_1 _12996_ (.A2(_04125_),
    .A1(net4955),
    .B1(net4763),
    .X(_04425_));
 sg13g2_a21oi_1 _12997_ (.A1(net4776),
    .A2(_04424_),
    .Y(_04426_),
    .B1(_04425_));
 sg13g2_o21ai_1 _12998_ (.B1(net5172),
    .Y(_04427_),
    .A1(net5293),
    .A2(_03109_));
 sg13g2_or3_1 _12999_ (.A(_04419_),
    .B(_04426_),
    .C(_04427_),
    .X(_04428_));
 sg13g2_a21o_1 _13000_ (.A2(_03338_),
    .A1(_03105_),
    .B1(net5293),
    .X(_04429_));
 sg13g2_and2_1 _13001_ (.A(net5287),
    .B(_03107_),
    .X(_04430_));
 sg13g2_a21oi_1 _13002_ (.A1(_04429_),
    .A2(_04430_),
    .Y(_04431_),
    .B1(net5160));
 sg13g2_a21oi_1 _13003_ (.A1(_03109_),
    .A2(_04255_),
    .Y(_04432_),
    .B1(net5244));
 sg13g2_o21ai_1 _13004_ (.B1(_04432_),
    .Y(_04433_),
    .A1(_03109_),
    .A2(_04255_));
 sg13g2_o21ai_1 _13005_ (.B1(_03102_),
    .Y(_04434_),
    .A1(_03342_),
    .A2(_04263_));
 sg13g2_a21oi_1 _13006_ (.A1(_03339_),
    .A2(_04434_),
    .Y(_04435_),
    .B1(net5169));
 sg13g2_o21ai_1 _13007_ (.B1(_04435_),
    .Y(_04436_),
    .A1(_03339_),
    .A2(_04434_));
 sg13g2_a21o_1 _13008_ (.A2(_04436_),
    .A1(_04433_),
    .B1(net5293),
    .X(_04437_));
 sg13g2_a21oi_1 _13009_ (.A1(net5298),
    .A2(_03795_),
    .Y(_04438_),
    .B1(net4717));
 sg13g2_a22oi_1 _13010_ (.Y(_04439_),
    .B1(_04437_),
    .B2(_04438_),
    .A2(_04431_),
    .A1(_04428_));
 sg13g2_inv_1 _13011_ (.Y(_04440_),
    .A(_04439_));
 sg13g2_a22oi_1 _13012_ (.Y(_04441_),
    .B1(_03523_),
    .B2(\m_sys._m_uart_io_b_mem_rdata[11] ),
    .A2(net4497),
    .A1(\m_sys._m_ram_io_b_port_rdata[11] ));
 sg13g2_and2_1 _13013_ (.A(\m_sys._m_uart_io_b_mem_rdata[11] ),
    .B(net4882),
    .X(_04442_));
 sg13g2_mux2_1 _13014_ (.A0(\m_sys._m_ram_io_b_port_rdata[11] ),
    .A1(\m_sys._m_ram_io_b_port_rdata[19] ),
    .S(net5362),
    .X(_04443_));
 sg13g2_o21ai_1 _13015_ (.B1(net4883),
    .Y(_04444_),
    .A1(net5358),
    .A2(_04443_));
 sg13g2_a21oi_1 _13016_ (.A1(net5358),
    .A2(_03821_),
    .Y(_04445_),
    .B1(_04444_));
 sg13g2_o21ai_1 _13017_ (.B1(net5279),
    .Y(_04446_),
    .A1(_04442_),
    .A2(_04445_));
 sg13g2_o21ai_1 _13018_ (.B1(_04446_),
    .Y(_04447_),
    .A1(net4879),
    .A2(_04441_));
 sg13g2_nand2b_1 _13019_ (.Y(_04448_),
    .B(_04447_),
    .A_N(_04289_));
 sg13g2_a221oi_1 _13020_ (.B2(_04288_),
    .C1(net5094),
    .B1(_04448_),
    .A1(net5101),
    .Y(_04449_),
    .A2(_04439_));
 sg13g2_o21ai_1 _13021_ (.B1(net4958),
    .Y(_04450_),
    .A1(_04418_),
    .A2(_04449_));
 sg13g2_a22oi_1 _13022_ (.Y(_04451_),
    .B1(net5048),
    .B2(\m_sys.m_core.m_gpr._GEN[171] ),
    .A2(net5065),
    .A1(\m_sys.m_core.m_gpr._GEN[235] ));
 sg13g2_a221oi_1 _13023_ (.B2(\m_sys.m_core.m_gpr._GEN[203] ),
    .C1(net5181),
    .B1(net5055),
    .A1(\m_sys.m_core.m_gpr._GEN[139] ),
    .Y(_04452_),
    .A2(net5151));
 sg13g2_nand2_1 _13024_ (.Y(_04453_),
    .A(\m_sys.m_core.m_gpr._GEN[107] ),
    .B(net5065));
 sg13g2_a221oi_1 _13025_ (.B2(\m_sys.m_core.m_gpr._GEN[75] ),
    .C1(net5329),
    .B1(net5055),
    .A1(\m_sys.m_core.m_gpr._GEN[43] ),
    .Y(_04454_),
    .A2(net5186));
 sg13g2_a22oi_1 _13026_ (.Y(_04455_),
    .B1(_04453_),
    .B2(_04454_),
    .A2(_04452_),
    .A1(_04451_));
 sg13g2_nor2_2 _13027_ (.A(net5317),
    .B(_03552_),
    .Y(_04456_));
 sg13g2_nor3_2 _13028_ (.A(net5317),
    .B(net4960),
    .C(_03552_),
    .Y(_04457_));
 sg13g2_a221oi_1 _13029_ (.B2(net3083),
    .C1(net4721),
    .B1(_04457_),
    .A1(net4386),
    .Y(_04458_),
    .A2(_04455_));
 sg13g2_a22oi_1 _13030_ (.Y(_00216_),
    .B1(_04450_),
    .B2(_04458_),
    .A2(net4721),
    .A1(net5230));
 sg13g2_nor2_1 _13031_ (.A(net5298),
    .B(_03104_),
    .Y(_04459_));
 sg13g2_nand2_1 _13032_ (.Y(_04460_),
    .A(net4891),
    .B(_04308_));
 sg13g2_nand2_1 _13033_ (.Y(_04461_),
    .A(_03106_),
    .B(net4900));
 sg13g2_o21ai_1 _13034_ (.B1(_04461_),
    .Y(_04462_),
    .A1(_03100_),
    .A2(net4900));
 sg13g2_nand2_1 _13035_ (.Y(_04463_),
    .A(net4926),
    .B(_04462_));
 sg13g2_o21ai_1 _13036_ (.B1(_04463_),
    .Y(_04464_),
    .A1(net4926),
    .A2(_04380_));
 sg13g2_o21ai_1 _13037_ (.B1(_04460_),
    .Y(_04465_),
    .A1(net4891),
    .A2(_04464_));
 sg13g2_nand2_1 _13038_ (.Y(_04466_),
    .A(net4776),
    .B(_04465_));
 sg13g2_a21oi_1 _13039_ (.A1(net4953),
    .A2(_04160_),
    .Y(_04467_),
    .B1(net4761));
 sg13g2_a21oi_1 _13040_ (.A1(_04466_),
    .A2(_04467_),
    .Y(_04468_),
    .B1(_04459_));
 sg13g2_nor3_1 _13041_ (.A(net5287),
    .B(net4767),
    .C(_03851_),
    .Y(_04469_));
 sg13g2_a21oi_1 _13042_ (.A1(net5293),
    .A2(_03103_),
    .Y(_04470_),
    .B1(net5172));
 sg13g2_a22oi_1 _13043_ (.Y(_04471_),
    .B1(_04470_),
    .B2(_03341_),
    .A2(_04469_),
    .A1(_03853_));
 sg13g2_o21ai_1 _13044_ (.B1(_04471_),
    .Y(_04472_),
    .A1(net5287),
    .A2(_04468_));
 sg13g2_xor2_1 _13045_ (.B(_04263_),
    .A(_03342_),
    .X(_04473_));
 sg13g2_a21oi_1 _13046_ (.A1(_03104_),
    .A2(_03184_),
    .Y(_04474_),
    .B1(net5243));
 sg13g2_o21ai_1 _13047_ (.B1(_04474_),
    .Y(_04475_),
    .A1(_03104_),
    .A2(_03184_));
 sg13g2_a21oi_1 _13048_ (.A1(net5243),
    .A2(_04473_),
    .Y(_04476_),
    .B1(net5293));
 sg13g2_a221oi_1 _13049_ (.B2(_04476_),
    .C1(net4717),
    .B1(_04475_),
    .A1(net5293),
    .Y(_04477_),
    .A2(_03839_));
 sg13g2_a21o_2 _13050_ (.A2(_04472_),
    .A1(net5256),
    .B1(_04477_),
    .X(_04478_));
 sg13g2_a21o_1 _13051_ (.A2(_04478_),
    .A1(_02369_),
    .B1(net5097),
    .X(_04479_));
 sg13g2_a22oi_1 _13052_ (.Y(_04480_),
    .B1(_03523_),
    .B2(\m_sys._m_uart_io_b_mem_rdata[10] ),
    .A2(net4497),
    .A1(\m_sys._m_ram_io_b_port_rdata[10] ));
 sg13g2_inv_1 _13053_ (.Y(_04481_),
    .A(_04480_));
 sg13g2_nand2b_1 _13054_ (.Y(_04482_),
    .B(net5363),
    .A_N(\m_sys._m_ram_io_b_port_rdata[18] ));
 sg13g2_o21ai_1 _13055_ (.B1(_04482_),
    .Y(_04483_),
    .A1(\m_sys._m_ram_io_b_port_rdata[10] ),
    .A2(net5362));
 sg13g2_nand3b_1 _13056_ (.B(net5357),
    .C(\m_sys._m_ram_io_b_port_rdata[26] ),
    .Y(_04484_),
    .A_N(net5362));
 sg13g2_o21ai_1 _13057_ (.B1(_04484_),
    .Y(_04485_),
    .A1(net5357),
    .A2(_04483_));
 sg13g2_a22oi_1 _13058_ (.Y(_04486_),
    .B1(_04485_),
    .B2(net4883),
    .A2(net4882),
    .A1(\m_sys._m_uart_io_b_mem_rdata[10] ));
 sg13g2_inv_1 _13059_ (.Y(_04487_),
    .A(_04486_));
 sg13g2_a22oi_1 _13060_ (.Y(_04488_),
    .B1(_04487_),
    .B2(net5278),
    .A2(_04481_),
    .A1(net5069));
 sg13g2_o21ai_1 _13061_ (.B1(_04288_),
    .Y(_04489_),
    .A1(_04289_),
    .A2(_04488_));
 sg13g2_xor2_1 _13062_ (.B(_04415_),
    .A(\m_sys.m_core.m_bru.io_i_pc[10] ),
    .X(_04490_));
 sg13g2_nand2_1 _13063_ (.Y(_04491_),
    .A(net4958),
    .B(_04490_));
 sg13g2_a22oi_1 _13064_ (.Y(_04492_),
    .B1(_04491_),
    .B2(net4748),
    .A2(_04489_),
    .A1(_04479_));
 sg13g2_nand2_1 _13065_ (.Y(_04493_),
    .A(\m_sys.m_core.m_gpr._GEN[106] ),
    .B(net5062));
 sg13g2_a221oi_1 _13066_ (.B2(\m_sys.m_core.m_gpr._GEN[74] ),
    .C1(net5327),
    .B1(net5050),
    .A1(\m_sys.m_core.m_gpr._GEN[42] ),
    .Y(_04494_),
    .A2(net5185));
 sg13g2_mux4_1 _13067_ (.S0(net5324),
    .A0(\m_sys.m_core.m_gpr._GEN[138] ),
    .A1(\m_sys.m_core.m_gpr._GEN[170] ),
    .A2(\m_sys.m_core.m_gpr._GEN[202] ),
    .A3(\m_sys.m_core.m_gpr._GEN[234] ),
    .S1(net5326),
    .X(_04495_));
 sg13g2_inv_1 _13068_ (.Y(_04496_),
    .A(_04495_));
 sg13g2_a22oi_1 _13069_ (.Y(_04497_),
    .B1(_04496_),
    .B2(net5327),
    .A2(_04494_),
    .A1(_04493_));
 sg13g2_a221oi_1 _13070_ (.B2(net4492),
    .C1(net4959),
    .B1(_04497_),
    .A1(\m_sys.m_core.m_bru.io_i_pc[10] ),
    .Y(_04498_),
    .A2(_04456_));
 sg13g2_nor3_1 _13071_ (.A(net4720),
    .B(_04492_),
    .C(_04498_),
    .Y(_04499_));
 sg13g2_a21o_1 _13072_ (.A2(net4720),
    .A1(net3153),
    .B1(_04499_),
    .X(_00217_));
 sg13g2_nand2_1 _13073_ (.Y(_04500_),
    .A(net4891),
    .B(_04347_));
 sg13g2_nand2_1 _13074_ (.Y(_04501_),
    .A(net4905),
    .B(_03177_));
 sg13g2_o21ai_1 _13075_ (.B1(_04501_),
    .Y(_04502_),
    .A1(_03100_),
    .A2(net4904));
 sg13g2_nand2_1 _13076_ (.Y(_04503_),
    .A(net4925),
    .B(_04502_));
 sg13g2_o21ai_1 _13077_ (.B1(_04503_),
    .Y(_04504_),
    .A1(net4926),
    .A2(_04421_));
 sg13g2_o21ai_1 _13078_ (.B1(_04500_),
    .Y(_04505_),
    .A1(net4886),
    .A2(_04504_));
 sg13g2_a21oi_1 _13079_ (.A1(net4777),
    .A2(_04505_),
    .Y(_04506_),
    .B1(net4764));
 sg13g2_o21ai_1 _13080_ (.B1(_04506_),
    .Y(_04507_),
    .A1(net4777),
    .A2(_04198_));
 sg13g2_o21ai_1 _13081_ (.B1(_04507_),
    .Y(_04508_),
    .A1(net5298),
    .A2(_03181_));
 sg13g2_nand3_1 _13082_ (.B(net4770),
    .C(_03893_),
    .A(net5172),
    .Y(_04509_));
 sg13g2_a21oi_1 _13083_ (.A1(net5298),
    .A2(_03180_),
    .Y(_04510_),
    .B1(net5171));
 sg13g2_a22oi_1 _13084_ (.Y(_04511_),
    .B1(_04510_),
    .B2(_03346_),
    .A2(_04508_),
    .A1(net5171));
 sg13g2_o21ai_1 _13085_ (.B1(_04511_),
    .Y(_04512_),
    .A1(_03895_),
    .A2(_04509_));
 sg13g2_nand3_1 _13086_ (.B(_03352_),
    .C(_04261_),
    .A(_03347_),
    .Y(_04513_));
 sg13g2_nand4_1 _13087_ (.B(_03353_),
    .C(_04262_),
    .A(net5244),
    .Y(_04514_),
    .D(_04513_));
 sg13g2_nand2_1 _13088_ (.Y(_04515_),
    .A(_03171_),
    .B(_03175_));
 sg13g2_and2_1 _13089_ (.A(_03174_),
    .B(_03181_),
    .X(_04516_));
 sg13g2_o21ai_1 _13090_ (.B1(net5169),
    .Y(_04517_),
    .A1(_03174_),
    .A2(_03181_));
 sg13g2_a221oi_1 _13091_ (.B2(_04516_),
    .C1(_04517_),
    .B1(_04515_),
    .A1(_03171_),
    .Y(_04518_),
    .A2(_03182_));
 sg13g2_nor2_1 _13092_ (.A(net5298),
    .B(_04518_),
    .Y(_04519_));
 sg13g2_a221oi_1 _13093_ (.B2(_04519_),
    .C1(net4717),
    .B1(_04514_),
    .A1(net5299),
    .Y(_04520_),
    .A2(_03879_));
 sg13g2_a21o_2 _13094_ (.A2(_04512_),
    .A1(net5256),
    .B1(_04520_),
    .X(_04521_));
 sg13g2_a21oi_1 _13095_ (.A1(_02369_),
    .A2(_04521_),
    .Y(_04522_),
    .B1(net5098));
 sg13g2_a22oi_1 _13096_ (.Y(_04523_),
    .B1(net4387),
    .B2(\m_sys._m_uart_io_b_mem_rdata[9] ),
    .A2(net4497),
    .A1(\m_sys._m_ram_io_b_port_rdata[9] ));
 sg13g2_inv_1 _13097_ (.Y(_04524_),
    .A(_04523_));
 sg13g2_mux2_1 _13098_ (.A0(\m_sys._m_ram_io_b_port_rdata[9] ),
    .A1(\m_sys._m_ram_io_b_port_rdata[17] ),
    .S(net5362),
    .X(_04525_));
 sg13g2_o21ai_1 _13099_ (.B1(net4883),
    .Y(_04526_),
    .A1(net5357),
    .A2(_04525_));
 sg13g2_a21oi_1 _13100_ (.A1(net5358),
    .A2(_03904_),
    .Y(_04527_),
    .B1(_04526_));
 sg13g2_a21o_1 _13101_ (.A2(net4882),
    .A1(\m_sys._m_uart_io_b_mem_rdata[9] ),
    .B1(_04527_),
    .X(_04528_));
 sg13g2_a22oi_1 _13102_ (.Y(_04529_),
    .B1(_04528_),
    .B2(net5278),
    .A2(_04524_),
    .A1(_03533_));
 sg13g2_o21ai_1 _13103_ (.B1(_04288_),
    .Y(_04530_),
    .A1(_04289_),
    .A2(_04529_));
 sg13g2_nand2b_1 _13104_ (.Y(_04531_),
    .B(_04530_),
    .A_N(_04522_));
 sg13g2_nor3_1 _13105_ (.A(_00109_),
    .B(_04412_),
    .C(_04413_),
    .Y(_04532_));
 sg13g2_xor2_1 _13106_ (.B(_04532_),
    .A(net3337),
    .X(_04533_));
 sg13g2_a21oi_1 _13107_ (.A1(net5094),
    .A2(_04533_),
    .Y(_04534_),
    .B1(net4971));
 sg13g2_nor2b_1 _13108_ (.A(net5325),
    .B_N(\m_sys.m_core.m_gpr._GEN[41] ),
    .Y(_04535_));
 sg13g2_a221oi_1 _13109_ (.B2(\m_sys.m_core.m_gpr._GEN[73] ),
    .C1(_04535_),
    .B1(net5053),
    .A1(\m_sys.m_core.m_gpr._GEN[105] ),
    .Y(_04536_),
    .A2(net5062));
 sg13g2_nand2b_1 _13110_ (.Y(_04537_),
    .B(net5148),
    .A_N(\m_sys.m_core.m_gpr._GEN[137] ));
 sg13g2_nand2b_1 _13111_ (.Y(_04538_),
    .B(net5049),
    .A_N(\m_sys.m_core.m_gpr._GEN[169] ));
 sg13g2_a22oi_1 _13112_ (.Y(_04539_),
    .B1(net5052),
    .B2(_02441_),
    .A2(net5061),
    .A1(_02442_));
 sg13g2_nand4_1 _13113_ (.B(_04537_),
    .C(_04538_),
    .A(net5327),
    .Y(_04540_),
    .D(_04539_));
 sg13g2_o21ai_1 _13114_ (.B1(_04540_),
    .Y(_04541_),
    .A1(\m_sys.m_core._m_decoder_io_o_rs1[2] ),
    .A2(_04536_));
 sg13g2_a22oi_1 _13115_ (.Y(_04542_),
    .B1(_04541_),
    .B2(net4492),
    .A2(_04456_),
    .A1(net3337));
 sg13g2_a221oi_1 _13116_ (.B2(net4971),
    .C1(net4718),
    .B1(_04542_),
    .A1(_04531_),
    .Y(_04543_),
    .A2(_04534_));
 sg13g2_a21o_1 _13117_ (.A2(net4720),
    .A1(net3445),
    .B1(_04543_),
    .X(_00218_));
 sg13g2_xor2_1 _13118_ (.B(_04414_),
    .A(\m_sys.m_core.m_bru.io_i_pc[8] ),
    .X(_04544_));
 sg13g2_nand2_1 _13119_ (.Y(_04545_),
    .A(net5245),
    .B(_03333_));
 sg13g2_o21ai_1 _13120_ (.B1(_04545_),
    .Y(_04546_),
    .A1(net5245),
    .A2(_03171_));
 sg13g2_xnor2_1 _13121_ (.Y(_04547_),
    .A(_03176_),
    .B(_04546_));
 sg13g2_nand2_1 _13122_ (.Y(_04548_),
    .A(net5161),
    .B(_04547_));
 sg13g2_a21oi_1 _13123_ (.A1(net5299),
    .A2(_03923_),
    .Y(_04549_),
    .B1(net4716));
 sg13g2_nand2_1 _13124_ (.Y(_04550_),
    .A(net4950),
    .B(_04233_));
 sg13g2_a21oi_1 _13125_ (.A1(net4896),
    .A2(_03177_),
    .Y(_04551_),
    .B1(_03591_));
 sg13g2_nor2_1 _13126_ (.A(net4925),
    .B(_04462_),
    .Y(_04552_));
 sg13g2_a21oi_1 _13127_ (.A1(net4924),
    .A2(_04551_),
    .Y(_04553_),
    .B1(_04552_));
 sg13g2_nor2_1 _13128_ (.A(net4886),
    .B(_04553_),
    .Y(_04554_));
 sg13g2_a21oi_1 _13129_ (.A1(net4891),
    .A2(_04382_),
    .Y(_04555_),
    .B1(_04554_));
 sg13g2_a21oi_1 _13130_ (.A1(net4779),
    .A2(_04555_),
    .Y(_04556_),
    .B1(net5162));
 sg13g2_a21oi_1 _13131_ (.A1(_04550_),
    .A2(_04556_),
    .Y(_04557_),
    .B1(net4769));
 sg13g2_nor3_1 _13132_ (.A(net4892),
    .B(_03935_),
    .C(_03936_),
    .Y(_04558_));
 sg13g2_nor2_1 _13133_ (.A(_04557_),
    .B(_04558_),
    .Y(_04559_));
 sg13g2_a21o_1 _13134_ (.A2(_03176_),
    .A1(net5161),
    .B1(net5288),
    .X(_04560_));
 sg13g2_nand2_1 _13135_ (.Y(_04561_),
    .A(net5298),
    .B(_03174_));
 sg13g2_nand3_1 _13136_ (.B(_03175_),
    .C(_04561_),
    .A(net5288),
    .Y(_04562_));
 sg13g2_o21ai_1 _13137_ (.B1(_04562_),
    .Y(_04563_),
    .A1(_04559_),
    .A2(_04560_));
 sg13g2_a22oi_1 _13138_ (.Y(_04564_),
    .B1(_04563_),
    .B2(net5255),
    .A2(_04549_),
    .A1(_04548_));
 sg13g2_o21ai_1 _13139_ (.B1(net5101),
    .Y(_04565_),
    .A1(net5309),
    .A2(_04564_));
 sg13g2_a22oi_1 _13140_ (.Y(_04566_),
    .B1(net4387),
    .B2(\m_sys._m_uart_io_b_mem_rdata[8] ),
    .A2(net4493),
    .A1(\m_sys._m_ram_io_b_port_rdata[8] ));
 sg13g2_inv_1 _13141_ (.Y(_04567_),
    .A(_04566_));
 sg13g2_mux2_1 _13142_ (.A0(\m_sys._m_ram_io_b_port_rdata[8] ),
    .A1(\m_sys._m_ram_io_b_port_rdata[16] ),
    .S(net5362),
    .X(_04568_));
 sg13g2_o21ai_1 _13143_ (.B1(net4883),
    .Y(_04569_),
    .A1(net5357),
    .A2(_04568_));
 sg13g2_a21oi_1 _13144_ (.A1(net5357),
    .A2(_03944_),
    .Y(_04570_),
    .B1(_04569_));
 sg13g2_a21o_1 _13145_ (.A2(net4882),
    .A1(\m_sys._m_uart_io_b_mem_rdata[8] ),
    .B1(_04570_),
    .X(_04571_));
 sg13g2_a22oi_1 _13146_ (.Y(_04572_),
    .B1(_04571_),
    .B2(net5278),
    .A2(_04567_),
    .A1(net5069));
 sg13g2_o21ai_1 _13147_ (.B1(_04288_),
    .Y(_04573_),
    .A1(_04289_),
    .A2(_04572_));
 sg13g2_a22oi_1 _13148_ (.Y(_04574_),
    .B1(_04565_),
    .B2(_04573_),
    .A2(_04544_),
    .A1(net5094));
 sg13g2_a22oi_1 _13149_ (.Y(_04575_),
    .B1(net5047),
    .B2(\m_sys.m_core.m_gpr._GEN[168] ),
    .A2(net5066),
    .A1(\m_sys.m_core.m_gpr._GEN[232] ));
 sg13g2_a221oi_1 _13150_ (.B2(\m_sys.m_core.m_gpr._GEN[200] ),
    .C1(net5182),
    .B1(net5057),
    .A1(\m_sys.m_core.m_gpr._GEN[136] ),
    .Y(_04576_),
    .A2(net5151));
 sg13g2_nand2_1 _13151_ (.Y(_04577_),
    .A(\m_sys.m_core.m_gpr._GEN[104] ),
    .B(net5066));
 sg13g2_a221oi_1 _13152_ (.B2(\m_sys.m_core.m_gpr._GEN[72] ),
    .C1(net5330),
    .B1(net5057),
    .A1(\m_sys.m_core.m_gpr._GEN[40] ),
    .Y(_04578_),
    .A2(net5189));
 sg13g2_a22oi_1 _13153_ (.Y(_04579_),
    .B1(_04577_),
    .B2(_04578_),
    .A2(_04576_),
    .A1(_04575_));
 sg13g2_a22oi_1 _13154_ (.Y(_04580_),
    .B1(_04579_),
    .B2(net4386),
    .A2(_04457_),
    .A1(net3447));
 sg13g2_o21ai_1 _13155_ (.B1(_04580_),
    .Y(_04581_),
    .A1(net4971),
    .A2(_04574_));
 sg13g2_mux2_1 _13156_ (.A0(_04581_),
    .A1(net5320),
    .S(net4718),
    .X(_00219_));
 sg13g2_nand2_1 _13157_ (.Y(_04582_),
    .A(_03119_),
    .B(_03170_));
 sg13g2_nor2_1 _13158_ (.A(_03167_),
    .B(_04582_),
    .Y(_04583_));
 sg13g2_nor2_1 _13159_ (.A(net5245),
    .B(_04583_),
    .Y(_04584_));
 sg13g2_a21oi_1 _13160_ (.A1(_03311_),
    .A2(_03325_),
    .Y(_04585_),
    .B1(_03329_));
 sg13g2_a21o_1 _13161_ (.A2(_03307_),
    .A1(_03119_),
    .B1(_04585_),
    .X(_04586_));
 sg13g2_nand2_1 _13162_ (.Y(_04587_),
    .A(_03330_),
    .B(_04586_));
 sg13g2_a22oi_1 _13163_ (.Y(_04588_),
    .B1(_04587_),
    .B2(net5245),
    .A2(_04584_),
    .A1(_03119_));
 sg13g2_a21oi_1 _13164_ (.A1(_03305_),
    .A2(_04588_),
    .Y(_04589_),
    .B1(net5297));
 sg13g2_o21ai_1 _13165_ (.B1(_04589_),
    .Y(_04590_),
    .A1(_03305_),
    .A2(_04588_));
 sg13g2_a21oi_1 _13166_ (.A1(net5297),
    .A2(_03970_),
    .Y(_04591_),
    .B1(net4716));
 sg13g2_nor3_2 _13167_ (.A(net4768),
    .B(_03977_),
    .C(_03979_),
    .Y(_04592_));
 sg13g2_and2_1 _13168_ (.A(_03419_),
    .B(_03435_),
    .X(_04593_));
 sg13g2_nor2_1 _13169_ (.A(net4925),
    .B(_04502_),
    .Y(_04594_));
 sg13g2_a21oi_1 _13170_ (.A1(net4924),
    .A2(_04593_),
    .Y(_04595_),
    .B1(_04594_));
 sg13g2_nand2_1 _13171_ (.Y(_04596_),
    .A(net4774),
    .B(_04595_));
 sg13g2_a21oi_1 _13172_ (.A1(net4886),
    .A2(_04423_),
    .Y(_04597_),
    .B1(net4946));
 sg13g2_a221oi_1 _13173_ (.B2(_04597_),
    .C1(net4764),
    .B1(_04596_),
    .A1(net4946),
    .Y(_04598_),
    .A2(_04277_));
 sg13g2_o21ai_1 _13174_ (.B1(net5170),
    .Y(_04599_),
    .A1(net5297),
    .A2(_03305_));
 sg13g2_nor3_1 _13175_ (.A(_04592_),
    .B(_04598_),
    .C(_04599_),
    .Y(_04600_));
 sg13g2_a21oi_1 _13176_ (.A1(net5161),
    .A2(_03115_),
    .Y(_04601_),
    .B1(net5170));
 sg13g2_a21oi_1 _13177_ (.A1(_03113_),
    .A2(_04601_),
    .Y(_04602_),
    .B1(_04600_));
 sg13g2_a22oi_1 _13178_ (.Y(_04603_),
    .B1(_04602_),
    .B2(net5255),
    .A2(_04591_),
    .A1(_04590_));
 sg13g2_a21oi_1 _13179_ (.A1(net5232),
    .A2(_04603_),
    .Y(_04604_),
    .B1(net5097));
 sg13g2_o21ai_1 _13180_ (.B1(net5097),
    .Y(_04605_),
    .A1(_03538_),
    .A2(_03548_));
 sg13g2_nor2_1 _13181_ (.A(_03519_),
    .B(_04605_),
    .Y(_04606_));
 sg13g2_nor2_1 _13182_ (.A(_00023_),
    .B(_04412_),
    .Y(_04607_));
 sg13g2_xnor2_1 _13183_ (.Y(_04608_),
    .A(net3313),
    .B(_04607_));
 sg13g2_a21oi_1 _13184_ (.A1(net5095),
    .A2(_04608_),
    .Y(_04609_),
    .B1(net4971));
 sg13g2_o21ai_1 _13185_ (.B1(_04609_),
    .Y(_04610_),
    .A1(_04604_),
    .A2(_04606_));
 sg13g2_a22oi_1 _13186_ (.Y(_04611_),
    .B1(net5049),
    .B2(\m_sys.m_core.m_gpr._GEN[167] ),
    .A2(net5061),
    .A1(\m_sys.m_core.m_gpr._GEN[231] ));
 sg13g2_a221oi_1 _13187_ (.B2(\m_sys.m_core.m_gpr._GEN[199] ),
    .C1(net5179),
    .B1(net5052),
    .A1(\m_sys.m_core.m_gpr._GEN[135] ),
    .Y(_04612_),
    .A2(net5149));
 sg13g2_nand2_1 _13188_ (.Y(_04613_),
    .A(\m_sys.m_core.m_gpr._GEN[103] ),
    .B(net5061));
 sg13g2_a221oi_1 _13189_ (.B2(\m_sys.m_core.m_gpr._GEN[71] ),
    .C1(net5327),
    .B1(net5052),
    .A1(\m_sys.m_core.m_gpr._GEN[39] ),
    .Y(_04614_),
    .A2(net5185));
 sg13g2_a22oi_1 _13190_ (.Y(_04615_),
    .B1(_04613_),
    .B2(_04614_),
    .A2(_04612_),
    .A1(_04611_));
 sg13g2_a221oi_1 _13191_ (.B2(net4386),
    .C1(net4718),
    .B1(_04615_),
    .A1(net3313),
    .Y(_04616_),
    .A2(_04457_));
 sg13g2_a22oi_1 _13192_ (.Y(_00220_),
    .B1(_04610_),
    .B2(_04616_),
    .A2(net4718),
    .A1(net5227));
 sg13g2_nand2_1 _13193_ (.Y(_04617_),
    .A(net3433),
    .B(net4719));
 sg13g2_xnor2_1 _13194_ (.Y(_04618_),
    .A(_03308_),
    .B(_04585_));
 sg13g2_nand2_1 _13195_ (.Y(_04619_),
    .A(_03167_),
    .B(_04582_));
 sg13g2_a221oi_1 _13196_ (.B2(_04584_),
    .C1(net5297),
    .B1(_04619_),
    .A1(net5245),
    .Y(_04620_),
    .A2(_04618_));
 sg13g2_inv_1 _13197_ (.Y(_04621_),
    .A(_04620_));
 sg13g2_a21oi_1 _13198_ (.A1(net5297),
    .A2(_04004_),
    .Y(_04622_),
    .B1(net4716));
 sg13g2_nor3_2 _13199_ (.A(_03410_),
    .B(_04011_),
    .C(_04014_),
    .Y(_04623_));
 sg13g2_o21ai_1 _13200_ (.B1(_03590_),
    .Y(_04624_),
    .A1(_03118_),
    .A2(net4896));
 sg13g2_nor2_1 _13201_ (.A(net4912),
    .B(_04624_),
    .Y(_04625_));
 sg13g2_a21oi_1 _13202_ (.A1(net4915),
    .A2(_04551_),
    .Y(_04626_),
    .B1(_04625_));
 sg13g2_nand2_1 _13203_ (.Y(_04627_),
    .A(net4774),
    .B(_04626_));
 sg13g2_a21oi_1 _13204_ (.A1(net4886),
    .A2(_04464_),
    .Y(_04628_),
    .B1(net4946));
 sg13g2_a221oi_1 _13205_ (.B2(_04628_),
    .C1(net4764),
    .B1(_04627_),
    .A1(net4946),
    .Y(_04629_),
    .A2(_04309_));
 sg13g2_o21ai_1 _13206_ (.B1(net5171),
    .Y(_04630_),
    .A1(net5297),
    .A2(_04582_));
 sg13g2_nor3_1 _13207_ (.A(_04623_),
    .B(_04629_),
    .C(_04630_),
    .Y(_04631_));
 sg13g2_nand2_1 _13208_ (.Y(_04632_),
    .A(net5161),
    .B(_03307_));
 sg13g2_nand3_1 _13209_ (.B(_03119_),
    .C(_04632_),
    .A(net5288),
    .Y(_04633_));
 sg13g2_nor2_1 _13210_ (.A(net5160),
    .B(_04631_),
    .Y(_04634_));
 sg13g2_a22oi_1 _13211_ (.Y(_04635_),
    .B1(_04633_),
    .B2(_04634_),
    .A2(_04622_),
    .A1(_04621_));
 sg13g2_mux2_1 _13212_ (.A0(_00134_),
    .A1(_00133_),
    .S(_03498_),
    .X(_04636_));
 sg13g2_mux2_1 _13213_ (.A0(_00060_),
    .A1(_04636_),
    .S(_02698_),
    .X(_04637_));
 sg13g2_mux2_1 _13214_ (.A0(_00060_),
    .A1(_00061_),
    .S(net5361),
    .X(_04638_));
 sg13g2_a21oi_1 _13215_ (.A1(net5355),
    .A2(_04022_),
    .Y(_04639_),
    .B1(net5072));
 sg13g2_o21ai_1 _13216_ (.B1(_04639_),
    .Y(_04640_),
    .A1(net5355),
    .A2(_04638_));
 sg13g2_a22oi_1 _13217_ (.Y(_04641_),
    .B1(net4882),
    .B2(_00134_),
    .A2(_03511_),
    .A1(_00133_));
 sg13g2_nand2_1 _13218_ (.Y(_04642_),
    .A(_04640_),
    .B(_04641_));
 sg13g2_a221oi_1 _13219_ (.B2(net5276),
    .C1(_04605_),
    .B1(_04642_),
    .A1(net5069),
    .Y(_04643_),
    .A2(_04637_));
 sg13g2_nor2_1 _13220_ (.A(net4748),
    .B(_04643_),
    .Y(_04644_));
 sg13g2_o21ai_1 _13221_ (.B1(_04644_),
    .Y(_04645_),
    .A1(net5097),
    .A2(_04635_));
 sg13g2_mux4_1 _13222_ (.S0(net5324),
    .A0(\m_sys.m_core.m_gpr._GEN[134] ),
    .A1(\m_sys.m_core.m_gpr._GEN[166] ),
    .A2(\m_sys.m_core.m_gpr._GEN[198] ),
    .A3(\m_sys.m_core.m_gpr._GEN[230] ),
    .S1(net5326),
    .X(_04646_));
 sg13g2_nand2b_1 _13223_ (.Y(_04647_),
    .B(net5052),
    .A_N(\m_sys.m_core.m_gpr._GEN[70] ));
 sg13g2_o21ai_1 _13224_ (.B1(_04647_),
    .Y(_04648_),
    .A1(\m_sys.m_core.m_gpr._GEN[38] ),
    .A2(net5326));
 sg13g2_a21oi_1 _13225_ (.A1(_02435_),
    .A2(net5061),
    .Y(_04649_),
    .B1(_04648_));
 sg13g2_mux2_2 _13226_ (.A0(_04646_),
    .A1(_04649_),
    .S(net5179),
    .X(_04650_));
 sg13g2_a221oi_1 _13227_ (.B2(net4492),
    .C1(net4960),
    .B1(_04650_),
    .A1(net3250),
    .Y(_04651_),
    .A2(_04456_));
 sg13g2_xor2_1 _13228_ (.B(_04412_),
    .A(\m_sys.m_core.m_bru.io_i_pc[6] ),
    .X(_04652_));
 sg13g2_a21oi_1 _13229_ (.A1(net5095),
    .A2(_04652_),
    .Y(_04653_),
    .B1(net4719));
 sg13g2_nand2_1 _13230_ (.Y(_04654_),
    .A(_04645_),
    .B(_04653_));
 sg13g2_o21ai_1 _13231_ (.B1(_04617_),
    .Y(_00221_),
    .A1(_04651_),
    .A2(_04654_));
 sg13g2_a22oi_1 _13232_ (.Y(_04655_),
    .B1(net4387),
    .B2(_00132_),
    .A2(net4494),
    .A1(_00058_));
 sg13g2_or2_1 _13233_ (.X(_04656_),
    .B(_04655_),
    .A(net4879));
 sg13g2_nor2_1 _13234_ (.A(_03498_),
    .B(net4878),
    .Y(_04657_));
 sg13g2_a21oi_2 _13235_ (.B1(_04657_),
    .Y(_04658_),
    .A2(_04323_),
    .A1(net5276));
 sg13g2_mux2_1 _13236_ (.A0(_00058_),
    .A1(_00059_),
    .S(net5361),
    .X(_04659_));
 sg13g2_a21oi_1 _13237_ (.A1(net5355),
    .A2(_04061_),
    .Y(_04660_),
    .B1(net5073));
 sg13g2_o21ai_1 _13238_ (.B1(_04660_),
    .Y(_04661_),
    .A1(net5356),
    .A2(_04659_));
 sg13g2_o21ai_1 _13239_ (.B1(_04661_),
    .Y(_04662_),
    .A1(_02500_),
    .A2(net4881));
 sg13g2_a221oi_1 _13240_ (.B2(net5280),
    .C1(_04605_),
    .B1(_04662_),
    .A1(_00131_),
    .Y(_04663_),
    .A2(_04658_));
 sg13g2_a21oi_1 _13241_ (.A1(_03150_),
    .A2(_03156_),
    .Y(_04664_),
    .B1(_03154_));
 sg13g2_o21ai_1 _13242_ (.B1(net5169),
    .Y(_04665_),
    .A1(_03163_),
    .A2(_04664_));
 sg13g2_a21oi_1 _13243_ (.A1(_03163_),
    .A2(_04664_),
    .Y(_04666_),
    .B1(_04665_));
 sg13g2_or2_1 _13244_ (.X(_04667_),
    .B(_03327_),
    .A(_03325_));
 sg13g2_o21ai_1 _13245_ (.B1(net5246),
    .Y(_04668_),
    .A1(_03311_),
    .A2(_04667_));
 sg13g2_a21oi_1 _13246_ (.A1(_03311_),
    .A2(_04667_),
    .Y(_04669_),
    .B1(_04668_));
 sg13g2_or3_1 _13247_ (.A(net5296),
    .B(_04666_),
    .C(_04669_),
    .X(_04670_));
 sg13g2_a21oi_1 _13248_ (.A1(net5299),
    .A2(_04040_),
    .Y(_04671_),
    .B1(net4716));
 sg13g2_a21oi_1 _13249_ (.A1(net5246),
    .A2(_04051_),
    .Y(_04672_),
    .B1(net4767));
 sg13g2_nor2_1 _13250_ (.A(net4779),
    .B(_04349_),
    .Y(_04673_));
 sg13g2_nand2_1 _13251_ (.Y(_04674_),
    .A(net4904),
    .B(_03159_));
 sg13g2_o21ai_1 _13252_ (.B1(_04674_),
    .Y(_04675_),
    .A1(_03118_),
    .A2(net4904));
 sg13g2_nand2_1 _13253_ (.Y(_04676_),
    .A(net4913),
    .B(_04593_));
 sg13g2_o21ai_1 _13254_ (.B1(_04676_),
    .Y(_04677_),
    .A1(net4912),
    .A2(_04675_));
 sg13g2_o21ai_1 _13255_ (.B1(net4777),
    .Y(_04678_),
    .A1(net4885),
    .A2(_04677_));
 sg13g2_a21oi_1 _13256_ (.A1(net4886),
    .A2(_04504_),
    .Y(_04679_),
    .B1(_04678_));
 sg13g2_nor2_1 _13257_ (.A(_04673_),
    .B(_04679_),
    .Y(_04680_));
 sg13g2_o21ai_1 _13258_ (.B1(net5171),
    .Y(_04681_),
    .A1(net5297),
    .A2(_03163_));
 sg13g2_a221oi_1 _13259_ (.B2(net4765),
    .C1(_04681_),
    .B1(_04680_),
    .A1(_04054_),
    .Y(_04682_),
    .A2(_04672_));
 sg13g2_a21oi_1 _13260_ (.A1(_03158_),
    .A2(_03310_),
    .Y(_04683_),
    .B1(net5297));
 sg13g2_nand2_1 _13261_ (.Y(_04684_),
    .A(net5288),
    .B(_03160_));
 sg13g2_o21ai_1 _13262_ (.B1(net5255),
    .Y(_04685_),
    .A1(_04683_),
    .A2(_04684_));
 sg13g2_nor2_1 _13263_ (.A(_04682_),
    .B(_04685_),
    .Y(_04686_));
 sg13g2_a21oi_2 _13264_ (.B1(_04686_),
    .Y(_04687_),
    .A2(_04671_),
    .A1(_04670_));
 sg13g2_nand2_1 _13265_ (.Y(_04688_),
    .A(net5232),
    .B(_04687_));
 sg13g2_a22oi_1 _13266_ (.Y(_04689_),
    .B1(_04688_),
    .B2(net5101),
    .A2(_04663_),
    .A1(_04656_));
 sg13g2_nor2_1 _13267_ (.A(_00009_),
    .B(_04411_),
    .Y(_04690_));
 sg13g2_xor2_1 _13268_ (.B(_04690_),
    .A(\m_sys.m_core.m_bru.io_i_pc[5] ),
    .X(_04691_));
 sg13g2_o21ai_1 _13269_ (.B1(net4960),
    .Y(_04692_),
    .A1(net5093),
    .A2(_04691_));
 sg13g2_a22oi_1 _13270_ (.Y(_04693_),
    .B1(net5046),
    .B2(\m_sys.m_core.m_gpr._GEN[165] ),
    .A2(net5059),
    .A1(\m_sys.m_core.m_gpr._GEN[229] ));
 sg13g2_a221oi_1 _13271_ (.B2(\m_sys.m_core.m_gpr._GEN[197] ),
    .C1(net5178),
    .B1(net5050),
    .A1(\m_sys.m_core.m_gpr._GEN[133] ),
    .Y(_04694_),
    .A2(net5149));
 sg13g2_nand2_1 _13272_ (.Y(_04695_),
    .A(\m_sys.m_core.m_gpr._GEN[101] ),
    .B(net5059));
 sg13g2_a221oi_1 _13273_ (.B2(\m_sys.m_core.m_gpr._GEN[69] ),
    .C1(net5328),
    .B1(net5050),
    .A1(\m_sys.m_core.m_gpr._GEN[37] ),
    .Y(_04696_),
    .A2(net5184));
 sg13g2_a22oi_1 _13274_ (.Y(_04697_),
    .B1(_04695_),
    .B2(_04696_),
    .A2(_04694_),
    .A1(_04693_));
 sg13g2_a22oi_1 _13275_ (.Y(_04698_),
    .B1(_04697_),
    .B2(net4386),
    .A2(_04457_),
    .A1(net3446));
 sg13g2_o21ai_1 _13276_ (.B1(_04698_),
    .Y(_04699_),
    .A1(_04689_),
    .A2(_04692_));
 sg13g2_mux2_1 _13277_ (.A0(_04699_),
    .A1(net5318),
    .S(net4718),
    .X(_00222_));
 sg13g2_nand2_1 _13278_ (.Y(_04700_),
    .A(net5315),
    .B(net4718));
 sg13g2_mux2_1 _13279_ (.A0(_03150_),
    .A1(_03324_),
    .S(net5245),
    .X(_04701_));
 sg13g2_o21ai_1 _13280_ (.B1(net5161),
    .Y(_04702_),
    .A1(_03157_),
    .A2(_04701_));
 sg13g2_a21oi_1 _13281_ (.A1(_03157_),
    .A2(_04701_),
    .Y(_04703_),
    .B1(_04702_));
 sg13g2_nor2_1 _13282_ (.A(net5161),
    .B(_04077_),
    .Y(_04704_));
 sg13g2_nor3_1 _13283_ (.A(net4716),
    .B(_04703_),
    .C(_04704_),
    .Y(_04705_));
 sg13g2_nor3_2 _13284_ (.A(net4768),
    .B(_04088_),
    .C(_04090_),
    .Y(_04706_));
 sg13g2_nand2b_1 _13285_ (.Y(_04707_),
    .B(net4885),
    .A_N(_04553_));
 sg13g2_a21oi_1 _13286_ (.A1(net4896),
    .A2(_03159_),
    .Y(_04708_),
    .B1(_03578_));
 sg13g2_nand2_1 _13287_ (.Y(_04709_),
    .A(net4912),
    .B(_04624_));
 sg13g2_o21ai_1 _13288_ (.B1(_04709_),
    .Y(_04710_),
    .A1(net4912),
    .A2(_04708_));
 sg13g2_o21ai_1 _13289_ (.B1(_04707_),
    .Y(_04711_),
    .A1(net4885),
    .A2(_04710_));
 sg13g2_o21ai_1 _13290_ (.B1(net4766),
    .Y(_04712_),
    .A1(net4780),
    .A2(_04384_));
 sg13g2_a21oi_1 _13291_ (.A1(net4777),
    .A2(_04711_),
    .Y(_04713_),
    .B1(_04712_));
 sg13g2_o21ai_1 _13292_ (.B1(net5170),
    .Y(_04714_),
    .A1(net5296),
    .A2(_03157_));
 sg13g2_nor3_1 _13293_ (.A(_04706_),
    .B(_04713_),
    .C(_04714_),
    .Y(_04715_));
 sg13g2_a21oi_1 _13294_ (.A1(net5161),
    .A2(_03156_),
    .Y(_04716_),
    .B1(net5170));
 sg13g2_a21oi_1 _13295_ (.A1(_03155_),
    .A2(_04716_),
    .Y(_04717_),
    .B1(_04715_));
 sg13g2_a21oi_2 _13296_ (.B1(_04705_),
    .Y(_04718_),
    .A2(_04717_),
    .A1(net5255));
 sg13g2_mux2_1 _13297_ (.A0(_00130_),
    .A1(_00129_),
    .S(_03498_),
    .X(_04719_));
 sg13g2_mux2_1 _13298_ (.A0(_00056_),
    .A1(_04719_),
    .S(_02698_),
    .X(_04720_));
 sg13g2_mux2_1 _13299_ (.A0(_00056_),
    .A1(_00057_),
    .S(net5361),
    .X(_04721_));
 sg13g2_a21oi_1 _13300_ (.A1(net5355),
    .A2(_04098_),
    .Y(_04722_),
    .B1(net5072));
 sg13g2_o21ai_1 _13301_ (.B1(_04722_),
    .Y(_04723_),
    .A1(net5354),
    .A2(_04721_));
 sg13g2_a22oi_1 _13302_ (.Y(_04724_),
    .B1(net4882),
    .B2(_00130_),
    .A2(_03511_),
    .A1(_00129_));
 sg13g2_nand2_1 _13303_ (.Y(_04725_),
    .A(_04723_),
    .B(_04724_));
 sg13g2_a221oi_1 _13304_ (.B2(net5276),
    .C1(_04605_),
    .B1(_04725_),
    .A1(net5069),
    .Y(_04726_),
    .A2(_04720_));
 sg13g2_nor2_1 _13305_ (.A(net4748),
    .B(_04726_),
    .Y(_04727_));
 sg13g2_o21ai_1 _13306_ (.B1(_04727_),
    .Y(_04728_),
    .A1(net5097),
    .A2(_04718_));
 sg13g2_mux4_1 _13307_ (.S0(net5324),
    .A0(\m_sys.m_core.m_gpr._GEN[132] ),
    .A1(\m_sys.m_core.m_gpr._GEN[164] ),
    .A2(\m_sys.m_core.m_gpr._GEN[196] ),
    .A3(\m_sys.m_core.m_gpr._GEN[228] ),
    .S1(net5326),
    .X(_04729_));
 sg13g2_nand2b_1 _13308_ (.Y(_04730_),
    .B(net5061),
    .A_N(\m_sys.m_core.m_gpr._GEN[100] ));
 sg13g2_o21ai_1 _13309_ (.B1(_04730_),
    .Y(_04731_),
    .A1(\m_sys.m_core.m_gpr._GEN[36] ),
    .A2(net5325));
 sg13g2_a21oi_1 _13310_ (.A1(_02431_),
    .A2(net5052),
    .Y(_04732_),
    .B1(_04731_));
 sg13g2_mux2_2 _13311_ (.A0(_04729_),
    .A1(_04732_),
    .S(net5179),
    .X(_04733_));
 sg13g2_a221oi_1 _13312_ (.B2(net4492),
    .C1(net4960),
    .B1(_04733_),
    .A1(net3385),
    .Y(_04734_),
    .A2(_04456_));
 sg13g2_xnor2_1 _13313_ (.Y(_04735_),
    .A(_02362_),
    .B(_04411_));
 sg13g2_a21oi_1 _13314_ (.A1(net5095),
    .A2(_04735_),
    .Y(_04736_),
    .B1(net4718));
 sg13g2_nand2_1 _13315_ (.Y(_04737_),
    .A(_04728_),
    .B(_04736_));
 sg13g2_o21ai_1 _13316_ (.B1(_04700_),
    .Y(_00223_),
    .A1(_04734_),
    .A2(_04737_));
 sg13g2_nand2_1 _13317_ (.Y(_04738_),
    .A(net5313),
    .B(net4719));
 sg13g2_xnor2_1 _13318_ (.Y(_04739_),
    .A(\m_sys.m_core.m_bru.io_i_pc[3] ),
    .B(\m_sys.m_core.m_bru.io_i_pc[2] ));
 sg13g2_nor4_2 _13319_ (.A(net5292),
    .B(net4768),
    .C(_04128_),
    .Y(_04740_),
    .D(_04131_));
 sg13g2_nor2_1 _13320_ (.A(net5170),
    .B(_03125_),
    .Y(_04741_));
 sg13g2_o21ai_1 _13321_ (.B1(_04741_),
    .Y(_04742_),
    .A1(net5161),
    .A2(_03126_));
 sg13g2_nor2_1 _13322_ (.A(net5295),
    .B(_03322_),
    .Y(_04743_));
 sg13g2_nor2_1 _13323_ (.A(_03426_),
    .B(_03432_),
    .Y(_04744_));
 sg13g2_a21oi_1 _13324_ (.A1(net4927),
    .A2(_04744_),
    .Y(_04745_),
    .B1(net4887));
 sg13g2_o21ai_1 _13325_ (.B1(_04745_),
    .Y(_04746_),
    .A1(net4927),
    .A2(_04675_));
 sg13g2_a21oi_1 _13326_ (.A1(net4885),
    .A2(_04595_),
    .Y(_04747_),
    .B1(net4946));
 sg13g2_a221oi_1 _13327_ (.B2(_04747_),
    .C1(net4764),
    .B1(_04746_),
    .A1(net4946),
    .Y(_04748_),
    .A2(_04424_));
 sg13g2_o21ai_1 _13328_ (.B1(net5170),
    .Y(_04749_),
    .A1(_04743_),
    .A2(_04748_));
 sg13g2_nand2_1 _13329_ (.Y(_04750_),
    .A(_04742_),
    .B(_04749_));
 sg13g2_o21ai_1 _13330_ (.B1(net5255),
    .Y(_04751_),
    .A1(_04740_),
    .A2(_04750_));
 sg13g2_o21ai_1 _13331_ (.B1(net5246),
    .Y(_04752_),
    .A1(_03315_),
    .A2(_03320_));
 sg13g2_nand2b_1 _13332_ (.Y(_04753_),
    .B(_03144_),
    .A_N(_04752_));
 sg13g2_o21ai_1 _13333_ (.B1(_04753_),
    .Y(_04754_),
    .A1(net5246),
    .A2(_03148_));
 sg13g2_a21oi_1 _13334_ (.A1(net5296),
    .A2(_04119_),
    .Y(_04755_),
    .B1(net4716));
 sg13g2_xnor2_1 _13335_ (.Y(_04756_),
    .A(_03322_),
    .B(_04754_));
 sg13g2_o21ai_1 _13336_ (.B1(_04755_),
    .Y(_04757_),
    .A1(net5295),
    .A2(_04756_));
 sg13g2_nand2_2 _13337_ (.Y(_04758_),
    .A(_04751_),
    .B(_04757_));
 sg13g2_a22oi_1 _13338_ (.Y(_04759_),
    .B1(net4387),
    .B2(_00128_),
    .A2(net4494),
    .A1(_00054_));
 sg13g2_or2_1 _13339_ (.X(_04760_),
    .B(_04759_),
    .A(net4879));
 sg13g2_mux2_1 _13340_ (.A0(_00054_),
    .A1(_00055_),
    .S(net5360),
    .X(_04761_));
 sg13g2_a21oi_1 _13341_ (.A1(net5355),
    .A2(_04138_),
    .Y(_04762_),
    .B1(net5072));
 sg13g2_o21ai_1 _13342_ (.B1(_04762_),
    .Y(_04763_),
    .A1(net5354),
    .A2(_04761_));
 sg13g2_o21ai_1 _13343_ (.B1(_04763_),
    .Y(_04764_),
    .A1(_02499_),
    .A2(net4881));
 sg13g2_a221oi_1 _13344_ (.B2(net5275),
    .C1(_04605_),
    .B1(_04764_),
    .A1(_00127_),
    .Y(_04765_),
    .A2(_04658_));
 sg13g2_a221oi_1 _13345_ (.B2(_04765_),
    .C1(net5094),
    .B1(_04760_),
    .A1(net5101),
    .Y(_04766_),
    .A2(_04758_));
 sg13g2_a21oi_1 _13346_ (.A1(net5095),
    .A2(_04739_),
    .Y(_04767_),
    .B1(_04766_));
 sg13g2_nor2b_1 _13347_ (.A(net5326),
    .B_N(\m_sys.m_core.m_gpr._GEN[35] ),
    .Y(_04768_));
 sg13g2_a221oi_1 _13348_ (.B2(\m_sys.m_core.m_gpr._GEN[67] ),
    .C1(_04768_),
    .B1(net5057),
    .A1(\m_sys.m_core.m_gpr._GEN[99] ),
    .Y(_04769_),
    .A2(net5066));
 sg13g2_nand2b_1 _13349_ (.Y(_04770_),
    .B(net5151),
    .A_N(\m_sys.m_core.m_gpr._GEN[131] ));
 sg13g2_nand2b_1 _13350_ (.Y(_04771_),
    .B(net5066),
    .A_N(\m_sys.m_core.m_gpr._GEN[227] ));
 sg13g2_a22oi_1 _13351_ (.Y(_04772_),
    .B1(net5047),
    .B2(_02428_),
    .A2(net5057),
    .A1(_02429_));
 sg13g2_nand4_1 _13352_ (.B(_04770_),
    .C(_04771_),
    .A(net5330),
    .Y(_04773_),
    .D(_04772_));
 sg13g2_o21ai_1 _13353_ (.B1(_04773_),
    .Y(_04774_),
    .A1(net5330),
    .A2(_04769_));
 sg13g2_a22oi_1 _13354_ (.Y(_04775_),
    .B1(_04774_),
    .B2(net4492),
    .A2(_04456_),
    .A1(\m_sys.m_core.m_bru.io_i_pc[3] ));
 sg13g2_a21oi_1 _13355_ (.A1(net4971),
    .A2(_04775_),
    .Y(_04776_),
    .B1(net4719));
 sg13g2_o21ai_1 _13356_ (.B1(_04776_),
    .Y(_04777_),
    .A1(net4971),
    .A2(_04767_));
 sg13g2_nand2_1 _13357_ (.Y(_00224_),
    .A(_04738_),
    .B(_04777_));
 sg13g2_a21o_1 _13358_ (.A2(_03320_),
    .A1(_03315_),
    .B1(_04752_),
    .X(_04778_));
 sg13g2_nor2_1 _13359_ (.A(_03142_),
    .B(_03146_),
    .Y(_04779_));
 sg13g2_nor3_1 _13360_ (.A(net5245),
    .B(_03147_),
    .C(_04779_),
    .Y(_04780_));
 sg13g2_nor2_1 _13361_ (.A(net5295),
    .B(_04780_),
    .Y(_04781_));
 sg13g2_a221oi_1 _13362_ (.B2(_04781_),
    .C1(net4716),
    .B1(_04778_),
    .A1(net5295),
    .Y(_04782_),
    .A2(_04155_));
 sg13g2_a21oi_1 _13363_ (.A1(net5250),
    .A2(_04162_),
    .Y(_04783_),
    .B1(_04165_));
 sg13g2_a21oi_1 _13364_ (.A1(_03129_),
    .A2(net4774),
    .Y(_04784_),
    .B1(net5295));
 sg13g2_nor3_1 _13365_ (.A(net5170),
    .B(_03130_),
    .C(_04784_),
    .Y(_04785_));
 sg13g2_nor2_1 _13366_ (.A(net5295),
    .B(_03146_),
    .Y(_04786_));
 sg13g2_or3_1 _13367_ (.A(net4912),
    .B(_03577_),
    .C(_03583_),
    .X(_04787_));
 sg13g2_a21oi_1 _13368_ (.A1(net4912),
    .A2(_04708_),
    .Y(_04788_),
    .B1(net4885));
 sg13g2_a22oi_1 _13369_ (.Y(_04789_),
    .B1(_04787_),
    .B2(_04788_),
    .A2(_04626_),
    .A1(net4885));
 sg13g2_mux2_1 _13370_ (.A0(_04465_),
    .A1(_04789_),
    .S(net4776),
    .X(_04790_));
 sg13g2_a21oi_1 _13371_ (.A1(net4765),
    .A2(_04790_),
    .Y(_04791_),
    .B1(_04786_));
 sg13g2_o21ai_1 _13372_ (.B1(_04791_),
    .Y(_04792_),
    .A1(net4767),
    .A2(_04783_));
 sg13g2_a21oi_1 _13373_ (.A1(net5170),
    .A2(_04792_),
    .Y(_04793_),
    .B1(_04785_));
 sg13g2_a21oi_2 _13374_ (.B1(_04782_),
    .Y(_04794_),
    .A2(_04793_),
    .A1(net5255));
 sg13g2_a22oi_1 _13375_ (.Y(_04795_),
    .B1(net4387),
    .B2(_00126_),
    .A2(net4494),
    .A1(_00052_));
 sg13g2_or2_1 _13376_ (.X(_04796_),
    .B(_04795_),
    .A(net4878));
 sg13g2_mux2_1 _13377_ (.A0(_00052_),
    .A1(_00053_),
    .S(net5360),
    .X(_04797_));
 sg13g2_a21oi_1 _13378_ (.A1(net5355),
    .A2(_04174_),
    .Y(_04798_),
    .B1(net5072));
 sg13g2_o21ai_1 _13379_ (.B1(_04798_),
    .Y(_04799_),
    .A1(net5354),
    .A2(_04797_));
 sg13g2_o21ai_1 _13380_ (.B1(_04799_),
    .Y(_04800_),
    .A1(_02498_),
    .A2(net4881));
 sg13g2_a221oi_1 _13381_ (.B2(net5275),
    .C1(_04605_),
    .B1(_04800_),
    .A1(_00125_),
    .Y(_04801_),
    .A2(_04658_));
 sg13g2_a21oi_2 _13382_ (.B1(net5094),
    .Y(_04802_),
    .A2(_04801_),
    .A1(_04796_));
 sg13g2_o21ai_1 _13383_ (.B1(_04802_),
    .Y(_04803_),
    .A1(net5097),
    .A2(_04794_));
 sg13g2_a21oi_1 _13384_ (.A1(_02372_),
    .A2(net5094),
    .Y(_04804_),
    .B1(net4971));
 sg13g2_nand2_1 _13385_ (.Y(_04805_),
    .A(_04803_),
    .B(_04804_));
 sg13g2_a22oi_1 _13386_ (.Y(_04806_),
    .B1(net5047),
    .B2(\m_sys.m_core.m_gpr._GEN[162] ),
    .A2(net5066),
    .A1(\m_sys.m_core.m_gpr._GEN[226] ));
 sg13g2_a221oi_1 _13387_ (.B2(\m_sys.m_core.m_gpr._GEN[194] ),
    .C1(net5182),
    .B1(net5057),
    .A1(\m_sys.m_core.m_gpr._GEN[130] ),
    .Y(_04807_),
    .A2(net5151));
 sg13g2_nand2_1 _13388_ (.Y(_04808_),
    .A(\m_sys.m_core.m_gpr._GEN[98] ),
    .B(net5066));
 sg13g2_a221oi_1 _13389_ (.B2(\m_sys.m_core.m_gpr._GEN[66] ),
    .C1(net5330),
    .B1(net5057),
    .A1(\m_sys.m_core.m_gpr._GEN[34] ),
    .Y(_04809_),
    .A2(net5189));
 sg13g2_a22oi_1 _13390_ (.Y(_04810_),
    .B1(_04808_),
    .B2(_04809_),
    .A2(_04807_),
    .A1(_04806_));
 sg13g2_a221oi_1 _13391_ (.B2(net4386),
    .C1(net4718),
    .B1(_04810_),
    .A1(net3366),
    .Y(_04811_),
    .A2(_04457_));
 sg13g2_a22oi_1 _13392_ (.Y(_00225_),
    .B1(_04805_),
    .B2(_04811_),
    .A2(net4719),
    .A1(net5231));
 sg13g2_nand2_1 _13393_ (.Y(_04812_),
    .A(net5312),
    .B(net4721));
 sg13g2_xnor2_1 _13394_ (.Y(_04813_),
    .A(_03312_),
    .B(_03313_));
 sg13g2_nor2_1 _13395_ (.A(net5245),
    .B(net4904),
    .Y(_04814_));
 sg13g2_xnor2_1 _13396_ (.Y(_04815_),
    .A(_04813_),
    .B(_04814_));
 sg13g2_a21oi_1 _13397_ (.A1(net5296),
    .A2(_04191_),
    .Y(_04816_),
    .B1(net4716));
 sg13g2_o21ai_1 _13398_ (.B1(_04816_),
    .Y(_04817_),
    .A1(net5295),
    .A2(_04815_));
 sg13g2_a21oi_1 _13399_ (.A1(net5253),
    .A2(_04200_),
    .Y(_04818_),
    .B1(net4768));
 sg13g2_nor2b_1 _13400_ (.A(_04203_),
    .B_N(_04818_),
    .Y(_04819_));
 sg13g2_nor2_1 _13401_ (.A(net4912),
    .B(_03428_),
    .Y(_04820_));
 sg13g2_a221oi_1 _13402_ (.B2(_03425_),
    .C1(net4887),
    .B1(_04820_),
    .A1(net4912),
    .Y(_04821_),
    .A2(_04744_));
 sg13g2_o21ai_1 _13403_ (.B1(net4785),
    .Y(_04822_),
    .A1(net4774),
    .A2(_04677_));
 sg13g2_a21oi_1 _13404_ (.A1(net4946),
    .A2(_04505_),
    .Y(_04823_),
    .B1(net4764));
 sg13g2_o21ai_1 _13405_ (.B1(_04823_),
    .Y(_04824_),
    .A1(_04821_),
    .A2(_04822_));
 sg13g2_o21ai_1 _13406_ (.B1(_04824_),
    .Y(_04825_),
    .A1(net5296),
    .A2(_03312_));
 sg13g2_nor3_1 _13407_ (.A(net5288),
    .B(_04819_),
    .C(_04825_),
    .Y(_04826_));
 sg13g2_o21ai_1 _13408_ (.B1(net5288),
    .Y(_04827_),
    .A1(net5295),
    .A2(_03141_));
 sg13g2_o21ai_1 _13409_ (.B1(net5255),
    .Y(_04828_),
    .A1(_03134_),
    .A2(_04827_));
 sg13g2_o21ai_1 _13410_ (.B1(_04817_),
    .Y(_04829_),
    .A1(_04826_),
    .A2(_04828_));
 sg13g2_o21ai_1 _13411_ (.B1(net5101),
    .Y(_04830_),
    .A1(\m_sys.m_core.m_fsm.r_cstate[1] ),
    .A2(_04829_));
 sg13g2_a22oi_1 _13412_ (.Y(_04831_),
    .B1(net4387),
    .B2(_00124_),
    .A2(net4493),
    .A1(_00050_));
 sg13g2_mux2_1 _13413_ (.A0(_00050_),
    .A1(_00051_),
    .S(net5360),
    .X(_04832_));
 sg13g2_a21oi_1 _13414_ (.A1(net5354),
    .A2(_04211_),
    .Y(_04833_),
    .B1(net5072));
 sg13g2_o21ai_1 _13415_ (.B1(_04833_),
    .Y(_04834_),
    .A1(net5355),
    .A2(_04832_));
 sg13g2_o21ai_1 _13416_ (.B1(_04834_),
    .Y(_04835_),
    .A1(_02497_),
    .A2(net4880));
 sg13g2_a221oi_1 _13417_ (.B2(net5275),
    .C1(_04605_),
    .B1(_04835_),
    .A1(_00123_),
    .Y(_04836_),
    .A2(_04658_));
 sg13g2_o21ai_1 _13418_ (.B1(_04836_),
    .Y(_04837_),
    .A1(net4878),
    .A2(_04831_));
 sg13g2_a22oi_1 _13419_ (.Y(_04838_),
    .B1(_04830_),
    .B2(_04837_),
    .A2(net5094),
    .A1(_02323_));
 sg13g2_nor2b_1 _13420_ (.A(net5326),
    .B_N(\m_sys.m_core.m_gpr._GEN[33] ),
    .Y(_04839_));
 sg13g2_a221oi_1 _13421_ (.B2(\m_sys.m_core.m_gpr._GEN[65] ),
    .C1(_04839_),
    .B1(net5052),
    .A1(\m_sys.m_core.m_gpr._GEN[97] ),
    .Y(_04840_),
    .A2(net5061));
 sg13g2_mux4_1 _13422_ (.S0(net5324),
    .A0(\m_sys.m_core.m_gpr._GEN[129] ),
    .A1(\m_sys.m_core.m_gpr._GEN[161] ),
    .A2(\m_sys.m_core.m_gpr._GEN[193] ),
    .A3(\m_sys.m_core.m_gpr._GEN[225] ),
    .S1(net5326),
    .X(_04841_));
 sg13g2_nor2_1 _13423_ (.A(net5179),
    .B(_04841_),
    .Y(_04842_));
 sg13g2_a21oi_2 _13424_ (.B1(_04842_),
    .Y(_04843_),
    .A2(_04840_),
    .A1(net5179));
 sg13g2_a221oi_1 _13425_ (.B2(net4492),
    .C1(net4959),
    .B1(_04843_),
    .A1(\m_sys.m_core._m_bru_io_o_res[1] ),
    .Y(_04844_),
    .A2(_04456_));
 sg13g2_nor2_1 _13426_ (.A(net4720),
    .B(_04844_),
    .Y(_04845_));
 sg13g2_o21ai_1 _13427_ (.B1(_04845_),
    .Y(_04846_),
    .A1(net4972),
    .A2(_04838_));
 sg13g2_nand2_1 _13428_ (.Y(_00226_),
    .A(_04812_),
    .B(_04846_));
 sg13g2_nor2_1 _13429_ (.A(net5169),
    .B(_03407_),
    .Y(_04847_));
 sg13g2_a22oi_1 _13430_ (.Y(_04848_),
    .B1(net4884),
    .B2(_03403_),
    .A2(_03071_),
    .A1(_03070_));
 sg13g2_a22oi_1 _13431_ (.Y(_04849_),
    .B1(_04848_),
    .B2(_03398_),
    .A2(_03404_),
    .A1(net5083));
 sg13g2_nor3_1 _13432_ (.A(net5172),
    .B(net5301),
    .C(net5255),
    .Y(_04850_));
 sg13g2_xnor2_1 _13433_ (.Y(_04851_),
    .A(_04847_),
    .B(_04849_));
 sg13g2_nand3b_1 _13434_ (.B(_03585_),
    .C(net4924),
    .Y(_04852_),
    .A_N(_03582_));
 sg13g2_nor3_1 _13435_ (.A(net4927),
    .B(_03577_),
    .C(_03583_),
    .Y(_04853_));
 sg13g2_nor2_1 _13436_ (.A(net4885),
    .B(_04853_),
    .Y(_04854_));
 sg13g2_a22oi_1 _13437_ (.Y(_04855_),
    .B1(_04852_),
    .B2(_04854_),
    .A2(_04710_),
    .A1(net4885));
 sg13g2_a21oi_1 _13438_ (.A1(net4949),
    .A2(_04555_),
    .Y(_04856_),
    .B1(net4895));
 sg13g2_o21ai_1 _13439_ (.B1(_04856_),
    .Y(_04857_),
    .A1(net4947),
    .A2(_04855_));
 sg13g2_a21oi_1 _13440_ (.A1(net4895),
    .A2(_04235_),
    .Y(_04858_),
    .B1(_03653_));
 sg13g2_a21oi_1 _13441_ (.A1(_03313_),
    .A2(_03585_),
    .Y(_04859_),
    .B1(net5301));
 sg13g2_a22oi_1 _13442_ (.Y(_04860_),
    .B1(_04857_),
    .B2(_04858_),
    .A2(_03139_),
    .A1(net5288));
 sg13g2_nand2b_1 _13443_ (.Y(_04861_),
    .B(_04860_),
    .A_N(_04859_));
 sg13g2_a21oi_1 _13444_ (.A1(net4765),
    .A2(_04226_),
    .Y(_04862_),
    .B1(_04859_));
 sg13g2_nor2_1 _13445_ (.A(_03443_),
    .B(_04862_),
    .Y(_04863_));
 sg13g2_a221oi_1 _13446_ (.B2(net5256),
    .C1(_04863_),
    .B1(_04861_),
    .A1(_04850_),
    .Y(_04864_),
    .A2(_04851_));
 sg13g2_mux2_1 _13447_ (.A0(_00122_),
    .A1(_00121_),
    .S(_03498_),
    .X(_04865_));
 sg13g2_mux2_1 _13448_ (.A0(_00048_),
    .A1(_04865_),
    .S(_02698_),
    .X(_04866_));
 sg13g2_mux2_1 _13449_ (.A0(_00048_),
    .A1(_00049_),
    .S(net5360),
    .X(_04867_));
 sg13g2_a21oi_1 _13450_ (.A1(net5354),
    .A2(_04244_),
    .Y(_04868_),
    .B1(net5072));
 sg13g2_o21ai_1 _13451_ (.B1(_04868_),
    .Y(_04869_),
    .A1(net5354),
    .A2(_04867_));
 sg13g2_a22oi_1 _13452_ (.Y(_04870_),
    .B1(net4882),
    .B2(_00122_),
    .A2(_03511_),
    .A1(_00121_));
 sg13g2_nand2_1 _13453_ (.Y(_04871_),
    .A(_04869_),
    .B(_04870_));
 sg13g2_a221oi_1 _13454_ (.B2(net5274),
    .C1(_04605_),
    .B1(_04871_),
    .A1(net5069),
    .Y(_04872_),
    .A2(_04866_));
 sg13g2_nor2_1 _13455_ (.A(net5094),
    .B(_04872_),
    .Y(_04873_));
 sg13g2_o21ai_1 _13456_ (.B1(_04873_),
    .Y(_04874_),
    .A1(net5097),
    .A2(_04864_));
 sg13g2_nand2_1 _13457_ (.Y(_04875_),
    .A(_02324_),
    .B(net5096));
 sg13g2_a21oi_1 _13458_ (.A1(_04874_),
    .A2(_04875_),
    .Y(_04876_),
    .B1(net4972));
 sg13g2_nand2b_1 _13459_ (.Y(_04877_),
    .B(net5061),
    .A_N(\m_sys.m_core.m_gpr._GEN[224] ));
 sg13g2_nand2b_1 _13460_ (.Y(_04878_),
    .B(net5148),
    .A_N(\m_sys.m_core.m_gpr._GEN[128] ));
 sg13g2_a22oi_1 _13461_ (.Y(_04879_),
    .B1(net5049),
    .B2(_02485_),
    .A2(net5052),
    .A1(_02486_));
 sg13g2_nand4_1 _13462_ (.B(_04877_),
    .C(_04878_),
    .A(net5327),
    .Y(_04880_),
    .D(_04879_));
 sg13g2_nor2b_1 _13463_ (.A(net5325),
    .B_N(\m_sys.m_core.m_gpr._GEN[32] ),
    .Y(_04881_));
 sg13g2_a221oi_1 _13464_ (.B2(\m_sys.m_core.m_gpr._GEN[64] ),
    .C1(_04881_),
    .B1(net5052),
    .A1(\m_sys.m_core.m_gpr._GEN[96] ),
    .Y(_04882_),
    .A2(net5061));
 sg13g2_o21ai_1 _13465_ (.B1(_04880_),
    .Y(_04883_),
    .A1(net5327),
    .A2(_04882_));
 sg13g2_a221oi_1 _13466_ (.B2(net4492),
    .C1(net4961),
    .B1(_04883_),
    .A1(\m_sys.m_core._m_bru_io_o_res[0] ),
    .Y(_04884_),
    .A2(_04456_));
 sg13g2_or2_1 _13467_ (.X(_04885_),
    .B(_04884_),
    .A(net4720));
 sg13g2_nand2_1 _13468_ (.Y(_04886_),
    .A(net3412),
    .B(net4720));
 sg13g2_o21ai_1 _13469_ (.B1(_04886_),
    .Y(_00227_),
    .A1(_04876_),
    .A2(_04885_));
 sg13g2_nand2b_2 _13470_ (.Y(_04887_),
    .B(\m_sys.m_uart.m_tx.r_cstate[1] ),
    .A_N(net2884));
 sg13g2_inv_1 _13471_ (.Y(_04888_),
    .A(_04887_));
 sg13g2_nand4_1 _13472_ (.B(\m_sys.m_uart.m_tx.r_bit_cnt[1] ),
    .C(\m_sys.m_uart.m_tx.r_bit_cnt[0] ),
    .A(\m_sys.m_uart.m_tx.r_bit_cnt[2] ),
    .Y(_04889_),
    .D(_00014_));
 sg13g2_a21oi_1 _13473_ (.A1(_04888_),
    .A2(_04889_),
    .Y(_04890_),
    .B1(_02526_));
 sg13g2_a21oi_1 _13474_ (.A1(net3206),
    .A2(_04887_),
    .Y(_04891_),
    .B1(_04890_));
 sg13g2_nor2_1 _13475_ (.A(net2884),
    .B(\m_sys.m_uart.m_tx.r_cstate[1] ),
    .Y(_04892_));
 sg13g2_nor2_1 _13476_ (.A(net5282),
    .B(net5283),
    .Y(_04893_));
 sg13g2_inv_1 _13477_ (.Y(_04894_),
    .A(_04893_));
 sg13g2_nor4_2 _13478_ (.A(\m_sys.m_bootloader.r_cstate[1] ),
    .B(net5285),
    .C(_00024_),
    .Y(_04895_),
    .D(_04894_));
 sg13g2_nand2_1 _13479_ (.Y(_04896_),
    .A(\m_sys.m_bootloader.r_cstate[1] ),
    .B(net5285));
 sg13g2_nor3_2 _13480_ (.A(net5283),
    .B(_02361_),
    .C(_02706_),
    .Y(_04897_));
 sg13g2_and2_1 _13481_ (.A(net5282),
    .B(_04897_),
    .X(_04898_));
 sg13g2_nand2_1 _13482_ (.Y(_04899_),
    .A(net5282),
    .B(_04897_));
 sg13g2_o21ai_1 _13483_ (.B1(net5271),
    .Y(_04900_),
    .A1(_04895_),
    .A2(_04898_));
 sg13g2_nand3_1 _13484_ (.B(_02696_),
    .C(_02703_),
    .A(_02693_),
    .Y(_04901_));
 sg13g2_a21oi_2 _13485_ (.B1(net5272),
    .Y(_04902_),
    .A2(_03548_),
    .A1(_02721_));
 sg13g2_a21oi_1 _13486_ (.A1(net5268),
    .A2(_00025_),
    .Y(_04903_),
    .B1(_04902_));
 sg13g2_o21ai_1 _13487_ (.B1(net5234),
    .Y(_04904_),
    .A1(_02676_),
    .A2(_04901_));
 sg13g2_nand2_1 _13488_ (.Y(_04905_),
    .A(_04903_),
    .B(_04904_));
 sg13g2_nand2_1 _13489_ (.Y(_04906_),
    .A(net4663),
    .B(_02669_));
 sg13g2_o21ai_1 _13490_ (.B1(_04900_),
    .Y(_04907_),
    .A1(_04905_),
    .A2(_04906_));
 sg13g2_inv_1 _13491_ (.Y(_04908_),
    .A(_04907_));
 sg13g2_a21oi_1 _13492_ (.A1(net5146),
    .A2(_04908_),
    .Y(_04909_),
    .B1(_04891_));
 sg13g2_nor2_1 _13493_ (.A(\m_sys.m_uart.m_tx.r_cstate[1] ),
    .B(net3206),
    .Y(_04910_));
 sg13g2_nor2b_1 _13494_ (.A(_02526_),
    .B_N(_04910_),
    .Y(_04911_));
 sg13g2_nor2_1 _13495_ (.A(_02526_),
    .B(_04887_),
    .Y(_04912_));
 sg13g2_and2_1 _13496_ (.A(net3302),
    .B(_04912_),
    .X(_04913_));
 sg13g2_and2_1 _13497_ (.A(net3208),
    .B(_04913_),
    .X(_04914_));
 sg13g2_nand2_1 _13498_ (.Y(_04915_),
    .A(net3161),
    .B(_04914_));
 sg13g2_nand2b_1 _13499_ (.Y(_04916_),
    .B(_04915_),
    .A_N(_04911_));
 sg13g2_a22oi_1 _13500_ (.Y(_04917_),
    .B1(_04909_),
    .B2(_04916_),
    .A2(_04891_),
    .A1(net3353));
 sg13g2_nor2_1 _13501_ (.A(net5376),
    .B(_04917_),
    .Y(_00228_));
 sg13g2_o21ai_1 _13502_ (.B1(_04915_),
    .Y(_04918_),
    .A1(_02527_),
    .A2(_04908_));
 sg13g2_a22oi_1 _13503_ (.Y(_04919_),
    .B1(_04909_),
    .B2(_04918_),
    .A2(_04891_),
    .A1(net2884));
 sg13g2_nor2_1 _13504_ (.A(net5376),
    .B(net2885),
    .Y(_00229_));
 sg13g2_nor2_1 _13505_ (.A(net3380),
    .B(_02365_),
    .Y(_04920_));
 sg13g2_nand3_1 _13506_ (.B(\m_sys.m_uart.m_rx.r_bit_cnt[1] ),
    .C(\m_sys.m_uart.m_rx.r_bit_cnt[0] ),
    .A(net2828),
    .Y(_04921_));
 sg13g2_nand2_1 _13507_ (.Y(_04922_),
    .A(net2903),
    .B(net3125));
 sg13g2_nor2_2 _13508_ (.A(net2903),
    .B(\m_sys.m_uart.m_rx.r_cstate[1] ),
    .Y(_04923_));
 sg13g2_nor3_1 _13509_ (.A(net3148),
    .B(_02364_),
    .C(net3408),
    .Y(_04924_));
 sg13g2_nor3_1 _13510_ (.A(_02602_),
    .B(_04920_),
    .C(_04924_),
    .Y(_04925_));
 sg13g2_nor3_1 _13511_ (.A(net5368),
    .B(_02579_),
    .C(_04925_),
    .Y(_00230_));
 sg13g2_a221oi_1 _13512_ (.B2(net3292),
    .C1(_02602_),
    .B1(_04920_),
    .A1(net3148),
    .Y(_04926_),
    .A2(_02365_));
 sg13g2_o21ai_1 _13513_ (.B1(net5379),
    .Y(_04927_),
    .A1(net2903),
    .A2(_04926_));
 sg13g2_a21oi_1 _13514_ (.A1(net2903),
    .A2(net4368),
    .Y(_00231_),
    .B1(_04927_));
 sg13g2_a22oi_1 _13515_ (.Y(_04928_),
    .B1(net5158),
    .B2(_02728_),
    .A2(net5311),
    .A1(net5240));
 sg13g2_nor2b_1 _13516_ (.A(_02681_),
    .B_N(_02677_),
    .Y(_04929_));
 sg13g2_nand2_1 _13517_ (.Y(_04930_),
    .A(_02671_),
    .B(_04929_));
 sg13g2_nor2_2 _13518_ (.A(_02647_),
    .B(net4490),
    .Y(_04931_));
 sg13g2_or2_1 _13519_ (.X(_04932_),
    .B(_02719_),
    .A(net5159));
 sg13g2_nor3_2 _13520_ (.A(_02685_),
    .B(_04902_),
    .C(_04932_),
    .Y(_04933_));
 sg13g2_nand2_1 _13521_ (.Y(_04934_),
    .A(_04931_),
    .B(net4327));
 sg13g2_nand2_1 _13522_ (.Y(_04935_),
    .A(net2400),
    .B(net4307));
 sg13g2_o21ai_1 _13523_ (.B1(_04935_),
    .Y(_00232_),
    .A1(net5045),
    .A2(_04934_));
 sg13g2_a22oi_1 _13524_ (.Y(_04936_),
    .B1(net5158),
    .B2(_02731_),
    .A2(\m_sys._m_core_io_b_mem_wdata[1] ),
    .A1(net5241));
 sg13g2_nand2_1 _13525_ (.Y(_04937_),
    .A(net1844),
    .B(net4306));
 sg13g2_o21ai_1 _13526_ (.B1(_04937_),
    .Y(_00233_),
    .A1(net4306),
    .A2(net4876));
 sg13g2_a22oi_1 _13527_ (.Y(_04938_),
    .B1(net5158),
    .B2(_02734_),
    .A2(\m_sys._m_core_io_b_mem_wdata[2] ),
    .A1(net5240));
 sg13g2_nand2_1 _13528_ (.Y(_04939_),
    .A(net2049),
    .B(net4307));
 sg13g2_o21ai_1 _13529_ (.B1(_04939_),
    .Y(_00234_),
    .A1(net4307),
    .A2(net5035));
 sg13g2_a22oi_1 _13530_ (.Y(_04940_),
    .B1(net5158),
    .B2(_02737_),
    .A2(\m_sys._m_core_io_b_mem_wdata[3] ),
    .A1(net5241));
 sg13g2_nand2_1 _13531_ (.Y(_04941_),
    .A(net2171),
    .B(net4307));
 sg13g2_o21ai_1 _13532_ (.B1(_04941_),
    .Y(_00235_),
    .A1(net4307),
    .A2(net4870));
 sg13g2_a22oi_1 _13533_ (.Y(_04942_),
    .B1(net5158),
    .B2(_02740_),
    .A2(\m_sys._m_core_io_b_mem_wdata[4] ),
    .A1(net5239));
 sg13g2_nand2_1 _13534_ (.Y(_04943_),
    .A(net1889),
    .B(net4306));
 sg13g2_o21ai_1 _13535_ (.B1(_04943_),
    .Y(_00236_),
    .A1(net4306),
    .A2(net5034));
 sg13g2_a22oi_1 _13536_ (.Y(_04944_),
    .B1(net5158),
    .B2(_02743_),
    .A2(\m_sys._m_core_io_b_mem_wdata[5] ),
    .A1(net5239));
 sg13g2_nand2_1 _13537_ (.Y(_04945_),
    .A(net2151),
    .B(net4307));
 sg13g2_o21ai_1 _13538_ (.B1(_04945_),
    .Y(_00237_),
    .A1(net4307),
    .A2(net4865));
 sg13g2_a22oi_1 _13539_ (.Y(_04946_),
    .B1(net5158),
    .B2(_02746_),
    .A2(\m_sys._m_core_io_b_mem_wdata[6] ),
    .A1(net5239));
 sg13g2_nand2_1 _13540_ (.Y(_04947_),
    .A(net1897),
    .B(net4306));
 sg13g2_o21ai_1 _13541_ (.B1(_04947_),
    .Y(_00238_),
    .A1(net4306),
    .A2(net5028));
 sg13g2_a22oi_1 _13542_ (.Y(_04948_),
    .B1(net5158),
    .B2(_02749_),
    .A2(\m_sys._m_core_io_b_mem_wdata[7] ),
    .A1(net5239));
 sg13g2_nand2_1 _13543_ (.Y(_04949_),
    .A(net2555),
    .B(net4306));
 sg13g2_o21ai_1 _13544_ (.B1(_04949_),
    .Y(_00239_),
    .A1(net4306),
    .A2(net4862));
 sg13g2_and2_2 _13545_ (.A(net5266),
    .B(_02723_),
    .X(_04950_));
 sg13g2_nor2b_2 _13546_ (.A(net5273),
    .B_N(\m_sys._m_core_io_b_mem_wdata[8] ),
    .Y(_04951_));
 sg13g2_a21oi_2 _13547_ (.B1(_04951_),
    .Y(_04952_),
    .A2(_04950_),
    .A1(\m_sys._m_bootloader_io_b_mem_wdata[0] ));
 sg13g2_a21oi_2 _13548_ (.B1(net5234),
    .Y(_04953_),
    .A2(\m_sys._m_bootloader_io_b_mem_wen[0] ),
    .A1(net5267));
 sg13g2_and3_1 _13549_ (.X(_04954_),
    .A(_02721_),
    .B(_03548_),
    .C(_04286_));
 sg13g2_nor2_1 _13550_ (.A(net5270),
    .B(_04954_),
    .Y(_04955_));
 sg13g2_nor3_2 _13551_ (.A(_04932_),
    .B(_04953_),
    .C(_04955_),
    .Y(_04956_));
 sg13g2_nand2_1 _13552_ (.Y(_04957_),
    .A(_04931_),
    .B(net4321));
 sg13g2_nand2_1 _13553_ (.Y(_04958_),
    .A(net2052),
    .B(net4305));
 sg13g2_o21ai_1 _13554_ (.B1(_04958_),
    .Y(_00240_),
    .A1(net4853),
    .A2(net4305));
 sg13g2_nor2_2 _13555_ (.A(net5273),
    .B(_02408_),
    .Y(_04959_));
 sg13g2_a21oi_2 _13556_ (.B1(_04959_),
    .Y(_04960_),
    .A2(_04950_),
    .A1(\m_sys._m_bootloader_io_b_mem_wdata[1] ));
 sg13g2_nand2_1 _13557_ (.Y(_04961_),
    .A(net1719),
    .B(net4305));
 sg13g2_o21ai_1 _13558_ (.B1(_04961_),
    .Y(_00241_),
    .A1(net4305),
    .A2(net4847));
 sg13g2_nand2_2 _13559_ (.Y(_04962_),
    .A(net5241),
    .B(net3407));
 sg13g2_a22oi_1 _13560_ (.Y(_04963_),
    .B1(_04950_),
    .B2(\m_sys._m_bootloader_io_b_mem_wdata[2] ),
    .A2(\m_sys._m_core_io_b_mem_wdata[10] ),
    .A1(net5241));
 sg13g2_nand2_1 _13561_ (.Y(_04964_),
    .A(net1902),
    .B(net4305));
 sg13g2_o21ai_1 _13562_ (.B1(_04964_),
    .Y(_00242_),
    .A1(net4305),
    .A2(net4842));
 sg13g2_nor2_2 _13563_ (.A(net5273),
    .B(_02410_),
    .Y(_04965_));
 sg13g2_a21oi_2 _13564_ (.B1(_04965_),
    .Y(_04966_),
    .A2(_04950_),
    .A1(\m_sys._m_bootloader_io_b_mem_wdata[3] ));
 sg13g2_nand2_1 _13565_ (.Y(_04967_),
    .A(net2097),
    .B(net4304));
 sg13g2_o21ai_1 _13566_ (.B1(_04967_),
    .Y(_00243_),
    .A1(net4304),
    .A2(net4838));
 sg13g2_nand2_1 _13567_ (.Y(_04968_),
    .A(net5233),
    .B(net3401));
 sg13g2_a22oi_1 _13568_ (.Y(_04969_),
    .B1(_04950_),
    .B2(\m_sys._m_bootloader_io_b_mem_wdata[4] ),
    .A2(\m_sys._m_core_io_b_mem_wdata[12] ),
    .A1(net5240));
 sg13g2_nand2_1 _13569_ (.Y(_04970_),
    .A(net1737),
    .B(net4304));
 sg13g2_o21ai_1 _13570_ (.B1(_04970_),
    .Y(_00244_),
    .A1(net4304),
    .A2(net4832));
 sg13g2_nor2b_2 _13571_ (.A(net5272),
    .B_N(\m_sys._m_core_io_b_mem_wdata[13] ),
    .Y(_04971_));
 sg13g2_a21oi_2 _13572_ (.B1(_04971_),
    .Y(_04972_),
    .A2(_04950_),
    .A1(\m_sys._m_bootloader_io_b_mem_wdata[5] ));
 sg13g2_nand2_1 _13573_ (.Y(_04973_),
    .A(net1817),
    .B(net4304));
 sg13g2_o21ai_1 _13574_ (.B1(_04973_),
    .Y(_00245_),
    .A1(net4304),
    .A2(net4826));
 sg13g2_nor2b_2 _13575_ (.A(net5272),
    .B_N(net3156),
    .Y(_04974_));
 sg13g2_a21oi_1 _13576_ (.A1(\m_sys._m_bootloader_io_b_mem_wdata[6] ),
    .A2(_04950_),
    .Y(_04975_),
    .B1(_04974_));
 sg13g2_nand2_1 _13577_ (.Y(_04976_),
    .A(net1698),
    .B(net4305));
 sg13g2_o21ai_1 _13578_ (.B1(_04976_),
    .Y(_00246_),
    .A1(net4305),
    .A2(net4821));
 sg13g2_nor2b_2 _13579_ (.A(net5272),
    .B_N(\m_sys._m_core_io_b_mem_wdata[15] ),
    .Y(_04977_));
 sg13g2_a21oi_2 _13580_ (.B1(_04977_),
    .Y(_04978_),
    .A2(_04950_),
    .A1(\m_sys._m_bootloader_io_b_mem_wdata[7] ));
 sg13g2_nand2_1 _13581_ (.Y(_04979_),
    .A(net1704),
    .B(net4304));
 sg13g2_o21ai_1 _13582_ (.B1(_04979_),
    .Y(_00247_),
    .A1(net4304),
    .A2(net4815));
 sg13g2_nor2b_1 _13583_ (.A(net4333),
    .B_N(_04931_),
    .Y(_04980_));
 sg13g2_nor2_1 _13584_ (.A(net2335),
    .B(net4303),
    .Y(_04981_));
 sg13g2_a21oi_1 _13585_ (.A1(net5138),
    .A2(net4303),
    .Y(_00248_),
    .B1(_04981_));
 sg13g2_nor2_1 _13586_ (.A(net2639),
    .B(_04980_),
    .Y(_04982_));
 sg13g2_a21oi_1 _13587_ (.A1(net4996),
    .A2(net4303),
    .Y(_00249_),
    .B1(_04982_));
 sg13g2_nor2_1 _13588_ (.A(net2326),
    .B(net4302),
    .Y(_04983_));
 sg13g2_a21oi_1 _13589_ (.A1(net5132),
    .A2(net4302),
    .Y(_00250_),
    .B1(_04983_));
 sg13g2_nor2_1 _13590_ (.A(net2424),
    .B(net4303),
    .Y(_04984_));
 sg13g2_a21oi_1 _13591_ (.A1(net4991),
    .A2(net4303),
    .Y(_00251_),
    .B1(_04984_));
 sg13g2_nor2_1 _13592_ (.A(net2221),
    .B(net4302),
    .Y(_04985_));
 sg13g2_a21oi_1 _13593_ (.A1(net5126),
    .A2(net4302),
    .Y(_00252_),
    .B1(_04985_));
 sg13g2_nor2_1 _13594_ (.A(net2659),
    .B(net4303),
    .Y(_04986_));
 sg13g2_a21oi_1 _13595_ (.A1(net4987),
    .A2(net4303),
    .Y(_00253_),
    .B1(_04986_));
 sg13g2_nor2_1 _13596_ (.A(net2402),
    .B(net4302),
    .Y(_04987_));
 sg13g2_a21oi_1 _13597_ (.A1(net5121),
    .A2(net4302),
    .Y(_00254_),
    .B1(_04987_));
 sg13g2_nor2_1 _13598_ (.A(net2881),
    .B(net4302),
    .Y(_04988_));
 sg13g2_a21oi_1 _13599_ (.A1(net4980),
    .A2(net4302),
    .Y(_00255_),
    .B1(_04988_));
 sg13g2_nor2_2 _13600_ (.A(_02644_),
    .B(net4487),
    .Y(_04989_));
 sg13g2_nand2_1 _13601_ (.Y(_04990_),
    .A(net4326),
    .B(_04989_));
 sg13g2_nand2_1 _13602_ (.Y(_04991_),
    .A(net2357),
    .B(net4301));
 sg13g2_o21ai_1 _13603_ (.B1(_04991_),
    .Y(_00256_),
    .A1(net5042),
    .A2(_04990_));
 sg13g2_nand2_1 _13604_ (.Y(_04992_),
    .A(net1898),
    .B(net4300));
 sg13g2_o21ai_1 _13605_ (.B1(_04992_),
    .Y(_00257_),
    .A1(net4876),
    .A2(net4300));
 sg13g2_nand2_1 _13606_ (.Y(_04993_),
    .A(net1787),
    .B(net4301));
 sg13g2_o21ai_1 _13607_ (.B1(_04993_),
    .Y(_00258_),
    .A1(net5035),
    .A2(net4301));
 sg13g2_nand2_1 _13608_ (.Y(_04994_),
    .A(net2051),
    .B(net4301));
 sg13g2_o21ai_1 _13609_ (.B1(_04994_),
    .Y(_00259_),
    .A1(net4870),
    .A2(net4301));
 sg13g2_nand2_1 _13610_ (.Y(_04995_),
    .A(net1762),
    .B(net4300));
 sg13g2_o21ai_1 _13611_ (.B1(_04995_),
    .Y(_00260_),
    .A1(net5034),
    .A2(net4300));
 sg13g2_nand2_1 _13612_ (.Y(_04996_),
    .A(net1891),
    .B(net4301));
 sg13g2_o21ai_1 _13613_ (.B1(_04996_),
    .Y(_00261_),
    .A1(net4865),
    .A2(net4301));
 sg13g2_nand2_1 _13614_ (.Y(_04997_),
    .A(net1928),
    .B(net4300));
 sg13g2_o21ai_1 _13615_ (.B1(_04997_),
    .Y(_00262_),
    .A1(net5028),
    .A2(net4300));
 sg13g2_nand2_1 _13616_ (.Y(_04998_),
    .A(net2161),
    .B(net4300));
 sg13g2_o21ai_1 _13617_ (.B1(_04998_),
    .Y(_00263_),
    .A1(net4862),
    .A2(net4300));
 sg13g2_a21oi_1 _13618_ (.A1(_02700_),
    .A2(net4958),
    .Y(_00264_),
    .B1(net5376));
 sg13g2_nand2_1 _13619_ (.Y(_04999_),
    .A(net5353),
    .B(_02475_));
 sg13g2_nand2b_1 _13620_ (.Y(_05000_),
    .B(\m_sys.m_core.m_bru.io_i_s1[30] ),
    .A_N(\m_sys.m_core.m_bru.io_i_s2[30] ));
 sg13g2_a21oi_1 _13621_ (.A1(_04999_),
    .A2(_05000_),
    .Y(_05001_),
    .B1(_03404_));
 sg13g2_a22oi_1 _13622_ (.Y(_05002_),
    .B1(_02477_),
    .B2(\m_sys.m_core.m_bru.io_i_s1[28] ),
    .A2(_02476_),
    .A1(\m_sys.m_core.m_bru.io_i_s1[29] ));
 sg13g2_nor2b_2 _13623_ (.A(_03404_),
    .B_N(_04999_),
    .Y(_05003_));
 sg13g2_nand2_1 _13624_ (.Y(_05004_),
    .A(_02443_),
    .B(\m_sys.m_core.m_bru.io_i_s2[30] ));
 sg13g2_nor2_1 _13625_ (.A(\m_sys.m_core.m_bru.io_i_s1[29] ),
    .B(_02476_),
    .Y(_05005_));
 sg13g2_nand3_1 _13626_ (.B(_05003_),
    .C(_05004_),
    .A(_05000_),
    .Y(_05006_));
 sg13g2_nor3_1 _13627_ (.A(_05002_),
    .B(_05005_),
    .C(_05006_),
    .Y(_05007_));
 sg13g2_o21ai_1 _13628_ (.B1(_05002_),
    .Y(_05008_),
    .A1(\m_sys.m_core.m_bru.io_i_s1[28] ),
    .A2(_02477_));
 sg13g2_or3_2 _13629_ (.A(_05005_),
    .B(_05006_),
    .C(_05008_),
    .X(_05009_));
 sg13g2_a22oi_1 _13630_ (.Y(_05010_),
    .B1(_02479_),
    .B2(\m_sys.m_core.m_bru.io_i_s1[26] ),
    .A2(_02478_),
    .A1(\m_sys.m_core.m_bru.io_i_s1[27] ));
 sg13g2_a22oi_1 _13631_ (.Y(_05011_),
    .B1(\m_sys.m_core.m_bru.io_i_s2[25] ),
    .B2(net5195),
    .A2(\m_sys.m_core.m_bru.io_i_s2[26] ),
    .A1(net5194));
 sg13g2_nand2_1 _13632_ (.Y(_05012_),
    .A(\m_sys.m_core.m_bru.io_i_s1[24] ),
    .B(_02480_));
 sg13g2_o21ai_1 _13633_ (.B1(_05012_),
    .Y(_05013_),
    .A1(net5195),
    .A2(\m_sys.m_core.m_bru.io_i_s2[25] ));
 sg13g2_nor2_1 _13634_ (.A(\m_sys.m_core.m_bru.io_i_s1[24] ),
    .B(_02480_),
    .Y(_05014_));
 sg13g2_a22oi_1 _13635_ (.Y(_05015_),
    .B1(_02482_),
    .B2(net5352),
    .A2(_02481_),
    .A1(\m_sys.m_core.m_bru.io_i_s1[23] ));
 sg13g2_a22oi_1 _13636_ (.Y(_05016_),
    .B1(\m_sys.m_core.m_bru.io_i_s2[21] ),
    .B2(net5218),
    .A2(\m_sys.m_core.m_bru.io_i_s2[22] ),
    .A1(net5208));
 sg13g2_a22oi_1 _13637_ (.Y(_05017_),
    .B1(\m_sys.m_core.m_bru.io_i_s2[19] ),
    .B2(net5176),
    .A2(\m_sys.m_core.m_bru.io_i_s2[20] ),
    .A1(net5199));
 sg13g2_nor2_1 _13638_ (.A(net5176),
    .B(\m_sys.m_core.m_bru.io_i_s2[19] ),
    .Y(_05018_));
 sg13g2_a22oi_1 _13639_ (.Y(_05019_),
    .B1(_02484_),
    .B2(net5327),
    .A2(_02483_),
    .A1(\m_sys.m_core.m_bru.io_i_s1[18] ));
 sg13g2_nand2_1 _13640_ (.Y(_05020_),
    .A(_02448_),
    .B(\m_sys.m_core.m_bru.io_i_s2[17] ));
 sg13g2_nand3b_1 _13641_ (.B(_05020_),
    .C(net5325),
    .Y(_05021_),
    .A_N(\m_sys.m_core.m_bru.io_i_s2[16] ));
 sg13g2_a22oi_1 _13642_ (.Y(_05022_),
    .B1(_05019_),
    .B2(_05021_),
    .A2(\m_sys.m_core.m_bru.io_i_s2[18] ),
    .A1(net5177));
 sg13g2_o21ai_1 _13643_ (.B1(_05017_),
    .Y(_05023_),
    .A1(_05018_),
    .A2(_05022_));
 sg13g2_nand2b_1 _13644_ (.Y(_05024_),
    .B(net5332),
    .A_N(\m_sys.m_core.m_bru.io_i_s2[20] ));
 sg13g2_nand2b_1 _13645_ (.Y(_05025_),
    .B(net5341),
    .A_N(\m_sys.m_core.m_bru.io_i_s2[21] ));
 sg13g2_nand3_1 _13646_ (.B(_05024_),
    .C(_05025_),
    .A(_05023_),
    .Y(_05026_));
 sg13g2_nand2_1 _13647_ (.Y(_05027_),
    .A(_05016_),
    .B(_05026_));
 sg13g2_a221oi_1 _13648_ (.B2(_05027_),
    .C1(_05014_),
    .B1(_05015_),
    .A1(net5197),
    .Y(_05028_),
    .A2(\m_sys.m_core.m_bru.io_i_s2[23] ));
 sg13g2_o21ai_1 _13649_ (.B1(_05011_),
    .Y(_05029_),
    .A1(_05013_),
    .A2(_05028_));
 sg13g2_a22oi_1 _13650_ (.Y(_05030_),
    .B1(\m_sys.m_core.m_bru.io_i_s2[13] ),
    .B2(net5224),
    .A2(\m_sys.m_core.m_bru.io_i_s2[14] ),
    .A1(net5222));
 sg13g2_a22oi_1 _13651_ (.Y(_05031_),
    .B1(_02471_),
    .B2(\m_sys.m_core.m_bru.io_i_s1[11] ),
    .A2(_02470_),
    .A1(net5322));
 sg13g2_a22oi_1 _13652_ (.Y(_05032_),
    .B1(_02468_),
    .B2(\m_sys.m_core.m_bru.io_i_s1[14] ),
    .A2(_02467_),
    .A1(net5324));
 sg13g2_a22oi_1 _13653_ (.Y(_05033_),
    .B1(_02474_),
    .B2(net5320),
    .A2(_02473_),
    .A1(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[2] ));
 sg13g2_nand4_1 _13654_ (.B(_05031_),
    .C(_05032_),
    .A(_05030_),
    .Y(_05034_),
    .D(_05033_));
 sg13g2_nor2_1 _13655_ (.A(net5229),
    .B(\m_sys.m_core.m_bru.io_i_s2[10] ),
    .Y(_05035_));
 sg13g2_nor2_1 _13656_ (.A(net5224),
    .B(\m_sys.m_core.m_bru.io_i_s2[13] ),
    .Y(_05036_));
 sg13g2_nor2_1 _13657_ (.A(net5320),
    .B(_02474_),
    .Y(_05037_));
 sg13g2_nor2_2 _13658_ (.A(net5324),
    .B(_02467_),
    .Y(_05038_));
 sg13g2_nor4_1 _13659_ (.A(_05035_),
    .B(_05036_),
    .C(_05037_),
    .D(_05038_),
    .Y(_05039_));
 sg13g2_a22oi_1 _13660_ (.Y(_05040_),
    .B1(\m_sys.m_core.m_bru.io_i_s2[10] ),
    .B2(net5229),
    .A2(\m_sys.m_core.m_bru.io_i_s2[11] ),
    .A1(net5230));
 sg13g2_nor2_1 _13661_ (.A(net5322),
    .B(_02470_),
    .Y(_05041_));
 sg13g2_nor2_1 _13662_ (.A(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[2] ),
    .B(_02473_),
    .Y(_05042_));
 sg13g2_nor2_1 _13663_ (.A(_05041_),
    .B(_05042_),
    .Y(_05043_));
 sg13g2_nand3_1 _13664_ (.B(_05040_),
    .C(_05043_),
    .A(_05039_),
    .Y(_05044_));
 sg13g2_or2_2 _13665_ (.X(_05045_),
    .B(_05044_),
    .A(_05034_));
 sg13g2_nor2_1 _13666_ (.A(net5227),
    .B(\m_sys.m_core.m_bru.io_i_s2[7] ),
    .Y(_05046_));
 sg13g2_a22oi_1 _13667_ (.Y(_05047_),
    .B1(\m_sys.m_core.m_bru.io_i_s2[6] ),
    .B2(net5226),
    .A2(\m_sys.m_core.m_bru.io_i_s2[7] ),
    .A1(net5227));
 sg13g2_a22oi_1 _13668_ (.Y(_05048_),
    .B1(_02465_),
    .B2(net5318),
    .A2(_02464_),
    .A1(\m_sys.m_core.m_bru.io_i_s1[6] ));
 sg13g2_nand2b_1 _13669_ (.Y(_05049_),
    .B(\m_sys.m_core.m_bru.io_i_s2[4] ),
    .A_N(net5315));
 sg13g2_o21ai_1 _13670_ (.B1(_05049_),
    .Y(_05050_),
    .A1(net5318),
    .A2(_02465_));
 sg13g2_a22oi_1 _13671_ (.Y(_05051_),
    .B1(_02463_),
    .B2(\m_sys.m_core.m_bru.io_i_s1[2] ),
    .A2(_02462_),
    .A1(net5313));
 sg13g2_nor2_1 _13672_ (.A(net5313),
    .B(_02462_),
    .Y(_05052_));
 sg13g2_a21oi_1 _13673_ (.A1(net5231),
    .A2(\m_sys.m_core.m_bru.io_i_s2[2] ),
    .Y(_05053_),
    .B1(_05052_));
 sg13g2_nand2b_1 _13674_ (.Y(_05054_),
    .B(_05051_),
    .A_N(_05052_));
 sg13g2_nand2_1 _13675_ (.Y(_05055_),
    .A(net5312),
    .B(_02461_));
 sg13g2_nand2_1 _13676_ (.Y(_05056_),
    .A(_02397_),
    .B(\m_sys.m_core.m_bru.io_i_s2[0] ));
 sg13g2_nand2b_1 _13677_ (.Y(_05057_),
    .B(\m_sys.m_core.m_bru.io_i_s2[1] ),
    .A_N(net5312));
 sg13g2_nand2_1 _13678_ (.Y(_05058_),
    .A(_05056_),
    .B(_05057_));
 sg13g2_a221oi_1 _13679_ (.B2(_05058_),
    .C1(_05054_),
    .B1(_05055_),
    .A1(net5231),
    .Y(_05059_),
    .A2(\m_sys.m_core.m_bru.io_i_s2[2] ));
 sg13g2_nor2_1 _13680_ (.A(_05051_),
    .B(_05052_),
    .Y(_05060_));
 sg13g2_nor2b_1 _13681_ (.A(\m_sys.m_core.m_bru.io_i_s2[4] ),
    .B_N(net5315),
    .Y(_05061_));
 sg13g2_nor3_1 _13682_ (.A(_05059_),
    .B(_05060_),
    .C(_05061_),
    .Y(_05062_));
 sg13g2_o21ai_1 _13683_ (.B1(_05048_),
    .Y(_05063_),
    .A1(_05050_),
    .A2(_05062_));
 sg13g2_a21oi_2 _13684_ (.B1(_05046_),
    .Y(_05064_),
    .A2(_05063_),
    .A1(_05047_));
 sg13g2_nor2_1 _13685_ (.A(_05033_),
    .B(_05042_),
    .Y(_05065_));
 sg13g2_o21ai_1 _13686_ (.B1(_05040_),
    .Y(_05066_),
    .A1(_05035_),
    .A2(_05065_));
 sg13g2_a21oi_1 _13687_ (.A1(_05031_),
    .A2(_05066_),
    .Y(_05067_),
    .B1(_05041_));
 sg13g2_o21ai_1 _13688_ (.B1(_05030_),
    .Y(_05068_),
    .A1(_05036_),
    .A2(_05067_));
 sg13g2_a21o_1 _13689_ (.A2(_05068_),
    .A1(_05032_),
    .B1(_05038_),
    .X(_05069_));
 sg13g2_o21ai_1 _13690_ (.B1(_05069_),
    .Y(_05070_),
    .A1(_05045_),
    .A2(_05064_));
 sg13g2_nand2_1 _13691_ (.Y(_05071_),
    .A(net5184),
    .B(\m_sys.m_core.m_bru.io_i_s2[16] ));
 sg13g2_nand2b_1 _13692_ (.Y(_05072_),
    .B(_05020_),
    .A_N(_05018_));
 sg13g2_nand3_1 _13693_ (.B(_05015_),
    .C(_05016_),
    .A(_05010_),
    .Y(_05073_));
 sg13g2_a221oi_1 _13694_ (.B2(net5177),
    .C1(_05072_),
    .B1(\m_sys.m_core.m_bru.io_i_s2[18] ),
    .A1(net5197),
    .Y(_05074_),
    .A2(\m_sys.m_core.m_bru.io_i_s2[23] ));
 sg13g2_o21ai_1 _13695_ (.B1(_05025_),
    .Y(_05075_),
    .A1(net5184),
    .A2(\m_sys.m_core.m_bru.io_i_s2[16] ));
 sg13g2_a221oi_1 _13696_ (.B2(net5196),
    .C1(_05075_),
    .B1(\m_sys.m_core.m_bru.io_i_s2[24] ),
    .A1(net5193),
    .Y(_05076_),
    .A2(\m_sys.m_core.m_bru.io_i_s2[27] ));
 sg13g2_and4_1 _13697_ (.A(_05019_),
    .B(_05024_),
    .C(_05071_),
    .D(_05076_),
    .X(_05077_));
 sg13g2_nand4_1 _13698_ (.B(_05017_),
    .C(_05074_),
    .A(_05011_),
    .Y(_05078_),
    .D(_05077_));
 sg13g2_nor4_2 _13699_ (.A(_05009_),
    .B(_05013_),
    .C(_05073_),
    .Y(_05079_),
    .D(_05078_));
 sg13g2_and2_1 _13700_ (.A(_05070_),
    .B(_05079_),
    .X(_05080_));
 sg13g2_a221oi_1 _13701_ (.B2(_05029_),
    .C1(_05009_),
    .B1(_05010_),
    .A1(net5193),
    .Y(_05081_),
    .A2(\m_sys.m_core.m_bru.io_i_s2[27] ));
 sg13g2_or4_2 _13702_ (.A(_05001_),
    .B(_05007_),
    .C(_05080_),
    .D(_05081_),
    .X(_05082_));
 sg13g2_nand2b_1 _13703_ (.Y(_05083_),
    .B(\m_sys.m_core.m_bru.io_i_uop[1] ),
    .A_N(\m_sys.m_core.m_bru.io_i_uop[0] ));
 sg13g2_xor2_1 _13704_ (.B(_05003_),
    .A(_00087_),
    .X(_05084_));
 sg13g2_o21ai_1 _13705_ (.B1(_05083_),
    .Y(_05085_),
    .A1(\m_sys.m_core.m_bru.io_i_uop[1] ),
    .A2(_05084_));
 sg13g2_a21oi_1 _13706_ (.A1(_05082_),
    .A2(_05085_),
    .Y(_05086_),
    .B1(_02459_));
 sg13g2_o21ai_1 _13707_ (.B1(_05086_),
    .Y(_05087_),
    .A1(_05082_),
    .A2(_05085_));
 sg13g2_nand3_1 _13708_ (.B(_05056_),
    .C(_05057_),
    .A(_05047_),
    .Y(_05088_));
 sg13g2_nor2_1 _13709_ (.A(_05050_),
    .B(_05088_),
    .Y(_05089_));
 sg13g2_nand2_1 _13710_ (.Y(_05090_),
    .A(_05048_),
    .B(_05089_));
 sg13g2_o21ai_1 _13711_ (.B1(_05055_),
    .Y(_05091_),
    .A1(_02397_),
    .A2(\m_sys.m_core.m_bru.io_i_s2[0] ));
 sg13g2_nor3_1 _13712_ (.A(_05046_),
    .B(_05061_),
    .C(_05091_),
    .Y(_05092_));
 sg13g2_nand3_1 _13713_ (.B(_05053_),
    .C(_05092_),
    .A(_05051_),
    .Y(_05093_));
 sg13g2_nor3_2 _13714_ (.A(_05045_),
    .B(_05090_),
    .C(_05093_),
    .Y(_05094_));
 sg13g2_a21oi_1 _13715_ (.A1(_05079_),
    .A2(_05094_),
    .Y(_05095_),
    .B1(\m_sys.m_core.m_bru.io_i_uop[1] ));
 sg13g2_xor2_1 _13716_ (.B(_05095_),
    .A(\m_sys.m_core.m_bru.io_i_uop[0] ),
    .X(_05096_));
 sg13g2_o21ai_1 _13717_ (.B1(_05087_),
    .Y(_05097_),
    .A1(\m_sys.m_core.m_bru.io_i_uop[2] ),
    .A2(_05096_));
 sg13g2_nand3_1 _13718_ (.B(net4961),
    .C(_05097_),
    .A(net3365),
    .Y(_05098_));
 sg13g2_a21oi_1 _13719_ (.A1(net5199),
    .A2(_02486_),
    .Y(_05099_),
    .B1(net5220));
 sg13g2_o21ai_1 _13720_ (.B1(_05099_),
    .Y(_05100_),
    .A1(net5199),
    .A2(\m_sys.m_core.m_gpr._GEN[224] ));
 sg13g2_a221oi_1 _13721_ (.B2(\m_sys.m_core.m_gpr._GEN[160] ),
    .C1(net5211),
    .B1(net5113),
    .A1(\m_sys.m_core.m_gpr._GEN[128] ),
    .Y(_05101_),
    .A2(net5153));
 sg13g2_mux2_1 _13722_ (.A0(\m_sys.m_core.m_gpr._GEN[64] ),
    .A1(\m_sys.m_core.m_gpr._GEN[96] ),
    .S(net5334),
    .X(_05102_));
 sg13g2_a22oi_1 _13723_ (.Y(_05103_),
    .B1(_05102_),
    .B2(net5343),
    .A2(net5113),
    .A1(\m_sys.m_core.m_gpr._GEN[32] ));
 sg13g2_a221oi_1 _13724_ (.B2(net5211),
    .C1(net5108),
    .B1(_05103_),
    .A1(_05100_),
    .Y(_05104_),
    .A2(_05101_));
 sg13g2_a21oi_1 _13725_ (.A1(net4733),
    .A2(_05104_),
    .Y(_05105_),
    .B1(net4735));
 sg13g2_a22oi_1 _13726_ (.Y(_00265_),
    .B1(_05098_),
    .B2(_05105_),
    .A2(net4735),
    .A1(net5221));
 sg13g2_nand2_1 _13727_ (.Y(_05106_),
    .A(_02677_),
    .B(_02681_));
 sg13g2_or2_1 _13728_ (.X(_05107_),
    .B(_05106_),
    .A(_02671_));
 sg13g2_nor2_2 _13729_ (.A(_02647_),
    .B(net4482),
    .Y(_05108_));
 sg13g2_nand2_1 _13730_ (.Y(_05109_),
    .A(net4326),
    .B(_05108_));
 sg13g2_nand2_1 _13731_ (.Y(_05110_),
    .A(net1687),
    .B(net4298));
 sg13g2_o21ai_1 _13732_ (.B1(_05110_),
    .Y(_00266_),
    .A1(net5042),
    .A2(net4298));
 sg13g2_nand2_1 _13733_ (.Y(_05111_),
    .A(net2215),
    .B(net4299));
 sg13g2_o21ai_1 _13734_ (.B1(_05111_),
    .Y(_00267_),
    .A1(net4877),
    .A2(net4299));
 sg13g2_nand2_1 _13735_ (.Y(_05112_),
    .A(net1747),
    .B(net4298));
 sg13g2_o21ai_1 _13736_ (.B1(_05112_),
    .Y(_00268_),
    .A1(net5035),
    .A2(net4298));
 sg13g2_nand2_1 _13737_ (.Y(_05113_),
    .A(net2268),
    .B(net4299));
 sg13g2_o21ai_1 _13738_ (.B1(_05113_),
    .Y(_00269_),
    .A1(net4869),
    .A2(net4299));
 sg13g2_nand2_1 _13739_ (.Y(_05114_),
    .A(net2199),
    .B(net4299));
 sg13g2_o21ai_1 _13740_ (.B1(_05114_),
    .Y(_00270_),
    .A1(net5031),
    .A2(net4299));
 sg13g2_nand2_1 _13741_ (.Y(_05115_),
    .A(net1915),
    .B(net4298));
 sg13g2_o21ai_1 _13742_ (.B1(_05115_),
    .Y(_00271_),
    .A1(net4864),
    .A2(net4298));
 sg13g2_nand2_1 _13743_ (.Y(_05116_),
    .A(net1724),
    .B(net4298));
 sg13g2_o21ai_1 _13744_ (.B1(_05116_),
    .Y(_00272_),
    .A1(net5029),
    .A2(net4298));
 sg13g2_nand2_1 _13745_ (.Y(_05117_),
    .A(net2148),
    .B(net4299));
 sg13g2_o21ai_1 _13746_ (.B1(_05117_),
    .Y(_00273_),
    .A1(net4863),
    .A2(net4299));
 sg13g2_nand2_1 _13747_ (.Y(_05118_),
    .A(net4320),
    .B(_05108_));
 sg13g2_nand2_1 _13748_ (.Y(_05119_),
    .A(net2024),
    .B(net4297));
 sg13g2_o21ai_1 _13749_ (.B1(_05119_),
    .Y(_00274_),
    .A1(net4854),
    .A2(net4297));
 sg13g2_nand2_1 _13750_ (.Y(_05120_),
    .A(net1943),
    .B(net4296));
 sg13g2_o21ai_1 _13751_ (.B1(_05120_),
    .Y(_00275_),
    .A1(net4847),
    .A2(net4296));
 sg13g2_nand2_1 _13752_ (.Y(_05121_),
    .A(net2084),
    .B(net4297));
 sg13g2_o21ai_1 _13753_ (.B1(_05121_),
    .Y(_00276_),
    .A1(net4843),
    .A2(net4297));
 sg13g2_nand2_1 _13754_ (.Y(_05122_),
    .A(net1852),
    .B(_05118_));
 sg13g2_o21ai_1 _13755_ (.B1(_05122_),
    .Y(_00277_),
    .A1(net4837),
    .A2(net4297));
 sg13g2_nand2_1 _13756_ (.Y(_05123_),
    .A(net2004),
    .B(net4296));
 sg13g2_o21ai_1 _13757_ (.B1(_05123_),
    .Y(_00278_),
    .A1(net4831),
    .A2(net4296));
 sg13g2_nand2_1 _13758_ (.Y(_05124_),
    .A(net1836),
    .B(net4297));
 sg13g2_o21ai_1 _13759_ (.B1(_05124_),
    .Y(_00279_),
    .A1(net4825),
    .A2(net4297));
 sg13g2_nand2_1 _13760_ (.Y(_05125_),
    .A(net1696),
    .B(net4296));
 sg13g2_o21ai_1 _13761_ (.B1(_05125_),
    .Y(_00280_),
    .A1(net4821),
    .A2(net4296));
 sg13g2_nand2_1 _13762_ (.Y(_05126_),
    .A(net2138),
    .B(net4296));
 sg13g2_o21ai_1 _13763_ (.B1(_05126_),
    .Y(_00281_),
    .A1(net4816),
    .A2(net4296));
 sg13g2_nand2b_2 _13764_ (.Y(_05127_),
    .B(_02724_),
    .A_N(_04953_));
 sg13g2_nor3_1 _13765_ (.A(net4597),
    .B(net4481),
    .C(net4317),
    .Y(_05128_));
 sg13g2_nor2_1 _13766_ (.A(net2915),
    .B(net4293),
    .Y(_05129_));
 sg13g2_and2_1 _13767_ (.A(net5270),
    .B(\m_sys._m_bootloader_io_b_mem_wdata[0] ),
    .X(_05130_));
 sg13g2_and2_1 _13768_ (.A(\m_sys._m_bootloader_io_b_mem_addr[1] ),
    .B(net5267),
    .X(_05131_));
 sg13g2_a22oi_1 _13769_ (.Y(_05132_),
    .B1(_05130_),
    .B2(net5143),
    .A2(\m_sys._m_core_io_b_mem_wdata[24] ),
    .A1(net5233));
 sg13g2_a21oi_1 _13770_ (.A1(net4293),
    .A2(net5025),
    .Y(_00282_),
    .B1(_05129_));
 sg13g2_nor2_1 _13771_ (.A(net2840),
    .B(net4293),
    .Y(_05133_));
 sg13g2_nor2_1 _13772_ (.A(net5237),
    .B(_02404_),
    .Y(_05134_));
 sg13g2_a22oi_1 _13773_ (.Y(_05135_),
    .B1(net5144),
    .B2(_05134_),
    .A2(\m_sys._m_core_io_b_mem_wdata[25] ),
    .A1(net5237));
 sg13g2_a21oi_1 _13774_ (.A1(net4293),
    .A2(net4811),
    .Y(_00283_),
    .B1(_05133_));
 sg13g2_nor2_1 _13775_ (.A(net2618),
    .B(net4295),
    .Y(_05136_));
 sg13g2_and2_1 _13776_ (.A(net5270),
    .B(\m_sys._m_bootloader_io_b_mem_wdata[2] ),
    .X(_05137_));
 sg13g2_a22oi_1 _13777_ (.Y(_05138_),
    .B1(net5143),
    .B2(_05137_),
    .A2(\m_sys._m_core_io_b_mem_wdata[26] ),
    .A1(net5233));
 sg13g2_a21oi_1 _13778_ (.A1(net4295),
    .A2(net5019),
    .Y(_00284_),
    .B1(_05136_));
 sg13g2_nor2_1 _13779_ (.A(net2661),
    .B(net4295),
    .Y(_05139_));
 sg13g2_nor2_1 _13780_ (.A(net5237),
    .B(_02405_),
    .Y(_05140_));
 sg13g2_a22oi_1 _13781_ (.Y(_05141_),
    .B1(net5144),
    .B2(_05140_),
    .A2(\m_sys._m_core_io_b_mem_wdata[27] ),
    .A1(net5237));
 sg13g2_a21oi_1 _13782_ (.A1(net4295),
    .A2(net4808),
    .Y(_00285_),
    .B1(_05139_));
 sg13g2_nor2_1 _13783_ (.A(net2671),
    .B(net4293),
    .Y(_05142_));
 sg13g2_and2_1 _13784_ (.A(net5270),
    .B(\m_sys._m_bootloader_io_b_mem_wdata[4] ),
    .X(_05143_));
 sg13g2_a22oi_1 _13785_ (.Y(_05144_),
    .B1(net5143),
    .B2(_05143_),
    .A2(\m_sys._m_core_io_b_mem_wdata[28] ),
    .A1(net5233));
 sg13g2_a21oi_1 _13786_ (.A1(net4293),
    .A2(net5011),
    .Y(_00286_),
    .B1(_05142_));
 sg13g2_nor2_1 _13787_ (.A(net2865),
    .B(net4294),
    .Y(_05145_));
 sg13g2_nor2_1 _13788_ (.A(net5238),
    .B(_02406_),
    .Y(_05146_));
 sg13g2_a22oi_1 _13789_ (.Y(_05147_),
    .B1(net5144),
    .B2(_05146_),
    .A2(\m_sys._m_core_io_b_mem_wdata[29] ),
    .A1(net5237));
 sg13g2_a21oi_1 _13790_ (.A1(net4294),
    .A2(net4801),
    .Y(_00287_),
    .B1(_05145_));
 sg13g2_nor2_1 _13791_ (.A(net2358),
    .B(net4293),
    .Y(_05148_));
 sg13g2_and2_1 _13792_ (.A(net5271),
    .B(\m_sys._m_bootloader_io_b_mem_wdata[6] ),
    .X(_05149_));
 sg13g2_a22oi_1 _13793_ (.Y(_05150_),
    .B1(net5143),
    .B2(_05149_),
    .A2(\m_sys._m_core_io_b_mem_wdata[30] ),
    .A1(net5233));
 sg13g2_a21oi_1 _13794_ (.A1(net4293),
    .A2(net5005),
    .Y(_00288_),
    .B1(_05148_));
 sg13g2_nor2_1 _13795_ (.A(net2638),
    .B(net4294),
    .Y(_05151_));
 sg13g2_nor2_1 _13796_ (.A(net5238),
    .B(_02407_),
    .Y(_05152_));
 sg13g2_a22oi_1 _13797_ (.Y(_05153_),
    .B1(net5144),
    .B2(_05152_),
    .A2(\m_sys._m_core_io_b_mem_wdata[31] ),
    .A1(net5237));
 sg13g2_a21oi_1 _13798_ (.A1(net4294),
    .A2(net4798),
    .Y(_00289_),
    .B1(_05151_));
 sg13g2_nand2_1 _13799_ (.Y(_05154_),
    .A(_02670_),
    .B(_04929_));
 sg13g2_nor2_2 _13800_ (.A(net4551),
    .B(net4475),
    .Y(_05155_));
 sg13g2_nand2_1 _13801_ (.Y(_05156_),
    .A(net4330),
    .B(_05155_));
 sg13g2_nand2_1 _13802_ (.Y(_05157_),
    .A(net1998),
    .B(net4291));
 sg13g2_o21ai_1 _13803_ (.B1(_05157_),
    .Y(_00290_),
    .A1(net5041),
    .A2(net4291));
 sg13g2_nand2_1 _13804_ (.Y(_05158_),
    .A(net2076),
    .B(net4292));
 sg13g2_o21ai_1 _13805_ (.B1(_05158_),
    .Y(_00291_),
    .A1(net4876),
    .A2(net4292));
 sg13g2_nand2_1 _13806_ (.Y(_05159_),
    .A(net2430),
    .B(net4291));
 sg13g2_o21ai_1 _13807_ (.B1(_05159_),
    .Y(_00292_),
    .A1(net5037),
    .A2(net4291));
 sg13g2_nand2_1 _13808_ (.Y(_05160_),
    .A(net1778),
    .B(net4292));
 sg13g2_o21ai_1 _13809_ (.B1(_05160_),
    .Y(_00293_),
    .A1(net4873),
    .A2(net4292));
 sg13g2_nand2_1 _13810_ (.Y(_05161_),
    .A(net1811),
    .B(net4291));
 sg13g2_o21ai_1 _13811_ (.B1(_05161_),
    .Y(_00294_),
    .A1(net5030),
    .A2(net4291));
 sg13g2_nand2_1 _13812_ (.Y(_05162_),
    .A(net1796),
    .B(net4291));
 sg13g2_o21ai_1 _13813_ (.B1(_05162_),
    .Y(_00295_),
    .A1(net4865),
    .A2(net4291));
 sg13g2_nand2_1 _13814_ (.Y(_05163_),
    .A(net2065),
    .B(net4292));
 sg13g2_o21ai_1 _13815_ (.B1(_05163_),
    .Y(_00296_),
    .A1(net5028),
    .A2(net4292));
 sg13g2_nand2_1 _13816_ (.Y(_05164_),
    .A(net1918),
    .B(net4292));
 sg13g2_o21ai_1 _13817_ (.B1(_05164_),
    .Y(_00297_),
    .A1(net4862),
    .A2(net4292));
 sg13g2_nand2_1 _13818_ (.Y(_05165_),
    .A(net4325),
    .B(_05155_));
 sg13g2_nand2_1 _13819_ (.Y(_05166_),
    .A(net1812),
    .B(net4290));
 sg13g2_o21ai_1 _13820_ (.B1(_05166_),
    .Y(_00298_),
    .A1(net4858),
    .A2(net4290));
 sg13g2_nand2_1 _13821_ (.Y(_05167_),
    .A(net2220),
    .B(net4289));
 sg13g2_o21ai_1 _13822_ (.B1(_05167_),
    .Y(_00299_),
    .A1(net4851),
    .A2(net4289));
 sg13g2_nand2_1 _13823_ (.Y(_05168_),
    .A(net2192),
    .B(net4290));
 sg13g2_o21ai_1 _13824_ (.B1(_05168_),
    .Y(_00300_),
    .A1(net4845),
    .A2(_05165_));
 sg13g2_nand2_1 _13825_ (.Y(_05169_),
    .A(net2026),
    .B(net4289));
 sg13g2_o21ai_1 _13826_ (.B1(_05169_),
    .Y(_00301_),
    .A1(net4839),
    .A2(net4289));
 sg13g2_nand2_1 _13827_ (.Y(_05170_),
    .A(net1953),
    .B(net4290));
 sg13g2_o21ai_1 _13828_ (.B1(_05170_),
    .Y(_00302_),
    .A1(net4833),
    .A2(net4290));
 sg13g2_nand2_1 _13829_ (.Y(_05171_),
    .A(net1839),
    .B(net4289));
 sg13g2_o21ai_1 _13830_ (.B1(_05171_),
    .Y(_00303_),
    .A1(net4829),
    .A2(net4289));
 sg13g2_nand2_1 _13831_ (.Y(_05172_),
    .A(net2067),
    .B(net4290));
 sg13g2_o21ai_1 _13832_ (.B1(_05172_),
    .Y(_00304_),
    .A1(net4820),
    .A2(net4290));
 sg13g2_nand2_1 _13833_ (.Y(_05173_),
    .A(net1985),
    .B(net4289));
 sg13g2_o21ai_1 _13834_ (.B1(_05173_),
    .Y(_00305_),
    .A1(net4819),
    .A2(net4289));
 sg13g2_nor2b_1 _13835_ (.A(net4331),
    .B_N(_05155_),
    .Y(_05174_));
 sg13g2_nor2_1 _13836_ (.A(net2876),
    .B(net4288),
    .Y(_05175_));
 sg13g2_a21oi_1 _13837_ (.A1(net5135),
    .A2(net4288),
    .Y(_00306_),
    .B1(_05175_));
 sg13g2_nor2_1 _13838_ (.A(net2574),
    .B(net4288),
    .Y(_05176_));
 sg13g2_a21oi_1 _13839_ (.A1(net4993),
    .A2(net4288),
    .Y(_00307_),
    .B1(_05176_));
 sg13g2_nor2_1 _13840_ (.A(net2476),
    .B(net4287),
    .Y(_05177_));
 sg13g2_a21oi_1 _13841_ (.A1(net5130),
    .A2(net4287),
    .Y(_00308_),
    .B1(_05177_));
 sg13g2_nor2_1 _13842_ (.A(net2345),
    .B(net4288),
    .Y(_05178_));
 sg13g2_a21oi_1 _13843_ (.A1(net4988),
    .A2(net4288),
    .Y(_00309_),
    .B1(_05178_));
 sg13g2_nor2_1 _13844_ (.A(net2405),
    .B(net4287),
    .Y(_05179_));
 sg13g2_a21oi_1 _13845_ (.A1(net5127),
    .A2(net4287),
    .Y(_00310_),
    .B1(_05179_));
 sg13g2_nor2_1 _13846_ (.A(net2325),
    .B(net4288),
    .Y(_05180_));
 sg13g2_a21oi_1 _13847_ (.A1(net4983),
    .A2(net4288),
    .Y(_00311_),
    .B1(_05180_));
 sg13g2_nor2_1 _13848_ (.A(net2731),
    .B(net4287),
    .Y(_05181_));
 sg13g2_a21oi_1 _13849_ (.A1(net5121),
    .A2(net4287),
    .Y(_00312_),
    .B1(_05181_));
 sg13g2_nor2_1 _13850_ (.A(net2579),
    .B(net4287),
    .Y(_05182_));
 sg13g2_a21oi_1 _13851_ (.A1(net4978),
    .A2(net4287),
    .Y(_00313_),
    .B1(_05182_));
 sg13g2_nor2_2 _13852_ (.A(_02675_),
    .B(net4479),
    .Y(_05183_));
 sg13g2_nand2_1 _13853_ (.Y(_05184_),
    .A(net4330),
    .B(_05183_));
 sg13g2_nand2_1 _13854_ (.Y(_05185_),
    .A(net1788),
    .B(net4286));
 sg13g2_o21ai_1 _13855_ (.B1(_05185_),
    .Y(_00314_),
    .A1(net5041),
    .A2(net4286));
 sg13g2_nand2_1 _13856_ (.Y(_05186_),
    .A(net1829),
    .B(net4285));
 sg13g2_o21ai_1 _13857_ (.B1(_05186_),
    .Y(_00315_),
    .A1(net4876),
    .A2(net4285));
 sg13g2_nand2_1 _13858_ (.Y(_05187_),
    .A(net2118),
    .B(net4286));
 sg13g2_o21ai_1 _13859_ (.B1(_05187_),
    .Y(_00316_),
    .A1(net5037),
    .A2(net4286));
 sg13g2_nand2_1 _13860_ (.Y(_05188_),
    .A(net2126),
    .B(net4285));
 sg13g2_o21ai_1 _13861_ (.B1(_05188_),
    .Y(_00317_),
    .A1(net4873),
    .A2(net4285));
 sg13g2_nand2_1 _13862_ (.Y(_05189_),
    .A(net2113),
    .B(net4285));
 sg13g2_o21ai_1 _13863_ (.B1(_05189_),
    .Y(_00318_),
    .A1(net5034),
    .A2(net4285));
 sg13g2_nand2_1 _13864_ (.Y(_05190_),
    .A(net2129),
    .B(net4286));
 sg13g2_o21ai_1 _13865_ (.B1(_05190_),
    .Y(_00319_),
    .A1(net4865),
    .A2(net4286));
 sg13g2_nand2_1 _13866_ (.Y(_05191_),
    .A(net2047),
    .B(net4286));
 sg13g2_o21ai_1 _13867_ (.B1(_05191_),
    .Y(_00320_),
    .A1(net5028),
    .A2(_05184_));
 sg13g2_nand2_1 _13868_ (.Y(_05192_),
    .A(net2231),
    .B(net4285));
 sg13g2_o21ai_1 _13869_ (.B1(_05192_),
    .Y(_00321_),
    .A1(net4862),
    .A2(net4285));
 sg13g2_nand2_1 _13870_ (.Y(_05193_),
    .A(net4325),
    .B(_05183_));
 sg13g2_nand2_1 _13871_ (.Y(_05194_),
    .A(net2081),
    .B(net4284));
 sg13g2_o21ai_1 _13872_ (.B1(_05194_),
    .Y(_00322_),
    .A1(net4855),
    .A2(net4284));
 sg13g2_nand2_1 _13873_ (.Y(_05195_),
    .A(net2107),
    .B(net4283));
 sg13g2_o21ai_1 _13874_ (.B1(_05195_),
    .Y(_00323_),
    .A1(net4851),
    .A2(net4283));
 sg13g2_nand2_1 _13875_ (.Y(_05196_),
    .A(net2119),
    .B(net4283));
 sg13g2_o21ai_1 _13876_ (.B1(_05196_),
    .Y(_00324_),
    .A1(net4845),
    .A2(net4283));
 sg13g2_nand2_1 _13877_ (.Y(_05197_),
    .A(net2092),
    .B(net4283));
 sg13g2_o21ai_1 _13878_ (.B1(_05197_),
    .Y(_00325_),
    .A1(net4841),
    .A2(net4283));
 sg13g2_nand2_1 _13879_ (.Y(_05198_),
    .A(net2168),
    .B(net4284));
 sg13g2_o21ai_1 _13880_ (.B1(_05198_),
    .Y(_00326_),
    .A1(net4833),
    .A2(net4284));
 sg13g2_nand2_1 _13881_ (.Y(_05199_),
    .A(net2036),
    .B(net4283));
 sg13g2_o21ai_1 _13882_ (.B1(_05199_),
    .Y(_00327_),
    .A1(net4829),
    .A2(net4283));
 sg13g2_nand2_1 _13883_ (.Y(_05200_),
    .A(net2106),
    .B(net4284));
 sg13g2_o21ai_1 _13884_ (.B1(_05200_),
    .Y(_00328_),
    .A1(net4820),
    .A2(net4284));
 sg13g2_nand2_1 _13885_ (.Y(_05201_),
    .A(net1905),
    .B(net4284));
 sg13g2_o21ai_1 _13886_ (.B1(_05201_),
    .Y(_00329_),
    .A1(net4819),
    .A2(_05193_));
 sg13g2_nor2b_1 _13887_ (.A(net4331),
    .B_N(_05183_),
    .Y(_05202_));
 sg13g2_nor2_1 _13888_ (.A(net2368),
    .B(net4282),
    .Y(_05203_));
 sg13g2_a21oi_1 _13889_ (.A1(net5135),
    .A2(net4282),
    .Y(_00330_),
    .B1(_05203_));
 sg13g2_nor2_1 _13890_ (.A(net2566),
    .B(net4282),
    .Y(_05204_));
 sg13g2_a21oi_1 _13891_ (.A1(net4993),
    .A2(net4282),
    .Y(_00331_),
    .B1(_05204_));
 sg13g2_nor2_1 _13892_ (.A(net2218),
    .B(net4281),
    .Y(_05205_));
 sg13g2_a21oi_1 _13893_ (.A1(net5130),
    .A2(net4281),
    .Y(_00332_),
    .B1(_05205_));
 sg13g2_nor2_1 _13894_ (.A(net2485),
    .B(net4282),
    .Y(_05206_));
 sg13g2_a21oi_1 _13895_ (.A1(net4988),
    .A2(net4282),
    .Y(_00333_),
    .B1(_05206_));
 sg13g2_nor2_1 _13896_ (.A(net2376),
    .B(net4281),
    .Y(_05207_));
 sg13g2_a21oi_1 _13897_ (.A1(net5127),
    .A2(net4281),
    .Y(_00334_),
    .B1(_05207_));
 sg13g2_nor2_1 _13898_ (.A(net2657),
    .B(net4282),
    .Y(_05208_));
 sg13g2_a21oi_1 _13899_ (.A1(net4983),
    .A2(net4282),
    .Y(_00335_),
    .B1(_05208_));
 sg13g2_nor2_1 _13900_ (.A(net2532),
    .B(net4281),
    .Y(_05209_));
 sg13g2_a21oi_1 _13901_ (.A1(net5121),
    .A2(net4281),
    .Y(_00336_),
    .B1(_05209_));
 sg13g2_nor2_1 _13902_ (.A(net2481),
    .B(net4281),
    .Y(_05210_));
 sg13g2_a21oi_1 _13903_ (.A1(net4978),
    .A2(net4281),
    .Y(_00337_),
    .B1(_05210_));
 sg13g2_nand2_1 _13904_ (.Y(_05211_),
    .A(net4321),
    .B(_04989_));
 sg13g2_nand2_1 _13905_ (.Y(_05212_),
    .A(net2040),
    .B(net4280));
 sg13g2_o21ai_1 _13906_ (.B1(_05212_),
    .Y(_00338_),
    .A1(net4853),
    .A2(net4280));
 sg13g2_nand2_1 _13907_ (.Y(_05213_),
    .A(net1859),
    .B(net4280));
 sg13g2_o21ai_1 _13908_ (.B1(_05213_),
    .Y(_00339_),
    .A1(net4847),
    .A2(net4280));
 sg13g2_nand2_1 _13909_ (.Y(_05214_),
    .A(net1910),
    .B(net4280));
 sg13g2_o21ai_1 _13910_ (.B1(_05214_),
    .Y(_00340_),
    .A1(net4842),
    .A2(net4280));
 sg13g2_nand2_1 _13911_ (.Y(_05215_),
    .A(net2074),
    .B(net4279));
 sg13g2_o21ai_1 _13912_ (.B1(_05215_),
    .Y(_00341_),
    .A1(net4838),
    .A2(net4279));
 sg13g2_nand2_1 _13913_ (.Y(_05216_),
    .A(net1984),
    .B(net4279));
 sg13g2_o21ai_1 _13914_ (.B1(_05216_),
    .Y(_00342_),
    .A1(net4831),
    .A2(net4279));
 sg13g2_nand2_1 _13915_ (.Y(_05217_),
    .A(net2053),
    .B(net4279));
 sg13g2_o21ai_1 _13916_ (.B1(_05217_),
    .Y(_00343_),
    .A1(net4826),
    .A2(net4279));
 sg13g2_nand2_1 _13917_ (.Y(_05218_),
    .A(net2042),
    .B(net4280));
 sg13g2_o21ai_1 _13918_ (.B1(_05218_),
    .Y(_00344_),
    .A1(net4824),
    .A2(net4280));
 sg13g2_nand2_1 _13919_ (.Y(_05219_),
    .A(net2103),
    .B(net4279));
 sg13g2_o21ai_1 _13920_ (.B1(_05219_),
    .Y(_00345_),
    .A1(net4816),
    .A2(net4279));
 sg13g2_nor2b_1 _13921_ (.A(net4332),
    .B_N(_04989_),
    .Y(_05220_));
 sg13g2_nor2_1 _13922_ (.A(net2149),
    .B(net4278),
    .Y(_05221_));
 sg13g2_a21oi_1 _13923_ (.A1(net5138),
    .A2(net4278),
    .Y(_00346_),
    .B1(_05221_));
 sg13g2_nor2_1 _13924_ (.A(net2369),
    .B(_05220_),
    .Y(_05222_));
 sg13g2_a21oi_1 _13925_ (.A1(net4995),
    .A2(net4278),
    .Y(_00347_),
    .B1(_05222_));
 sg13g2_nor2_1 _13926_ (.A(net2346),
    .B(net4277),
    .Y(_05223_));
 sg13g2_a21oi_1 _13927_ (.A1(net5132),
    .A2(net4277),
    .Y(_00348_),
    .B1(_05223_));
 sg13g2_nor2_1 _13928_ (.A(net2758),
    .B(net4278),
    .Y(_05224_));
 sg13g2_a21oi_1 _13929_ (.A1(net4991),
    .A2(net4278),
    .Y(_00349_),
    .B1(_05224_));
 sg13g2_nor2_1 _13930_ (.A(net2289),
    .B(net4277),
    .Y(_05225_));
 sg13g2_a21oi_1 _13931_ (.A1(net5125),
    .A2(net4277),
    .Y(_00350_),
    .B1(_05225_));
 sg13g2_nor2_1 _13932_ (.A(net2678),
    .B(net4278),
    .Y(_05226_));
 sg13g2_a21oi_1 _13933_ (.A1(net4986),
    .A2(net4278),
    .Y(_00351_),
    .B1(_05226_));
 sg13g2_nor2_1 _13934_ (.A(net2625),
    .B(net4277),
    .Y(_05227_));
 sg13g2_a21oi_1 _13935_ (.A1(net5120),
    .A2(net4277),
    .Y(_00352_),
    .B1(_05227_));
 sg13g2_nor2_1 _13936_ (.A(net2349),
    .B(net4277),
    .Y(_05228_));
 sg13g2_a21oi_1 _13937_ (.A1(net4980),
    .A2(net4277),
    .Y(_00353_),
    .B1(_05228_));
 sg13g2_nor2_2 _13938_ (.A(_02650_),
    .B(net4487),
    .Y(_05229_));
 sg13g2_nand2_1 _13939_ (.Y(_05230_),
    .A(net4327),
    .B(_05229_));
 sg13g2_nand2_1 _13940_ (.Y(_05231_),
    .A(net1834),
    .B(net4275));
 sg13g2_o21ai_1 _13941_ (.B1(_05231_),
    .Y(_00354_),
    .A1(net5042),
    .A2(net4275));
 sg13g2_nand2_1 _13942_ (.Y(_05232_),
    .A(net2100),
    .B(net4275));
 sg13g2_o21ai_1 _13943_ (.B1(_05232_),
    .Y(_00355_),
    .A1(net4876),
    .A2(net4275));
 sg13g2_nand2_1 _13944_ (.Y(_05233_),
    .A(net2088),
    .B(net4276));
 sg13g2_o21ai_1 _13945_ (.B1(_05233_),
    .Y(_00356_),
    .A1(net5035),
    .A2(net4276));
 sg13g2_nand2_1 _13946_ (.Y(_05234_),
    .A(net2175),
    .B(net4276));
 sg13g2_o21ai_1 _13947_ (.B1(_05234_),
    .Y(_00357_),
    .A1(net4870),
    .A2(net4276));
 sg13g2_nand2_1 _13948_ (.Y(_05235_),
    .A(net2214),
    .B(net4275));
 sg13g2_o21ai_1 _13949_ (.B1(_05235_),
    .Y(_00358_),
    .A1(net5034),
    .A2(net4275));
 sg13g2_nand2_1 _13950_ (.Y(_05236_),
    .A(net2140),
    .B(net4276));
 sg13g2_o21ai_1 _13951_ (.B1(_05236_),
    .Y(_00359_),
    .A1(net4865),
    .A2(net4276));
 sg13g2_nand2_1 _13952_ (.Y(_05237_),
    .A(net1901),
    .B(net4276));
 sg13g2_o21ai_1 _13953_ (.B1(_05237_),
    .Y(_00360_),
    .A1(net5028),
    .A2(_05230_));
 sg13g2_nand2_1 _13954_ (.Y(_05238_),
    .A(net2054),
    .B(net4275));
 sg13g2_o21ai_1 _13955_ (.B1(_05238_),
    .Y(_00361_),
    .A1(net4862),
    .A2(net4275));
 sg13g2_nand2_1 _13956_ (.Y(_05239_),
    .A(net4321),
    .B(_05229_));
 sg13g2_nand2_1 _13957_ (.Y(_05240_),
    .A(net1825),
    .B(net4273));
 sg13g2_o21ai_1 _13958_ (.B1(_05240_),
    .Y(_00362_),
    .A1(net4853),
    .A2(net4273));
 sg13g2_nand2_1 _13959_ (.Y(_05241_),
    .A(net1820),
    .B(net4274));
 sg13g2_o21ai_1 _13960_ (.B1(_05241_),
    .Y(_00363_),
    .A1(net4847),
    .A2(net4274));
 sg13g2_nand2_1 _13961_ (.Y(_05242_),
    .A(net2006),
    .B(net4273));
 sg13g2_o21ai_1 _13962_ (.B1(_05242_),
    .Y(_00364_),
    .A1(net4842),
    .A2(net4273));
 sg13g2_nand2_1 _13963_ (.Y(_05243_),
    .A(net1726),
    .B(net4273));
 sg13g2_o21ai_1 _13964_ (.B1(_05243_),
    .Y(_00365_),
    .A1(net4838),
    .A2(net4273));
 sg13g2_nand2_1 _13965_ (.Y(_05244_),
    .A(net2015),
    .B(net4273));
 sg13g2_o21ai_1 _13966_ (.B1(_05244_),
    .Y(_00366_),
    .A1(net4831),
    .A2(net4273));
 sg13g2_nand2_1 _13967_ (.Y(_05245_),
    .A(net1711),
    .B(net4274));
 sg13g2_o21ai_1 _13968_ (.B1(_05245_),
    .Y(_00367_),
    .A1(net4826),
    .A2(net4274));
 sg13g2_nand2_1 _13969_ (.Y(_05246_),
    .A(net1764),
    .B(net4274));
 sg13g2_o21ai_1 _13970_ (.B1(_05246_),
    .Y(_00368_),
    .A1(net4820),
    .A2(net4274));
 sg13g2_nand2_1 _13971_ (.Y(_05247_),
    .A(net1994),
    .B(net4274));
 sg13g2_o21ai_1 _13972_ (.B1(_05247_),
    .Y(_00369_),
    .A1(net4816),
    .A2(net4274));
 sg13g2_nor2b_1 _13973_ (.A(net4335),
    .B_N(_05229_),
    .Y(_05248_));
 sg13g2_nor2_1 _13974_ (.A(net2433),
    .B(net4272),
    .Y(_05249_));
 sg13g2_a21oi_1 _13975_ (.A1(net5138),
    .A2(net4272),
    .Y(_00370_),
    .B1(_05249_));
 sg13g2_nor2_1 _13976_ (.A(net2291),
    .B(net4272),
    .Y(_05250_));
 sg13g2_a21oi_1 _13977_ (.A1(net4994),
    .A2(net4272),
    .Y(_00371_),
    .B1(_05250_));
 sg13g2_nor2_1 _13978_ (.A(net2819),
    .B(net4271),
    .Y(_05251_));
 sg13g2_a21oi_1 _13979_ (.A1(net5132),
    .A2(net4271),
    .Y(_00372_),
    .B1(_05251_));
 sg13g2_nor2_1 _13980_ (.A(net2388),
    .B(net4272),
    .Y(_05252_));
 sg13g2_a21oi_1 _13981_ (.A1(net4991),
    .A2(net4272),
    .Y(_00373_),
    .B1(_05252_));
 sg13g2_nor2_1 _13982_ (.A(net2841),
    .B(net4271),
    .Y(_05253_));
 sg13g2_a21oi_1 _13983_ (.A1(net5126),
    .A2(net4271),
    .Y(_00374_),
    .B1(_05253_));
 sg13g2_nor2_1 _13984_ (.A(net2428),
    .B(net4272),
    .Y(_05254_));
 sg13g2_a21oi_1 _13985_ (.A1(net4986),
    .A2(net4272),
    .Y(_00375_),
    .B1(_05254_));
 sg13g2_nor2_1 _13986_ (.A(net2723),
    .B(net4271),
    .Y(_05255_));
 sg13g2_a21oi_1 _13987_ (.A1(net5120),
    .A2(net4271),
    .Y(_00376_),
    .B1(_05255_));
 sg13g2_nor2_1 _13988_ (.A(net2341),
    .B(net4271),
    .Y(_05256_));
 sg13g2_a21oi_1 _13989_ (.A1(net4980),
    .A2(net4271),
    .Y(_00377_),
    .B1(_05256_));
 sg13g2_nor2_2 _13990_ (.A(_02675_),
    .B(net4490),
    .Y(_05257_));
 sg13g2_nand2_1 _13991_ (.Y(_05258_),
    .A(net4326),
    .B(_05257_));
 sg13g2_nand2_1 _13992_ (.Y(_05259_),
    .A(net2159),
    .B(net4270));
 sg13g2_o21ai_1 _13993_ (.B1(_05259_),
    .Y(_00378_),
    .A1(net5042),
    .A2(net4270));
 sg13g2_nand2_1 _13994_ (.Y(_05260_),
    .A(net1987),
    .B(net4269));
 sg13g2_o21ai_1 _13995_ (.B1(_05260_),
    .Y(_00379_),
    .A1(net4876),
    .A2(net4269));
 sg13g2_nand2_1 _13996_ (.Y(_05261_),
    .A(net1963),
    .B(net4270));
 sg13g2_o21ai_1 _13997_ (.B1(_05261_),
    .Y(_00380_),
    .A1(net5035),
    .A2(net4270));
 sg13g2_nand2_1 _13998_ (.Y(_05262_),
    .A(net1966),
    .B(net4270));
 sg13g2_o21ai_1 _13999_ (.B1(_05262_),
    .Y(_00381_),
    .A1(net4870),
    .A2(net4270));
 sg13g2_nand2_1 _14000_ (.Y(_05263_),
    .A(net2063),
    .B(net4269));
 sg13g2_o21ai_1 _14001_ (.B1(_05263_),
    .Y(_00382_),
    .A1(net5034),
    .A2(net4269));
 sg13g2_nand2_1 _14002_ (.Y(_05264_),
    .A(net2136),
    .B(net4270));
 sg13g2_o21ai_1 _14003_ (.B1(_05264_),
    .Y(_00383_),
    .A1(net4864),
    .A2(net4270));
 sg13g2_nand2_1 _14004_ (.Y(_05265_),
    .A(net2104),
    .B(net4269));
 sg13g2_o21ai_1 _14005_ (.B1(_05265_),
    .Y(_00384_),
    .A1(net5028),
    .A2(net4269));
 sg13g2_nand2_1 _14006_ (.Y(_05266_),
    .A(net1777),
    .B(net4269));
 sg13g2_o21ai_1 _14007_ (.B1(_05266_),
    .Y(_00385_),
    .A1(net4862),
    .A2(net4269));
 sg13g2_nand2_1 _14008_ (.Y(_05267_),
    .A(net4320),
    .B(_05257_));
 sg13g2_nand2_1 _14009_ (.Y(_05268_),
    .A(net1821),
    .B(net4267));
 sg13g2_o21ai_1 _14010_ (.B1(_05268_),
    .Y(_00386_),
    .A1(net4853),
    .A2(net4267));
 sg13g2_nand2_1 _14011_ (.Y(_05269_),
    .A(net1826),
    .B(net4268));
 sg13g2_o21ai_1 _14012_ (.B1(_05269_),
    .Y(_00387_),
    .A1(net4847),
    .A2(net4268));
 sg13g2_nand2_1 _14013_ (.Y(_05270_),
    .A(net2072),
    .B(net4267));
 sg13g2_o21ai_1 _14014_ (.B1(_05270_),
    .Y(_00388_),
    .A1(net4842),
    .A2(net4267));
 sg13g2_nand2_1 _14015_ (.Y(_05271_),
    .A(net2062),
    .B(net4267));
 sg13g2_o21ai_1 _14016_ (.B1(_05271_),
    .Y(_00389_),
    .A1(net4837),
    .A2(net4267));
 sg13g2_nand2_1 _14017_ (.Y(_05272_),
    .A(net2059),
    .B(net4267));
 sg13g2_o21ai_1 _14018_ (.B1(_05272_),
    .Y(_00390_),
    .A1(net4832),
    .A2(net4267));
 sg13g2_nand2_1 _14019_ (.Y(_05273_),
    .A(net1931),
    .B(net4268));
 sg13g2_o21ai_1 _14020_ (.B1(_05273_),
    .Y(_00391_),
    .A1(net4825),
    .A2(net4268));
 sg13g2_nand2_1 _14021_ (.Y(_05274_),
    .A(net2122),
    .B(net4268));
 sg13g2_o21ai_1 _14022_ (.B1(_05274_),
    .Y(_00392_),
    .A1(net4820),
    .A2(net4268));
 sg13g2_nand2_1 _14023_ (.Y(_05275_),
    .A(net1877),
    .B(net4268));
 sg13g2_o21ai_1 _14024_ (.B1(_05275_),
    .Y(_00393_),
    .A1(net4815),
    .A2(net4268));
 sg13g2_nor2b_1 _14025_ (.A(net4335),
    .B_N(_05257_),
    .Y(_05276_));
 sg13g2_nor2_1 _14026_ (.A(net2775),
    .B(net4266),
    .Y(_05277_));
 sg13g2_a21oi_1 _14027_ (.A1(net5138),
    .A2(net4266),
    .Y(_00394_),
    .B1(_05277_));
 sg13g2_nor2_1 _14028_ (.A(net2295),
    .B(net4266),
    .Y(_05278_));
 sg13g2_a21oi_1 _14029_ (.A1(net4994),
    .A2(net4266),
    .Y(_00395_),
    .B1(_05278_));
 sg13g2_nor2_1 _14030_ (.A(net2519),
    .B(net4265),
    .Y(_05279_));
 sg13g2_a21oi_1 _14031_ (.A1(net5132),
    .A2(net4265),
    .Y(_00396_),
    .B1(_05279_));
 sg13g2_nor2_1 _14032_ (.A(net2866),
    .B(net4266),
    .Y(_05280_));
 sg13g2_a21oi_1 _14033_ (.A1(net4991),
    .A2(net4266),
    .Y(_00397_),
    .B1(_05280_));
 sg13g2_nor2_1 _14034_ (.A(net2821),
    .B(net4265),
    .Y(_05281_));
 sg13g2_a21oi_1 _14035_ (.A1(net5126),
    .A2(net4265),
    .Y(_00398_),
    .B1(_05281_));
 sg13g2_nor2_1 _14036_ (.A(net2550),
    .B(net4266),
    .Y(_05282_));
 sg13g2_a21oi_1 _14037_ (.A1(net4986),
    .A2(net4266),
    .Y(_00399_),
    .B1(_05282_));
 sg13g2_nor2_1 _14038_ (.A(net2886),
    .B(net4265),
    .Y(_05283_));
 sg13g2_a21oi_1 _14039_ (.A1(net5120),
    .A2(net4265),
    .Y(_00400_),
    .B1(_05283_));
 sg13g2_nor2_1 _14040_ (.A(net2712),
    .B(net4265),
    .Y(_05284_));
 sg13g2_a21oi_1 _14041_ (.A1(net4980),
    .A2(net4265),
    .Y(_00401_),
    .B1(_05284_));
 sg13g2_nor2_1 _14042_ (.A(net5322),
    .B(\m_sys.m_core.m_bru.io_i_s1[14] ),
    .Y(_05285_));
 sg13g2_a21oi_2 _14043_ (.B1(_05285_),
    .Y(_05286_),
    .A2(_00026_),
    .A1(net5322));
 sg13g2_nand2_1 _14044_ (.Y(_05287_),
    .A(net5323),
    .B(_05286_));
 sg13g2_nand2_1 _14045_ (.Y(_05288_),
    .A(net5322),
    .B(\m_sys.m_core.m_bru.io_i_s1[14] ));
 sg13g2_nand2b_1 _14046_ (.Y(_05289_),
    .B(net5224),
    .A_N(_05288_));
 sg13g2_or2_1 _14047_ (.X(_05290_),
    .B(_00026_),
    .A(net5322));
 sg13g2_a21oi_1 _14048_ (.A1(_05288_),
    .A2(_05290_),
    .Y(_05291_),
    .B1(net5323));
 sg13g2_nand2b_1 _14049_ (.Y(_05292_),
    .B(_05287_),
    .A_N(_05291_));
 sg13g2_nor3_2 _14050_ (.A(net5323),
    .B(net5322),
    .C(\m_sys.m_core.m_bru.io_i_s1[14] ),
    .Y(_05293_));
 sg13g2_nand3_1 _14051_ (.B(net5322),
    .C(_00026_),
    .A(net5224),
    .Y(_05294_));
 sg13g2_nor2_1 _14052_ (.A(net5323),
    .B(_05286_),
    .Y(_05295_));
 sg13g2_o21ai_1 _14053_ (.B1(net4957),
    .Y(_05296_),
    .A1(_05292_),
    .A2(_05295_));
 sg13g2_nor3_1 _14054_ (.A(_02368_),
    .B(net5102),
    .C(_03556_),
    .Y(_05297_));
 sg13g2_nand2_1 _14055_ (.Y(_05298_),
    .A(_05296_),
    .B(_05297_));
 sg13g2_a21oi_1 _14056_ (.A1(_02755_),
    .A2(_05298_),
    .Y(_05299_),
    .B1(_02701_));
 sg13g2_nor2_1 _14057_ (.A(net5376),
    .B(_05299_),
    .Y(_00402_));
 sg13g2_a21oi_1 _14058_ (.A1(_05288_),
    .A2(_05294_),
    .Y(_05300_),
    .B1(net4962));
 sg13g2_a22oi_1 _14059_ (.Y(_05301_),
    .B1(net4957),
    .B2(_05300_),
    .A2(net4962),
    .A1(net3085));
 sg13g2_inv_1 _14060_ (.Y(_00403_),
    .A(_05301_));
 sg13g2_nor2b_1 _14061_ (.A(_05293_),
    .B_N(net4957),
    .Y(_05302_));
 sg13g2_nand3_1 _14062_ (.B(net4957),
    .C(_05286_),
    .A(net5323),
    .Y(_05303_));
 sg13g2_nor3_1 _14063_ (.A(net4962),
    .B(net5102),
    .C(_03556_),
    .Y(_05304_));
 sg13g2_a22oi_1 _14064_ (.Y(_00404_),
    .B1(_05303_),
    .B2(_05304_),
    .A2(net4962),
    .A1(_02458_));
 sg13g2_and2_1 _14065_ (.A(net5315),
    .B(_02772_),
    .X(_05305_));
 sg13g2_nand2_1 _14066_ (.Y(_05306_),
    .A(net5315),
    .B(_02772_));
 sg13g2_nor2_1 _14067_ (.A(_05293_),
    .B(_05306_),
    .Y(_05307_));
 sg13g2_a22oi_1 _14068_ (.Y(_05308_),
    .B1(_05300_),
    .B2(_05307_),
    .A2(net4962),
    .A1(net5302));
 sg13g2_inv_1 _14069_ (.Y(_00405_),
    .A(_05308_));
 sg13g2_nand2_1 _14070_ (.Y(_05309_),
    .A(net4974),
    .B(_05305_));
 sg13g2_nand3_1 _14071_ (.B(net5223),
    .C(_00026_),
    .A(\m_sys.m_core.m_bru.io_i_s1[13] ),
    .Y(_05310_));
 sg13g2_nand3_1 _14072_ (.B(_05288_),
    .C(_05290_),
    .A(net5323),
    .Y(_05311_));
 sg13g2_a21oi_1 _14073_ (.A1(_05287_),
    .A2(_05311_),
    .Y(_05312_),
    .B1(_05309_));
 sg13g2_a21o_1 _14074_ (.A2(net4964),
    .A1(net5287),
    .B1(_05312_),
    .X(_00406_));
 sg13g2_nor3_1 _14075_ (.A(net4643),
    .B(net4488),
    .C(net4317),
    .Y(_05313_));
 sg13g2_nor2_1 _14076_ (.A(net2228),
    .B(net4263),
    .Y(_05314_));
 sg13g2_a21oi_1 _14077_ (.A1(net5022),
    .A2(net4263),
    .Y(_00407_),
    .B1(_05314_));
 sg13g2_nor2_1 _14078_ (.A(net2392),
    .B(net4263),
    .Y(_05315_));
 sg13g2_a21oi_1 _14079_ (.A1(net4811),
    .A2(net4263),
    .Y(_00408_),
    .B1(_05315_));
 sg13g2_nor2_1 _14080_ (.A(net2386),
    .B(_05313_),
    .Y(_05316_));
 sg13g2_a21oi_1 _14081_ (.A1(net5019),
    .A2(net4264),
    .Y(_00409_),
    .B1(_05316_));
 sg13g2_nor2_1 _14082_ (.A(net2282),
    .B(net4264),
    .Y(_05317_));
 sg13g2_a21oi_1 _14083_ (.A1(net4808),
    .A2(net4264),
    .Y(_00410_),
    .B1(_05317_));
 sg13g2_nor2_1 _14084_ (.A(net2242),
    .B(net4263),
    .Y(_05318_));
 sg13g2_a21oi_1 _14085_ (.A1(net5011),
    .A2(net4263),
    .Y(_00411_),
    .B1(_05318_));
 sg13g2_nor2_1 _14086_ (.A(net2627),
    .B(net4263),
    .Y(_05319_));
 sg13g2_a21oi_1 _14087_ (.A1(net4801),
    .A2(net4263),
    .Y(_00412_),
    .B1(_05319_));
 sg13g2_nor2_1 _14088_ (.A(net2299),
    .B(net4264),
    .Y(_05320_));
 sg13g2_a21oi_1 _14089_ (.A1(net5005),
    .A2(net4264),
    .Y(_00413_),
    .B1(_05320_));
 sg13g2_nor2_1 _14090_ (.A(net2374),
    .B(net4264),
    .Y(_05321_));
 sg13g2_a21oi_1 _14091_ (.A1(net4798),
    .A2(net4264),
    .Y(_00414_),
    .B1(_05321_));
 sg13g2_nor2b_1 _14092_ (.A(_02677_),
    .B_N(_02681_),
    .Y(_05322_));
 sg13g2_nand2_1 _14093_ (.Y(_05323_),
    .A(_02671_),
    .B(_05322_));
 sg13g2_nor2_2 _14094_ (.A(net4551),
    .B(net4469),
    .Y(_05324_));
 sg13g2_nand2_1 _14095_ (.Y(_05325_),
    .A(net4326),
    .B(_05324_));
 sg13g2_nand2_1 _14096_ (.Y(_05326_),
    .A(net1886),
    .B(net4261));
 sg13g2_o21ai_1 _14097_ (.B1(_05326_),
    .Y(_00415_),
    .A1(net5041),
    .A2(net4262));
 sg13g2_nand2_1 _14098_ (.Y(_05327_),
    .A(net2410),
    .B(net4261));
 sg13g2_o21ai_1 _14099_ (.B1(_05327_),
    .Y(_00416_),
    .A1(net4877),
    .A2(net4261));
 sg13g2_nand2_1 _14100_ (.Y(_05328_),
    .A(net1874),
    .B(net4262));
 sg13g2_o21ai_1 _14101_ (.B1(_05328_),
    .Y(_00417_),
    .A1(net5036),
    .A2(net4262));
 sg13g2_nand2_1 _14102_ (.Y(_05329_),
    .A(net2008),
    .B(net4262));
 sg13g2_o21ai_1 _14103_ (.B1(_05329_),
    .Y(_00418_),
    .A1(net4869),
    .A2(net4262));
 sg13g2_nand2_1 _14104_ (.Y(_05330_),
    .A(net1798),
    .B(net4261));
 sg13g2_o21ai_1 _14105_ (.B1(_05330_),
    .Y(_00419_),
    .A1(net5030),
    .A2(net4261));
 sg13g2_nand2_1 _14106_ (.Y(_05331_),
    .A(net1870),
    .B(net4262));
 sg13g2_o21ai_1 _14107_ (.B1(_05331_),
    .Y(_00420_),
    .A1(net4864),
    .A2(net4262));
 sg13g2_nand2_1 _14108_ (.Y(_05332_),
    .A(net2364),
    .B(_05325_));
 sg13g2_o21ai_1 _14109_ (.B1(_05332_),
    .Y(_00421_),
    .A1(net5029),
    .A2(net4261));
 sg13g2_nand2_1 _14110_ (.Y(_05333_),
    .A(net2498),
    .B(net4261));
 sg13g2_o21ai_1 _14111_ (.B1(_05333_),
    .Y(_00422_),
    .A1(net4863),
    .A2(net4261));
 sg13g2_nor2b_1 _14112_ (.A(net4317),
    .B_N(_05229_),
    .Y(_05334_));
 sg13g2_nor2_1 _14113_ (.A(net2781),
    .B(net4259),
    .Y(_05335_));
 sg13g2_a21oi_1 _14114_ (.A1(net5022),
    .A2(net4259),
    .Y(_00423_),
    .B1(_05335_));
 sg13g2_nor2_1 _14115_ (.A(net2387),
    .B(net4259),
    .Y(_05336_));
 sg13g2_a21oi_1 _14116_ (.A1(net4811),
    .A2(net4259),
    .Y(_00424_),
    .B1(_05336_));
 sg13g2_nor2_1 _14117_ (.A(net2856),
    .B(_05334_),
    .Y(_05337_));
 sg13g2_a21oi_1 _14118_ (.A1(net5019),
    .A2(net4260),
    .Y(_00425_),
    .B1(_05337_));
 sg13g2_nor2_1 _14119_ (.A(net2528),
    .B(net4260),
    .Y(_05338_));
 sg13g2_a21oi_1 _14120_ (.A1(net4808),
    .A2(net4260),
    .Y(_00426_),
    .B1(_05338_));
 sg13g2_nor2_1 _14121_ (.A(net2463),
    .B(net4259),
    .Y(_05339_));
 sg13g2_a21oi_1 _14122_ (.A1(net5011),
    .A2(net4259),
    .Y(_00427_),
    .B1(_05339_));
 sg13g2_nor2_1 _14123_ (.A(net2540),
    .B(net4259),
    .Y(_05340_));
 sg13g2_a21oi_1 _14124_ (.A1(net4801),
    .A2(net4259),
    .Y(_00428_),
    .B1(_05340_));
 sg13g2_nor2_1 _14125_ (.A(net2743),
    .B(net4260),
    .Y(_05341_));
 sg13g2_a21oi_1 _14126_ (.A1(net5005),
    .A2(net4260),
    .Y(_00429_),
    .B1(_05341_));
 sg13g2_nor2_1 _14127_ (.A(net2303),
    .B(net4260),
    .Y(_05342_));
 sg13g2_a21oi_1 _14128_ (.A1(net4798),
    .A2(net4260),
    .Y(_00430_),
    .B1(_05342_));
 sg13g2_nand2_1 _14129_ (.Y(_05343_),
    .A(net4320),
    .B(_05324_));
 sg13g2_nand2_1 _14130_ (.Y(_05344_),
    .A(net2102),
    .B(net4258));
 sg13g2_o21ai_1 _14131_ (.B1(_05344_),
    .Y(_00431_),
    .A1(net4853),
    .A2(net4257));
 sg13g2_nand2_1 _14132_ (.Y(_05345_),
    .A(net1938),
    .B(net4258));
 sg13g2_o21ai_1 _14133_ (.B1(_05345_),
    .Y(_00432_),
    .A1(net4848),
    .A2(net4258));
 sg13g2_nand2_1 _14134_ (.Y(_05346_),
    .A(net2141),
    .B(net4257));
 sg13g2_o21ai_1 _14135_ (.B1(_05346_),
    .Y(_00433_),
    .A1(net4842),
    .A2(net4257));
 sg13g2_nand2_1 _14136_ (.Y(_05347_),
    .A(net1896),
    .B(net4258));
 sg13g2_o21ai_1 _14137_ (.B1(_05347_),
    .Y(_00434_),
    .A1(net4837),
    .A2(net4257));
 sg13g2_nand2_1 _14138_ (.Y(_05348_),
    .A(net2028),
    .B(net4257));
 sg13g2_o21ai_1 _14139_ (.B1(_05348_),
    .Y(_00435_),
    .A1(net4832),
    .A2(net4257));
 sg13g2_nand2_1 _14140_ (.Y(_05349_),
    .A(net2132),
    .B(_05343_));
 sg13g2_o21ai_1 _14141_ (.B1(_05349_),
    .Y(_00436_),
    .A1(net4825),
    .A2(net4258));
 sg13g2_nand2_1 _14142_ (.Y(_05350_),
    .A(net2073),
    .B(net4257));
 sg13g2_o21ai_1 _14143_ (.B1(_05350_),
    .Y(_00437_),
    .A1(net4821),
    .A2(net4257));
 sg13g2_nand2_1 _14144_ (.Y(_05351_),
    .A(net2068),
    .B(net4258));
 sg13g2_o21ai_1 _14145_ (.B1(_05351_),
    .Y(_00438_),
    .A1(net4815),
    .A2(net4258));
 sg13g2_nor2b_1 _14146_ (.A(net4317),
    .B_N(_05257_),
    .Y(_05352_));
 sg13g2_nor2_1 _14147_ (.A(net2544),
    .B(net4255),
    .Y(_05353_));
 sg13g2_a21oi_1 _14148_ (.A1(net5022),
    .A2(net4255),
    .Y(_00439_),
    .B1(_05353_));
 sg13g2_nor2_1 _14149_ (.A(net2592),
    .B(net4255),
    .Y(_05354_));
 sg13g2_a21oi_1 _14150_ (.A1(net4811),
    .A2(net4255),
    .Y(_00440_),
    .B1(_05354_));
 sg13g2_nor2_1 _14151_ (.A(net2417),
    .B(_05352_),
    .Y(_05355_));
 sg13g2_a21oi_1 _14152_ (.A1(net5018),
    .A2(net4256),
    .Y(_00441_),
    .B1(_05355_));
 sg13g2_nor2_1 _14153_ (.A(net2741),
    .B(net4256),
    .Y(_05356_));
 sg13g2_a21oi_1 _14154_ (.A1(net4808),
    .A2(net4256),
    .Y(_00442_),
    .B1(_05356_));
 sg13g2_nor2_1 _14155_ (.A(net2523),
    .B(net4255),
    .Y(_05357_));
 sg13g2_a21oi_1 _14156_ (.A1(net5011),
    .A2(net4255),
    .Y(_00443_),
    .B1(_05357_));
 sg13g2_nor2_1 _14157_ (.A(net2450),
    .B(net4255),
    .Y(_05358_));
 sg13g2_a21oi_1 _14158_ (.A1(net4801),
    .A2(net4255),
    .Y(_00444_),
    .B1(_05358_));
 sg13g2_nor2_1 _14159_ (.A(net2852),
    .B(net4256),
    .Y(_05359_));
 sg13g2_a21oi_1 _14160_ (.A1(net5005),
    .A2(net4256),
    .Y(_00445_),
    .B1(_05359_));
 sg13g2_nor2_1 _14161_ (.A(net2298),
    .B(net4256),
    .Y(_05360_));
 sg13g2_a21oi_1 _14162_ (.A1(net4798),
    .A2(net4256),
    .Y(_00446_),
    .B1(_05360_));
 sg13g2_nor2b_1 _14163_ (.A(net4331),
    .B_N(_05324_),
    .Y(_05361_));
 sg13g2_nor2_1 _14164_ (.A(net2720),
    .B(net4254),
    .Y(_05362_));
 sg13g2_a21oi_1 _14165_ (.A1(net5137),
    .A2(net4254),
    .Y(_00447_),
    .B1(_05362_));
 sg13g2_nor2_1 _14166_ (.A(net2692),
    .B(net4254),
    .Y(_05363_));
 sg13g2_a21oi_1 _14167_ (.A1(net4993),
    .A2(net4254),
    .Y(_00448_),
    .B1(_05363_));
 sg13g2_nor2_1 _14168_ (.A(net2531),
    .B(net4253),
    .Y(_05364_));
 sg13g2_a21oi_1 _14169_ (.A1(net5130),
    .A2(net4253),
    .Y(_00449_),
    .B1(_05364_));
 sg13g2_nor2_1 _14170_ (.A(net2414),
    .B(net4254),
    .Y(_05365_));
 sg13g2_a21oi_1 _14171_ (.A1(net4988),
    .A2(net4254),
    .Y(_00450_),
    .B1(_05365_));
 sg13g2_nor2_1 _14172_ (.A(net2434),
    .B(net4253),
    .Y(_05366_));
 sg13g2_a21oi_1 _14173_ (.A1(net5125),
    .A2(net4253),
    .Y(_00451_),
    .B1(_05366_));
 sg13g2_nor2_1 _14174_ (.A(net2360),
    .B(net4254),
    .Y(_05367_));
 sg13g2_a21oi_1 _14175_ (.A1(net4984),
    .A2(net4254),
    .Y(_00452_),
    .B1(_05367_));
 sg13g2_nor2_1 _14176_ (.A(net2873),
    .B(net4253),
    .Y(_05368_));
 sg13g2_a21oi_1 _14177_ (.A1(net5121),
    .A2(net4253),
    .Y(_00453_),
    .B1(_05368_));
 sg13g2_nor2_1 _14178_ (.A(net2628),
    .B(net4253),
    .Y(_05369_));
 sg13g2_a21oi_1 _14179_ (.A1(net4978),
    .A2(net4253),
    .Y(_00454_),
    .B1(_05369_));
 sg13g2_nand2_2 _14180_ (.Y(_05370_),
    .A(_02670_),
    .B(_05322_));
 sg13g2_nor2_2 _14181_ (.A(net4597),
    .B(net4463),
    .Y(_05371_));
 sg13g2_nor2b_1 _14182_ (.A(net4318),
    .B_N(_05371_),
    .Y(_05372_));
 sg13g2_nor2_1 _14183_ (.A(net2816),
    .B(net4251),
    .Y(_05373_));
 sg13g2_a21oi_1 _14184_ (.A1(net5023),
    .A2(net4251),
    .Y(_00455_),
    .B1(_05373_));
 sg13g2_nor2_1 _14185_ (.A(net2760),
    .B(_05372_),
    .Y(_05374_));
 sg13g2_a21oi_1 _14186_ (.A1(net4814),
    .A2(net4252),
    .Y(_00456_),
    .B1(_05374_));
 sg13g2_nor2_1 _14187_ (.A(net2667),
    .B(net4251),
    .Y(_05375_));
 sg13g2_a21oi_1 _14188_ (.A1(net5018),
    .A2(net4251),
    .Y(_00457_),
    .B1(_05375_));
 sg13g2_nor2_1 _14189_ (.A(net2454),
    .B(net4251),
    .Y(_05376_));
 sg13g2_a21oi_1 _14190_ (.A1(net4809),
    .A2(net4251),
    .Y(_00458_),
    .B1(_05376_));
 sg13g2_nor2_1 _14191_ (.A(net2643),
    .B(net4252),
    .Y(_05377_));
 sg13g2_a21oi_1 _14192_ (.A1(net5014),
    .A2(net4252),
    .Y(_00459_),
    .B1(_05377_));
 sg13g2_nor2_1 _14193_ (.A(net2513),
    .B(net4252),
    .Y(_05378_));
 sg13g2_a21oi_1 _14194_ (.A1(net4803),
    .A2(net4252),
    .Y(_00460_),
    .B1(_05378_));
 sg13g2_nor2_1 _14195_ (.A(net2586),
    .B(net4252),
    .Y(_05379_));
 sg13g2_a21oi_1 _14196_ (.A1(net5007),
    .A2(net4252),
    .Y(_00461_),
    .B1(_05379_));
 sg13g2_nor2_1 _14197_ (.A(net2339),
    .B(net4251),
    .Y(_05380_));
 sg13g2_a21oi_1 _14198_ (.A1(net4799),
    .A2(net4251),
    .Y(_00462_),
    .B1(_05380_));
 sg13g2_nor2_2 _14199_ (.A(net4506),
    .B(net4471),
    .Y(_05381_));
 sg13g2_nand2_1 _14200_ (.Y(_05382_),
    .A(net4327),
    .B(_05381_));
 sg13g2_nand2_1 _14201_ (.Y(_05383_),
    .A(net1838),
    .B(net4250));
 sg13g2_o21ai_1 _14202_ (.B1(_05383_),
    .Y(_00463_),
    .A1(net5041),
    .A2(net4250));
 sg13g2_nand2_1 _14203_ (.Y(_05384_),
    .A(net2018),
    .B(net4250));
 sg13g2_o21ai_1 _14204_ (.B1(_05384_),
    .Y(_00464_),
    .A1(net4877),
    .A2(net4250));
 sg13g2_nand2_1 _14205_ (.Y(_05385_),
    .A(net1979),
    .B(net4249));
 sg13g2_o21ai_1 _14206_ (.B1(_05385_),
    .Y(_00465_),
    .A1(net5036),
    .A2(net4249));
 sg13g2_nand2_1 _14207_ (.Y(_05386_),
    .A(net2249),
    .B(net4249));
 sg13g2_o21ai_1 _14208_ (.B1(_05386_),
    .Y(_00466_),
    .A1(net4869),
    .A2(net4249));
 sg13g2_nand2_1 _14209_ (.Y(_05387_),
    .A(net1790),
    .B(net4249));
 sg13g2_o21ai_1 _14210_ (.B1(_05387_),
    .Y(_00467_),
    .A1(net5030),
    .A2(net4249));
 sg13g2_nand2_1 _14211_ (.Y(_05388_),
    .A(net2353),
    .B(net4249));
 sg13g2_o21ai_1 _14212_ (.B1(_05388_),
    .Y(_00468_),
    .A1(_04944_),
    .A2(net4249));
 sg13g2_nand2_1 _14213_ (.Y(_05389_),
    .A(net1765),
    .B(net4250));
 sg13g2_o21ai_1 _14214_ (.B1(_05389_),
    .Y(_00469_),
    .A1(net5029),
    .A2(net4250));
 sg13g2_nand2_1 _14215_ (.Y(_05390_),
    .A(net2193),
    .B(net4250));
 sg13g2_o21ai_1 _14216_ (.B1(_05390_),
    .Y(_00470_),
    .A1(net4863),
    .A2(net4250));
 sg13g2_nor2_2 _14217_ (.A(_02644_),
    .B(net4463),
    .Y(_05391_));
 sg13g2_nor2b_1 _14218_ (.A(net4318),
    .B_N(_05391_),
    .Y(_05392_));
 sg13g2_nor2_1 _14219_ (.A(net2217),
    .B(net4246),
    .Y(_05393_));
 sg13g2_a21oi_1 _14220_ (.A1(net5023),
    .A2(net4246),
    .Y(_00471_),
    .B1(_05393_));
 sg13g2_nor2_1 _14221_ (.A(net2390),
    .B(net4248),
    .Y(_05394_));
 sg13g2_a21oi_1 _14222_ (.A1(net4814),
    .A2(net4248),
    .Y(_00472_),
    .B1(_05394_));
 sg13g2_nor2_1 _14223_ (.A(net2754),
    .B(net4246),
    .Y(_05395_));
 sg13g2_a21oi_1 _14224_ (.A1(_05138_),
    .A2(net4246),
    .Y(_00473_),
    .B1(_05395_));
 sg13g2_nor2_1 _14225_ (.A(net2564),
    .B(net4246),
    .Y(_05396_));
 sg13g2_a21oi_1 _14226_ (.A1(net4809),
    .A2(net4246),
    .Y(_00474_),
    .B1(_05396_));
 sg13g2_nor2_1 _14227_ (.A(net2408),
    .B(net4248),
    .Y(_05397_));
 sg13g2_a21oi_1 _14228_ (.A1(net5014),
    .A2(net4248),
    .Y(_00475_),
    .B1(_05397_));
 sg13g2_nor2_1 _14229_ (.A(net2194),
    .B(net4247),
    .Y(_05398_));
 sg13g2_a21oi_1 _14230_ (.A1(net4803),
    .A2(net4247),
    .Y(_00476_),
    .B1(_05398_));
 sg13g2_nor2_1 _14231_ (.A(net2624),
    .B(net4246),
    .Y(_05399_));
 sg13g2_a21oi_1 _14232_ (.A1(net5007),
    .A2(net4246),
    .Y(_00477_),
    .B1(_05399_));
 sg13g2_nor2_1 _14233_ (.A(net2785),
    .B(net4247),
    .Y(_05400_));
 sg13g2_a21oi_1 _14234_ (.A1(net4799),
    .A2(net4247),
    .Y(_00478_),
    .B1(_05400_));
 sg13g2_nand2_1 _14235_ (.Y(_05401_),
    .A(net4320),
    .B(_05381_));
 sg13g2_nand2_1 _14236_ (.Y(_05402_),
    .A(net1797),
    .B(net4245));
 sg13g2_o21ai_1 _14237_ (.B1(_05402_),
    .Y(_00479_),
    .A1(net4853),
    .A2(net4244));
 sg13g2_nand2_1 _14238_ (.Y(_05403_),
    .A(net2020),
    .B(net4245));
 sg13g2_o21ai_1 _14239_ (.B1(_05403_),
    .Y(_00480_),
    .A1(net4848),
    .A2(net4245));
 sg13g2_nand2_1 _14240_ (.Y(_05404_),
    .A(net1906),
    .B(net4244));
 sg13g2_o21ai_1 _14241_ (.B1(_05404_),
    .Y(_00481_),
    .A1(net4842),
    .A2(net4244));
 sg13g2_nand2_1 _14242_ (.Y(_05405_),
    .A(net1872),
    .B(net4244));
 sg13g2_o21ai_1 _14243_ (.B1(_05405_),
    .Y(_00482_),
    .A1(net4837),
    .A2(net4244));
 sg13g2_nand2_1 _14244_ (.Y(_05406_),
    .A(net2060),
    .B(net4244));
 sg13g2_o21ai_1 _14245_ (.B1(_05406_),
    .Y(_00483_),
    .A1(net4831),
    .A2(net4244));
 sg13g2_nand2_1 _14246_ (.Y(_05407_),
    .A(net1887),
    .B(net4245));
 sg13g2_o21ai_1 _14247_ (.B1(_05407_),
    .Y(_00484_),
    .A1(net4825),
    .A2(net4245));
 sg13g2_nand2_1 _14248_ (.Y(_05408_),
    .A(net1795),
    .B(_05401_));
 sg13g2_o21ai_1 _14249_ (.B1(_05408_),
    .Y(_00485_),
    .A1(net4820),
    .A2(net4244));
 sg13g2_nand2_1 _14250_ (.Y(_05409_),
    .A(net1862),
    .B(net4245));
 sg13g2_o21ai_1 _14251_ (.B1(_05409_),
    .Y(_00486_),
    .A1(net4815),
    .A2(net4245));
 sg13g2_nor2_2 _14252_ (.A(net4643),
    .B(net4470),
    .Y(_05410_));
 sg13g2_nor2b_1 _14253_ (.A(net4331),
    .B_N(_05410_),
    .Y(_05411_));
 sg13g2_nor2_1 _14254_ (.A(net2426),
    .B(net4243),
    .Y(_05412_));
 sg13g2_a21oi_1 _14255_ (.A1(net5137),
    .A2(net4243),
    .Y(_00487_),
    .B1(_05412_));
 sg13g2_nor2_1 _14256_ (.A(net2622),
    .B(net4243),
    .Y(_05413_));
 sg13g2_a21oi_1 _14257_ (.A1(net4993),
    .A2(net4243),
    .Y(_00488_),
    .B1(_05413_));
 sg13g2_nor2_1 _14258_ (.A(net2286),
    .B(net4242),
    .Y(_05414_));
 sg13g2_a21oi_1 _14259_ (.A1(net5130),
    .A2(net4242),
    .Y(_00489_),
    .B1(_05414_));
 sg13g2_nor2_1 _14260_ (.A(net2637),
    .B(net4242),
    .Y(_05415_));
 sg13g2_a21oi_1 _14261_ (.A1(net4989),
    .A2(net4242),
    .Y(_00490_),
    .B1(_05415_));
 sg13g2_nor2_1 _14262_ (.A(net2362),
    .B(net4243),
    .Y(_05416_));
 sg13g2_a21oi_1 _14263_ (.A1(net5125),
    .A2(net4243),
    .Y(_00491_),
    .B1(_05416_));
 sg13g2_nor2_1 _14264_ (.A(net2174),
    .B(net4242),
    .Y(_05417_));
 sg13g2_a21oi_1 _14265_ (.A1(net4984),
    .A2(net4242),
    .Y(_00492_),
    .B1(_05417_));
 sg13g2_nor2_1 _14266_ (.A(net2269),
    .B(net4243),
    .Y(_05418_));
 sg13g2_a21oi_1 _14267_ (.A1(net5121),
    .A2(net4243),
    .Y(_00493_),
    .B1(_05418_));
 sg13g2_nor2_1 _14268_ (.A(net2422),
    .B(net4242),
    .Y(_05419_));
 sg13g2_a21oi_1 _14269_ (.A1(net4978),
    .A2(net4242),
    .Y(_00494_),
    .B1(_05419_));
 sg13g2_nor2_2 _14270_ (.A(net4551),
    .B(net4462),
    .Y(_05420_));
 sg13g2_nor2b_1 _14271_ (.A(net4318),
    .B_N(_05420_),
    .Y(_05421_));
 sg13g2_nor2_1 _14272_ (.A(net2165),
    .B(net4240),
    .Y(_05422_));
 sg13g2_a21oi_1 _14273_ (.A1(net5023),
    .A2(net4240),
    .Y(_00495_),
    .B1(_05422_));
 sg13g2_nor2_1 _14274_ (.A(net2783),
    .B(_05421_),
    .Y(_05423_));
 sg13g2_a21oi_1 _14275_ (.A1(net4814),
    .A2(net4241),
    .Y(_00496_),
    .B1(_05423_));
 sg13g2_nor2_1 _14276_ (.A(net2263),
    .B(net4240),
    .Y(_05424_));
 sg13g2_a21oi_1 _14277_ (.A1(net5018),
    .A2(net4240),
    .Y(_00497_),
    .B1(_05424_));
 sg13g2_nor2_1 _14278_ (.A(net2864),
    .B(net4240),
    .Y(_05425_));
 sg13g2_a21oi_1 _14279_ (.A1(net4808),
    .A2(net4240),
    .Y(_00498_),
    .B1(_05425_));
 sg13g2_nor2_1 _14280_ (.A(net2875),
    .B(net4241),
    .Y(_05426_));
 sg13g2_a21oi_1 _14281_ (.A1(net5014),
    .A2(net4241),
    .Y(_00499_),
    .B1(_05426_));
 sg13g2_nor2_1 _14282_ (.A(net2518),
    .B(net4241),
    .Y(_05427_));
 sg13g2_a21oi_1 _14283_ (.A1(net4803),
    .A2(net4241),
    .Y(_00500_),
    .B1(_05427_));
 sg13g2_nor2_1 _14284_ (.A(net2832),
    .B(net4241),
    .Y(_05428_));
 sg13g2_a21oi_1 _14285_ (.A1(net5007),
    .A2(net4241),
    .Y(_00501_),
    .B1(_05428_));
 sg13g2_nor2_1 _14286_ (.A(net2347),
    .B(net4240),
    .Y(_05429_));
 sg13g2_a21oi_1 _14287_ (.A1(net4799),
    .A2(net4240),
    .Y(_00502_),
    .B1(_05429_));
 sg13g2_nor2b_1 _14288_ (.A(net4331),
    .B_N(_05381_),
    .Y(_05430_));
 sg13g2_nor2_1 _14289_ (.A(net2634),
    .B(net4239),
    .Y(_05431_));
 sg13g2_a21oi_1 _14290_ (.A1(net5137),
    .A2(net4239),
    .Y(_00503_),
    .B1(_05431_));
 sg13g2_nor2_1 _14291_ (.A(net2468),
    .B(net4239),
    .Y(_05432_));
 sg13g2_a21oi_1 _14292_ (.A1(net4994),
    .A2(net4239),
    .Y(_00504_),
    .B1(_05432_));
 sg13g2_nor2_1 _14293_ (.A(net2395),
    .B(net4238),
    .Y(_05433_));
 sg13g2_a21oi_1 _14294_ (.A1(net5130),
    .A2(net4238),
    .Y(_00505_),
    .B1(_05433_));
 sg13g2_nor2_1 _14295_ (.A(net2251),
    .B(net4238),
    .Y(_05434_));
 sg13g2_a21oi_1 _14296_ (.A1(net4989),
    .A2(net4238),
    .Y(_00506_),
    .B1(_05434_));
 sg13g2_nor2_1 _14297_ (.A(net2797),
    .B(net4239),
    .Y(_05435_));
 sg13g2_a21oi_1 _14298_ (.A1(net5125),
    .A2(net4239),
    .Y(_00507_),
    .B1(_05435_));
 sg13g2_nor2_1 _14299_ (.A(net2746),
    .B(net4238),
    .Y(_05436_));
 sg13g2_a21oi_1 _14300_ (.A1(net4984),
    .A2(net4238),
    .Y(_00508_),
    .B1(_05436_));
 sg13g2_nor2_1 _14301_ (.A(net2794),
    .B(net4239),
    .Y(_05437_));
 sg13g2_a21oi_1 _14302_ (.A1(net5120),
    .A2(net4239),
    .Y(_00509_),
    .B1(_05437_));
 sg13g2_nor2_1 _14303_ (.A(net2704),
    .B(net4238),
    .Y(_05438_));
 sg13g2_a21oi_1 _14304_ (.A1(net4978),
    .A2(net4238),
    .Y(_00510_),
    .B1(_05438_));
 sg13g2_nor2_2 _14305_ (.A(net4643),
    .B(net4481),
    .Y(_05439_));
 sg13g2_nor2b_1 _14306_ (.A(net4317),
    .B_N(_05439_),
    .Y(_05440_));
 sg13g2_nor2_1 _14307_ (.A(net2596),
    .B(net4236),
    .Y(_05441_));
 sg13g2_a21oi_1 _14308_ (.A1(net5025),
    .A2(net4236),
    .Y(_00511_),
    .B1(_05441_));
 sg13g2_nor2_1 _14309_ (.A(net2766),
    .B(net4236),
    .Y(_05442_));
 sg13g2_a21oi_1 _14310_ (.A1(net4811),
    .A2(net4236),
    .Y(_00512_),
    .B1(_05442_));
 sg13g2_nor2_1 _14311_ (.A(net2470),
    .B(net4237),
    .Y(_05443_));
 sg13g2_a21oi_1 _14312_ (.A1(net5018),
    .A2(net4237),
    .Y(_00513_),
    .B1(_05443_));
 sg13g2_nor2_1 _14313_ (.A(net2317),
    .B(net4237),
    .Y(_05444_));
 sg13g2_a21oi_1 _14314_ (.A1(net4808),
    .A2(net4237),
    .Y(_00514_),
    .B1(_05444_));
 sg13g2_nor2_1 _14315_ (.A(net2642),
    .B(net4236),
    .Y(_05445_));
 sg13g2_a21oi_1 _14316_ (.A1(net5011),
    .A2(net4236),
    .Y(_00515_),
    .B1(_05445_));
 sg13g2_nor2_1 _14317_ (.A(net2293),
    .B(net4237),
    .Y(_05446_));
 sg13g2_a21oi_1 _14318_ (.A1(net4801),
    .A2(net4237),
    .Y(_00516_),
    .B1(_05446_));
 sg13g2_nor2_1 _14319_ (.A(net2292),
    .B(net4236),
    .Y(_05447_));
 sg13g2_a21oi_1 _14320_ (.A1(net5005),
    .A2(net4236),
    .Y(_00517_),
    .B1(_05447_));
 sg13g2_nor2_1 _14321_ (.A(net2583),
    .B(net4237),
    .Y(_05448_));
 sg13g2_a21oi_1 _14322_ (.A1(net4798),
    .A2(net4237),
    .Y(_00518_),
    .B1(_05448_));
 sg13g2_nor2_2 _14323_ (.A(net4597),
    .B(net4499),
    .Y(_05449_));
 sg13g2_nand2_1 _14324_ (.Y(_05450_),
    .A(net4329),
    .B(_05449_));
 sg13g2_nand2_1 _14325_ (.Y(_05451_),
    .A(net2180),
    .B(net4234));
 sg13g2_o21ai_1 _14326_ (.B1(_05451_),
    .Y(_00519_),
    .A1(net5044),
    .A2(net4234));
 sg13g2_nand2_1 _14327_ (.Y(_05452_),
    .A(net1883),
    .B(net4235));
 sg13g2_o21ai_1 _14328_ (.B1(_05452_),
    .Y(_00520_),
    .A1(net4874),
    .A2(net4235));
 sg13g2_nand2_1 _14329_ (.Y(_05453_),
    .A(net2157),
    .B(net4235));
 sg13g2_o21ai_1 _14330_ (.B1(_05453_),
    .Y(_00521_),
    .A1(net5039),
    .A2(_05450_));
 sg13g2_nand2_1 _14331_ (.Y(_05454_),
    .A(net2056),
    .B(net4234));
 sg13g2_o21ai_1 _14332_ (.B1(_05454_),
    .Y(_00522_),
    .A1(net4872),
    .A2(net4234));
 sg13g2_nand2_1 _14333_ (.Y(_05455_),
    .A(net1892),
    .B(net4234));
 sg13g2_o21ai_1 _14334_ (.B1(_05455_),
    .Y(_00523_),
    .A1(net5033),
    .A2(net4234));
 sg13g2_nand2_1 _14335_ (.Y(_05456_),
    .A(net2096),
    .B(net4234));
 sg13g2_o21ai_1 _14336_ (.B1(_05456_),
    .Y(_00524_),
    .A1(net4867),
    .A2(net4234));
 sg13g2_nand2_1 _14337_ (.Y(_05457_),
    .A(net1842),
    .B(net4235));
 sg13g2_o21ai_1 _14338_ (.B1(_05457_),
    .Y(_00525_),
    .A1(net5026),
    .A2(net4235));
 sg13g2_nand2_1 _14339_ (.Y(_05458_),
    .A(net1843),
    .B(net4235));
 sg13g2_o21ai_1 _14340_ (.B1(_05458_),
    .Y(_00526_),
    .A1(net4861),
    .A2(net4235));
 sg13g2_nor2_2 _14341_ (.A(net4597),
    .B(net4470),
    .Y(_05459_));
 sg13g2_nor2b_1 _14342_ (.A(net4316),
    .B_N(_05459_),
    .Y(_05460_));
 sg13g2_nor2_1 _14343_ (.A(net2261),
    .B(net4233),
    .Y(_05461_));
 sg13g2_a21oi_1 _14344_ (.A1(net5021),
    .A2(net4233),
    .Y(_00527_),
    .B1(_05461_));
 sg13g2_nor2_1 _14345_ (.A(net2499),
    .B(net4232),
    .Y(_05462_));
 sg13g2_a21oi_1 _14346_ (.A1(net4810),
    .A2(net4232),
    .Y(_00528_),
    .B1(_05462_));
 sg13g2_nor2_1 _14347_ (.A(net2230),
    .B(net4233),
    .Y(_05463_));
 sg13g2_a21oi_1 _14348_ (.A1(net5015),
    .A2(_05460_),
    .Y(_00529_),
    .B1(_05463_));
 sg13g2_nor2_1 _14349_ (.A(net2342),
    .B(net4233),
    .Y(_05464_));
 sg13g2_a21oi_1 _14350_ (.A1(net4805),
    .A2(net4233),
    .Y(_00530_),
    .B1(_05464_));
 sg13g2_nor2_1 _14351_ (.A(net2240),
    .B(net4232),
    .Y(_05465_));
 sg13g2_a21oi_1 _14352_ (.A1(net5010),
    .A2(net4232),
    .Y(_00531_),
    .B1(_05465_));
 sg13g2_nor2_1 _14353_ (.A(net2955),
    .B(net4232),
    .Y(_05466_));
 sg13g2_a21oi_1 _14354_ (.A1(net4800),
    .A2(net4232),
    .Y(_00532_),
    .B1(_05466_));
 sg13g2_nor2_1 _14355_ (.A(net2607),
    .B(net4233),
    .Y(_05467_));
 sg13g2_a21oi_1 _14356_ (.A1(net5006),
    .A2(net4233),
    .Y(_00533_),
    .B1(_05467_));
 sg13g2_nor2_1 _14357_ (.A(net2569),
    .B(net4232),
    .Y(_05468_));
 sg13g2_a21oi_1 _14358_ (.A1(net4795),
    .A2(net4232),
    .Y(_00534_),
    .B1(_05468_));
 sg13g2_nand2_1 _14359_ (.Y(_05469_),
    .A(net4323),
    .B(_05449_));
 sg13g2_nand2_1 _14360_ (.Y(_05470_),
    .A(net1685),
    .B(net4231));
 sg13g2_o21ai_1 _14361_ (.B1(_05470_),
    .Y(_00535_),
    .A1(net4857),
    .A2(net4231));
 sg13g2_nand2_1 _14362_ (.Y(_05471_),
    .A(net2021),
    .B(net4230));
 sg13g2_o21ai_1 _14363_ (.B1(_05471_),
    .Y(_00536_),
    .A1(net4849),
    .A2(net4230));
 sg13g2_nand2_1 _14364_ (.Y(_05472_),
    .A(net1837),
    .B(net4231));
 sg13g2_o21ai_1 _14365_ (.B1(_05472_),
    .Y(_00537_),
    .A1(net4846),
    .A2(net4231));
 sg13g2_nand2_1 _14366_ (.Y(_05473_),
    .A(net1754),
    .B(net4230));
 sg13g2_o21ai_1 _14367_ (.B1(_05473_),
    .Y(_00538_),
    .A1(net4841),
    .A2(net4230));
 sg13g2_nand2_1 _14368_ (.Y(_05474_),
    .A(net1941),
    .B(net4231));
 sg13g2_o21ai_1 _14369_ (.B1(_05474_),
    .Y(_00539_),
    .A1(net4835),
    .A2(net4231));
 sg13g2_nand2_1 _14370_ (.Y(_05475_),
    .A(net1925),
    .B(net4230));
 sg13g2_o21ai_1 _14371_ (.B1(_05475_),
    .Y(_00540_),
    .A1(net4827),
    .A2(net4230));
 sg13g2_nand2_1 _14372_ (.Y(_05476_),
    .A(net2170),
    .B(net4231));
 sg13g2_o21ai_1 _14373_ (.B1(_05476_),
    .Y(_00541_),
    .A1(net4823),
    .A2(net4231));
 sg13g2_nand2_1 _14374_ (.Y(_05477_),
    .A(net1752),
    .B(net4230));
 sg13g2_o21ai_1 _14375_ (.B1(_05477_),
    .Y(_00542_),
    .A1(net4817),
    .A2(net4230));
 sg13g2_nor2b_1 _14376_ (.A(net4316),
    .B_N(_05410_),
    .Y(_05478_));
 sg13g2_nor2_1 _14377_ (.A(net2545),
    .B(net4229),
    .Y(_05479_));
 sg13g2_a21oi_1 _14378_ (.A1(net5021),
    .A2(net4229),
    .Y(_00543_),
    .B1(_05479_));
 sg13g2_nor2_1 _14379_ (.A(net2146),
    .B(net4228),
    .Y(_05480_));
 sg13g2_a21oi_1 _14380_ (.A1(net4810),
    .A2(net4228),
    .Y(_00544_),
    .B1(_05480_));
 sg13g2_nor2_1 _14381_ (.A(net2223),
    .B(net4229),
    .Y(_05481_));
 sg13g2_a21oi_1 _14382_ (.A1(net5015),
    .A2(net4229),
    .Y(_00545_),
    .B1(_05481_));
 sg13g2_nor2_1 _14383_ (.A(net2216),
    .B(net4229),
    .Y(_05482_));
 sg13g2_a21oi_1 _14384_ (.A1(net4805),
    .A2(_05478_),
    .Y(_00546_),
    .B1(_05482_));
 sg13g2_nor2_1 _14385_ (.A(net2258),
    .B(net4228),
    .Y(_05483_));
 sg13g2_a21oi_1 _14386_ (.A1(net5010),
    .A2(net4228),
    .Y(_00547_),
    .B1(_05483_));
 sg13g2_nor2_1 _14387_ (.A(net2259),
    .B(net4228),
    .Y(_05484_));
 sg13g2_a21oi_1 _14388_ (.A1(net4800),
    .A2(net4228),
    .Y(_00548_),
    .B1(_05484_));
 sg13g2_nor2_1 _14389_ (.A(net2535),
    .B(net4229),
    .Y(_05485_));
 sg13g2_a21oi_1 _14390_ (.A1(net5006),
    .A2(net4229),
    .Y(_00549_),
    .B1(_05485_));
 sg13g2_nor2_1 _14391_ (.A(net2296),
    .B(net4228),
    .Y(_05486_));
 sg13g2_a21oi_1 _14392_ (.A1(net4795),
    .A2(net4228),
    .Y(_00550_),
    .B1(_05486_));
 sg13g2_nor2b_1 _14393_ (.A(net4333),
    .B_N(_05449_),
    .Y(_05487_));
 sg13g2_nor2_1 _14394_ (.A(net2745),
    .B(net4226),
    .Y(_05488_));
 sg13g2_a21oi_1 _14395_ (.A1(net5135),
    .A2(net4226),
    .Y(_00551_),
    .B1(_05488_));
 sg13g2_nor2_1 _14396_ (.A(net2660),
    .B(net4226),
    .Y(_05489_));
 sg13g2_a21oi_1 _14397_ (.A1(net4997),
    .A2(net4226),
    .Y(_00552_),
    .B1(_05489_));
 sg13g2_nor2_1 _14398_ (.A(net2710),
    .B(net4227),
    .Y(_05490_));
 sg13g2_a21oi_1 _14399_ (.A1(net5133),
    .A2(net4227),
    .Y(_00553_),
    .B1(_05490_));
 sg13g2_nor2_1 _14400_ (.A(net2363),
    .B(net4226),
    .Y(_05491_));
 sg13g2_a21oi_1 _14401_ (.A1(net4988),
    .A2(net4226),
    .Y(_00554_),
    .B1(_05491_));
 sg13g2_nor2_1 _14402_ (.A(net2184),
    .B(net4227),
    .Y(_05492_));
 sg13g2_a21oi_1 _14403_ (.A1(net5128),
    .A2(net4227),
    .Y(_00555_),
    .B1(_05492_));
 sg13g2_nor2_1 _14404_ (.A(net2206),
    .B(net4226),
    .Y(_05493_));
 sg13g2_a21oi_1 _14405_ (.A1(net4983),
    .A2(net4226),
    .Y(_00556_),
    .B1(_05493_));
 sg13g2_nor2_1 _14406_ (.A(net2288),
    .B(net4227),
    .Y(_05494_));
 sg13g2_a21oi_1 _14407_ (.A1(net5122),
    .A2(net4227),
    .Y(_00557_),
    .B1(_05494_));
 sg13g2_nor2_1 _14408_ (.A(net2857),
    .B(net4227),
    .Y(_05495_));
 sg13g2_a21oi_1 _14409_ (.A1(net4981),
    .A2(net4227),
    .Y(_00558_),
    .B1(_05495_));
 sg13g2_nor2b_1 _14410_ (.A(net4316),
    .B_N(_05324_),
    .Y(_05496_));
 sg13g2_nor2_1 _14411_ (.A(net2636),
    .B(_05496_),
    .Y(_05497_));
 sg13g2_a21oi_1 _14412_ (.A1(net5021),
    .A2(net4225),
    .Y(_00559_),
    .B1(_05497_));
 sg13g2_nor2_1 _14413_ (.A(net2274),
    .B(net4224),
    .Y(_05498_));
 sg13g2_a21oi_1 _14414_ (.A1(net4810),
    .A2(net4224),
    .Y(_00560_),
    .B1(_05498_));
 sg13g2_nor2_1 _14415_ (.A(net2560),
    .B(net4225),
    .Y(_05499_));
 sg13g2_a21oi_1 _14416_ (.A1(net5015),
    .A2(net4225),
    .Y(_00561_),
    .B1(_05499_));
 sg13g2_nor2_1 _14417_ (.A(net2820),
    .B(net4225),
    .Y(_05500_));
 sg13g2_a21oi_1 _14418_ (.A1(net4805),
    .A2(net4225),
    .Y(_00562_),
    .B1(_05500_));
 sg13g2_nor2_1 _14419_ (.A(net2782),
    .B(net4224),
    .Y(_05501_));
 sg13g2_a21oi_1 _14420_ (.A1(net5010),
    .A2(net4224),
    .Y(_00563_),
    .B1(_05501_));
 sg13g2_nor2_1 _14421_ (.A(net2779),
    .B(net4224),
    .Y(_05502_));
 sg13g2_a21oi_1 _14422_ (.A1(net4800),
    .A2(net4224),
    .Y(_00564_),
    .B1(_05502_));
 sg13g2_nor2_1 _14423_ (.A(net2790),
    .B(net4225),
    .Y(_05503_));
 sg13g2_a21oi_1 _14424_ (.A1(net5006),
    .A2(net4225),
    .Y(_00565_),
    .B1(_05503_));
 sg13g2_nor2_1 _14425_ (.A(net2229),
    .B(net4224),
    .Y(_05504_));
 sg13g2_a21oi_1 _14426_ (.A1(net4795),
    .A2(net4224),
    .Y(_00566_),
    .B1(_05504_));
 sg13g2_nor2_2 _14427_ (.A(_02644_),
    .B(net4500),
    .Y(_05505_));
 sg13g2_nand2_1 _14428_ (.Y(_05506_),
    .A(net4329),
    .B(_05505_));
 sg13g2_nand2_1 _14429_ (.Y(_05507_),
    .A(net1878),
    .B(net4222));
 sg13g2_o21ai_1 _14430_ (.B1(_05507_),
    .Y(_00567_),
    .A1(net5044),
    .A2(_05506_));
 sg13g2_nand2_1 _14431_ (.Y(_05508_),
    .A(net1804),
    .B(net4223));
 sg13g2_o21ai_1 _14432_ (.B1(_05508_),
    .Y(_00568_),
    .A1(net4874),
    .A2(net4223));
 sg13g2_nand2_1 _14433_ (.Y(_05509_),
    .A(net1673),
    .B(net4222));
 sg13g2_o21ai_1 _14434_ (.B1(_05509_),
    .Y(_00569_),
    .A1(net5039),
    .A2(net4222));
 sg13g2_nand2_1 _14435_ (.Y(_05510_),
    .A(net1710),
    .B(net4222));
 sg13g2_o21ai_1 _14436_ (.B1(_05510_),
    .Y(_00570_),
    .A1(net4872),
    .A2(net4222));
 sg13g2_nand2_1 _14437_ (.Y(_05511_),
    .A(net1999),
    .B(net4222));
 sg13g2_o21ai_1 _14438_ (.B1(_05511_),
    .Y(_00571_),
    .A1(net5033),
    .A2(net4223));
 sg13g2_nand2_1 _14439_ (.Y(_05512_),
    .A(net2469),
    .B(net4222));
 sg13g2_o21ai_1 _14440_ (.B1(_05512_),
    .Y(_00572_),
    .A1(net4867),
    .A2(net4222));
 sg13g2_nand2_1 _14441_ (.Y(_05513_),
    .A(net1971),
    .B(net4223));
 sg13g2_o21ai_1 _14442_ (.B1(_05513_),
    .Y(_00573_),
    .A1(net5026),
    .A2(net4223));
 sg13g2_nand2_1 _14443_ (.Y(_05514_),
    .A(net1743),
    .B(net4223));
 sg13g2_o21ai_1 _14444_ (.B1(_05514_),
    .Y(_00574_),
    .A1(net4861),
    .A2(net4223));
 sg13g2_nor2b_1 _14445_ (.A(net4316),
    .B_N(_05381_),
    .Y(_05515_));
 sg13g2_nor2_1 _14446_ (.A(net2909),
    .B(net4220),
    .Y(_05516_));
 sg13g2_a21oi_1 _14447_ (.A1(net5021),
    .A2(net4220),
    .Y(_00575_),
    .B1(_05516_));
 sg13g2_nor2_1 _14448_ (.A(net2620),
    .B(net4219),
    .Y(_05517_));
 sg13g2_a21oi_1 _14449_ (.A1(net4810),
    .A2(net4219),
    .Y(_00576_),
    .B1(_05517_));
 sg13g2_nor2_1 _14450_ (.A(net2907),
    .B(net4221),
    .Y(_05518_));
 sg13g2_a21oi_1 _14451_ (.A1(net5015),
    .A2(net4221),
    .Y(_00577_),
    .B1(_05518_));
 sg13g2_nor2_1 _14452_ (.A(net2319),
    .B(net4221),
    .Y(_05519_));
 sg13g2_a21oi_1 _14453_ (.A1(net4805),
    .A2(net4221),
    .Y(_00578_),
    .B1(_05519_));
 sg13g2_nor2_1 _14454_ (.A(net2839),
    .B(net4219),
    .Y(_05520_));
 sg13g2_a21oi_1 _14455_ (.A1(net5010),
    .A2(net4219),
    .Y(_00579_),
    .B1(_05520_));
 sg13g2_nor2_1 _14456_ (.A(net2604),
    .B(net4219),
    .Y(_05521_));
 sg13g2_a21oi_1 _14457_ (.A1(net4800),
    .A2(net4219),
    .Y(_00580_),
    .B1(_05521_));
 sg13g2_nor2_1 _14458_ (.A(net2654),
    .B(net4219),
    .Y(_05522_));
 sg13g2_a21oi_1 _14459_ (.A1(net5006),
    .A2(net4219),
    .Y(_00581_),
    .B1(_05522_));
 sg13g2_nor2_1 _14460_ (.A(net2798),
    .B(net4220),
    .Y(_05523_));
 sg13g2_a21oi_1 _14461_ (.A1(net4795),
    .A2(net4220),
    .Y(_00582_),
    .B1(_05523_));
 sg13g2_nand2_1 _14462_ (.Y(_05524_),
    .A(net4323),
    .B(_05505_));
 sg13g2_nand2_1 _14463_ (.Y(_05525_),
    .A(net2022),
    .B(net4218));
 sg13g2_o21ai_1 _14464_ (.B1(_05525_),
    .Y(_00583_),
    .A1(net4857),
    .A2(net4218));
 sg13g2_nand2_1 _14465_ (.Y(_05526_),
    .A(net1840),
    .B(net4217));
 sg13g2_o21ai_1 _14466_ (.B1(_05526_),
    .Y(_00584_),
    .A1(net4850),
    .A2(net4217));
 sg13g2_nand2_1 _14467_ (.Y(_05527_),
    .A(net1697),
    .B(net4218));
 sg13g2_o21ai_1 _14468_ (.B1(_05527_),
    .Y(_00585_),
    .A1(net4846),
    .A2(net4218));
 sg13g2_nand2_1 _14469_ (.Y(_05528_),
    .A(net1757),
    .B(net4217));
 sg13g2_o21ai_1 _14470_ (.B1(_05528_),
    .Y(_00586_),
    .A1(net4841),
    .A2(net4217));
 sg13g2_nand2_1 _14471_ (.Y(_05529_),
    .A(net1895),
    .B(net4218));
 sg13g2_o21ai_1 _14472_ (.B1(_05529_),
    .Y(_00587_),
    .A1(net4835),
    .A2(net4218));
 sg13g2_nand2_1 _14473_ (.Y(_05530_),
    .A(net1728),
    .B(net4217));
 sg13g2_o21ai_1 _14474_ (.B1(_05530_),
    .Y(_00588_),
    .A1(net4827),
    .A2(net4217));
 sg13g2_nand2_1 _14475_ (.Y(_05531_),
    .A(net2237),
    .B(net4218));
 sg13g2_o21ai_1 _14476_ (.B1(_05531_),
    .Y(_00589_),
    .A1(net4823),
    .A2(net4218));
 sg13g2_nand2_1 _14477_ (.Y(_05532_),
    .A(net1734),
    .B(net4217));
 sg13g2_o21ai_1 _14478_ (.B1(_05532_),
    .Y(_00590_),
    .A1(net4817),
    .A2(net4217));
 sg13g2_nor2b_1 _14479_ (.A(net4314),
    .B_N(_05449_),
    .Y(_05533_));
 sg13g2_nor2_1 _14480_ (.A(net2572),
    .B(net4215),
    .Y(_05534_));
 sg13g2_a21oi_1 _14481_ (.A1(net5023),
    .A2(net4215),
    .Y(_00591_),
    .B1(_05534_));
 sg13g2_nor2_1 _14482_ (.A(net2810),
    .B(net4216),
    .Y(_05535_));
 sg13g2_a21oi_1 _14483_ (.A1(net4812),
    .A2(net4216),
    .Y(_00592_),
    .B1(_05535_));
 sg13g2_nor2_1 _14484_ (.A(net2337),
    .B(net4214),
    .Y(_05536_));
 sg13g2_a21oi_1 _14485_ (.A1(net5017),
    .A2(net4214),
    .Y(_00593_),
    .B1(_05536_));
 sg13g2_nor2_1 _14486_ (.A(net2582),
    .B(net4214),
    .Y(_05537_));
 sg13g2_a21oi_1 _14487_ (.A1(net4807),
    .A2(net4214),
    .Y(_00594_),
    .B1(_05537_));
 sg13g2_nor2_1 _14488_ (.A(net2761),
    .B(net4216),
    .Y(_05538_));
 sg13g2_a21oi_1 _14489_ (.A1(net5012),
    .A2(net4216),
    .Y(_00595_),
    .B1(_05538_));
 sg13g2_nor2_1 _14490_ (.A(net2399),
    .B(net4214),
    .Y(_05539_));
 sg13g2_a21oi_1 _14491_ (.A1(net4802),
    .A2(net4214),
    .Y(_00596_),
    .B1(_05539_));
 sg13g2_nor2_1 _14492_ (.A(net2195),
    .B(net4214),
    .Y(_05540_));
 sg13g2_a21oi_1 _14493_ (.A1(net5008),
    .A2(net4214),
    .Y(_00597_),
    .B1(_05540_));
 sg13g2_nor2_1 _14494_ (.A(net2813),
    .B(net4215),
    .Y(_05541_));
 sg13g2_a21oi_1 _14495_ (.A1(net4796),
    .A2(net4215),
    .Y(_00598_),
    .B1(_05541_));
 sg13g2_nor2b_1 _14496_ (.A(net4332),
    .B_N(_05505_),
    .Y(_05542_));
 sg13g2_nor2_1 _14497_ (.A(net2457),
    .B(net4212),
    .Y(_05543_));
 sg13g2_a21oi_1 _14498_ (.A1(net5135),
    .A2(net4212),
    .Y(_00599_),
    .B1(_05543_));
 sg13g2_nor2_1 _14499_ (.A(net2371),
    .B(net4212),
    .Y(_05544_));
 sg13g2_a21oi_1 _14500_ (.A1(net4994),
    .A2(net4212),
    .Y(_00600_),
    .B1(_05544_));
 sg13g2_nor2_1 _14501_ (.A(net2328),
    .B(net4213),
    .Y(_05545_));
 sg13g2_a21oi_1 _14502_ (.A1(net5133),
    .A2(net4213),
    .Y(_00601_),
    .B1(_05545_));
 sg13g2_nor2_1 _14503_ (.A(net2530),
    .B(net4212),
    .Y(_05546_));
 sg13g2_a21oi_1 _14504_ (.A1(net4988),
    .A2(net4212),
    .Y(_00602_),
    .B1(_05546_));
 sg13g2_nor2_1 _14505_ (.A(net2330),
    .B(net4213),
    .Y(_05547_));
 sg13g2_a21oi_1 _14506_ (.A1(net5128),
    .A2(net4213),
    .Y(_00603_),
    .B1(_05547_));
 sg13g2_nor2_1 _14507_ (.A(net2219),
    .B(net4212),
    .Y(_05548_));
 sg13g2_a21oi_1 _14508_ (.A1(net4983),
    .A2(net4212),
    .Y(_00604_),
    .B1(_05548_));
 sg13g2_nor2_1 _14509_ (.A(net2323),
    .B(net4213),
    .Y(_05549_));
 sg13g2_a21oi_1 _14510_ (.A1(net5122),
    .A2(net4213),
    .Y(_00605_),
    .B1(_05549_));
 sg13g2_nor2_1 _14511_ (.A(net2382),
    .B(net4213),
    .Y(_05550_));
 sg13g2_a21oi_1 _14512_ (.A1(net4981),
    .A2(net4213),
    .Y(_00606_),
    .B1(_05550_));
 sg13g2_nor2_2 _14513_ (.A(net4506),
    .B(net4463),
    .Y(_05551_));
 sg13g2_nor2b_1 _14514_ (.A(net4334),
    .B_N(_05551_),
    .Y(_05552_));
 sg13g2_nor2_1 _14515_ (.A(net2688),
    .B(net4211),
    .Y(_05553_));
 sg13g2_a21oi_1 _14516_ (.A1(net5139),
    .A2(net4211),
    .Y(_00607_),
    .B1(_05553_));
 sg13g2_nor2_1 _14517_ (.A(net2751),
    .B(net4211),
    .Y(_05554_));
 sg13g2_a21oi_1 _14518_ (.A1(net4996),
    .A2(net4211),
    .Y(_00608_),
    .B1(_05554_));
 sg13g2_nor2_1 _14519_ (.A(net2773),
    .B(net4210),
    .Y(_05555_));
 sg13g2_a21oi_1 _14520_ (.A1(net5134),
    .A2(net4210),
    .Y(_00609_),
    .B1(_05555_));
 sg13g2_nor2_1 _14521_ (.A(net2803),
    .B(net4210),
    .Y(_05556_));
 sg13g2_a21oi_1 _14522_ (.A1(net4992),
    .A2(net4211),
    .Y(_00610_),
    .B1(_05556_));
 sg13g2_nor2_1 _14523_ (.A(net2494),
    .B(_05552_),
    .Y(_05557_));
 sg13g2_a21oi_1 _14524_ (.A1(net5129),
    .A2(net4210),
    .Y(_00611_),
    .B1(_05557_));
 sg13g2_nor2_1 _14525_ (.A(net2874),
    .B(net4211),
    .Y(_05558_));
 sg13g2_a21oi_1 _14526_ (.A1(net4985),
    .A2(net4211),
    .Y(_00612_),
    .B1(_05558_));
 sg13g2_nor2_1 _14527_ (.A(net2744),
    .B(net4210),
    .Y(_05559_));
 sg13g2_a21oi_1 _14528_ (.A1(net5123),
    .A2(net4210),
    .Y(_00613_),
    .B1(_05559_));
 sg13g2_nor2_1 _14529_ (.A(net2568),
    .B(net4210),
    .Y(_05560_));
 sg13g2_a21oi_1 _14530_ (.A1(net4982),
    .A2(net4210),
    .Y(_00614_),
    .B1(_05560_));
 sg13g2_nand2_1 _14531_ (.Y(_05561_),
    .A(_02671_),
    .B(_02682_));
 sg13g2_nor2_2 _14532_ (.A(net4551),
    .B(net4457),
    .Y(_05562_));
 sg13g2_nor2b_1 _14533_ (.A(net4315),
    .B_N(_05562_),
    .Y(_05563_));
 sg13g2_nor2_1 _14534_ (.A(net2658),
    .B(net4208),
    .Y(_05564_));
 sg13g2_a21oi_1 _14535_ (.A1(net5020),
    .A2(net4208),
    .Y(_00615_),
    .B1(_05564_));
 sg13g2_nor2_1 _14536_ (.A(net2765),
    .B(net4209),
    .Y(_05565_));
 sg13g2_a21oi_1 _14537_ (.A1(net4813),
    .A2(net4209),
    .Y(_00616_),
    .B1(_05565_));
 sg13g2_nor2_1 _14538_ (.A(net2606),
    .B(net4208),
    .Y(_05566_));
 sg13g2_a21oi_1 _14539_ (.A1(net5016),
    .A2(net4208),
    .Y(_00617_),
    .B1(_05566_));
 sg13g2_nor2_1 _14540_ (.A(net2616),
    .B(net4208),
    .Y(_05567_));
 sg13g2_a21oi_1 _14541_ (.A1(net4806),
    .A2(net4208),
    .Y(_00618_),
    .B1(_05567_));
 sg13g2_nor2_1 _14542_ (.A(net2267),
    .B(net4209),
    .Y(_05568_));
 sg13g2_a21oi_1 _14543_ (.A1(net5012),
    .A2(net4209),
    .Y(_00619_),
    .B1(_05568_));
 sg13g2_nor2_1 _14544_ (.A(net2497),
    .B(net4209),
    .Y(_05569_));
 sg13g2_a21oi_1 _14545_ (.A1(net4802),
    .A2(_05563_),
    .Y(_00620_),
    .B1(_05569_));
 sg13g2_nor2_1 _14546_ (.A(net2772),
    .B(net4209),
    .Y(_05570_));
 sg13g2_a21oi_1 _14547_ (.A1(net5008),
    .A2(net4209),
    .Y(_00621_),
    .B1(_05570_));
 sg13g2_nor2_1 _14548_ (.A(net2804),
    .B(net4208),
    .Y(_05571_));
 sg13g2_a21oi_1 _14549_ (.A1(net4795),
    .A2(net4208),
    .Y(_00622_),
    .B1(_05571_));
 sg13g2_nor3_1 _14550_ (.A(net4597),
    .B(net4486),
    .C(net4317),
    .Y(_05572_));
 sg13g2_nor2_1 _14551_ (.A(net2700),
    .B(net4207),
    .Y(_05573_));
 sg13g2_a21oi_1 _14552_ (.A1(net5022),
    .A2(net4207),
    .Y(_00623_),
    .B1(_05573_));
 sg13g2_nor2_1 _14553_ (.A(net2747),
    .B(net4206),
    .Y(_05574_));
 sg13g2_a21oi_1 _14554_ (.A1(net4811),
    .A2(net4206),
    .Y(_00624_),
    .B1(_05574_));
 sg13g2_nor2_1 _14555_ (.A(net2333),
    .B(_05572_),
    .Y(_05575_));
 sg13g2_a21oi_1 _14556_ (.A1(net5018),
    .A2(net4207),
    .Y(_00625_),
    .B1(_05575_));
 sg13g2_nor2_1 _14557_ (.A(net2211),
    .B(net4207),
    .Y(_05576_));
 sg13g2_a21oi_1 _14558_ (.A1(net4808),
    .A2(net4207),
    .Y(_00626_),
    .B1(_05576_));
 sg13g2_nor2_1 _14559_ (.A(net2198),
    .B(net4206),
    .Y(_05577_));
 sg13g2_a21oi_1 _14560_ (.A1(net5011),
    .A2(net4206),
    .Y(_00627_),
    .B1(_05577_));
 sg13g2_nor2_1 _14561_ (.A(net2738),
    .B(net4206),
    .Y(_05578_));
 sg13g2_a21oi_1 _14562_ (.A1(net4801),
    .A2(net4206),
    .Y(_00628_),
    .B1(_05578_));
 sg13g2_nor2_1 _14563_ (.A(net2271),
    .B(net4207),
    .Y(_05579_));
 sg13g2_a21oi_1 _14564_ (.A1(net5005),
    .A2(net4207),
    .Y(_00629_),
    .B1(_05579_));
 sg13g2_nor2_1 _14565_ (.A(net2719),
    .B(net4206),
    .Y(_05580_));
 sg13g2_a21oi_1 _14566_ (.A1(net4798),
    .A2(net4206),
    .Y(_00630_),
    .B1(_05580_));
 sg13g2_nor2_2 _14567_ (.A(net4643),
    .B(net4476),
    .Y(_05581_));
 sg13g2_nor2b_1 _14568_ (.A(net4316),
    .B_N(_05581_),
    .Y(_05582_));
 sg13g2_nor2_1 _14569_ (.A(net2304),
    .B(net4203),
    .Y(_05583_));
 sg13g2_a21oi_1 _14570_ (.A1(net5020),
    .A2(net4203),
    .Y(_00631_),
    .B1(_05583_));
 sg13g2_nor2_1 _14571_ (.A(net2266),
    .B(net4203),
    .Y(_05584_));
 sg13g2_a21oi_1 _14572_ (.A1(net4810),
    .A2(net4203),
    .Y(_00632_),
    .B1(_05584_));
 sg13g2_nor2_1 _14573_ (.A(net2334),
    .B(net4205),
    .Y(_05585_));
 sg13g2_a21oi_1 _14574_ (.A1(net5016),
    .A2(net4205),
    .Y(_00633_),
    .B1(_05585_));
 sg13g2_nor2_1 _14575_ (.A(net2461),
    .B(net4204),
    .Y(_05586_));
 sg13g2_a21oi_1 _14576_ (.A1(net4806),
    .A2(net4204),
    .Y(_00634_),
    .B1(_05586_));
 sg13g2_nor2_1 _14577_ (.A(net2127),
    .B(net4203),
    .Y(_05587_));
 sg13g2_a21oi_1 _14578_ (.A1(net5010),
    .A2(net4203),
    .Y(_00635_),
    .B1(_05587_));
 sg13g2_nor2_1 _14579_ (.A(net3039),
    .B(net4203),
    .Y(_05588_));
 sg13g2_a21oi_1 _14580_ (.A1(net4800),
    .A2(net4203),
    .Y(_00636_),
    .B1(_05588_));
 sg13g2_nor2_1 _14581_ (.A(net2477),
    .B(net4205),
    .Y(_05589_));
 sg13g2_a21oi_1 _14582_ (.A1(net5007),
    .A2(net4205),
    .Y(_00637_),
    .B1(_05589_));
 sg13g2_nor2_1 _14583_ (.A(net2529),
    .B(net4204),
    .Y(_05590_));
 sg13g2_a21oi_1 _14584_ (.A1(net4795),
    .A2(net4204),
    .Y(_00638_),
    .B1(_05590_));
 sg13g2_nand2_1 _14585_ (.Y(_05591_),
    .A(net4330),
    .B(_05371_));
 sg13g2_nand2_1 _14586_ (.Y(_05592_),
    .A(net1783),
    .B(net4201));
 sg13g2_o21ai_1 _14587_ (.B1(_05592_),
    .Y(_00639_),
    .A1(net5045),
    .A2(net4201));
 sg13g2_nand2_1 _14588_ (.Y(_05593_),
    .A(net1750),
    .B(net4201));
 sg13g2_o21ai_1 _14589_ (.B1(_05593_),
    .Y(_00640_),
    .A1(net4874),
    .A2(net4201));
 sg13g2_nand2_1 _14590_ (.Y(_05594_),
    .A(net1863),
    .B(net4202));
 sg13g2_o21ai_1 _14591_ (.B1(_05594_),
    .Y(_00641_),
    .A1(net5040),
    .A2(net4202));
 sg13g2_nand2_1 _14592_ (.Y(_05595_),
    .A(net2086),
    .B(net4202));
 sg13g2_o21ai_1 _14593_ (.B1(_05595_),
    .Y(_00642_),
    .A1(net4870),
    .A2(net4202));
 sg13g2_nand2_1 _14594_ (.Y(_05596_),
    .A(net2203),
    .B(net4202));
 sg13g2_o21ai_1 _14595_ (.B1(_05596_),
    .Y(_00643_),
    .A1(net5031),
    .A2(net4202));
 sg13g2_nand2_1 _14596_ (.Y(_05597_),
    .A(net1736),
    .B(net4201));
 sg13g2_o21ai_1 _14597_ (.B1(_05597_),
    .Y(_00644_),
    .A1(net4868),
    .A2(net4201));
 sg13g2_nand2_1 _14598_ (.Y(_05598_),
    .A(net1982),
    .B(net4202));
 sg13g2_o21ai_1 _14599_ (.B1(_05598_),
    .Y(_00645_),
    .A1(net5027),
    .A2(_05591_));
 sg13g2_nand2_1 _14600_ (.Y(_05599_),
    .A(net2079),
    .B(net4201));
 sg13g2_o21ai_1 _14601_ (.B1(_05599_),
    .Y(_00646_),
    .A1(net4859),
    .A2(net4201));
 sg13g2_nand2_1 _14602_ (.Y(_05600_),
    .A(_02684_),
    .B(net4329));
 sg13g2_nand2_1 _14603_ (.Y(_05601_),
    .A(net2188),
    .B(net4199));
 sg13g2_o21ai_1 _14604_ (.B1(_05601_),
    .Y(_00647_),
    .A1(net5044),
    .A2(net4199));
 sg13g2_nand2_1 _14605_ (.Y(_05602_),
    .A(net1935),
    .B(net4200));
 sg13g2_o21ai_1 _14606_ (.B1(_05602_),
    .Y(_00648_),
    .A1(net4874),
    .A2(net4200));
 sg13g2_nand2_1 _14607_ (.Y(_05603_),
    .A(net2098),
    .B(net4200));
 sg13g2_o21ai_1 _14608_ (.B1(_05603_),
    .Y(_00649_),
    .A1(net5039),
    .A2(_05600_));
 sg13g2_nand2_1 _14609_ (.Y(_05604_),
    .A(net1991),
    .B(net4199));
 sg13g2_o21ai_1 _14610_ (.B1(_05604_),
    .Y(_00650_),
    .A1(net4872),
    .A2(net4199));
 sg13g2_nand2_1 _14611_ (.Y(_05605_),
    .A(net2163),
    .B(net4199));
 sg13g2_o21ai_1 _14612_ (.B1(_05605_),
    .Y(_00651_),
    .A1(net5033),
    .A2(net4199));
 sg13g2_nand2_1 _14613_ (.Y(_05606_),
    .A(net2099),
    .B(net4199));
 sg13g2_o21ai_1 _14614_ (.B1(_05606_),
    .Y(_00652_),
    .A1(net4867),
    .A2(net4199));
 sg13g2_nand2_1 _14615_ (.Y(_05607_),
    .A(net1819),
    .B(net4200));
 sg13g2_o21ai_1 _14616_ (.B1(_05607_),
    .Y(_00653_),
    .A1(net5026),
    .A2(net4200));
 sg13g2_nand2_1 _14617_ (.Y(_05608_),
    .A(net1950),
    .B(net4200));
 sg13g2_o21ai_1 _14618_ (.B1(_05608_),
    .Y(_00654_),
    .A1(net4861),
    .A2(net4200));
 sg13g2_nor2_2 _14619_ (.A(_02699_),
    .B(_02753_),
    .Y(_05609_));
 sg13g2_or2_2 _14620_ (.X(_05610_),
    .B(_02753_),
    .A(_02699_));
 sg13g2_nand2_1 _14621_ (.Y(_05611_),
    .A(\m_sys._m_core_io_b_mem_wdata[0] ),
    .B(net3348));
 sg13g2_o21ai_1 _14622_ (.B1(_05611_),
    .Y(_05612_),
    .A1(_02372_),
    .A2(net5310));
 sg13g2_o21ai_1 _14623_ (.B1(net5384),
    .Y(_05613_),
    .A1(_05610_),
    .A2(_05612_));
 sg13g2_a21oi_1 _14624_ (.A1(_02363_),
    .A2(net4793),
    .Y(_00655_),
    .B1(_05613_));
 sg13g2_nand2_1 _14625_ (.Y(_05614_),
    .A(_02402_),
    .B(_04739_));
 sg13g2_a21oi_1 _14626_ (.A1(net5310),
    .A2(_02462_),
    .Y(_05615_),
    .B1(net4793));
 sg13g2_a22oi_1 _14627_ (.Y(_05616_),
    .B1(_05614_),
    .B2(_05615_),
    .A2(net4793),
    .A1(net3343));
 sg13g2_nor2_1 _14628_ (.A(net5376),
    .B(net3344),
    .Y(_00656_));
 sg13g2_nand2b_1 _14629_ (.Y(_05617_),
    .B(net5221),
    .A_N(_04735_));
 sg13g2_a21oi_1 _14630_ (.A1(net5310),
    .A2(net3298),
    .Y(_05618_),
    .B1(net4793));
 sg13g2_a221oi_1 _14631_ (.B2(_05618_),
    .C1(net5376),
    .B1(_05617_),
    .A1(_02362_),
    .Y(_00657_),
    .A2(net4793));
 sg13g2_nand2_1 _14632_ (.Y(_05619_),
    .A(net5221),
    .B(_04691_));
 sg13g2_a21oi_1 _14633_ (.A1(net5311),
    .A2(net3251),
    .Y(_05620_),
    .B1(net4793));
 sg13g2_o21ai_1 _14634_ (.B1(net5384),
    .Y(_05621_),
    .A1(\m_sys.m_core.m_bru.io_i_pc[5] ),
    .A2(_05609_));
 sg13g2_a21oi_1 _14635_ (.A1(_05619_),
    .A2(_05620_),
    .Y(_00658_),
    .B1(_05621_));
 sg13g2_nand2_1 _14636_ (.Y(_05622_),
    .A(net5221),
    .B(_04652_));
 sg13g2_a21oi_1 _14637_ (.A1(net5310),
    .A2(_02464_),
    .Y(_05623_),
    .B1(net4793));
 sg13g2_a22oi_1 _14638_ (.Y(_05624_),
    .B1(_05622_),
    .B2(_05623_),
    .A2(net4793),
    .A1(net3250));
 sg13g2_nor2_1 _14639_ (.A(net5376),
    .B(_05624_),
    .Y(_00659_));
 sg13g2_or2_1 _14640_ (.X(_05625_),
    .B(_04608_),
    .A(net5310));
 sg13g2_a21oi_1 _14641_ (.A1(net5310),
    .A2(net3178),
    .Y(_05626_),
    .B1(net4794));
 sg13g2_o21ai_1 _14642_ (.B1(net5384),
    .Y(_05627_),
    .A1(net3313),
    .A2(_05609_));
 sg13g2_a21oi_1 _14643_ (.A1(_05625_),
    .A2(_05626_),
    .Y(_00660_),
    .B1(_05627_));
 sg13g2_o21ai_1 _14644_ (.B1(net5384),
    .Y(_05628_),
    .A1(\m_sys.m_core.m_bru.io_i_pc[8] ),
    .A2(_05609_));
 sg13g2_nand2_1 _14645_ (.Y(_05629_),
    .A(net5221),
    .B(_04544_));
 sg13g2_a21oi_1 _14646_ (.A1(net5310),
    .A2(net3296),
    .Y(_05630_),
    .B1(net4794));
 sg13g2_a21oi_1 _14647_ (.A1(_05629_),
    .A2(_05630_),
    .Y(_00661_),
    .B1(_05628_));
 sg13g2_nand2_1 _14648_ (.Y(_05631_),
    .A(net5221),
    .B(_04533_));
 sg13g2_a21oi_1 _14649_ (.A1(net5311),
    .A2(net3028),
    .Y(_05632_),
    .B1(net4794));
 sg13g2_o21ai_1 _14650_ (.B1(net5384),
    .Y(_05633_),
    .A1(net3337),
    .A2(_05609_));
 sg13g2_a21oi_1 _14651_ (.A1(_05631_),
    .A2(_05632_),
    .Y(_00662_),
    .B1(_05633_));
 sg13g2_nand2_1 _14652_ (.Y(_05634_),
    .A(net5221),
    .B(_04490_));
 sg13g2_a21oi_1 _14653_ (.A1(net5311),
    .A2(_02472_),
    .Y(_05635_),
    .B1(net4794));
 sg13g2_a22oi_1 _14654_ (.Y(_05636_),
    .B1(_05634_),
    .B2(_05635_),
    .A2(net4794),
    .A1(net3257));
 sg13g2_nor2_1 _14655_ (.A(net5377),
    .B(_05636_),
    .Y(_00663_));
 sg13g2_nand2_1 _14656_ (.Y(_05637_),
    .A(net5221),
    .B(_04417_));
 sg13g2_a21oi_1 _14657_ (.A1(\m_sys._m_core_io_b_mem_wdata[0] ),
    .A2(_02471_),
    .Y(_05638_),
    .B1(net4794));
 sg13g2_a22oi_1 _14658_ (.Y(_05639_),
    .B1(_05637_),
    .B2(_05638_),
    .A2(net4794),
    .A1(net3083));
 sg13g2_nor2_1 _14659_ (.A(net5377),
    .B(net3084),
    .Y(_00664_));
 sg13g2_nor2_2 _14660_ (.A(net4597),
    .B(net4456),
    .Y(_05640_));
 sg13g2_nor2b_1 _14661_ (.A(net4334),
    .B_N(_05640_),
    .Y(_05641_));
 sg13g2_nor2_1 _14662_ (.A(net2763),
    .B(net4198),
    .Y(_05642_));
 sg13g2_a21oi_1 _14663_ (.A1(net5137),
    .A2(net4198),
    .Y(_00665_),
    .B1(_05642_));
 sg13g2_nor2_1 _14664_ (.A(net2381),
    .B(net4198),
    .Y(_05643_));
 sg13g2_a21oi_1 _14665_ (.A1(net4995),
    .A2(net4198),
    .Y(_00666_),
    .B1(_05643_));
 sg13g2_nor2_1 _14666_ (.A(net2706),
    .B(net4197),
    .Y(_05644_));
 sg13g2_a21oi_1 _14667_ (.A1(net5131),
    .A2(net4197),
    .Y(_00667_),
    .B1(_05644_));
 sg13g2_nor2_1 _14668_ (.A(net2427),
    .B(net4198),
    .Y(_05645_));
 sg13g2_a21oi_1 _14669_ (.A1(net4990),
    .A2(net4198),
    .Y(_00668_),
    .B1(_05645_));
 sg13g2_nor2_1 _14670_ (.A(net2256),
    .B(net4197),
    .Y(_05646_));
 sg13g2_a21oi_1 _14671_ (.A1(net5128),
    .A2(net4197),
    .Y(_00669_),
    .B1(_05646_));
 sg13g2_nor2_1 _14672_ (.A(net2548),
    .B(_05641_),
    .Y(_05647_));
 sg13g2_a21oi_1 _14673_ (.A1(net4986),
    .A2(net4198),
    .Y(_00670_),
    .B1(_05647_));
 sg13g2_nor2_1 _14674_ (.A(net2580),
    .B(net4197),
    .Y(_05648_));
 sg13g2_a21oi_1 _14675_ (.A1(net5122),
    .A2(net4197),
    .Y(_00671_),
    .B1(_05648_));
 sg13g2_nor2_1 _14676_ (.A(net2418),
    .B(net4197),
    .Y(_05649_));
 sg13g2_a21oi_1 _14677_ (.A1(net4979),
    .A2(net4197),
    .Y(_00672_),
    .B1(_05649_));
 sg13g2_nand2_1 _14678_ (.Y(_05650_),
    .A(net4326),
    .B(_05410_));
 sg13g2_nand2_1 _14679_ (.Y(_05651_),
    .A(net1921),
    .B(net4195));
 sg13g2_o21ai_1 _14680_ (.B1(_05651_),
    .Y(_00673_),
    .A1(net5041),
    .A2(net4196));
 sg13g2_nand2_1 _14681_ (.Y(_05652_),
    .A(net1663),
    .B(net4195));
 sg13g2_o21ai_1 _14682_ (.B1(_05652_),
    .Y(_00674_),
    .A1(net4877),
    .A2(_05650_));
 sg13g2_nand2_1 _14683_ (.Y(_05653_),
    .A(net1768),
    .B(net4196));
 sg13g2_o21ai_1 _14684_ (.B1(_05653_),
    .Y(_00675_),
    .A1(net5036),
    .A2(net4196));
 sg13g2_nand2_1 _14685_ (.Y(_05654_),
    .A(net1678),
    .B(net4196));
 sg13g2_o21ai_1 _14686_ (.B1(_05654_),
    .Y(_00676_),
    .A1(net4869),
    .A2(net4196));
 sg13g2_nand2_1 _14687_ (.Y(_05655_),
    .A(net1695),
    .B(net4195));
 sg13g2_o21ai_1 _14688_ (.B1(_05655_),
    .Y(_00677_),
    .A1(net5030),
    .A2(net4195));
 sg13g2_nand2_1 _14689_ (.Y(_05656_),
    .A(net1890),
    .B(net4196));
 sg13g2_o21ai_1 _14690_ (.B1(_05656_),
    .Y(_00678_),
    .A1(net4864),
    .A2(net4196));
 sg13g2_nand2_1 _14691_ (.Y(_05657_),
    .A(net1706),
    .B(net4195));
 sg13g2_o21ai_1 _14692_ (.B1(_05657_),
    .Y(_00679_),
    .A1(net5029),
    .A2(net4195));
 sg13g2_nand2_1 _14693_ (.Y(_05658_),
    .A(net1923),
    .B(net4195));
 sg13g2_o21ai_1 _14694_ (.B1(_05658_),
    .Y(_00680_),
    .A1(net4863),
    .A2(net4195));
 sg13g2_nand2_1 _14695_ (.Y(_05659_),
    .A(_02684_),
    .B(net4323));
 sg13g2_nand2_1 _14696_ (.Y(_05660_),
    .A(net1779),
    .B(net4194));
 sg13g2_o21ai_1 _14697_ (.B1(_05660_),
    .Y(_00681_),
    .A1(net4857),
    .A2(net4194));
 sg13g2_nand2_1 _14698_ (.Y(_05661_),
    .A(net1948),
    .B(net4193));
 sg13g2_o21ai_1 _14699_ (.B1(_05661_),
    .Y(_00682_),
    .A1(net4849),
    .A2(net4193));
 sg13g2_nand2_1 _14700_ (.Y(_05662_),
    .A(net1946),
    .B(net4194));
 sg13g2_o21ai_1 _14701_ (.B1(_05662_),
    .Y(_00683_),
    .A1(net4846),
    .A2(net4194));
 sg13g2_nand2_1 _14702_ (.Y(_05663_),
    .A(net2027),
    .B(net4193));
 sg13g2_o21ai_1 _14703_ (.B1(_05663_),
    .Y(_00684_),
    .A1(net4840),
    .A2(net4193));
 sg13g2_nand2_1 _14704_ (.Y(_05664_),
    .A(net1753),
    .B(net4194));
 sg13g2_o21ai_1 _14705_ (.B1(_05664_),
    .Y(_00685_),
    .A1(net4835),
    .A2(net4194));
 sg13g2_nand2_1 _14706_ (.Y(_05665_),
    .A(net1858),
    .B(net4193));
 sg13g2_o21ai_1 _14707_ (.B1(_05665_),
    .Y(_00686_),
    .A1(net4827),
    .A2(net4193));
 sg13g2_nand2_1 _14708_ (.Y(_05666_),
    .A(net1989),
    .B(net4194));
 sg13g2_o21ai_1 _14709_ (.B1(_05666_),
    .Y(_00687_),
    .A1(net4823),
    .A2(net4194));
 sg13g2_nand2_1 _14710_ (.Y(_05667_),
    .A(net1775),
    .B(net4193));
 sg13g2_o21ai_1 _14711_ (.B1(_05667_),
    .Y(_00688_),
    .A1(net4817),
    .A2(net4193));
 sg13g2_nor2_2 _14712_ (.A(net4551),
    .B(net4481),
    .Y(_05668_));
 sg13g2_nor2b_1 _14713_ (.A(net4317),
    .B_N(_05668_),
    .Y(_05669_));
 sg13g2_nor2_1 _14714_ (.A(net2233),
    .B(net4191),
    .Y(_05670_));
 sg13g2_a21oi_1 _14715_ (.A1(net5022),
    .A2(net4191),
    .Y(_00689_),
    .B1(_05670_));
 sg13g2_nor2_1 _14716_ (.A(net2672),
    .B(net4191),
    .Y(_05671_));
 sg13g2_a21oi_1 _14717_ (.A1(net4811),
    .A2(net4191),
    .Y(_00690_),
    .B1(_05671_));
 sg13g2_nor2_1 _14718_ (.A(net2338),
    .B(net4192),
    .Y(_05672_));
 sg13g2_a21oi_1 _14719_ (.A1(net5018),
    .A2(net4192),
    .Y(_00691_),
    .B1(_05672_));
 sg13g2_nor2_1 _14720_ (.A(net2686),
    .B(_05669_),
    .Y(_05673_));
 sg13g2_a21oi_1 _14721_ (.A1(net4808),
    .A2(net4192),
    .Y(_00692_),
    .B1(_05673_));
 sg13g2_nor2_1 _14722_ (.A(net2920),
    .B(net4191),
    .Y(_05674_));
 sg13g2_a21oi_1 _14723_ (.A1(net5011),
    .A2(net4191),
    .Y(_00693_),
    .B1(_05674_));
 sg13g2_nor2_1 _14724_ (.A(net2235),
    .B(net4192),
    .Y(_05675_));
 sg13g2_a21oi_1 _14725_ (.A1(net4801),
    .A2(net4192),
    .Y(_00694_),
    .B1(_05675_));
 sg13g2_nor2_1 _14726_ (.A(net2340),
    .B(net4191),
    .Y(_05676_));
 sg13g2_a21oi_1 _14727_ (.A1(net5005),
    .A2(net4191),
    .Y(_00695_),
    .B1(_05676_));
 sg13g2_nor2_1 _14728_ (.A(net2736),
    .B(net4192),
    .Y(_05677_));
 sg13g2_a21oi_1 _14729_ (.A1(net4798),
    .A2(net4192),
    .Y(_00696_),
    .B1(_05677_));
 sg13g2_nor2_2 _14730_ (.A(net4551),
    .B(net4500),
    .Y(_05678_));
 sg13g2_nor2b_1 _14731_ (.A(net4332),
    .B_N(_05678_),
    .Y(_05679_));
 sg13g2_nor2_1 _14732_ (.A(net2739),
    .B(net4189),
    .Y(_05680_));
 sg13g2_a21oi_1 _14733_ (.A1(net5135),
    .A2(net4189),
    .Y(_00697_),
    .B1(_05680_));
 sg13g2_nor2_1 _14734_ (.A(net2455),
    .B(net4189),
    .Y(_05681_));
 sg13g2_a21oi_1 _14735_ (.A1(net4993),
    .A2(net4189),
    .Y(_00698_),
    .B1(_05681_));
 sg13g2_nor2_1 _14736_ (.A(net2209),
    .B(net4190),
    .Y(_05682_));
 sg13g2_a21oi_1 _14737_ (.A1(net5133),
    .A2(net4190),
    .Y(_00699_),
    .B1(_05682_));
 sg13g2_nor2_1 _14738_ (.A(net2391),
    .B(net4189),
    .Y(_05683_));
 sg13g2_a21oi_1 _14739_ (.A1(net4988),
    .A2(net4189),
    .Y(_00700_),
    .B1(_05683_));
 sg13g2_nor2_1 _14740_ (.A(net2647),
    .B(net4190),
    .Y(_05684_));
 sg13g2_a21oi_1 _14741_ (.A1(net5128),
    .A2(net4190),
    .Y(_00701_),
    .B1(_05684_));
 sg13g2_nor2_1 _14742_ (.A(net2780),
    .B(net4189),
    .Y(_05685_));
 sg13g2_a21oi_1 _14743_ (.A1(net4983),
    .A2(net4189),
    .Y(_00702_),
    .B1(_05685_));
 sg13g2_nor2_1 _14744_ (.A(net2641),
    .B(net4190),
    .Y(_05686_));
 sg13g2_a21oi_1 _14745_ (.A1(net5122),
    .A2(net4190),
    .Y(_00703_),
    .B1(_05686_));
 sg13g2_nor2_1 _14746_ (.A(net2182),
    .B(net4190),
    .Y(_05687_));
 sg13g2_a21oi_1 _14747_ (.A1(net4981),
    .A2(net4190),
    .Y(_00704_),
    .B1(_05687_));
 sg13g2_nor3_1 _14748_ (.A(net4506),
    .B(net4500),
    .C(net4314),
    .Y(_05688_));
 sg13g2_nor2_1 _14749_ (.A(net2812),
    .B(_05688_),
    .Y(_05689_));
 sg13g2_a21oi_1 _14750_ (.A1(net5023),
    .A2(net4188),
    .Y(_00705_),
    .B1(_05689_));
 sg13g2_nor2_1 _14751_ (.A(net2301),
    .B(net4188),
    .Y(_05690_));
 sg13g2_a21oi_1 _14752_ (.A1(net4812),
    .A2(net4188),
    .Y(_00706_),
    .B1(_05690_));
 sg13g2_nor2_1 _14753_ (.A(net2423),
    .B(net4188),
    .Y(_05691_));
 sg13g2_a21oi_1 _14754_ (.A1(net5017),
    .A2(net4187),
    .Y(_00707_),
    .B1(_05691_));
 sg13g2_nor2_1 _14755_ (.A(net2570),
    .B(net4187),
    .Y(_05692_));
 sg13g2_a21oi_1 _14756_ (.A1(net4807),
    .A2(net4187),
    .Y(_00708_),
    .B1(_05692_));
 sg13g2_nor2_1 _14757_ (.A(net2705),
    .B(net4188),
    .Y(_05693_));
 sg13g2_a21oi_1 _14758_ (.A1(net5012),
    .A2(net4188),
    .Y(_00709_),
    .B1(_05693_));
 sg13g2_nor2_1 _14759_ (.A(net2380),
    .B(net4187),
    .Y(_05694_));
 sg13g2_a21oi_1 _14760_ (.A1(net4802),
    .A2(net4187),
    .Y(_00710_),
    .B1(_05694_));
 sg13g2_nor2_1 _14761_ (.A(net2492),
    .B(net4187),
    .Y(_05695_));
 sg13g2_a21oi_1 _14762_ (.A1(net5008),
    .A2(net4187),
    .Y(_00711_),
    .B1(_05695_));
 sg13g2_nor2_1 _14763_ (.A(net2356),
    .B(net4187),
    .Y(_05696_));
 sg13g2_a21oi_1 _14764_ (.A1(net4796),
    .A2(net4188),
    .Y(_00712_),
    .B1(_05696_));
 sg13g2_nor2b_1 _14765_ (.A(net4316),
    .B_N(_05183_),
    .Y(_05697_));
 sg13g2_nor2_1 _14766_ (.A(net2742),
    .B(net4184),
    .Y(_05698_));
 sg13g2_a21oi_1 _14767_ (.A1(net5020),
    .A2(net4184),
    .Y(_00713_),
    .B1(_05698_));
 sg13g2_nor2_1 _14768_ (.A(net2587),
    .B(net4184),
    .Y(_05699_));
 sg13g2_a21oi_1 _14769_ (.A1(net4810),
    .A2(net4184),
    .Y(_00714_),
    .B1(_05699_));
 sg13g2_nor2_1 _14770_ (.A(net2756),
    .B(net4186),
    .Y(_05700_));
 sg13g2_a21oi_1 _14771_ (.A1(net5015),
    .A2(net4186),
    .Y(_00715_),
    .B1(_05700_));
 sg13g2_nor2_1 _14772_ (.A(net2609),
    .B(net4185),
    .Y(_05701_));
 sg13g2_a21oi_1 _14773_ (.A1(net4806),
    .A2(net4185),
    .Y(_00716_),
    .B1(_05701_));
 sg13g2_nor2_1 _14774_ (.A(net2655),
    .B(net4184),
    .Y(_05702_));
 sg13g2_a21oi_1 _14775_ (.A1(net5010),
    .A2(net4184),
    .Y(_00717_),
    .B1(_05702_));
 sg13g2_nor2_1 _14776_ (.A(net2789),
    .B(net4184),
    .Y(_05703_));
 sg13g2_a21oi_1 _14777_ (.A1(net4800),
    .A2(net4184),
    .Y(_00718_),
    .B1(_05703_));
 sg13g2_nor2_1 _14778_ (.A(net2817),
    .B(net4186),
    .Y(_05704_));
 sg13g2_a21oi_1 _14779_ (.A1(net5009),
    .A2(net4186),
    .Y(_00719_),
    .B1(_05704_));
 sg13g2_nor2_1 _14780_ (.A(net2365),
    .B(net4185),
    .Y(_05705_));
 sg13g2_a21oi_1 _14781_ (.A1(net4795),
    .A2(net4185),
    .Y(_00720_),
    .B1(_05705_));
 sg13g2_nand2_1 _14782_ (.Y(_05706_),
    .A(net4323),
    .B(_05678_));
 sg13g2_nand2_1 _14783_ (.Y(_05707_),
    .A(net2164),
    .B(net4183));
 sg13g2_o21ai_1 _14784_ (.B1(_05707_),
    .Y(_00721_),
    .A1(net4857),
    .A2(net4183));
 sg13g2_nand2_1 _14785_ (.Y(_05708_),
    .A(net2101),
    .B(net4182));
 sg13g2_o21ai_1 _14786_ (.B1(_05708_),
    .Y(_00722_),
    .A1(net4849),
    .A2(net4182));
 sg13g2_nand2_1 _14787_ (.Y(_05709_),
    .A(net1962),
    .B(net4183));
 sg13g2_o21ai_1 _14788_ (.B1(_05709_),
    .Y(_00723_),
    .A1(net4846),
    .A2(net4183));
 sg13g2_nand2_1 _14789_ (.Y(_05710_),
    .A(net1707),
    .B(net4182));
 sg13g2_o21ai_1 _14790_ (.B1(_05710_),
    .Y(_00724_),
    .A1(net4840),
    .A2(net4182));
 sg13g2_nand2_1 _14791_ (.Y(_05711_),
    .A(net1956),
    .B(net4183));
 sg13g2_o21ai_1 _14792_ (.B1(_05711_),
    .Y(_00725_),
    .A1(net4835),
    .A2(net4183));
 sg13g2_nand2_1 _14793_ (.Y(_05712_),
    .A(net1717),
    .B(net4182));
 sg13g2_o21ai_1 _14794_ (.B1(_05712_),
    .Y(_00726_),
    .A1(net4827),
    .A2(net4182));
 sg13g2_nand2_1 _14795_ (.Y(_05713_),
    .A(net1969),
    .B(net4183));
 sg13g2_o21ai_1 _14796_ (.B1(_05713_),
    .Y(_00727_),
    .A1(net4823),
    .A2(net4183));
 sg13g2_nand2_1 _14797_ (.Y(_05714_),
    .A(net1793),
    .B(net4182));
 sg13g2_o21ai_1 _14798_ (.B1(_05714_),
    .Y(_00728_),
    .A1(net4817),
    .A2(net4182));
 sg13g2_o21ai_1 _14799_ (.B1(_02527_),
    .Y(_05715_),
    .A1(_02526_),
    .A2(_04887_));
 sg13g2_a21o_2 _14800_ (.A2(\m_sys._m_core_io_b_mem_wdata[7] ),
    .A1(net5237),
    .B1(_05152_),
    .X(_05716_));
 sg13g2_nand3_1 _14801_ (.B(net4454),
    .C(_05716_),
    .A(net5145),
    .Y(_05717_));
 sg13g2_o21ai_1 _14802_ (.B1(_05717_),
    .Y(_00729_),
    .A1(_02421_),
    .A2(net4454));
 sg13g2_nor2b_1 _14803_ (.A(net4314),
    .B_N(_05678_),
    .Y(_05718_));
 sg13g2_nor2_1 _14804_ (.A(net2311),
    .B(net4181),
    .Y(_05719_));
 sg13g2_a21oi_1 _14805_ (.A1(net5023),
    .A2(net4181),
    .Y(_00730_),
    .B1(_05719_));
 sg13g2_nor2_1 _14806_ (.A(net2831),
    .B(net4181),
    .Y(_05720_));
 sg13g2_a21oi_1 _14807_ (.A1(net4812),
    .A2(net4181),
    .Y(_00731_),
    .B1(_05720_));
 sg13g2_nor2_1 _14808_ (.A(net2172),
    .B(net4181),
    .Y(_05721_));
 sg13g2_a21oi_1 _14809_ (.A1(net5017),
    .A2(net4181),
    .Y(_00732_),
    .B1(_05721_));
 sg13g2_nor2_1 _14810_ (.A(net2407),
    .B(net4180),
    .Y(_05722_));
 sg13g2_a21oi_1 _14811_ (.A1(net4805),
    .A2(net4180),
    .Y(_00733_),
    .B1(_05722_));
 sg13g2_nor2_1 _14812_ (.A(net2467),
    .B(net4181),
    .Y(_05723_));
 sg13g2_a21oi_1 _14813_ (.A1(net5012),
    .A2(net4181),
    .Y(_00734_),
    .B1(_05723_));
 sg13g2_nor2_1 _14814_ (.A(net2547),
    .B(net4180),
    .Y(_05724_));
 sg13g2_a21oi_1 _14815_ (.A1(net4802),
    .A2(net4180),
    .Y(_00735_),
    .B1(_05724_));
 sg13g2_nor2_1 _14816_ (.A(net2442),
    .B(net4180),
    .Y(_05725_));
 sg13g2_a21oi_1 _14817_ (.A1(net5006),
    .A2(net4180),
    .Y(_00736_),
    .B1(_05725_));
 sg13g2_nor2_1 _14818_ (.A(net2713),
    .B(net4180),
    .Y(_05726_));
 sg13g2_a21oi_1 _14819_ (.A1(net4796),
    .A2(net4180),
    .Y(_00737_),
    .B1(_05726_));
 sg13g2_nand2_1 _14820_ (.Y(_05727_),
    .A(net4320),
    .B(_05410_));
 sg13g2_nand2_1 _14821_ (.Y(_05728_),
    .A(net1702),
    .B(net4179));
 sg13g2_o21ai_1 _14822_ (.B1(_05728_),
    .Y(_00738_),
    .A1(net4853),
    .A2(net4179));
 sg13g2_nand2_1 _14823_ (.Y(_05729_),
    .A(net1727),
    .B(net4179));
 sg13g2_o21ai_1 _14824_ (.B1(_05729_),
    .Y(_00739_),
    .A1(net4848),
    .A2(net4179));
 sg13g2_nand2_1 _14825_ (.Y(_05730_),
    .A(net1880),
    .B(net4178));
 sg13g2_o21ai_1 _14826_ (.B1(_05730_),
    .Y(_00740_),
    .A1(net4842),
    .A2(net4178));
 sg13g2_nand2_1 _14827_ (.Y(_05731_),
    .A(net1773),
    .B(net4178));
 sg13g2_o21ai_1 _14828_ (.B1(_05731_),
    .Y(_00741_),
    .A1(net4838),
    .A2(net4178));
 sg13g2_nand2_1 _14829_ (.Y(_05732_),
    .A(net1733),
    .B(net4178));
 sg13g2_o21ai_1 _14830_ (.B1(_05732_),
    .Y(_00742_),
    .A1(net4831),
    .A2(net4178));
 sg13g2_nand2_1 _14831_ (.Y(_05733_),
    .A(net2095),
    .B(_05727_));
 sg13g2_o21ai_1 _14832_ (.B1(_05733_),
    .Y(_00743_),
    .A1(net4826),
    .A2(net4179));
 sg13g2_nand2_1 _14833_ (.Y(_05734_),
    .A(net1690),
    .B(net4178));
 sg13g2_o21ai_1 _14834_ (.B1(_05734_),
    .Y(_00744_),
    .A1(net4821),
    .A2(net4178));
 sg13g2_nand2_1 _14835_ (.Y(_05735_),
    .A(net1721),
    .B(net4179));
 sg13g2_o21ai_1 _14836_ (.B1(_05735_),
    .Y(_00745_),
    .A1(net4815),
    .A2(net4179));
 sg13g2_nor2b_1 _14837_ (.A(net4314),
    .B_N(_05505_),
    .Y(_05736_));
 sg13g2_nor2_1 _14838_ (.A(net2691),
    .B(_05736_),
    .Y(_05737_));
 sg13g2_a21oi_1 _14839_ (.A1(net5023),
    .A2(net4177),
    .Y(_00746_),
    .B1(_05737_));
 sg13g2_nor2_1 _14840_ (.A(net2440),
    .B(net4177),
    .Y(_05738_));
 sg13g2_a21oi_1 _14841_ (.A1(net4812),
    .A2(net4177),
    .Y(_00747_),
    .B1(_05738_));
 sg13g2_nor2_1 _14842_ (.A(net2189),
    .B(net4177),
    .Y(_05739_));
 sg13g2_a21oi_1 _14843_ (.A1(net5015),
    .A2(net4177),
    .Y(_00748_),
    .B1(_05739_));
 sg13g2_nor2_1 _14844_ (.A(net2156),
    .B(net4176),
    .Y(_05740_));
 sg13g2_a21oi_1 _14845_ (.A1(net4805),
    .A2(net4176),
    .Y(_00749_),
    .B1(_05740_));
 sg13g2_nor2_1 _14846_ (.A(net2147),
    .B(net4177),
    .Y(_05741_));
 sg13g2_a21oi_1 _14847_ (.A1(net5012),
    .A2(net4177),
    .Y(_00750_),
    .B1(_05741_));
 sg13g2_nor2_1 _14848_ (.A(net2205),
    .B(net4176),
    .Y(_05742_));
 sg13g2_a21oi_1 _14849_ (.A1(net4802),
    .A2(net4176),
    .Y(_00751_),
    .B1(_05742_));
 sg13g2_nor2_1 _14850_ (.A(net2793),
    .B(net4176),
    .Y(_05743_));
 sg13g2_a21oi_1 _14851_ (.A1(net5006),
    .A2(net4176),
    .Y(_00752_),
    .B1(_05743_));
 sg13g2_nor2_1 _14852_ (.A(net2489),
    .B(net4176),
    .Y(_05744_));
 sg13g2_a21oi_1 _14853_ (.A1(net4796),
    .A2(net4176),
    .Y(_00753_),
    .B1(_05744_));
 sg13g2_nand2_1 _14854_ (.Y(_05745_),
    .A(net4329),
    .B(_05678_));
 sg13g2_nand2_1 _14855_ (.Y(_05746_),
    .A(net1784),
    .B(net4175));
 sg13g2_o21ai_1 _14856_ (.B1(_05746_),
    .Y(_00754_),
    .A1(net5044),
    .A2(_05745_));
 sg13g2_nand2_1 _14857_ (.Y(_05747_),
    .A(net1972),
    .B(net4175));
 sg13g2_o21ai_1 _14858_ (.B1(_05747_),
    .Y(_00755_),
    .A1(net4874),
    .A2(net4175));
 sg13g2_nand2_1 _14859_ (.Y(_05748_),
    .A(net1738),
    .B(net4174));
 sg13g2_o21ai_1 _14860_ (.B1(_05748_),
    .Y(_00756_),
    .A1(net5039),
    .A2(net4174));
 sg13g2_nand2_1 _14861_ (.Y(_05749_),
    .A(net1967),
    .B(net4174));
 sg13g2_o21ai_1 _14862_ (.B1(_05749_),
    .Y(_00757_),
    .A1(net4872),
    .A2(net4174));
 sg13g2_nand2_1 _14863_ (.Y(_05750_),
    .A(net1900),
    .B(net4174));
 sg13g2_o21ai_1 _14864_ (.B1(_05750_),
    .Y(_00758_),
    .A1(net5033),
    .A2(net4174));
 sg13g2_nand2_1 _14865_ (.Y(_05751_),
    .A(net1933),
    .B(net4174));
 sg13g2_o21ai_1 _14866_ (.B1(_05751_),
    .Y(_00759_),
    .A1(net4867),
    .A2(net4174));
 sg13g2_nand2_1 _14867_ (.Y(_05752_),
    .A(net1806),
    .B(net4175));
 sg13g2_o21ai_1 _14868_ (.B1(_05752_),
    .Y(_00760_),
    .A1(net5026),
    .A2(net4175));
 sg13g2_nand2_1 _14869_ (.Y(_05753_),
    .A(net2152),
    .B(net4175));
 sg13g2_o21ai_1 _14870_ (.B1(_05753_),
    .Y(_00761_),
    .A1(net4861),
    .A2(net4175));
 sg13g2_nor2b_1 _14871_ (.A(net4331),
    .B_N(_05581_),
    .Y(_05754_));
 sg13g2_nor2_1 _14872_ (.A(net2549),
    .B(net4173),
    .Y(_05755_));
 sg13g2_a21oi_1 _14873_ (.A1(net5135),
    .A2(net4173),
    .Y(_00762_),
    .B1(_05755_));
 sg13g2_nor2_1 _14874_ (.A(net2509),
    .B(net4173),
    .Y(_05756_));
 sg13g2_a21oi_1 _14875_ (.A1(net4993),
    .A2(net4173),
    .Y(_00763_),
    .B1(_05756_));
 sg13g2_nor2_1 _14876_ (.A(net2478),
    .B(net4172),
    .Y(_05757_));
 sg13g2_a21oi_1 _14877_ (.A1(net5130),
    .A2(net4172),
    .Y(_00764_),
    .B1(_05757_));
 sg13g2_nor2_1 _14878_ (.A(net2300),
    .B(net4173),
    .Y(_05758_));
 sg13g2_a21oi_1 _14879_ (.A1(net4988),
    .A2(net4173),
    .Y(_00765_),
    .B1(_05758_));
 sg13g2_nor2_1 _14880_ (.A(net2599),
    .B(net4172),
    .Y(_05759_));
 sg13g2_a21oi_1 _14881_ (.A1(net5127),
    .A2(net4172),
    .Y(_00766_),
    .B1(_05759_));
 sg13g2_nor2_1 _14882_ (.A(net2305),
    .B(net4173),
    .Y(_05760_));
 sg13g2_a21oi_1 _14883_ (.A1(net4983),
    .A2(net4173),
    .Y(_00767_),
    .B1(_05760_));
 sg13g2_nor2_1 _14884_ (.A(net2732),
    .B(net4172),
    .Y(_05761_));
 sg13g2_a21oi_1 _14885_ (.A1(net5121),
    .A2(net4172),
    .Y(_00768_),
    .B1(_05761_));
 sg13g2_nor2_1 _14886_ (.A(net2626),
    .B(net4172),
    .Y(_05762_));
 sg13g2_a21oi_1 _14887_ (.A1(net4978),
    .A2(net4172),
    .Y(_00769_),
    .B1(_05762_));
 sg13g2_nand2_1 _14888_ (.Y(_05763_),
    .A(net4322),
    .B(_05371_));
 sg13g2_nand2_1 _14889_ (.Y(_05764_),
    .A(net1809),
    .B(net4170));
 sg13g2_o21ai_1 _14890_ (.B1(_05764_),
    .Y(_00770_),
    .A1(net4855),
    .A2(net4170));
 sg13g2_nand2_1 _14891_ (.Y(_05765_),
    .A(net1899),
    .B(net4171));
 sg13g2_o21ai_1 _14892_ (.B1(_05765_),
    .Y(_00771_),
    .A1(net4851),
    .A2(net4171));
 sg13g2_nand2_1 _14893_ (.Y(_05766_),
    .A(net2108),
    .B(net4170));
 sg13g2_o21ai_1 _14894_ (.B1(_05766_),
    .Y(_00772_),
    .A1(net4844),
    .A2(net4170));
 sg13g2_nand2_1 _14895_ (.Y(_05767_),
    .A(net1693),
    .B(net4171));
 sg13g2_o21ai_1 _14896_ (.B1(_05767_),
    .Y(_00773_),
    .A1(net4839),
    .A2(net4171));
 sg13g2_nand2_1 _14897_ (.Y(_05768_),
    .A(net1814),
    .B(net4170));
 sg13g2_o21ai_1 _14898_ (.B1(_05768_),
    .Y(_00774_),
    .A1(net4833),
    .A2(net4170));
 sg13g2_nand2_1 _14899_ (.Y(_05769_),
    .A(net1756),
    .B(net4171));
 sg13g2_o21ai_1 _14900_ (.B1(_05769_),
    .Y(_00775_),
    .A1(net4829),
    .A2(net4171));
 sg13g2_nand2_1 _14901_ (.Y(_05770_),
    .A(net1740),
    .B(net4171));
 sg13g2_o21ai_1 _14902_ (.B1(_05770_),
    .Y(_00776_),
    .A1(net4822),
    .A2(net4171));
 sg13g2_nand2_1 _14903_ (.Y(_05771_),
    .A(net1893),
    .B(net4170));
 sg13g2_o21ai_1 _14904_ (.B1(_05771_),
    .Y(_00777_),
    .A1(net4816),
    .A2(net4170));
 sg13g2_nor2_1 _14905_ (.A(net2567),
    .B(_04887_),
    .Y(_05772_));
 sg13g2_o21ai_1 _14906_ (.B1(net5385),
    .Y(_00778_),
    .A1(net3207),
    .A2(_05772_));
 sg13g2_nand2b_1 _14907_ (.Y(_05773_),
    .B(_02671_),
    .A_N(_05106_));
 sg13g2_nor2_2 _14908_ (.A(net4597),
    .B(net4449),
    .Y(_05774_));
 sg13g2_nor2b_1 _14909_ (.A(net4315),
    .B_N(_05774_),
    .Y(_05775_));
 sg13g2_nor2_1 _14910_ (.A(net2584),
    .B(net4168),
    .Y(_05776_));
 sg13g2_a21oi_1 _14911_ (.A1(net5024),
    .A2(net4168),
    .Y(_00779_),
    .B1(_05776_));
 sg13g2_nor2_1 _14912_ (.A(net2757),
    .B(net4168),
    .Y(_05777_));
 sg13g2_a21oi_1 _14913_ (.A1(net4813),
    .A2(net4168),
    .Y(_00780_),
    .B1(_05777_));
 sg13g2_nor2_1 _14914_ (.A(net2558),
    .B(net4169),
    .Y(_05778_));
 sg13g2_a21oi_1 _14915_ (.A1(net5019),
    .A2(net4169),
    .Y(_00781_),
    .B1(_05778_));
 sg13g2_nor2_1 _14916_ (.A(net2538),
    .B(net4169),
    .Y(_05779_));
 sg13g2_a21oi_1 _14917_ (.A1(_05141_),
    .A2(net4169),
    .Y(_00782_),
    .B1(_05779_));
 sg13g2_nor2_1 _14918_ (.A(net2591),
    .B(net4168),
    .Y(_05780_));
 sg13g2_a21oi_1 _14919_ (.A1(net5012),
    .A2(net4168),
    .Y(_00783_),
    .B1(_05780_));
 sg13g2_nor2_1 _14920_ (.A(net2201),
    .B(net4169),
    .Y(_05781_));
 sg13g2_a21oi_1 _14921_ (.A1(net4803),
    .A2(net4169),
    .Y(_00784_),
    .B1(_05781_));
 sg13g2_nor2_1 _14922_ (.A(net2853),
    .B(net4169),
    .Y(_05782_));
 sg13g2_a21oi_1 _14923_ (.A1(net5008),
    .A2(net4169),
    .Y(_00785_),
    .B1(_05782_));
 sg13g2_nor2_1 _14924_ (.A(net2187),
    .B(net4168),
    .Y(_05783_));
 sg13g2_a21oi_1 _14925_ (.A1(net4797),
    .A2(net4168),
    .Y(_00786_),
    .B1(_05783_));
 sg13g2_nand2_2 _14926_ (.Y(_05784_),
    .A(net4322),
    .B(_05581_));
 sg13g2_nand2_1 _14927_ (.Y(_05785_),
    .A(net1776),
    .B(net4167));
 sg13g2_o21ai_1 _14928_ (.B1(_05785_),
    .Y(_00787_),
    .A1(net4858),
    .A2(net4167));
 sg13g2_nand2_1 _14929_ (.Y(_05786_),
    .A(net1672),
    .B(net4166));
 sg13g2_o21ai_1 _14930_ (.B1(_05786_),
    .Y(_00788_),
    .A1(net4851),
    .A2(net4166));
 sg13g2_nand2_1 _14931_ (.Y(_05787_),
    .A(net1937),
    .B(_05784_));
 sg13g2_o21ai_1 _14932_ (.B1(_05787_),
    .Y(_00789_),
    .A1(net4845),
    .A2(net4166));
 sg13g2_nand2_1 _14933_ (.Y(_05788_),
    .A(net1961),
    .B(net4166));
 sg13g2_o21ai_1 _14934_ (.B1(_05788_),
    .Y(_00790_),
    .A1(net4841),
    .A2(net4166));
 sg13g2_nand2_1 _14935_ (.Y(_05789_),
    .A(net2016),
    .B(net4167));
 sg13g2_o21ai_1 _14936_ (.B1(_05789_),
    .Y(_00791_),
    .A1(net4833),
    .A2(net4167));
 sg13g2_nand2_1 _14937_ (.Y(_05790_),
    .A(net2005),
    .B(net4166));
 sg13g2_o21ai_1 _14938_ (.B1(_05790_),
    .Y(_00792_),
    .A1(net4829),
    .A2(net4166));
 sg13g2_nand2_1 _14939_ (.Y(_05791_),
    .A(net2125),
    .B(net4167));
 sg13g2_o21ai_1 _14940_ (.B1(_05791_),
    .Y(_00793_),
    .A1(net4820),
    .A2(net4167));
 sg13g2_nand2_1 _14941_ (.Y(_05792_),
    .A(net1888),
    .B(net4166));
 sg13g2_o21ai_1 _14942_ (.B1(_05792_),
    .Y(_00794_),
    .A1(net4819),
    .A2(net4167));
 sg13g2_nor2b_1 _14943_ (.A(net4334),
    .B_N(_05371_),
    .Y(_05793_));
 sg13g2_nor2_1 _14944_ (.A(net2505),
    .B(net4164),
    .Y(_05794_));
 sg13g2_a21oi_1 _14945_ (.A1(net5139),
    .A2(net4164),
    .Y(_00795_),
    .B1(_05794_));
 sg13g2_nor2_1 _14946_ (.A(net2815),
    .B(net4164),
    .Y(_05795_));
 sg13g2_a21oi_1 _14947_ (.A1(net4996),
    .A2(net4164),
    .Y(_00796_),
    .B1(_05795_));
 sg13g2_nor2_1 _14948_ (.A(net2788),
    .B(net4165),
    .Y(_05796_));
 sg13g2_a21oi_1 _14949_ (.A1(net5134),
    .A2(net4165),
    .Y(_00797_),
    .B1(_05796_));
 sg13g2_nor2_1 _14950_ (.A(net2436),
    .B(net4164),
    .Y(_05797_));
 sg13g2_a21oi_1 _14951_ (.A1(net4992),
    .A2(net4164),
    .Y(_00798_),
    .B1(_05797_));
 sg13g2_nor2_1 _14952_ (.A(net2404),
    .B(net4165),
    .Y(_05798_));
 sg13g2_a21oi_1 _14953_ (.A1(net5129),
    .A2(net4165),
    .Y(_00799_),
    .B1(_05798_));
 sg13g2_nor2_1 _14954_ (.A(net2279),
    .B(net4164),
    .Y(_05799_));
 sg13g2_a21oi_1 _14955_ (.A1(net4985),
    .A2(net4164),
    .Y(_00800_),
    .B1(_05799_));
 sg13g2_nor2_1 _14956_ (.A(net2690),
    .B(net4165),
    .Y(_05800_));
 sg13g2_a21oi_1 _14957_ (.A1(net5123),
    .A2(net4165),
    .Y(_00801_),
    .B1(_05800_));
 sg13g2_nor2_1 _14958_ (.A(net2354),
    .B(net4165),
    .Y(_05801_));
 sg13g2_a21oi_1 _14959_ (.A1(net4982),
    .A2(net4165),
    .Y(_00802_),
    .B1(_05801_));
 sg13g2_nor2_2 _14960_ (.A(net4551),
    .B(net4448),
    .Y(_05802_));
 sg13g2_nor2b_1 _14961_ (.A(net4314),
    .B_N(_05802_),
    .Y(_05803_));
 sg13g2_nor2_1 _14962_ (.A(net2435),
    .B(net4162),
    .Y(_05804_));
 sg13g2_a21oi_1 _14963_ (.A1(net5024),
    .A2(net4162),
    .Y(_00803_),
    .B1(_05804_));
 sg13g2_nor2_1 _14964_ (.A(net2177),
    .B(net4162),
    .Y(_05805_));
 sg13g2_a21oi_1 _14965_ (.A1(net4813),
    .A2(net4162),
    .Y(_00804_),
    .B1(_05805_));
 sg13g2_nor2_1 _14966_ (.A(net2610),
    .B(net4163),
    .Y(_05806_));
 sg13g2_a21oi_1 _14967_ (.A1(net5019),
    .A2(net4163),
    .Y(_00805_),
    .B1(_05806_));
 sg13g2_nor2_1 _14968_ (.A(net2666),
    .B(net4163),
    .Y(_05807_));
 sg13g2_a21oi_1 _14969_ (.A1(net4809),
    .A2(net4163),
    .Y(_00806_),
    .B1(_05807_));
 sg13g2_nor2_1 _14970_ (.A(net2154),
    .B(net4162),
    .Y(_05808_));
 sg13g2_a21oi_1 _14971_ (.A1(net5013),
    .A2(net4162),
    .Y(_00807_),
    .B1(_05808_));
 sg13g2_nor2_1 _14972_ (.A(net2650),
    .B(net4163),
    .Y(_05809_));
 sg13g2_a21oi_1 _14973_ (.A1(net4803),
    .A2(net4163),
    .Y(_00808_),
    .B1(_05809_));
 sg13g2_nor2_1 _14974_ (.A(net2202),
    .B(net4163),
    .Y(_05810_));
 sg13g2_a21oi_1 _14975_ (.A1(net5008),
    .A2(net4163),
    .Y(_00809_),
    .B1(_05810_));
 sg13g2_nor2_1 _14976_ (.A(net2438),
    .B(net4162),
    .Y(_05811_));
 sg13g2_a21oi_1 _14977_ (.A1(net4796),
    .A2(net4162),
    .Y(_00810_),
    .B1(_05811_));
 sg13g2_nor2b_1 _14978_ (.A(net4335),
    .B_N(_05439_),
    .Y(_05812_));
 sg13g2_nor2_1 _14979_ (.A(net2730),
    .B(net4160),
    .Y(_05813_));
 sg13g2_a21oi_1 _14980_ (.A1(net5138),
    .A2(net4161),
    .Y(_00811_),
    .B1(_05813_));
 sg13g2_nor2_1 _14981_ (.A(net2673),
    .B(net4160),
    .Y(_05814_));
 sg13g2_a21oi_1 _14982_ (.A1(net4995),
    .A2(net4160),
    .Y(_00812_),
    .B1(_05814_));
 sg13g2_nor2_1 _14983_ (.A(net2662),
    .B(_05812_),
    .Y(_05815_));
 sg13g2_a21oi_1 _14984_ (.A1(net5134),
    .A2(net4160),
    .Y(_00813_),
    .B1(_05815_));
 sg13g2_nor2_1 _14985_ (.A(net2158),
    .B(net4161),
    .Y(_05816_));
 sg13g2_a21oi_1 _14986_ (.A1(net4991),
    .A2(net4161),
    .Y(_00814_),
    .B1(_05816_));
 sg13g2_nor2_1 _14987_ (.A(net2197),
    .B(net4161),
    .Y(_05817_));
 sg13g2_a21oi_1 _14988_ (.A1(net5126),
    .A2(net4161),
    .Y(_00815_),
    .B1(_05817_));
 sg13g2_nor2_1 _14989_ (.A(net2336),
    .B(net4160),
    .Y(_05818_));
 sg13g2_a21oi_1 _14990_ (.A1(net4985),
    .A2(net4160),
    .Y(_00816_),
    .B1(_05818_));
 sg13g2_nor2_1 _14991_ (.A(net2597),
    .B(net4161),
    .Y(_05819_));
 sg13g2_a21oi_1 _14992_ (.A1(net5120),
    .A2(net4161),
    .Y(_00817_),
    .B1(_05819_));
 sg13g2_nor2_1 _14993_ (.A(net2649),
    .B(net4160),
    .Y(_05820_));
 sg13g2_a21oi_1 _14994_ (.A1(net4982),
    .A2(net4160),
    .Y(_00818_),
    .B1(_05820_));
 sg13g2_nand2_1 _14995_ (.Y(_05821_),
    .A(net4327),
    .B(_05581_));
 sg13g2_nand2_1 _14996_ (.Y(_05822_),
    .A(net1761),
    .B(net4158));
 sg13g2_o21ai_1 _14997_ (.B1(_05822_),
    .Y(_00819_),
    .A1(net5041),
    .A2(net4158));
 sg13g2_nand2_1 _14998_ (.Y(_05823_),
    .A(net1744),
    .B(net4159));
 sg13g2_o21ai_1 _14999_ (.B1(_05823_),
    .Y(_00820_),
    .A1(net4876),
    .A2(net4159));
 sg13g2_nand2_1 _15000_ (.Y(_05824_),
    .A(net1805),
    .B(net4158));
 sg13g2_o21ai_1 _15001_ (.B1(_05824_),
    .Y(_00821_),
    .A1(net5037),
    .A2(net4158));
 sg13g2_nand2_1 _15002_ (.Y(_05825_),
    .A(net1722),
    .B(net4159));
 sg13g2_o21ai_1 _15003_ (.B1(_05825_),
    .Y(_00822_),
    .A1(net4873),
    .A2(net4159));
 sg13g2_nand2_1 _15004_ (.Y(_05826_),
    .A(net1909),
    .B(net4158));
 sg13g2_o21ai_1 _15005_ (.B1(_05826_),
    .Y(_00823_),
    .A1(net5030),
    .A2(net4158));
 sg13g2_nand2_1 _15006_ (.Y(_05827_),
    .A(net1723),
    .B(net4158));
 sg13g2_o21ai_1 _15007_ (.B1(_05827_),
    .Y(_00824_),
    .A1(net4865),
    .A2(net4158));
 sg13g2_nand2_1 _15008_ (.Y(_05828_),
    .A(net1936),
    .B(net4159));
 sg13g2_o21ai_1 _15009_ (.B1(_05828_),
    .Y(_00825_),
    .A1(net5028),
    .A2(net4159));
 sg13g2_nand2_1 _15010_ (.Y(_05829_),
    .A(net1705),
    .B(net4159));
 sg13g2_o21ai_1 _15011_ (.B1(_05829_),
    .Y(_00826_),
    .A1(net4862),
    .A2(net4159));
 sg13g2_nand2_1 _15012_ (.Y(_05830_),
    .A(net4330),
    .B(_05391_));
 sg13g2_nand2_1 _15013_ (.Y(_05831_),
    .A(net2087),
    .B(net4155));
 sg13g2_o21ai_1 _15014_ (.B1(_05831_),
    .Y(_00827_),
    .A1(net5045),
    .A2(net4155));
 sg13g2_nand2_1 _15015_ (.Y(_05832_),
    .A(net1885),
    .B(net4155));
 sg13g2_o21ai_1 _15016_ (.B1(_05832_),
    .Y(_00828_),
    .A1(net4874),
    .A2(net4155));
 sg13g2_nand2_1 _15017_ (.Y(_05833_),
    .A(net1861),
    .B(net4156));
 sg13g2_o21ai_1 _15018_ (.B1(_05833_),
    .Y(_00829_),
    .A1(net5040),
    .A2(net4156));
 sg13g2_nand2_1 _15019_ (.Y(_05834_),
    .A(net1975),
    .B(net4157));
 sg13g2_o21ai_1 _15020_ (.B1(_05834_),
    .Y(_00830_),
    .A1(net4870),
    .A2(net4157));
 sg13g2_nand2_1 _15021_ (.Y(_05835_),
    .A(net1755),
    .B(net4157));
 sg13g2_o21ai_1 _15022_ (.B1(_05835_),
    .Y(_00831_),
    .A1(net5031),
    .A2(net4157));
 sg13g2_nand2_1 _15023_ (.Y(_05836_),
    .A(net1912),
    .B(net4155));
 sg13g2_o21ai_1 _15024_ (.B1(_05836_),
    .Y(_00832_),
    .A1(net4868),
    .A2(net4155));
 sg13g2_nand2_1 _15025_ (.Y(_05837_),
    .A(net1714),
    .B(net4156));
 sg13g2_o21ai_1 _15026_ (.B1(_05837_),
    .Y(_00833_),
    .A1(net5027),
    .A2(net4156));
 sg13g2_nand2_1 _15027_ (.Y(_05838_),
    .A(net1662),
    .B(net4155));
 sg13g2_o21ai_1 _15028_ (.B1(_05838_),
    .Y(_00834_),
    .A1(net4859),
    .A2(net4155));
 sg13g2_nand2_1 _15029_ (.Y(_05839_),
    .A(net4321),
    .B(_05439_));
 sg13g2_nand2_1 _15030_ (.Y(_05840_),
    .A(net1856),
    .B(net4154));
 sg13g2_o21ai_1 _15031_ (.B1(_05840_),
    .Y(_00835_),
    .A1(net4854),
    .A2(net4154));
 sg13g2_nand2_1 _15032_ (.Y(_05841_),
    .A(net1708),
    .B(net4153));
 sg13g2_o21ai_1 _15033_ (.B1(_05841_),
    .Y(_00836_),
    .A1(net4847),
    .A2(net4153));
 sg13g2_nand2_1 _15034_ (.Y(_05842_),
    .A(net1677),
    .B(net4154));
 sg13g2_o21ai_1 _15035_ (.B1(_05842_),
    .Y(_00837_),
    .A1(net4843),
    .A2(net4154));
 sg13g2_nand2_1 _15036_ (.Y(_05843_),
    .A(net1670),
    .B(net4154));
 sg13g2_o21ai_1 _15037_ (.B1(_05843_),
    .Y(_00838_),
    .A1(net4837),
    .A2(net4154));
 sg13g2_nand2_1 _15038_ (.Y(_05844_),
    .A(net1731),
    .B(net4153));
 sg13g2_o21ai_1 _15039_ (.B1(_05844_),
    .Y(_00839_),
    .A1(net4831),
    .A2(net4153));
 sg13g2_nand2_1 _15040_ (.Y(_05845_),
    .A(net1674),
    .B(net4154));
 sg13g2_o21ai_1 _15041_ (.B1(_05845_),
    .Y(_00840_),
    .A1(net4825),
    .A2(net4154));
 sg13g2_nand2_1 _15042_ (.Y(_05846_),
    .A(net1920),
    .B(net4153));
 sg13g2_o21ai_1 _15043_ (.B1(_05846_),
    .Y(_00841_),
    .A1(net4821),
    .A2(net4153));
 sg13g2_nand2_1 _15044_ (.Y(_05847_),
    .A(net1675),
    .B(net4153));
 sg13g2_o21ai_1 _15045_ (.B1(_05847_),
    .Y(_00842_),
    .A1(net4816),
    .A2(net4153));
 sg13g2_nor2_2 _15046_ (.A(net4643),
    .B(net4448),
    .Y(_05848_));
 sg13g2_nor2b_1 _15047_ (.A(net4314),
    .B_N(_05848_),
    .Y(_05849_));
 sg13g2_nor2_1 _15048_ (.A(net2306),
    .B(net4151),
    .Y(_05850_));
 sg13g2_a21oi_1 _15049_ (.A1(net5024),
    .A2(net4151),
    .Y(_00843_),
    .B1(_05850_));
 sg13g2_nor2_1 _15050_ (.A(net2411),
    .B(net4152),
    .Y(_05851_));
 sg13g2_a21oi_1 _15051_ (.A1(net4812),
    .A2(net4152),
    .Y(_00844_),
    .B1(_05851_));
 sg13g2_nor2_1 _15052_ (.A(net2431),
    .B(net4151),
    .Y(_05852_));
 sg13g2_a21oi_1 _15053_ (.A1(net5019),
    .A2(_05849_),
    .Y(_00845_),
    .B1(_05852_));
 sg13g2_nor2_1 _15054_ (.A(net2272),
    .B(net4151),
    .Y(_05853_));
 sg13g2_a21oi_1 _15055_ (.A1(net4809),
    .A2(net4151),
    .Y(_00846_),
    .B1(_05853_));
 sg13g2_nor2_1 _15056_ (.A(net2398),
    .B(net4152),
    .Y(_05854_));
 sg13g2_a21oi_1 _15057_ (.A1(net5012),
    .A2(net4152),
    .Y(_00847_),
    .B1(_05854_));
 sg13g2_nor2_1 _15058_ (.A(net2396),
    .B(net4151),
    .Y(_05855_));
 sg13g2_a21oi_1 _15059_ (.A1(net4803),
    .A2(net4151),
    .Y(_00848_),
    .B1(_05855_));
 sg13g2_nor2_1 _15060_ (.A(net2493),
    .B(net4151),
    .Y(_05856_));
 sg13g2_a21oi_1 _15061_ (.A1(net5007),
    .A2(net4152),
    .Y(_00849_),
    .B1(_05856_));
 sg13g2_nor2_1 _15062_ (.A(net2290),
    .B(net4152),
    .Y(_05857_));
 sg13g2_a21oi_1 _15063_ (.A1(net4796),
    .A2(net4152),
    .Y(_00850_),
    .B1(_05857_));
 sg13g2_nand2_1 _15064_ (.Y(_05858_),
    .A(net4326),
    .B(_05439_));
 sg13g2_nand2_1 _15065_ (.Y(_05859_),
    .A(net1873),
    .B(net4149));
 sg13g2_o21ai_1 _15066_ (.B1(_05859_),
    .Y(_00851_),
    .A1(net5042),
    .A2(net4149));
 sg13g2_nand2_1 _15067_ (.Y(_05860_),
    .A(net1692),
    .B(_05858_));
 sg13g2_o21ai_1 _15068_ (.B1(_05860_),
    .Y(_00852_),
    .A1(net4877),
    .A2(net4150));
 sg13g2_nand2_1 _15069_ (.Y(_05861_),
    .A(net1794),
    .B(net4150));
 sg13g2_o21ai_1 _15070_ (.B1(_05861_),
    .Y(_00853_),
    .A1(net5035),
    .A2(net4150));
 sg13g2_nand2_1 _15071_ (.Y(_05862_),
    .A(net1815),
    .B(net4150));
 sg13g2_o21ai_1 _15072_ (.B1(_05862_),
    .Y(_00854_),
    .A1(net4869),
    .A2(net4150));
 sg13g2_nand2_1 _15073_ (.Y(_05863_),
    .A(net1986),
    .B(net4149));
 sg13g2_o21ai_1 _15074_ (.B1(_05863_),
    .Y(_00855_),
    .A1(net5031),
    .A2(net4149));
 sg13g2_nand2_1 _15075_ (.Y(_05864_),
    .A(net1741),
    .B(net4150));
 sg13g2_o21ai_1 _15076_ (.B1(_05864_),
    .Y(_00856_),
    .A1(net4864),
    .A2(net4150));
 sg13g2_nand2_1 _15077_ (.Y(_05865_),
    .A(net1700),
    .B(net4149));
 sg13g2_o21ai_1 _15078_ (.B1(_05865_),
    .Y(_00857_),
    .A1(net5029),
    .A2(net4149));
 sg13g2_nand2_1 _15079_ (.Y(_05866_),
    .A(net2046),
    .B(net4149));
 sg13g2_o21ai_1 _15080_ (.B1(_05866_),
    .Y(_00858_),
    .A1(net4863),
    .A2(net4149));
 sg13g2_nor2_2 _15081_ (.A(net4597),
    .B(net4474),
    .Y(_05867_));
 sg13g2_nor2b_1 _15082_ (.A(net4331),
    .B_N(_05867_),
    .Y(_05868_));
 sg13g2_nor2_1 _15083_ (.A(net2355),
    .B(net4148),
    .Y(_05869_));
 sg13g2_a21oi_1 _15084_ (.A1(net5135),
    .A2(net4148),
    .Y(_00859_),
    .B1(_05869_));
 sg13g2_nor2_1 _15085_ (.A(net2605),
    .B(net4148),
    .Y(_05870_));
 sg13g2_a21oi_1 _15086_ (.A1(net4993),
    .A2(net4148),
    .Y(_00860_),
    .B1(_05870_));
 sg13g2_nor2_1 _15087_ (.A(net2372),
    .B(net4147),
    .Y(_05871_));
 sg13g2_a21oi_1 _15088_ (.A1(net5130),
    .A2(net4147),
    .Y(_00861_),
    .B1(_05871_));
 sg13g2_nor2_1 _15089_ (.A(net2373),
    .B(net4148),
    .Y(_05872_));
 sg13g2_a21oi_1 _15090_ (.A1(net4988),
    .A2(net4148),
    .Y(_00862_),
    .B1(_05872_));
 sg13g2_nor2_1 _15091_ (.A(net2343),
    .B(net4147),
    .Y(_05873_));
 sg13g2_a21oi_1 _15092_ (.A1(net5127),
    .A2(net4147),
    .Y(_00863_),
    .B1(_05873_));
 sg13g2_nor2_1 _15093_ (.A(net2367),
    .B(net4148),
    .Y(_05874_));
 sg13g2_a21oi_1 _15094_ (.A1(net4983),
    .A2(net4148),
    .Y(_00864_),
    .B1(_05874_));
 sg13g2_nor2_1 _15095_ (.A(net2166),
    .B(net4147),
    .Y(_05875_));
 sg13g2_a21oi_1 _15096_ (.A1(net5121),
    .A2(net4147),
    .Y(_00865_),
    .B1(_05875_));
 sg13g2_nor2_1 _15097_ (.A(net2361),
    .B(net4147),
    .Y(_05876_));
 sg13g2_a21oi_1 _15098_ (.A1(net4978),
    .A2(net4147),
    .Y(_00866_),
    .B1(_05876_));
 sg13g2_nand2_1 _15099_ (.Y(_05877_),
    .A(net4322),
    .B(_05391_));
 sg13g2_nand2_1 _15100_ (.Y(_05878_),
    .A(net2037),
    .B(net4145));
 sg13g2_o21ai_1 _15101_ (.B1(_05878_),
    .Y(_00867_),
    .A1(net4855),
    .A2(net4145));
 sg13g2_nand2_1 _15102_ (.Y(_05879_),
    .A(net1772),
    .B(net4146));
 sg13g2_o21ai_1 _15103_ (.B1(_05879_),
    .Y(_00868_),
    .A1(net4851),
    .A2(net4146));
 sg13g2_nand2_1 _15104_ (.Y(_05880_),
    .A(net2150),
    .B(net4146));
 sg13g2_o21ai_1 _15105_ (.B1(_05880_),
    .Y(_00869_),
    .A1(net4844),
    .A2(net4146));
 sg13g2_nand2_1 _15106_ (.Y(_05881_),
    .A(net1746),
    .B(_05877_));
 sg13g2_o21ai_1 _15107_ (.B1(_05881_),
    .Y(_00870_),
    .A1(net4839),
    .A2(net4146));
 sg13g2_nand2_1 _15108_ (.Y(_05882_),
    .A(net2061),
    .B(net4145));
 sg13g2_o21ai_1 _15109_ (.B1(_05882_),
    .Y(_00871_),
    .A1(net4833),
    .A2(net4145));
 sg13g2_nand2_1 _15110_ (.Y(_05883_),
    .A(net1911),
    .B(net4145));
 sg13g2_o21ai_1 _15111_ (.B1(_05883_),
    .Y(_00872_),
    .A1(net4829),
    .A2(net4145));
 sg13g2_nand2_1 _15112_ (.Y(_05884_),
    .A(net2071),
    .B(net4146));
 sg13g2_o21ai_1 _15113_ (.B1(_05884_),
    .Y(_00873_),
    .A1(net4822),
    .A2(net4146));
 sg13g2_nand2_1 _15114_ (.Y(_05885_),
    .A(net1824),
    .B(net4145));
 sg13g2_o21ai_1 _15115_ (.B1(_05885_),
    .Y(_00874_),
    .A1(_04978_),
    .A2(net4145));
 sg13g2_nor2_2 _15116_ (.A(net4506),
    .B(net4457),
    .Y(_05886_));
 sg13g2_nor2b_1 _15117_ (.A(net4332),
    .B_N(_05886_),
    .Y(_05887_));
 sg13g2_nor2_1 _15118_ (.A(net2553),
    .B(net4143),
    .Y(_05888_));
 sg13g2_a21oi_1 _15119_ (.A1(net5137),
    .A2(net4143),
    .Y(_00875_),
    .B1(_05888_));
 sg13g2_nor2_1 _15120_ (.A(net2571),
    .B(net4144),
    .Y(_05889_));
 sg13g2_a21oi_1 _15121_ (.A1(net4995),
    .A2(net4144),
    .Y(_00876_),
    .B1(_05889_));
 sg13g2_nor2_1 _15122_ (.A(net2320),
    .B(net4143),
    .Y(_05890_));
 sg13g2_a21oi_1 _15123_ (.A1(net5131),
    .A2(net4143),
    .Y(_00877_),
    .B1(_05890_));
 sg13g2_nor2_1 _15124_ (.A(net2689),
    .B(net4144),
    .Y(_05891_));
 sg13g2_a21oi_1 _15125_ (.A1(net4990),
    .A2(net4144),
    .Y(_00878_),
    .B1(_05891_));
 sg13g2_nor2_1 _15126_ (.A(net2767),
    .B(net4144),
    .Y(_05892_));
 sg13g2_a21oi_1 _15127_ (.A1(net5128),
    .A2(net4144),
    .Y(_00879_),
    .B1(_05892_));
 sg13g2_nor2_1 _15128_ (.A(net2601),
    .B(net4143),
    .Y(_05893_));
 sg13g2_a21oi_1 _15129_ (.A1(net4986),
    .A2(net4143),
    .Y(_00880_),
    .B1(_05893_));
 sg13g2_nor2_1 _15130_ (.A(net2615),
    .B(net4144),
    .Y(_05894_));
 sg13g2_a21oi_1 _15131_ (.A1(net5122),
    .A2(net4144),
    .Y(_00881_),
    .B1(_05894_));
 sg13g2_nor2_1 _15132_ (.A(net2776),
    .B(net4143),
    .Y(_05895_));
 sg13g2_a21oi_1 _15133_ (.A1(net4979),
    .A2(net4143),
    .Y(_00882_),
    .B1(_05895_));
 sg13g2_nand2_1 _15134_ (.Y(_05896_),
    .A(net4324),
    .B(_05886_));
 sg13g2_nand2_1 _15135_ (.Y(_05897_),
    .A(net1709),
    .B(net4142));
 sg13g2_o21ai_1 _15136_ (.B1(_05897_),
    .Y(_00883_),
    .A1(net4856),
    .A2(net4142));
 sg13g2_nand2_1 _15137_ (.Y(_05898_),
    .A(net2009),
    .B(net4142));
 sg13g2_o21ai_1 _15138_ (.B1(_05898_),
    .Y(_00884_),
    .A1(net4849),
    .A2(net4142));
 sg13g2_nand2_1 _15139_ (.Y(_05899_),
    .A(net1831),
    .B(net4142));
 sg13g2_o21ai_1 _15140_ (.B1(_05899_),
    .Y(_00885_),
    .A1(net4845),
    .A2(net4142));
 sg13g2_nand2_1 _15141_ (.Y(_05900_),
    .A(net1926),
    .B(net4142));
 sg13g2_o21ai_1 _15142_ (.B1(_05900_),
    .Y(_00886_),
    .A1(net4840),
    .A2(net4142));
 sg13g2_nand2_1 _15143_ (.Y(_05901_),
    .A(net1997),
    .B(net4141));
 sg13g2_o21ai_1 _15144_ (.B1(_05901_),
    .Y(_00887_),
    .A1(net4834),
    .A2(net4141));
 sg13g2_nand2_1 _15145_ (.Y(_05902_),
    .A(net2117),
    .B(net4141));
 sg13g2_o21ai_1 _15146_ (.B1(_05902_),
    .Y(_00888_),
    .A1(net4828),
    .A2(net4141));
 sg13g2_nand2_1 _15147_ (.Y(_05903_),
    .A(net1851),
    .B(net4141));
 sg13g2_o21ai_1 _15148_ (.B1(_05903_),
    .Y(_00889_),
    .A1(net4822),
    .A2(net4141));
 sg13g2_nand2_1 _15149_ (.Y(_05904_),
    .A(net1810),
    .B(net4141));
 sg13g2_o21ai_1 _15150_ (.B1(_05904_),
    .Y(_00890_),
    .A1(net4817),
    .A2(net4141));
 sg13g2_nand2_1 _15151_ (.Y(_05905_),
    .A(net4328),
    .B(_05886_));
 sg13g2_nand2_1 _15152_ (.Y(_05906_),
    .A(net2105),
    .B(_05905_));
 sg13g2_o21ai_1 _15153_ (.B1(_05906_),
    .Y(_00891_),
    .A1(net5043),
    .A2(net4140));
 sg13g2_nand2_1 _15154_ (.Y(_05907_),
    .A(net1853),
    .B(net4140));
 sg13g2_o21ai_1 _15155_ (.B1(_05907_),
    .Y(_00892_),
    .A1(_04936_),
    .A2(net4140));
 sg13g2_nand2_1 _15156_ (.Y(_05908_),
    .A(net1947),
    .B(net4139));
 sg13g2_o21ai_1 _15157_ (.B1(_05908_),
    .Y(_00893_),
    .A1(net5038),
    .A2(net4139));
 sg13g2_nand2_1 _15158_ (.Y(_05909_),
    .A(net1930),
    .B(net4139));
 sg13g2_o21ai_1 _15159_ (.B1(_05909_),
    .Y(_00894_),
    .A1(net4871),
    .A2(net4139));
 sg13g2_nand2_1 _15160_ (.Y(_05910_),
    .A(net2029),
    .B(net4139));
 sg13g2_o21ai_1 _15161_ (.B1(_05910_),
    .Y(_00895_),
    .A1(net5032),
    .A2(net4139));
 sg13g2_nand2_1 _15162_ (.Y(_05911_),
    .A(net2055),
    .B(net4139));
 sg13g2_o21ai_1 _15163_ (.B1(_05911_),
    .Y(_00896_),
    .A1(net4866),
    .A2(net4139));
 sg13g2_nand2_1 _15164_ (.Y(_05912_),
    .A(net1977),
    .B(net4140));
 sg13g2_o21ai_1 _15165_ (.B1(_05912_),
    .Y(_00897_),
    .A1(_04946_),
    .A2(net4140));
 sg13g2_nand2_1 _15166_ (.Y(_05913_),
    .A(net1791),
    .B(net4140));
 sg13g2_o21ai_1 _15167_ (.B1(_05913_),
    .Y(_00898_),
    .A1(net4859),
    .A2(net4140));
 sg13g2_nor2b_1 _15168_ (.A(net4334),
    .B_N(_05562_),
    .Y(_05914_));
 sg13g2_nor2_1 _15169_ (.A(net2280),
    .B(net4138),
    .Y(_05915_));
 sg13g2_a21oi_1 _15170_ (.A1(net5137),
    .A2(net4138),
    .Y(_00899_),
    .B1(_05915_));
 sg13g2_nor2_1 _15171_ (.A(net2516),
    .B(net4137),
    .Y(_05916_));
 sg13g2_a21oi_1 _15172_ (.A1(net4995),
    .A2(net4137),
    .Y(_00900_),
    .B1(_05916_));
 sg13g2_nor2_1 _15173_ (.A(net2244),
    .B(net4138),
    .Y(_05917_));
 sg13g2_a21oi_1 _15174_ (.A1(net5131),
    .A2(net4138),
    .Y(_00901_),
    .B1(_05917_));
 sg13g2_nor2_1 _15175_ (.A(net2680),
    .B(net4137),
    .Y(_05918_));
 sg13g2_a21oi_1 _15176_ (.A1(net4990),
    .A2(net4137),
    .Y(_00902_),
    .B1(_05918_));
 sg13g2_nor2_1 _15177_ (.A(net2695),
    .B(net4137),
    .Y(_05919_));
 sg13g2_a21oi_1 _15178_ (.A1(net5128),
    .A2(net4137),
    .Y(_00903_),
    .B1(_05919_));
 sg13g2_nor2_1 _15179_ (.A(net2409),
    .B(_05914_),
    .Y(_05920_));
 sg13g2_a21oi_1 _15180_ (.A1(net4986),
    .A2(net4138),
    .Y(_00904_),
    .B1(_05920_));
 sg13g2_nor2_1 _15181_ (.A(net2167),
    .B(net4137),
    .Y(_05921_));
 sg13g2_a21oi_1 _15182_ (.A1(net5122),
    .A2(net4137),
    .Y(_00905_),
    .B1(_05921_));
 sg13g2_nor2_1 _15183_ (.A(net2669),
    .B(net4138),
    .Y(_05922_));
 sg13g2_a21oi_1 _15184_ (.A1(net4979),
    .A2(net4138),
    .Y(_00906_),
    .B1(_05922_));
 sg13g2_nand2_1 _15185_ (.Y(_05923_),
    .A(net4324),
    .B(_05562_));
 sg13g2_nand2_1 _15186_ (.Y(_05924_),
    .A(net1760),
    .B(net4136));
 sg13g2_o21ai_1 _15187_ (.B1(_05924_),
    .Y(_00907_),
    .A1(net4856),
    .A2(net4136));
 sg13g2_nand2_1 _15188_ (.Y(_05925_),
    .A(net2111),
    .B(net4136));
 sg13g2_o21ai_1 _15189_ (.B1(_05925_),
    .Y(_00908_),
    .A1(net4850),
    .A2(net4136));
 sg13g2_nand2_1 _15190_ (.Y(_05926_),
    .A(net1742),
    .B(net4136));
 sg13g2_o21ai_1 _15191_ (.B1(_05926_),
    .Y(_00909_),
    .A1(net4845),
    .A2(net4136));
 sg13g2_nand2_1 _15192_ (.Y(_05927_),
    .A(net1786),
    .B(net4136));
 sg13g2_o21ai_1 _15193_ (.B1(_05927_),
    .Y(_00910_),
    .A1(net4840),
    .A2(net4136));
 sg13g2_nand2_1 _15194_ (.Y(_05928_),
    .A(net1875),
    .B(net4135));
 sg13g2_o21ai_1 _15195_ (.B1(_05928_),
    .Y(_00911_),
    .A1(net4834),
    .A2(net4135));
 sg13g2_nand2_1 _15196_ (.Y(_05929_),
    .A(net1841),
    .B(net4135));
 sg13g2_o21ai_1 _15197_ (.B1(_05929_),
    .Y(_00912_),
    .A1(net4828),
    .A2(net4135));
 sg13g2_nand2_1 _15198_ (.Y(_05930_),
    .A(net1682),
    .B(net4135));
 sg13g2_o21ai_1 _15199_ (.B1(_05930_),
    .Y(_00913_),
    .A1(net4822),
    .A2(net4135));
 sg13g2_nand2_1 _15200_ (.Y(_05931_),
    .A(net2112),
    .B(net4135));
 sg13g2_o21ai_1 _15201_ (.B1(_05931_),
    .Y(_00914_),
    .A1(net4817),
    .A2(net4135));
 sg13g2_nand2_1 _15202_ (.Y(_05932_),
    .A(net4328),
    .B(_05562_));
 sg13g2_nand2_1 _15203_ (.Y(_05933_),
    .A(net1904),
    .B(_05932_));
 sg13g2_o21ai_1 _15204_ (.B1(_05933_),
    .Y(_00915_),
    .A1(net5043),
    .A2(net4134));
 sg13g2_nand2_1 _15205_ (.Y(_05934_),
    .A(net1860),
    .B(net4134));
 sg13g2_o21ai_1 _15206_ (.B1(_05934_),
    .Y(_00916_),
    .A1(net4875),
    .A2(net4134));
 sg13g2_nand2_1 _15207_ (.Y(_05935_),
    .A(net1879),
    .B(net4133));
 sg13g2_o21ai_1 _15208_ (.B1(_05935_),
    .Y(_00917_),
    .A1(net5038),
    .A2(net4133));
 sg13g2_nand2_1 _15209_ (.Y(_05936_),
    .A(net1919),
    .B(net4133));
 sg13g2_o21ai_1 _15210_ (.B1(_05936_),
    .Y(_00918_),
    .A1(net4871),
    .A2(net4133));
 sg13g2_nand2_1 _15211_ (.Y(_05937_),
    .A(net2094),
    .B(net4133));
 sg13g2_o21ai_1 _15212_ (.B1(_05937_),
    .Y(_00919_),
    .A1(net5032),
    .A2(net4133));
 sg13g2_nand2_1 _15213_ (.Y(_05938_),
    .A(net1927),
    .B(net4133));
 sg13g2_o21ai_1 _15214_ (.B1(_05938_),
    .Y(_00920_),
    .A1(net4866),
    .A2(net4133));
 sg13g2_nand2_1 _15215_ (.Y(_05939_),
    .A(net2091),
    .B(net4134));
 sg13g2_o21ai_1 _15216_ (.B1(_05939_),
    .Y(_00921_),
    .A1(net5026),
    .A2(net4134));
 sg13g2_nand2_1 _15217_ (.Y(_05940_),
    .A(net2058),
    .B(net4134));
 sg13g2_o21ai_1 _15218_ (.B1(_05940_),
    .Y(_00922_),
    .A1(net4860),
    .A2(net4134));
 sg13g2_nor2b_1 _15219_ (.A(net4332),
    .B_N(_05668_),
    .Y(_05941_));
 sg13g2_nor2_1 _15220_ (.A(net2842),
    .B(net4131),
    .Y(_05942_));
 sg13g2_a21oi_1 _15221_ (.A1(net5138),
    .A2(net4131),
    .Y(_00923_),
    .B1(_05942_));
 sg13g2_nor2_1 _15222_ (.A(net2526),
    .B(net4131),
    .Y(_05943_));
 sg13g2_a21oi_1 _15223_ (.A1(net4995),
    .A2(net4131),
    .Y(_00924_),
    .B1(_05943_));
 sg13g2_nor2_1 _15224_ (.A(net2644),
    .B(net4132),
    .Y(_05944_));
 sg13g2_a21oi_1 _15225_ (.A1(_02735_),
    .A2(_05941_),
    .Y(_00925_),
    .B1(_05944_));
 sg13g2_nor2_1 _15226_ (.A(net2581),
    .B(net4132),
    .Y(_05945_));
 sg13g2_a21oi_1 _15227_ (.A1(net4991),
    .A2(net4132),
    .Y(_00926_),
    .B1(_05945_));
 sg13g2_nor2_1 _15228_ (.A(net2287),
    .B(net4132),
    .Y(_05946_));
 sg13g2_a21oi_1 _15229_ (.A1(net5125),
    .A2(net4132),
    .Y(_00927_),
    .B1(_05946_));
 sg13g2_nor2_1 _15230_ (.A(net2253),
    .B(net4131),
    .Y(_05947_));
 sg13g2_a21oi_1 _15231_ (.A1(net4985),
    .A2(net4131),
    .Y(_00928_),
    .B1(_05947_));
 sg13g2_nor2_1 _15232_ (.A(net2495),
    .B(net4132),
    .Y(_05948_));
 sg13g2_a21oi_1 _15233_ (.A1(net5120),
    .A2(net4132),
    .Y(_00929_),
    .B1(_05948_));
 sg13g2_nor2_1 _15234_ (.A(net2651),
    .B(net4131),
    .Y(_05949_));
 sg13g2_a21oi_1 _15235_ (.A1(net4982),
    .A2(net4131),
    .Y(_00930_),
    .B1(_05949_));
 sg13g2_nand2_1 _15236_ (.Y(_05950_),
    .A(net4320),
    .B(_05668_));
 sg13g2_nand2_1 _15237_ (.Y(_05951_),
    .A(net1881),
    .B(net4130));
 sg13g2_o21ai_1 _15238_ (.B1(_05951_),
    .Y(_00931_),
    .A1(net4854),
    .A2(net4130));
 sg13g2_nand2_1 _15239_ (.Y(_05952_),
    .A(net1712),
    .B(net4129));
 sg13g2_o21ai_1 _15240_ (.B1(_05952_),
    .Y(_00932_),
    .A1(net4847),
    .A2(net4129));
 sg13g2_nand2_1 _15241_ (.Y(_05953_),
    .A(net2003),
    .B(net4130));
 sg13g2_o21ai_1 _15242_ (.B1(_05953_),
    .Y(_00933_),
    .A1(net4843),
    .A2(net4130));
 sg13g2_nand2_1 _15243_ (.Y(_05954_),
    .A(net1849),
    .B(net4130));
 sg13g2_o21ai_1 _15244_ (.B1(_05954_),
    .Y(_00934_),
    .A1(net4837),
    .A2(_05950_));
 sg13g2_nand2_1 _15245_ (.Y(_05955_),
    .A(net1781),
    .B(net4129));
 sg13g2_o21ai_1 _15246_ (.B1(_05955_),
    .Y(_00935_),
    .A1(net4831),
    .A2(net4129));
 sg13g2_nand2_1 _15247_ (.Y(_05956_),
    .A(net1688),
    .B(net4129));
 sg13g2_o21ai_1 _15248_ (.B1(_05956_),
    .Y(_00936_),
    .A1(net4825),
    .A2(net4130));
 sg13g2_nand2_1 _15249_ (.Y(_05957_),
    .A(net2043),
    .B(net4130));
 sg13g2_o21ai_1 _15250_ (.B1(_05957_),
    .Y(_00937_),
    .A1(net4821),
    .A2(net4129));
 sg13g2_nand2_1 _15251_ (.Y(_05958_),
    .A(net1759),
    .B(net4129));
 sg13g2_o21ai_1 _15252_ (.B1(_05958_),
    .Y(_00938_),
    .A1(net4816),
    .A2(net4129));
 sg13g2_nand2_1 _15253_ (.Y(_05959_),
    .A(net4326),
    .B(_05668_));
 sg13g2_nand2_1 _15254_ (.Y(_05960_),
    .A(net2085),
    .B(net4127));
 sg13g2_o21ai_1 _15255_ (.B1(_05960_),
    .Y(_00939_),
    .A1(net5042),
    .A2(net4127));
 sg13g2_nand2_1 _15256_ (.Y(_05961_),
    .A(net2017),
    .B(net4128));
 sg13g2_o21ai_1 _15257_ (.B1(_05961_),
    .Y(_00940_),
    .A1(net4877),
    .A2(_05959_));
 sg13g2_nand2_1 _15258_ (.Y(_05962_),
    .A(net2030),
    .B(net4128));
 sg13g2_o21ai_1 _15259_ (.B1(_05962_),
    .Y(_00941_),
    .A1(net5035),
    .A2(net4128));
 sg13g2_nand2_1 _15260_ (.Y(_05963_),
    .A(net2179),
    .B(net4128));
 sg13g2_o21ai_1 _15261_ (.B1(_05963_),
    .Y(_00942_),
    .A1(net4869),
    .A2(net4128));
 sg13g2_nand2_1 _15262_ (.Y(_05964_),
    .A(net1884),
    .B(net4127));
 sg13g2_o21ai_1 _15263_ (.B1(_05964_),
    .Y(_00943_),
    .A1(net5031),
    .A2(net4127));
 sg13g2_nand2_1 _15264_ (.Y(_05965_),
    .A(net2034),
    .B(net4128));
 sg13g2_o21ai_1 _15265_ (.B1(_05965_),
    .Y(_00944_),
    .A1(net4864),
    .A2(net4128));
 sg13g2_nand2_1 _15266_ (.Y(_05966_),
    .A(net1846),
    .B(net4127));
 sg13g2_o21ai_1 _15267_ (.B1(_05966_),
    .Y(_00945_),
    .A1(net5029),
    .A2(net4127));
 sg13g2_nand2_1 _15268_ (.Y(_05967_),
    .A(net1869),
    .B(net4127));
 sg13g2_o21ai_1 _15269_ (.B1(_05967_),
    .Y(_00946_),
    .A1(net4863),
    .A2(net4127));
 sg13g2_nor2_2 _15270_ (.A(net4643),
    .B(net4456),
    .Y(_05968_));
 sg13g2_nor2b_1 _15271_ (.A(net4332),
    .B_N(_05968_),
    .Y(_05969_));
 sg13g2_nor2_1 _15272_ (.A(net2681),
    .B(net4126),
    .Y(_05970_));
 sg13g2_a21oi_1 _15273_ (.A1(net5137),
    .A2(net4126),
    .Y(_00947_),
    .B1(_05970_));
 sg13g2_nor2_1 _15274_ (.A(net2479),
    .B(net4125),
    .Y(_05971_));
 sg13g2_a21oi_1 _15275_ (.A1(net4995),
    .A2(_05969_),
    .Y(_00948_),
    .B1(_05971_));
 sg13g2_nor2_1 _15276_ (.A(net2255),
    .B(net4126),
    .Y(_05972_));
 sg13g2_a21oi_1 _15277_ (.A1(net5131),
    .A2(net4126),
    .Y(_00949_),
    .B1(_05972_));
 sg13g2_nor2_1 _15278_ (.A(net2632),
    .B(net4125),
    .Y(_05973_));
 sg13g2_a21oi_1 _15279_ (.A1(net4989),
    .A2(net4125),
    .Y(_00950_),
    .B1(_05973_));
 sg13g2_nor2_1 _15280_ (.A(net2608),
    .B(net4125),
    .Y(_05974_));
 sg13g2_a21oi_1 _15281_ (.A1(net5127),
    .A2(net4125),
    .Y(_00951_),
    .B1(_05974_));
 sg13g2_nor2_1 _15282_ (.A(net2314),
    .B(net4125),
    .Y(_05975_));
 sg13g2_a21oi_1 _15283_ (.A1(net4986),
    .A2(net4126),
    .Y(_00952_),
    .B1(_05975_));
 sg13g2_nor2_1 _15284_ (.A(net2764),
    .B(net4125),
    .Y(_05976_));
 sg13g2_a21oi_1 _15285_ (.A1(net5122),
    .A2(net4125),
    .Y(_00953_),
    .B1(_05976_));
 sg13g2_nor2_1 _15286_ (.A(net2250),
    .B(net4126),
    .Y(_05977_));
 sg13g2_a21oi_1 _15287_ (.A1(net4979),
    .A2(net4126),
    .Y(_00954_),
    .B1(_05977_));
 sg13g2_nand2_1 _15288_ (.Y(_05978_),
    .A(net4324),
    .B(_05968_));
 sg13g2_nand2_1 _15289_ (.Y(_05979_),
    .A(net1716),
    .B(net4124));
 sg13g2_o21ai_1 _15290_ (.B1(_05979_),
    .Y(_00955_),
    .A1(net4856),
    .A2(net4124));
 sg13g2_nand2_1 _15291_ (.Y(_05980_),
    .A(net1802),
    .B(net4124));
 sg13g2_o21ai_1 _15292_ (.B1(_05980_),
    .Y(_00956_),
    .A1(net4850),
    .A2(net4124));
 sg13g2_nand2_1 _15293_ (.Y(_05981_),
    .A(net1894),
    .B(net4124));
 sg13g2_o21ai_1 _15294_ (.B1(_05981_),
    .Y(_00957_),
    .A1(net4845),
    .A2(net4124));
 sg13g2_nand2_1 _15295_ (.Y(_05982_),
    .A(net2239),
    .B(net4124));
 sg13g2_o21ai_1 _15296_ (.B1(_05982_),
    .Y(_00958_),
    .A1(net4839),
    .A2(net4124));
 sg13g2_nand2_1 _15297_ (.Y(_05983_),
    .A(net1739),
    .B(net4123));
 sg13g2_o21ai_1 _15298_ (.B1(_05983_),
    .Y(_00959_),
    .A1(net4834),
    .A2(net4123));
 sg13g2_nand2_1 _15299_ (.Y(_05984_),
    .A(net2190),
    .B(net4123));
 sg13g2_o21ai_1 _15300_ (.B1(_05984_),
    .Y(_00960_),
    .A1(net4828),
    .A2(net4123));
 sg13g2_nand2_1 _15301_ (.Y(_05985_),
    .A(net1828),
    .B(net4123));
 sg13g2_o21ai_1 _15302_ (.B1(_05985_),
    .Y(_00961_),
    .A1(net4822),
    .A2(net4123));
 sg13g2_nand2_1 _15303_ (.Y(_05986_),
    .A(net1691),
    .B(net4123));
 sg13g2_o21ai_1 _15304_ (.B1(_05986_),
    .Y(_00962_),
    .A1(net4817),
    .A2(net4123));
 sg13g2_nand2_1 _15305_ (.Y(_05987_),
    .A(net4328),
    .B(_05968_));
 sg13g2_nand2_1 _15306_ (.Y(_05988_),
    .A(net1684),
    .B(net4122));
 sg13g2_o21ai_1 _15307_ (.B1(_05988_),
    .Y(_00963_),
    .A1(net5043),
    .A2(net4122));
 sg13g2_nand2_1 _15308_ (.Y(_05989_),
    .A(net1680),
    .B(net4121));
 sg13g2_o21ai_1 _15309_ (.B1(_05989_),
    .Y(_00964_),
    .A1(net4875),
    .A2(net4121));
 sg13g2_nand2_1 _15310_ (.Y(_05990_),
    .A(net2252),
    .B(net4122));
 sg13g2_o21ai_1 _15311_ (.B1(_05990_),
    .Y(_00965_),
    .A1(net5038),
    .A2(net4122));
 sg13g2_nand2_1 _15312_ (.Y(_05991_),
    .A(net1785),
    .B(net4122));
 sg13g2_o21ai_1 _15313_ (.B1(_05991_),
    .Y(_00966_),
    .A1(net4871),
    .A2(net4122));
 sg13g2_nand2_1 _15314_ (.Y(_05992_),
    .A(net1666),
    .B(net4121));
 sg13g2_o21ai_1 _15315_ (.B1(_05992_),
    .Y(_00967_),
    .A1(net5032),
    .A2(net4121));
 sg13g2_nand2_1 _15316_ (.Y(_05993_),
    .A(net1960),
    .B(net4122));
 sg13g2_o21ai_1 _15317_ (.B1(_05993_),
    .Y(_00968_),
    .A1(net4866),
    .A2(net4122));
 sg13g2_nand2_1 _15318_ (.Y(_05994_),
    .A(net1833),
    .B(net4121));
 sg13g2_o21ai_1 _15319_ (.B1(_05994_),
    .Y(_00969_),
    .A1(net5026),
    .A2(net4121));
 sg13g2_nand2_1 _15320_ (.Y(_05995_),
    .A(net1855),
    .B(net4121));
 sg13g2_o21ai_1 _15321_ (.B1(_05995_),
    .Y(_00970_),
    .A1(net4860),
    .A2(net4121));
 sg13g2_nand2_1 _15322_ (.Y(_05996_),
    .A(net4324),
    .B(_05640_));
 sg13g2_nand2_1 _15323_ (.Y(_05997_),
    .A(net1816),
    .B(net4120));
 sg13g2_o21ai_1 _15324_ (.B1(_05997_),
    .Y(_00971_),
    .A1(net4856),
    .A2(net4120));
 sg13g2_nand2_1 _15325_ (.Y(_05998_),
    .A(net1807),
    .B(net4120));
 sg13g2_o21ai_1 _15326_ (.B1(_05998_),
    .Y(_00972_),
    .A1(net4850),
    .A2(net4120));
 sg13g2_nand2_1 _15327_ (.Y(_05999_),
    .A(net1995),
    .B(net4120));
 sg13g2_o21ai_1 _15328_ (.B1(_05999_),
    .Y(_00973_),
    .A1(net4845),
    .A2(net4120));
 sg13g2_nand2_1 _15329_ (.Y(_06000_),
    .A(net2139),
    .B(net4120));
 sg13g2_o21ai_1 _15330_ (.B1(_06000_),
    .Y(_00974_),
    .A1(net4839),
    .A2(net4120));
 sg13g2_nand2_1 _15331_ (.Y(_06001_),
    .A(net2213),
    .B(net4119));
 sg13g2_o21ai_1 _15332_ (.B1(_06001_),
    .Y(_00975_),
    .A1(net4834),
    .A2(net4119));
 sg13g2_nand2_1 _15333_ (.Y(_06002_),
    .A(net2038),
    .B(net4119));
 sg13g2_o21ai_1 _15334_ (.B1(_06002_),
    .Y(_00976_),
    .A1(net4828),
    .A2(net4119));
 sg13g2_nand2_1 _15335_ (.Y(_06003_),
    .A(net1725),
    .B(net4119));
 sg13g2_o21ai_1 _15336_ (.B1(_06003_),
    .Y(_00977_),
    .A1(net4822),
    .A2(net4119));
 sg13g2_nand2_1 _15337_ (.Y(_06004_),
    .A(net1942),
    .B(net4119));
 sg13g2_o21ai_1 _15338_ (.B1(_06004_),
    .Y(_00978_),
    .A1(net4817),
    .A2(net4119));
 sg13g2_nand2_2 _15339_ (.Y(_06005_),
    .A(net4328),
    .B(_05640_));
 sg13g2_nand2_1 _15340_ (.Y(_06006_),
    .A(net2048),
    .B(net4118));
 sg13g2_o21ai_1 _15341_ (.B1(_06006_),
    .Y(_00979_),
    .A1(net5043),
    .A2(net4118));
 sg13g2_nand2_1 _15342_ (.Y(_06007_),
    .A(net1845),
    .B(net4117));
 sg13g2_o21ai_1 _15343_ (.B1(_06007_),
    .Y(_00980_),
    .A1(net4874),
    .A2(net4117));
 sg13g2_nand2_1 _15344_ (.Y(_06008_),
    .A(net1686),
    .B(net4118));
 sg13g2_o21ai_1 _15345_ (.B1(_06008_),
    .Y(_00981_),
    .A1(net5038),
    .A2(net4118));
 sg13g2_nand2_1 _15346_ (.Y(_06009_),
    .A(net1758),
    .B(net4118));
 sg13g2_o21ai_1 _15347_ (.B1(_06009_),
    .Y(_00982_),
    .A1(net4871),
    .A2(net4118));
 sg13g2_nand2_1 _15348_ (.Y(_06010_),
    .A(net1718),
    .B(net4117));
 sg13g2_o21ai_1 _15349_ (.B1(_06010_),
    .Y(_00983_),
    .A1(net5032),
    .A2(net4117));
 sg13g2_nand2_1 _15350_ (.Y(_06011_),
    .A(net1958),
    .B(net4118));
 sg13g2_o21ai_1 _15351_ (.B1(_06011_),
    .Y(_00984_),
    .A1(net4866),
    .A2(net4118));
 sg13g2_nand2_1 _15352_ (.Y(_06012_),
    .A(net1770),
    .B(net4117));
 sg13g2_o21ai_1 _15353_ (.B1(_06012_),
    .Y(_00985_),
    .A1(net5026),
    .A2(net4117));
 sg13g2_nand2_1 _15354_ (.Y(_06013_),
    .A(net1848),
    .B(net4117));
 sg13g2_o21ai_1 _15355_ (.B1(_06013_),
    .Y(_00986_),
    .A1(net4859),
    .A2(net4117));
 sg13g2_nor2b_1 _15356_ (.A(net5146),
    .B_N(net2556),
    .Y(_06014_));
 sg13g2_a21o_2 _15357_ (.A2(net5310),
    .A1(net5233),
    .B1(_05130_),
    .X(_06015_));
 sg13g2_a21oi_1 _15358_ (.A1(net5146),
    .A2(_06015_),
    .Y(_06016_),
    .B1(_06014_));
 sg13g2_nor2_1 _15359_ (.A(net2567),
    .B(net4455),
    .Y(_06017_));
 sg13g2_a21oi_1 _15360_ (.A1(net4455),
    .A2(_06016_),
    .Y(_00987_),
    .B1(_06017_));
 sg13g2_nor2b_1 _15361_ (.A(net5146),
    .B_N(\m_sys.m_uart.m_tx.r_data[2] ),
    .Y(_06018_));
 sg13g2_a21o_2 _15362_ (.A2(\m_sys._m_core_io_b_mem_wdata[1] ),
    .A1(net5238),
    .B1(_05134_),
    .X(_06019_));
 sg13g2_a21oi_1 _15363_ (.A1(net5146),
    .A2(_06019_),
    .Y(_06020_),
    .B1(_06018_));
 sg13g2_nor2_1 _15364_ (.A(net2556),
    .B(net4455),
    .Y(_06021_));
 sg13g2_a21oi_1 _15365_ (.A1(net4455),
    .A2(_06020_),
    .Y(_00988_),
    .B1(_06021_));
 sg13g2_nor2b_1 _15366_ (.A(net5146),
    .B_N(net2737),
    .Y(_06022_));
 sg13g2_a21o_2 _15367_ (.A2(\m_sys._m_core_io_b_mem_wdata[2] ),
    .A1(net5236),
    .B1(_05137_),
    .X(_06023_));
 sg13g2_a21oi_1 _15368_ (.A1(net5146),
    .A2(_06023_),
    .Y(_06024_),
    .B1(_06022_));
 sg13g2_nor2_1 _15369_ (.A(net2916),
    .B(net4455),
    .Y(_06025_));
 sg13g2_a21oi_1 _15370_ (.A1(net4455),
    .A2(_06024_),
    .Y(_00989_),
    .B1(_06025_));
 sg13g2_nor2b_1 _15371_ (.A(net5145),
    .B_N(net2702),
    .Y(_06026_));
 sg13g2_a21o_2 _15372_ (.A2(\m_sys._m_core_io_b_mem_wdata[3] ),
    .A1(net5238),
    .B1(_05140_),
    .X(_06027_));
 sg13g2_a21oi_1 _15373_ (.A1(net5146),
    .A2(_06027_),
    .Y(_06028_),
    .B1(_06026_));
 sg13g2_nor2_1 _15374_ (.A(net2737),
    .B(net4455),
    .Y(_06029_));
 sg13g2_a21oi_1 _15375_ (.A1(net4455),
    .A2(_06028_),
    .Y(_00990_),
    .B1(_06029_));
 sg13g2_nor2b_1 _15376_ (.A(net5145),
    .B_N(\m_sys.m_uart.m_tx.r_data[5] ),
    .Y(_06030_));
 sg13g2_a21o_2 _15377_ (.A2(\m_sys._m_core_io_b_mem_wdata[4] ),
    .A1(net5233),
    .B1(_05143_),
    .X(_06031_));
 sg13g2_a21oi_1 _15378_ (.A1(net5145),
    .A2(_06031_),
    .Y(_06032_),
    .B1(_06030_));
 sg13g2_nor2_1 _15379_ (.A(net2702),
    .B(net4454),
    .Y(_06033_));
 sg13g2_a21oi_1 _15380_ (.A1(net4454),
    .A2(_06032_),
    .Y(_00991_),
    .B1(_06033_));
 sg13g2_nor2b_1 _15381_ (.A(net5145),
    .B_N(net2284),
    .Y(_06034_));
 sg13g2_a21o_2 _15382_ (.A2(\m_sys._m_core_io_b_mem_wdata[5] ),
    .A1(net5237),
    .B1(_05146_),
    .X(_06035_));
 sg13g2_a21oi_1 _15383_ (.A1(net5145),
    .A2(_06035_),
    .Y(_06036_),
    .B1(_06034_));
 sg13g2_nor2_1 _15384_ (.A(net2715),
    .B(net4454),
    .Y(_06037_));
 sg13g2_a21oi_1 _15385_ (.A1(net4454),
    .A2(_06036_),
    .Y(_00992_),
    .B1(_06037_));
 sg13g2_nor2b_1 _15386_ (.A(net5145),
    .B_N(\m_sys.m_uart.m_tx.r_data[7] ),
    .Y(_06038_));
 sg13g2_a21o_2 _15387_ (.A2(\m_sys._m_core_io_b_mem_wdata[6] ),
    .A1(net5233),
    .B1(_05149_),
    .X(_06039_));
 sg13g2_a21oi_1 _15388_ (.A1(net5145),
    .A2(_06039_),
    .Y(_06040_),
    .B1(_06038_));
 sg13g2_nor2_1 _15389_ (.A(net2284),
    .B(net4454),
    .Y(_06041_));
 sg13g2_a21oi_1 _15390_ (.A1(net4454),
    .A2(_06040_),
    .Y(_00993_),
    .B1(_06041_));
 sg13g2_nor2b_1 _15391_ (.A(net4318),
    .B_N(_05551_),
    .Y(_06042_));
 sg13g2_nor2_1 _15392_ (.A(net2464),
    .B(net4114),
    .Y(_06043_));
 sg13g2_a21oi_1 _15393_ (.A1(net5023),
    .A2(net4114),
    .Y(_00994_),
    .B1(_06043_));
 sg13g2_nor2_1 _15394_ (.A(net2483),
    .B(net4116),
    .Y(_06044_));
 sg13g2_a21oi_1 _15395_ (.A1(net4814),
    .A2(net4116),
    .Y(_00995_),
    .B1(_06044_));
 sg13g2_nor2_1 _15396_ (.A(net2432),
    .B(net4114),
    .Y(_06045_));
 sg13g2_a21oi_1 _15397_ (.A1(net5018),
    .A2(net4114),
    .Y(_00996_),
    .B1(_06045_));
 sg13g2_nor2_1 _15398_ (.A(net2818),
    .B(net4114),
    .Y(_06046_));
 sg13g2_a21oi_1 _15399_ (.A1(net4809),
    .A2(net4114),
    .Y(_00997_),
    .B1(_06046_));
 sg13g2_nor2_1 _15400_ (.A(net2755),
    .B(net4116),
    .Y(_06047_));
 sg13g2_a21oi_1 _15401_ (.A1(net5014),
    .A2(net4116),
    .Y(_00998_),
    .B1(_06047_));
 sg13g2_nor2_1 _15402_ (.A(net2264),
    .B(net4114),
    .Y(_06048_));
 sg13g2_a21oi_1 _15403_ (.A1(net4803),
    .A2(net4115),
    .Y(_00999_),
    .B1(_06048_));
 sg13g2_nor2_1 _15404_ (.A(net2389),
    .B(net4115),
    .Y(_06049_));
 sg13g2_a21oi_1 _15405_ (.A1(net5007),
    .A2(net4114),
    .Y(_01000_),
    .B1(_06049_));
 sg13g2_nor2_1 _15406_ (.A(net2504),
    .B(net4115),
    .Y(_06050_));
 sg13g2_a21oi_1 _15407_ (.A1(net4799),
    .A2(net4115),
    .Y(_01001_),
    .B1(_06050_));
 sg13g2_nor2b_1 _15408_ (.A(net4334),
    .B_N(_05420_),
    .Y(_06051_));
 sg13g2_nor2_1 _15409_ (.A(net2517),
    .B(net4113),
    .Y(_06052_));
 sg13g2_a21oi_1 _15410_ (.A1(net5139),
    .A2(net4113),
    .Y(_01002_),
    .B1(_06052_));
 sg13g2_nor2_1 _15411_ (.A(net2717),
    .B(net4113),
    .Y(_06053_));
 sg13g2_a21oi_1 _15412_ (.A1(net4996),
    .A2(net4113),
    .Y(_01003_),
    .B1(_06053_));
 sg13g2_nor2_1 _15413_ (.A(net2623),
    .B(net4112),
    .Y(_06054_));
 sg13g2_a21oi_1 _15414_ (.A1(net5134),
    .A2(net4112),
    .Y(_01004_),
    .B1(_06054_));
 sg13g2_nor2_1 _15415_ (.A(net2351),
    .B(net4112),
    .Y(_06055_));
 sg13g2_a21oi_1 _15416_ (.A1(net4992),
    .A2(net4112),
    .Y(_01005_),
    .B1(_06055_));
 sg13g2_nor2_1 _15417_ (.A(net2370),
    .B(_06051_),
    .Y(_06056_));
 sg13g2_a21oi_1 _15418_ (.A1(net5129),
    .A2(net4113),
    .Y(_01006_),
    .B1(_06056_));
 sg13g2_nor2_1 _15419_ (.A(net2488),
    .B(net4113),
    .Y(_06057_));
 sg13g2_a21oi_1 _15420_ (.A1(net4985),
    .A2(net4113),
    .Y(_01007_),
    .B1(_06057_));
 sg13g2_nor2_1 _15421_ (.A(net2617),
    .B(net4112),
    .Y(_06058_));
 sg13g2_a21oi_1 _15422_ (.A1(net5123),
    .A2(net4112),
    .Y(_01008_),
    .B1(_06058_));
 sg13g2_nor2_1 _15423_ (.A(net2327),
    .B(net4112),
    .Y(_06059_));
 sg13g2_a21oi_1 _15424_ (.A1(net4982),
    .A2(net4112),
    .Y(_01009_),
    .B1(_06059_));
 sg13g2_nor2b_1 _15425_ (.A(net4315),
    .B_N(_05968_),
    .Y(_06060_));
 sg13g2_nor2_1 _15426_ (.A(net2260),
    .B(net4110),
    .Y(_06061_));
 sg13g2_a21oi_1 _15427_ (.A1(net5020),
    .A2(net4110),
    .Y(_01010_),
    .B1(_06061_));
 sg13g2_nor2_1 _15428_ (.A(net2698),
    .B(_06060_),
    .Y(_06062_));
 sg13g2_a21oi_1 _15429_ (.A1(net4812),
    .A2(net4111),
    .Y(_01011_),
    .B1(_06062_));
 sg13g2_nor2_1 _15430_ (.A(net2718),
    .B(net4110),
    .Y(_06063_));
 sg13g2_a21oi_1 _15431_ (.A1(net5016),
    .A2(net4110),
    .Y(_01012_),
    .B1(_06063_));
 sg13g2_nor2_1 _15432_ (.A(net2191),
    .B(net4110),
    .Y(_06064_));
 sg13g2_a21oi_1 _15433_ (.A1(net4806),
    .A2(net4110),
    .Y(_01013_),
    .B1(_06064_));
 sg13g2_nor2_1 _15434_ (.A(net2254),
    .B(net4111),
    .Y(_06065_));
 sg13g2_a21oi_1 _15435_ (.A1(net5012),
    .A2(net4111),
    .Y(_01014_),
    .B1(_06065_));
 sg13g2_nor2_1 _15436_ (.A(net2595),
    .B(net4111),
    .Y(_06066_));
 sg13g2_a21oi_1 _15437_ (.A1(net4802),
    .A2(net4111),
    .Y(_01015_),
    .B1(_06066_));
 sg13g2_nor2_1 _15438_ (.A(net2419),
    .B(net4111),
    .Y(_06067_));
 sg13g2_a21oi_1 _15439_ (.A1(net5006),
    .A2(net4110),
    .Y(_01016_),
    .B1(_06067_));
 sg13g2_nor2_1 _15440_ (.A(net2656),
    .B(net4111),
    .Y(_06068_));
 sg13g2_a21oi_1 _15441_ (.A1(net4795),
    .A2(net4110),
    .Y(_01017_),
    .B1(_06068_));
 sg13g2_nand2_1 _15442_ (.Y(_06069_),
    .A(net4330),
    .B(_05551_));
 sg13g2_nand2_1 _15443_ (.Y(_06070_),
    .A(net2080),
    .B(net4108));
 sg13g2_o21ai_1 _15444_ (.B1(_06070_),
    .Y(_01018_),
    .A1(net5045),
    .A2(net4108));
 sg13g2_nand2_1 _15445_ (.Y(_06071_),
    .A(net1955),
    .B(net4108));
 sg13g2_o21ai_1 _15446_ (.B1(_06071_),
    .Y(_01019_),
    .A1(net4874),
    .A2(net4108));
 sg13g2_nand2_1 _15447_ (.Y(_06072_),
    .A(net1751),
    .B(net4107));
 sg13g2_o21ai_1 _15448_ (.B1(_06072_),
    .Y(_01020_),
    .A1(net5040),
    .A2(net4107));
 sg13g2_nand2_1 _15449_ (.Y(_06073_),
    .A(net1932),
    .B(net4109));
 sg13g2_o21ai_1 _15450_ (.B1(_06073_),
    .Y(_01021_),
    .A1(net4870),
    .A2(net4109));
 sg13g2_nand2_1 _15451_ (.Y(_06074_),
    .A(net2110),
    .B(net4109));
 sg13g2_o21ai_1 _15452_ (.B1(_06074_),
    .Y(_01022_),
    .A1(net5030),
    .A2(net4109));
 sg13g2_nand2_1 _15453_ (.Y(_06075_),
    .A(net1803),
    .B(net4107));
 sg13g2_o21ai_1 _15454_ (.B1(_06075_),
    .Y(_01023_),
    .A1(net4868),
    .A2(net4107));
 sg13g2_nand2_1 _15455_ (.Y(_06076_),
    .A(net1827),
    .B(net4107));
 sg13g2_o21ai_1 _15456_ (.B1(_06076_),
    .Y(_01024_),
    .A1(net5027),
    .A2(net4107));
 sg13g2_nand2_1 _15457_ (.Y(_06077_),
    .A(net1813),
    .B(net4107));
 sg13g2_o21ai_1 _15458_ (.B1(_06077_),
    .Y(_01025_),
    .A1(net4859),
    .A2(net4107));
 sg13g2_nand3_1 _15459_ (.B(net5283),
    .C(_02709_),
    .A(net5282),
    .Y(_06078_));
 sg13g2_nand2_2 _15460_ (.Y(_06079_),
    .A(_02360_),
    .B(net5283));
 sg13g2_nor2_1 _15461_ (.A(_02706_),
    .B(_06079_),
    .Y(_06080_));
 sg13g2_or2_2 _15462_ (.X(_06081_),
    .B(_06079_),
    .A(_02706_));
 sg13g2_and2_2 _15463_ (.A(net5004),
    .B(_06081_),
    .X(_06082_));
 sg13g2_nand2_2 _15464_ (.Y(_06083_),
    .A(net5004),
    .B(_06081_));
 sg13g2_or2_1 _15465_ (.X(_06084_),
    .B(_04922_),
    .A(_02600_));
 sg13g2_inv_1 _15466_ (.Y(_06085_),
    .A(_06084_));
 sg13g2_nor4_1 _15467_ (.A(\m_sys.m_bootloader.r_byte_cnt[4] ),
    .B(\m_sys.m_bootloader.r_byte_cnt[5] ),
    .C(\m_sys.m_bootloader.r_byte_cnt[6] ),
    .D(\m_sys.m_bootloader.r_byte_cnt[7] ),
    .Y(_06086_));
 sg13g2_nor4_1 _15468_ (.A(_02401_),
    .B(\m_sys.m_bootloader.r_byte_cnt[1] ),
    .C(\m_sys.m_bootloader.r_byte_cnt[2] ),
    .D(\m_sys.m_bootloader.r_byte_cnt[3] ),
    .Y(_06087_));
 sg13g2_nand2_1 _15469_ (.Y(_06088_),
    .A(_06086_),
    .B(_06087_));
 sg13g2_or4_1 _15470_ (.A(\m_sys.m_bootloader.r_byte_cnt[8] ),
    .B(\m_sys.m_bootloader.r_byte_cnt[9] ),
    .C(\m_sys.m_bootloader.r_byte_cnt[10] ),
    .D(\m_sys.m_bootloader.r_byte_cnt[11] ),
    .X(_06089_));
 sg13g2_or4_1 _15471_ (.A(\m_sys.m_bootloader.r_byte_cnt[12] ),
    .B(\m_sys.m_bootloader.r_byte_cnt[13] ),
    .C(\m_sys.m_bootloader.r_byte_cnt[14] ),
    .D(\m_sys.m_bootloader.r_byte_cnt[15] ),
    .X(_06090_));
 sg13g2_nor3_1 _15472_ (.A(_06088_),
    .B(_06089_),
    .C(_06090_),
    .Y(_06091_));
 sg13g2_nor2_1 _15473_ (.A(_02401_),
    .B(\m_sys.m_bootloader.r_byte_cnt[3] ),
    .Y(_06092_));
 sg13g2_nor3_1 _15474_ (.A(\m_sys.m_bootloader.r_byte_cnt[8] ),
    .B(\m_sys.m_bootloader.r_byte_cnt[11] ),
    .C(_06090_),
    .Y(_06093_));
 sg13g2_nor4_1 _15475_ (.A(\m_sys.m_bootloader.r_byte_cnt[1] ),
    .B(\m_sys.m_bootloader.r_byte_cnt[2] ),
    .C(\m_sys.m_bootloader.r_byte_cnt[9] ),
    .D(\m_sys.m_bootloader.r_byte_cnt[10] ),
    .Y(_06094_));
 sg13g2_and4_1 _15476_ (.A(_06086_),
    .B(_06092_),
    .C(_06093_),
    .D(_06094_),
    .X(_06095_));
 sg13g2_nor2b_2 _15477_ (.A(net4715),
    .B_N(_06095_),
    .Y(_06096_));
 sg13g2_nand2_2 _15478_ (.Y(_06097_),
    .A(_06085_),
    .B(_06095_));
 sg13g2_nand3_1 _15479_ (.B(_02713_),
    .C(_02715_),
    .A(net5268),
    .Y(_06098_));
 sg13g2_nand2_1 _15480_ (.Y(_06099_),
    .A(net5147),
    .B(_04895_));
 sg13g2_nor2_1 _15481_ (.A(_02706_),
    .B(_02712_),
    .Y(_06100_));
 sg13g2_or2_1 _15482_ (.X(_06101_),
    .B(_02712_),
    .A(_02706_));
 sg13g2_nand4_1 _15483_ (.B(net5283),
    .C(\m_sys.m_bootloader.r_cstate[1] ),
    .A(net5282),
    .Y(_06102_),
    .D(net5286));
 sg13g2_inv_1 _15484_ (.Y(_06103_),
    .A(_06102_));
 sg13g2_nor2_2 _15485_ (.A(\m_sys.m_bootloader.r_cstate[4] ),
    .B(_06102_),
    .Y(_06104_));
 sg13g2_nand2_1 _15486_ (.Y(_06105_),
    .A(_02359_),
    .B(_06103_));
 sg13g2_nand2_1 _15487_ (.Y(_06106_),
    .A(_02709_),
    .B(_04893_));
 sg13g2_nor2_2 _15488_ (.A(net5284),
    .B(_06106_),
    .Y(_06107_));
 sg13g2_nor4_1 _15489_ (.A(_06083_),
    .B(_06100_),
    .C(_06104_),
    .D(_06107_),
    .Y(_06108_));
 sg13g2_nor3_2 _15490_ (.A(net5282),
    .B(net5284),
    .C(_02706_),
    .Y(_06109_));
 sg13g2_nor2b_2 _15491_ (.A(net5283),
    .B_N(_06109_),
    .Y(_06110_));
 sg13g2_nand2_1 _15492_ (.Y(_06111_),
    .A(_02707_),
    .B(_04893_));
 sg13g2_nor3_1 _15493_ (.A(net5284),
    .B(_02710_),
    .C(_02712_),
    .Y(_06112_));
 sg13g2_nand3b_1 _15494_ (.B(_02361_),
    .C(_02709_),
    .Y(_06113_),
    .A_N(_02712_));
 sg13g2_nand2_1 _15495_ (.Y(_06114_),
    .A(_06111_),
    .B(_06113_));
 sg13g2_nor2_1 _15496_ (.A(_02711_),
    .B(_04894_),
    .Y(_06115_));
 sg13g2_nand3_1 _15497_ (.B(_02709_),
    .C(_04893_),
    .A(net5284),
    .Y(_06116_));
 sg13g2_nand3_1 _15498_ (.B(_06113_),
    .C(_06116_),
    .A(net4789),
    .Y(_06117_));
 sg13g2_nor2_1 _15499_ (.A(_02711_),
    .B(_06079_),
    .Y(_06118_));
 sg13g2_and2_1 _15500_ (.A(_02360_),
    .B(_04897_),
    .X(_06119_));
 sg13g2_nor2_1 _15501_ (.A(_06118_),
    .B(_06119_),
    .Y(_06120_));
 sg13g2_nor2b_1 _15502_ (.A(_06117_),
    .B_N(_06120_),
    .Y(_06121_));
 sg13g2_nand4_1 _15503_ (.B(_06099_),
    .C(_06108_),
    .A(_06098_),
    .Y(_06122_),
    .D(_06121_));
 sg13g2_nor3_2 _15504_ (.A(net5284),
    .B(_02710_),
    .C(_06079_),
    .Y(_06123_));
 sg13g2_nand2b_1 _15505_ (.Y(_06124_),
    .B(_04897_),
    .A_N(net5147));
 sg13g2_a22oi_1 _15506_ (.Y(_06125_),
    .B1(_06117_),
    .B2(net4715),
    .A2(_06097_),
    .A1(_06083_));
 sg13g2_nand3_1 _15507_ (.B(_06124_),
    .C(_06125_),
    .A(_06122_),
    .Y(_06126_));
 sg13g2_a21oi_1 _15508_ (.A1(net1),
    .A2(_06107_),
    .Y(_06127_),
    .B1(net4347));
 sg13g2_nand2_2 _15509_ (.Y(_06128_),
    .A(net5285),
    .B(net4792));
 sg13g2_nand2_1 _15510_ (.Y(_06129_),
    .A(_02708_),
    .B(net5004));
 sg13g2_xnor2_1 _15511_ (.Y(_06130_),
    .A(\m_sys.m_bootloader.r_num_cnt[3] ),
    .B(\m_sys.m_bootloader.r_num[3] ));
 sg13g2_xnor2_1 _15512_ (.Y(_06131_),
    .A(\m_sys.m_bootloader.r_num_cnt[0] ),
    .B(\m_sys.m_bootloader.r_num[0] ));
 sg13g2_xor2_1 _15513_ (.B(\m_sys.m_bootloader.r_num[6] ),
    .A(\m_sys.m_bootloader.r_num_cnt[6] ),
    .X(_06132_));
 sg13g2_xnor2_1 _15514_ (.Y(_06133_),
    .A(\m_sys.m_bootloader.r_num_cnt[4] ),
    .B(\m_sys.m_bootloader.r_num[4] ));
 sg13g2_xnor2_1 _15515_ (.Y(_06134_),
    .A(\m_sys.m_bootloader.r_num_cnt[7] ),
    .B(\m_sys.m_bootloader.r_num[7] ));
 sg13g2_xnor2_1 _15516_ (.Y(_06135_),
    .A(\m_sys.m_bootloader.r_num_cnt[5] ),
    .B(\m_sys.m_bootloader.r_num[5] ));
 sg13g2_xnor2_1 _15517_ (.Y(_06136_),
    .A(\m_sys.m_bootloader.r_num_cnt[2] ),
    .B(\m_sys.m_bootloader.r_num[2] ));
 sg13g2_xnor2_1 _15518_ (.Y(_06137_),
    .A(\m_sys.m_bootloader.r_num_cnt[1] ),
    .B(\m_sys.m_bootloader.r_num[1] ));
 sg13g2_nand3_1 _15519_ (.B(_06135_),
    .C(_06136_),
    .A(_06134_),
    .Y(_06138_));
 sg13g2_nand4_1 _15520_ (.B(_06131_),
    .C(_06133_),
    .A(_06130_),
    .Y(_06139_),
    .D(_06137_));
 sg13g2_nor3_2 _15521_ (.A(_06132_),
    .B(_06138_),
    .C(_06139_),
    .Y(_06140_));
 sg13g2_nor3_1 _15522_ (.A(\m_sys.m_bootloader.r_offset_0[0] ),
    .B(\m_sys.m_bootloader.r_offset_0[1] ),
    .C(\m_sys.m_bootloader.r_offset_0[2] ),
    .Y(_06141_));
 sg13g2_or4_2 _15523_ (.A(\m_sys.m_bootloader.r_offset_0[0] ),
    .B(\m_sys.m_bootloader.r_offset_0[1] ),
    .C(\m_sys.m_bootloader.r_offset_0[2] ),
    .D(\m_sys.m_bootloader.r_offset_0[3] ),
    .X(_06142_));
 sg13g2_or3_1 _15524_ (.A(\m_sys.m_bootloader.r_offset_0[4] ),
    .B(\m_sys.m_bootloader.r_offset_0[5] ),
    .C(_06142_),
    .X(_06143_));
 sg13g2_or2_1 _15525_ (.X(_06144_),
    .B(\m_sys.m_bootloader.r_offset_0[7] ),
    .A(\m_sys.m_bootloader.r_offset_0[6] ));
 sg13g2_nor4_2 _15526_ (.A(\m_sys.m_bootloader.r_offset_0[4] ),
    .B(\m_sys.m_bootloader.r_offset_0[5] ),
    .C(_06142_),
    .Y(_06145_),
    .D(_06144_));
 sg13g2_nand2b_1 _15527_ (.Y(_06146_),
    .B(_06145_),
    .A_N(\m_sys.m_bootloader.r_offset_1[0] ));
 sg13g2_or4_2 _15528_ (.A(\m_sys.m_bootloader.r_offset_1[0] ),
    .B(\m_sys.m_bootloader.r_offset_1[1] ),
    .C(_06143_),
    .D(_06144_),
    .X(_06147_));
 sg13g2_nor3_1 _15529_ (.A(\m_sys.m_bootloader.r_offset_1[2] ),
    .B(\m_sys.m_bootloader.r_offset_1[3] ),
    .C(_06147_),
    .Y(_06148_));
 sg13g2_nor4_2 _15530_ (.A(\m_sys.m_bootloader.r_offset_1[2] ),
    .B(\m_sys.m_bootloader.r_offset_1[3] ),
    .C(\m_sys.m_bootloader.r_offset_1[4] ),
    .Y(_06149_),
    .D(_06147_));
 sg13g2_nor2b_1 _15531_ (.A(\m_sys.m_bootloader.r_offset_1[5] ),
    .B_N(_06149_),
    .Y(_06150_));
 sg13g2_nand2b_1 _15532_ (.Y(_06151_),
    .B(_06150_),
    .A_N(\m_sys.m_bootloader.r_offset_1[6] ));
 sg13g2_xnor2_1 _15533_ (.Y(_06152_),
    .A(\m_sys.m_bootloader.r_offset_1[7] ),
    .B(_00042_));
 sg13g2_xnor2_1 _15534_ (.Y(_06153_),
    .A(_06151_),
    .B(_06152_));
 sg13g2_xor2_1 _15535_ (.B(_06149_),
    .A(\m_sys.m_bootloader.r_offset_1[5] ),
    .X(_06154_));
 sg13g2_xnor2_1 _15536_ (.Y(_06155_),
    .A(_00040_),
    .B(_06154_));
 sg13g2_xnor2_1 _15537_ (.Y(_06156_),
    .A(\m_sys.m_bootloader.r_offset_1[6] ),
    .B(_06150_));
 sg13g2_nand2b_1 _15538_ (.Y(_06157_),
    .B(_00041_),
    .A_N(_06156_));
 sg13g2_nand2b_1 _15539_ (.Y(_06158_),
    .B(_06156_),
    .A_N(_00041_));
 sg13g2_o21ai_1 _15540_ (.B1(\m_sys.m_bootloader.r_offset_1[3] ),
    .Y(_06159_),
    .A1(\m_sys.m_bootloader.r_offset_1[2] ),
    .A2(_06147_));
 sg13g2_nand2b_1 _15541_ (.Y(_06160_),
    .B(_06159_),
    .A_N(_06148_));
 sg13g2_xnor2_1 _15542_ (.Y(_06161_),
    .A(_00038_),
    .B(_06160_));
 sg13g2_xor2_1 _15543_ (.B(_06147_),
    .A(\m_sys.m_bootloader.r_offset_1[2] ),
    .X(_06162_));
 sg13g2_nand2b_1 _15544_ (.Y(_06163_),
    .B(_00037_),
    .A_N(_06162_));
 sg13g2_xnor2_1 _15545_ (.Y(_06164_),
    .A(\m_sys.m_bootloader.r_offset_1[0] ),
    .B(_06145_));
 sg13g2_nor2b_1 _15546_ (.A(_06164_),
    .B_N(_00035_),
    .Y(_06165_));
 sg13g2_o21ai_1 _15547_ (.B1(\m_sys.m_bootloader.r_offset_0[2] ),
    .Y(_06166_),
    .A1(\m_sys.m_bootloader.r_offset_0[0] ),
    .A2(\m_sys.m_bootloader.r_offset_0[1] ));
 sg13g2_nor2b_1 _15548_ (.A(_06141_),
    .B_N(_06166_),
    .Y(_06167_));
 sg13g2_xnor2_1 _15549_ (.Y(_06168_),
    .A(\m_sys.m_bootloader.r_offset_0[1] ),
    .B(\m_sys.m_bootloader.r_byte_cnt[1] ));
 sg13g2_nand3_1 _15550_ (.B(\m_sys.m_bootloader.r_offset_0[0] ),
    .C(_06168_),
    .A(_02401_),
    .Y(_06169_));
 sg13g2_nand2b_1 _15551_ (.Y(_06170_),
    .B(\m_sys.m_bootloader.r_byte_cnt[0] ),
    .A_N(\m_sys.m_bootloader.r_offset_0[0] ));
 sg13g2_o21ai_1 _15552_ (.B1(_06169_),
    .Y(_06171_),
    .A1(_06168_),
    .A2(_06170_));
 sg13g2_xnor2_1 _15553_ (.Y(_06172_),
    .A(_00028_),
    .B(_06167_));
 sg13g2_xnor2_1 _15554_ (.Y(_06173_),
    .A(\m_sys.m_bootloader.r_offset_0[3] ),
    .B(_06141_));
 sg13g2_xnor2_1 _15555_ (.Y(_06174_),
    .A(_00029_),
    .B(_06173_));
 sg13g2_xor2_1 _15556_ (.B(_06142_),
    .A(\m_sys.m_bootloader.r_offset_0[4] ),
    .X(_06175_));
 sg13g2_xnor2_1 _15557_ (.Y(_06176_),
    .A(_00030_),
    .B(_06175_));
 sg13g2_nand4_1 _15558_ (.B(_06172_),
    .C(_06174_),
    .A(_06171_),
    .Y(_06177_),
    .D(_06176_));
 sg13g2_o21ai_1 _15559_ (.B1(\m_sys.m_bootloader.r_offset_0[5] ),
    .Y(_06178_),
    .A1(\m_sys.m_bootloader.r_offset_0[4] ),
    .A2(_06142_));
 sg13g2_nand2_1 _15560_ (.Y(_06179_),
    .A(_06143_),
    .B(_06178_));
 sg13g2_xnor2_1 _15561_ (.Y(_06180_),
    .A(_00031_),
    .B(_06179_));
 sg13g2_nor3_1 _15562_ (.A(_06165_),
    .B(_06177_),
    .C(_06180_),
    .Y(_06181_));
 sg13g2_nand2b_1 _15563_ (.Y(_06182_),
    .B(_06164_),
    .A_N(_00035_));
 sg13g2_xnor2_1 _15564_ (.Y(_06183_),
    .A(\m_sys.m_bootloader.r_offset_0[7] ),
    .B(_00034_));
 sg13g2_nand2b_1 _15565_ (.Y(_06184_),
    .B(_00033_),
    .A_N(_00032_));
 sg13g2_o21ai_1 _15566_ (.B1(_06184_),
    .Y(_06185_),
    .A1(_06143_),
    .A2(_06183_));
 sg13g2_a21oi_1 _15567_ (.A1(_02403_),
    .A2(_00032_),
    .Y(_06186_),
    .B1(_06183_));
 sg13g2_nor2_1 _15568_ (.A(_06143_),
    .B(_06186_),
    .Y(_06187_));
 sg13g2_mux2_1 _15569_ (.A0(_06186_),
    .A1(_06187_),
    .S(_06185_),
    .X(_06188_));
 sg13g2_nand4_1 _15570_ (.B(_06181_),
    .C(_06182_),
    .A(_06163_),
    .Y(_06189_),
    .D(_06188_));
 sg13g2_xnor2_1 _15571_ (.Y(_06190_),
    .A(\m_sys.m_bootloader.r_offset_1[1] ),
    .B(_06146_));
 sg13g2_xnor2_1 _15572_ (.Y(_06191_),
    .A(_00036_),
    .B(_06190_));
 sg13g2_nor2b_1 _15573_ (.A(_00037_),
    .B_N(_06162_),
    .Y(_06192_));
 sg13g2_nor4_1 _15574_ (.A(_06161_),
    .B(_06189_),
    .C(_06191_),
    .D(_06192_),
    .Y(_06193_));
 sg13g2_xnor2_1 _15575_ (.Y(_06194_),
    .A(\m_sys.m_bootloader.r_offset_1[4] ),
    .B(_06148_));
 sg13g2_xnor2_1 _15576_ (.Y(_06195_),
    .A(_00039_),
    .B(_06194_));
 sg13g2_nand4_1 _15577_ (.B(_06158_),
    .C(_06193_),
    .A(_06157_),
    .Y(_06196_),
    .D(_06195_));
 sg13g2_nor3_2 _15578_ (.A(_06153_),
    .B(_06155_),
    .C(_06196_),
    .Y(_06197_));
 sg13g2_inv_1 _15579_ (.Y(_06198_),
    .A(_06197_));
 sg13g2_and2_1 _15580_ (.A(_06140_),
    .B(_06197_),
    .X(_06199_));
 sg13g2_nand2_1 _15581_ (.Y(_06200_),
    .A(_06140_),
    .B(_06197_));
 sg13g2_a21oi_1 _15582_ (.A1(_06105_),
    .A2(_06199_),
    .Y(_06201_),
    .B1(_06129_));
 sg13g2_o21ai_1 _15583_ (.B1(_06101_),
    .Y(_06202_),
    .A1(_02360_),
    .A2(_02711_));
 sg13g2_o21ai_1 _15584_ (.B1(_06113_),
    .Y(_06203_),
    .A1(_06201_),
    .A2(_06202_));
 sg13g2_a21o_1 _15585_ (.A2(_06203_),
    .A1(_06128_),
    .B1(_06109_),
    .X(_06204_));
 sg13g2_or4_1 _15586_ (.A(\m_sys._m_uart_io_o_bl_data[7] ),
    .B(net5261),
    .C(\m_sys._m_uart_io_o_bl_data[5] ),
    .D(net5263),
    .X(_06205_));
 sg13g2_nor3_2 _15587_ (.A(\m_sys._m_uart_io_o_bl_data[3] ),
    .B(net5265),
    .C(_06205_),
    .Y(_06206_));
 sg13g2_nand3_1 _15588_ (.B(_06110_),
    .C(_06206_),
    .A(\m_sys._m_uart_io_o_bl_data[0] ),
    .Y(_06207_));
 sg13g2_nand4_1 _15589_ (.B(_06120_),
    .C(_06204_),
    .A(_06106_),
    .Y(_06208_),
    .D(_06207_));
 sg13g2_a221oi_1 _15590_ (.B2(_06208_),
    .C1(net5369),
    .B1(_06127_),
    .A1(_02361_),
    .Y(_01026_),
    .A2(net4347));
 sg13g2_nor3_1 _15591_ (.A(net5285),
    .B(_02706_),
    .C(_02712_),
    .Y(_06209_));
 sg13g2_o21ai_1 _15592_ (.B1(_06100_),
    .Y(_06210_),
    .A1(_02361_),
    .A2(_06140_));
 sg13g2_nor2_1 _15593_ (.A(net5286),
    .B(net5004),
    .Y(_06211_));
 sg13g2_nor2_1 _15594_ (.A(_06104_),
    .B(_06211_),
    .Y(_06212_));
 sg13g2_nand2_1 _15595_ (.Y(_06213_),
    .A(_06210_),
    .B(_06212_));
 sg13g2_nand2_1 _15596_ (.Y(_06214_),
    .A(_06197_),
    .B(_06209_));
 sg13g2_o21ai_1 _15597_ (.B1(_06213_),
    .Y(_06215_),
    .A1(_06140_),
    .A2(_06214_));
 sg13g2_a21oi_1 _15598_ (.A1(_06118_),
    .A2(_06140_),
    .Y(_06216_),
    .B1(_06119_));
 sg13g2_nor3_1 _15599_ (.A(\m_sys._m_uart_io_o_bl_data[1] ),
    .B(\m_sys._m_uart_io_o_bl_data[0] ),
    .C(_06116_),
    .Y(_06217_));
 sg13g2_a21oi_1 _15600_ (.A1(_06206_),
    .A2(_06217_),
    .Y(_06218_),
    .B1(_06107_));
 sg13g2_nand3_1 _15601_ (.B(\m_sys._m_uart_io_o_bl_data[0] ),
    .C(_06110_),
    .A(\m_sys._m_uart_io_o_bl_data[1] ),
    .Y(_06219_));
 sg13g2_o21ai_1 _15602_ (.B1(_06206_),
    .Y(_06220_),
    .A1(\m_sys._m_uart_io_o_bl_data[1] ),
    .A2(\m_sys._m_uart_io_o_bl_data[0] ));
 sg13g2_a221oi_1 _15603_ (.B2(_06220_),
    .C1(_06112_),
    .B1(_06110_),
    .A1(net5284),
    .Y(_06221_),
    .A2(net4792));
 sg13g2_nand4_1 _15604_ (.B(_06218_),
    .C(_06219_),
    .A(_06216_),
    .Y(_06222_),
    .D(_06221_));
 sg13g2_a21o_1 _15605_ (.A2(_06206_),
    .A1(\m_sys._m_uart_io_o_bl_data[1] ),
    .B1(net4789),
    .X(_06223_));
 sg13g2_o21ai_1 _15606_ (.B1(_06223_),
    .Y(_06224_),
    .A1(_02342_),
    .A2(net4789));
 sg13g2_nor2_1 _15607_ (.A(_06126_),
    .B(_06222_),
    .Y(_06225_));
 sg13g2_a22oi_1 _15608_ (.Y(_06226_),
    .B1(_06215_),
    .B2(_06225_),
    .A2(net4347),
    .A1(net3410));
 sg13g2_nor2_1 _15609_ (.A(net5369),
    .B(_06226_),
    .Y(_01027_));
 sg13g2_nor2_2 _15610_ (.A(net5286),
    .B(_06081_),
    .Y(_06227_));
 sg13g2_nor2_1 _15611_ (.A(_06104_),
    .B(_06197_),
    .Y(_06228_));
 sg13g2_o21ai_1 _15612_ (.B1(_04899_),
    .Y(_06229_),
    .A1(_06129_),
    .A2(_06228_));
 sg13g2_nand2_1 _15613_ (.Y(_06230_),
    .A(_06210_),
    .B(_06229_));
 sg13g2_o21ai_1 _15614_ (.B1(_06128_),
    .Y(_06231_),
    .A1(_02710_),
    .A2(_02712_));
 sg13g2_a21oi_1 _15615_ (.A1(_06200_),
    .A2(_06209_),
    .Y(_06232_),
    .B1(_06231_));
 sg13g2_a21oi_1 _15616_ (.A1(_06230_),
    .A2(_06232_),
    .Y(_06233_),
    .B1(_06227_));
 sg13g2_o21ai_1 _15617_ (.B1(_06216_),
    .Y(_06234_),
    .A1(_06118_),
    .A2(_06233_));
 sg13g2_a21oi_1 _15618_ (.A1(net4789),
    .A2(_06234_),
    .Y(_06235_),
    .B1(_06224_));
 sg13g2_o21ai_1 _15619_ (.B1(_06218_),
    .Y(_06236_),
    .A1(_06115_),
    .A2(_06235_));
 sg13g2_a22oi_1 _15620_ (.Y(_06237_),
    .B1(_06127_),
    .B2(_06236_),
    .A2(net4347),
    .A1(net5283));
 sg13g2_nor2_1 _15621_ (.A(net5369),
    .B(_06237_),
    .Y(_01028_));
 sg13g2_nand2b_1 _15622_ (.Y(_06238_),
    .B(_06229_),
    .A_N(_06231_));
 sg13g2_a21oi_1 _15623_ (.A1(_06120_),
    .A2(_06238_),
    .Y(_06239_),
    .B1(_06109_));
 sg13g2_nand2_1 _15624_ (.Y(_06240_),
    .A(_06106_),
    .B(_06223_));
 sg13g2_nor3_1 _15625_ (.A(_06227_),
    .B(_06239_),
    .C(_06240_),
    .Y(_06241_));
 sg13g2_o21ai_1 _15626_ (.B1(net5383),
    .Y(_06242_),
    .A1(net4347),
    .A2(_06241_));
 sg13g2_a21oi_1 _15627_ (.A1(_02360_),
    .A2(net4347),
    .Y(_01029_),
    .B1(_06242_));
 sg13g2_o21ai_1 _15628_ (.B1(net5383),
    .Y(_06243_),
    .A1(_06103_),
    .A2(net4347));
 sg13g2_a21oi_1 _15629_ (.A1(_02359_),
    .A2(net4347),
    .Y(_01030_),
    .B1(_06243_));
 sg13g2_nor2_1 _15630_ (.A(net4714),
    .B(net4789),
    .Y(_06244_));
 sg13g2_mux2_1 _15631_ (.A0(\m_sys.m_bootloader.r_num_cnt[0] ),
    .A1(net3210),
    .S(_06244_),
    .X(_06245_));
 sg13g2_nor2b_1 _15632_ (.A(net4790),
    .B_N(net3211),
    .Y(_01031_));
 sg13g2_a21oi_1 _15633_ (.A1(\m_sys.m_bootloader.r_num_cnt[0] ),
    .A2(_06244_),
    .Y(_06246_),
    .B1(net2877));
 sg13g2_and3_1 _15634_ (.X(_06247_),
    .A(net2877),
    .B(\m_sys.m_bootloader.r_num_cnt[0] ),
    .C(_06244_));
 sg13g2_nor3_1 _15635_ (.A(net4790),
    .B(net2878),
    .C(_06247_),
    .Y(_01032_));
 sg13g2_nor2_1 _15636_ (.A(net3107),
    .B(_06247_),
    .Y(_06248_));
 sg13g2_and2_1 _15637_ (.A(net3107),
    .B(_06247_),
    .X(_06249_));
 sg13g2_nor3_1 _15638_ (.A(net4790),
    .B(net3108),
    .C(_06249_),
    .Y(_01033_));
 sg13g2_nor2_1 _15639_ (.A(net3137),
    .B(_06249_),
    .Y(_06250_));
 sg13g2_and2_1 _15640_ (.A(net3137),
    .B(_06249_),
    .X(_06251_));
 sg13g2_nor3_1 _15641_ (.A(net4790),
    .B(_06250_),
    .C(_06251_),
    .Y(_01034_));
 sg13g2_nor2_1 _15642_ (.A(net3181),
    .B(_06251_),
    .Y(_06252_));
 sg13g2_and2_1 _15643_ (.A(net3181),
    .B(_06251_),
    .X(_06253_));
 sg13g2_nor3_1 _15644_ (.A(net4790),
    .B(_06252_),
    .C(_06253_),
    .Y(_01035_));
 sg13g2_nor2_1 _15645_ (.A(net3123),
    .B(_06253_),
    .Y(_06254_));
 sg13g2_and2_1 _15646_ (.A(net3123),
    .B(_06253_),
    .X(_06255_));
 sg13g2_nor3_1 _15647_ (.A(net4790),
    .B(net3124),
    .C(_06255_),
    .Y(_01036_));
 sg13g2_nor2_1 _15648_ (.A(net3121),
    .B(_06255_),
    .Y(_06256_));
 sg13g2_and2_1 _15649_ (.A(net3121),
    .B(_06255_),
    .X(_06257_));
 sg13g2_nor3_1 _15650_ (.A(net4790),
    .B(net3122),
    .C(_06257_),
    .Y(_01037_));
 sg13g2_a21oi_1 _15651_ (.A1(net3171),
    .A2(_06257_),
    .Y(_06258_),
    .B1(net4790));
 sg13g2_o21ai_1 _15652_ (.B1(_06258_),
    .Y(_06259_),
    .A1(net3171),
    .A2(_06257_));
 sg13g2_inv_1 _15653_ (.Y(_01038_),
    .A(_06259_));
 sg13g2_nand2b_1 _15654_ (.Y(_06260_),
    .B(_06098_),
    .A_N(_02704_));
 sg13g2_and3_1 _15655_ (.X(_01039_),
    .A(net5384),
    .B(net1654),
    .C(_06260_));
 sg13g2_a21oi_1 _15656_ (.A1(net4715),
    .A2(_06114_),
    .Y(_06261_),
    .B1(_06224_));
 sg13g2_o21ai_1 _15657_ (.B1(_06261_),
    .Y(_06262_),
    .A1(_06104_),
    .A2(_06114_));
 sg13g2_nor2_2 _15658_ (.A(_06110_),
    .B(net4382),
    .Y(_06263_));
 sg13g2_nand2b_1 _15659_ (.Y(_06264_),
    .B(net4789),
    .A_N(net4382));
 sg13g2_nor2_1 _15660_ (.A(\m_sys._m_gpio8_io_b_mem_rdata[0] ),
    .B(_03512_),
    .Y(_06265_));
 sg13g2_o21ai_1 _15661_ (.B1(_04869_),
    .Y(_06266_),
    .A1(\m_sys._m_uart_io_b_mem_rdata[0] ),
    .A2(net4880));
 sg13g2_o21ai_1 _15662_ (.B1(net5274),
    .Y(_06267_),
    .A1(_06265_),
    .A2(_06266_));
 sg13g2_nand3_1 _15663_ (.B(_02389_),
    .C(_02715_),
    .A(\m_sys._m_bootloader_io_b_mem_addr[11] ),
    .Y(_06268_));
 sg13g2_nand2b_1 _15664_ (.Y(_06269_),
    .B(net4998),
    .A_N(\m_sys._m_uart_io_b_mem_rdata[0] ));
 sg13g2_o21ai_1 _15665_ (.B1(_06269_),
    .Y(_06270_),
    .A1(\m_sys._m_gpio8_io_b_mem_rdata[0] ),
    .A2(net4998));
 sg13g2_a21oi_1 _15666_ (.A1(\m_sys._m_ram_io_b_port_rdata[0] ),
    .A2(net5140),
    .Y(_06271_),
    .B1(net4878));
 sg13g2_o21ai_1 _15667_ (.B1(_06271_),
    .Y(_06272_),
    .A1(net5140),
    .A2(_06270_));
 sg13g2_a21o_1 _15668_ (.A2(_06272_),
    .A1(_06267_),
    .B1(net5001),
    .X(_06273_));
 sg13g2_o21ai_1 _15669_ (.B1(_06273_),
    .Y(_06274_),
    .A1(\m_sys._m_uart_io_o_bl_data[0] ),
    .A2(_06113_));
 sg13g2_nand2_1 _15670_ (.Y(_06275_),
    .A(net3326),
    .B(net4382));
 sg13g2_o21ai_1 _15671_ (.B1(_06275_),
    .Y(_01040_),
    .A1(_06264_),
    .A2(_06274_));
 sg13g2_mux2_1 _15672_ (.A0(\m_sys._m_gpio8_io_b_mem_rdata[1] ),
    .A1(\m_sys._m_uart_io_b_mem_rdata[1] ),
    .S(net4999),
    .X(_06276_));
 sg13g2_nand2_1 _15673_ (.Y(_06277_),
    .A(_02717_),
    .B(_06276_));
 sg13g2_a21oi_1 _15674_ (.A1(\m_sys._m_ram_io_b_port_rdata[1] ),
    .A2(_02716_),
    .Y(_06278_),
    .B1(net4879));
 sg13g2_nor2_1 _15675_ (.A(\m_sys._m_gpio8_io_b_mem_rdata[1] ),
    .B(_03512_),
    .Y(_06279_));
 sg13g2_o21ai_1 _15676_ (.B1(_04834_),
    .Y(_06280_),
    .A1(\m_sys._m_uart_io_b_mem_rdata[1] ),
    .A2(net4880));
 sg13g2_o21ai_1 _15677_ (.B1(net5275),
    .Y(_06281_),
    .A1(_06279_),
    .A2(_06280_));
 sg13g2_a21oi_1 _15678_ (.A1(_06277_),
    .A2(_06278_),
    .Y(_06282_),
    .B1(net5000));
 sg13g2_a22oi_1 _15679_ (.Y(_06283_),
    .B1(_06281_),
    .B2(_06282_),
    .A2(net5000),
    .A1(\m_sys._m_uart_io_o_bl_data[1] ));
 sg13g2_a22oi_1 _15680_ (.Y(_01041_),
    .B1(_06263_),
    .B2(_06283_),
    .A2(_06262_),
    .A1(_02404_));
 sg13g2_nor2_1 _15681_ (.A(\m_sys._m_gpio8_io_b_mem_rdata[2] ),
    .B(_03512_),
    .Y(_06284_));
 sg13g2_o21ai_1 _15682_ (.B1(_04799_),
    .Y(_06285_),
    .A1(\m_sys._m_uart_io_b_mem_rdata[2] ),
    .A2(net4881));
 sg13g2_o21ai_1 _15683_ (.B1(net5276),
    .Y(_06286_),
    .A1(_06284_),
    .A2(_06285_));
 sg13g2_nor2b_1 _15684_ (.A(\m_sys._m_uart_io_b_mem_rdata[2] ),
    .B_N(net4999),
    .Y(_06287_));
 sg13g2_o21ai_1 _15685_ (.B1(_02717_),
    .Y(_06288_),
    .A1(\m_sys._m_gpio8_io_b_mem_rdata[2] ),
    .A2(net4999));
 sg13g2_a21oi_1 _15686_ (.A1(\m_sys._m_ram_io_b_port_rdata[2] ),
    .A2(_02716_),
    .Y(_06289_),
    .B1(net4879));
 sg13g2_o21ai_1 _15687_ (.B1(_06289_),
    .Y(_06290_),
    .A1(_06287_),
    .A2(_06288_));
 sg13g2_a21oi_1 _15688_ (.A1(_06286_),
    .A2(_06290_),
    .Y(_06291_),
    .B1(net5001));
 sg13g2_o21ai_1 _15689_ (.B1(_06263_),
    .Y(_06292_),
    .A1(net5265),
    .A2(_06113_));
 sg13g2_nand2_1 _15690_ (.Y(_06293_),
    .A(net3339),
    .B(_06262_));
 sg13g2_o21ai_1 _15691_ (.B1(_06293_),
    .Y(_01042_),
    .A1(_06291_),
    .A2(_06292_));
 sg13g2_mux2_1 _15692_ (.A0(\m_sys._m_gpio8_io_b_mem_rdata[3] ),
    .A1(\m_sys._m_uart_io_b_mem_rdata[3] ),
    .S(net4999),
    .X(_06294_));
 sg13g2_nand2_1 _15693_ (.Y(_06295_),
    .A(_02717_),
    .B(_06294_));
 sg13g2_a21oi_1 _15694_ (.A1(\m_sys._m_ram_io_b_port_rdata[3] ),
    .A2(net5140),
    .Y(_06296_),
    .B1(net4878));
 sg13g2_nor2_1 _15695_ (.A(\m_sys._m_gpio8_io_b_mem_rdata[3] ),
    .B(_03512_),
    .Y(_06297_));
 sg13g2_o21ai_1 _15696_ (.B1(_04763_),
    .Y(_06298_),
    .A1(\m_sys._m_uart_io_b_mem_rdata[3] ),
    .A2(net4880));
 sg13g2_o21ai_1 _15697_ (.B1(net5275),
    .Y(_06299_),
    .A1(_06297_),
    .A2(_06298_));
 sg13g2_a21oi_1 _15698_ (.A1(_06295_),
    .A2(_06296_),
    .Y(_06300_),
    .B1(net5000));
 sg13g2_a22oi_1 _15699_ (.Y(_06301_),
    .B1(_06299_),
    .B2(_06300_),
    .A2(net5000),
    .A1(net5264));
 sg13g2_a22oi_1 _15700_ (.Y(_01043_),
    .B1(_06263_),
    .B2(_06301_),
    .A2(net4382),
    .A1(_02405_));
 sg13g2_nor2_1 _15701_ (.A(\m_sys._m_gpio8_io_b_mem_rdata[4] ),
    .B(_03512_),
    .Y(_06302_));
 sg13g2_o21ai_1 _15702_ (.B1(_04723_),
    .Y(_06303_),
    .A1(\m_sys._m_uart_io_b_mem_rdata[4] ),
    .A2(net4880));
 sg13g2_o21ai_1 _15703_ (.B1(net5275),
    .Y(_06304_),
    .A1(_06302_),
    .A2(_06303_));
 sg13g2_nor2b_1 _15704_ (.A(\m_sys._m_uart_io_b_mem_rdata[4] ),
    .B_N(net4999),
    .Y(_06305_));
 sg13g2_o21ai_1 _15705_ (.B1(_02717_),
    .Y(_06306_),
    .A1(\m_sys._m_gpio8_io_b_mem_rdata[4] ),
    .A2(net4998));
 sg13g2_a21oi_1 _15706_ (.A1(\m_sys._m_ram_io_b_port_rdata[4] ),
    .A2(net5140),
    .Y(_06307_),
    .B1(net4878));
 sg13g2_o21ai_1 _15707_ (.B1(_06307_),
    .Y(_06308_),
    .A1(_06305_),
    .A2(_06306_));
 sg13g2_a21oi_1 _15708_ (.A1(_06304_),
    .A2(_06308_),
    .Y(_06309_),
    .B1(net5001));
 sg13g2_o21ai_1 _15709_ (.B1(_06263_),
    .Y(_06310_),
    .A1(net5263),
    .A2(_06113_));
 sg13g2_nand2_1 _15710_ (.Y(_06311_),
    .A(net3244),
    .B(net4382));
 sg13g2_o21ai_1 _15711_ (.B1(_06311_),
    .Y(_01044_),
    .A1(_06309_),
    .A2(_06310_));
 sg13g2_mux2_1 _15712_ (.A0(\m_sys._m_gpio8_io_b_mem_rdata[5] ),
    .A1(\m_sys._m_uart_io_b_mem_rdata[5] ),
    .S(net4998),
    .X(_06312_));
 sg13g2_nand2_1 _15713_ (.Y(_06313_),
    .A(_02717_),
    .B(_06312_));
 sg13g2_a21oi_1 _15714_ (.A1(\m_sys._m_ram_io_b_port_rdata[5] ),
    .A2(net5140),
    .Y(_06314_),
    .B1(net4878));
 sg13g2_nor2_1 _15715_ (.A(\m_sys._m_gpio8_io_b_mem_rdata[5] ),
    .B(_03512_),
    .Y(_06315_));
 sg13g2_o21ai_1 _15716_ (.B1(_04661_),
    .Y(_06316_),
    .A1(\m_sys._m_uart_io_b_mem_rdata[5] ),
    .A2(net4880));
 sg13g2_o21ai_1 _15717_ (.B1(net5275),
    .Y(_06317_),
    .A1(_06315_),
    .A2(_06316_));
 sg13g2_a21oi_1 _15718_ (.A1(_06313_),
    .A2(_06314_),
    .Y(_06318_),
    .B1(net5000));
 sg13g2_a22oi_1 _15719_ (.Y(_06319_),
    .B1(_06317_),
    .B2(_06318_),
    .A2(net5000),
    .A1(net5262));
 sg13g2_a22oi_1 _15720_ (.Y(_01045_),
    .B1(_06263_),
    .B2(_06319_),
    .A2(net4382),
    .A1(_02406_));
 sg13g2_nor2_1 _15721_ (.A(\m_sys._m_gpio8_io_b_mem_rdata[6] ),
    .B(_03512_),
    .Y(_06320_));
 sg13g2_o21ai_1 _15722_ (.B1(_04640_),
    .Y(_06321_),
    .A1(\m_sys._m_uart_io_b_mem_rdata[6] ),
    .A2(net4880));
 sg13g2_o21ai_1 _15723_ (.B1(net5275),
    .Y(_06322_),
    .A1(_06320_),
    .A2(_06321_));
 sg13g2_nor2b_1 _15724_ (.A(\m_sys._m_uart_io_b_mem_rdata[6] ),
    .B_N(net4998),
    .Y(_06323_));
 sg13g2_o21ai_1 _15725_ (.B1(_02717_),
    .Y(_06324_),
    .A1(\m_sys._m_gpio8_io_b_mem_rdata[6] ),
    .A2(net4998));
 sg13g2_a21oi_1 _15726_ (.A1(\m_sys._m_ram_io_b_port_rdata[6] ),
    .A2(net5140),
    .Y(_06325_),
    .B1(net4878));
 sg13g2_o21ai_1 _15727_ (.B1(_06325_),
    .Y(_06326_),
    .A1(_06323_),
    .A2(_06324_));
 sg13g2_a21oi_1 _15728_ (.A1(_06322_),
    .A2(_06326_),
    .Y(_06327_),
    .B1(net5001));
 sg13g2_o21ai_1 _15729_ (.B1(_06263_),
    .Y(_06328_),
    .A1(net5261),
    .A2(_06113_));
 sg13g2_nand2_1 _15730_ (.Y(_06329_),
    .A(net3286),
    .B(net4382));
 sg13g2_o21ai_1 _15731_ (.B1(_06329_),
    .Y(_01046_),
    .A1(_06327_),
    .A2(_06328_));
 sg13g2_nand2b_1 _15732_ (.Y(_06330_),
    .B(_02418_),
    .A_N(net4998));
 sg13g2_a21oi_1 _15733_ (.A1(_02417_),
    .A2(net4998),
    .Y(_06331_),
    .B1(net5140));
 sg13g2_a22oi_1 _15734_ (.Y(_06332_),
    .B1(_06330_),
    .B2(_06331_),
    .A2(net5140),
    .A1(\m_sys._m_ram_io_b_port_rdata[7] ));
 sg13g2_a21oi_1 _15735_ (.A1(_02418_),
    .A2(_03511_),
    .Y(_06333_),
    .B1(_03509_));
 sg13g2_o21ai_1 _15736_ (.B1(_06333_),
    .Y(_06334_),
    .A1(\m_sys._m_uart_io_b_mem_rdata[7] ),
    .A2(net4880));
 sg13g2_o21ai_1 _15737_ (.B1(_06334_),
    .Y(_06335_),
    .A1(net5274),
    .A2(_06332_));
 sg13g2_a21oi_1 _15738_ (.A1(_03501_),
    .A2(_06332_),
    .Y(_06336_),
    .B1(net5000));
 sg13g2_a221oi_1 _15739_ (.B2(_06336_),
    .C1(_06264_),
    .B1(_06335_),
    .A1(net5260),
    .Y(_06337_),
    .A2(net5000));
 sg13g2_a21oi_1 _15740_ (.A1(_02407_),
    .A2(net4382),
    .Y(_01047_),
    .B1(_06337_));
 sg13g2_nor2_1 _15741_ (.A(net4715),
    .B(_06116_),
    .Y(_06338_));
 sg13g2_nor2_1 _15742_ (.A(net2905),
    .B(_06338_),
    .Y(_06339_));
 sg13g2_a21oi_1 _15743_ (.A1(_02342_),
    .A2(net4447),
    .Y(_01048_),
    .B1(_06339_));
 sg13g2_nor2_1 _15744_ (.A(net2970),
    .B(_06338_),
    .Y(_06340_));
 sg13g2_a21oi_1 _15745_ (.A1(_02341_),
    .A2(net4447),
    .Y(_01049_),
    .B1(_06340_));
 sg13g2_mux2_1 _15746_ (.A0(net2882),
    .A1(net5265),
    .S(net4447),
    .X(_01050_));
 sg13g2_mux2_1 _15747_ (.A0(net2854),
    .A1(net5264),
    .S(net4447),
    .X(_01051_));
 sg13g2_mux2_1 _15748_ (.A0(net2799),
    .A1(net5263),
    .S(net4447),
    .X(_01052_));
 sg13g2_mux2_1 _15749_ (.A0(net2890),
    .A1(net5262),
    .S(net4447),
    .X(_01053_));
 sg13g2_mux2_1 _15750_ (.A0(net2891),
    .A1(net5261),
    .S(net4447),
    .X(_01054_));
 sg13g2_mux2_1 _15751_ (.A0(net2897),
    .A1(net5260),
    .S(net4447),
    .X(_01055_));
 sg13g2_nor2_1 _15752_ (.A(\m_sys.m_bootloader.r_byte_cnt[0] ),
    .B(net4715),
    .Y(_06341_));
 sg13g2_nand3_1 _15753_ (.B(_06083_),
    .C(_06341_),
    .A(_02361_),
    .Y(_06342_));
 sg13g2_nand2_1 _15754_ (.Y(_06343_),
    .A(net2044),
    .B(net4381));
 sg13g2_o21ai_1 _15755_ (.B1(_06343_),
    .Y(_01056_),
    .A1(_02342_),
    .A2(net4381));
 sg13g2_nand2_1 _15756_ (.Y(_06344_),
    .A(net1992),
    .B(net4381));
 sg13g2_o21ai_1 _15757_ (.B1(_06344_),
    .Y(_01057_),
    .A1(_02341_),
    .A2(net4381));
 sg13g2_mux2_1 _15758_ (.A0(net5265),
    .A1(net2917),
    .S(_06342_),
    .X(_01058_));
 sg13g2_mux2_1 _15759_ (.A0(net5264),
    .A1(net3041),
    .S(net4381),
    .X(_01059_));
 sg13g2_mux2_1 _15760_ (.A0(net5263),
    .A1(net3049),
    .S(net4381),
    .X(_01060_));
 sg13g2_mux2_1 _15761_ (.A0(net5262),
    .A1(net3072),
    .S(net4381),
    .X(_01061_));
 sg13g2_mux2_1 _15762_ (.A0(net5261),
    .A1(net3056),
    .S(net4381),
    .X(_01062_));
 sg13g2_mux2_1 _15763_ (.A0(net5260),
    .A1(net3045),
    .S(_06342_),
    .X(_01063_));
 sg13g2_nand2_1 _15764_ (.Y(_06345_),
    .A(\m_sys.m_bootloader.r_byte_cnt[0] ),
    .B(_06085_));
 sg13g2_nor3_2 _15765_ (.A(net5286),
    .B(_06082_),
    .C(_06345_),
    .Y(_06346_));
 sg13g2_nor2_1 _15766_ (.A(net2932),
    .B(_06346_),
    .Y(_06347_));
 sg13g2_a21oi_1 _15767_ (.A1(_02342_),
    .A2(_06346_),
    .Y(_01064_),
    .B1(_06347_));
 sg13g2_nor2_1 _15768_ (.A(net2578),
    .B(_06346_),
    .Y(_06348_));
 sg13g2_a21oi_1 _15769_ (.A1(_02341_),
    .A2(_06346_),
    .Y(_01065_),
    .B1(_06348_));
 sg13g2_mux2_1 _15770_ (.A0(net2613),
    .A1(net5265),
    .S(_06346_),
    .X(_01066_));
 sg13g2_mux2_1 _15771_ (.A0(net2896),
    .A1(net5264),
    .S(_06346_),
    .X(_01067_));
 sg13g2_nor2_2 _15772_ (.A(_02361_),
    .B(_06082_),
    .Y(_06349_));
 sg13g2_nand2_1 _15773_ (.Y(_06350_),
    .A(net5286),
    .B(_06083_));
 sg13g2_nand2_1 _15774_ (.Y(_06351_),
    .A(_06341_),
    .B(_06349_));
 sg13g2_nand2_1 _15775_ (.Y(_06352_),
    .A(net3144),
    .B(net4380));
 sg13g2_o21ai_1 _15776_ (.B1(_06352_),
    .Y(_01068_),
    .A1(_02342_),
    .A2(_06351_));
 sg13g2_nand2_1 _15777_ (.Y(_06353_),
    .A(net3151),
    .B(net4380));
 sg13g2_o21ai_1 _15778_ (.B1(_06353_),
    .Y(_01069_),
    .A1(_02341_),
    .A2(_06351_));
 sg13g2_mux2_1 _15779_ (.A0(net5265),
    .A1(net3184),
    .S(net4380),
    .X(_01070_));
 sg13g2_mux2_1 _15780_ (.A0(net5264),
    .A1(net3212),
    .S(net4380),
    .X(_01071_));
 sg13g2_mux2_1 _15781_ (.A0(net5263),
    .A1(net3369),
    .S(net4380),
    .X(_01072_));
 sg13g2_mux2_1 _15782_ (.A0(net5262),
    .A1(net3239),
    .S(net4380),
    .X(_01073_));
 sg13g2_mux2_1 _15783_ (.A0(net5261),
    .A1(net2948),
    .S(net4380),
    .X(_01074_));
 sg13g2_mux2_1 _15784_ (.A0(net5260),
    .A1(net3188),
    .S(net4380),
    .X(_01075_));
 sg13g2_nor2_2 _15785_ (.A(_06345_),
    .B(_06350_),
    .Y(_06354_));
 sg13g2_nor2_1 _15786_ (.A(net3067),
    .B(net4354),
    .Y(_06355_));
 sg13g2_a21oi_1 _15787_ (.A1(_02342_),
    .A2(_06354_),
    .Y(_01076_),
    .B1(_06355_));
 sg13g2_nor2_1 _15788_ (.A(net3087),
    .B(_06354_),
    .Y(_06356_));
 sg13g2_a21oi_1 _15789_ (.A1(_02341_),
    .A2(net4354),
    .Y(_01077_),
    .B1(_06356_));
 sg13g2_mux2_1 _15790_ (.A0(net3280),
    .A1(net5265),
    .S(net4354),
    .X(_01078_));
 sg13g2_mux2_1 _15791_ (.A0(net3160),
    .A1(net5264),
    .S(net4354),
    .X(_01079_));
 sg13g2_mux2_1 _15792_ (.A0(net3154),
    .A1(net5263),
    .S(net4354),
    .X(_01080_));
 sg13g2_mux2_1 _15793_ (.A0(net3088),
    .A1(net5262),
    .S(net4354),
    .X(_01081_));
 sg13g2_mux2_1 _15794_ (.A0(net3091),
    .A1(net5261),
    .S(net4354),
    .X(_01082_));
 sg13g2_mux2_1 _15795_ (.A0(net2927),
    .A1(net5260),
    .S(net4354),
    .X(_01083_));
 sg13g2_o21ai_1 _15796_ (.B1(net5384),
    .Y(_01084_),
    .A1(net5234),
    .A2(_06123_));
 sg13g2_nor2_2 _15797_ (.A(net4715),
    .B(_06207_),
    .Y(_06357_));
 sg13g2_nor2_1 _15798_ (.A(net3195),
    .B(_06357_),
    .Y(_06358_));
 sg13g2_a21oi_1 _15799_ (.A1(net2522),
    .A2(_06357_),
    .Y(_01085_),
    .B1(net3196));
 sg13g2_nor3_1 _15800_ (.A(_06100_),
    .B(_06211_),
    .C(_06349_),
    .Y(_06359_));
 sg13g2_o21ai_1 _15801_ (.B1(_06359_),
    .Y(_06360_),
    .A1(_06099_),
    .A2(_06197_));
 sg13g2_nor2_1 _15802_ (.A(_04898_),
    .B(_06211_),
    .Y(_06361_));
 sg13g2_nand3_1 _15803_ (.B(_06360_),
    .C(_06361_),
    .A(_06214_),
    .Y(_06362_));
 sg13g2_nand2_1 _15804_ (.Y(_06363_),
    .A(net5267),
    .B(net4310));
 sg13g2_o21ai_1 _15805_ (.B1(net4712),
    .Y(_06364_),
    .A1(\m_sys.m_bootloader._GEN_22[0] ),
    .A2(net4383));
 sg13g2_a21oi_1 _15806_ (.A1(_02367_),
    .A2(net4383),
    .Y(_06365_),
    .B1(_06364_));
 sg13g2_a21oi_1 _15807_ (.A1(net1866),
    .A2(net4709),
    .Y(_06366_),
    .B1(_06365_));
 sg13g2_o21ai_1 _15808_ (.B1(_06363_),
    .Y(_01086_),
    .A1(net4310),
    .A2(net1867));
 sg13g2_nor2_1 _15809_ (.A(net1992),
    .B(net4383),
    .Y(_06367_));
 sg13g2_o21ai_1 _15810_ (.B1(net4711),
    .Y(_06368_),
    .A1(\m_sys._m_bootloader_io_b_mem_addr[1] ),
    .A2(_06096_));
 sg13g2_nor2_1 _15811_ (.A(net5143),
    .B(net4711),
    .Y(_06369_));
 sg13g2_o21ai_1 _15812_ (.B1(_06369_),
    .Y(_06370_),
    .A1(net3248),
    .A2(net5267));
 sg13g2_o21ai_1 _15813_ (.B1(_06370_),
    .Y(_06371_),
    .A1(_06367_),
    .A2(_06368_));
 sg13g2_mux2_1 _15814_ (.A0(_06371_),
    .A1(net3248),
    .S(net4310),
    .X(_01087_));
 sg13g2_nand2b_1 _15815_ (.Y(_06372_),
    .B(_06096_),
    .A_N(net2917));
 sg13g2_a21oi_1 _15816_ (.A1(_02373_),
    .A2(net4383),
    .Y(_06373_),
    .B1(net4710));
 sg13g2_xnor2_1 _15817_ (.Y(_06374_),
    .A(_02373_),
    .B(net5143));
 sg13g2_a221oi_1 _15818_ (.B2(net4710),
    .C1(net4311),
    .B1(_06374_),
    .A1(_06372_),
    .Y(_06375_),
    .A2(_06373_));
 sg13g2_a21oi_1 _15819_ (.A1(_02373_),
    .A2(net4311),
    .Y(_01088_),
    .B1(_06375_));
 sg13g2_mux2_1 _15820_ (.A0(\m_sys._m_bootloader_io_b_mem_addr[3] ),
    .A1(net3041),
    .S(_06096_),
    .X(_06376_));
 sg13g2_and3_1 _15821_ (.X(_06377_),
    .A(\m_sys._m_bootloader_io_b_mem_addr[2] ),
    .B(\m_sys._m_bootloader_io_b_mem_addr[3] ),
    .C(net5143));
 sg13g2_a21oi_1 _15822_ (.A1(\m_sys._m_bootloader_io_b_mem_addr[2] ),
    .A2(net5143),
    .Y(_06378_),
    .B1(net3101));
 sg13g2_nor3_1 _15823_ (.A(net4712),
    .B(_06377_),
    .C(_06378_),
    .Y(_06379_));
 sg13g2_a21oi_1 _15824_ (.A1(net4712),
    .A2(_06376_),
    .Y(_06380_),
    .B1(_06379_));
 sg13g2_nand2_1 _15825_ (.Y(_06381_),
    .A(net3101),
    .B(net4311));
 sg13g2_o21ai_1 _15826_ (.B1(_06381_),
    .Y(_01089_),
    .A1(net4311),
    .A2(_06380_));
 sg13g2_a21oi_1 _15827_ (.A1(_02370_),
    .A2(net4383),
    .Y(_06382_),
    .B1(net4709));
 sg13g2_o21ai_1 _15828_ (.B1(_06382_),
    .Y(_06383_),
    .A1(net3049),
    .A2(net4384));
 sg13g2_and2_1 _15829_ (.A(\m_sys._m_bootloader_io_b_mem_addr[4] ),
    .B(_06377_),
    .X(_06384_));
 sg13g2_o21ai_1 _15830_ (.B1(net4709),
    .Y(_06385_),
    .A1(\m_sys._m_bootloader_io_b_mem_addr[4] ),
    .A2(_06377_));
 sg13g2_o21ai_1 _15831_ (.B1(_06383_),
    .Y(_06386_),
    .A1(_06384_),
    .A2(_06385_));
 sg13g2_mux2_1 _15832_ (.A0(_06386_),
    .A1(net3370),
    .S(net4310),
    .X(_01090_));
 sg13g2_mux2_1 _15833_ (.A0(\m_sys._m_bootloader_io_b_mem_addr[5] ),
    .A1(net3072),
    .S(_06096_),
    .X(_06387_));
 sg13g2_nand2_2 _15834_ (.Y(_06388_),
    .A(\m_sys._m_bootloader_io_b_mem_addr[5] ),
    .B(_06384_));
 sg13g2_o21ai_1 _15835_ (.B1(net4709),
    .Y(_06389_),
    .A1(net3133),
    .A2(_06384_));
 sg13g2_nor2b_1 _15836_ (.A(_06389_),
    .B_N(_06388_),
    .Y(_06390_));
 sg13g2_a21oi_1 _15837_ (.A1(net4711),
    .A2(_06387_),
    .Y(_06391_),
    .B1(_06390_));
 sg13g2_nand2_1 _15838_ (.Y(_06392_),
    .A(net3133),
    .B(net4312));
 sg13g2_o21ai_1 _15839_ (.B1(_06392_),
    .Y(_01091_),
    .A1(net4310),
    .A2(_06391_));
 sg13g2_o21ai_1 _15840_ (.B1(net4711),
    .Y(_06393_),
    .A1(\m_sys.m_bootloader._GEN_22[6] ),
    .A2(net4383));
 sg13g2_a21oi_1 _15841_ (.A1(_02389_),
    .A2(net4384),
    .Y(_06394_),
    .B1(_06393_));
 sg13g2_nor2_1 _15842_ (.A(_02389_),
    .B(_06388_),
    .Y(_06395_));
 sg13g2_xnor2_1 _15843_ (.Y(_06396_),
    .A(net3037),
    .B(_06388_));
 sg13g2_a21oi_1 _15844_ (.A1(net4709),
    .A2(_06396_),
    .Y(_06397_),
    .B1(_06394_));
 sg13g2_nand2_1 _15845_ (.Y(_06398_),
    .A(net3037),
    .B(net4310));
 sg13g2_o21ai_1 _15846_ (.B1(_06398_),
    .Y(_01092_),
    .A1(net4310),
    .A2(_06397_));
 sg13g2_nand2_1 _15847_ (.Y(_06399_),
    .A(net3375),
    .B(net4384));
 sg13g2_a21oi_1 _15848_ (.A1(net3045),
    .A2(_06096_),
    .Y(_06400_),
    .B1(net4710));
 sg13g2_nor2_1 _15849_ (.A(_00045_),
    .B(_06388_),
    .Y(_06401_));
 sg13g2_xnor2_1 _15850_ (.Y(_06402_),
    .A(\m_sys._m_bootloader_io_b_mem_addr[7] ),
    .B(_06401_));
 sg13g2_a221oi_1 _15851_ (.B2(net4709),
    .C1(net4312),
    .B1(_06402_),
    .A1(_06399_),
    .Y(_06403_),
    .A2(_06400_));
 sg13g2_a21o_1 _15852_ (.A2(net4311),
    .A1(net3375),
    .B1(_06403_),
    .X(_01093_));
 sg13g2_mux2_1 _15853_ (.A0(\m_sys._m_bootloader_io_b_mem_addr[8] ),
    .A1(net2932),
    .S(_06096_),
    .X(_06404_));
 sg13g2_and3_1 _15854_ (.X(_06405_),
    .A(\m_sys._m_bootloader_io_b_mem_addr[8] ),
    .B(\m_sys._m_bootloader_io_b_mem_addr[7] ),
    .C(_06395_));
 sg13g2_a21oi_1 _15855_ (.A1(net3452),
    .A2(_06395_),
    .Y(_06406_),
    .B1(net3197));
 sg13g2_nor3_1 _15856_ (.A(net4711),
    .B(_06405_),
    .C(_06406_),
    .Y(_06407_));
 sg13g2_a21oi_1 _15857_ (.A1(net4711),
    .A2(_06404_),
    .Y(_06408_),
    .B1(_06407_));
 sg13g2_nand2_1 _15858_ (.Y(_06409_),
    .A(net3197),
    .B(net4311));
 sg13g2_o21ai_1 _15859_ (.B1(_06409_),
    .Y(_01094_),
    .A1(net4312),
    .A2(_06408_));
 sg13g2_nand2b_1 _15860_ (.Y(_06410_),
    .B(_06096_),
    .A_N(net2578));
 sg13g2_a21oi_1 _15861_ (.A1(_02388_),
    .A2(net4383),
    .Y(_06411_),
    .B1(net4710));
 sg13g2_xnor2_1 _15862_ (.Y(_06412_),
    .A(_02388_),
    .B(_06405_));
 sg13g2_a221oi_1 _15863_ (.B2(net4710),
    .C1(net4311),
    .B1(_06412_),
    .A1(_06410_),
    .Y(_06413_),
    .A2(_06411_));
 sg13g2_a21oi_1 _15864_ (.A1(_02388_),
    .A2(net4312),
    .Y(_01095_),
    .B1(_06413_));
 sg13g2_a21o_1 _15865_ (.A2(_06405_),
    .A1(\m_sys._m_bootloader_io_b_mem_addr[9] ),
    .B1(\m_sys._m_bootloader_io_b_mem_addr[10] ),
    .X(_06414_));
 sg13g2_nand3_1 _15866_ (.B(\m_sys._m_bootloader_io_b_mem_addr[9] ),
    .C(_06405_),
    .A(\m_sys._m_bootloader_io_b_mem_addr[10] ),
    .Y(_06415_));
 sg13g2_a21oi_1 _15867_ (.A1(_06414_),
    .A2(_06415_),
    .Y(_06416_),
    .B1(net4711));
 sg13g2_nand2_1 _15868_ (.Y(_06417_),
    .A(net2613),
    .B(_06096_));
 sg13g2_a21oi_1 _15869_ (.A1(\m_sys._m_bootloader_io_b_mem_addr[10] ),
    .A2(net4384),
    .Y(_06418_),
    .B1(net4709));
 sg13g2_a21oi_1 _15870_ (.A1(_06417_),
    .A2(_06418_),
    .Y(_06419_),
    .B1(_06416_));
 sg13g2_mux2_1 _15871_ (.A0(_06419_),
    .A1(net3354),
    .S(net4311),
    .X(_01096_));
 sg13g2_nand2_1 _15872_ (.Y(_06420_),
    .A(net3245),
    .B(net4313));
 sg13g2_o21ai_1 _15873_ (.B1(net4711),
    .Y(_06421_),
    .A1(net2896),
    .A2(net4383));
 sg13g2_a21oi_1 _15874_ (.A1(_02387_),
    .A2(net4384),
    .Y(_06422_),
    .B1(_06421_));
 sg13g2_xnor2_1 _15875_ (.Y(_06423_),
    .A(\m_sys._m_bootloader_io_b_mem_addr[11] ),
    .B(_06415_));
 sg13g2_a21oi_1 _15876_ (.A1(net4709),
    .A2(_06423_),
    .Y(_06424_),
    .B1(_06422_));
 sg13g2_o21ai_1 _15877_ (.B1(_06420_),
    .Y(_01097_),
    .A1(net4310),
    .A2(_06424_));
 sg13g2_a22oi_1 _15878_ (.Y(_06425_),
    .B1(net4581),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][0] ),
    .A2(net4674),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][0] ));
 sg13g2_a22oi_1 _15879_ (.Y(_06426_),
    .B1(net4536),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][0] ),
    .A2(net4629),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][0] ));
 sg13g2_a21oi_1 _15880_ (.A1(_06425_),
    .A2(_06426_),
    .Y(_06427_),
    .B1(net4478));
 sg13g2_a22oi_1 _15881_ (.Y(_06428_),
    .B1(net4639),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][0] ),
    .A2(net4688),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][0] ));
 sg13g2_a22oi_1 _15882_ (.Y(_06429_),
    .B1(net4547),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][0] ),
    .A2(net4592),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][0] ));
 sg13g2_a21oi_2 _15883_ (.B1(net4504),
    .Y(_06430_),
    .A2(_06429_),
    .A1(_06428_));
 sg13g2_a22oi_1 _15884_ (.Y(_06431_),
    .B1(net4580),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][0] ),
    .A2(net4677),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][0] ));
 sg13g2_a22oi_1 _15885_ (.Y(_06432_),
    .B1(net4536),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][0] ),
    .A2(net4628),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][0] ));
 sg13g2_a21oi_1 _15886_ (.A1(_06431_),
    .A2(_06432_),
    .Y(_06433_),
    .B1(net4473));
 sg13g2_nor3_2 _15887_ (.A(_06427_),
    .B(_06430_),
    .C(_06433_),
    .Y(_06434_));
 sg13g2_a22oi_1 _15888_ (.Y(_06435_),
    .B1(net4531),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][0] ),
    .A2(net4623),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][0] ));
 sg13g2_a22oi_1 _15889_ (.Y(_06436_),
    .B1(net4576),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][0] ),
    .A2(net4676),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][0] ));
 sg13g2_a21o_1 _15890_ (.A2(_06436_),
    .A1(_06435_),
    .B1(net4483),
    .X(_06437_));
 sg13g2_a22oi_1 _15891_ (.Y(_06438_),
    .B1(net4587),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][0] ),
    .A2(net4681),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][0] ));
 sg13g2_a22oi_1 _15892_ (.Y(_06439_),
    .B1(net4542),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][0] ),
    .A2(net4634),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][0] ));
 sg13g2_a21oi_1 _15893_ (.A1(_06438_),
    .A2(_06439_),
    .Y(_06440_),
    .B1(net4466));
 sg13g2_a22oi_1 _15894_ (.Y(_06441_),
    .B1(net4541),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][0] ),
    .A2(net4586),
    .A1(\m_sys.m_ram.m_ram.r_mem[14][0] ));
 sg13g2_a22oi_1 _15895_ (.Y(_06442_),
    .B1(net4633),
    .B2(\m_sys.m_ram.m_ram.r_mem[12][0] ),
    .A2(net4689),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][0] ));
 sg13g2_a21oi_2 _15896_ (.B1(net4491),
    .Y(_06443_),
    .A2(_06442_),
    .A1(_06441_));
 sg13g2_a22oi_1 _15897_ (.Y(_06444_),
    .B1(net4546),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][0] ),
    .A2(net4591),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][0] ));
 sg13g2_a22oi_1 _15898_ (.Y(_06445_),
    .B1(net4638),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][0] ),
    .A2(net4686),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][0] ));
 sg13g2_a21oi_2 _15899_ (.B1(net4452),
    .Y(_06446_),
    .A2(_06445_),
    .A1(_06444_));
 sg13g2_a22oi_1 _15900_ (.Y(_06447_),
    .B1(net4546),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][0] ),
    .A2(net4591),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][0] ));
 sg13g2_a22oi_1 _15901_ (.Y(_06448_),
    .B1(net4638),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][0] ),
    .A2(net4686),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][0] ));
 sg13g2_a21oi_2 _15902_ (.B1(net4460),
    .Y(_06449_),
    .A2(_06448_),
    .A1(_06447_));
 sg13g2_nor4_2 _15903_ (.A(_06440_),
    .B(_06443_),
    .C(_06446_),
    .Y(_06450_),
    .D(_06449_));
 sg13g2_nand4_1 _15904_ (.B(_06434_),
    .C(_06437_),
    .A(net4365),
    .Y(_06451_),
    .D(_06450_));
 sg13g2_o21ai_1 _15905_ (.B1(_06451_),
    .Y(_06452_),
    .A1(net3308),
    .A2(net4359));
 sg13g2_nor2_1 _15906_ (.A(net5371),
    .B(_06452_),
    .Y(_01098_));
 sg13g2_a22oi_1 _15907_ (.Y(_06453_),
    .B1(net4593),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][1] ),
    .A2(net4688),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][1] ));
 sg13g2_a22oi_1 _15908_ (.Y(_06454_),
    .B1(net4548),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][1] ),
    .A2(net4640),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][1] ));
 sg13g2_a21oi_1 _15909_ (.A1(_06453_),
    .A2(_06454_),
    .Y(_06455_),
    .B1(net4504));
 sg13g2_a22oi_1 _15910_ (.Y(_06456_),
    .B1(net4623),
    .B2(\m_sys.m_ram.m_ram.r_mem[0][1] ),
    .A2(net4676),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][1] ));
 sg13g2_a22oi_1 _15911_ (.Y(_06457_),
    .B1(net4531),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][1] ),
    .A2(net4577),
    .A1(\m_sys.m_ram.m_ram.r_mem[2][1] ));
 sg13g2_a21oi_2 _15912_ (.B1(net4483),
    .Y(_06458_),
    .A2(_06457_),
    .A1(_06456_));
 sg13g2_a22oi_1 _15913_ (.Y(_06459_),
    .B1(net4586),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][1] ),
    .A2(net4681),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][1] ));
 sg13g2_a22oi_1 _15914_ (.Y(_06460_),
    .B1(net4541),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][1] ),
    .A2(net4633),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][1] ));
 sg13g2_a21oi_1 _15915_ (.A1(_06459_),
    .A2(_06460_),
    .Y(_06461_),
    .B1(net4478));
 sg13g2_a22oi_1 _15916_ (.Y(_06462_),
    .B1(net4593),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][1] ),
    .A2(net4688),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][1] ));
 sg13g2_a22oi_1 _15917_ (.Y(_06463_),
    .B1(net4548),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][1] ),
    .A2(net4640),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][1] ));
 sg13g2_a21oi_1 _15918_ (.A1(_06462_),
    .A2(_06463_),
    .Y(_06464_),
    .B1(net4460));
 sg13g2_a22oi_1 _15919_ (.Y(_06465_),
    .B1(net4587),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][1] ),
    .A2(net4689),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][1] ));
 sg13g2_a22oi_1 _15920_ (.Y(_06466_),
    .B1(net4542),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][1] ),
    .A2(net4634),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][1] ));
 sg13g2_a21oi_1 _15921_ (.A1(_06465_),
    .A2(_06466_),
    .Y(_06467_),
    .B1(net4466));
 sg13g2_a22oi_1 _15922_ (.Y(_06468_),
    .B1(net4541),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][1] ),
    .A2(net4689),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][1] ));
 sg13g2_a22oi_1 _15923_ (.Y(_06469_),
    .B1(net4587),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][1] ),
    .A2(net4633),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][1] ));
 sg13g2_a21o_1 _15924_ (.A2(_06469_),
    .A1(_06468_),
    .B1(net4491),
    .X(_06470_));
 sg13g2_a22oi_1 _15925_ (.Y(_06471_),
    .B1(net4548),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][1] ),
    .A2(net4593),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][1] ));
 sg13g2_a22oi_1 _15926_ (.Y(_06472_),
    .B1(net4640),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][1] ),
    .A2(net4685),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][1] ));
 sg13g2_a21oi_2 _15927_ (.B1(net4452),
    .Y(_06473_),
    .A2(_06472_),
    .A1(_06471_));
 sg13g2_a22oi_1 _15928_ (.Y(_06474_),
    .B1(net4580),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][1] ),
    .A2(net4677),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][1] ));
 sg13g2_a22oi_1 _15929_ (.Y(_06475_),
    .B1(net4535),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][1] ),
    .A2(net4628),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][1] ));
 sg13g2_a21oi_2 _15930_ (.B1(net4473),
    .Y(_06476_),
    .A2(_06475_),
    .A1(_06474_));
 sg13g2_nor3_2 _15931_ (.A(_06455_),
    .B(_06458_),
    .C(_06473_),
    .Y(_06477_));
 sg13g2_nor4_1 _15932_ (.A(_06461_),
    .B(_06464_),
    .C(_06467_),
    .D(_06476_),
    .Y(_06478_));
 sg13g2_nand4_1 _15933_ (.B(_06470_),
    .C(_06477_),
    .A(net4364),
    .Y(_06479_),
    .D(_06478_));
 sg13g2_o21ai_1 _15934_ (.B1(_06479_),
    .Y(_06480_),
    .A1(net3342),
    .A2(net4358));
 sg13g2_nor2_1 _15935_ (.A(net5371),
    .B(_06480_),
    .Y(_01099_));
 sg13g2_a22oi_1 _15936_ (.Y(_06481_),
    .B1(net4532),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][2] ),
    .A2(net4669),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][2] ));
 sg13g2_a22oi_1 _15937_ (.Y(_06482_),
    .B1(net4577),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][2] ),
    .A2(net4624),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][2] ));
 sg13g2_a21oi_1 _15938_ (.A1(_06481_),
    .A2(_06482_),
    .Y(_06483_),
    .B1(net4472));
 sg13g2_a22oi_1 _15939_ (.Y(_06484_),
    .B1(net4637),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][2] ),
    .A2(net4686),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][2] ));
 sg13g2_a22oi_1 _15940_ (.Y(_06485_),
    .B1(net4545),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][2] ),
    .A2(net4591),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][2] ));
 sg13g2_a21oi_1 _15941_ (.A1(_06484_),
    .A2(_06485_),
    .Y(_06486_),
    .B1(net4453));
 sg13g2_a22oi_1 _15942_ (.Y(_06487_),
    .B1(net4580),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][2] ),
    .A2(net4673),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][2] ));
 sg13g2_a22oi_1 _15943_ (.Y(_06488_),
    .B1(net4535),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][2] ),
    .A2(net4628),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][2] ));
 sg13g2_a21oi_2 _15944_ (.B1(net4478),
    .Y(_06489_),
    .A2(_06488_),
    .A1(_06487_));
 sg13g2_a22oi_1 _15945_ (.Y(_06490_),
    .B1(net4546),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][2] ),
    .A2(net4638),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][2] ));
 sg13g2_a22oi_1 _15946_ (.Y(_06491_),
    .B1(net4591),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][2] ),
    .A2(net4685),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][2] ));
 sg13g2_a21oi_1 _15947_ (.A1(_06490_),
    .A2(_06491_),
    .Y(_06492_),
    .B1(net4460));
 sg13g2_a22oi_1 _15948_ (.Y(_06493_),
    .B1(net4571),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][2] ),
    .A2(net4663),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][2] ));
 sg13g2_a22oi_1 _15949_ (.Y(_06494_),
    .B1(net4531),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][2] ),
    .A2(net4623),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][2] ));
 sg13g2_a21oi_2 _15950_ (.B1(net4483),
    .Y(_06495_),
    .A2(_06494_),
    .A1(_06493_));
 sg13g2_a22oi_1 _15951_ (.Y(_06496_),
    .B1(net4541),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][2] ),
    .A2(net4586),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][2] ));
 sg13g2_a22oi_1 _15952_ (.Y(_06497_),
    .B1(net4633),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][2] ),
    .A2(net4681),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][2] ));
 sg13g2_a21o_1 _15953_ (.A2(_06497_),
    .A1(_06496_),
    .B1(net4466),
    .X(_06498_));
 sg13g2_a22oi_1 _15954_ (.Y(_06499_),
    .B1(net4547),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][2] ),
    .A2(net4592),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][2] ));
 sg13g2_a22oi_1 _15955_ (.Y(_06500_),
    .B1(net4639),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][2] ),
    .A2(net4688),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][2] ));
 sg13g2_a21oi_1 _15956_ (.A1(_06499_),
    .A2(_06500_),
    .Y(_06501_),
    .B1(net4504));
 sg13g2_a22oi_1 _15957_ (.Y(_06502_),
    .B1(net4577),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][2] ),
    .A2(net4676),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][2] ));
 sg13g2_a22oi_1 _15958_ (.Y(_06503_),
    .B1(net4532),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][2] ),
    .A2(net4624),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][2] ));
 sg13g2_a21oi_1 _15959_ (.A1(_06502_),
    .A2(_06503_),
    .Y(_06504_),
    .B1(net4490));
 sg13g2_nor3_2 _15960_ (.A(_06486_),
    .B(_06492_),
    .C(_06501_),
    .Y(_06505_));
 sg13g2_nor4_2 _15961_ (.A(_06483_),
    .B(_06489_),
    .C(_06495_),
    .Y(_06506_),
    .D(_06504_));
 sg13g2_nand4_1 _15962_ (.B(_06498_),
    .C(_06505_),
    .A(net4363),
    .Y(_06507_),
    .D(_06506_));
 sg13g2_o21ai_1 _15963_ (.B1(_06507_),
    .Y(_06508_),
    .A1(net3324),
    .A2(net4358));
 sg13g2_nor2_1 _15964_ (.A(net5371),
    .B(_06508_),
    .Y(_01100_));
 sg13g2_a22oi_1 _15965_ (.Y(_06509_),
    .B1(net4586),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][3] ),
    .A2(net4681),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][3] ));
 sg13g2_a22oi_1 _15966_ (.Y(_06510_),
    .B1(net4541),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][3] ),
    .A2(net4633),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][3] ));
 sg13g2_a21oi_2 _15967_ (.B1(net4478),
    .Y(_06511_),
    .A2(_06510_),
    .A1(_06509_));
 sg13g2_a22oi_1 _15968_ (.Y(_06512_),
    .B1(net4591),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][3] ),
    .A2(net4685),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][3] ));
 sg13g2_a22oi_1 _15969_ (.Y(_06513_),
    .B1(net4546),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][3] ),
    .A2(net4638),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][3] ));
 sg13g2_a21oi_1 _15970_ (.A1(_06512_),
    .A2(_06513_),
    .Y(_06514_),
    .B1(net4460));
 sg13g2_a22oi_1 _15971_ (.Y(_06515_),
    .B1(net4546),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][3] ),
    .A2(net4688),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][3] ));
 sg13g2_a22oi_1 _15972_ (.Y(_06516_),
    .B1(net4591),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][3] ),
    .A2(net4638),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][3] ));
 sg13g2_a21oi_1 _15973_ (.A1(_06515_),
    .A2(_06516_),
    .Y(_06517_),
    .B1(net4504));
 sg13g2_nor3_2 _15974_ (.A(_06511_),
    .B(_06514_),
    .C(_06517_),
    .Y(_06518_));
 sg13g2_a22oi_1 _15975_ (.Y(_06519_),
    .B1(net4571),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][3] ),
    .A2(net4663),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][3] ));
 sg13g2_a22oi_1 _15976_ (.Y(_06520_),
    .B1(net4526),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][3] ),
    .A2(net4619),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][3] ));
 sg13g2_a21o_1 _15977_ (.A2(_06520_),
    .A1(_06519_),
    .B1(net4482),
    .X(_06521_));
 sg13g2_a22oi_1 _15978_ (.Y(_06522_),
    .B1(net4548),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][3] ),
    .A2(net4593),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][3] ));
 sg13g2_a22oi_1 _15979_ (.Y(_06523_),
    .B1(net4640),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][3] ),
    .A2(net4685),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][3] ));
 sg13g2_a21oi_2 _15980_ (.B1(net4451),
    .Y(_06524_),
    .A2(_06523_),
    .A1(_06522_));
 sg13g2_a22oi_1 _15981_ (.Y(_06525_),
    .B1(net4577),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][3] ),
    .A2(net4676),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][3] ));
 sg13g2_a22oi_1 _15982_ (.Y(_06526_),
    .B1(net4532),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][3] ),
    .A2(net4624),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][3] ));
 sg13g2_a21oi_2 _15983_ (.B1(net4472),
    .Y(_06527_),
    .A2(_06526_),
    .A1(_06525_));
 sg13g2_a22oi_1 _15984_ (.Y(_06528_),
    .B1(net4628),
    .B2(\m_sys.m_ram.m_ram.r_mem[12][3] ),
    .A2(net4677),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][3] ));
 sg13g2_a22oi_1 _15985_ (.Y(_06529_),
    .B1(net4535),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][3] ),
    .A2(net4580),
    .A1(\m_sys.m_ram.m_ram.r_mem[14][3] ));
 sg13g2_a21oi_1 _15986_ (.A1(_06528_),
    .A2(_06529_),
    .Y(_06530_),
    .B1(net4489));
 sg13g2_a22oi_1 _15987_ (.Y(_06531_),
    .B1(net4536),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][3] ),
    .A2(net4581),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][3] ));
 sg13g2_a22oi_1 _15988_ (.Y(_06532_),
    .B1(net4629),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][3] ),
    .A2(net4677),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][3] ));
 sg13g2_a21oi_1 _15989_ (.A1(_06531_),
    .A2(_06532_),
    .Y(_06533_),
    .B1(net4465));
 sg13g2_nor4_2 _15990_ (.A(_06524_),
    .B(_06527_),
    .C(_06530_),
    .Y(_06534_),
    .D(_06533_));
 sg13g2_nand4_1 _15991_ (.B(_06518_),
    .C(_06521_),
    .A(net4365),
    .Y(_06535_),
    .D(_06534_));
 sg13g2_o21ai_1 _15992_ (.B1(_06535_),
    .Y(_06536_),
    .A1(net3318),
    .A2(net4358));
 sg13g2_nor2_1 _15993_ (.A(net5371),
    .B(_06536_),
    .Y(_01101_));
 sg13g2_a22oi_1 _15994_ (.Y(_06537_),
    .B1(net4586),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][4] ),
    .A2(net4689),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][4] ));
 sg13g2_a22oi_1 _15995_ (.Y(_06538_),
    .B1(net4541),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][4] ),
    .A2(net4633),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][4] ));
 sg13g2_a21oi_2 _15996_ (.B1(net4489),
    .Y(_06539_),
    .A2(_06538_),
    .A1(_06537_));
 sg13g2_a22oi_1 _15997_ (.Y(_06540_),
    .B1(net4546),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][4] ),
    .A2(net4638),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][4] ));
 sg13g2_a22oi_1 _15998_ (.Y(_06541_),
    .B1(net4592),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][4] ),
    .A2(net4690),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][4] ));
 sg13g2_a21oi_1 _15999_ (.A1(_06540_),
    .A2(_06541_),
    .Y(_06542_),
    .B1(net4504));
 sg13g2_a22oi_1 _16000_ (.Y(_06543_),
    .B1(net4592),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][4] ),
    .A2(net4688),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][4] ));
 sg13g2_a22oi_1 _16001_ (.Y(_06544_),
    .B1(net4547),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][4] ),
    .A2(net4639),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][4] ));
 sg13g2_a21oi_1 _16002_ (.A1(_06543_),
    .A2(_06544_),
    .Y(_06545_),
    .B1(net4460));
 sg13g2_nor3_2 _16003_ (.A(_06539_),
    .B(_06542_),
    .C(_06545_),
    .Y(_06546_));
 sg13g2_a22oi_1 _16004_ (.Y(_06547_),
    .B1(net4576),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][4] ),
    .A2(net4676),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][4] ));
 sg13g2_a22oi_1 _16005_ (.Y(_06548_),
    .B1(net4526),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][4] ),
    .A2(net4618),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][4] ));
 sg13g2_a21o_1 _16006_ (.A2(_06548_),
    .A1(_06547_),
    .B1(net4482),
    .X(_06549_));
 sg13g2_a22oi_1 _16007_ (.Y(_06550_),
    .B1(net4536),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][4] ),
    .A2(net4581),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][4] ));
 sg13g2_a22oi_1 _16008_ (.Y(_06551_),
    .B1(net4629),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][4] ),
    .A2(net4677),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][4] ));
 sg13g2_a21oi_1 _16009_ (.A1(_06550_),
    .A2(_06551_),
    .Y(_06552_),
    .B1(net4465));
 sg13g2_a22oi_1 _16010_ (.Y(_06553_),
    .B1(net4535),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][4] ),
    .A2(net4673),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][4] ));
 sg13g2_a22oi_1 _16011_ (.Y(_06554_),
    .B1(net4580),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][4] ),
    .A2(net4628),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][4] ));
 sg13g2_a21oi_1 _16012_ (.A1(_06553_),
    .A2(_06554_),
    .Y(_06555_),
    .B1(net4472));
 sg13g2_a22oi_1 _16013_ (.Y(_06556_),
    .B1(net4581),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][4] ),
    .A2(net4674),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][4] ));
 sg13g2_a22oi_1 _16014_ (.Y(_06557_),
    .B1(net4536),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][4] ),
    .A2(net4629),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][4] ));
 sg13g2_a21oi_1 _16015_ (.A1(_06556_),
    .A2(_06557_),
    .Y(_06558_),
    .B1(net4479));
 sg13g2_a22oi_1 _16016_ (.Y(_06559_),
    .B1(net4546),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][4] ),
    .A2(net4685),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][4] ));
 sg13g2_a22oi_1 _16017_ (.Y(_06560_),
    .B1(net4591),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][4] ),
    .A2(net4636),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][4] ));
 sg13g2_a21oi_2 _16018_ (.B1(net4451),
    .Y(_06561_),
    .A2(_06560_),
    .A1(_06559_));
 sg13g2_nor4_2 _16019_ (.A(_06552_),
    .B(_06555_),
    .C(_06558_),
    .Y(_06562_),
    .D(_06561_));
 sg13g2_nand4_1 _16020_ (.B(_06546_),
    .C(_06549_),
    .A(net4364),
    .Y(_06563_),
    .D(_06562_));
 sg13g2_o21ai_1 _16021_ (.B1(_06563_),
    .Y(_06564_),
    .A1(net3258),
    .A2(net4358));
 sg13g2_nor2_1 _16022_ (.A(net5371),
    .B(_06564_),
    .Y(_01102_));
 sg13g2_a22oi_1 _16023_ (.Y(_06565_),
    .B1(net4639),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][5] ),
    .A2(net4690),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][5] ));
 sg13g2_a22oi_1 _16024_ (.Y(_06566_),
    .B1(net4547),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][5] ),
    .A2(net4592),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][5] ));
 sg13g2_a21oi_1 _16025_ (.A1(_06565_),
    .A2(_06566_),
    .Y(_06567_),
    .B1(net4503));
 sg13g2_a22oi_1 _16026_ (.Y(_06568_),
    .B1(net4577),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][5] ),
    .A2(net4677),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][5] ));
 sg13g2_a22oi_1 _16027_ (.Y(_06569_),
    .B1(net4531),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][5] ),
    .A2(net4624),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][5] ));
 sg13g2_a21oi_1 _16028_ (.A1(_06568_),
    .A2(_06569_),
    .Y(_06570_),
    .B1(net4490));
 sg13g2_a22oi_1 _16029_ (.Y(_06571_),
    .B1(net4577),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][5] ),
    .A2(net4676),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][5] ));
 sg13g2_a22oi_1 _16030_ (.Y(_06572_),
    .B1(net4532),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][5] ),
    .A2(net4624),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][5] ));
 sg13g2_a21oi_1 _16031_ (.A1(_06571_),
    .A2(_06572_),
    .Y(_06573_),
    .B1(net4472));
 sg13g2_a22oi_1 _16032_ (.Y(_06574_),
    .B1(net4591),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][5] ),
    .A2(net4685),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][5] ));
 sg13g2_a22oi_1 _16033_ (.Y(_06575_),
    .B1(net4546),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][5] ),
    .A2(net4638),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][5] ));
 sg13g2_a21oi_1 _16034_ (.A1(_06574_),
    .A2(_06575_),
    .Y(_06576_),
    .B1(net4451));
 sg13g2_a22oi_1 _16035_ (.Y(_06577_),
    .B1(net4547),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][5] ),
    .A2(net4592),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][5] ));
 sg13g2_a22oi_1 _16036_ (.Y(_06578_),
    .B1(net4638),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][5] ),
    .A2(net4688),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][5] ));
 sg13g2_a21oi_1 _16037_ (.A1(_06577_),
    .A2(_06578_),
    .Y(_06579_),
    .B1(net4460));
 sg13g2_a22oi_1 _16038_ (.Y(_06580_),
    .B1(net4581),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][5] ),
    .A2(net4629),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][5] ));
 sg13g2_a22oi_1 _16039_ (.Y(_06581_),
    .B1(net4535),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][5] ),
    .A2(net4673),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][5] ));
 sg13g2_a21oi_2 _16040_ (.B1(net4478),
    .Y(_06582_),
    .A2(_06581_),
    .A1(_06580_));
 sg13g2_a22oi_1 _16041_ (.Y(_06583_),
    .B1(net4571),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][5] ),
    .A2(net4663),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][5] ));
 sg13g2_a22oi_1 _16042_ (.Y(_06584_),
    .B1(net4526),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][5] ),
    .A2(net4618),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][5] ));
 sg13g2_a21oi_2 _16043_ (.B1(net4482),
    .Y(_06585_),
    .A2(_06584_),
    .A1(_06583_));
 sg13g2_a22oi_1 _16044_ (.Y(_06586_),
    .B1(net4542),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][5] ),
    .A2(net4689),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][5] ));
 sg13g2_a22oi_1 _16045_ (.Y(_06587_),
    .B1(net4586),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][5] ),
    .A2(net4633),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][5] ));
 sg13g2_a21o_1 _16046_ (.A2(_06587_),
    .A1(_06586_),
    .B1(net4466),
    .X(_06588_));
 sg13g2_nor3_2 _16047_ (.A(_06567_),
    .B(_06576_),
    .C(_06579_),
    .Y(_06589_));
 sg13g2_nor4_2 _16048_ (.A(_06570_),
    .B(_06573_),
    .C(_06582_),
    .Y(_06590_),
    .D(_06585_));
 sg13g2_nand4_1 _16049_ (.B(_06588_),
    .C(_06589_),
    .A(net4364),
    .Y(_06591_),
    .D(_06590_));
 sg13g2_o21ai_1 _16050_ (.B1(_06591_),
    .Y(_06592_),
    .A1(net3362),
    .A2(net4358));
 sg13g2_nor2_1 _16051_ (.A(net5372),
    .B(_06592_),
    .Y(_01103_));
 sg13g2_a22oi_1 _16052_ (.Y(_06593_),
    .B1(net4640),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][6] ),
    .A2(net4688),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][6] ));
 sg13g2_a22oi_1 _16053_ (.Y(_06594_),
    .B1(net4548),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][6] ),
    .A2(net4593),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][6] ));
 sg13g2_a21oi_2 _16054_ (.B1(net4503),
    .Y(_06595_),
    .A2(_06594_),
    .A1(_06593_));
 sg13g2_a22oi_1 _16055_ (.Y(_06596_),
    .B1(net4535),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][6] ),
    .A2(net4678),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][6] ));
 sg13g2_a22oi_1 _16056_ (.Y(_06597_),
    .B1(net4580),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][6] ),
    .A2(net4628),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][6] ));
 sg13g2_a21oi_1 _16057_ (.A1(_06596_),
    .A2(_06597_),
    .Y(_06598_),
    .B1(net4472));
 sg13g2_a22oi_1 _16058_ (.Y(_06599_),
    .B1(net4586),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][6] ),
    .A2(net4689),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][6] ));
 sg13g2_a22oi_1 _16059_ (.Y(_06600_),
    .B1(net4541),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][6] ),
    .A2(net4629),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][6] ));
 sg13g2_a21oi_1 _16060_ (.A1(_06599_),
    .A2(_06600_),
    .Y(_06601_),
    .B1(net4489));
 sg13g2_a22oi_1 _16061_ (.Y(_06602_),
    .B1(net4531),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][6] ),
    .A2(net4623),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][6] ));
 sg13g2_a22oi_1 _16062_ (.Y(_06603_),
    .B1(net4576),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][6] ),
    .A2(net4676),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][6] ));
 sg13g2_a21oi_2 _16063_ (.B1(net4482),
    .Y(_06604_),
    .A2(_06603_),
    .A1(_06602_));
 sg13g2_a22oi_1 _16064_ (.Y(_06605_),
    .B1(net4542),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][6] ),
    .A2(net4587),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][6] ));
 sg13g2_a22oi_1 _16065_ (.Y(_06606_),
    .B1(net4634),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][6] ),
    .A2(net4682),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][6] ));
 sg13g2_a21oi_2 _16066_ (.B1(net4452),
    .Y(_06607_),
    .A2(_06606_),
    .A1(_06605_));
 sg13g2_a22oi_1 _16067_ (.Y(_06608_),
    .B1(net4593),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][6] ),
    .A2(net4685),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][6] ));
 sg13g2_a22oi_1 _16068_ (.Y(_06609_),
    .B1(net4548),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][6] ),
    .A2(net4640),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][6] ));
 sg13g2_a21oi_2 _16069_ (.B1(net4460),
    .Y(_06610_),
    .A2(_06609_),
    .A1(_06608_));
 sg13g2_a22oi_1 _16070_ (.Y(_06611_),
    .B1(net4581),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][6] ),
    .A2(net4673),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][6] ));
 sg13g2_a22oi_1 _16071_ (.Y(_06612_),
    .B1(net4536),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][6] ),
    .A2(net4629),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][6] ));
 sg13g2_a21oi_1 _16072_ (.A1(_06611_),
    .A2(_06612_),
    .Y(_06613_),
    .B1(net4477));
 sg13g2_a22oi_1 _16073_ (.Y(_06614_),
    .B1(net4542),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][6] ),
    .A2(net4587),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][6] ));
 sg13g2_a22oi_1 _16074_ (.Y(_06615_),
    .B1(net4634),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][6] ),
    .A2(net4689),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][6] ));
 sg13g2_a21o_1 _16075_ (.A2(_06615_),
    .A1(_06614_),
    .B1(net4466),
    .X(_06616_));
 sg13g2_nor3_1 _16076_ (.A(_06595_),
    .B(_06604_),
    .C(_06607_),
    .Y(_06617_));
 sg13g2_nor4_1 _16077_ (.A(_06598_),
    .B(_06601_),
    .C(_06610_),
    .D(_06613_),
    .Y(_06618_));
 sg13g2_nand4_1 _16078_ (.B(_06616_),
    .C(_06617_),
    .A(net4364),
    .Y(_06619_),
    .D(_06618_));
 sg13g2_o21ai_1 _16079_ (.B1(_06619_),
    .Y(_06620_),
    .A1(net3325),
    .A2(net4358));
 sg13g2_nor2_1 _16080_ (.A(net5371),
    .B(_06620_),
    .Y(_01104_));
 sg13g2_a22oi_1 _16081_ (.Y(_06621_),
    .B1(net4629),
    .B2(\m_sys.m_ram.m_ram.r_mem[12][7] ),
    .A2(net4677),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][7] ));
 sg13g2_a22oi_1 _16082_ (.Y(_06622_),
    .B1(net4536),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][7] ),
    .A2(net4581),
    .A1(\m_sys.m_ram.m_ram.r_mem[14][7] ));
 sg13g2_a21oi_1 _16083_ (.A1(_06621_),
    .A2(_06622_),
    .Y(_06623_),
    .B1(net4489));
 sg13g2_a22oi_1 _16084_ (.Y(_06624_),
    .B1(net4576),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][7] ),
    .A2(net4676),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][7] ));
 sg13g2_a22oi_1 _16085_ (.Y(_06625_),
    .B1(net4531),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][7] ),
    .A2(net4623),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][7] ));
 sg13g2_a21oi_2 _16086_ (.B1(net4482),
    .Y(_06626_),
    .A2(_06625_),
    .A1(_06624_));
 sg13g2_a22oi_1 _16087_ (.Y(_06627_),
    .B1(net4593),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][7] ),
    .A2(net4685),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][7] ));
 sg13g2_a22oi_1 _16088_ (.Y(_06628_),
    .B1(net4548),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][7] ),
    .A2(net4640),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][7] ));
 sg13g2_a21oi_2 _16089_ (.B1(net4460),
    .Y(_06629_),
    .A2(_06628_),
    .A1(_06627_));
 sg13g2_nor3_1 _16090_ (.A(_06623_),
    .B(_06626_),
    .C(_06629_),
    .Y(_06630_));
 sg13g2_a22oi_1 _16091_ (.Y(_06631_),
    .B1(net4634),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][7] ),
    .A2(net4689),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][7] ));
 sg13g2_a22oi_1 _16092_ (.Y(_06632_),
    .B1(net4542),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][7] ),
    .A2(net4587),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][7] ));
 sg13g2_a21o_1 _16093_ (.A2(_06632_),
    .A1(_06631_),
    .B1(net4505),
    .X(_06633_));
 sg13g2_a22oi_1 _16094_ (.Y(_06634_),
    .B1(net4586),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][7] ),
    .A2(net4681),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][7] ));
 sg13g2_a22oi_1 _16095_ (.Y(_06635_),
    .B1(net4541),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][7] ),
    .A2(net4633),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][7] ));
 sg13g2_a21oi_1 _16096_ (.A1(_06634_),
    .A2(_06635_),
    .Y(_06636_),
    .B1(net4477));
 sg13g2_a22oi_1 _16097_ (.Y(_06637_),
    .B1(net4542),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][7] ),
    .A2(net4588),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][7] ));
 sg13g2_a22oi_1 _16098_ (.Y(_06638_),
    .B1(net4634),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][7] ),
    .A2(net4682),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][7] ));
 sg13g2_a21oi_1 _16099_ (.A1(_06637_),
    .A2(_06638_),
    .Y(_06639_),
    .B1(net4466));
 sg13g2_a22oi_1 _16100_ (.Y(_06640_),
    .B1(net4542),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][7] ),
    .A2(net4587),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][7] ));
 sg13g2_a22oi_1 _16101_ (.Y(_06641_),
    .B1(net4634),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][7] ),
    .A2(net4682),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][7] ));
 sg13g2_a21oi_1 _16102_ (.A1(_06640_),
    .A2(_06641_),
    .Y(_06642_),
    .B1(net4452));
 sg13g2_a22oi_1 _16103_ (.Y(_06643_),
    .B1(net4580),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][7] ),
    .A2(net4673),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][7] ));
 sg13g2_a22oi_1 _16104_ (.Y(_06644_),
    .B1(net4535),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][7] ),
    .A2(net4628),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][7] ));
 sg13g2_a21oi_2 _16105_ (.B1(net4472),
    .Y(_06645_),
    .A2(_06644_),
    .A1(_06643_));
 sg13g2_nor4_2 _16106_ (.A(_06636_),
    .B(_06639_),
    .C(_06642_),
    .Y(_06646_),
    .D(_06645_));
 sg13g2_nand4_1 _16107_ (.B(_06630_),
    .C(_06633_),
    .A(net4363),
    .Y(_06647_),
    .D(_06646_));
 sg13g2_o21ai_1 _16108_ (.B1(_06647_),
    .Y(_06648_),
    .A1(net3309),
    .A2(net4358));
 sg13g2_nor2_1 _16109_ (.A(net5371),
    .B(_06648_),
    .Y(_01105_));
 sg13g2_a22oi_1 _16110_ (.Y(_06649_),
    .B1(net4538),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][8] ),
    .A2(net4682),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][8] ));
 sg13g2_a22oi_1 _16111_ (.Y(_06650_),
    .B1(net4585),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][8] ),
    .A2(net4632),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][8] ));
 sg13g2_a21oi_1 _16112_ (.A1(_06649_),
    .A2(_06650_),
    .Y(_06651_),
    .B1(net4459));
 sg13g2_a22oi_1 _16113_ (.Y(_06652_),
    .B1(net4574),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][8] ),
    .A2(net4668),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][8] ));
 sg13g2_a22oi_1 _16114_ (.Y(_06653_),
    .B1(net4529),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][8] ),
    .A2(net4622),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][8] ));
 sg13g2_a21oi_2 _16115_ (.B1(net4471),
    .Y(_06654_),
    .A2(_06653_),
    .A1(_06652_));
 sg13g2_a22oi_1 _16116_ (.Y(_06655_),
    .B1(net4574),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][8] ),
    .A2(net4670),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][8] ));
 sg13g2_a22oi_1 _16117_ (.Y(_06656_),
    .B1(net4529),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][8] ),
    .A2(net4622),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][8] ));
 sg13g2_a21oi_1 _16118_ (.A1(_06655_),
    .A2(_06656_),
    .Y(_06657_),
    .B1(net4490));
 sg13g2_a22oi_1 _16119_ (.Y(_06658_),
    .B1(net4545),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][8] ),
    .A2(net4637),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][8] ));
 sg13g2_a22oi_1 _16120_ (.Y(_06659_),
    .B1(net4590),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][8] ),
    .A2(net4686),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][8] ));
 sg13g2_a21oi_1 _16121_ (.A1(_06658_),
    .A2(_06659_),
    .Y(_06660_),
    .B1(net4503));
 sg13g2_a22oi_1 _16122_ (.Y(_06661_),
    .B1(net4545),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][8] ),
    .A2(net4589),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][8] ));
 sg13g2_a22oi_1 _16123_ (.Y(_06662_),
    .B1(net4636),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][8] ),
    .A2(net4684),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][8] ));
 sg13g2_a21oi_1 _16124_ (.A1(_06661_),
    .A2(_06662_),
    .Y(_06663_),
    .B1(net4451));
 sg13g2_a22oi_1 _16125_ (.Y(_06664_),
    .B1(net4576),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][8] ),
    .A2(net4669),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][8] ));
 sg13g2_a22oi_1 _16126_ (.Y(_06665_),
    .B1(net4532),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][8] ),
    .A2(net4623),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][8] ));
 sg13g2_a21oi_2 _16127_ (.B1(net4483),
    .Y(_06666_),
    .A2(_06665_),
    .A1(_06664_));
 sg13g2_a22oi_1 _16128_ (.Y(_06667_),
    .B1(net4579),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][8] ),
    .A2(net4672),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][8] ));
 sg13g2_a22oi_1 _16129_ (.Y(_06668_),
    .B1(net4534),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][8] ),
    .A2(net4627),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][8] ));
 sg13g2_a21oi_2 _16130_ (.B1(net4478),
    .Y(_06669_),
    .A2(_06668_),
    .A1(_06667_));
 sg13g2_a22oi_1 _16131_ (.Y(_06670_),
    .B1(net4534),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][8] ),
    .A2(net4674),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][8] ));
 sg13g2_a22oi_1 _16132_ (.Y(_06671_),
    .B1(net4579),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][8] ),
    .A2(net4627),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][8] ));
 sg13g2_a21o_1 _16133_ (.A2(_06671_),
    .A1(_06670_),
    .B1(net4465),
    .X(_06672_));
 sg13g2_nor3_2 _16134_ (.A(_06651_),
    .B(_06660_),
    .C(_06663_),
    .Y(_06673_));
 sg13g2_nor4_2 _16135_ (.A(_06654_),
    .B(_06657_),
    .C(_06666_),
    .Y(_06674_),
    .D(_06669_));
 sg13g2_nand4_1 _16136_ (.B(_06672_),
    .C(_06673_),
    .A(net4363),
    .Y(_06675_),
    .D(_06674_));
 sg13g2_o21ai_1 _16137_ (.B1(_06675_),
    .Y(_06676_),
    .A1(net3242),
    .A2(net4359));
 sg13g2_nor2_1 _16138_ (.A(net5372),
    .B(_06676_),
    .Y(_01106_));
 sg13g2_a22oi_1 _16139_ (.Y(_06677_),
    .B1(net4578),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][9] ),
    .A2(net4673),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][9] ));
 sg13g2_a22oi_1 _16140_ (.Y(_06678_),
    .B1(net4534),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][9] ),
    .A2(net4627),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][9] ));
 sg13g2_a21oi_2 _16141_ (.B1(net4489),
    .Y(_06679_),
    .A2(_06678_),
    .A1(_06677_));
 sg13g2_a22oi_1 _16142_ (.Y(_06680_),
    .B1(net4544),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][9] ),
    .A2(net4635),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][9] ));
 sg13g2_a22oi_1 _16143_ (.Y(_06681_),
    .B1(net4585),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][9] ),
    .A2(net4682),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][9] ));
 sg13g2_a21oi_1 _16144_ (.A1(_06680_),
    .A2(_06681_),
    .Y(_06682_),
    .B1(net4505));
 sg13g2_a22oi_1 _16145_ (.Y(_06683_),
    .B1(net4584),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][9] ),
    .A2(net4681),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][9] ));
 sg13g2_a22oi_1 _16146_ (.Y(_06684_),
    .B1(net4540),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][9] ),
    .A2(net4635),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][9] ));
 sg13g2_a21oi_1 _16147_ (.A1(_06683_),
    .A2(_06684_),
    .Y(_06685_),
    .B1(net4459));
 sg13g2_nor3_1 _16148_ (.A(_06679_),
    .B(_06682_),
    .C(_06685_),
    .Y(_06686_));
 sg13g2_a22oi_1 _16149_ (.Y(_06687_),
    .B1(net4579),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][9] ),
    .A2(net4674),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][9] ));
 sg13g2_a22oi_1 _16150_ (.Y(_06688_),
    .B1(net4539),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][9] ),
    .A2(net4631),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][9] ));
 sg13g2_a21o_1 _16151_ (.A2(_06688_),
    .A1(_06687_),
    .B1(net4465),
    .X(_06689_));
 sg13g2_a22oi_1 _16152_ (.Y(_06690_),
    .B1(net4530),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][9] ),
    .A2(net4575),
    .A1(\m_sys.m_ram.m_ram.r_mem[2][9] ));
 sg13g2_a22oi_1 _16153_ (.Y(_06691_),
    .B1(net4621),
    .B2(\m_sys.m_ram.m_ram.r_mem[0][9] ),
    .A2(net4667),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][9] ));
 sg13g2_a21oi_2 _16154_ (.B1(net4484),
    .Y(_06692_),
    .A2(_06691_),
    .A1(_06690_));
 sg13g2_a22oi_1 _16155_ (.Y(_06693_),
    .B1(net4533),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][9] ),
    .A2(net4671),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][9] ));
 sg13g2_a22oi_1 _16156_ (.Y(_06694_),
    .B1(net4578),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][9] ),
    .A2(net4626),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][9] ));
 sg13g2_a21oi_1 _16157_ (.A1(_06693_),
    .A2(_06694_),
    .Y(_06695_),
    .B1(net4471));
 sg13g2_a22oi_1 _16158_ (.Y(_06696_),
    .B1(net4584),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][9] ),
    .A2(net4679),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][9] ));
 sg13g2_a22oi_1 _16159_ (.Y(_06697_),
    .B1(net4539),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][9] ),
    .A2(net4627),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][9] ));
 sg13g2_a21oi_1 _16160_ (.A1(_06696_),
    .A2(_06697_),
    .Y(_06698_),
    .B1(net4477));
 sg13g2_a22oi_1 _16161_ (.Y(_06699_),
    .B1(net4538),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][9] ),
    .A2(net4680),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][9] ));
 sg13g2_a22oi_1 _16162_ (.Y(_06700_),
    .B1(net4583),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][9] ),
    .A2(net4632),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][9] ));
 sg13g2_a21oi_2 _16163_ (.B1(net4452),
    .Y(_06701_),
    .A2(_06700_),
    .A1(_06699_));
 sg13g2_nor4_2 _16164_ (.A(_06692_),
    .B(_06695_),
    .C(_06698_),
    .Y(_06702_),
    .D(_06701_));
 sg13g2_nand4_1 _16165_ (.B(_06686_),
    .C(_06689_),
    .A(net4363),
    .Y(_06703_),
    .D(_06702_));
 sg13g2_o21ai_1 _16166_ (.B1(_06703_),
    .Y(_06704_),
    .A1(net3305),
    .A2(net4360));
 sg13g2_nor2_1 _16167_ (.A(net5372),
    .B(_06704_),
    .Y(_01107_));
 sg13g2_a22oi_1 _16168_ (.Y(_06705_),
    .B1(net4584),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][10] ),
    .A2(net4679),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][10] ));
 sg13g2_a22oi_1 _16169_ (.Y(_06706_),
    .B1(net4539),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][10] ),
    .A2(net4631),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][10] ));
 sg13g2_a21oi_2 _16170_ (.B1(net4477),
    .Y(_06707_),
    .A2(_06706_),
    .A1(_06705_));
 sg13g2_a22oi_1 _16171_ (.Y(_06708_),
    .B1(net4637),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][10] ),
    .A2(net4687),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][10] ));
 sg13g2_a22oi_1 _16172_ (.Y(_06709_),
    .B1(net4544),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][10] ),
    .A2(net4589),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][10] ));
 sg13g2_a21oi_1 _16173_ (.A1(_06708_),
    .A2(_06709_),
    .Y(_06710_),
    .B1(net4451));
 sg13g2_a22oi_1 _16174_ (.Y(_06711_),
    .B1(net4545),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][10] ),
    .A2(net4590),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][10] ));
 sg13g2_a22oi_1 _16175_ (.Y(_06712_),
    .B1(net4637),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][10] ),
    .A2(net4684),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][10] ));
 sg13g2_a21oi_1 _16176_ (.A1(_06711_),
    .A2(_06712_),
    .Y(_06713_),
    .B1(net4503));
 sg13g2_nor3_2 _16177_ (.A(_06707_),
    .B(_06710_),
    .C(_06713_),
    .Y(_06714_));
 sg13g2_a22oi_1 _16178_ (.Y(_06715_),
    .B1(net4531),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][10] ),
    .A2(net4576),
    .A1(\m_sys.m_ram.m_ram.r_mem[2][10] ));
 sg13g2_a22oi_1 _16179_ (.Y(_06716_),
    .B1(net4621),
    .B2(\m_sys.m_ram.m_ram.r_mem[0][10] ),
    .A2(net4669),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][10] ));
 sg13g2_a21o_1 _16180_ (.A2(_06716_),
    .A1(_06715_),
    .B1(net4484),
    .X(_06717_));
 sg13g2_a22oi_1 _16181_ (.Y(_06718_),
    .B1(net4577),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][10] ),
    .A2(net4669),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][10] ));
 sg13g2_a22oi_1 _16182_ (.Y(_06719_),
    .B1(net4532),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][10] ),
    .A2(net4624),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][10] ));
 sg13g2_a21oi_1 _16183_ (.A1(_06718_),
    .A2(_06719_),
    .Y(_06720_),
    .B1(net4490));
 sg13g2_a22oi_1 _16184_ (.Y(_06721_),
    .B1(net4533),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][10] ),
    .A2(net4578),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][10] ));
 sg13g2_a22oi_1 _16185_ (.Y(_06722_),
    .B1(net4626),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][10] ),
    .A2(net4673),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][10] ));
 sg13g2_a21oi_1 _16186_ (.A1(_06721_),
    .A2(_06722_),
    .Y(_06723_),
    .B1(net4467));
 sg13g2_a22oi_1 _16187_ (.Y(_06724_),
    .B1(net4540),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][10] ),
    .A2(net4583),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][10] ));
 sg13g2_a22oi_1 _16188_ (.Y(_06725_),
    .B1(net4631),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][10] ),
    .A2(net4681),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][10] ));
 sg13g2_a21oi_2 _16189_ (.B1(net4459),
    .Y(_06726_),
    .A2(_06725_),
    .A1(_06724_));
 sg13g2_a22oi_1 _16190_ (.Y(_06727_),
    .B1(net4574),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][10] ),
    .A2(net4667),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][10] ));
 sg13g2_a22oi_1 _16191_ (.Y(_06728_),
    .B1(net4529),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][10] ),
    .A2(net4622),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][10] ));
 sg13g2_a21oi_2 _16192_ (.B1(net4471),
    .Y(_06729_),
    .A2(_06728_),
    .A1(_06727_));
 sg13g2_nor4_1 _16193_ (.A(_06720_),
    .B(_06723_),
    .C(_06726_),
    .D(_06729_),
    .Y(_06730_));
 sg13g2_nand4_1 _16194_ (.B(_06714_),
    .C(_06717_),
    .A(net4365),
    .Y(_06731_),
    .D(_06730_));
 sg13g2_o21ai_1 _16195_ (.B1(_06731_),
    .Y(_06732_),
    .A1(net3271),
    .A2(net4359));
 sg13g2_nor2_1 _16196_ (.A(net5372),
    .B(_06732_),
    .Y(_01108_));
 sg13g2_a22oi_1 _16197_ (.Y(_06733_),
    .B1(net4584),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][11] ),
    .A2(net4681),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][11] ));
 sg13g2_a22oi_1 _16198_ (.Y(_06734_),
    .B1(net4539),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][11] ),
    .A2(net4632),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][11] ));
 sg13g2_a21oi_1 _16199_ (.A1(_06733_),
    .A2(_06734_),
    .Y(_06735_),
    .B1(net4465));
 sg13g2_a22oi_1 _16200_ (.Y(_06736_),
    .B1(net4631),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][11] ),
    .A2(net4679),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][11] ));
 sg13g2_a22oi_1 _16201_ (.Y(_06737_),
    .B1(net4540),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][11] ),
    .A2(net4583),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][11] ));
 sg13g2_a21oi_2 _16202_ (.B1(net4459),
    .Y(_06738_),
    .A2(_06737_),
    .A1(_06736_));
 sg13g2_a22oi_1 _16203_ (.Y(_06739_),
    .B1(net4589),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][11] ),
    .A2(net4684),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][11] ));
 sg13g2_a22oi_1 _16204_ (.Y(_06740_),
    .B1(net4544),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][11] ),
    .A2(net4636),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][11] ));
 sg13g2_a21oi_2 _16205_ (.B1(net4452),
    .Y(_06741_),
    .A2(_06740_),
    .A1(_06739_));
 sg13g2_a22oi_1 _16206_ (.Y(_06742_),
    .B1(net4584),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][11] ),
    .A2(net4679),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][11] ));
 sg13g2_a22oi_1 _16207_ (.Y(_06743_),
    .B1(net4539),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][11] ),
    .A2(net4631),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][11] ));
 sg13g2_a21oi_1 _16208_ (.A1(_06742_),
    .A2(_06743_),
    .Y(_06744_),
    .B1(net4477));
 sg13g2_a22oi_1 _16209_ (.Y(_06745_),
    .B1(net4622),
    .B2(\m_sys.m_ram.m_ram.r_mem[12][11] ),
    .A2(net4667),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][11] ));
 sg13g2_a22oi_1 _16210_ (.Y(_06746_),
    .B1(net4529),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][11] ),
    .A2(net4575),
    .A1(\m_sys.m_ram.m_ram.r_mem[14][11] ));
 sg13g2_a21oi_1 _16211_ (.A1(_06745_),
    .A2(_06746_),
    .Y(_06747_),
    .B1(net4490));
 sg13g2_a22oi_1 _16212_ (.Y(_06748_),
    .B1(net4621),
    .B2(\m_sys.m_ram.m_ram.r_mem[0][11] ),
    .A2(net4669),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][11] ));
 sg13g2_a22oi_1 _16213_ (.Y(_06749_),
    .B1(net4530),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][11] ),
    .A2(net4575),
    .A1(\m_sys.m_ram.m_ram.r_mem[2][11] ));
 sg13g2_a21oi_1 _16214_ (.A1(_06748_),
    .A2(_06749_),
    .Y(_06750_),
    .B1(net4484));
 sg13g2_a22oi_1 _16215_ (.Y(_06751_),
    .B1(net4544),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][11] ),
    .A2(net4589),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][11] ));
 sg13g2_a22oi_1 _16216_ (.Y(_06752_),
    .B1(net4636),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][11] ),
    .A2(net4684),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][11] ));
 sg13g2_a21oi_2 _16217_ (.B1(net4503),
    .Y(_06753_),
    .A2(_06752_),
    .A1(_06751_));
 sg13g2_a22oi_1 _16218_ (.Y(_06754_),
    .B1(net4574),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][11] ),
    .A2(net4668),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][11] ));
 sg13g2_a22oi_1 _16219_ (.Y(_06755_),
    .B1(net4529),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][11] ),
    .A2(net4622),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][11] ));
 sg13g2_a21o_1 _16220_ (.A2(_06755_),
    .A1(_06754_),
    .B1(net4471),
    .X(_06756_));
 sg13g2_nor3_2 _16221_ (.A(_06735_),
    .B(_06744_),
    .C(_06753_),
    .Y(_06757_));
 sg13g2_nor4_1 _16222_ (.A(_06738_),
    .B(_06741_),
    .C(_06747_),
    .D(_06750_),
    .Y(_06758_));
 sg13g2_nand4_1 _16223_ (.B(_06756_),
    .C(_06757_),
    .A(net4365),
    .Y(_06759_),
    .D(_06758_));
 sg13g2_o21ai_1 _16224_ (.B1(_06759_),
    .Y(_06760_),
    .A1(net3238),
    .A2(net4360));
 sg13g2_nor2_1 _16225_ (.A(net5373),
    .B(_06760_),
    .Y(_01109_));
 sg13g2_a22oi_1 _16226_ (.Y(_06761_),
    .B1(net4574),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][12] ),
    .A2(net4668),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][12] ));
 sg13g2_a22oi_1 _16227_ (.Y(_06762_),
    .B1(net4529),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][12] ),
    .A2(net4622),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][12] ));
 sg13g2_a21oi_1 _16228_ (.A1(_06761_),
    .A2(_06762_),
    .Y(_06763_),
    .B1(net4471));
 sg13g2_a22oi_1 _16229_ (.Y(_06764_),
    .B1(net4538),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][12] ),
    .A2(net4632),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][12] ));
 sg13g2_a22oi_1 _16230_ (.Y(_06765_),
    .B1(net4583),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][12] ),
    .A2(net4680),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][12] ));
 sg13g2_a21oi_2 _16231_ (.B1(net4459),
    .Y(_06766_),
    .A2(_06765_),
    .A1(_06764_));
 sg13g2_a22oi_1 _16232_ (.Y(_06767_),
    .B1(net4574),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][12] ),
    .A2(net4667),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][12] ));
 sg13g2_a22oi_1 _16233_ (.Y(_06768_),
    .B1(net4529),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][12] ),
    .A2(net4622),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][12] ));
 sg13g2_a21oi_1 _16234_ (.A1(_06767_),
    .A2(_06768_),
    .Y(_06769_),
    .B1(net4490));
 sg13g2_a22oi_1 _16235_ (.Y(_06770_),
    .B1(net4590),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][12] ),
    .A2(net4637),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][12] ));
 sg13g2_a22oi_1 _16236_ (.Y(_06771_),
    .B1(net4545),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][12] ),
    .A2(net4687),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][12] ));
 sg13g2_a21oi_1 _16237_ (.A1(_06770_),
    .A2(_06771_),
    .Y(_06772_),
    .B1(net4451));
 sg13g2_a22oi_1 _16238_ (.Y(_06773_),
    .B1(net4545),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][12] ),
    .A2(net4590),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][12] ));
 sg13g2_a22oi_1 _16239_ (.Y(_06774_),
    .B1(net4637),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][12] ),
    .A2(net4687),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][12] ));
 sg13g2_a21oi_1 _16240_ (.A1(_06773_),
    .A2(_06774_),
    .Y(_06775_),
    .B1(net4503));
 sg13g2_a22oi_1 _16241_ (.Y(_06776_),
    .B1(net4579),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][12] ),
    .A2(net4672),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][12] ));
 sg13g2_a22oi_1 _16242_ (.Y(_06777_),
    .B1(net4534),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][12] ),
    .A2(net4627),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][12] ));
 sg13g2_a21oi_2 _16243_ (.B1(net4477),
    .Y(_06778_),
    .A2(_06777_),
    .A1(_06776_));
 sg13g2_a22oi_1 _16244_ (.Y(_06779_),
    .B1(net4621),
    .B2(\m_sys.m_ram.m_ram.r_mem[0][12] ),
    .A2(net4667),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][12] ));
 sg13g2_a22oi_1 _16245_ (.Y(_06780_),
    .B1(net4530),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][12] ),
    .A2(net4575),
    .A1(\m_sys.m_ram.m_ram.r_mem[2][12] ));
 sg13g2_a21oi_2 _16246_ (.B1(net4484),
    .Y(_06781_),
    .A2(_06780_),
    .A1(_06779_));
 sg13g2_a22oi_1 _16247_ (.Y(_06782_),
    .B1(net4533),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][12] ),
    .A2(net4578),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][12] ));
 sg13g2_a22oi_1 _16248_ (.Y(_06783_),
    .B1(net4626),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][12] ),
    .A2(net4671),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][12] ));
 sg13g2_a21o_1 _16249_ (.A2(_06783_),
    .A1(_06782_),
    .B1(net4467),
    .X(_06784_));
 sg13g2_nor3_2 _16250_ (.A(_06766_),
    .B(_06772_),
    .C(_06775_),
    .Y(_06785_));
 sg13g2_nor4_2 _16251_ (.A(_06763_),
    .B(_06769_),
    .C(_06778_),
    .Y(_06786_),
    .D(_06781_));
 sg13g2_nand4_1 _16252_ (.B(_06784_),
    .C(_06785_),
    .A(net4363),
    .Y(_06787_),
    .D(_06786_));
 sg13g2_o21ai_1 _16253_ (.B1(_06787_),
    .Y(_06788_),
    .A1(net3191),
    .A2(net4365));
 sg13g2_nor2_1 _16254_ (.A(net5374),
    .B(_06788_),
    .Y(_01110_));
 sg13g2_a22oi_1 _16255_ (.Y(_06789_),
    .B1(net4533),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][13] ),
    .A2(net4578),
    .A1(\m_sys.m_ram.m_ram.r_mem[22][13] ));
 sg13g2_a22oi_1 _16256_ (.Y(_06790_),
    .B1(net4626),
    .B2(\m_sys.m_ram.m_ram.r_mem[20][13] ),
    .A2(net4671),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][13] ));
 sg13g2_a21oi_1 _16257_ (.A1(_06789_),
    .A2(_06790_),
    .Y(_06791_),
    .B1(net4472));
 sg13g2_a22oi_1 _16258_ (.Y(_06792_),
    .B1(net4626),
    .B2(\m_sys.m_ram.m_ram.r_mem[12][13] ),
    .A2(net4671),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][13] ));
 sg13g2_a22oi_1 _16259_ (.Y(_06793_),
    .B1(net4533),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][13] ),
    .A2(net4578),
    .A1(\m_sys.m_ram.m_ram.r_mem[14][13] ));
 sg13g2_a21oi_1 _16260_ (.A1(_06792_),
    .A2(_06793_),
    .Y(_06794_),
    .B1(net4489));
 sg13g2_a22oi_1 _16261_ (.Y(_06795_),
    .B1(net4584),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][13] ),
    .A2(net4679),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][13] ));
 sg13g2_a22oi_1 _16262_ (.Y(_06796_),
    .B1(net4539),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][13] ),
    .A2(net4631),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][13] ));
 sg13g2_a21oi_1 _16263_ (.A1(_06795_),
    .A2(_06796_),
    .Y(_06797_),
    .B1(net4477));
 sg13g2_a22oi_1 _16264_ (.Y(_06798_),
    .B1(net4621),
    .B2(\m_sys.m_ram.m_ram.r_mem[0][13] ),
    .A2(net4667),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][13] ));
 sg13g2_a22oi_1 _16265_ (.Y(_06799_),
    .B1(net4530),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][13] ),
    .A2(net4575),
    .A1(\m_sys.m_ram.m_ram.r_mem[2][13] ));
 sg13g2_a21oi_2 _16266_ (.B1(net4484),
    .Y(_06800_),
    .A2(_06799_),
    .A1(_06798_));
 sg13g2_a22oi_1 _16267_ (.Y(_06801_),
    .B1(net4583),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][13] ),
    .A2(net4680),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][13] ));
 sg13g2_a22oi_1 _16268_ (.Y(_06802_),
    .B1(net4538),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][13] ),
    .A2(net4632),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][13] ));
 sg13g2_a21oi_2 _16269_ (.B1(net4452),
    .Y(_06803_),
    .A2(_06802_),
    .A1(_06801_));
 sg13g2_a22oi_1 _16270_ (.Y(_06804_),
    .B1(net4538),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][13] ),
    .A2(net4585),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][13] ));
 sg13g2_a22oi_1 _16271_ (.Y(_06805_),
    .B1(net4632),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][13] ),
    .A2(net4680),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][13] ));
 sg13g2_a21o_1 _16272_ (.A2(_06805_),
    .A1(_06804_),
    .B1(net4505),
    .X(_06806_));
 sg13g2_a22oi_1 _16273_ (.Y(_06807_),
    .B1(net4538),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][13] ),
    .A2(net4583),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][13] ));
 sg13g2_a22oi_1 _16274_ (.Y(_06808_),
    .B1(net4631),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][13] ),
    .A2(net4679),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][13] ));
 sg13g2_a21oi_1 _16275_ (.A1(_06807_),
    .A2(_06808_),
    .Y(_06809_),
    .B1(net4459));
 sg13g2_a22oi_1 _16276_ (.Y(_06810_),
    .B1(net4579),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][13] ),
    .A2(net4671),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][13] ));
 sg13g2_a22oi_1 _16277_ (.Y(_06811_),
    .B1(net4534),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][13] ),
    .A2(net4627),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][13] ));
 sg13g2_a21oi_1 _16278_ (.A1(_06810_),
    .A2(_06811_),
    .Y(_06812_),
    .B1(net4465));
 sg13g2_nor3_1 _16279_ (.A(_06794_),
    .B(_06800_),
    .C(_06809_),
    .Y(_06813_));
 sg13g2_nor4_1 _16280_ (.A(_06791_),
    .B(_06797_),
    .C(_06803_),
    .D(_06812_),
    .Y(_06814_));
 sg13g2_nand4_1 _16281_ (.B(_06806_),
    .C(_06813_),
    .A(net4363),
    .Y(_06815_),
    .D(_06814_));
 sg13g2_o21ai_1 _16282_ (.B1(_06815_),
    .Y(_06816_),
    .A1(net3096),
    .A2(net4360));
 sg13g2_nor2_1 _16283_ (.A(net5373),
    .B(_06816_),
    .Y(_01111_));
 sg13g2_a22oi_1 _16284_ (.Y(_06817_),
    .B1(net4631),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][14] ),
    .A2(net4679),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][14] ));
 sg13g2_a22oi_1 _16285_ (.Y(_06818_),
    .B1(net4538),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][14] ),
    .A2(net4583),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][14] ));
 sg13g2_a21oi_2 _16286_ (.B1(net4459),
    .Y(_06819_),
    .A2(_06818_),
    .A1(_06817_));
 sg13g2_a22oi_1 _16287_ (.Y(_06820_),
    .B1(net4579),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][14] ),
    .A2(net4672),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][14] ));
 sg13g2_a22oi_1 _16288_ (.Y(_06821_),
    .B1(net4534),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][14] ),
    .A2(net4630),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][14] ));
 sg13g2_a21oi_1 _16289_ (.A1(_06820_),
    .A2(_06821_),
    .Y(_06822_),
    .B1(net4478));
 sg13g2_a22oi_1 _16290_ (.Y(_06823_),
    .B1(net4574),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][14] ),
    .A2(net4668),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][14] ));
 sg13g2_a22oi_1 _16291_ (.Y(_06824_),
    .B1(net4533),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][14] ),
    .A2(net4626),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][14] ));
 sg13g2_a21oi_1 _16292_ (.A1(_06823_),
    .A2(_06824_),
    .Y(_06825_),
    .B1(net4471));
 sg13g2_nor3_1 _16293_ (.A(_06819_),
    .B(_06822_),
    .C(_06825_),
    .Y(_06826_));
 sg13g2_a22oi_1 _16294_ (.Y(_06827_),
    .B1(net4580),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][14] ),
    .A2(net4673),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][14] ));
 sg13g2_a22oi_1 _16295_ (.Y(_06828_),
    .B1(net4535),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][14] ),
    .A2(net4628),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][14] ));
 sg13g2_a21o_1 _16296_ (.A2(_06828_),
    .A1(_06827_),
    .B1(net4489),
    .X(_06829_));
 sg13g2_a22oi_1 _16297_ (.Y(_06830_),
    .B1(net4575),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][14] ),
    .A2(net4667),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][14] ));
 sg13g2_a22oi_1 _16298_ (.Y(_06831_),
    .B1(net4530),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][14] ),
    .A2(net4621),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][14] ));
 sg13g2_a21oi_2 _16299_ (.B1(net4484),
    .Y(_06832_),
    .A2(_06831_),
    .A1(_06830_));
 sg13g2_a22oi_1 _16300_ (.Y(_06833_),
    .B1(net4539),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][14] ),
    .A2(net4679),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][14] ));
 sg13g2_a22oi_1 _16301_ (.Y(_06834_),
    .B1(net4584),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][14] ),
    .A2(net4632),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][14] ));
 sg13g2_a21oi_1 _16302_ (.A1(_06833_),
    .A2(_06834_),
    .Y(_06835_),
    .B1(net4465));
 sg13g2_a22oi_1 _16303_ (.Y(_06836_),
    .B1(net4544),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][14] ),
    .A2(net4589),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][14] ));
 sg13g2_a22oi_1 _16304_ (.Y(_06837_),
    .B1(net4636),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][14] ),
    .A2(net4684),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][14] ));
 sg13g2_a21oi_2 _16305_ (.B1(net4451),
    .Y(_06838_),
    .A2(_06837_),
    .A1(_06836_));
 sg13g2_a22oi_1 _16306_ (.Y(_06839_),
    .B1(net4636),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][14] ),
    .A2(net4684),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][14] ));
 sg13g2_a22oi_1 _16307_ (.Y(_06840_),
    .B1(net4544),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][14] ),
    .A2(net4589),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][14] ));
 sg13g2_a21oi_2 _16308_ (.B1(net4503),
    .Y(_06841_),
    .A2(_06840_),
    .A1(_06839_));
 sg13g2_nor4_2 _16309_ (.A(_06832_),
    .B(_06835_),
    .C(_06838_),
    .Y(_06842_),
    .D(_06841_));
 sg13g2_nand4_1 _16310_ (.B(_06826_),
    .C(_06829_),
    .A(net4363),
    .Y(_06843_),
    .D(_06842_));
 sg13g2_o21ai_1 _16311_ (.B1(_06843_),
    .Y(_06844_),
    .A1(net3158),
    .A2(net4365));
 sg13g2_nor2_1 _16312_ (.A(net5373),
    .B(_06844_),
    .Y(_01112_));
 sg13g2_a22oi_1 _16313_ (.Y(_06845_),
    .B1(net4589),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][15] ),
    .A2(net4684),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][15] ));
 sg13g2_a22oi_1 _16314_ (.Y(_06846_),
    .B1(net4544),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][15] ),
    .A2(net4636),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][15] ));
 sg13g2_a21oi_2 _16315_ (.B1(net4503),
    .Y(_06847_),
    .A2(_06846_),
    .A1(_06845_));
 sg13g2_a22oi_1 _16316_ (.Y(_06848_),
    .B1(net4621),
    .B2(\m_sys.m_ram.m_ram.r_mem[0][15] ),
    .A2(net4667),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][15] ));
 sg13g2_a22oi_1 _16317_ (.Y(_06849_),
    .B1(net4529),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][15] ),
    .A2(net4574),
    .A1(\m_sys.m_ram.m_ram.r_mem[2][15] ));
 sg13g2_a21oi_2 _16318_ (.B1(net4484),
    .Y(_06850_),
    .A2(_06849_),
    .A1(_06848_));
 sg13g2_a22oi_1 _16319_ (.Y(_06851_),
    .B1(net4578),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][15] ),
    .A2(net4671),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][15] ));
 sg13g2_a22oi_1 _16320_ (.Y(_06852_),
    .B1(net4533),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][15] ),
    .A2(net4626),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][15] ));
 sg13g2_a21oi_1 _16321_ (.A1(_06851_),
    .A2(_06852_),
    .Y(_06853_),
    .B1(net4489));
 sg13g2_a22oi_1 _16322_ (.Y(_06854_),
    .B1(net4578),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][15] ),
    .A2(net4671),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][15] ));
 sg13g2_a22oi_1 _16323_ (.Y(_06855_),
    .B1(net4533),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][15] ),
    .A2(net4626),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][15] ));
 sg13g2_a21oi_1 _16324_ (.A1(_06854_),
    .A2(_06855_),
    .Y(_06856_),
    .B1(net4471));
 sg13g2_a22oi_1 _16325_ (.Y(_06857_),
    .B1(net4534),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][15] ),
    .A2(net4671),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][15] ));
 sg13g2_a22oi_1 _16326_ (.Y(_06858_),
    .B1(net4579),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][15] ),
    .A2(net4627),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][15] ));
 sg13g2_a21oi_1 _16327_ (.A1(_06857_),
    .A2(_06858_),
    .Y(_06859_),
    .B1(net4465));
 sg13g2_a22oi_1 _16328_ (.Y(_06860_),
    .B1(net4589),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][15] ),
    .A2(net4684),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][15] ));
 sg13g2_a22oi_1 _16329_ (.Y(_06861_),
    .B1(net4544),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][15] ),
    .A2(net4636),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][15] ));
 sg13g2_a21oi_2 _16330_ (.B1(net4451),
    .Y(_06862_),
    .A2(_06861_),
    .A1(_06860_));
 sg13g2_a22oi_1 _16331_ (.Y(_06863_),
    .B1(net4583),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][15] ),
    .A2(net4680),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][15] ));
 sg13g2_a22oi_1 _16332_ (.Y(_06864_),
    .B1(net4538),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][15] ),
    .A2(net4635),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][15] ));
 sg13g2_a21oi_2 _16333_ (.B1(net4459),
    .Y(_06865_),
    .A2(_06864_),
    .A1(_06863_));
 sg13g2_a22oi_1 _16334_ (.Y(_06866_),
    .B1(net4539),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][15] ),
    .A2(net4584),
    .A1(\m_sys.m_ram.m_ram.r_mem[10][15] ));
 sg13g2_a22oi_1 _16335_ (.Y(_06867_),
    .B1(net4630),
    .B2(\m_sys.m_ram.m_ram.r_mem[8][15] ),
    .A2(net4672),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][15] ));
 sg13g2_a21o_1 _16336_ (.A2(_06867_),
    .A1(_06866_),
    .B1(net4477),
    .X(_06868_));
 sg13g2_nor3_1 _16337_ (.A(_06847_),
    .B(_06856_),
    .C(_06859_),
    .Y(_06869_));
 sg13g2_nor4_1 _16338_ (.A(_06850_),
    .B(_06853_),
    .C(_06862_),
    .D(_06865_),
    .Y(_06870_));
 sg13g2_nand4_1 _16339_ (.B(_06868_),
    .C(_06869_),
    .A(net4363),
    .Y(_06871_),
    .D(_06870_));
 sg13g2_o21ai_1 _16340_ (.B1(_06871_),
    .Y(_06872_),
    .A1(net3136),
    .A2(net4365));
 sg13g2_nor2_1 _16341_ (.A(net5373),
    .B(_06872_),
    .Y(_01113_));
 sg13g2_a22oi_1 _16342_ (.Y(_06873_),
    .B1(net4611),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][16] ),
    .A2(net4656),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][16] ));
 sg13g2_a22oi_1 _16343_ (.Y(_06874_),
    .B1(net4520),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][16] ),
    .A2(net4565),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][16] ));
 sg13g2_a21oi_1 _16344_ (.A1(_06873_),
    .A2(_06874_),
    .Y(_06875_),
    .B1(net4458));
 sg13g2_a22oi_1 _16345_ (.Y(_06876_),
    .B1(net4566),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][16] ),
    .A2(net4612),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][16] ));
 sg13g2_a22oi_1 _16346_ (.Y(_06877_),
    .B1(net4521),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][16] ),
    .A2(net4657),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][16] ));
 sg13g2_a21oi_1 _16347_ (.A1(_06876_),
    .A2(_06877_),
    .Y(_06878_),
    .B1(net4469));
 sg13g2_a22oi_1 _16348_ (.Y(_06879_),
    .B1(net4566),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][16] ),
    .A2(net4657),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][16] ));
 sg13g2_a22oi_1 _16349_ (.Y(_06880_),
    .B1(net4521),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][16] ),
    .A2(net4612),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][16] ));
 sg13g2_a21oi_1 _16350_ (.A1(_06879_),
    .A2(_06880_),
    .Y(_06881_),
    .B1(net4487));
 sg13g2_nor3_1 _16351_ (.A(_06875_),
    .B(_06878_),
    .C(_06881_),
    .Y(_06882_));
 sg13g2_a22oi_1 _16352_ (.Y(_06883_),
    .B1(net4572),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][16] ),
    .A2(net4664),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][16] ));
 sg13g2_a22oi_1 _16353_ (.Y(_06884_),
    .B1(net4527),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][16] ),
    .A2(net4618),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][16] ));
 sg13g2_a21o_1 _16354_ (.A2(_06884_),
    .A1(_06883_),
    .B1(net4485),
    .X(_06885_));
 sg13g2_a22oi_1 _16355_ (.Y(_06886_),
    .B1(net4524),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][16] ),
    .A2(net4569),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][16] ));
 sg13g2_a22oi_1 _16356_ (.Y(_06887_),
    .B1(net4616),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][16] ),
    .A2(net4660),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][16] ));
 sg13g2_a21oi_1 _16357_ (.A1(_06886_),
    .A2(_06887_),
    .Y(_06888_),
    .B1(net4450));
 sg13g2_a22oi_1 _16358_ (.Y(_06889_),
    .B1(net4568),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][16] ),
    .A2(net4659),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][16] ));
 sg13g2_a22oi_1 _16359_ (.Y(_06890_),
    .B1(net4523),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][16] ),
    .A2(net4614),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][16] ));
 sg13g2_a21oi_1 _16360_ (.A1(_06889_),
    .A2(_06890_),
    .Y(_06891_),
    .B1(net4501));
 sg13g2_a22oi_1 _16361_ (.Y(_06892_),
    .B1(net4563),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][16] ),
    .A2(net4655),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][16] ));
 sg13g2_a22oi_1 _16362_ (.Y(_06893_),
    .B1(net4519),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][16] ),
    .A2(net4609),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][16] ));
 sg13g2_a21oi_2 _16363_ (.B1(net4476),
    .Y(_06894_),
    .A2(_06893_),
    .A1(_06892_));
 sg13g2_a22oi_1 _16364_ (.Y(_06895_),
    .B1(net4524),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][16] ),
    .A2(net4569),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][16] ));
 sg13g2_a22oi_1 _16365_ (.Y(_06896_),
    .B1(net4616),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][16] ),
    .A2(net4662),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][16] ));
 sg13g2_a21oi_2 _16366_ (.B1(net4464),
    .Y(_06897_),
    .A2(_06896_),
    .A1(_06895_));
 sg13g2_nor4_2 _16367_ (.A(_06888_),
    .B(_06891_),
    .C(_06894_),
    .Y(_06898_),
    .D(_06897_));
 sg13g2_nand4_1 _16368_ (.B(_06882_),
    .C(_06885_),
    .A(net4362),
    .Y(_06899_),
    .D(_06898_));
 sg13g2_o21ai_1 _16369_ (.B1(_06899_),
    .Y(_06900_),
    .A1(net3336),
    .A2(net4360));
 sg13g2_nor2_1 _16370_ (.A(net5373),
    .B(_06900_),
    .Y(_01114_));
 sg13g2_a22oi_1 _16371_ (.Y(_06901_),
    .B1(net4572),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][17] ),
    .A2(net4664),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][17] ));
 sg13g2_a22oi_1 _16372_ (.Y(_06902_),
    .B1(net4527),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][17] ),
    .A2(net4618),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][17] ));
 sg13g2_a21oi_2 _16373_ (.B1(net4485),
    .Y(_06903_),
    .A2(_06902_),
    .A1(_06901_));
 sg13g2_a22oi_1 _16374_ (.Y(_06904_),
    .B1(net4563),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][17] ),
    .A2(net4655),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][17] ));
 sg13g2_a22oi_1 _16375_ (.Y(_06905_),
    .B1(net4519),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][17] ),
    .A2(net4609),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][17] ));
 sg13g2_a21oi_2 _16376_ (.B1(net4475),
    .Y(_06906_),
    .A2(_06905_),
    .A1(_06904_));
 sg13g2_a22oi_1 _16377_ (.Y(_06907_),
    .B1(net4568),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][17] ),
    .A2(net4654),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][17] ));
 sg13g2_a22oi_1 _16378_ (.Y(_06908_),
    .B1(net4523),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][17] ),
    .A2(net4614),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][17] ));
 sg13g2_a21oi_1 _16379_ (.A1(_06907_),
    .A2(_06908_),
    .Y(_06909_),
    .B1(net4501));
 sg13g2_nor3_2 _16380_ (.A(_06903_),
    .B(_06906_),
    .C(_06909_),
    .Y(_06910_));
 sg13g2_a22oi_1 _16381_ (.Y(_06911_),
    .B1(net4572),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][17] ),
    .A2(net4661),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][17] ));
 sg13g2_a22oi_1 _16382_ (.Y(_06912_),
    .B1(net4527),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][17] ),
    .A2(net4618),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][17] ));
 sg13g2_a21o_1 _16383_ (.A2(_06912_),
    .A1(_06911_),
    .B1(net4458),
    .X(_06913_));
 sg13g2_a22oi_1 _16384_ (.Y(_06914_),
    .B1(net4567),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][17] ),
    .A2(net4657),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][17] ));
 sg13g2_a22oi_1 _16385_ (.Y(_06915_),
    .B1(net4521),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][17] ),
    .A2(net4609),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][17] ));
 sg13g2_a21oi_2 _16386_ (.B1(net4469),
    .Y(_06916_),
    .A2(_06915_),
    .A1(_06914_));
 sg13g2_a22oi_1 _16387_ (.Y(_06917_),
    .B1(net4526),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][17] ),
    .A2(net4662),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][17] ));
 sg13g2_a22oi_1 _16388_ (.Y(_06918_),
    .B1(net4571),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][17] ),
    .A2(net4619),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][17] ));
 sg13g2_a21oi_1 _16389_ (.A1(_06917_),
    .A2(_06918_),
    .Y(_06919_),
    .B1(net4464));
 sg13g2_a22oi_1 _16390_ (.Y(_06920_),
    .B1(net4524),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][17] ),
    .A2(net4570),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][17] ));
 sg13g2_a22oi_1 _16391_ (.Y(_06921_),
    .B1(net4617),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][17] ),
    .A2(net4660),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][17] ));
 sg13g2_a21oi_2 _16392_ (.B1(net4450),
    .Y(_06922_),
    .A2(_06921_),
    .A1(_06920_));
 sg13g2_a22oi_1 _16393_ (.Y(_06923_),
    .B1(net4618),
    .B2(\m_sys.m_ram.m_ram.r_mem[12][17] ),
    .A2(net4661),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][17] ));
 sg13g2_a22oi_1 _16394_ (.Y(_06924_),
    .B1(net4527),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][17] ),
    .A2(net4572),
    .A1(\m_sys.m_ram.m_ram.r_mem[14][17] ));
 sg13g2_a21oi_1 _16395_ (.A1(_06923_),
    .A2(_06924_),
    .Y(_06925_),
    .B1(net4488));
 sg13g2_nor4_1 _16396_ (.A(_06916_),
    .B(_06919_),
    .C(_06922_),
    .D(_06925_),
    .Y(_06926_));
 sg13g2_nand4_1 _16397_ (.B(_06910_),
    .C(_06913_),
    .A(net4362),
    .Y(_06927_),
    .D(_06926_));
 sg13g2_o21ai_1 _16398_ (.B1(_06927_),
    .Y(_06928_),
    .A1(net3314),
    .A2(net4360));
 sg13g2_nor2_1 _16399_ (.A(net5373),
    .B(_06928_),
    .Y(_01115_));
 sg13g2_a22oi_1 _16400_ (.Y(_06929_),
    .B1(net4564),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][18] ),
    .A2(net4610),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][18] ));
 sg13g2_a22oi_1 _16401_ (.Y(_06930_),
    .B1(net4518),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][18] ),
    .A2(net4656),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][18] ));
 sg13g2_a21oi_1 _16402_ (.A1(_06929_),
    .A2(_06930_),
    .Y(_06931_),
    .B1(net4469));
 sg13g2_a22oi_1 _16403_ (.Y(_06932_),
    .B1(net4616),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][18] ),
    .A2(net4660),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][18] ));
 sg13g2_a22oi_1 _16404_ (.Y(_06933_),
    .B1(net4524),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][18] ),
    .A2(net4569),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][18] ));
 sg13g2_a21oi_1 _16405_ (.A1(_06932_),
    .A2(_06933_),
    .Y(_06934_),
    .B1(net4450));
 sg13g2_a22oi_1 _16406_ (.Y(_06935_),
    .B1(net4564),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][18] ),
    .A2(net4654),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][18] ));
 sg13g2_a22oi_1 _16407_ (.Y(_06936_),
    .B1(net4518),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][18] ),
    .A2(net4610),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][18] ));
 sg13g2_a21oi_2 _16408_ (.B1(net4475),
    .Y(_06937_),
    .A2(_06936_),
    .A1(_06935_));
 sg13g2_a22oi_1 _16409_ (.Y(_06938_),
    .B1(net4573),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][18] ),
    .A2(net4663),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][18] ));
 sg13g2_a22oi_1 _16410_ (.Y(_06939_),
    .B1(net4528),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][18] ),
    .A2(net4619),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][18] ));
 sg13g2_a21oi_2 _16411_ (.B1(net4482),
    .Y(_06940_),
    .A2(_06939_),
    .A1(_06938_));
 sg13g2_a22oi_1 _16412_ (.Y(_06941_),
    .B1(net4523),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][18] ),
    .A2(net4568),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][18] ));
 sg13g2_a22oi_1 _16413_ (.Y(_06942_),
    .B1(net4614),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][18] ),
    .A2(net4659),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][18] ));
 sg13g2_a21oi_1 _16414_ (.A1(_06941_),
    .A2(_06942_),
    .Y(_06943_),
    .B1(net4502));
 sg13g2_a22oi_1 _16415_ (.Y(_06944_),
    .B1(net4565),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][18] ),
    .A2(net4656),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][18] ));
 sg13g2_a22oi_1 _16416_ (.Y(_06945_),
    .B1(net4520),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][18] ),
    .A2(net4611),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][18] ));
 sg13g2_a21oi_1 _16417_ (.A1(_06944_),
    .A2(_06945_),
    .Y(_06946_),
    .B1(net4487));
 sg13g2_a22oi_1 _16418_ (.Y(_06947_),
    .B1(net4563),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][18] ),
    .A2(net4657),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][18] ));
 sg13g2_a22oi_1 _16419_ (.Y(_06948_),
    .B1(net4519),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][18] ),
    .A2(net4609),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][18] ));
 sg13g2_a21oi_1 _16420_ (.A1(_06947_),
    .A2(_06948_),
    .Y(_06949_),
    .B1(net4461));
 sg13g2_a22oi_1 _16421_ (.Y(_06950_),
    .B1(net4530),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][18] ),
    .A2(net4576),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][18] ));
 sg13g2_a22oi_1 _16422_ (.Y(_06951_),
    .B1(net4621),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][18] ),
    .A2(net4669),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][18] ));
 sg13g2_a21o_1 _16423_ (.A2(_06951_),
    .A1(_06950_),
    .B1(net4467),
    .X(_06952_));
 sg13g2_nor3_1 _16424_ (.A(_06934_),
    .B(_06940_),
    .C(_06943_),
    .Y(_06953_));
 sg13g2_nor4_2 _16425_ (.A(_06931_),
    .B(_06937_),
    .C(_06946_),
    .Y(_06954_),
    .D(_06949_));
 sg13g2_nand4_1 _16426_ (.B(_06952_),
    .C(_06953_),
    .A(net4362),
    .Y(_06955_),
    .D(_06954_));
 sg13g2_o21ai_1 _16427_ (.B1(_06955_),
    .Y(_06956_),
    .A1(net3220),
    .A2(net4361));
 sg13g2_nor2_1 _16428_ (.A(net5374),
    .B(_06956_),
    .Y(_01116_));
 sg13g2_a22oi_1 _16429_ (.Y(_06957_),
    .B1(net4570),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][19] ),
    .A2(net4661),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][19] ));
 sg13g2_a22oi_1 _16430_ (.Y(_06958_),
    .B1(net4523),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][19] ),
    .A2(net4615),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][19] ));
 sg13g2_a21oi_1 _16431_ (.A1(_06957_),
    .A2(_06958_),
    .Y(_06959_),
    .B1(net4458));
 sg13g2_a22oi_1 _16432_ (.Y(_06960_),
    .B1(net4563),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][19] ),
    .A2(net4609),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][19] ));
 sg13g2_a22oi_1 _16433_ (.Y(_06961_),
    .B1(net4519),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][19] ),
    .A2(net4657),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][19] ));
 sg13g2_a21oi_1 _16434_ (.A1(_06960_),
    .A2(_06961_),
    .Y(_06962_),
    .B1(net4469));
 sg13g2_a22oi_1 _16435_ (.Y(_06963_),
    .B1(net4569),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][19] ),
    .A2(net4660),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][19] ));
 sg13g2_a22oi_1 _16436_ (.Y(_06964_),
    .B1(net4525),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][19] ),
    .A2(net4616),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][19] ));
 sg13g2_a21oi_2 _16437_ (.B1(net4450),
    .Y(_06965_),
    .A2(_06964_),
    .A1(_06963_));
 sg13g2_nor3_2 _16438_ (.A(_06959_),
    .B(_06962_),
    .C(_06965_),
    .Y(_06966_));
 sg13g2_a22oi_1 _16439_ (.Y(_06967_),
    .B1(net4619),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][19] ),
    .A2(net4662),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][19] ));
 sg13g2_a22oi_1 _16440_ (.Y(_06968_),
    .B1(net4526),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][19] ),
    .A2(net4571),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][19] ));
 sg13g2_a21o_1 _16441_ (.A2(_06968_),
    .A1(_06967_),
    .B1(net4464),
    .X(_06969_));
 sg13g2_a22oi_1 _16442_ (.Y(_06970_),
    .B1(net4563),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][19] ),
    .A2(net4654),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][19] ));
 sg13g2_a22oi_1 _16443_ (.Y(_06971_),
    .B1(net4523),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][19] ),
    .A2(net4614),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][19] ));
 sg13g2_a21oi_2 _16444_ (.B1(net4501),
    .Y(_06972_),
    .A2(_06971_),
    .A1(_06970_));
 sg13g2_a22oi_1 _16445_ (.Y(_06973_),
    .B1(net4521),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][19] ),
    .A2(net4663),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][19] ));
 sg13g2_a22oi_1 _16446_ (.Y(_06974_),
    .B1(net4566),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][19] ),
    .A2(net4612),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][19] ));
 sg13g2_a21oi_1 _16447_ (.A1(_06973_),
    .A2(_06974_),
    .Y(_06975_),
    .B1(net4485));
 sg13g2_a22oi_1 _16448_ (.Y(_06976_),
    .B1(net4521),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][19] ),
    .A2(net4566),
    .A1(\m_sys.m_ram.m_ram.r_mem[14][19] ));
 sg13g2_a22oi_1 _16449_ (.Y(_06977_),
    .B1(net4612),
    .B2(\m_sys.m_ram.m_ram.r_mem[12][19] ),
    .A2(net4657),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][19] ));
 sg13g2_a21oi_1 _16450_ (.A1(_06976_),
    .A2(_06977_),
    .Y(_06978_),
    .B1(net4487));
 sg13g2_a22oi_1 _16451_ (.Y(_06979_),
    .B1(net4563),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][19] ),
    .A2(net4655),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][19] ));
 sg13g2_a22oi_1 _16452_ (.Y(_06980_),
    .B1(net4519),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][19] ),
    .A2(net4609),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][19] ));
 sg13g2_a21oi_2 _16453_ (.B1(net4475),
    .Y(_06981_),
    .A2(_06980_),
    .A1(_06979_));
 sg13g2_nor4_1 _16454_ (.A(_06972_),
    .B(_06975_),
    .C(_06978_),
    .D(_06981_),
    .Y(_06982_));
 sg13g2_nand4_1 _16455_ (.B(_06966_),
    .C(_06969_),
    .A(net4362),
    .Y(_06983_),
    .D(_06982_));
 sg13g2_o21ai_1 _16456_ (.B1(_06983_),
    .Y(_06984_),
    .A1(net3311),
    .A2(net4360));
 sg13g2_nor2_1 _16457_ (.A(net5373),
    .B(_06984_),
    .Y(_01117_));
 sg13g2_a22oi_1 _16458_ (.Y(_06985_),
    .B1(net4564),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][20] ),
    .A2(net4610),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][20] ));
 sg13g2_a22oi_1 _16459_ (.Y(_06986_),
    .B1(net4518),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][20] ),
    .A2(net4656),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][20] ));
 sg13g2_a21oi_2 _16460_ (.B1(net4470),
    .Y(_06987_),
    .A2(_06986_),
    .A1(_06985_));
 sg13g2_a22oi_1 _16461_ (.Y(_06988_),
    .B1(net4616),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][20] ),
    .A2(net4660),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][20] ));
 sg13g2_a22oi_1 _16462_ (.Y(_06989_),
    .B1(net4524),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][20] ),
    .A2(net4569),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][20] ));
 sg13g2_a21oi_1 _16463_ (.A1(_06988_),
    .A2(_06989_),
    .Y(_06990_),
    .B1(net4450));
 sg13g2_a22oi_1 _16464_ (.Y(_06991_),
    .B1(net4565),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][20] ),
    .A2(net4656),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][20] ));
 sg13g2_a22oi_1 _16465_ (.Y(_06992_),
    .B1(net4520),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][20] ),
    .A2(net4611),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][20] ));
 sg13g2_a21oi_1 _16466_ (.A1(_06991_),
    .A2(_06992_),
    .Y(_06993_),
    .B1(net4487));
 sg13g2_a22oi_1 _16467_ (.Y(_06994_),
    .B1(net4523),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][20] ),
    .A2(net4614),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][20] ));
 sg13g2_a22oi_1 _16468_ (.Y(_06995_),
    .B1(net4568),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][20] ),
    .A2(net4659),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][20] ));
 sg13g2_a21oi_1 _16469_ (.A1(_06994_),
    .A2(_06995_),
    .Y(_06996_),
    .B1(net4501));
 sg13g2_a22oi_1 _16470_ (.Y(_06997_),
    .B1(net4525),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][20] ),
    .A2(net4568),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][20] ));
 sg13g2_a22oi_1 _16471_ (.Y(_06998_),
    .B1(net4615),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][20] ),
    .A2(net4659),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][20] ));
 sg13g2_a21oi_1 _16472_ (.A1(_06997_),
    .A2(_06998_),
    .Y(_06999_),
    .B1(net4458));
 sg13g2_a22oi_1 _16473_ (.Y(_07000_),
    .B1(net4564),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][20] ),
    .A2(net4654),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][20] ));
 sg13g2_a22oi_1 _16474_ (.Y(_07001_),
    .B1(net4518),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][20] ),
    .A2(net4610),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][20] ));
 sg13g2_a21oi_2 _16475_ (.B1(net4475),
    .Y(_07002_),
    .A2(_07001_),
    .A1(_07000_));
 sg13g2_a22oi_1 _16476_ (.Y(_07003_),
    .B1(net4565),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][20] ),
    .A2(net4663),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][20] ));
 sg13g2_a22oi_1 _16477_ (.Y(_07004_),
    .B1(net4520),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][20] ),
    .A2(net4611),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][20] ));
 sg13g2_a21oi_1 _16478_ (.A1(_07003_),
    .A2(_07004_),
    .Y(_07005_),
    .B1(net4481));
 sg13g2_a22oi_1 _16479_ (.Y(_07006_),
    .B1(net4526),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][20] ),
    .A2(net4571),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][20] ));
 sg13g2_a22oi_1 _16480_ (.Y(_07007_),
    .B1(net4623),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][20] ),
    .A2(net4669),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][20] ));
 sg13g2_a21o_1 _16481_ (.A2(_07007_),
    .A1(_07006_),
    .B1(net4467),
    .X(_07008_));
 sg13g2_nor3_2 _16482_ (.A(_06990_),
    .B(_06996_),
    .C(_06999_),
    .Y(_07009_));
 sg13g2_nor4_2 _16483_ (.A(_06987_),
    .B(_06993_),
    .C(_07002_),
    .Y(_07010_),
    .D(_07005_));
 sg13g2_nand4_1 _16484_ (.B(_07008_),
    .C(_07009_),
    .A(net4362),
    .Y(_07011_),
    .D(_07010_));
 sg13g2_o21ai_1 _16485_ (.B1(_07011_),
    .Y(_07012_),
    .A1(net3155),
    .A2(net4360));
 sg13g2_nor2_1 _16486_ (.A(net5374),
    .B(_07012_),
    .Y(_01118_));
 sg13g2_a22oi_1 _16487_ (.Y(_07013_),
    .B1(net4616),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][21] ),
    .A2(net4660),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][21] ));
 sg13g2_a22oi_1 _16488_ (.Y(_07014_),
    .B1(net4524),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][21] ),
    .A2(net4569),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][21] ));
 sg13g2_a21oi_2 _16489_ (.B1(net4453),
    .Y(_07015_),
    .A2(_07014_),
    .A1(_07013_));
 sg13g2_a22oi_1 _16490_ (.Y(_07016_),
    .B1(net4568),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][21] ),
    .A2(net4614),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][21] ));
 sg13g2_a22oi_1 _16491_ (.Y(_07017_),
    .B1(net4523),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][21] ),
    .A2(net4659),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][21] ));
 sg13g2_a21oi_1 _16492_ (.A1(_07016_),
    .A2(_07017_),
    .Y(_07018_),
    .B1(net4501));
 sg13g2_a22oi_1 _16493_ (.Y(_07019_),
    .B1(net4567),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][21] ),
    .A2(net4655),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][21] ));
 sg13g2_a22oi_1 _16494_ (.Y(_07020_),
    .B1(net4519),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][21] ),
    .A2(net4613),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][21] ));
 sg13g2_a21oi_1 _16495_ (.A1(_07019_),
    .A2(_07020_),
    .Y(_07021_),
    .B1(net4469));
 sg13g2_nor3_2 _16496_ (.A(_07015_),
    .B(_07018_),
    .C(_07021_),
    .Y(_07022_));
 sg13g2_a22oi_1 _16497_ (.Y(_07023_),
    .B1(net4572),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][21] ),
    .A2(net4664),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][21] ));
 sg13g2_a22oi_1 _16498_ (.Y(_07024_),
    .B1(net4527),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][21] ),
    .A2(net4618),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][21] ));
 sg13g2_a21o_1 _16499_ (.A2(_07024_),
    .A1(_07023_),
    .B1(net4485),
    .X(_07025_));
 sg13g2_a22oi_1 _16500_ (.Y(_07026_),
    .B1(net4563),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][21] ),
    .A2(net4654),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][21] ));
 sg13g2_a22oi_1 _16501_ (.Y(_07027_),
    .B1(net4519),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][21] ),
    .A2(net4609),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][21] ));
 sg13g2_a21oi_2 _16502_ (.B1(net4475),
    .Y(_07028_),
    .A2(_07027_),
    .A1(_07026_));
 sg13g2_a22oi_1 _16503_ (.Y(_07029_),
    .B1(net4527),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][21] ),
    .A2(net4572),
    .A1(\m_sys.m_ram.m_ram.r_mem[14][21] ));
 sg13g2_a22oi_1 _16504_ (.Y(_07030_),
    .B1(net4618),
    .B2(\m_sys.m_ram.m_ram.r_mem[12][21] ),
    .A2(net4661),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][21] ));
 sg13g2_a21oi_1 _16505_ (.A1(_07029_),
    .A2(_07030_),
    .Y(_07031_),
    .B1(net4488));
 sg13g2_a22oi_1 _16506_ (.Y(_07032_),
    .B1(net4527),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][21] ),
    .A2(net4572),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][21] ));
 sg13g2_a22oi_1 _16507_ (.Y(_07033_),
    .B1(net4615),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][21] ),
    .A2(net4661),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][21] ));
 sg13g2_a21oi_1 _16508_ (.A1(_07032_),
    .A2(_07033_),
    .Y(_07034_),
    .B1(net4458));
 sg13g2_a22oi_1 _16509_ (.Y(_07035_),
    .B1(net4571),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][21] ),
    .A2(net4661),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][21] ));
 sg13g2_a22oi_1 _16510_ (.Y(_07036_),
    .B1(net4526),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][21] ),
    .A2(net4619),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][21] ));
 sg13g2_a21oi_1 _16511_ (.A1(_07035_),
    .A2(_07036_),
    .Y(_07037_),
    .B1(net4464));
 sg13g2_nor4_1 _16512_ (.A(_07028_),
    .B(_07031_),
    .C(_07034_),
    .D(_07037_),
    .Y(_07038_));
 sg13g2_nand4_1 _16513_ (.B(_07022_),
    .C(_07025_),
    .A(net4362),
    .Y(_07039_),
    .D(_07038_));
 sg13g2_o21ai_1 _16514_ (.B1(_07039_),
    .Y(_07040_),
    .A1(net3190),
    .A2(net4360));
 sg13g2_nor2_1 _16515_ (.A(net5373),
    .B(_07040_),
    .Y(_01119_));
 sg13g2_a22oi_1 _16516_ (.Y(_07041_),
    .B1(net4565),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][22] ),
    .A2(net4663),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][22] ));
 sg13g2_a22oi_1 _16517_ (.Y(_07042_),
    .B1(net4520),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][22] ),
    .A2(net4611),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][22] ));
 sg13g2_a21oi_1 _16518_ (.A1(_07041_),
    .A2(_07042_),
    .Y(_07043_),
    .B1(net4485));
 sg13g2_a22oi_1 _16519_ (.Y(_07044_),
    .B1(net4565),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][22] ),
    .A2(net4656),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][22] ));
 sg13g2_a22oi_1 _16520_ (.Y(_07045_),
    .B1(net4520),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][22] ),
    .A2(net4611),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][22] ));
 sg13g2_a21oi_1 _16521_ (.A1(_07044_),
    .A2(_07045_),
    .Y(_07046_),
    .B1(net4487));
 sg13g2_a22oi_1 _16522_ (.Y(_07047_),
    .B1(net4564),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][22] ),
    .A2(net4654),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][22] ));
 sg13g2_a22oi_1 _16523_ (.Y(_07048_),
    .B1(net4518),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][22] ),
    .A2(net4610),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][22] ));
 sg13g2_a21oi_2 _16524_ (.B1(net4475),
    .Y(_07049_),
    .A2(_07048_),
    .A1(_07047_));
 sg13g2_nor3_1 _16525_ (.A(_07043_),
    .B(_07046_),
    .C(_07049_),
    .Y(_07050_));
 sg13g2_a22oi_1 _16526_ (.Y(_07051_),
    .B1(net4565),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][22] ),
    .A2(net4611),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][22] ));
 sg13g2_a22oi_1 _16527_ (.Y(_07052_),
    .B1(net4520),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][22] ),
    .A2(net4656),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][22] ));
 sg13g2_a21o_1 _16528_ (.A2(_07052_),
    .A1(_07051_),
    .B1(net4469),
    .X(_07053_));
 sg13g2_a22oi_1 _16529_ (.Y(_07054_),
    .B1(net4570),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][22] ),
    .A2(net4659),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][22] ));
 sg13g2_a22oi_1 _16530_ (.Y(_07055_),
    .B1(net4525),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][22] ),
    .A2(net4614),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][22] ));
 sg13g2_a21oi_2 _16531_ (.B1(net4501),
    .Y(_07056_),
    .A2(_07055_),
    .A1(_07054_));
 sg13g2_a22oi_1 _16532_ (.Y(_07057_),
    .B1(net4524),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][22] ),
    .A2(net4569),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][22] ));
 sg13g2_a22oi_1 _16533_ (.Y(_07058_),
    .B1(net4616),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][22] ),
    .A2(net4661),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][22] ));
 sg13g2_a21oi_1 _16534_ (.A1(_07057_),
    .A2(_07058_),
    .Y(_07059_),
    .B1(net4464));
 sg13g2_a22oi_1 _16535_ (.Y(_07060_),
    .B1(net4525),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][22] ),
    .A2(net4568),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][22] ));
 sg13g2_a22oi_1 _16536_ (.Y(_07061_),
    .B1(net4615),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][22] ),
    .A2(net4661),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][22] ));
 sg13g2_a21oi_1 _16537_ (.A1(_07060_),
    .A2(_07061_),
    .Y(_07062_),
    .B1(net4458));
 sg13g2_a22oi_1 _16538_ (.Y(_07063_),
    .B1(net4616),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][22] ),
    .A2(net4659),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][22] ));
 sg13g2_a22oi_1 _16539_ (.Y(_07064_),
    .B1(net4524),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][22] ),
    .A2(net4569),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][22] ));
 sg13g2_a21oi_2 _16540_ (.B1(net4450),
    .Y(_07065_),
    .A2(_07064_),
    .A1(_07063_));
 sg13g2_nor4_2 _16541_ (.A(_07056_),
    .B(_07059_),
    .C(_07062_),
    .Y(_07066_),
    .D(_07065_));
 sg13g2_nand4_1 _16542_ (.B(_07050_),
    .C(_07053_),
    .A(net4362),
    .Y(_07067_),
    .D(_07066_));
 sg13g2_o21ai_1 _16543_ (.B1(_07067_),
    .Y(_07068_),
    .A1(net3270),
    .A2(net4358));
 sg13g2_nor2_1 _16544_ (.A(net5371),
    .B(_07068_),
    .Y(_01120_));
 sg13g2_a22oi_1 _16545_ (.Y(_07069_),
    .B1(net4525),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][23] ),
    .A2(net4617),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][23] ));
 sg13g2_a22oi_1 _16546_ (.Y(_07070_),
    .B1(net4570),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][23] ),
    .A2(net4660),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][23] ));
 sg13g2_a21oi_1 _16547_ (.A1(_07069_),
    .A2(_07070_),
    .Y(_07071_),
    .B1(net4450));
 sg13g2_a22oi_1 _16548_ (.Y(_07072_),
    .B1(net4564),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][23] ),
    .A2(net4654),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][23] ));
 sg13g2_a22oi_1 _16549_ (.Y(_07073_),
    .B1(net4518),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][23] ),
    .A2(net4610),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][23] ));
 sg13g2_a21oi_2 _16550_ (.B1(net4475),
    .Y(_07074_),
    .A2(_07073_),
    .A1(_07072_));
 sg13g2_a22oi_1 _16551_ (.Y(_07075_),
    .B1(net4564),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][23] ),
    .A2(net4654),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][23] ));
 sg13g2_a22oi_1 _16552_ (.Y(_07076_),
    .B1(net4518),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][23] ),
    .A2(net4610),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][23] ));
 sg13g2_a21oi_1 _16553_ (.A1(_07075_),
    .A2(_07076_),
    .Y(_07077_),
    .B1(net4469));
 sg13g2_a22oi_1 _16554_ (.Y(_07078_),
    .B1(net4611),
    .B2(\m_sys.m_ram.m_ram.r_mem[12][23] ),
    .A2(net4656),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][23] ));
 sg13g2_a22oi_1 _16555_ (.Y(_07079_),
    .B1(net4520),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][23] ),
    .A2(net4565),
    .A1(\m_sys.m_ram.m_ram.r_mem[14][23] ));
 sg13g2_a21oi_1 _16556_ (.A1(_07078_),
    .A2(_07079_),
    .Y(_07080_),
    .B1(net4487));
 sg13g2_a22oi_1 _16557_ (.Y(_07081_),
    .B1(net4526),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][23] ),
    .A2(net4571),
    .A1(\m_sys.m_ram.m_ram.r_mem[2][23] ));
 sg13g2_a22oi_1 _16558_ (.Y(_07082_),
    .B1(net4619),
    .B2(\m_sys.m_ram.m_ram.r_mem[0][23] ),
    .A2(net4664),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][23] ));
 sg13g2_a21oi_2 _16559_ (.B1(net4482),
    .Y(_07083_),
    .A2(_07082_),
    .A1(_07081_));
 sg13g2_a22oi_1 _16560_ (.Y(_07084_),
    .B1(net4614),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][23] ),
    .A2(net4659),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][23] ));
 sg13g2_a22oi_1 _16561_ (.Y(_07085_),
    .B1(net4523),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][23] ),
    .A2(net4568),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][23] ));
 sg13g2_a21oi_2 _16562_ (.B1(net4501),
    .Y(_07086_),
    .A2(_07085_),
    .A1(_07084_));
 sg13g2_a22oi_1 _16563_ (.Y(_07087_),
    .B1(net4563),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][23] ),
    .A2(net4657),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][23] ));
 sg13g2_a22oi_1 _16564_ (.Y(_07088_),
    .B1(net4518),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][23] ),
    .A2(net4609),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][23] ));
 sg13g2_a21oi_1 _16565_ (.A1(_07087_),
    .A2(_07088_),
    .Y(_07089_),
    .B1(net4461));
 sg13g2_a22oi_1 _16566_ (.Y(_07090_),
    .B1(net4531),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][23] ),
    .A2(net4576),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][23] ));
 sg13g2_a22oi_1 _16567_ (.Y(_07091_),
    .B1(net4623),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][23] ),
    .A2(net4669),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][23] ));
 sg13g2_a21o_1 _16568_ (.A2(_07091_),
    .A1(_07090_),
    .B1(net4467),
    .X(_07092_));
 sg13g2_nor3_1 _16569_ (.A(_07071_),
    .B(_07083_),
    .C(_07086_),
    .Y(_07093_));
 sg13g2_nor4_2 _16570_ (.A(_07074_),
    .B(_07077_),
    .C(_07080_),
    .Y(_07094_),
    .D(_07089_));
 sg13g2_nand4_1 _16571_ (.B(_07092_),
    .C(_07093_),
    .A(net4362),
    .Y(_07095_),
    .D(_07094_));
 sg13g2_o21ai_1 _16572_ (.B1(_07095_),
    .Y(_07096_),
    .A1(net3159),
    .A2(net4361));
 sg13g2_nor2_1 _16573_ (.A(net5374),
    .B(_07096_),
    .Y(_01121_));
 sg13g2_a22oi_1 _16574_ (.Y(_07097_),
    .B1(net4554),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][24] ),
    .A2(net4645),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][24] ));
 sg13g2_a22oi_1 _16575_ (.Y(_07098_),
    .B1(net4508),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][24] ),
    .A2(net4599),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][24] ));
 sg13g2_a21oi_1 _16576_ (.A1(_07097_),
    .A2(_07098_),
    .Y(_07099_),
    .B1(net4456));
 sg13g2_a22oi_1 _16577_ (.Y(_07100_),
    .B1(net4603),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][24] ),
    .A2(net4649),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][24] ));
 sg13g2_a22oi_1 _16578_ (.Y(_07101_),
    .B1(net4514),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][24] ),
    .A2(net4559),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][24] ));
 sg13g2_a21oi_2 _16579_ (.B1(net4499),
    .Y(_07102_),
    .A2(_07101_),
    .A1(_07100_));
 sg13g2_a22oi_1 _16580_ (.Y(_07103_),
    .B1(net4555),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][24] ),
    .A2(net4652),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][24] ));
 sg13g2_a22oi_1 _16581_ (.Y(_07104_),
    .B1(net4509),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][24] ),
    .A2(net4601),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][24] ));
 sg13g2_a21oi_2 _16582_ (.B1(net4486),
    .Y(_07105_),
    .A2(_07104_),
    .A1(_07103_));
 sg13g2_a22oi_1 _16583_ (.Y(_07106_),
    .B1(net4509),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][24] ),
    .A2(net4555),
    .A1(\m_sys.m_ram.m_ram.r_mem[2][24] ));
 sg13g2_a22oi_1 _16584_ (.Y(_07107_),
    .B1(net4600),
    .B2(\m_sys.m_ram.m_ram.r_mem[0][24] ),
    .A2(net4646),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][24] ));
 sg13g2_a21oi_2 _16585_ (.B1(net4480),
    .Y(_07108_),
    .A2(_07107_),
    .A1(_07106_));
 sg13g2_a22oi_1 _16586_ (.Y(_07109_),
    .B1(net4516),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][24] ),
    .A2(net4561),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][24] ));
 sg13g2_a22oi_1 _16587_ (.Y(_07110_),
    .B1(net4603),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][24] ),
    .A2(net4650),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][24] ));
 sg13g2_a21oi_1 _16588_ (.A1(_07109_),
    .A2(_07110_),
    .Y(_07111_),
    .B1(net4448));
 sg13g2_a22oi_1 _16589_ (.Y(_07112_),
    .B1(net4552),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][24] ),
    .A2(net4646),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][24] ));
 sg13g2_a22oi_1 _16590_ (.Y(_07113_),
    .B1(net4508),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][24] ),
    .A2(net4598),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][24] ));
 sg13g2_a21oi_1 _16591_ (.A1(_07112_),
    .A2(_07113_),
    .Y(_07114_),
    .B1(net4474));
 sg13g2_a22oi_1 _16592_ (.Y(_07115_),
    .B1(net4507),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][24] ),
    .A2(net4644),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][24] ));
 sg13g2_a22oi_1 _16593_ (.Y(_07116_),
    .B1(net4553),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][24] ),
    .A2(net4599),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][24] ));
 sg13g2_a21oi_2 _16594_ (.B1(net4468),
    .Y(_07117_),
    .A2(_07116_),
    .A1(_07115_));
 sg13g2_a22oi_1 _16595_ (.Y(_07118_),
    .B1(net4515),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][24] ),
    .A2(net4560),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][24] ));
 sg13g2_a22oi_1 _16596_ (.Y(_07119_),
    .B1(net4605),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][24] ),
    .A2(net4650),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][24] ));
 sg13g2_a21o_1 _16597_ (.A2(_07119_),
    .A1(_07118_),
    .B1(net4462),
    .X(_07120_));
 sg13g2_nor3_1 _16598_ (.A(_07102_),
    .B(_07108_),
    .C(_07111_),
    .Y(_07121_));
 sg13g2_nor4_2 _16599_ (.A(_07099_),
    .B(_07105_),
    .C(_07114_),
    .Y(_07122_),
    .D(_07117_));
 sg13g2_nand4_1 _16600_ (.B(_07120_),
    .C(_07121_),
    .A(net4357),
    .Y(_07123_),
    .D(_07122_));
 sg13g2_o21ai_1 _16601_ (.B1(_07123_),
    .Y(_07124_),
    .A1(net3404),
    .A2(net4355));
 sg13g2_nor2_1 _16602_ (.A(net5368),
    .B(_07124_),
    .Y(_01122_));
 sg13g2_a22oi_1 _16603_ (.Y(_07125_),
    .B1(net4514),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][25] ),
    .A2(net4604),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][25] ));
 sg13g2_a22oi_1 _16604_ (.Y(_07126_),
    .B1(net4558),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][25] ),
    .A2(net4649),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][25] ));
 sg13g2_a21oi_1 _16605_ (.A1(_07125_),
    .A2(_07126_),
    .Y(_07127_),
    .B1(net4457));
 sg13g2_a22oi_1 _16606_ (.Y(_07128_),
    .B1(net4556),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][25] ),
    .A2(net4652),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][25] ));
 sg13g2_a22oi_1 _16607_ (.Y(_07129_),
    .B1(net4510),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][25] ),
    .A2(net4601),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][25] ));
 sg13g2_a21oi_1 _16608_ (.A1(_07128_),
    .A2(_07129_),
    .Y(_07130_),
    .B1(net4486));
 sg13g2_a22oi_1 _16609_ (.Y(_07131_),
    .B1(net4552),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][25] ),
    .A2(net4644),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][25] ));
 sg13g2_a22oi_1 _16610_ (.Y(_07132_),
    .B1(net4507),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][25] ),
    .A2(net4598),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][25] ));
 sg13g2_a21oi_2 _16611_ (.B1(net4468),
    .Y(_07133_),
    .A2(_07132_),
    .A1(_07131_));
 sg13g2_a22oi_1 _16612_ (.Y(_07134_),
    .B1(net4559),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][25] ),
    .A2(net4651),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][25] ));
 sg13g2_a22oi_1 _16613_ (.Y(_07135_),
    .B1(net4514),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][25] ),
    .A2(net4607),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][25] ));
 sg13g2_a21oi_1 _16614_ (.A1(_07134_),
    .A2(_07135_),
    .Y(_07136_),
    .B1(net4499));
 sg13g2_a22oi_1 _16615_ (.Y(_07137_),
    .B1(net4514),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][25] ),
    .A2(net4558),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][25] ));
 sg13g2_a22oi_1 _16616_ (.Y(_07138_),
    .B1(net4604),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][25] ),
    .A2(net4649),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][25] ));
 sg13g2_a21oi_1 _16617_ (.A1(_07137_),
    .A2(_07138_),
    .Y(_07139_),
    .B1(net4449));
 sg13g2_a22oi_1 _16618_ (.Y(_07140_),
    .B1(net4552),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][25] ),
    .A2(net4646),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][25] ));
 sg13g2_a22oi_1 _16619_ (.Y(_07141_),
    .B1(net4508),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][25] ),
    .A2(net4598),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][25] ));
 sg13g2_a21oi_1 _16620_ (.A1(_07140_),
    .A2(_07141_),
    .Y(_07142_),
    .B1(net4474));
 sg13g2_a22oi_1 _16621_ (.Y(_07143_),
    .B1(net4555),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][25] ),
    .A2(net4600),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][25] ));
 sg13g2_a22oi_1 _16622_ (.Y(_07144_),
    .B1(net4509),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][25] ),
    .A2(net4646),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][25] ));
 sg13g2_a21oi_1 _16623_ (.A1(_07143_),
    .A2(_07144_),
    .Y(_07145_),
    .B1(net4480));
 sg13g2_a22oi_1 _16624_ (.Y(_07146_),
    .B1(net4516),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][25] ),
    .A2(net4653),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][25] ));
 sg13g2_a22oi_1 _16625_ (.Y(_07147_),
    .B1(net4561),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][25] ),
    .A2(net4606),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][25] ));
 sg13g2_a21o_1 _16626_ (.A2(_07147_),
    .A1(_07146_),
    .B1(net4462),
    .X(_07148_));
 sg13g2_nor3_2 _16627_ (.A(_07127_),
    .B(_07136_),
    .C(_07139_),
    .Y(_07149_));
 sg13g2_nor4_2 _16628_ (.A(_07130_),
    .B(_07133_),
    .C(_07142_),
    .Y(_07150_),
    .D(_07145_));
 sg13g2_nand4_1 _16629_ (.B(_07148_),
    .C(_07149_),
    .A(net4356),
    .Y(_07151_),
    .D(_07150_));
 sg13g2_o21ai_1 _16630_ (.B1(_07151_),
    .Y(_07152_),
    .A1(net3398),
    .A2(net4356));
 sg13g2_nor2_1 _16631_ (.A(net5367),
    .B(_07152_),
    .Y(_01123_));
 sg13g2_a22oi_1 _16632_ (.Y(_07153_),
    .B1(net4561),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][26] ),
    .A2(net4651),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][26] ));
 sg13g2_a22oi_1 _16633_ (.Y(_07154_),
    .B1(net4516),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][26] ),
    .A2(net4606),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][26] ));
 sg13g2_a21oi_1 _16634_ (.A1(_07153_),
    .A2(_07154_),
    .Y(_07155_),
    .B1(net4448));
 sg13g2_a22oi_1 _16635_ (.Y(_07156_),
    .B1(net4603),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][26] ),
    .A2(net4649),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][26] ));
 sg13g2_a22oi_1 _16636_ (.Y(_07157_),
    .B1(net4513),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][26] ),
    .A2(net4558),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][26] ));
 sg13g2_a21oi_2 _16637_ (.B1(net4499),
    .Y(_07158_),
    .A2(_07157_),
    .A1(_07156_));
 sg13g2_a22oi_1 _16638_ (.Y(_07159_),
    .B1(net4560),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][26] ),
    .A2(net4653),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][26] ));
 sg13g2_a22oi_1 _16639_ (.Y(_07160_),
    .B1(net4511),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][26] ),
    .A2(net4602),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][26] ));
 sg13g2_a21oi_1 _16640_ (.A1(_07159_),
    .A2(_07160_),
    .Y(_07161_),
    .B1(net4488));
 sg13g2_nor3_1 _16641_ (.A(_07155_),
    .B(_07158_),
    .C(_07161_),
    .Y(_07162_));
 sg13g2_a22oi_1 _16642_ (.Y(_07163_),
    .B1(net4556),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][26] ),
    .A2(net4646),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][26] ));
 sg13g2_a22oi_1 _16643_ (.Y(_07164_),
    .B1(net4511),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][26] ),
    .A2(net4602),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][26] ));
 sg13g2_a21o_1 _16644_ (.A2(_07164_),
    .A1(_07163_),
    .B1(net4474),
    .X(_07165_));
 sg13g2_a22oi_1 _16645_ (.Y(_07166_),
    .B1(net4508),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][26] ),
    .A2(net4553),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][26] ));
 sg13g2_a22oi_1 _16646_ (.Y(_07167_),
    .B1(net4599),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][26] ),
    .A2(net4647),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][26] ));
 sg13g2_a21oi_1 _16647_ (.A1(_07166_),
    .A2(_07167_),
    .Y(_07168_),
    .B1(net4456));
 sg13g2_a22oi_1 _16648_ (.Y(_07169_),
    .B1(net4557),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][26] ),
    .A2(net4647),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][26] ));
 sg13g2_a22oi_1 _16649_ (.Y(_07170_),
    .B1(net4511),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][26] ),
    .A2(net4602),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][26] ));
 sg13g2_a21oi_1 _16650_ (.A1(_07169_),
    .A2(_07170_),
    .Y(_07171_),
    .B1(net4480));
 sg13g2_a22oi_1 _16651_ (.Y(_07172_),
    .B1(net4553),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][26] ),
    .A2(net4599),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][26] ));
 sg13g2_a22oi_1 _16652_ (.Y(_07173_),
    .B1(net4512),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][26] ),
    .A2(net4645),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][26] ));
 sg13g2_a21oi_2 _16653_ (.B1(net4468),
    .Y(_07174_),
    .A2(_07173_),
    .A1(_07172_));
 sg13g2_a22oi_1 _16654_ (.Y(_07175_),
    .B1(net4515),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][26] ),
    .A2(net4560),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][26] ));
 sg13g2_a22oi_1 _16655_ (.Y(_07176_),
    .B1(net4605),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][26] ),
    .A2(net4650),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][26] ));
 sg13g2_a21oi_1 _16656_ (.A1(_07175_),
    .A2(_07176_),
    .Y(_07177_),
    .B1(net4462));
 sg13g2_nor4_1 _16657_ (.A(_07168_),
    .B(_07171_),
    .C(_07174_),
    .D(_07177_),
    .Y(_07178_));
 sg13g2_nand4_1 _16658_ (.B(_07162_),
    .C(_07165_),
    .A(net4357),
    .Y(_07179_),
    .D(_07178_));
 sg13g2_o21ai_1 _16659_ (.B1(_07179_),
    .Y(_07180_),
    .A1(net3431),
    .A2(net4356));
 sg13g2_nor2_1 _16660_ (.A(net5367),
    .B(_07180_),
    .Y(_01124_));
 sg13g2_a22oi_1 _16661_ (.Y(_07181_),
    .B1(net4556),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][27] ),
    .A2(net4647),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][27] ));
 sg13g2_a22oi_1 _16662_ (.Y(_07182_),
    .B1(net4511),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][27] ),
    .A2(net4602),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][27] ));
 sg13g2_a21oi_1 _16663_ (.A1(_07181_),
    .A2(_07182_),
    .Y(_07183_),
    .B1(net4480));
 sg13g2_a22oi_1 _16664_ (.Y(_07184_),
    .B1(net4553),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][27] ),
    .A2(net4645),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][27] ));
 sg13g2_a22oi_1 _16665_ (.Y(_07185_),
    .B1(net4508),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][27] ),
    .A2(net4608),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][27] ));
 sg13g2_a21oi_2 _16666_ (.B1(net4468),
    .Y(_07186_),
    .A2(_07185_),
    .A1(_07184_));
 sg13g2_a22oi_1 _16667_ (.Y(_07187_),
    .B1(net4516),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][27] ),
    .A2(net4561),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][27] ));
 sg13g2_a22oi_1 _16668_ (.Y(_07188_),
    .B1(net4605),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][27] ),
    .A2(net4650),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][27] ));
 sg13g2_a21oi_1 _16669_ (.A1(_07187_),
    .A2(_07188_),
    .Y(_07189_),
    .B1(net4448));
 sg13g2_nor3_1 _16670_ (.A(_07183_),
    .B(_07186_),
    .C(_07189_),
    .Y(_07190_));
 sg13g2_a22oi_1 _16671_ (.Y(_07191_),
    .B1(net4557),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][27] ),
    .A2(net4653),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][27] ));
 sg13g2_a22oi_1 _16672_ (.Y(_07192_),
    .B1(net4511),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][27] ),
    .A2(net4602),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][27] ));
 sg13g2_a21o_1 _16673_ (.A2(_07192_),
    .A1(_07191_),
    .B1(net4486),
    .X(_07193_));
 sg13g2_a22oi_1 _16674_ (.Y(_07194_),
    .B1(net4507),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][27] ),
    .A2(net4552),
    .A1(\m_sys.m_ram.m_ram.r_mem[10][27] ));
 sg13g2_a22oi_1 _16675_ (.Y(_07195_),
    .B1(net4598),
    .B2(\m_sys.m_ram.m_ram.r_mem[8][27] ),
    .A2(net4646),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][27] ));
 sg13g2_a21oi_1 _16676_ (.A1(_07194_),
    .A2(_07195_),
    .Y(_07196_),
    .B1(net4474));
 sg13g2_a22oi_1 _16677_ (.Y(_07197_),
    .B1(net4599),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][27] ),
    .A2(net4647),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][27] ));
 sg13g2_a22oi_1 _16678_ (.Y(_07198_),
    .B1(net4508),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][27] ),
    .A2(net4553),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][27] ));
 sg13g2_a21oi_1 _16679_ (.A1(_07197_),
    .A2(_07198_),
    .Y(_07199_),
    .B1(net4456));
 sg13g2_a22oi_1 _16680_ (.Y(_07200_),
    .B1(net4553),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][27] ),
    .A2(net4645),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][27] ));
 sg13g2_a22oi_1 _16681_ (.Y(_07201_),
    .B1(net4513),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][27] ),
    .A2(net4603),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][27] ));
 sg13g2_a21oi_2 _16682_ (.B1(net4499),
    .Y(_07202_),
    .A2(_07201_),
    .A1(_07200_));
 sg13g2_a22oi_1 _16683_ (.Y(_07203_),
    .B1(net4515),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][27] ),
    .A2(net4650),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][27] ));
 sg13g2_a22oi_1 _16684_ (.Y(_07204_),
    .B1(net4560),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][27] ),
    .A2(net4605),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][27] ));
 sg13g2_a21oi_2 _16685_ (.B1(net4462),
    .Y(_07205_),
    .A2(_07204_),
    .A1(_07203_));
 sg13g2_nor4_2 _16686_ (.A(_07196_),
    .B(_07199_),
    .C(_07202_),
    .Y(_07206_),
    .D(_07205_));
 sg13g2_nand4_1 _16687_ (.B(_07190_),
    .C(_07193_),
    .A(net4355),
    .Y(_07207_),
    .D(_07206_));
 sg13g2_o21ai_1 _16688_ (.B1(_07207_),
    .Y(_07208_),
    .A1(net3420),
    .A2(net4355));
 sg13g2_nor2_1 _16689_ (.A(net5368),
    .B(_07208_),
    .Y(_01125_));
 sg13g2_a22oi_1 _16690_ (.Y(_07209_),
    .B1(net4514),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][28] ),
    .A2(net4559),
    .A1(\m_sys.m_ram.m_ram.r_mem[26][28] ));
 sg13g2_a22oi_1 _16691_ (.Y(_07210_),
    .B1(net4607),
    .B2(\m_sys.m_ram.m_ram.r_mem[24][28] ),
    .A2(net4649),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][28] ));
 sg13g2_a21oi_1 _16692_ (.A1(_07209_),
    .A2(_07210_),
    .Y(_07211_),
    .B1(net4500));
 sg13g2_a22oi_1 _16693_ (.Y(_07212_),
    .B1(net4513),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][28] ),
    .A2(net4604),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][28] ));
 sg13g2_a22oi_1 _16694_ (.Y(_07213_),
    .B1(net4559),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][28] ),
    .A2(net4649),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][28] ));
 sg13g2_a21oi_1 _16695_ (.A1(_07212_),
    .A2(_07213_),
    .Y(_07214_),
    .B1(net4457));
 sg13g2_a22oi_1 _16696_ (.Y(_07215_),
    .B1(net4554),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][28] ),
    .A2(net4644),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][28] ));
 sg13g2_a22oi_1 _16697_ (.Y(_07216_),
    .B1(net4507),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][28] ),
    .A2(net4598),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][28] ));
 sg13g2_a21oi_2 _16698_ (.B1(net4468),
    .Y(_07217_),
    .A2(_07216_),
    .A1(_07215_));
 sg13g2_a22oi_1 _16699_ (.Y(_07218_),
    .B1(net4556),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][28] ),
    .A2(net4652),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][28] ));
 sg13g2_a22oi_1 _16700_ (.Y(_07219_),
    .B1(net4510),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][28] ),
    .A2(net4600),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][28] ));
 sg13g2_a21oi_1 _16701_ (.A1(_07218_),
    .A2(_07219_),
    .Y(_07220_),
    .B1(net4480));
 sg13g2_a22oi_1 _16702_ (.Y(_07221_),
    .B1(net4514),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][28] ),
    .A2(net4558),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][28] ));
 sg13g2_a22oi_1 _16703_ (.Y(_07222_),
    .B1(net4604),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][28] ),
    .A2(net4649),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][28] ));
 sg13g2_a21oi_1 _16704_ (.A1(_07221_),
    .A2(_07222_),
    .Y(_07223_),
    .B1(net4449));
 sg13g2_a22oi_1 _16705_ (.Y(_07224_),
    .B1(net4555),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][28] ),
    .A2(net4652),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][28] ));
 sg13g2_a22oi_1 _16706_ (.Y(_07225_),
    .B1(net4510),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][28] ),
    .A2(net4601),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][28] ));
 sg13g2_a21oi_1 _16707_ (.A1(_07224_),
    .A2(_07225_),
    .Y(_07226_),
    .B1(net4486));
 sg13g2_a22oi_1 _16708_ (.Y(_07227_),
    .B1(net4600),
    .B2(\m_sys.m_ram.m_ram.r_mem[8][28] ),
    .A2(net4646),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][28] ));
 sg13g2_a22oi_1 _16709_ (.Y(_07228_),
    .B1(net4509),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][28] ),
    .A2(net4555),
    .A1(\m_sys.m_ram.m_ram.r_mem[10][28] ));
 sg13g2_a21oi_1 _16710_ (.A1(_07227_),
    .A2(_07228_),
    .Y(_07229_),
    .B1(net4474));
 sg13g2_a22oi_1 _16711_ (.Y(_07230_),
    .B1(net4516),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][28] ),
    .A2(net4561),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][28] ));
 sg13g2_a22oi_1 _16712_ (.Y(_07231_),
    .B1(net4606),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][28] ),
    .A2(net4653),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][28] ));
 sg13g2_a21o_1 _16713_ (.A2(_07231_),
    .A1(_07230_),
    .B1(net4463),
    .X(_07232_));
 sg13g2_nor3_2 _16714_ (.A(_07211_),
    .B(_07214_),
    .C(_07223_),
    .Y(_07233_));
 sg13g2_nor4_2 _16715_ (.A(_07217_),
    .B(_07220_),
    .C(_07226_),
    .Y(_07234_),
    .D(_07229_));
 sg13g2_nand4_1 _16716_ (.B(_07232_),
    .C(_07233_),
    .A(net4356),
    .Y(_07235_),
    .D(_07234_));
 sg13g2_o21ai_1 _16717_ (.B1(_07235_),
    .Y(_07236_),
    .A1(net3427),
    .A2(net4356));
 sg13g2_nor2_1 _16718_ (.A(net5367),
    .B(_07236_),
    .Y(_01126_));
 sg13g2_a22oi_1 _16719_ (.Y(_07237_),
    .B1(net4509),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][29] ),
    .A2(net4556),
    .A1(\m_sys.m_ram.m_ram.r_mem[2][29] ));
 sg13g2_a22oi_1 _16720_ (.Y(_07238_),
    .B1(net4600),
    .B2(\m_sys.m_ram.m_ram.r_mem[0][29] ),
    .A2(net4647),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][29] ));
 sg13g2_a21oi_1 _16721_ (.A1(_07237_),
    .A2(_07238_),
    .Y(_07239_),
    .B1(net4480));
 sg13g2_a22oi_1 _16722_ (.Y(_07240_),
    .B1(net4553),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][29] ),
    .A2(net4645),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][29] ));
 sg13g2_a22oi_1 _16723_ (.Y(_07241_),
    .B1(net4513),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][29] ),
    .A2(net4603),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][29] ));
 sg13g2_a21oi_2 _16724_ (.B1(net4499),
    .Y(_07242_),
    .A2(_07241_),
    .A1(_07240_));
 sg13g2_a22oi_1 _16725_ (.Y(_07243_),
    .B1(net4555),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][29] ),
    .A2(net4652),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][29] ));
 sg13g2_a22oi_1 _16726_ (.Y(_07244_),
    .B1(net4509),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][29] ),
    .A2(net4601),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][29] ));
 sg13g2_a21oi_2 _16727_ (.B1(net4486),
    .Y(_07245_),
    .A2(_07244_),
    .A1(_07243_));
 sg13g2_a22oi_1 _16728_ (.Y(_07246_),
    .B1(net4561),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][29] ),
    .A2(net4651),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][29] ));
 sg13g2_a22oi_1 _16729_ (.Y(_07247_),
    .B1(net4515),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][29] ),
    .A2(net4606),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][29] ));
 sg13g2_a21oi_1 _16730_ (.A1(_07246_),
    .A2(_07247_),
    .Y(_07248_),
    .B1(net4448));
 sg13g2_a22oi_1 _16731_ (.Y(_07249_),
    .B1(net4552),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][29] ),
    .A2(net4599),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][29] ));
 sg13g2_a22oi_1 _16732_ (.Y(_07250_),
    .B1(net4508),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][29] ),
    .A2(net4644),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][29] ));
 sg13g2_a21oi_1 _16733_ (.A1(_07249_),
    .A2(_07250_),
    .Y(_07251_),
    .B1(net4474));
 sg13g2_a22oi_1 _16734_ (.Y(_07252_),
    .B1(net4515),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][29] ),
    .A2(net4653),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][29] ));
 sg13g2_a22oi_1 _16735_ (.Y(_07253_),
    .B1(net4560),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][29] ),
    .A2(net4605),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][29] ));
 sg13g2_a21o_1 _16736_ (.A2(_07253_),
    .A1(_07252_),
    .B1(net4462),
    .X(_07254_));
 sg13g2_a22oi_1 _16737_ (.Y(_07255_),
    .B1(net4513),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][29] ),
    .A2(net4558),
    .A1(\m_sys.m_ram.m_ram.r_mem[30][29] ));
 sg13g2_a22oi_1 _16738_ (.Y(_07256_),
    .B1(net4603),
    .B2(\m_sys.m_ram.m_ram.r_mem[28][29] ),
    .A2(net4650),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][29] ));
 sg13g2_a21oi_2 _16739_ (.B1(net4456),
    .Y(_07257_),
    .A2(_07256_),
    .A1(_07255_));
 sg13g2_a22oi_1 _16740_ (.Y(_07258_),
    .B1(net4552),
    .B2(\m_sys.m_ram.m_ram.r_mem[22][29] ),
    .A2(net4644),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][29] ));
 sg13g2_a22oi_1 _16741_ (.Y(_07259_),
    .B1(net4507),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][29] ),
    .A2(net4598),
    .A1(\m_sys.m_ram.m_ram.r_mem[20][29] ));
 sg13g2_a21oi_1 _16742_ (.A1(_07258_),
    .A2(_07259_),
    .Y(_07260_),
    .B1(net4468));
 sg13g2_nor3_1 _16743_ (.A(_07239_),
    .B(_07248_),
    .C(_07257_),
    .Y(_07261_));
 sg13g2_nor4_2 _16744_ (.A(_07242_),
    .B(_07245_),
    .C(_07251_),
    .Y(_07262_),
    .D(_07260_));
 sg13g2_nand4_1 _16745_ (.B(_07254_),
    .C(_07261_),
    .A(net4355),
    .Y(_07263_),
    .D(_07262_));
 sg13g2_o21ai_1 _16746_ (.B1(_07263_),
    .Y(_07264_),
    .A1(net3432),
    .A2(net4355));
 sg13g2_nor2_1 _16747_ (.A(net5367),
    .B(_07264_),
    .Y(_01127_));
 sg13g2_a22oi_1 _16748_ (.Y(_07265_),
    .B1(net4598),
    .B2(\m_sys.m_ram.m_ram.r_mem[20][30] ),
    .A2(net4644),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][30] ));
 sg13g2_a22oi_1 _16749_ (.Y(_07266_),
    .B1(net4507),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][30] ),
    .A2(net4552),
    .A1(\m_sys.m_ram.m_ram.r_mem[22][30] ));
 sg13g2_a21oi_2 _16750_ (.B1(net4468),
    .Y(_07267_),
    .A2(_07266_),
    .A1(_07265_));
 sg13g2_a22oi_1 _16751_ (.Y(_07268_),
    .B1(net4555),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][30] ),
    .A2(net4646),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][30] ));
 sg13g2_a22oi_1 _16752_ (.Y(_07269_),
    .B1(net4509),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][30] ),
    .A2(net4600),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][30] ));
 sg13g2_a21oi_1 _16753_ (.A1(_07268_),
    .A2(_07269_),
    .Y(_07270_),
    .B1(net4480));
 sg13g2_a22oi_1 _16754_ (.Y(_07271_),
    .B1(net4553),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][30] ),
    .A2(net4645),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][30] ));
 sg13g2_a22oi_1 _16755_ (.Y(_07272_),
    .B1(net4513),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][30] ),
    .A2(net4603),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][30] ));
 sg13g2_a21oi_2 _16756_ (.B1(net4499),
    .Y(_07273_),
    .A2(_07272_),
    .A1(_07271_));
 sg13g2_nor3_1 _16757_ (.A(_07267_),
    .B(_07270_),
    .C(_07273_),
    .Y(_07274_));
 sg13g2_a22oi_1 _16758_ (.Y(_07275_),
    .B1(net4512),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][30] ),
    .A2(net4647),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][30] ));
 sg13g2_a22oi_1 _16759_ (.Y(_07276_),
    .B1(net4558),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][30] ),
    .A2(net4604),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][30] ));
 sg13g2_a21o_1 _16760_ (.A2(_07276_),
    .A1(_07275_),
    .B1(net4456),
    .X(_07277_));
 sg13g2_a22oi_1 _16761_ (.Y(_07278_),
    .B1(net4560),
    .B2(\m_sys.m_ram.m_ram.r_mem[18][30] ),
    .A2(net4653),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][30] ));
 sg13g2_a22oi_1 _16762_ (.Y(_07279_),
    .B1(net4515),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][30] ),
    .A2(net4605),
    .A1(\m_sys.m_ram.m_ram.r_mem[16][30] ));
 sg13g2_a21oi_1 _16763_ (.A1(_07278_),
    .A2(_07279_),
    .Y(_07280_),
    .B1(net4462));
 sg13g2_a22oi_1 _16764_ (.Y(_07281_),
    .B1(net4515),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][30] ),
    .A2(net4560),
    .A1(\m_sys.m_ram.m_ram.r_mem[10][30] ));
 sg13g2_a22oi_1 _16765_ (.Y(_07282_),
    .B1(net4605),
    .B2(\m_sys.m_ram.m_ram.r_mem[8][30] ),
    .A2(net4650),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][30] ));
 sg13g2_a21oi_1 _16766_ (.A1(_07281_),
    .A2(_07282_),
    .Y(_07283_),
    .B1(net4476));
 sg13g2_a22oi_1 _16767_ (.Y(_07284_),
    .B1(net4516),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][30] ),
    .A2(net4561),
    .A1(\m_sys.m_ram.m_ram.r_mem[6][30] ));
 sg13g2_a22oi_1 _16768_ (.Y(_07285_),
    .B1(net4606),
    .B2(\m_sys.m_ram.m_ram.r_mem[4][30] ),
    .A2(net4651),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][30] ));
 sg13g2_a21oi_1 _16769_ (.A1(_07284_),
    .A2(_07285_),
    .Y(_07286_),
    .B1(net4448));
 sg13g2_a22oi_1 _16770_ (.Y(_07287_),
    .B1(net4556),
    .B2(\m_sys.m_ram.m_ram.r_mem[14][30] ),
    .A2(net4652),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][30] ));
 sg13g2_a22oi_1 _16771_ (.Y(_07288_),
    .B1(net4511),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][30] ),
    .A2(net4602),
    .A1(\m_sys.m_ram.m_ram.r_mem[12][30] ));
 sg13g2_a21oi_2 _16772_ (.B1(net4486),
    .Y(_07289_),
    .A2(_07288_),
    .A1(_07287_));
 sg13g2_nor4_1 _16773_ (.A(_07280_),
    .B(_07283_),
    .C(_07286_),
    .D(_07289_),
    .Y(_07290_));
 sg13g2_nand4_1 _16774_ (.B(_07274_),
    .C(_07277_),
    .A(net4357),
    .Y(_07291_),
    .D(_07290_));
 sg13g2_o21ai_1 _16775_ (.B1(_07291_),
    .Y(_07292_),
    .A1(net3403),
    .A2(net4355));
 sg13g2_nor2_1 _16776_ (.A(net5367),
    .B(_07292_),
    .Y(_01128_));
 sg13g2_a22oi_1 _16777_ (.Y(_07293_),
    .B1(net4515),
    .B2(\m_sys.m_ram.m_ram.r_mem[19][31] ),
    .A2(net4560),
    .A1(\m_sys.m_ram.m_ram.r_mem[18][31] ));
 sg13g2_a22oi_1 _16778_ (.Y(_07294_),
    .B1(net4605),
    .B2(\m_sys.m_ram.m_ram.r_mem[16][31] ),
    .A2(net4653),
    .A1(\m_sys.m_ram.m_ram.r_mem[17][31] ));
 sg13g2_a21oi_1 _16779_ (.A1(_07293_),
    .A2(_07294_),
    .Y(_07295_),
    .B1(net4462));
 sg13g2_a22oi_1 _16780_ (.Y(_07296_),
    .B1(net4507),
    .B2(\m_sys.m_ram.m_ram.r_mem[23][31] ),
    .A2(net4552),
    .A1(\m_sys.m_ram.m_ram.r_mem[22][31] ));
 sg13g2_a22oi_1 _16781_ (.Y(_07297_),
    .B1(net4598),
    .B2(\m_sys.m_ram.m_ram.r_mem[20][31] ),
    .A2(net4644),
    .A1(\m_sys.m_ram.m_ram.r_mem[21][31] ));
 sg13g2_a21oi_2 _16782_ (.B1(net4468),
    .Y(_07298_),
    .A2(_07297_),
    .A1(_07296_));
 sg13g2_a22oi_1 _16783_ (.Y(_07299_),
    .B1(net4554),
    .B2(\m_sys.m_ram.m_ram.r_mem[30][31] ),
    .A2(net4645),
    .A1(\m_sys.m_ram.m_ram.r_mem[29][31] ));
 sg13g2_a22oi_1 _16784_ (.Y(_07300_),
    .B1(net4513),
    .B2(\m_sys.m_ram.m_ram.r_mem[31][31] ),
    .A2(net4604),
    .A1(\m_sys.m_ram.m_ram.r_mem[28][31] ));
 sg13g2_a21oi_1 _16785_ (.A1(_07299_),
    .A2(_07300_),
    .Y(_07301_),
    .B1(net4456));
 sg13g2_a22oi_1 _16786_ (.Y(_07302_),
    .B1(net4554),
    .B2(\m_sys.m_ram.m_ram.r_mem[10][31] ),
    .A2(net4644),
    .A1(\m_sys.m_ram.m_ram.r_mem[9][31] ));
 sg13g2_a22oi_1 _16787_ (.Y(_07303_),
    .B1(net4507),
    .B2(\m_sys.m_ram.m_ram.r_mem[11][31] ),
    .A2(net4599),
    .A1(\m_sys.m_ram.m_ram.r_mem[8][31] ));
 sg13g2_a21oi_2 _16788_ (.B1(net4474),
    .Y(_07304_),
    .A2(_07303_),
    .A1(_07302_));
 sg13g2_a22oi_1 _16789_ (.Y(_07305_),
    .B1(net4558),
    .B2(\m_sys.m_ram.m_ram.r_mem[6][31] ),
    .A2(net4650),
    .A1(\m_sys.m_ram.m_ram.r_mem[5][31] ));
 sg13g2_a22oi_1 _16790_ (.Y(_07306_),
    .B1(net4514),
    .B2(\m_sys.m_ram.m_ram.r_mem[7][31] ),
    .A2(net4604),
    .A1(\m_sys.m_ram.m_ram.r_mem[4][31] ));
 sg13g2_a21oi_1 _16791_ (.A1(_07305_),
    .A2(_07306_),
    .Y(_07307_),
    .B1(net4448));
 sg13g2_a22oi_1 _16792_ (.Y(_07308_),
    .B1(net4509),
    .B2(\m_sys.m_ram.m_ram.r_mem[3][31] ),
    .A2(net4652),
    .A1(\m_sys.m_ram.m_ram.r_mem[1][31] ));
 sg13g2_a22oi_1 _16793_ (.Y(_07309_),
    .B1(net4555),
    .B2(\m_sys.m_ram.m_ram.r_mem[2][31] ),
    .A2(net4600),
    .A1(\m_sys.m_ram.m_ram.r_mem[0][31] ));
 sg13g2_a21o_1 _16794_ (.A2(_07309_),
    .A1(_07308_),
    .B1(net4480),
    .X(_07310_));
 sg13g2_a22oi_1 _16795_ (.Y(_07311_),
    .B1(net4510),
    .B2(\m_sys.m_ram.m_ram.r_mem[15][31] ),
    .A2(net4556),
    .A1(\m_sys.m_ram.m_ram.r_mem[14][31] ));
 sg13g2_a22oi_1 _16796_ (.Y(_07312_),
    .B1(net4600),
    .B2(\m_sys.m_ram.m_ram.r_mem[12][31] ),
    .A2(net4652),
    .A1(\m_sys.m_ram.m_ram.r_mem[13][31] ));
 sg13g2_a21oi_1 _16797_ (.A1(_07311_),
    .A2(_07312_),
    .Y(_07313_),
    .B1(net4486));
 sg13g2_a22oi_1 _16798_ (.Y(_07314_),
    .B1(net4558),
    .B2(\m_sys.m_ram.m_ram.r_mem[26][31] ),
    .A2(net4649),
    .A1(\m_sys.m_ram.m_ram.r_mem[25][31] ));
 sg13g2_a22oi_1 _16799_ (.Y(_07315_),
    .B1(net4513),
    .B2(\m_sys.m_ram.m_ram.r_mem[27][31] ),
    .A2(net4603),
    .A1(\m_sys.m_ram.m_ram.r_mem[24][31] ));
 sg13g2_a21oi_2 _16800_ (.B1(net4499),
    .Y(_07316_),
    .A2(_07315_),
    .A1(_07314_));
 sg13g2_nor3_1 _16801_ (.A(_07295_),
    .B(_07298_),
    .C(_07313_),
    .Y(_07317_));
 sg13g2_nor4_2 _16802_ (.A(_07301_),
    .B(_07304_),
    .C(_07307_),
    .Y(_07318_),
    .D(_07316_));
 sg13g2_nand4_1 _16803_ (.B(_07310_),
    .C(_07317_),
    .A(net4355),
    .Y(_07319_),
    .D(_07318_));
 sg13g2_o21ai_1 _16804_ (.B1(_07319_),
    .Y(_07320_),
    .A1(net3430),
    .A2(net4355));
 sg13g2_nor2_1 _16805_ (.A(net5367),
    .B(_07320_),
    .Y(_01129_));
 sg13g2_nor2_2 _16806_ (.A(net4506),
    .B(net4485),
    .Y(_07321_));
 sg13g2_nor2b_1 _16807_ (.A(net4317),
    .B_N(_07321_),
    .Y(_07322_));
 sg13g2_nor2_1 _16808_ (.A(net2310),
    .B(net4105),
    .Y(_07323_));
 sg13g2_a21oi_1 _16809_ (.A1(net5022),
    .A2(net4105),
    .Y(_01130_),
    .B1(_07323_));
 sg13g2_nor2_1 _16810_ (.A(net2377),
    .B(net4105),
    .Y(_07324_));
 sg13g2_a21oi_1 _16811_ (.A1(net4811),
    .A2(net4105),
    .Y(_01131_),
    .B1(_07324_));
 sg13g2_nor2_1 _16812_ (.A(net2393),
    .B(net4106),
    .Y(_07325_));
 sg13g2_a21oi_1 _16813_ (.A1(net5018),
    .A2(net4106),
    .Y(_01132_),
    .B1(_07325_));
 sg13g2_nor2_1 _16814_ (.A(net2652),
    .B(net4106),
    .Y(_07326_));
 sg13g2_a21oi_1 _16815_ (.A1(net4809),
    .A2(net4106),
    .Y(_01133_),
    .B1(_07326_));
 sg13g2_nor2_1 _16816_ (.A(net2851),
    .B(net4105),
    .Y(_07327_));
 sg13g2_a21oi_1 _16817_ (.A1(net5011),
    .A2(net4105),
    .Y(_01134_),
    .B1(_07327_));
 sg13g2_nor2_1 _16818_ (.A(net2753),
    .B(net4106),
    .Y(_07328_));
 sg13g2_a21oi_1 _16819_ (.A1(net4801),
    .A2(net4106),
    .Y(_01135_),
    .B1(_07328_));
 sg13g2_nor2_1 _16820_ (.A(net2443),
    .B(net4105),
    .Y(_07329_));
 sg13g2_a21oi_1 _16821_ (.A1(net5005),
    .A2(net4105),
    .Y(_01136_),
    .B1(_07329_));
 sg13g2_nor2_1 _16822_ (.A(net2675),
    .B(net4106),
    .Y(_07330_));
 sg13g2_a21oi_1 _16823_ (.A1(net4798),
    .A2(net4106),
    .Y(_01137_),
    .B1(_07330_));
 sg13g2_nand4_1 _16824_ (.B(\m_sys._m_bootloader_io_b_mem_addr[6] ),
    .C(_02713_),
    .A(\m_sys._m_bootloader_io_b_mem_addr[11] ),
    .Y(_07331_),
    .D(_02715_));
 sg13g2_nand2_1 _16825_ (.Y(_07332_),
    .A(net5268),
    .B(_07331_));
 sg13g2_nand4_1 _16826_ (.B(net4390),
    .C(_04954_),
    .A(net3263),
    .Y(_07333_),
    .D(_07332_));
 sg13g2_or2_1 _16827_ (.X(_07334_),
    .B(_07333_),
    .A(_04905_));
 sg13g2_o21ai_1 _16828_ (.B1(net5380),
    .Y(_07335_),
    .A1(_06015_),
    .A2(net4343));
 sg13g2_a21oi_1 _16829_ (.A1(_02358_),
    .A2(net4343),
    .Y(_01138_),
    .B1(_07335_));
 sg13g2_o21ai_1 _16830_ (.B1(net5380),
    .Y(_07336_),
    .A1(_06019_),
    .A2(net4346));
 sg13g2_a21oi_1 _16831_ (.A1(_02357_),
    .A2(_07334_),
    .Y(_01139_),
    .B1(_07336_));
 sg13g2_o21ai_1 _16832_ (.B1(net5379),
    .Y(_07337_),
    .A1(_06023_),
    .A2(net4341));
 sg13g2_a21oi_1 _16833_ (.A1(_02356_),
    .A2(net4342),
    .Y(_01140_),
    .B1(_07337_));
 sg13g2_nand2b_1 _16834_ (.Y(_07338_),
    .B(_06027_),
    .A_N(net4342));
 sg13g2_a21oi_1 _16835_ (.A1(net3414),
    .A2(net4344),
    .Y(_07339_),
    .B1(net5368));
 sg13g2_nand2_1 _16836_ (.Y(_01141_),
    .A(_07338_),
    .B(_07339_));
 sg13g2_nand2b_1 _16837_ (.Y(_07340_),
    .B(_06031_),
    .A_N(net4342));
 sg13g2_a21oi_1 _16838_ (.A1(net3152),
    .A2(net4342),
    .Y(_07341_),
    .B1(net5368));
 sg13g2_nand2_1 _16839_ (.Y(_01142_),
    .A(_07340_),
    .B(_07341_));
 sg13g2_o21ai_1 _16840_ (.B1(net5380),
    .Y(_07342_),
    .A1(_06035_),
    .A2(net4346));
 sg13g2_a21oi_1 _16841_ (.A1(_02353_),
    .A2(net4346),
    .Y(_01143_),
    .B1(_07342_));
 sg13g2_nand2b_1 _16842_ (.Y(_07343_),
    .B(_06039_),
    .A_N(net4344));
 sg13g2_a21oi_1 _16843_ (.A1(net3381),
    .A2(net4344),
    .Y(_07344_),
    .B1(net5368));
 sg13g2_nand2_1 _16844_ (.Y(_01144_),
    .A(_07343_),
    .B(_07344_));
 sg13g2_o21ai_1 _16845_ (.B1(net5380),
    .Y(_07345_),
    .A1(_05716_),
    .A2(net4343));
 sg13g2_a21oi_1 _16846_ (.A1(_02351_),
    .A2(net4343),
    .Y(_01145_),
    .B1(_07345_));
 sg13g2_o21ai_1 _16847_ (.B1(net5379),
    .Y(_07346_),
    .A1(_04951_),
    .A2(net4341));
 sg13g2_a21oi_1 _16848_ (.A1(_02350_),
    .A2(net4341),
    .Y(_01146_),
    .B1(_07346_));
 sg13g2_o21ai_1 _16849_ (.B1(net5379),
    .Y(_07347_),
    .A1(_04959_),
    .A2(net4341));
 sg13g2_a21oi_1 _16850_ (.A1(_02349_),
    .A2(net4341),
    .Y(_01147_),
    .B1(_07347_));
 sg13g2_a21oi_1 _16851_ (.A1(net3076),
    .A2(net4346),
    .Y(_07348_),
    .B1(net5367));
 sg13g2_o21ai_1 _16852_ (.B1(_07348_),
    .Y(_01148_),
    .A1(_04962_),
    .A2(net4346));
 sg13g2_o21ai_1 _16853_ (.B1(net5380),
    .Y(_07349_),
    .A1(_04965_),
    .A2(net4343));
 sg13g2_a21oi_1 _16854_ (.A1(_02348_),
    .A2(net4343),
    .Y(_01149_),
    .B1(_07349_));
 sg13g2_a21oi_1 _16855_ (.A1(net3319),
    .A2(net4346),
    .Y(_07350_),
    .B1(net5367));
 sg13g2_o21ai_1 _16856_ (.B1(_07350_),
    .Y(_01150_),
    .A1(_04968_),
    .A2(net4346));
 sg13g2_o21ai_1 _16857_ (.B1(net5379),
    .Y(_07351_),
    .A1(_04971_),
    .A2(net4343));
 sg13g2_a21oi_1 _16858_ (.A1(_02346_),
    .A2(net4343),
    .Y(_01151_),
    .B1(_07351_));
 sg13g2_o21ai_1 _16859_ (.B1(net5379),
    .Y(_07352_),
    .A1(_04974_),
    .A2(net4341));
 sg13g2_a21oi_1 _16860_ (.A1(_02345_),
    .A2(net4341),
    .Y(_01152_),
    .B1(_07352_));
 sg13g2_o21ai_1 _16861_ (.B1(net5379),
    .Y(_07353_),
    .A1(_04977_),
    .A2(net4344));
 sg13g2_a21oi_1 _16862_ (.A1(_02344_),
    .A2(net4341),
    .Y(_01153_),
    .B1(_07353_));
 sg13g2_a21oi_1 _16863_ (.A1(_02340_),
    .A2(net9),
    .Y(_07354_),
    .B1(net1));
 sg13g2_nor2_1 _16864_ (.A(net5370),
    .B(_07354_),
    .Y(_01154_));
 sg13g2_a21oi_1 _16865_ (.A1(_02339_),
    .A2(net10),
    .Y(_07355_),
    .B1(net2));
 sg13g2_nor2_1 _16866_ (.A(net5370),
    .B(_07355_),
    .Y(_01155_));
 sg13g2_a21oi_1 _16867_ (.A1(_02338_),
    .A2(net11),
    .Y(_07356_),
    .B1(net3));
 sg13g2_nor2_1 _16868_ (.A(net5370),
    .B(_07356_),
    .Y(_01156_));
 sg13g2_a21oi_1 _16869_ (.A1(_02337_),
    .A2(net12),
    .Y(_07357_),
    .B1(net4));
 sg13g2_nor2_1 _16870_ (.A(net5369),
    .B(_07357_),
    .Y(_01157_));
 sg13g2_a21oi_1 _16871_ (.A1(_02336_),
    .A2(net13),
    .Y(_07358_),
    .B1(net5));
 sg13g2_nor2_1 _16872_ (.A(net5369),
    .B(_07358_),
    .Y(_01158_));
 sg13g2_a21oi_1 _16873_ (.A1(_02335_),
    .A2(net14),
    .Y(_07359_),
    .B1(net6));
 sg13g2_nor2_1 _16874_ (.A(net5369),
    .B(_07359_),
    .Y(_01159_));
 sg13g2_a21oi_1 _16875_ (.A1(_02334_),
    .A2(net15),
    .Y(_07360_),
    .B1(net7));
 sg13g2_nor2_1 _16876_ (.A(net5369),
    .B(_07360_),
    .Y(_01160_));
 sg13g2_a21oi_1 _16877_ (.A1(_02333_),
    .A2(net16),
    .Y(_07361_),
    .B1(net8));
 sg13g2_nor2_1 _16878_ (.A(net5369),
    .B(_07361_),
    .Y(_01161_));
 sg13g2_nor2_2 _16879_ (.A(net5271),
    .B(net4715),
    .Y(_07362_));
 sg13g2_nor2_1 _16880_ (.A(_02648_),
    .B(_02670_),
    .Y(_07363_));
 sg13g2_inv_1 _16881_ (.Y(_07364_),
    .A(net4353));
 sg13g2_a21oi_1 _16882_ (.A1(net2533),
    .A2(_07364_),
    .Y(_07365_),
    .B1(net4446));
 sg13g2_nor2_1 _16883_ (.A(net5368),
    .B(_07365_),
    .Y(_01162_));
 sg13g2_nand2b_2 _16884_ (.Y(_07366_),
    .B(_04920_),
    .A_N(_02600_));
 sg13g2_inv_1 _16885_ (.Y(_07367_),
    .A(net4708));
 sg13g2_a21oi_1 _16886_ (.A1(net3357),
    .A2(net3125),
    .Y(_07368_),
    .B1(net4445));
 sg13g2_a21o_1 _16887_ (.A2(net4445),
    .A1(net3357),
    .B1(_07368_),
    .X(_07369_));
 sg13g2_inv_1 _16888_ (.Y(_01163_),
    .A(_07369_));
 sg13g2_a21o_1 _16889_ (.A2(net4445),
    .A1(net3357),
    .B1(net3291),
    .X(_07370_));
 sg13g2_nand3_1 _16890_ (.B(net3357),
    .C(net4445),
    .A(net3291),
    .Y(_07371_));
 sg13g2_and3_1 _16891_ (.X(_01164_),
    .A(net3125),
    .B(_07370_),
    .C(_07371_));
 sg13g2_o21ai_1 _16892_ (.B1(\m_sys.m_uart.m_rx.r_cstate[1] ),
    .Y(_07372_),
    .A1(_02343_),
    .A2(_07371_));
 sg13g2_a21oi_1 _16893_ (.A1(_02343_),
    .A2(_07371_),
    .Y(_01165_),
    .B1(_07372_));
 sg13g2_nor2_1 _16894_ (.A(net2522),
    .B(net4708),
    .Y(_07373_));
 sg13g2_a221oi_1 _16895_ (.B2(_02342_),
    .C1(_07373_),
    .B1(_07366_),
    .A1(_02364_),
    .Y(_01166_),
    .A2(_02365_));
 sg13g2_nor2_1 _16896_ (.A(net5265),
    .B(net4708),
    .Y(_07374_));
 sg13g2_a221oi_1 _16897_ (.B2(_02341_),
    .C1(_07374_),
    .B1(net4708),
    .A1(_02364_),
    .Y(_01167_),
    .A2(_02365_));
 sg13g2_nor2_1 _16898_ (.A(net5264),
    .B(net4708),
    .Y(_07375_));
 sg13g2_nor2_1 _16899_ (.A(net2752),
    .B(_07367_),
    .Y(_07376_));
 sg13g2_nor3_1 _16900_ (.A(net3126),
    .B(_07375_),
    .C(_07376_),
    .Y(_01168_));
 sg13g2_nor2_1 _16901_ (.A(net5263),
    .B(net4708),
    .Y(_07377_));
 sg13g2_nor2_1 _16902_ (.A(net5264),
    .B(_07367_),
    .Y(_07378_));
 sg13g2_nor3_1 _16903_ (.A(net3126),
    .B(_07377_),
    .C(_07378_),
    .Y(_01169_));
 sg13g2_nor2_1 _16904_ (.A(net3003),
    .B(net4445),
    .Y(_07379_));
 sg13g2_nor2_1 _16905_ (.A(net5262),
    .B(_07366_),
    .Y(_07380_));
 sg13g2_nor3_1 _16906_ (.A(_04923_),
    .B(_07379_),
    .C(_07380_),
    .Y(_01170_));
 sg13g2_nor2_1 _16907_ (.A(net2663),
    .B(_07366_),
    .Y(_07381_));
 sg13g2_nor2_1 _16908_ (.A(net5262),
    .B(net4445),
    .Y(_07382_));
 sg13g2_nor3_1 _16909_ (.A(_04923_),
    .B(_07381_),
    .C(_07382_),
    .Y(_01171_));
 sg13g2_nor2_1 _16910_ (.A(net5260),
    .B(net4708),
    .Y(_07383_));
 sg13g2_nor2_1 _16911_ (.A(net5261),
    .B(net4445),
    .Y(_07384_));
 sg13g2_nor3_1 _16912_ (.A(net3126),
    .B(_07383_),
    .C(_07384_),
    .Y(_01172_));
 sg13g2_nor2_1 _16913_ (.A(net3148),
    .B(net4708),
    .Y(_07385_));
 sg13g2_nor2_1 _16914_ (.A(net5260),
    .B(net4445),
    .Y(_07386_));
 sg13g2_nor3_1 _16915_ (.A(net3126),
    .B(_07385_),
    .C(_07386_),
    .Y(_01173_));
 sg13g2_nor2_1 _16916_ (.A(net2862),
    .B(net4446),
    .Y(_07387_));
 sg13g2_a21oi_1 _16917_ (.A1(_02342_),
    .A2(net4446),
    .Y(_01174_),
    .B1(_07387_));
 sg13g2_nor2_1 _16918_ (.A(net2010),
    .B(net4446),
    .Y(_07388_));
 sg13g2_a21oi_1 _16919_ (.A1(_02341_),
    .A2(net4446),
    .Y(_01175_),
    .B1(_07388_));
 sg13g2_mux2_1 _16920_ (.A0(net2378),
    .A1(net2752),
    .S(net4446),
    .X(_01176_));
 sg13g2_mux2_1 _16921_ (.A0(net2123),
    .A1(net2846),
    .S(_07362_),
    .X(_01177_));
 sg13g2_mux2_1 _16922_ (.A0(net2445),
    .A1(net5263),
    .S(net4446),
    .X(_01178_));
 sg13g2_mux2_1 _16923_ (.A0(net1659),
    .A1(net5262),
    .S(_07362_),
    .X(_01179_));
 sg13g2_mux2_1 _16924_ (.A0(net1657),
    .A1(net5261),
    .S(_07362_),
    .X(_01180_));
 sg13g2_mux2_1 _16925_ (.A0(net2120),
    .A1(net5260),
    .S(net4446),
    .X(_01181_));
 sg13g2_nand2_1 _16926_ (.Y(_07389_),
    .A(net5274),
    .B(net3138));
 sg13g2_o21ai_1 _16927_ (.B1(_07389_),
    .Y(_01182_),
    .A1(net5274),
    .A2(_02677_));
 sg13g2_nand2_1 _16928_ (.Y(_07390_),
    .A(net5235),
    .B(_02692_));
 sg13g2_a21oi_1 _16929_ (.A1(net5269),
    .A2(\m_sys._m_bootloader_io_b_mem_addr[7] ),
    .Y(_07391_),
    .B1(net5280));
 sg13g2_a22oi_1 _16930_ (.Y(_01183_),
    .B1(_07390_),
    .B2(_07391_),
    .A2(_02416_),
    .A1(net5281));
 sg13g2_nand2_1 _16931_ (.Y(_07392_),
    .A(net5235),
    .B(_02688_));
 sg13g2_a21oi_1 _16932_ (.A1(net5269),
    .A2(\m_sys._m_bootloader_io_b_mem_addr[8] ),
    .Y(_07393_),
    .B1(net5280));
 sg13g2_a22oi_1 _16933_ (.Y(_01184_),
    .B1(_07392_),
    .B2(_07393_),
    .A2(_02412_),
    .A1(net5281));
 sg13g2_nand2_1 _16934_ (.Y(_07394_),
    .A(net5235),
    .B(_02690_));
 sg13g2_a21oi_1 _16935_ (.A1(net5269),
    .A2(\m_sys._m_bootloader_io_b_mem_addr[9] ),
    .Y(_07395_),
    .B1(net5280));
 sg13g2_a22oi_1 _16936_ (.Y(_01185_),
    .B1(_07394_),
    .B2(_07395_),
    .A2(_02413_),
    .A1(net5281));
 sg13g2_nand2_1 _16937_ (.Y(_07396_),
    .A(net5235),
    .B(_02687_));
 sg13g2_a21oi_1 _16938_ (.A1(net5269),
    .A2(\m_sys._m_bootloader_io_b_mem_addr[10] ),
    .Y(_07397_),
    .B1(net5280));
 sg13g2_a22oi_1 _16939_ (.Y(_01186_),
    .B1(_07396_),
    .B2(_07397_),
    .A2(_02415_),
    .A1(net5280));
 sg13g2_nand2_1 _16940_ (.Y(_07398_),
    .A(net5235),
    .B(_02696_));
 sg13g2_a21oi_1 _16941_ (.A1(net5270),
    .A2(net3245),
    .Y(_07399_),
    .B1(net5280));
 sg13g2_a22oi_1 _16942_ (.Y(_01187_),
    .B1(_07398_),
    .B2(_07399_),
    .A2(_02414_),
    .A1(net5280));
 sg13g2_nor2_2 _16943_ (.A(net4506),
    .B(net4449),
    .Y(_07400_));
 sg13g2_nor2b_1 _16944_ (.A(net4314),
    .B_N(_07400_),
    .Y(_07401_));
 sg13g2_nor2_1 _16945_ (.A(net2629),
    .B(net4103),
    .Y(_07402_));
 sg13g2_a21oi_1 _16946_ (.A1(net5024),
    .A2(net4103),
    .Y(_01188_),
    .B1(_07402_));
 sg13g2_nor2_1 _16947_ (.A(net2453),
    .B(net4103),
    .Y(_07403_));
 sg13g2_a21oi_1 _16948_ (.A1(net4813),
    .A2(net4103),
    .Y(_01189_),
    .B1(_07403_));
 sg13g2_nor2_1 _16949_ (.A(net2366),
    .B(net4104),
    .Y(_07404_));
 sg13g2_a21oi_1 _16950_ (.A1(net5019),
    .A2(net4104),
    .Y(_01190_),
    .B1(_07404_));
 sg13g2_nor2_1 _16951_ (.A(net2777),
    .B(net4104),
    .Y(_07405_));
 sg13g2_a21oi_1 _16952_ (.A1(net4809),
    .A2(net4104),
    .Y(_01191_),
    .B1(_07405_));
 sg13g2_nor2_1 _16953_ (.A(net2415),
    .B(net4103),
    .Y(_07406_));
 sg13g2_a21oi_1 _16954_ (.A1(net5013),
    .A2(net4103),
    .Y(_01192_),
    .B1(_07406_));
 sg13g2_nor2_1 _16955_ (.A(net2273),
    .B(net4104),
    .Y(_07407_));
 sg13g2_a21oi_1 _16956_ (.A1(net4803),
    .A2(net4104),
    .Y(_01193_),
    .B1(_07407_));
 sg13g2_nor2_1 _16957_ (.A(net2858),
    .B(net4104),
    .Y(_07408_));
 sg13g2_a21oi_1 _16958_ (.A1(net5007),
    .A2(net4104),
    .Y(_01194_),
    .B1(_07408_));
 sg13g2_nor2_1 _16959_ (.A(net2861),
    .B(net4103),
    .Y(_07409_));
 sg13g2_a21oi_1 _16960_ (.A1(net4797),
    .A2(net4103),
    .Y(_01195_),
    .B1(_07409_));
 sg13g2_nand3_1 _16961_ (.B(net4392),
    .C(_02670_),
    .A(net2533),
    .Y(_07410_));
 sg13g2_a21oi_1 _16962_ (.A1(\m_sys.m_uart.r_rx_data[0] ),
    .A2(net4353),
    .Y(_07411_),
    .B1(net4390));
 sg13g2_a22oi_1 _16963_ (.Y(_01196_),
    .B1(_07410_),
    .B2(_07411_),
    .A2(net4388),
    .A1(_02358_));
 sg13g2_a22oi_1 _16964_ (.Y(_07412_),
    .B1(net4353),
    .B2(net2010),
    .A2(net4390),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[1] ));
 sg13g2_inv_1 _16965_ (.Y(_01197_),
    .A(net2011));
 sg13g2_a22oi_1 _16966_ (.Y(_07413_),
    .B1(net4353),
    .B2(net2378),
    .A2(net4389),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[2] ));
 sg13g2_inv_1 _16967_ (.Y(_01198_),
    .A(net2379));
 sg13g2_a22oi_1 _16968_ (.Y(_07414_),
    .B1(_07363_),
    .B2(net2123),
    .A2(net4389),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[3] ));
 sg13g2_inv_1 _16969_ (.Y(_01199_),
    .A(net2124));
 sg13g2_nand3_1 _16970_ (.B(_02670_),
    .C(net5147),
    .A(net4392),
    .Y(_07415_));
 sg13g2_a21oi_1 _16971_ (.A1(net2445),
    .A2(net4353),
    .Y(_07416_),
    .B1(net4389));
 sg13g2_a22oi_1 _16972_ (.Y(_01200_),
    .B1(_07415_),
    .B2(_07416_),
    .A2(net4389),
    .A1(_02354_));
 sg13g2_a22oi_1 _16973_ (.Y(_07417_),
    .B1(net4353),
    .B2(net1659),
    .A2(net4389),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[5] ));
 sg13g2_inv_1 _16974_ (.Y(_01201_),
    .A(net1660));
 sg13g2_a22oi_1 _16975_ (.Y(_07418_),
    .B1(net4353),
    .B2(net1657),
    .A2(net4389),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[6] ));
 sg13g2_inv_1 _16976_ (.Y(_01202_),
    .A(net1658));
 sg13g2_a22oi_1 _16977_ (.Y(_07419_),
    .B1(net4353),
    .B2(net2120),
    .A2(net4389),
    .A1(\m_sys.m_uart.m_rx.io_i_ncycle[7] ));
 sg13g2_inv_1 _16978_ (.Y(_01203_),
    .A(net2121));
 sg13g2_nand2_1 _16979_ (.Y(_07420_),
    .A(net4327),
    .B(_05459_));
 sg13g2_nand2_1 _16980_ (.Y(_07421_),
    .A(net1865),
    .B(_07420_));
 sg13g2_o21ai_1 _16981_ (.B1(_07421_),
    .Y(_01204_),
    .A1(net5041),
    .A2(net4101));
 sg13g2_nand2_1 _16982_ (.Y(_07422_),
    .A(net2090),
    .B(net4102));
 sg13g2_o21ai_1 _16983_ (.B1(_07422_),
    .Y(_01205_),
    .A1(net4877),
    .A2(net4101));
 sg13g2_nand2_1 _16984_ (.Y(_07423_),
    .A(net2162),
    .B(net4102));
 sg13g2_o21ai_1 _16985_ (.B1(_07423_),
    .Y(_01206_),
    .A1(net5036),
    .A2(net4102));
 sg13g2_nand2_1 _16986_ (.Y(_07424_),
    .A(net1671),
    .B(net4102));
 sg13g2_o21ai_1 _16987_ (.B1(_07424_),
    .Y(_01207_),
    .A1(net4869),
    .A2(net4102));
 sg13g2_nand2_1 _16988_ (.Y(_07425_),
    .A(net1929),
    .B(net4101));
 sg13g2_o21ai_1 _16989_ (.B1(_07425_),
    .Y(_01208_),
    .A1(net5030),
    .A2(net4101));
 sg13g2_nand2_1 _16990_ (.Y(_07426_),
    .A(net1667),
    .B(net4102));
 sg13g2_o21ai_1 _16991_ (.B1(_07426_),
    .Y(_01209_),
    .A1(net4864),
    .A2(net4102));
 sg13g2_nand2_1 _16992_ (.Y(_07427_),
    .A(net1689),
    .B(net4101));
 sg13g2_o21ai_1 _16993_ (.B1(_07427_),
    .Y(_01210_),
    .A1(net5029),
    .A2(net4101));
 sg13g2_nand2_1 _16994_ (.Y(_07428_),
    .A(net1823),
    .B(net4101));
 sg13g2_o21ai_1 _16995_ (.B1(_07428_),
    .Y(_01211_),
    .A1(net4863),
    .A2(net4101));
 sg13g2_a21oi_1 _16996_ (.A1(net3302),
    .A2(\m_sys.m_uart.m_tx.r_cstate[1] ),
    .Y(_07429_),
    .B1(_04912_));
 sg13g2_or2_1 _16997_ (.X(_07430_),
    .B(net3303),
    .A(_04913_));
 sg13g2_inv_1 _16998_ (.Y(_01212_),
    .A(_07430_));
 sg13g2_o21ai_1 _16999_ (.B1(\m_sys.m_uart.m_tx.r_cstate[1] ),
    .Y(_07431_),
    .A1(net3208),
    .A2(_04913_));
 sg13g2_nor2_1 _17000_ (.A(_04914_),
    .B(net3209),
    .Y(_01213_));
 sg13g2_o21ai_1 _17001_ (.B1(\m_sys.m_uart.m_tx.r_cstate[1] ),
    .Y(_07432_),
    .A1(net3161),
    .A2(_04914_));
 sg13g2_nor2b_1 _17002_ (.A(net3162),
    .B_N(_04915_),
    .Y(_01214_));
 sg13g2_nand2_1 _17003_ (.Y(_07433_),
    .A(_02364_),
    .B(net4));
 sg13g2_nand3_1 _17004_ (.B(_04922_),
    .C(_07433_),
    .A(net5379),
    .Y(_01215_));
 sg13g2_nor2b_2 _17005_ (.A(net4315),
    .B_N(_05640_),
    .Y(_07434_));
 sg13g2_nor2_1 _17006_ (.A(net2397),
    .B(net4099),
    .Y(_07435_));
 sg13g2_a21oi_1 _17007_ (.A1(net5020),
    .A2(net4099),
    .Y(_01216_),
    .B1(_07435_));
 sg13g2_nor2_1 _17008_ (.A(net2210),
    .B(net4100),
    .Y(_07436_));
 sg13g2_a21oi_1 _17009_ (.A1(net4812),
    .A2(net4100),
    .Y(_01217_),
    .B1(_07436_));
 sg13g2_nor2_1 _17010_ (.A(net2508),
    .B(net4099),
    .Y(_07437_));
 sg13g2_a21oi_1 _17011_ (.A1(net5016),
    .A2(net4099),
    .Y(_01218_),
    .B1(_07437_));
 sg13g2_nor2_1 _17012_ (.A(net2448),
    .B(net4099),
    .Y(_07438_));
 sg13g2_a21oi_1 _17013_ (.A1(net4805),
    .A2(net4099),
    .Y(_01219_),
    .B1(_07438_));
 sg13g2_nor2_1 _17014_ (.A(net2226),
    .B(net4100),
    .Y(_07439_));
 sg13g2_a21oi_1 _17015_ (.A1(net5013),
    .A2(net4100),
    .Y(_01220_),
    .B1(_07439_));
 sg13g2_nor2_1 _17016_ (.A(net2465),
    .B(net4100),
    .Y(_07440_));
 sg13g2_a21oi_1 _17017_ (.A1(net4802),
    .A2(net4100),
    .Y(_01221_),
    .B1(_07440_));
 sg13g2_nor2_1 _17018_ (.A(net2679),
    .B(net4099),
    .Y(_07441_));
 sg13g2_a21oi_1 _17019_ (.A1(net5006),
    .A2(net4099),
    .Y(_01222_),
    .B1(_07441_));
 sg13g2_nor2_1 _17020_ (.A(net2640),
    .B(net4100),
    .Y(_07442_));
 sg13g2_a21oi_1 _17021_ (.A1(net4796),
    .A2(net4100),
    .Y(_01223_),
    .B1(_07442_));
 sg13g2_nand2_1 _17022_ (.Y(_07443_),
    .A(net4322),
    .B(_05420_));
 sg13g2_nand2_1 _17023_ (.Y(_07444_),
    .A(net2069),
    .B(net4098));
 sg13g2_o21ai_1 _17024_ (.B1(_07444_),
    .Y(_01224_),
    .A1(net4855),
    .A2(net4098));
 sg13g2_nand2_1 _17025_ (.Y(_07445_),
    .A(net2128),
    .B(net4097));
 sg13g2_o21ai_1 _17026_ (.B1(_07445_),
    .Y(_01225_),
    .A1(net4851),
    .A2(net4097));
 sg13g2_nand2_1 _17027_ (.Y(_07446_),
    .A(net1681),
    .B(net4098));
 sg13g2_o21ai_1 _17028_ (.B1(_07446_),
    .Y(_01226_),
    .A1(net4844),
    .A2(net4098));
 sg13g2_nand2_1 _17029_ (.Y(_07447_),
    .A(net1832),
    .B(net4097));
 sg13g2_o21ai_1 _17030_ (.B1(_07447_),
    .Y(_01227_),
    .A1(net4839),
    .A2(net4097));
 sg13g2_nand2_1 _17031_ (.Y(_07448_),
    .A(net2033),
    .B(net4098));
 sg13g2_o21ai_1 _17032_ (.B1(_07448_),
    .Y(_01228_),
    .A1(net4836),
    .A2(net4098));
 sg13g2_nand2_1 _17033_ (.Y(_07449_),
    .A(net2012),
    .B(net4097));
 sg13g2_o21ai_1 _17034_ (.B1(_07449_),
    .Y(_01229_),
    .A1(net4829),
    .A2(net4097));
 sg13g2_nand2_1 _17035_ (.Y(_07450_),
    .A(net1903),
    .B(net4097));
 sg13g2_o21ai_1 _17036_ (.B1(_07450_),
    .Y(_01230_),
    .A1(net4822),
    .A2(net4097));
 sg13g2_nand2_1 _17037_ (.Y(_07451_),
    .A(net2116),
    .B(net4098));
 sg13g2_o21ai_1 _17038_ (.B1(_07451_),
    .Y(_01231_),
    .A1(net4815),
    .A2(_07443_));
 sg13g2_nor2_1 _17039_ (.A(_02714_),
    .B(net4999),
    .Y(_07452_));
 sg13g2_a21oi_1 _17040_ (.A1(_02704_),
    .A2(_03498_),
    .Y(_07453_),
    .B1(_07452_));
 sg13g2_nor2b_2 _17041_ (.A(_07453_),
    .B_N(_04903_),
    .Y(_07454_));
 sg13g2_nand2b_1 _17042_ (.Y(_07455_),
    .B(_07454_),
    .A_N(net4393));
 sg13g2_o21ai_1 _17043_ (.B1(net5383),
    .Y(_07456_),
    .A1(_06015_),
    .A2(net4340));
 sg13g2_a21oi_1 _17044_ (.A1(_02340_),
    .A2(net4340),
    .Y(_01232_),
    .B1(_07456_));
 sg13g2_o21ai_1 _17045_ (.B1(net5383),
    .Y(_07457_),
    .A1(_06019_),
    .A2(net4340));
 sg13g2_a21oi_1 _17046_ (.A1(_02339_),
    .A2(net4340),
    .Y(_01233_),
    .B1(_07457_));
 sg13g2_o21ai_1 _17047_ (.B1(net5382),
    .Y(_07458_),
    .A1(_06023_),
    .A2(net4340));
 sg13g2_a21oi_1 _17048_ (.A1(_02338_),
    .A2(net4340),
    .Y(_01234_),
    .B1(_07458_));
 sg13g2_o21ai_1 _17049_ (.B1(net5382),
    .Y(_07459_),
    .A1(_06027_),
    .A2(net4340));
 sg13g2_a21oi_1 _17050_ (.A1(_02337_),
    .A2(net4340),
    .Y(_01235_),
    .B1(_07459_));
 sg13g2_o21ai_1 _17051_ (.B1(net5381),
    .Y(_07460_),
    .A1(_06031_),
    .A2(net4339));
 sg13g2_a21oi_1 _17052_ (.A1(_02336_),
    .A2(net4339),
    .Y(_01236_),
    .B1(_07460_));
 sg13g2_o21ai_1 _17053_ (.B1(net5381),
    .Y(_07461_),
    .A1(_06035_),
    .A2(net4339));
 sg13g2_a21oi_1 _17054_ (.A1(_02335_),
    .A2(net4339),
    .Y(_01237_),
    .B1(_07461_));
 sg13g2_o21ai_1 _17055_ (.B1(net5381),
    .Y(_07462_),
    .A1(_06039_),
    .A2(net4339));
 sg13g2_a21oi_1 _17056_ (.A1(_02334_),
    .A2(net4339),
    .Y(_01238_),
    .B1(_07462_));
 sg13g2_o21ai_1 _17057_ (.B1(net5381),
    .Y(_07463_),
    .A1(_05716_),
    .A2(net4339));
 sg13g2_a21oi_1 _17058_ (.A1(_02333_),
    .A2(net4339),
    .Y(_01239_),
    .B1(_07463_));
 sg13g2_nand2_2 _17059_ (.Y(_07464_),
    .A(\m_sys.m_core.r_ctrl_wb_en ),
    .B(_05609_));
 sg13g2_or2_1 _17060_ (.X(_07465_),
    .B(_07464_),
    .A(_00145_));
 sg13g2_nand2_1 _17061_ (.Y(_07466_),
    .A(\m_sys.m_core.m_gpr.io_b_write_addr[0] ),
    .B(\m_sys.m_core.m_gpr.io_b_write_addr[1] ));
 sg13g2_nor2_1 _17062_ (.A(_07465_),
    .B(_07466_),
    .Y(_07467_));
 sg13g2_nor2_1 _17063_ (.A(net2973),
    .B(net4437),
    .Y(_07468_));
 sg13g2_a21oi_1 _17064_ (.A1(_02397_),
    .A2(net4437),
    .Y(_01240_),
    .B1(_07468_));
 sg13g2_mux2_1 _17065_ (.A0(net3104),
    .A1(\m_sys.m_core.m_bru.io_i_s1[1] ),
    .S(net4438),
    .X(_01241_));
 sg13g2_nor2_1 _17066_ (.A(net3063),
    .B(net4443),
    .Y(_07469_));
 sg13g2_a21oi_1 _17067_ (.A1(_02371_),
    .A2(net4443),
    .Y(_01242_),
    .B1(_07469_));
 sg13g2_mux2_1 _17068_ (.A0(net3092),
    .A1(net5314),
    .S(net4443),
    .X(_01243_));
 sg13g2_mux2_1 _17069_ (.A0(net3110),
    .A1(\m_sys.m_core.m_bru.io_i_s1[4] ),
    .S(net4438),
    .X(_01244_));
 sg13g2_mux2_1 _17070_ (.A0(net2895),
    .A1(net5319),
    .S(net4435),
    .X(_01245_));
 sg13g2_nor2_1 _17071_ (.A(net2887),
    .B(net4437),
    .Y(_07470_));
 sg13g2_a21oi_1 _17072_ (.A1(_02386_),
    .A2(net4437),
    .Y(_01246_),
    .B1(_07470_));
 sg13g2_nor2_1 _17073_ (.A(net2808),
    .B(net4437),
    .Y(_07471_));
 sg13g2_a21oi_1 _17074_ (.A1(_02385_),
    .A2(net4437),
    .Y(_01247_),
    .B1(_07471_));
 sg13g2_mux2_1 _17075_ (.A0(net2962),
    .A1(net5321),
    .S(net4441),
    .X(_01248_));
 sg13g2_nor2_1 _17076_ (.A(net2996),
    .B(net4438),
    .Y(_07472_));
 sg13g2_a21oi_1 _17077_ (.A1(_02384_),
    .A2(net4437),
    .Y(_01249_),
    .B1(_07472_));
 sg13g2_nor2_1 _17078_ (.A(net3077),
    .B(net4438),
    .Y(_07473_));
 sg13g2_a21oi_1 _17079_ (.A1(_02383_),
    .A2(net4437),
    .Y(_01250_),
    .B1(_07473_));
 sg13g2_nor2_1 _17080_ (.A(net2956),
    .B(net4441),
    .Y(_07474_));
 sg13g2_a21oi_1 _17081_ (.A1(_02381_),
    .A2(net4441),
    .Y(_01251_),
    .B1(_07474_));
 sg13g2_nor2_1 _17082_ (.A(net2835),
    .B(net4440),
    .Y(_07475_));
 sg13g2_a21oi_1 _17083_ (.A1(_02399_),
    .A2(net4440),
    .Y(_01252_),
    .B1(_07475_));
 sg13g2_nor2_1 _17084_ (.A(net2943),
    .B(net4441),
    .Y(_07476_));
 sg13g2_a21oi_1 _17085_ (.A1(net5225),
    .A2(net4441),
    .Y(_01253_),
    .B1(_07476_));
 sg13g2_nor2_1 _17086_ (.A(net2979),
    .B(net4442),
    .Y(_07477_));
 sg13g2_a21oi_1 _17087_ (.A1(_02400_),
    .A2(net4442),
    .Y(_01254_),
    .B1(_07477_));
 sg13g2_nor2_1 _17088_ (.A(net2847),
    .B(net4443),
    .Y(_07478_));
 sg13g2_a21oi_1 _17089_ (.A1(_02445_),
    .A2(net4443),
    .Y(_01255_),
    .B1(_07478_));
 sg13g2_nor2_1 _17090_ (.A(net2941),
    .B(net4442),
    .Y(_07479_));
 sg13g2_a21oi_1 _17091_ (.A1(net5187),
    .A2(net4442),
    .Y(_01256_),
    .B1(_07479_));
 sg13g2_nor2_1 _17092_ (.A(net2908),
    .B(net4442),
    .Y(_07480_));
 sg13g2_a21oi_1 _17093_ (.A1(net5180),
    .A2(net4442),
    .Y(_01257_),
    .B1(_07480_));
 sg13g2_nor2_1 _17094_ (.A(net2958),
    .B(net4443),
    .Y(_07481_));
 sg13g2_a21oi_1 _17095_ (.A1(_02450_),
    .A2(net4443),
    .Y(_01258_),
    .B1(_07481_));
 sg13g2_nor2_1 _17096_ (.A(net3054),
    .B(net4442),
    .Y(_07482_));
 sg13g2_a21oi_1 _17097_ (.A1(_02452_),
    .A2(net4442),
    .Y(_01259_),
    .B1(_07482_));
 sg13g2_nor2_1 _17098_ (.A(net2928),
    .B(net4440),
    .Y(_07483_));
 sg13g2_a21oi_1 _17099_ (.A1(net5201),
    .A2(net4440),
    .Y(_01260_),
    .B1(_07483_));
 sg13g2_nor2_1 _17100_ (.A(net2975),
    .B(net4444),
    .Y(_07484_));
 sg13g2_a21oi_1 _17101_ (.A1(net5219),
    .A2(net4444),
    .Y(_01261_),
    .B1(_07484_));
 sg13g2_nor2_1 _17102_ (.A(net2902),
    .B(net4440),
    .Y(_07485_));
 sg13g2_a21oi_1 _17103_ (.A1(net5213),
    .A2(net4440),
    .Y(_01262_),
    .B1(_07485_));
 sg13g2_nor2_1 _17104_ (.A(net2892),
    .B(net4440),
    .Y(_07486_));
 sg13g2_a21oi_1 _17105_ (.A1(_02427_),
    .A2(net4440),
    .Y(_01263_),
    .B1(_07486_));
 sg13g2_nor2_1 _17106_ (.A(net2965),
    .B(net4436),
    .Y(_07487_));
 sg13g2_a21oi_1 _17107_ (.A1(_02430_),
    .A2(net4435),
    .Y(_01264_),
    .B1(_07487_));
 sg13g2_nor2_1 _17108_ (.A(net2983),
    .B(net4436),
    .Y(_07488_));
 sg13g2_a21oi_1 _17109_ (.A1(_02432_),
    .A2(net4436),
    .Y(_01265_),
    .B1(_07488_));
 sg13g2_nor2_1 _17110_ (.A(net2998),
    .B(net4435),
    .Y(_07489_));
 sg13g2_a21oi_1 _17111_ (.A1(_02434_),
    .A2(net4435),
    .Y(_01266_),
    .B1(_07489_));
 sg13g2_nor2_1 _17112_ (.A(net2925),
    .B(net4436),
    .Y(_07490_));
 sg13g2_a21oi_1 _17113_ (.A1(_02437_),
    .A2(net4436),
    .Y(_01267_),
    .B1(_07490_));
 sg13g2_nor2_1 _17114_ (.A(net2823),
    .B(net4436),
    .Y(_07491_));
 sg13g2_a21oi_1 _17115_ (.A1(_02439_),
    .A2(net4436),
    .Y(_01268_),
    .B1(_07491_));
 sg13g2_nor2_1 _17116_ (.A(net2934),
    .B(net4441),
    .Y(_07492_));
 sg13g2_a21oi_1 _17117_ (.A1(_02440_),
    .A2(net4441),
    .Y(_01269_),
    .B1(_07492_));
 sg13g2_nor2_1 _17118_ (.A(net3006),
    .B(net4435),
    .Y(_07493_));
 sg13g2_a21oi_1 _17119_ (.A1(_02443_),
    .A2(net4435),
    .Y(_01270_),
    .B1(_07493_));
 sg13g2_nor2_1 _17120_ (.A(net2939),
    .B(net4435),
    .Y(_07494_));
 sg13g2_a21oi_1 _17121_ (.A1(_02444_),
    .A2(net4435),
    .Y(_01271_),
    .B1(_07494_));
 sg13g2_nand2_1 _17122_ (.Y(_07495_),
    .A(net4392),
    .B(_07454_));
 sg13g2_o21ai_1 _17123_ (.B1(net5383),
    .Y(_07496_),
    .A1(_06015_),
    .A2(net4338));
 sg13g2_a21oi_1 _17124_ (.A1(_02332_),
    .A2(net4338),
    .Y(_01272_),
    .B1(_07496_));
 sg13g2_o21ai_1 _17125_ (.B1(net5383),
    .Y(_07497_),
    .A1(_06019_),
    .A2(net4338));
 sg13g2_a21oi_1 _17126_ (.A1(_02331_),
    .A2(net4338),
    .Y(_01273_),
    .B1(_07497_));
 sg13g2_o21ai_1 _17127_ (.B1(net5382),
    .Y(_07498_),
    .A1(_06023_),
    .A2(net4337));
 sg13g2_a21oi_1 _17128_ (.A1(_02330_),
    .A2(net4338),
    .Y(_01274_),
    .B1(_07498_));
 sg13g2_o21ai_1 _17129_ (.B1(net5382),
    .Y(_07499_),
    .A1(_06027_),
    .A2(net4338));
 sg13g2_a21oi_1 _17130_ (.A1(_02329_),
    .A2(_07495_),
    .Y(_01275_),
    .B1(_07499_));
 sg13g2_o21ai_1 _17131_ (.B1(net5381),
    .Y(_07500_),
    .A1(_06031_),
    .A2(net4337));
 sg13g2_a21oi_1 _17132_ (.A1(_02328_),
    .A2(net4337),
    .Y(_01276_),
    .B1(_07500_));
 sg13g2_o21ai_1 _17133_ (.B1(net5381),
    .Y(_07501_),
    .A1(_06035_),
    .A2(net4337));
 sg13g2_a21oi_1 _17134_ (.A1(_02327_),
    .A2(net4338),
    .Y(_01277_),
    .B1(_07501_));
 sg13g2_o21ai_1 _17135_ (.B1(net5381),
    .Y(_07502_),
    .A1(_06039_),
    .A2(net4337));
 sg13g2_a21oi_1 _17136_ (.A1(_02326_),
    .A2(net4337),
    .Y(_01278_),
    .B1(_07502_));
 sg13g2_o21ai_1 _17137_ (.B1(net5381),
    .Y(_07503_),
    .A1(_05716_),
    .A2(net4337));
 sg13g2_a21oi_1 _17138_ (.A1(_02325_),
    .A2(net4337),
    .Y(_01279_),
    .B1(_07503_));
 sg13g2_nand2_1 _17139_ (.Y(_07504_),
    .A(net4320),
    .B(_05459_));
 sg13g2_nand2_1 _17140_ (.Y(_07505_),
    .A(net1913),
    .B(net4096));
 sg13g2_o21ai_1 _17141_ (.B1(_07505_),
    .Y(_01280_),
    .A1(net4853),
    .A2(net4095));
 sg13g2_nand2_1 _17142_ (.Y(_07506_),
    .A(net1996),
    .B(net4096));
 sg13g2_o21ai_1 _17143_ (.B1(_07506_),
    .Y(_01281_),
    .A1(net4848),
    .A2(net4096));
 sg13g2_nand2_1 _17144_ (.Y(_07507_),
    .A(net1801),
    .B(net4095));
 sg13g2_o21ai_1 _17145_ (.B1(_07507_),
    .Y(_01282_),
    .A1(net4842),
    .A2(net4095));
 sg13g2_nand2_1 _17146_ (.Y(_07508_),
    .A(net1908),
    .B(net4095));
 sg13g2_o21ai_1 _17147_ (.B1(_07508_),
    .Y(_01283_),
    .A1(net4837),
    .A2(net4095));
 sg13g2_nand2_1 _17148_ (.Y(_07509_),
    .A(net2050),
    .B(net4095));
 sg13g2_o21ai_1 _17149_ (.B1(_07509_),
    .Y(_01284_),
    .A1(net4832),
    .A2(net4095));
 sg13g2_nand2_1 _17150_ (.Y(_07510_),
    .A(net1988),
    .B(net4096));
 sg13g2_o21ai_1 _17151_ (.B1(_07510_),
    .Y(_01285_),
    .A1(net4825),
    .A2(net4096));
 sg13g2_nand2_1 _17152_ (.Y(_07511_),
    .A(net1720),
    .B(_07504_));
 sg13g2_o21ai_1 _17153_ (.B1(_07511_),
    .Y(_01286_),
    .A1(net4820),
    .A2(net4095));
 sg13g2_nand2_1 _17154_ (.Y(_07512_),
    .A(net1701),
    .B(net4096));
 sg13g2_o21ai_1 _17155_ (.B1(_07512_),
    .Y(_01287_),
    .A1(net4815),
    .A2(net4096));
 sg13g2_nor2b_1 _17156_ (.A(net4333),
    .B_N(_05108_),
    .Y(_07513_));
 sg13g2_nor2_1 _17157_ (.A(net2270),
    .B(net4093),
    .Y(_07514_));
 sg13g2_a21oi_1 _17158_ (.A1(net5139),
    .A2(net4093),
    .Y(_01288_),
    .B1(_07514_));
 sg13g2_nor2_1 _17159_ (.A(net2602),
    .B(net4093),
    .Y(_07515_));
 sg13g2_a21oi_1 _17160_ (.A1(net4994),
    .A2(net4093),
    .Y(_01289_),
    .B1(_07515_));
 sg13g2_nor2_1 _17161_ (.A(net2559),
    .B(net4094),
    .Y(_07516_));
 sg13g2_a21oi_1 _17162_ (.A1(net5134),
    .A2(_07513_),
    .Y(_01290_),
    .B1(_07516_));
 sg13g2_nor2_1 _17163_ (.A(net2247),
    .B(net4094),
    .Y(_07517_));
 sg13g2_a21oi_1 _17164_ (.A1(net4991),
    .A2(net4094),
    .Y(_01291_),
    .B1(_07517_));
 sg13g2_nor2_1 _17165_ (.A(net2212),
    .B(net4094),
    .Y(_07518_));
 sg13g2_a21oi_1 _17166_ (.A1(net5125),
    .A2(net4094),
    .Y(_01292_),
    .B1(_07518_));
 sg13g2_nor2_1 _17167_ (.A(net2276),
    .B(net4093),
    .Y(_07519_));
 sg13g2_a21oi_1 _17168_ (.A1(net4985),
    .A2(net4093),
    .Y(_01293_),
    .B1(_07519_));
 sg13g2_nor2_1 _17169_ (.A(net2603),
    .B(net4094),
    .Y(_07520_));
 sg13g2_a21oi_1 _17170_ (.A1(net5120),
    .A2(net4094),
    .Y(_01294_),
    .B1(_07520_));
 sg13g2_nor2_1 _17171_ (.A(net2543),
    .B(net4093),
    .Y(_07521_));
 sg13g2_a21oi_1 _17172_ (.A1(net4982),
    .A2(net4093),
    .Y(_01295_),
    .B1(_07521_));
 sg13g2_nor2b_1 _17173_ (.A(net4331),
    .B_N(_05459_),
    .Y(_07522_));
 sg13g2_nor2_1 _17174_ (.A(net2403),
    .B(net4092),
    .Y(_07523_));
 sg13g2_a21oi_1 _17175_ (.A1(net5137),
    .A2(net4092),
    .Y(_01296_),
    .B1(_07523_));
 sg13g2_nor2_1 _17176_ (.A(net2778),
    .B(net4092),
    .Y(_07524_));
 sg13g2_a21oi_1 _17177_ (.A1(net4993),
    .A2(net4092),
    .Y(_01297_),
    .B1(_07524_));
 sg13g2_nor2_1 _17178_ (.A(net2665),
    .B(net4091),
    .Y(_07525_));
 sg13g2_a21oi_1 _17179_ (.A1(net5130),
    .A2(net4091),
    .Y(_01298_),
    .B1(_07525_));
 sg13g2_nor2_1 _17180_ (.A(net2621),
    .B(net4092),
    .Y(_07526_));
 sg13g2_a21oi_1 _17181_ (.A1(net4989),
    .A2(net4092),
    .Y(_01299_),
    .B1(_07526_));
 sg13g2_nor2_1 _17182_ (.A(net2693),
    .B(net4091),
    .Y(_07527_));
 sg13g2_a21oi_1 _17183_ (.A1(net5125),
    .A2(net4091),
    .Y(_01300_),
    .B1(_07527_));
 sg13g2_nor2_1 _17184_ (.A(net2770),
    .B(net4092),
    .Y(_07528_));
 sg13g2_a21oi_1 _17185_ (.A1(net4983),
    .A2(net4092),
    .Y(_01301_),
    .B1(_07528_));
 sg13g2_nor2_1 _17186_ (.A(net2512),
    .B(net4091),
    .Y(_07529_));
 sg13g2_a21oi_1 _17187_ (.A1(net5121),
    .A2(net4091),
    .Y(_01302_),
    .B1(_07529_));
 sg13g2_nor2_1 _17188_ (.A(net2729),
    .B(net4091),
    .Y(_07530_));
 sg13g2_a21oi_1 _17189_ (.A1(net4978),
    .A2(net4091),
    .Y(_01303_),
    .B1(_07530_));
 sg13g2_nor2b_1 _17190_ (.A(net4316),
    .B_N(_05155_),
    .Y(_07531_));
 sg13g2_nor2_1 _17191_ (.A(net2849),
    .B(net4088),
    .Y(_07532_));
 sg13g2_a21oi_1 _17192_ (.A1(net5020),
    .A2(net4088),
    .Y(_01304_),
    .B1(_07532_));
 sg13g2_nor2_1 _17193_ (.A(net2308),
    .B(net4088),
    .Y(_07533_));
 sg13g2_a21oi_1 _17194_ (.A1(net4810),
    .A2(net4088),
    .Y(_01305_),
    .B1(_07533_));
 sg13g2_nor2_1 _17195_ (.A(net2709),
    .B(net4090),
    .Y(_07534_));
 sg13g2_a21oi_1 _17196_ (.A1(net5016),
    .A2(net4090),
    .Y(_01306_),
    .B1(_07534_));
 sg13g2_nor2_1 _17197_ (.A(net2600),
    .B(net4089),
    .Y(_07535_));
 sg13g2_a21oi_1 _17198_ (.A1(net4806),
    .A2(net4089),
    .Y(_01307_),
    .B1(_07535_));
 sg13g2_nor2_1 _17199_ (.A(net2160),
    .B(net4088),
    .Y(_07536_));
 sg13g2_a21oi_1 _17200_ (.A1(net5010),
    .A2(net4088),
    .Y(_01308_),
    .B1(_07536_));
 sg13g2_nor2_1 _17201_ (.A(net2619),
    .B(net4088),
    .Y(_07537_));
 sg13g2_a21oi_1 _17202_ (.A1(net4800),
    .A2(net4088),
    .Y(_01309_),
    .B1(_07537_));
 sg13g2_nor2_1 _17203_ (.A(net2283),
    .B(net4090),
    .Y(_07538_));
 sg13g2_a21oi_1 _17204_ (.A1(net5009),
    .A2(net4090),
    .Y(_01310_),
    .B1(_07538_));
 sg13g2_nor2_1 _17205_ (.A(net2501),
    .B(net4089),
    .Y(_07539_));
 sg13g2_a21oi_1 _17206_ (.A1(net4797),
    .A2(net4089),
    .Y(_01311_),
    .B1(_07539_));
 sg13g2_a21oi_1 _17207_ (.A1(_02710_),
    .A2(_04896_),
    .Y(_07540_),
    .B1(_02712_));
 sg13g2_a21oi_1 _17208_ (.A1(net5147),
    .A2(_04895_),
    .Y(_07541_),
    .B1(_06109_));
 sg13g2_a21oi_1 _17209_ (.A1(_06359_),
    .A2(_07541_),
    .Y(_07542_),
    .B1(_07540_));
 sg13g2_nand2_1 _17210_ (.Y(_07543_),
    .A(net4789),
    .B(_07542_));
 sg13g2_nor2_1 _17211_ (.A(net4714),
    .B(_06220_),
    .Y(_07544_));
 sg13g2_o21ai_1 _17212_ (.B1(_07542_),
    .Y(_07545_),
    .A1(net4789),
    .A2(_07544_));
 sg13g2_nand2_1 _17213_ (.Y(_07546_),
    .A(net3364),
    .B(net4350));
 sg13g2_nor2_1 _17214_ (.A(_06083_),
    .B(net4336),
    .Y(_07547_));
 sg13g2_or2_2 _17215_ (.X(_07548_),
    .B(_07547_),
    .A(net4351));
 sg13g2_nor2_2 _17216_ (.A(_06082_),
    .B(_06085_),
    .Y(_07549_));
 sg13g2_xnor2_1 _17217_ (.Y(_07550_),
    .A(_02401_),
    .B(_07549_));
 sg13g2_o21ai_1 _17218_ (.B1(_07546_),
    .Y(_01312_),
    .A1(_07548_),
    .A2(_07550_));
 sg13g2_nand2_1 _17219_ (.Y(_07551_),
    .A(\m_sys.m_bootloader.r_byte_cnt[0] ),
    .B(\m_sys.m_bootloader.r_byte_cnt[1] ));
 sg13g2_xnor2_1 _17220_ (.Y(_07552_),
    .A(\m_sys.m_bootloader.r_byte_cnt[0] ),
    .B(\m_sys.m_bootloader.r_byte_cnt[1] ));
 sg13g2_inv_1 _17221_ (.Y(_07553_),
    .A(_07552_));
 sg13g2_nand3_1 _17222_ (.B(net4336),
    .C(_07553_),
    .A(net5003),
    .Y(_07554_));
 sg13g2_nor2_2 _17223_ (.A(net4713),
    .B(_06091_),
    .Y(_07555_));
 sg13g2_a22oi_1 _17224_ (.Y(_07556_),
    .B1(_07553_),
    .B2(_07555_),
    .A2(net4714),
    .A1(\m_sys.m_bootloader.r_byte_cnt[1] ));
 sg13g2_or2_1 _17225_ (.X(_07557_),
    .B(_07556_),
    .A(net5002));
 sg13g2_nand3_1 _17226_ (.B(_07554_),
    .C(_07557_),
    .A(_06081_),
    .Y(_07558_));
 sg13g2_a21oi_1 _17227_ (.A1(net4792),
    .A2(_07556_),
    .Y(_07559_),
    .B1(net4352));
 sg13g2_a22oi_1 _17228_ (.Y(_07560_),
    .B1(_07558_),
    .B2(_07559_),
    .A2(_07545_),
    .A1(net3417));
 sg13g2_inv_1 _17229_ (.Y(_01313_),
    .A(_07560_));
 sg13g2_nor2_1 _17230_ (.A(_00028_),
    .B(_07551_),
    .Y(_07561_));
 sg13g2_xnor2_1 _17231_ (.Y(_07562_),
    .A(_00028_),
    .B(_07551_));
 sg13g2_inv_1 _17232_ (.Y(_07563_),
    .A(_07562_));
 sg13g2_nand3_1 _17233_ (.B(_06198_),
    .C(_07563_),
    .A(net5003),
    .Y(_07564_));
 sg13g2_a22oi_1 _17234_ (.Y(_07565_),
    .B1(_07555_),
    .B2(_07563_),
    .A2(net4714),
    .A1(net3170));
 sg13g2_or2_1 _17235_ (.X(_07566_),
    .B(_07565_),
    .A(net5003));
 sg13g2_nand3_1 _17236_ (.B(_07564_),
    .C(_07566_),
    .A(_06081_),
    .Y(_07567_));
 sg13g2_a21oi_1 _17237_ (.A1(net4791),
    .A2(_07565_),
    .Y(_07568_),
    .B1(net4351));
 sg13g2_a22oi_1 _17238_ (.Y(_07569_),
    .B1(_07567_),
    .B2(_07568_),
    .A2(net4349),
    .A1(net3170));
 sg13g2_inv_1 _17239_ (.Y(_01314_),
    .A(_07569_));
 sg13g2_xnor2_1 _17240_ (.Y(_07570_),
    .A(_00029_),
    .B(_07561_));
 sg13g2_nand4_1 _17241_ (.B(_06128_),
    .C(net4336),
    .A(net5004),
    .Y(_07571_),
    .D(_07570_));
 sg13g2_a22oi_1 _17242_ (.Y(_07572_),
    .B1(_07555_),
    .B2(_07570_),
    .A2(net4713),
    .A1(\m_sys.m_bootloader.r_byte_cnt[3] ));
 sg13g2_nor2_1 _17243_ (.A(_06082_),
    .B(_07572_),
    .Y(_07573_));
 sg13g2_nor2_1 _17244_ (.A(_06227_),
    .B(_07573_),
    .Y(_07574_));
 sg13g2_a221oi_1 _17245_ (.B2(_07571_),
    .C1(net4351),
    .B1(_07574_),
    .A1(_06227_),
    .Y(_07575_),
    .A2(_07572_));
 sg13g2_a21oi_1 _17246_ (.A1(net3172),
    .A2(net4349),
    .Y(_07576_),
    .B1(_07575_));
 sg13g2_inv_1 _17247_ (.Y(_01315_),
    .A(_07576_));
 sg13g2_nand4_1 _17248_ (.B(\m_sys.m_bootloader.r_byte_cnt[1] ),
    .C(\m_sys.m_bootloader.r_byte_cnt[2] ),
    .A(\m_sys.m_bootloader.r_byte_cnt[0] ),
    .Y(_07577_),
    .D(\m_sys.m_bootloader.r_byte_cnt[3] ));
 sg13g2_nor2_1 _17249_ (.A(_00030_),
    .B(_07577_),
    .Y(_07578_));
 sg13g2_xnor2_1 _17250_ (.Y(_07579_),
    .A(_00030_),
    .B(_07577_));
 sg13g2_inv_1 _17251_ (.Y(_07580_),
    .A(_07579_));
 sg13g2_nand3_1 _17252_ (.B(net4336),
    .C(_07580_),
    .A(net5003),
    .Y(_07581_));
 sg13g2_a22oi_1 _17253_ (.Y(_07582_),
    .B1(_07555_),
    .B2(_07580_),
    .A2(net4713),
    .A1(net3079));
 sg13g2_or2_1 _17254_ (.X(_07583_),
    .B(_07582_),
    .A(net5002));
 sg13g2_nand3_1 _17255_ (.B(_07581_),
    .C(_07583_),
    .A(_06081_),
    .Y(_07584_));
 sg13g2_a21oi_1 _17256_ (.A1(net4791),
    .A2(_07582_),
    .Y(_07585_),
    .B1(net4351));
 sg13g2_a22oi_1 _17257_ (.Y(_07586_),
    .B1(_07584_),
    .B2(_07585_),
    .A2(net4349),
    .A1(net3079));
 sg13g2_inv_1 _17258_ (.Y(_01316_),
    .A(_07586_));
 sg13g2_xnor2_1 _17259_ (.Y(_07587_),
    .A(_00031_),
    .B(_07578_));
 sg13g2_nand3_1 _17260_ (.B(net4336),
    .C(_07587_),
    .A(net5002),
    .Y(_07588_));
 sg13g2_a22oi_1 _17261_ (.Y(_07589_),
    .B1(_07555_),
    .B2(_07587_),
    .A2(net4713),
    .A1(\m_sys.m_bootloader.r_byte_cnt[5] ));
 sg13g2_a21o_1 _17262_ (.A2(_07589_),
    .A1(_06081_),
    .B1(_06082_),
    .X(_07590_));
 sg13g2_a221oi_1 _17263_ (.B2(_07588_),
    .C1(net4351),
    .B1(_07590_),
    .A1(net4791),
    .Y(_07591_),
    .A2(_07589_));
 sg13g2_a21o_1 _17264_ (.A2(net4349),
    .A1(net3112),
    .B1(_07591_),
    .X(_01317_));
 sg13g2_nand2_1 _17265_ (.Y(_07592_),
    .A(net2880),
    .B(net4349));
 sg13g2_nand2_1 _17266_ (.Y(_07593_),
    .A(\m_sys.m_bootloader.r_byte_cnt[4] ),
    .B(\m_sys.m_bootloader.r_byte_cnt[5] ));
 sg13g2_nor2_1 _17267_ (.A(_07577_),
    .B(_07593_),
    .Y(_07594_));
 sg13g2_nor3_1 _17268_ (.A(_00032_),
    .B(_07577_),
    .C(_07593_),
    .Y(_07595_));
 sg13g2_xnor2_1 _17269_ (.Y(_07596_),
    .A(_00032_),
    .B(_07594_));
 sg13g2_nand3_1 _17270_ (.B(net4336),
    .C(_07596_),
    .A(net5002),
    .Y(_07597_));
 sg13g2_a22oi_1 _17271_ (.Y(_07598_),
    .B1(_07555_),
    .B2(_07596_),
    .A2(net4713),
    .A1(net2880));
 sg13g2_o21ai_1 _17272_ (.B1(_07597_),
    .Y(_07599_),
    .A1(net5002),
    .A2(_07598_));
 sg13g2_a21oi_1 _17273_ (.A1(net4791),
    .A2(_07598_),
    .Y(_07600_),
    .B1(net4351));
 sg13g2_o21ai_1 _17274_ (.B1(_07600_),
    .Y(_07601_),
    .A1(net4791),
    .A2(_07599_));
 sg13g2_nand2_1 _17275_ (.Y(_01318_),
    .A(_07592_),
    .B(_07601_));
 sg13g2_xnor2_1 _17276_ (.Y(_07602_),
    .A(_00034_),
    .B(_07595_));
 sg13g2_nand3_1 _17277_ (.B(net4336),
    .C(_07602_),
    .A(net5002),
    .Y(_07603_));
 sg13g2_a22oi_1 _17278_ (.Y(_07604_),
    .B1(_07555_),
    .B2(_07602_),
    .A2(net4713),
    .A1(\m_sys.m_bootloader.r_byte_cnt[7] ));
 sg13g2_a21o_1 _17279_ (.A2(_07604_),
    .A1(_06081_),
    .B1(_06082_),
    .X(_07605_));
 sg13g2_a221oi_1 _17280_ (.B2(_07603_),
    .C1(net4351),
    .B1(_07605_),
    .A1(net4791),
    .Y(_07606_),
    .A2(_07604_));
 sg13g2_a21o_1 _17281_ (.A2(net4349),
    .A1(net3135),
    .B1(_07606_),
    .X(_01319_));
 sg13g2_nand2_1 _17282_ (.Y(_07607_),
    .A(net3046),
    .B(net4349));
 sg13g2_nand3_1 _17283_ (.B(\m_sys.m_bootloader.r_byte_cnt[7] ),
    .C(_07594_),
    .A(\m_sys.m_bootloader.r_byte_cnt[6] ),
    .Y(_07608_));
 sg13g2_nor2_1 _17284_ (.A(_00035_),
    .B(_07608_),
    .Y(_07609_));
 sg13g2_xor2_1 _17285_ (.B(_07608_),
    .A(_00035_),
    .X(_07610_));
 sg13g2_nand3_1 _17286_ (.B(net4336),
    .C(_07610_),
    .A(net5002),
    .Y(_07611_));
 sg13g2_a22oi_1 _17287_ (.Y(_07612_),
    .B1(_07555_),
    .B2(_07610_),
    .A2(net4713),
    .A1(\m_sys.m_bootloader.r_byte_cnt[8] ));
 sg13g2_o21ai_1 _17288_ (.B1(_07611_),
    .Y(_07613_),
    .A1(net5002),
    .A2(_07612_));
 sg13g2_a21oi_1 _17289_ (.A1(net4791),
    .A2(_07612_),
    .Y(_07614_),
    .B1(net4351));
 sg13g2_o21ai_1 _17290_ (.B1(_07614_),
    .Y(_07615_),
    .A1(net4791),
    .A2(_07613_));
 sg13g2_nand2_1 _17291_ (.Y(_01320_),
    .A(_07607_),
    .B(_07615_));
 sg13g2_o21ai_1 _17292_ (.B1(_06083_),
    .Y(_07616_),
    .A1(net4713),
    .A2(_06091_));
 sg13g2_xnor2_1 _17293_ (.Y(_07617_),
    .A(_00036_),
    .B(_07609_));
 sg13g2_a22oi_1 _17294_ (.Y(_07618_),
    .B1(_07616_),
    .B2(_07617_),
    .A2(_07549_),
    .A1(net3022));
 sg13g2_nand2_1 _17295_ (.Y(_07619_),
    .A(net3022),
    .B(net4349));
 sg13g2_o21ai_1 _17296_ (.B1(_07619_),
    .Y(_01321_),
    .A1(_07548_),
    .A2(_07618_));
 sg13g2_nand2_1 _17297_ (.Y(_07620_),
    .A(net3061),
    .B(net4350));
 sg13g2_nor2b_2 _17298_ (.A(_07547_),
    .B_N(_07616_),
    .Y(_07621_));
 sg13g2_nand2_1 _17299_ (.Y(_07622_),
    .A(\m_sys.m_bootloader.r_byte_cnt[8] ),
    .B(\m_sys.m_bootloader.r_byte_cnt[9] ));
 sg13g2_nor2_1 _17300_ (.A(_07608_),
    .B(_07622_),
    .Y(_07623_));
 sg13g2_nor3_1 _17301_ (.A(_00037_),
    .B(_07608_),
    .C(_07622_),
    .Y(_07624_));
 sg13g2_xnor2_1 _17302_ (.Y(_07625_),
    .A(_00037_),
    .B(_07623_));
 sg13g2_a22oi_1 _17303_ (.Y(_07626_),
    .B1(_07621_),
    .B2(_07625_),
    .A2(_07549_),
    .A1(net3061));
 sg13g2_o21ai_1 _17304_ (.B1(_07620_),
    .Y(_01322_),
    .A1(net4352),
    .A2(_07626_));
 sg13g2_xnor2_1 _17305_ (.Y(_07627_),
    .A(_00038_),
    .B(_07624_));
 sg13g2_a22oi_1 _17306_ (.Y(_07628_),
    .B1(_07616_),
    .B2(_07627_),
    .A2(_07549_),
    .A1(net3001));
 sg13g2_nand2_1 _17307_ (.Y(_07629_),
    .A(net3001),
    .B(net4350));
 sg13g2_o21ai_1 _17308_ (.B1(_07629_),
    .Y(_01323_),
    .A1(_07548_),
    .A2(_07628_));
 sg13g2_nand3_1 _17309_ (.B(\m_sys.m_bootloader.r_byte_cnt[11] ),
    .C(_07623_),
    .A(\m_sys.m_bootloader.r_byte_cnt[10] ),
    .Y(_07630_));
 sg13g2_inv_1 _17310_ (.Y(_07631_),
    .A(_07630_));
 sg13g2_nor2_1 _17311_ (.A(_00039_),
    .B(_07630_),
    .Y(_07632_));
 sg13g2_xor2_1 _17312_ (.B(_07630_),
    .A(_00039_),
    .X(_07633_));
 sg13g2_a22oi_1 _17313_ (.Y(_07634_),
    .B1(_07616_),
    .B2(_07633_),
    .A2(_07549_),
    .A1(net2921));
 sg13g2_nand2_1 _17314_ (.Y(_07635_),
    .A(net2921),
    .B(net4350));
 sg13g2_o21ai_1 _17315_ (.B1(_07635_),
    .Y(_01324_),
    .A1(_07548_),
    .A2(_07634_));
 sg13g2_nand2_1 _17316_ (.Y(_07636_),
    .A(net2833),
    .B(net4350));
 sg13g2_xnor2_1 _17317_ (.Y(_07637_),
    .A(_00040_),
    .B(_07632_));
 sg13g2_a22oi_1 _17318_ (.Y(_07638_),
    .B1(_07621_),
    .B2(_07637_),
    .A2(_07549_),
    .A1(net2833));
 sg13g2_o21ai_1 _17319_ (.B1(_07636_),
    .Y(_01325_),
    .A1(net4352),
    .A2(_07638_));
 sg13g2_nand2_1 _17320_ (.Y(_07639_),
    .A(net2451),
    .B(net4350));
 sg13g2_nand3_1 _17321_ (.B(\m_sys.m_bootloader.r_byte_cnt[13] ),
    .C(_07631_),
    .A(\m_sys.m_bootloader.r_byte_cnt[12] ),
    .Y(_07640_));
 sg13g2_nor2_1 _17322_ (.A(_00041_),
    .B(_07640_),
    .Y(_07641_));
 sg13g2_xor2_1 _17323_ (.B(_07640_),
    .A(_00041_),
    .X(_07642_));
 sg13g2_a22oi_1 _17324_ (.Y(_01776_),
    .B1(_07621_),
    .B2(_07642_),
    .A2(_07549_),
    .A1(net2451));
 sg13g2_o21ai_1 _17325_ (.B1(_07639_),
    .Y(_01326_),
    .A1(net4352),
    .A2(_01776_));
 sg13g2_nand2_1 _17326_ (.Y(_01777_),
    .A(net2561),
    .B(net4350));
 sg13g2_xnor2_1 _17327_ (.Y(_01778_),
    .A(_00042_),
    .B(_07641_));
 sg13g2_a22oi_1 _17328_ (.Y(_01779_),
    .B1(_07621_),
    .B2(_01778_),
    .A2(_07549_),
    .A1(net2561));
 sg13g2_o21ai_1 _17329_ (.B1(_01777_),
    .Y(_01327_),
    .A1(net4352),
    .A2(_01779_));
 sg13g2_a21oi_2 _17330_ (.B1(net4957),
    .Y(_01780_),
    .A2(_05305_),
    .A1(net5317));
 sg13g2_a21o_2 _17331_ (.A2(_05305_),
    .A1(net5317),
    .B1(net4957),
    .X(_01781_));
 sg13g2_a21oi_2 _17332_ (.B1(_03556_),
    .Y(_01782_),
    .A2(_02773_),
    .A1(net5318));
 sg13g2_nor2_1 _17333_ (.A(_00018_),
    .B(_01782_),
    .Y(_01783_));
 sg13g2_nand2b_2 _17334_ (.Y(_01784_),
    .B(_02772_),
    .A_N(net5317));
 sg13g2_nor2_1 _17335_ (.A(_00078_),
    .B(_01784_),
    .Y(_01785_));
 sg13g2_o21ai_1 _17336_ (.B1(net4706),
    .Y(_01786_),
    .A1(_01783_),
    .A2(_01785_));
 sg13g2_a21oi_1 _17337_ (.A1(_05104_),
    .A2(net4703),
    .Y(_01787_),
    .B1(net4959));
 sg13g2_a22oi_1 _17338_ (.Y(_01788_),
    .B1(_01786_),
    .B2(_01787_),
    .A2(_04864_),
    .A1(net4959));
 sg13g2_nand2_1 _17339_ (.Y(_01789_),
    .A(net4750),
    .B(_01788_));
 sg13g2_o21ai_1 _17340_ (.B1(_01789_),
    .Y(_01328_),
    .A1(_02460_),
    .A2(net4750));
 sg13g2_nand2_1 _17341_ (.Y(_01790_),
    .A(net3202),
    .B(net4756));
 sg13g2_nor2_1 _17342_ (.A(_00066_),
    .B(_01782_),
    .Y(_01791_));
 sg13g2_nor2_1 _17343_ (.A(_00065_),
    .B(_01784_),
    .Y(_01792_));
 sg13g2_o21ai_1 _17344_ (.B1(net4706),
    .Y(_01793_),
    .A1(_01791_),
    .A2(_01792_));
 sg13g2_a21oi_1 _17345_ (.A1(_02769_),
    .A2(net4704),
    .Y(_01794_),
    .B1(net4959));
 sg13g2_nand2_1 _17346_ (.Y(_01795_),
    .A(_01793_),
    .B(_01794_));
 sg13g2_o21ai_1 _17347_ (.B1(_01795_),
    .Y(_01796_),
    .A1(net4972),
    .A2(_04829_));
 sg13g2_o21ai_1 _17348_ (.B1(_01790_),
    .Y(_01329_),
    .A1(net4755),
    .A2(_01796_));
 sg13g2_or2_1 _17349_ (.X(_01797_),
    .B(_01784_),
    .A(_00067_));
 sg13g2_o21ai_1 _17350_ (.B1(_01797_),
    .Y(_01798_),
    .A1(_00068_),
    .A2(_01782_));
 sg13g2_o21ai_1 _17351_ (.B1(net4972),
    .Y(_01799_),
    .A1(_02793_),
    .A2(net4706));
 sg13g2_a21oi_2 _17352_ (.B1(_01799_),
    .Y(_01800_),
    .A2(_01798_),
    .A1(net4706));
 sg13g2_a21oi_1 _17353_ (.A1(net4960),
    .A2(_04794_),
    .Y(_01801_),
    .B1(_01800_));
 sg13g2_nand2_1 _17354_ (.Y(_01802_),
    .A(net4749),
    .B(_01801_));
 sg13g2_o21ai_1 _17355_ (.B1(_01802_),
    .Y(_01330_),
    .A1(_02463_),
    .A2(net4749));
 sg13g2_nor2_1 _17356_ (.A(_00070_),
    .B(_01782_),
    .Y(_01803_));
 sg13g2_nor2_1 _17357_ (.A(_00069_),
    .B(_01784_),
    .Y(_01804_));
 sg13g2_o21ai_1 _17358_ (.B1(net4706),
    .Y(_01805_),
    .A1(_01803_),
    .A2(_01804_));
 sg13g2_a21oi_1 _17359_ (.A1(_02803_),
    .A2(net4703),
    .Y(_01806_),
    .B1(net4959));
 sg13g2_a21oi_1 _17360_ (.A1(_01805_),
    .A2(_01806_),
    .Y(_01807_),
    .B1(net4755));
 sg13g2_o21ai_1 _17361_ (.B1(_01807_),
    .Y(_01808_),
    .A1(net4971),
    .A2(_04758_));
 sg13g2_o21ai_1 _17362_ (.B1(_01808_),
    .Y(_01331_),
    .A1(_02462_),
    .A2(net4749));
 sg13g2_or2_1 _17363_ (.X(_01809_),
    .B(_01784_),
    .A(_00071_));
 sg13g2_o21ai_1 _17364_ (.B1(_01809_),
    .Y(_01810_),
    .A1(_00016_),
    .A2(_01782_));
 sg13g2_o21ai_1 _17365_ (.B1(net4972),
    .Y(_01811_),
    .A1(_02812_),
    .A2(net4706));
 sg13g2_a21oi_2 _17366_ (.B1(_01811_),
    .Y(_01812_),
    .A2(_01810_),
    .A1(net4706));
 sg13g2_a21oi_1 _17367_ (.A1(net4960),
    .A2(_04718_),
    .Y(_01813_),
    .B1(_01812_));
 sg13g2_nand2_1 _17368_ (.Y(_01814_),
    .A(net4749),
    .B(_01813_));
 sg13g2_o21ai_1 _17369_ (.B1(_01814_),
    .Y(_01332_),
    .A1(_02466_),
    .A2(net4749));
 sg13g2_nand2_1 _17370_ (.Y(_01815_),
    .A(net4960),
    .B(_04687_));
 sg13g2_a21oi_2 _17371_ (.B1(_02782_),
    .Y(_01816_),
    .A2(_01784_),
    .A1(_02774_));
 sg13g2_nor2_2 _17372_ (.A(_03556_),
    .B(_01816_),
    .Y(_01817_));
 sg13g2_a21oi_1 _17373_ (.A1(_02822_),
    .A2(net4703),
    .Y(_01818_),
    .B1(net4963));
 sg13g2_o21ai_1 _17374_ (.B1(_01818_),
    .Y(_01819_),
    .A1(_00072_),
    .A2(_01817_));
 sg13g2_nand3_1 _17375_ (.B(_01815_),
    .C(_01819_),
    .A(net4749),
    .Y(_01820_));
 sg13g2_o21ai_1 _17376_ (.B1(_01820_),
    .Y(_01333_),
    .A1(_02465_),
    .A2(net4749));
 sg13g2_nand2_1 _17377_ (.Y(_01821_),
    .A(net4959),
    .B(_04635_));
 sg13g2_a21oi_1 _17378_ (.A1(_02830_),
    .A2(net4703),
    .Y(_01822_),
    .B1(net4965));
 sg13g2_o21ai_1 _17379_ (.B1(_01822_),
    .Y(_01823_),
    .A1(net3232),
    .A2(_01817_));
 sg13g2_a21oi_1 _17380_ (.A1(_01821_),
    .A2(_01823_),
    .Y(_01824_),
    .B1(net4755));
 sg13g2_a21oi_1 _17381_ (.A1(_02464_),
    .A2(net4755),
    .Y(_01334_),
    .B1(_01824_));
 sg13g2_or2_1 _17382_ (.X(_01825_),
    .B(_01817_),
    .A(_00074_));
 sg13g2_a21oi_1 _17383_ (.A1(_02837_),
    .A2(net4703),
    .Y(_01826_),
    .B1(net4965));
 sg13g2_a22oi_1 _17384_ (.Y(_01827_),
    .B1(_01825_),
    .B2(_01826_),
    .A2(_04603_),
    .A1(net4965));
 sg13g2_mux2_1 _17385_ (.A0(net3178),
    .A1(_01827_),
    .S(net4749),
    .X(_01335_));
 sg13g2_nand2_1 _17386_ (.Y(_01828_),
    .A(net4959),
    .B(_04564_));
 sg13g2_a21oi_1 _17387_ (.A1(_02844_),
    .A2(net4703),
    .Y(_01829_),
    .B1(net4963));
 sg13g2_o21ai_1 _17388_ (.B1(_01829_),
    .Y(_01830_),
    .A1(net1799),
    .A2(_01817_));
 sg13g2_nand3_1 _17389_ (.B(_01828_),
    .C(_01830_),
    .A(net4750),
    .Y(_01831_));
 sg13g2_o21ai_1 _17390_ (.B1(_01831_),
    .Y(_01336_),
    .A1(_02474_),
    .A2(net4748));
 sg13g2_nand2_1 _17391_ (.Y(_01832_),
    .A(net3028),
    .B(net4756));
 sg13g2_a21oi_1 _17392_ (.A1(_02851_),
    .A2(net4704),
    .Y(_01833_),
    .B1(net4965));
 sg13g2_o21ai_1 _17393_ (.B1(_01833_),
    .Y(_01834_),
    .A1(net2471),
    .A2(_01817_));
 sg13g2_o21ai_1 _17394_ (.B1(_01834_),
    .Y(_01835_),
    .A1(net4972),
    .A2(_04521_));
 sg13g2_o21ai_1 _17395_ (.B1(_01832_),
    .Y(_01337_),
    .A1(net4756),
    .A2(_01835_));
 sg13g2_nand2_1 _17396_ (.Y(_01836_),
    .A(net3019),
    .B(net4755));
 sg13g2_a21oi_1 _17397_ (.A1(_02858_),
    .A2(net4703),
    .Y(_01837_),
    .B1(net4963));
 sg13g2_o21ai_1 _17398_ (.B1(_01837_),
    .Y(_01838_),
    .A1(net1655),
    .A2(_01817_));
 sg13g2_o21ai_1 _17399_ (.B1(_01838_),
    .Y(_01839_),
    .A1(net4974),
    .A2(_04478_));
 sg13g2_o21ai_1 _17400_ (.B1(_01836_),
    .Y(_01338_),
    .A1(net4755),
    .A2(_01839_));
 sg13g2_nor2_1 _17401_ (.A(_00080_),
    .B(_03556_),
    .Y(_01840_));
 sg13g2_a21oi_1 _17402_ (.A1(net5353),
    .A2(_03556_),
    .Y(_01841_),
    .B1(_01840_));
 sg13g2_a221oi_1 _17403_ (.B2(_01840_),
    .C1(net4704),
    .B1(_01816_),
    .A1(net5353),
    .Y(_01842_),
    .A2(_03556_));
 sg13g2_o21ai_1 _17404_ (.B1(net4707),
    .Y(_01843_),
    .A1(_01817_),
    .A2(_01841_));
 sg13g2_a21oi_1 _17405_ (.A1(_02868_),
    .A2(net4703),
    .Y(_01844_),
    .B1(net4963));
 sg13g2_a221oi_1 _17406_ (.B2(_01844_),
    .C1(net4756),
    .B1(net4348),
    .A1(net4963),
    .Y(_01845_),
    .A2(_04440_));
 sg13g2_a21oi_1 _17407_ (.A1(_02471_),
    .A2(net4755),
    .Y(_01339_),
    .B1(_01845_));
 sg13g2_nor2_1 _17408_ (.A(net4974),
    .B(_04391_),
    .Y(_01846_));
 sg13g2_nand2_1 _17409_ (.Y(_01847_),
    .A(\m_sys.m_core.m_bru.io_i_s1[12] ),
    .B(net4741));
 sg13g2_a221oi_1 _17410_ (.B2(_01847_),
    .C1(net4964),
    .B1(net4379),
    .A1(_02880_),
    .Y(_01848_),
    .A2(net4704));
 sg13g2_o21ai_1 _17411_ (.B1(net4754),
    .Y(_01849_),
    .A1(_01846_),
    .A2(_01848_));
 sg13g2_o21ai_1 _17412_ (.B1(_01849_),
    .Y(_01340_),
    .A1(_02470_),
    .A2(net4754));
 sg13g2_nor2_1 _17413_ (.A(net4974),
    .B(_04355_),
    .Y(_01850_));
 sg13g2_nand2_1 _17414_ (.Y(_01851_),
    .A(net5323),
    .B(net4741));
 sg13g2_a221oi_1 _17415_ (.B2(_01851_),
    .C1(net4964),
    .B1(net4379),
    .A1(_02893_),
    .Y(_01852_),
    .A2(net4704));
 sg13g2_nor3_1 _17416_ (.A(net4760),
    .B(_01850_),
    .C(_01852_),
    .Y(_01853_));
 sg13g2_a21oi_1 _17417_ (.A1(_02469_),
    .A2(net4756),
    .Y(_01341_),
    .B1(_01853_));
 sg13g2_a21oi_1 _17418_ (.A1(\m_sys.m_core.m_bru.io_i_s1[14] ),
    .A2(net4741),
    .Y(_01854_),
    .B1(net4348));
 sg13g2_a21o_1 _17419_ (.A2(net4704),
    .A1(_02903_),
    .B1(net4966),
    .X(_01855_));
 sg13g2_a22oi_1 _17420_ (.Y(_01856_),
    .B1(_04317_),
    .B2(net5096),
    .A2(net4756),
    .A1(net3405));
 sg13g2_o21ai_1 _17421_ (.B1(_01856_),
    .Y(_01342_),
    .A1(_01854_),
    .A2(_01855_));
 sg13g2_nand2_1 _17422_ (.Y(_01857_),
    .A(net4966),
    .B(_04285_));
 sg13g2_nand2_1 _17423_ (.Y(_01858_),
    .A(net5324),
    .B(net4741));
 sg13g2_a221oi_1 _17424_ (.B2(_01858_),
    .C1(net4966),
    .B1(net4379),
    .A1(_02915_),
    .Y(_01859_),
    .A2(net4705));
 sg13g2_nor2_1 _17425_ (.A(net4757),
    .B(_01859_),
    .Y(_01860_));
 sg13g2_a22oi_1 _17426_ (.Y(_01343_),
    .B1(_01857_),
    .B2(_01860_),
    .A2(net4757),
    .A1(_02467_));
 sg13g2_nand2_1 _17427_ (.Y(_01861_),
    .A(net5325),
    .B(net4743));
 sg13g2_a221oi_1 _17428_ (.B2(_01861_),
    .C1(net4969),
    .B1(_01842_),
    .A1(_02927_),
    .Y(_01862_),
    .A2(_01781_));
 sg13g2_a21oi_1 _17429_ (.A1(net3418),
    .A2(net4759),
    .Y(_01863_),
    .B1(_01862_));
 sg13g2_o21ai_1 _17430_ (.B1(_01863_),
    .Y(_01344_),
    .A1(_03067_),
    .A2(_04242_));
 sg13g2_nor2_1 _17431_ (.A(net4976),
    .B(_04210_),
    .Y(_01864_));
 sg13g2_nand2_1 _17432_ (.Y(_01865_),
    .A(net5327),
    .B(net4743));
 sg13g2_a221oi_1 _17433_ (.B2(_01865_),
    .C1(net4969),
    .B1(_01842_),
    .A1(_02939_),
    .Y(_01866_),
    .A2(net4705));
 sg13g2_nor3_1 _17434_ (.A(net4759),
    .B(_01864_),
    .C(_01866_),
    .Y(_01867_));
 sg13g2_a21oi_1 _17435_ (.A1(_02484_),
    .A2(net4759),
    .Y(_01345_),
    .B1(_01867_));
 sg13g2_nand2_1 _17436_ (.Y(_01868_),
    .A(\m_sys.m_core.m_bru.io_i_s1[18] ),
    .B(net4743));
 sg13g2_a221oi_1 _17437_ (.B2(_01868_),
    .C1(net4969),
    .B1(net4379),
    .A1(_02951_),
    .Y(_01869_),
    .A2(net4705));
 sg13g2_nand2_1 _17438_ (.Y(_01870_),
    .A(net4969),
    .B(_04172_));
 sg13g2_o21ai_1 _17439_ (.B1(_01870_),
    .Y(_01871_),
    .A1(net5096),
    .A2(_01869_));
 sg13g2_o21ai_1 _17440_ (.B1(_01871_),
    .Y(_01346_),
    .A1(_02483_),
    .A2(net4752));
 sg13g2_nand2_1 _17441_ (.Y(_01872_),
    .A(\m_sys.m_core.m_bru.io_i_s1[19] ),
    .B(net4743));
 sg13g2_a221oi_1 _17442_ (.B2(_01872_),
    .C1(net4968),
    .B1(net4379),
    .A1(_02961_),
    .Y(_01873_),
    .A2(net4705));
 sg13g2_a21oi_1 _17443_ (.A1(net4969),
    .A2(_04137_),
    .Y(_01874_),
    .B1(_01873_));
 sg13g2_nor2_1 _17444_ (.A(net3349),
    .B(net4752),
    .Y(_01875_));
 sg13g2_a21oi_1 _17445_ (.A1(net4752),
    .A2(_01874_),
    .Y(_01347_),
    .B1(_01875_));
 sg13g2_a21oi_1 _17446_ (.A1(net5332),
    .A2(net4742),
    .Y(_01876_),
    .B1(net4348));
 sg13g2_o21ai_1 _17447_ (.B1(net4975),
    .Y(_01877_),
    .A1(_02971_),
    .A2(net4707));
 sg13g2_or2_1 _17448_ (.X(_01878_),
    .B(_01877_),
    .A(_01876_));
 sg13g2_a22oi_1 _17449_ (.Y(_01879_),
    .B1(_01878_),
    .B2(net5093),
    .A2(_04097_),
    .A1(net4968));
 sg13g2_a21o_1 _17450_ (.A2(net4758),
    .A1(net3359),
    .B1(_01879_),
    .X(_01348_));
 sg13g2_or2_1 _17451_ (.X(_01880_),
    .B(_04060_),
    .A(net4975));
 sg13g2_a21oi_1 _17452_ (.A1(net5341),
    .A2(net4742),
    .Y(_01881_),
    .B1(net4348));
 sg13g2_o21ai_1 _17453_ (.B1(net4975),
    .Y(_01882_),
    .A1(_02978_),
    .A2(net4707));
 sg13g2_o21ai_1 _17454_ (.B1(_01880_),
    .Y(_01883_),
    .A1(_01881_),
    .A2(_01882_));
 sg13g2_mux2_1 _17455_ (.A0(net3304),
    .A1(_01883_),
    .S(net4751),
    .X(_01349_));
 sg13g2_a21oi_1 _17456_ (.A1(net5352),
    .A2(net4742),
    .Y(_01884_),
    .B1(net4348));
 sg13g2_o21ai_1 _17457_ (.B1(net4975),
    .Y(_01885_),
    .A1(_02986_),
    .A2(net4707));
 sg13g2_or2_1 _17458_ (.X(_01886_),
    .B(_01885_),
    .A(_01884_));
 sg13g2_a22oi_1 _17459_ (.Y(_01887_),
    .B1(_01886_),
    .B2(net5093),
    .A2(_04021_),
    .A1(net4968));
 sg13g2_a21o_1 _17460_ (.A2(net4758),
    .A1(net3262),
    .B1(_01887_),
    .X(_01350_));
 sg13g2_a21o_1 _17461_ (.A2(net4742),
    .A1(\m_sys.m_core.m_bru.io_i_s1[23] ),
    .B1(_01843_),
    .X(_01888_));
 sg13g2_a21oi_1 _17462_ (.A1(_02996_),
    .A2(net4705),
    .Y(_01889_),
    .B1(net4968));
 sg13g2_a221oi_1 _17463_ (.B2(_01889_),
    .C1(net4758),
    .B1(_01888_),
    .A1(net4968),
    .Y(_01890_),
    .A2(_03986_));
 sg13g2_a21oi_1 _17464_ (.A1(_02481_),
    .A2(net4758),
    .Y(_01351_),
    .B1(_01890_));
 sg13g2_nor2_1 _17465_ (.A(net4975),
    .B(_03943_),
    .Y(_01891_));
 sg13g2_nand2_1 _17466_ (.Y(_01892_),
    .A(\m_sys.m_core.m_bru.io_i_s1[24] ),
    .B(net4742));
 sg13g2_o21ai_1 _17467_ (.B1(net4975),
    .Y(_01893_),
    .A1(_03003_),
    .A2(_01780_));
 sg13g2_a21oi_1 _17468_ (.A1(net4379),
    .A2(_01892_),
    .Y(_01894_),
    .B1(_01893_));
 sg13g2_nor3_1 _17469_ (.A(net4758),
    .B(_01891_),
    .C(_01894_),
    .Y(_01895_));
 sg13g2_a21oi_1 _17470_ (.A1(_02480_),
    .A2(net4759),
    .Y(_01352_),
    .B1(_01895_));
 sg13g2_nand2_1 _17471_ (.Y(_01896_),
    .A(\m_sys.m_core.m_bru.io_i_s1[25] ),
    .B(net4742));
 sg13g2_a221oi_1 _17472_ (.B2(_01896_),
    .C1(net4967),
    .B1(net4379),
    .A1(_03013_),
    .Y(_01897_),
    .A2(net4705));
 sg13g2_a21oi_1 _17473_ (.A1(net4967),
    .A2(_03903_),
    .Y(_01898_),
    .B1(_01897_));
 sg13g2_nor2_1 _17474_ (.A(net3275),
    .B(net4751),
    .Y(_01899_));
 sg13g2_a21oi_1 _17475_ (.A1(net4751),
    .A2(_01898_),
    .Y(_01353_),
    .B1(_01899_));
 sg13g2_a21oi_1 _17476_ (.A1(\m_sys.m_core.m_bru.io_i_s1[26] ),
    .A2(net4742),
    .Y(_01900_),
    .B1(net4348));
 sg13g2_o21ai_1 _17477_ (.B1(net4977),
    .Y(_01901_),
    .A1(_03021_),
    .A2(net4707));
 sg13g2_or2_1 _17478_ (.X(_01902_),
    .B(_01901_),
    .A(_01900_));
 sg13g2_a22oi_1 _17479_ (.Y(_01903_),
    .B1(_01902_),
    .B2(net5093),
    .A2(_03860_),
    .A1(net4966));
 sg13g2_a21o_1 _17480_ (.A2(net4758),
    .A1(net3043),
    .B1(_01903_),
    .X(_01354_));
 sg13g2_a21o_1 _17481_ (.A2(net4742),
    .A1(\m_sys.m_core.m_bru.io_i_s1[27] ),
    .B1(_01843_),
    .X(_01904_));
 sg13g2_a21oi_1 _17482_ (.A1(_03031_),
    .A2(net4705),
    .Y(_01905_),
    .B1(net4968));
 sg13g2_a221oi_1 _17483_ (.B2(_01905_),
    .C1(net4759),
    .B1(_01904_),
    .A1(net4968),
    .Y(_01906_),
    .A2(_03818_));
 sg13g2_a21oi_1 _17484_ (.A1(_02478_),
    .A2(net4758),
    .Y(_01355_),
    .B1(_01906_));
 sg13g2_a21oi_1 _17485_ (.A1(\m_sys.m_core.m_bru.io_i_s1[28] ),
    .A2(net4741),
    .Y(_01907_),
    .B1(_01843_));
 sg13g2_o21ai_1 _17486_ (.B1(net4977),
    .Y(_01908_),
    .A1(_03039_),
    .A2(net4707));
 sg13g2_or2_1 _17487_ (.X(_01909_),
    .B(_01908_),
    .A(_01907_));
 sg13g2_a22oi_1 _17488_ (.Y(_01910_),
    .B1(_01909_),
    .B2(_03067_),
    .A2(_03769_),
    .A1(net4966));
 sg13g2_a21o_1 _17489_ (.A2(net4757),
    .A1(net3192),
    .B1(_01910_),
    .X(_01356_));
 sg13g2_nor2_1 _17490_ (.A(net4977),
    .B(_03715_),
    .Y(_01911_));
 sg13g2_nand2_1 _17491_ (.Y(_01912_),
    .A(\m_sys.m_core.m_bru.io_i_s1[29] ),
    .B(net4741));
 sg13g2_a221oi_1 _17492_ (.B2(_01912_),
    .C1(net4966),
    .B1(net4379),
    .A1(_03047_),
    .Y(_01913_),
    .A2(net4705));
 sg13g2_nor3_1 _17493_ (.A(net4757),
    .B(_01911_),
    .C(_01913_),
    .Y(_01914_));
 sg13g2_a21oi_1 _17494_ (.A1(_02476_),
    .A2(net4760),
    .Y(_01357_),
    .B1(_01914_));
 sg13g2_a21oi_1 _17495_ (.A1(\m_sys.m_core.m_bru.io_i_s1[30] ),
    .A2(net4741),
    .Y(_01915_),
    .B1(net4348));
 sg13g2_o21ai_1 _17496_ (.B1(net4977),
    .Y(_01916_),
    .A1(_03055_),
    .A2(net4706));
 sg13g2_or2_1 _17497_ (.X(_01917_),
    .B(_01916_),
    .A(_01915_));
 sg13g2_a22oi_1 _17498_ (.Y(_01918_),
    .B1(_01917_),
    .B2(net5093),
    .A2(_03658_),
    .A1(net4966));
 sg13g2_a21o_1 _17499_ (.A2(net4757),
    .A1(net3215),
    .B1(_01918_),
    .X(_01358_));
 sg13g2_a21oi_1 _17500_ (.A1(net5353),
    .A2(net4741),
    .Y(_01919_),
    .B1(net4348));
 sg13g2_o21ai_1 _17501_ (.B1(net4977),
    .Y(_01920_),
    .A1(_03062_),
    .A2(net4707));
 sg13g2_o21ai_1 _17502_ (.B1(net4753),
    .Y(_01921_),
    .A1(_01919_),
    .A2(_01920_));
 sg13g2_a21oi_1 _17503_ (.A1(net4966),
    .A2(_03495_),
    .Y(_01922_),
    .B1(_01921_));
 sg13g2_a21oi_1 _17504_ (.A1(_02475_),
    .A2(net4757),
    .Y(_01359_),
    .B1(_01922_));
 sg13g2_nor4_1 _17505_ (.A(net5222),
    .B(net3444),
    .C(net4962),
    .D(_05306_),
    .Y(_01923_));
 sg13g2_a21o_1 _17506_ (.A2(net4962),
    .A1(net5256),
    .B1(_01923_),
    .X(_01360_));
 sg13g2_nor2_1 _17507_ (.A(_00027_),
    .B(net4794),
    .Y(_01924_));
 sg13g2_nand2b_1 _17508_ (.Y(_01925_),
    .B(_05609_),
    .A_N(_00027_));
 sg13g2_nor2_1 _17509_ (.A(net3222),
    .B(_01924_),
    .Y(_01926_));
 sg13g2_a21oi_1 _17510_ (.A1(net5311),
    .A2(\m_sys.m_core.m_bru.io_i_s2[0] ),
    .Y(_01927_),
    .B1(_01925_));
 sg13g2_nor3_1 _17511_ (.A(net5377),
    .B(net3223),
    .C(_01927_),
    .Y(_01361_));
 sg13g2_nor2_1 _17512_ (.A(net3173),
    .B(_01924_),
    .Y(_01928_));
 sg13g2_a21oi_1 _17513_ (.A1(net5311),
    .A2(\m_sys.m_core.m_bru.io_i_s2[1] ),
    .Y(_01929_),
    .B1(_01925_));
 sg13g2_nor3_1 _17514_ (.A(net5377),
    .B(net3174),
    .C(_01929_),
    .Y(_01362_));
 sg13g2_nand4_1 _17515_ (.B(_05292_),
    .C(_05294_),
    .A(net4974),
    .Y(_01930_),
    .D(_05302_));
 sg13g2_o21ai_1 _17516_ (.B1(_01930_),
    .Y(_01363_),
    .A1(_02459_),
    .A2(net4974));
 sg13g2_o21ai_1 _17517_ (.B1(_05293_),
    .Y(_01931_),
    .A1(net5319),
    .A2(_05306_));
 sg13g2_nand2_1 _17518_ (.Y(_01932_),
    .A(_05289_),
    .B(_05310_));
 sg13g2_nand2_1 _17519_ (.Y(_01933_),
    .A(_05294_),
    .B(_01932_));
 sg13g2_nor4_1 _17520_ (.A(\m_sys.m_core.m_bru.io_i_s1[25] ),
    .B(\m_sys.m_core.m_bru.io_i_s1[26] ),
    .C(\m_sys.m_core.m_bru.io_i_s1[27] ),
    .D(\m_sys.m_core.m_bru.io_i_s1[28] ),
    .Y(_01934_));
 sg13g2_nand4_1 _17521_ (.B(\m_sys.m_core.m_bru.io_i_s1[30] ),
    .C(_00080_),
    .A(net5192),
    .Y(_01935_),
    .D(_01934_));
 sg13g2_a221oi_1 _17522_ (.B2(_05310_),
    .C1(_05309_),
    .B1(_01935_),
    .A1(_01931_),
    .Y(_01936_),
    .A2(_01933_));
 sg13g2_a21o_1 _17523_ (.A2(net4962),
    .A1(net5244),
    .B1(_01936_),
    .X(_01364_));
 sg13g2_o21ai_1 _17524_ (.B1(net4786),
    .Y(_01365_),
    .A1(_02488_),
    .A2(net4973));
 sg13g2_nand2_1 _17525_ (.Y(_01937_),
    .A(net4973),
    .B(_02773_));
 sg13g2_or2_1 _17526_ (.X(_01938_),
    .B(_01937_),
    .A(net4957));
 sg13g2_or3_1 _17527_ (.A(net5315),
    .B(_05289_),
    .C(_01784_),
    .X(_01939_));
 sg13g2_a21oi_1 _17528_ (.A1(_05294_),
    .A2(_01939_),
    .Y(_01940_),
    .B1(_01938_));
 sg13g2_a21o_1 _17529_ (.A2(net4958),
    .A1(net3312),
    .B1(_01940_),
    .X(_01366_));
 sg13g2_nand2_1 _17530_ (.Y(_01941_),
    .A(net3176),
    .B(net4958));
 sg13g2_o21ai_1 _17531_ (.B1(_01941_),
    .Y(_01367_),
    .A1(_05310_),
    .A2(_01938_));
 sg13g2_a21o_1 _17532_ (.A2(net4958),
    .A1(net2946),
    .B1(net4733),
    .X(_01368_));
 sg13g2_or4_1 _17533_ (.A(net5317),
    .B(net5323),
    .C(_05286_),
    .D(_01937_),
    .X(_01942_));
 sg13g2_o21ai_1 _17534_ (.B1(_01942_),
    .Y(_01369_),
    .A1(_02501_),
    .A2(net4973));
 sg13g2_a21oi_2 _17535_ (.B1(net4965),
    .Y(_01943_),
    .A2(_02775_),
    .A1(_02772_));
 sg13g2_a22oi_1 _17536_ (.Y(_01370_),
    .B1(_03557_),
    .B2(_01943_),
    .A2(net4967),
    .A1(_02503_));
 sg13g2_nor2_1 _17537_ (.A(net3185),
    .B(net4976),
    .Y(_01944_));
 sg13g2_a21oi_1 _17538_ (.A1(_02385_),
    .A2(net4976),
    .Y(_01371_),
    .B1(_01944_));
 sg13g2_mux2_1 _17539_ (.A0(net5321),
    .A1(net3329),
    .S(net4968),
    .X(_01372_));
 sg13g2_nor2_1 _17540_ (.A(net2931),
    .B(net4976),
    .Y(_01945_));
 sg13g2_a21oi_1 _17541_ (.A1(net5228),
    .A2(net4976),
    .Y(_01373_),
    .B1(_01945_));
 sg13g2_nand2b_1 _17542_ (.Y(_01946_),
    .B(_02699_),
    .A_N(_02634_));
 sg13g2_a21oi_1 _17543_ (.A1(_02754_),
    .A2(_01946_),
    .Y(_01374_),
    .B1(net5376));
 sg13g2_nor2b_1 _17544_ (.A(net4316),
    .B_N(_05867_),
    .Y(_01947_));
 sg13g2_nor2_1 _17545_ (.A(net2791),
    .B(net4085),
    .Y(_01948_));
 sg13g2_a21oi_1 _17546_ (.A1(net5020),
    .A2(net4085),
    .Y(_01375_),
    .B1(_01948_));
 sg13g2_nor2_1 _17547_ (.A(net2762),
    .B(net4085),
    .Y(_01949_));
 sg13g2_a21oi_1 _17548_ (.A1(net4810),
    .A2(net4085),
    .Y(_01376_),
    .B1(_01949_));
 sg13g2_nor2_1 _17549_ (.A(net2208),
    .B(net4087),
    .Y(_01950_));
 sg13g2_a21oi_1 _17550_ (.A1(net5015),
    .A2(net4087),
    .Y(_01377_),
    .B1(_01950_));
 sg13g2_nor2_1 _17551_ (.A(net2554),
    .B(net4086),
    .Y(_01951_));
 sg13g2_a21oi_1 _17552_ (.A1(net4806),
    .A2(net4086),
    .Y(_01378_),
    .B1(_01951_));
 sg13g2_nor2_1 _17553_ (.A(net2668),
    .B(net4085),
    .Y(_01952_));
 sg13g2_a21oi_1 _17554_ (.A1(net5010),
    .A2(net4085),
    .Y(_01379_),
    .B1(_01952_));
 sg13g2_nor2_1 _17555_ (.A(net2699),
    .B(net4085),
    .Y(_01953_));
 sg13g2_a21oi_1 _17556_ (.A1(net4800),
    .A2(net4085),
    .Y(_01380_),
    .B1(_01953_));
 sg13g2_nor2_1 _17557_ (.A(net2515),
    .B(net4087),
    .Y(_01954_));
 sg13g2_a21oi_1 _17558_ (.A1(net5007),
    .A2(net4087),
    .Y(_01381_),
    .B1(_01954_));
 sg13g2_nor2_1 _17559_ (.A(net2855),
    .B(net4086),
    .Y(_01955_));
 sg13g2_a21oi_1 _17560_ (.A1(net4797),
    .A2(net4086),
    .Y(_01382_),
    .B1(_01955_));
 sg13g2_nor2b_1 _17561_ (.A(net4334),
    .B_N(_05391_),
    .Y(_01956_));
 sg13g2_nor2_1 _17562_ (.A(net2200),
    .B(net4083),
    .Y(_01957_));
 sg13g2_a21oi_1 _17563_ (.A1(net5135),
    .A2(net4083),
    .Y(_01383_),
    .B1(_01957_));
 sg13g2_nor2_1 _17564_ (.A(net2539),
    .B(net4083),
    .Y(_01958_));
 sg13g2_a21oi_1 _17565_ (.A1(net4996),
    .A2(net4083),
    .Y(_01384_),
    .B1(_01958_));
 sg13g2_nor2_1 _17566_ (.A(net2593),
    .B(net4084),
    .Y(_01959_));
 sg13g2_a21oi_1 _17567_ (.A1(net5134),
    .A2(net4084),
    .Y(_01385_),
    .B1(_01959_));
 sg13g2_nor2_1 _17568_ (.A(net2546),
    .B(net4083),
    .Y(_01960_));
 sg13g2_a21oi_1 _17569_ (.A1(net4992),
    .A2(net4083),
    .Y(_01386_),
    .B1(_01960_));
 sg13g2_nor2_1 _17570_ (.A(net2506),
    .B(net4084),
    .Y(_01961_));
 sg13g2_a21oi_1 _17571_ (.A1(net5129),
    .A2(net4084),
    .Y(_01387_),
    .B1(_01961_));
 sg13g2_nor2_1 _17572_ (.A(net2316),
    .B(net4083),
    .Y(_01962_));
 sg13g2_a21oi_1 _17573_ (.A1(net4985),
    .A2(net4083),
    .Y(_01388_),
    .B1(_01962_));
 sg13g2_nor2_1 _17574_ (.A(net2480),
    .B(net4084),
    .Y(_01963_));
 sg13g2_a21oi_1 _17575_ (.A1(net5123),
    .A2(net4084),
    .Y(_01389_),
    .B1(_01963_));
 sg13g2_nor2_1 _17576_ (.A(net2674),
    .B(net4084),
    .Y(_01964_));
 sg13g2_a21oi_1 _17577_ (.A1(net4982),
    .A2(net4084),
    .Y(_01390_),
    .B1(_01964_));
 sg13g2_nand2_1 _17578_ (.Y(_01965_),
    .A(net4330),
    .B(_05420_));
 sg13g2_nand2_1 _17579_ (.Y(_01966_),
    .A(net2078),
    .B(net4081));
 sg13g2_o21ai_1 _17580_ (.B1(_01966_),
    .Y(_01391_),
    .A1(net5045),
    .A2(net4081));
 sg13g2_nand2_1 _17581_ (.Y(_01967_),
    .A(net1871),
    .B(net4080));
 sg13g2_o21ai_1 _17582_ (.B1(_01967_),
    .Y(_01392_),
    .A1(net4875),
    .A2(net4081));
 sg13g2_nand2_1 _17583_ (.Y(_01968_),
    .A(net1735),
    .B(net4080));
 sg13g2_o21ai_1 _17584_ (.B1(_01968_),
    .Y(_01393_),
    .A1(net5040),
    .A2(net4080));
 sg13g2_nand2_1 _17585_ (.Y(_01969_),
    .A(net2145),
    .B(net4082));
 sg13g2_o21ai_1 _17586_ (.B1(_01969_),
    .Y(_01394_),
    .A1(net4870),
    .A2(net4082));
 sg13g2_nand2_1 _17587_ (.Y(_01970_),
    .A(net1990),
    .B(net4082));
 sg13g2_o21ai_1 _17588_ (.B1(_01970_),
    .Y(_01395_),
    .A1(net5030),
    .A2(net4082));
 sg13g2_nand2_1 _17589_ (.Y(_01971_),
    .A(net1954),
    .B(net4080));
 sg13g2_o21ai_1 _17590_ (.B1(_01971_),
    .Y(_01396_),
    .A1(net4868),
    .A2(net4080));
 sg13g2_nand2_1 _17591_ (.Y(_01972_),
    .A(net1676),
    .B(net4080));
 sg13g2_o21ai_1 _17592_ (.B1(_01972_),
    .Y(_01397_),
    .A1(net5027),
    .A2(net4080));
 sg13g2_nand2_1 _17593_ (.Y(_01973_),
    .A(net1679),
    .B(net4081));
 sg13g2_o21ai_1 _17594_ (.B1(_01973_),
    .Y(_01398_),
    .A1(net4859),
    .A2(net4080));
 sg13g2_nand2_1 _17595_ (.Y(_01974_),
    .A(net4322),
    .B(_05551_));
 sg13g2_nand2_1 _17596_ (.Y(_01975_),
    .A(net1952),
    .B(net4078));
 sg13g2_o21ai_1 _17597_ (.B1(_01975_),
    .Y(_01399_),
    .A1(net4855),
    .A2(net4078));
 sg13g2_nand2_1 _17598_ (.Y(_01976_),
    .A(net1774),
    .B(net4079));
 sg13g2_o21ai_1 _17599_ (.B1(_01976_),
    .Y(_01400_),
    .A1(net4851),
    .A2(net4079));
 sg13g2_nand2_1 _17600_ (.Y(_01977_),
    .A(net2025),
    .B(net4078));
 sg13g2_o21ai_1 _17601_ (.B1(_01977_),
    .Y(_01401_),
    .A1(net4844),
    .A2(net4078));
 sg13g2_nand2_1 _17602_ (.Y(_01978_),
    .A(net2114),
    .B(net4079));
 sg13g2_o21ai_1 _17603_ (.B1(_01978_),
    .Y(_01402_),
    .A1(net4839),
    .A2(net4079));
 sg13g2_nand2_1 _17604_ (.Y(_01979_),
    .A(net1792),
    .B(net4078));
 sg13g2_o21ai_1 _17605_ (.B1(_01979_),
    .Y(_01403_),
    .A1(net4836),
    .A2(net4078));
 sg13g2_nand2_1 _17606_ (.Y(_01980_),
    .A(net1983),
    .B(net4079));
 sg13g2_o21ai_1 _17607_ (.B1(_01980_),
    .Y(_01404_),
    .A1(net4829),
    .A2(net4079));
 sg13g2_nand2_1 _17608_ (.Y(_01981_),
    .A(net2243),
    .B(net4079));
 sg13g2_o21ai_1 _17609_ (.B1(_01981_),
    .Y(_01405_),
    .A1(net4822),
    .A2(net4079));
 sg13g2_nand2_1 _17610_ (.Y(_01982_),
    .A(net2176),
    .B(net4078));
 sg13g2_o21ai_1 _17611_ (.B1(_01982_),
    .Y(_01406_),
    .A1(net4815),
    .A2(net4078));
 sg13g2_nor2b_1 _17612_ (.A(net4314),
    .B_N(_05886_),
    .Y(_01983_));
 sg13g2_nor2_1 _17613_ (.A(net2490),
    .B(net4076),
    .Y(_01984_));
 sg13g2_a21oi_1 _17614_ (.A1(net5020),
    .A2(net4076),
    .Y(_01407_),
    .B1(_01984_));
 sg13g2_nor2_1 _17615_ (.A(net2734),
    .B(net4077),
    .Y(_01985_));
 sg13g2_a21oi_1 _17616_ (.A1(net4812),
    .A2(net4077),
    .Y(_01408_),
    .B1(_01985_));
 sg13g2_nor2_1 _17617_ (.A(net2714),
    .B(net4076),
    .Y(_01986_));
 sg13g2_a21oi_1 _17618_ (.A1(net5015),
    .A2(net4076),
    .Y(_01409_),
    .B1(_01986_));
 sg13g2_nor2_1 _17619_ (.A(net2565),
    .B(net4076),
    .Y(_01987_));
 sg13g2_a21oi_1 _17620_ (.A1(net4805),
    .A2(net4076),
    .Y(_01410_),
    .B1(_01987_));
 sg13g2_nor2_1 _17621_ (.A(net2344),
    .B(net4077),
    .Y(_01988_));
 sg13g2_a21oi_1 _17622_ (.A1(net5013),
    .A2(net4077),
    .Y(_01411_),
    .B1(_01988_));
 sg13g2_nor2_1 _17623_ (.A(net2527),
    .B(net4077),
    .Y(_01989_));
 sg13g2_a21oi_1 _17624_ (.A1(net4802),
    .A2(_01983_),
    .Y(_01412_),
    .B1(_01989_));
 sg13g2_nor2_1 _17625_ (.A(net2318),
    .B(net4077),
    .Y(_01990_));
 sg13g2_a21oi_1 _17626_ (.A1(net5008),
    .A2(net4077),
    .Y(_01413_),
    .B1(_01990_));
 sg13g2_nor2_1 _17627_ (.A(net2315),
    .B(net4076),
    .Y(_01991_));
 sg13g2_a21oi_1 _17628_ (.A1(net4796),
    .A2(net4076),
    .Y(_01414_),
    .B1(_01991_));
 sg13g2_nand2_1 _17629_ (.Y(_01992_),
    .A(net4326),
    .B(_07321_));
 sg13g2_nand2_1 _17630_ (.Y(_01993_),
    .A(net2278),
    .B(net4075));
 sg13g2_o21ai_1 _17631_ (.B1(_01993_),
    .Y(_01415_),
    .A1(net5042),
    .A2(net4075));
 sg13g2_nand2_1 _17632_ (.Y(_01994_),
    .A(net2183),
    .B(net4075));
 sg13g2_o21ai_1 _17633_ (.B1(_01994_),
    .Y(_01416_),
    .A1(net4877),
    .A2(net4075));
 sg13g2_nand2_1 _17634_ (.Y(_01995_),
    .A(net2265),
    .B(net4074));
 sg13g2_o21ai_1 _17635_ (.B1(_01995_),
    .Y(_01417_),
    .A1(net5035),
    .A2(net4074));
 sg13g2_nand2_1 _17636_ (.Y(_01996_),
    .A(net2589),
    .B(net4074));
 sg13g2_o21ai_1 _17637_ (.B1(_01996_),
    .Y(_01418_),
    .A1(net4869),
    .A2(net4074));
 sg13g2_nand2_1 _17638_ (.Y(_01997_),
    .A(net2144),
    .B(net4074));
 sg13g2_o21ai_1 _17639_ (.B1(_01997_),
    .Y(_01419_),
    .A1(net5031),
    .A2(net4074));
 sg13g2_nand2_1 _17640_ (.Y(_01998_),
    .A(net2066),
    .B(net4074));
 sg13g2_o21ai_1 _17641_ (.B1(_01998_),
    .Y(_01420_),
    .A1(net4864),
    .A2(net4074));
 sg13g2_nand2_1 _17642_ (.Y(_01999_),
    .A(net1973),
    .B(net4075));
 sg13g2_o21ai_1 _17643_ (.B1(_01999_),
    .Y(_01421_),
    .A1(net5029),
    .A2(net4075));
 sg13g2_nand2_1 _17644_ (.Y(_02000_),
    .A(net2002),
    .B(net4075));
 sg13g2_o21ai_1 _17645_ (.B1(_02000_),
    .Y(_01422_),
    .A1(net4863),
    .A2(net4075));
 sg13g2_nand2_1 _17646_ (.Y(_02001_),
    .A(net4320),
    .B(_07321_));
 sg13g2_nand2_1 _17647_ (.Y(_02002_),
    .A(net1939),
    .B(net4073));
 sg13g2_o21ai_1 _17648_ (.B1(_02002_),
    .Y(_01423_),
    .A1(net4854),
    .A2(net4073));
 sg13g2_nand2_1 _17649_ (.Y(_02003_),
    .A(net1749),
    .B(net4072));
 sg13g2_o21ai_1 _17650_ (.B1(_02003_),
    .Y(_01424_),
    .A1(net4847),
    .A2(net4071));
 sg13g2_nand2_1 _17651_ (.Y(_02004_),
    .A(net2093),
    .B(net4073));
 sg13g2_o21ai_1 _17652_ (.B1(_02004_),
    .Y(_01425_),
    .A1(net4843),
    .A2(net4073));
 sg13g2_nand2_1 _17653_ (.Y(_02005_),
    .A(net2155),
    .B(net4072));
 sg13g2_o21ai_1 _17654_ (.B1(_02005_),
    .Y(_01426_),
    .A1(net4837),
    .A2(net4073));
 sg13g2_nand2_1 _17655_ (.Y(_02006_),
    .A(net1959),
    .B(net4071));
 sg13g2_o21ai_1 _17656_ (.B1(_02006_),
    .Y(_01427_),
    .A1(net4831),
    .A2(net4071));
 sg13g2_nand2_1 _17657_ (.Y(_02007_),
    .A(net1847),
    .B(net4071));
 sg13g2_o21ai_1 _17658_ (.B1(_02007_),
    .Y(_01428_),
    .A1(net4825),
    .A2(net4072));
 sg13g2_nand2_1 _17659_ (.Y(_02008_),
    .A(net2057),
    .B(net4071));
 sg13g2_o21ai_1 _17660_ (.B1(_02008_),
    .Y(_01429_),
    .A1(net4821),
    .A2(net4071));
 sg13g2_nand2_1 _17661_ (.Y(_02009_),
    .A(net1766),
    .B(net4071));
 sg13g2_o21ai_1 _17662_ (.B1(_02009_),
    .Y(_01430_),
    .A1(net4816),
    .A2(net4071));
 sg13g2_nor2b_1 _17663_ (.A(net4332),
    .B_N(_07321_),
    .Y(_02010_));
 sg13g2_nor2_1 _17664_ (.A(net2238),
    .B(net4069),
    .Y(_02011_));
 sg13g2_a21oi_1 _17665_ (.A1(net5139),
    .A2(net4069),
    .Y(_01431_),
    .B1(_02011_));
 sg13g2_nor2_1 _17666_ (.A(net2294),
    .B(net4069),
    .Y(_02012_));
 sg13g2_a21oi_1 _17667_ (.A1(net4995),
    .A2(net4069),
    .Y(_01432_),
    .B1(_02012_));
 sg13g2_nor2_1 _17668_ (.A(net2683),
    .B(net4069),
    .Y(_02013_));
 sg13g2_a21oi_1 _17669_ (.A1(net5134),
    .A2(net4069),
    .Y(_01433_),
    .B1(_02013_));
 sg13g2_nor2_1 _17670_ (.A(net2806),
    .B(net4070),
    .Y(_02014_));
 sg13g2_a21oi_1 _17671_ (.A1(net4991),
    .A2(net4070),
    .Y(_01434_),
    .B1(_02014_));
 sg13g2_nor2_1 _17672_ (.A(net2491),
    .B(net4070),
    .Y(_02015_));
 sg13g2_a21oi_1 _17673_ (.A1(net5125),
    .A2(net4070),
    .Y(_01435_),
    .B1(_02015_));
 sg13g2_nor2_1 _17674_ (.A(net2413),
    .B(net4069),
    .Y(_02016_));
 sg13g2_a21oi_1 _17675_ (.A1(net4985),
    .A2(net4070),
    .Y(_01436_),
    .B1(_02016_));
 sg13g2_nor2_1 _17676_ (.A(net2462),
    .B(net4070),
    .Y(_02017_));
 sg13g2_a21oi_1 _17677_ (.A1(net5120),
    .A2(net4070),
    .Y(_01437_),
    .B1(_02017_));
 sg13g2_nor2_1 _17678_ (.A(net2496),
    .B(net4069),
    .Y(_02018_));
 sg13g2_a21oi_1 _17679_ (.A1(net4982),
    .A2(_02010_),
    .Y(_01438_),
    .B1(_02018_));
 sg13g2_nand2_1 _17680_ (.Y(_02019_),
    .A(net4328),
    .B(_05774_));
 sg13g2_nand2_1 _17681_ (.Y(_02020_),
    .A(net2077),
    .B(net4067));
 sg13g2_o21ai_1 _17682_ (.B1(_02020_),
    .Y(_01439_),
    .A1(net5043),
    .A2(net4067));
 sg13g2_nand2_1 _17683_ (.Y(_02021_),
    .A(net2035),
    .B(net4068));
 sg13g2_o21ai_1 _17684_ (.B1(_02021_),
    .Y(_01440_),
    .A1(net4875),
    .A2(net4068));
 sg13g2_nand2_1 _17685_ (.Y(_02022_),
    .A(net2013),
    .B(net4068));
 sg13g2_o21ai_1 _17686_ (.B1(_02022_),
    .Y(_01441_),
    .A1(net5038),
    .A2(_02019_));
 sg13g2_nand2_1 _17687_ (.Y(_02023_),
    .A(net1945),
    .B(net4067));
 sg13g2_o21ai_1 _17688_ (.B1(_02023_),
    .Y(_01442_),
    .A1(net4871),
    .A2(net4067));
 sg13g2_nand2_1 _17689_ (.Y(_02024_),
    .A(net1830),
    .B(net4067));
 sg13g2_o21ai_1 _17690_ (.B1(_02024_),
    .Y(_01443_),
    .A1(net5032),
    .A2(net4067));
 sg13g2_nand2_1 _17691_ (.Y(_02025_),
    .A(net1665),
    .B(net4067));
 sg13g2_o21ai_1 _17692_ (.B1(_02025_),
    .Y(_01444_),
    .A1(net4866),
    .A2(net4067));
 sg13g2_nand2_1 _17693_ (.Y(_02026_),
    .A(net2225),
    .B(net4068));
 sg13g2_o21ai_1 _17694_ (.B1(_02026_),
    .Y(_01445_),
    .A1(net5027),
    .A2(net4068));
 sg13g2_nand2_1 _17695_ (.Y(_02027_),
    .A(net2023),
    .B(net4068));
 sg13g2_o21ai_1 _17696_ (.B1(_02027_),
    .Y(_01446_),
    .A1(net4860),
    .A2(net4068));
 sg13g2_nand2_1 _17697_ (.Y(_02028_),
    .A(net4323),
    .B(_05774_));
 sg13g2_nand2_1 _17698_ (.Y(_02029_),
    .A(net1767),
    .B(net4066));
 sg13g2_o21ai_1 _17699_ (.B1(_02029_),
    .Y(_01447_),
    .A1(net4856),
    .A2(net4066));
 sg13g2_nand2_1 _17700_ (.Y(_02030_),
    .A(net2169),
    .B(net4065));
 sg13g2_o21ai_1 _17701_ (.B1(_02030_),
    .Y(_01448_),
    .A1(net4849),
    .A2(net4065));
 sg13g2_nand2_1 _17702_ (.Y(_02031_),
    .A(net1882),
    .B(net4066));
 sg13g2_o21ai_1 _17703_ (.B1(_02031_),
    .Y(_01449_),
    .A1(net4846),
    .A2(net4066));
 sg13g2_nand2_1 _17704_ (.Y(_02032_),
    .A(net1949),
    .B(net4066));
 sg13g2_o21ai_1 _17705_ (.B1(_02032_),
    .Y(_01450_),
    .A1(net4840),
    .A2(net4065));
 sg13g2_nand2_1 _17706_ (.Y(_02033_),
    .A(net1782),
    .B(net4066));
 sg13g2_o21ai_1 _17707_ (.B1(_02033_),
    .Y(_01451_),
    .A1(net4834),
    .A2(net4066));
 sg13g2_nand2_1 _17708_ (.Y(_02034_),
    .A(net1944),
    .B(net4065));
 sg13g2_o21ai_1 _17709_ (.B1(_02034_),
    .Y(_01452_),
    .A1(net4827),
    .A2(net4065));
 sg13g2_nand2_1 _17710_ (.Y(_02035_),
    .A(net1907),
    .B(net4065));
 sg13g2_o21ai_1 _17711_ (.B1(_02035_),
    .Y(_01453_),
    .A1(net4823),
    .A2(net4065));
 sg13g2_nand2_1 _17712_ (.Y(_02036_),
    .A(net1729),
    .B(_02028_));
 sg13g2_o21ai_1 _17713_ (.B1(_02036_),
    .Y(_01454_),
    .A1(net4818),
    .A2(net4065));
 sg13g2_nor2b_1 _17714_ (.A(net4333),
    .B_N(_05774_),
    .Y(_02037_));
 sg13g2_nor2_1 _17715_ (.A(net2502),
    .B(net4063),
    .Y(_02038_));
 sg13g2_a21oi_1 _17716_ (.A1(net5136),
    .A2(net4063),
    .Y(_01455_),
    .B1(_02038_));
 sg13g2_nor2_1 _17717_ (.A(net2313),
    .B(net4064),
    .Y(_02039_));
 sg13g2_a21oi_1 _17718_ (.A1(net4997),
    .A2(net4064),
    .Y(_01456_),
    .B1(_02039_));
 sg13g2_nor2_1 _17719_ (.A(net2525),
    .B(net4063),
    .Y(_02040_));
 sg13g2_a21oi_1 _17720_ (.A1(net5133),
    .A2(net4063),
    .Y(_01457_),
    .B1(_02040_));
 sg13g2_nor2_1 _17721_ (.A(net2677),
    .B(net4064),
    .Y(_02041_));
 sg13g2_a21oi_1 _17722_ (.A1(net4990),
    .A2(net4064),
    .Y(_01458_),
    .B1(_02041_));
 sg13g2_nor2_1 _17723_ (.A(net2521),
    .B(net4063),
    .Y(_02042_));
 sg13g2_a21oi_1 _17724_ (.A1(net5129),
    .A2(net4063),
    .Y(_01459_),
    .B1(_02042_));
 sg13g2_nor2_1 _17725_ (.A(net2814),
    .B(net4063),
    .Y(_02043_));
 sg13g2_a21oi_1 _17726_ (.A1(net4984),
    .A2(net4063),
    .Y(_01460_),
    .B1(_02043_));
 sg13g2_nor2_1 _17727_ (.A(net2727),
    .B(net4064),
    .Y(_02044_));
 sg13g2_a21oi_1 _17728_ (.A1(net5123),
    .A2(net4064),
    .Y(_01461_),
    .B1(_02044_));
 sg13g2_nor2_1 _17729_ (.A(net2437),
    .B(net4064),
    .Y(_02045_));
 sg13g2_a21oi_1 _17730_ (.A1(net4981),
    .A2(net4064),
    .Y(_01462_),
    .B1(_02045_));
 sg13g2_nand2_1 _17731_ (.Y(_02046_),
    .A(net4328),
    .B(_05848_));
 sg13g2_nand2_1 _17732_ (.Y(_02047_),
    .A(net1669),
    .B(net4062));
 sg13g2_o21ai_1 _17733_ (.B1(_02047_),
    .Y(_01463_),
    .A1(net5043),
    .A2(net4061));
 sg13g2_nand2_1 _17734_ (.Y(_02048_),
    .A(net1808),
    .B(net4062));
 sg13g2_o21ai_1 _17735_ (.B1(_02048_),
    .Y(_01464_),
    .A1(net4875),
    .A2(net4062));
 sg13g2_nand2_1 _17736_ (.Y(_02049_),
    .A(net1683),
    .B(_02046_));
 sg13g2_o21ai_1 _17737_ (.B1(_02049_),
    .Y(_01465_),
    .A1(net5038),
    .A2(net4061));
 sg13g2_nand2_1 _17738_ (.Y(_02050_),
    .A(net2143),
    .B(net4061));
 sg13g2_o21ai_1 _17739_ (.B1(_02050_),
    .Y(_01466_),
    .A1(net4871),
    .A2(net4061));
 sg13g2_nand2_1 _17740_ (.Y(_02051_),
    .A(net1934),
    .B(net4061));
 sg13g2_o21ai_1 _17741_ (.B1(_02051_),
    .Y(_01467_),
    .A1(net5032),
    .A2(net4061));
 sg13g2_nand2_1 _17742_ (.Y(_02052_),
    .A(net1857),
    .B(net4061));
 sg13g2_o21ai_1 _17743_ (.B1(_02052_),
    .Y(_01468_),
    .A1(net4866),
    .A2(net4061));
 sg13g2_nand2_1 _17744_ (.Y(_02053_),
    .A(net2075),
    .B(net4062));
 sg13g2_o21ai_1 _17745_ (.B1(_02053_),
    .Y(_01469_),
    .A1(net5027),
    .A2(net4062));
 sg13g2_nand2_1 _17746_ (.Y(_02054_),
    .A(net1780),
    .B(net4062));
 sg13g2_o21ai_1 _17747_ (.B1(_02054_),
    .Y(_01470_),
    .A1(net4860),
    .A2(net4062));
 sg13g2_nor2_1 _17748_ (.A(\m_sys.m_core.m_gpr.io_b_write_addr[1] ),
    .B(_07465_),
    .Y(_02055_));
 sg13g2_nor3_1 _17749_ (.A(\m_sys.m_core.m_gpr.io_b_write_addr[0] ),
    .B(\m_sys.m_core.m_gpr.io_b_write_addr[1] ),
    .C(_07465_),
    .Y(_02056_));
 sg13g2_nor2_1 _17750_ (.A(net3117),
    .B(net4426),
    .Y(_02057_));
 sg13g2_a21oi_1 _17751_ (.A1(_02397_),
    .A2(net4426),
    .Y(_01471_),
    .B1(_02057_));
 sg13g2_mux2_1 _17752_ (.A0(net2988),
    .A1(\m_sys.m_core.m_bru.io_i_s1[1] ),
    .S(net4428),
    .X(_01472_));
 sg13g2_nor2_1 _17753_ (.A(net3050),
    .B(net4429),
    .Y(_02058_));
 sg13g2_a21oi_1 _17754_ (.A1(_02371_),
    .A2(net4429),
    .Y(_01473_),
    .B1(_02058_));
 sg13g2_mux2_1 _17755_ (.A0(net3069),
    .A1(net5314),
    .S(net4430),
    .X(_01474_));
 sg13g2_mux2_1 _17756_ (.A0(net2987),
    .A1(net5316),
    .S(net4425),
    .X(_01475_));
 sg13g2_mux2_1 _17757_ (.A0(net2981),
    .A1(\m_sys.m_core.m_bru.io_i_s1[5] ),
    .S(net4427),
    .X(_01476_));
 sg13g2_nor2_1 _17758_ (.A(net3048),
    .B(net4426),
    .Y(_02059_));
 sg13g2_a21oi_1 _17759_ (.A1(net5226),
    .A2(net4426),
    .Y(_01477_),
    .B1(_02059_));
 sg13g2_nor2_1 _17760_ (.A(net3082),
    .B(net4428),
    .Y(_02060_));
 sg13g2_a21oi_1 _17761_ (.A1(net5227),
    .A2(net4428),
    .Y(_01478_),
    .B1(_02060_));
 sg13g2_mux2_1 _17762_ (.A0(net3008),
    .A1(net5321),
    .S(net4430),
    .X(_01479_));
 sg13g2_nor2_1 _17763_ (.A(net3052),
    .B(net4428),
    .Y(_02061_));
 sg13g2_a21oi_1 _17764_ (.A1(net5228),
    .A2(net4425),
    .Y(_01480_),
    .B1(_02061_));
 sg13g2_nor2_1 _17765_ (.A(net2953),
    .B(net4428),
    .Y(_02062_));
 sg13g2_a21oi_1 _17766_ (.A1(_02383_),
    .A2(net4428),
    .Y(_01481_),
    .B1(_02062_));
 sg13g2_nor2_1 _17767_ (.A(net2944),
    .B(net4429),
    .Y(_02063_));
 sg13g2_a21oi_1 _17768_ (.A1(_02381_),
    .A2(net4429),
    .Y(_01482_),
    .B1(_02063_));
 sg13g2_nor2_1 _17769_ (.A(net2883),
    .B(net4431),
    .Y(_02064_));
 sg13g2_a21oi_1 _17770_ (.A1(net5223),
    .A2(net4431),
    .Y(_01483_),
    .B1(_02064_));
 sg13g2_nor2_1 _17771_ (.A(net2898),
    .B(net4429),
    .Y(_02065_));
 sg13g2_a21oi_1 _17772_ (.A1(net5225),
    .A2(net4429),
    .Y(_01484_),
    .B1(_02065_));
 sg13g2_nor2_1 _17773_ (.A(net2976),
    .B(net4432),
    .Y(_02066_));
 sg13g2_a21oi_1 _17774_ (.A1(_02400_),
    .A2(net4431),
    .Y(_01485_),
    .B1(_02066_));
 sg13g2_nor2_1 _17775_ (.A(net3187),
    .B(net4433),
    .Y(_02067_));
 sg13g2_a21oi_1 _17776_ (.A1(net5191),
    .A2(net4433),
    .Y(_01486_),
    .B1(_02067_));
 sg13g2_nor2_1 _17777_ (.A(net3047),
    .B(net4433),
    .Y(_02068_));
 sg13g2_a21oi_1 _17778_ (.A1(net5187),
    .A2(net4433),
    .Y(_01487_),
    .B1(_02068_));
 sg13g2_nor2_1 _17779_ (.A(net3036),
    .B(net4431),
    .Y(_02069_));
 sg13g2_a21oi_1 _17780_ (.A1(net5180),
    .A2(net4431),
    .Y(_01488_),
    .B1(_02069_));
 sg13g2_nor2_1 _17781_ (.A(net2960),
    .B(net4430),
    .Y(_02070_));
 sg13g2_a21oi_1 _17782_ (.A1(_02450_),
    .A2(net4430),
    .Y(_01489_),
    .B1(_02070_));
 sg13g2_nor2_1 _17783_ (.A(net2971),
    .B(net4433),
    .Y(_02071_));
 sg13g2_a21oi_1 _17784_ (.A1(_02452_),
    .A2(net4433),
    .Y(_01490_),
    .B1(_02071_));
 sg13g2_nor2_1 _17785_ (.A(net3081),
    .B(net4432),
    .Y(_02072_));
 sg13g2_a21oi_1 _17786_ (.A1(net5201),
    .A2(net4432),
    .Y(_01491_),
    .B1(_02072_));
 sg13g2_nor2_1 _17787_ (.A(net2914),
    .B(net4431),
    .Y(_02073_));
 sg13g2_a21oi_1 _17788_ (.A1(net5219),
    .A2(net4431),
    .Y(_01492_),
    .B1(_02073_));
 sg13g2_nor2_1 _17789_ (.A(net3005),
    .B(net4432),
    .Y(_02074_));
 sg13g2_a21oi_1 _17790_ (.A1(net5212),
    .A2(net4431),
    .Y(_01493_),
    .B1(_02074_));
 sg13g2_nor2_1 _17791_ (.A(net3073),
    .B(net4432),
    .Y(_02075_));
 sg13g2_a21oi_1 _17792_ (.A1(_02427_),
    .A2(net4432),
    .Y(_01494_),
    .B1(_02075_));
 sg13g2_nor2_1 _17793_ (.A(net2930),
    .B(net4427),
    .Y(_02076_));
 sg13g2_a21oi_1 _17794_ (.A1(net5196),
    .A2(net4427),
    .Y(_01495_),
    .B1(_02076_));
 sg13g2_nor2_1 _17795_ (.A(net3014),
    .B(net4428),
    .Y(_02077_));
 sg13g2_a21oi_1 _17796_ (.A1(_02432_),
    .A2(net4427),
    .Y(_01496_),
    .B1(_02077_));
 sg13g2_nor2_1 _17797_ (.A(net3058),
    .B(net4425),
    .Y(_02078_));
 sg13g2_a21oi_1 _17798_ (.A1(net5194),
    .A2(net4425),
    .Y(_01497_),
    .B1(_02078_));
 sg13g2_nor2_1 _17799_ (.A(net2942),
    .B(net4427),
    .Y(_02079_));
 sg13g2_a21oi_1 _17800_ (.A1(net5193),
    .A2(net4427),
    .Y(_01498_),
    .B1(_02079_));
 sg13g2_nor2_1 _17801_ (.A(net2949),
    .B(net4427),
    .Y(_02080_));
 sg13g2_a21oi_1 _17802_ (.A1(_02439_),
    .A2(net4427),
    .Y(_01499_),
    .B1(_02080_));
 sg13g2_nor2_1 _17803_ (.A(net2870),
    .B(net4429),
    .Y(_02081_));
 sg13g2_a21oi_1 _17804_ (.A1(net5192),
    .A2(net4429),
    .Y(_01500_),
    .B1(_02081_));
 sg13g2_nor2_1 _17805_ (.A(net2859),
    .B(net4425),
    .Y(_02082_));
 sg13g2_a21oi_1 _17806_ (.A1(_02443_),
    .A2(net4425),
    .Y(_01501_),
    .B1(_02082_));
 sg13g2_nor2_1 _17807_ (.A(net3034),
    .B(net4425),
    .Y(_02083_));
 sg13g2_a21oi_1 _17808_ (.A1(_02444_),
    .A2(net4425),
    .Y(_01502_),
    .B1(_02083_));
 sg13g2_nor2_1 _17809_ (.A(\m_sys.m_core.m_gpr.io_b_write_addr[2] ),
    .B(_07464_),
    .Y(_02084_));
 sg13g2_nor3_1 _17810_ (.A(\m_sys.m_core.m_gpr.io_b_write_addr[2] ),
    .B(_07464_),
    .C(_07466_),
    .Y(_02085_));
 sg13g2_nor2_1 _17811_ (.A(net3011),
    .B(net4695),
    .Y(_02086_));
 sg13g2_a21oi_1 _17812_ (.A1(_02397_),
    .A2(net4695),
    .Y(_01503_),
    .B1(_02086_));
 sg13g2_mux2_1 _17813_ (.A0(net3059),
    .A1(\m_sys.m_core.m_bru.io_i_s1[1] ),
    .S(net4695),
    .X(_01504_));
 sg13g2_nor2_1 _17814_ (.A(net2900),
    .B(net4700),
    .Y(_02087_));
 sg13g2_a21oi_1 _17815_ (.A1(_02371_),
    .A2(net4700),
    .Y(_01505_),
    .B1(_02087_));
 sg13g2_mux2_1 _17816_ (.A0(net3070),
    .A1(net5314),
    .S(net4700),
    .X(_01506_));
 sg13g2_mux2_1 _17817_ (.A0(net3065),
    .A1(net5316),
    .S(net4695),
    .X(_01507_));
 sg13g2_mux2_1 _17818_ (.A0(net3024),
    .A1(\m_sys.m_core.m_bru.io_i_s1[5] ),
    .S(net4693),
    .X(_01508_));
 sg13g2_nor2_1 _17819_ (.A(net2449),
    .B(net4695),
    .Y(_02088_));
 sg13g2_a21oi_1 _17820_ (.A1(net5226),
    .A2(net4695),
    .Y(_01509_),
    .B1(_02088_));
 sg13g2_nor2_1 _17821_ (.A(net2967),
    .B(net4696),
    .Y(_02089_));
 sg13g2_a21oi_1 _17822_ (.A1(net5227),
    .A2(net4696),
    .Y(_01510_),
    .B1(_02089_));
 sg13g2_mux2_1 _17823_ (.A0(net3042),
    .A1(net5321),
    .S(net4700),
    .X(_01511_));
 sg13g2_nor2_1 _17824_ (.A(net2910),
    .B(net4696),
    .Y(_02090_));
 sg13g2_a21oi_1 _17825_ (.A1(net5228),
    .A2(net4696),
    .Y(_01512_),
    .B1(_02090_));
 sg13g2_nor2_1 _17826_ (.A(net3009),
    .B(net4695),
    .Y(_02091_));
 sg13g2_a21oi_1 _17827_ (.A1(_02383_),
    .A2(net4695),
    .Y(_01513_),
    .B1(_02091_));
 sg13g2_nor2_1 _17828_ (.A(net2929),
    .B(net4698),
    .Y(_02092_));
 sg13g2_a21oi_1 _17829_ (.A1(net5230),
    .A2(net4698),
    .Y(_01514_),
    .B1(_02092_));
 sg13g2_nor2_1 _17830_ (.A(net3013),
    .B(net4697),
    .Y(_02093_));
 sg13g2_a21oi_1 _17831_ (.A1(net5223),
    .A2(net4697),
    .Y(_01515_),
    .B1(_02093_));
 sg13g2_nor2_1 _17832_ (.A(net2993),
    .B(net4698),
    .Y(_02094_));
 sg13g2_a21oi_1 _17833_ (.A1(net5225),
    .A2(net4698),
    .Y(_01516_),
    .B1(_02094_));
 sg13g2_nor2_1 _17834_ (.A(net2951),
    .B(net4699),
    .Y(_02095_));
 sg13g2_a21oi_1 _17835_ (.A1(net5222),
    .A2(net4699),
    .Y(_01517_),
    .B1(_02095_));
 sg13g2_nor2_1 _17836_ (.A(net2924),
    .B(net4699),
    .Y(_02096_));
 sg13g2_a21oi_1 _17837_ (.A1(net5191),
    .A2(net4699),
    .Y(_01518_),
    .B1(_02096_));
 sg13g2_nor2_1 _17838_ (.A(net2894),
    .B(net4699),
    .Y(_02097_));
 sg13g2_a21oi_1 _17839_ (.A1(net5188),
    .A2(net4700),
    .Y(_01519_),
    .B1(_02097_));
 sg13g2_nor2_1 _17840_ (.A(net3103),
    .B(net4699),
    .Y(_02098_));
 sg13g2_a21oi_1 _17841_ (.A1(net5181),
    .A2(net4699),
    .Y(_01520_),
    .B1(_02098_));
 sg13g2_nor2_1 _17842_ (.A(net2923),
    .B(net4700),
    .Y(_02099_));
 sg13g2_a21oi_1 _17843_ (.A1(net5177),
    .A2(net4700),
    .Y(_01521_),
    .B1(_02099_));
 sg13g2_nor2_1 _17844_ (.A(net2889),
    .B(net4701),
    .Y(_02100_));
 sg13g2_a21oi_1 _17845_ (.A1(net5176),
    .A2(net4699),
    .Y(_01522_),
    .B1(_02100_));
 sg13g2_nor2_1 _17846_ (.A(net3044),
    .B(net4697),
    .Y(_02101_));
 sg13g2_a21oi_1 _17847_ (.A1(net5201),
    .A2(net4697),
    .Y(_01523_),
    .B1(_02101_));
 sg13g2_nor2_1 _17848_ (.A(net2947),
    .B(net4697),
    .Y(_02102_));
 sg13g2_a21oi_1 _17849_ (.A1(net5219),
    .A2(net4697),
    .Y(_01524_),
    .B1(_02102_));
 sg13g2_nor2_1 _17850_ (.A(net3000),
    .B(net4698),
    .Y(_02103_));
 sg13g2_a21oi_1 _17851_ (.A1(net5212),
    .A2(net4701),
    .Y(_01525_),
    .B1(_02103_));
 sg13g2_nor2_1 _17852_ (.A(net2963),
    .B(net4697),
    .Y(_02104_));
 sg13g2_a21oi_1 _17853_ (.A1(net5197),
    .A2(net4697),
    .Y(_01526_),
    .B1(_02104_));
 sg13g2_nor2_1 _17854_ (.A(net2992),
    .B(net4694),
    .Y(_02105_));
 sg13g2_a21oi_1 _17855_ (.A1(net5196),
    .A2(net4694),
    .Y(_01527_),
    .B1(_02105_));
 sg13g2_nor2_1 _17856_ (.A(net3040),
    .B(net4694),
    .Y(_02106_));
 sg13g2_a21oi_1 _17857_ (.A1(net5195),
    .A2(net4694),
    .Y(_01528_),
    .B1(_02106_));
 sg13g2_nor2_1 _17858_ (.A(net3057),
    .B(net4693),
    .Y(_02107_));
 sg13g2_a21oi_1 _17859_ (.A1(net5194),
    .A2(net4693),
    .Y(_01529_),
    .B1(_02107_));
 sg13g2_nor2_1 _17860_ (.A(net3016),
    .B(net4694),
    .Y(_02108_));
 sg13g2_a21oi_1 _17861_ (.A1(net5193),
    .A2(net4693),
    .Y(_01530_),
    .B1(_02108_));
 sg13g2_nor2_1 _17862_ (.A(net3029),
    .B(net4694),
    .Y(_02109_));
 sg13g2_a21oi_1 _17863_ (.A1(_02439_),
    .A2(net4694),
    .Y(_01531_),
    .B1(_02109_));
 sg13g2_nor2_1 _17864_ (.A(net3017),
    .B(net4698),
    .Y(_02110_));
 sg13g2_a21oi_1 _17865_ (.A1(net5192),
    .A2(net4698),
    .Y(_01532_),
    .B1(_02110_));
 sg13g2_nor2_1 _17866_ (.A(net2968),
    .B(net4693),
    .Y(_02111_));
 sg13g2_a21oi_1 _17867_ (.A1(_02443_),
    .A2(net4693),
    .Y(_01533_),
    .B1(_02111_));
 sg13g2_nor2_1 _17868_ (.A(net2994),
    .B(net4693),
    .Y(_02112_));
 sg13g2_a21oi_1 _17869_ (.A1(_02444_),
    .A2(net4693),
    .Y(_01534_),
    .B1(_02112_));
 sg13g2_nor2b_1 _17870_ (.A(\m_sys.m_core.m_gpr.io_b_write_addr[0] ),
    .B_N(\m_sys.m_core.m_gpr.io_b_write_addr[1] ),
    .Y(_02113_));
 sg13g2_nand2_1 _17871_ (.Y(_02114_),
    .A(_02084_),
    .B(_02113_));
 sg13g2_nand2_1 _17872_ (.Y(_02115_),
    .A(net1980),
    .B(net4417));
 sg13g2_o21ai_1 _17873_ (.B1(_02115_),
    .Y(_01535_),
    .A1(_02397_),
    .A2(net4417));
 sg13g2_nor2_1 _17874_ (.A(net5312),
    .B(net4417),
    .Y(_02116_));
 sg13g2_a21oi_1 _17875_ (.A1(_02425_),
    .A2(net4417),
    .Y(_01536_),
    .B1(_02116_));
 sg13g2_nand2_1 _17876_ (.Y(_02117_),
    .A(net2748),
    .B(net4423));
 sg13g2_o21ai_1 _17877_ (.B1(_02117_),
    .Y(_01537_),
    .A1(net5231),
    .A2(net4423));
 sg13g2_mux2_1 _17878_ (.A0(net5314),
    .A1(net2978),
    .S(net4423),
    .X(_01538_));
 sg13g2_nor2_1 _17879_ (.A(net5316),
    .B(net4417),
    .Y(_02118_));
 sg13g2_a21oi_1 _17880_ (.A1(_02431_),
    .A2(net4417),
    .Y(_01539_),
    .B1(_02118_));
 sg13g2_mux2_1 _17881_ (.A0(net5319),
    .A1(net3021),
    .S(net4416),
    .X(_01540_));
 sg13g2_nand2_1 _17882_ (.Y(_02119_),
    .A(net2359),
    .B(net4417));
 sg13g2_o21ai_1 _17883_ (.B1(_02119_),
    .Y(_01541_),
    .A1(net5226),
    .A2(net4417));
 sg13g2_nand2_1 _17884_ (.Y(_02120_),
    .A(net2083),
    .B(net4418));
 sg13g2_o21ai_1 _17885_ (.B1(_02120_),
    .Y(_01542_),
    .A1(net5227),
    .A2(net4418));
 sg13g2_mux2_1 _17886_ (.A0(net5321),
    .A1(net3018),
    .S(net4423),
    .X(_01543_));
 sg13g2_nand2_1 _17887_ (.Y(_02121_),
    .A(net2542),
    .B(net4418));
 sg13g2_o21ai_1 _17888_ (.B1(_02121_),
    .Y(_01544_),
    .A1(net5228),
    .A2(net4418));
 sg13g2_nand2_1 _17889_ (.Y(_02122_),
    .A(net2331),
    .B(net4416));
 sg13g2_o21ai_1 _17890_ (.B1(_02122_),
    .Y(_01545_),
    .A1(net5229),
    .A2(net4416));
 sg13g2_nand2_1 _17891_ (.Y(_02123_),
    .A(net2447),
    .B(net4421));
 sg13g2_o21ai_1 _17892_ (.B1(_02123_),
    .Y(_01546_),
    .A1(net5230),
    .A2(net4421));
 sg13g2_nand2_1 _17893_ (.Y(_02124_),
    .A(net2350),
    .B(net4420));
 sg13g2_o21ai_1 _17894_ (.B1(_02124_),
    .Y(_01547_),
    .A1(net5223),
    .A2(net4420));
 sg13g2_nand2_1 _17895_ (.Y(_02125_),
    .A(net2421),
    .B(net4421));
 sg13g2_o21ai_1 _17896_ (.B1(_02125_),
    .Y(_01548_),
    .A1(net5225),
    .A2(net4421));
 sg13g2_nand2_1 _17897_ (.Y(_02126_),
    .A(net2329),
    .B(net4422));
 sg13g2_o21ai_1 _17898_ (.B1(_02126_),
    .Y(_01549_),
    .A1(net5222),
    .A2(net4422));
 sg13g2_nand2_1 _17899_ (.Y(_02127_),
    .A(net2708),
    .B(net4422));
 sg13g2_o21ai_1 _17900_ (.B1(_02127_),
    .Y(_01550_),
    .A1(net5191),
    .A2(net4422));
 sg13g2_nand2_1 _17901_ (.Y(_02128_),
    .A(net2670),
    .B(net4422));
 sg13g2_o21ai_1 _17902_ (.B1(_02128_),
    .Y(_01551_),
    .A1(net5187),
    .A2(net4422));
 sg13g2_nand2_1 _17903_ (.Y(_02129_),
    .A(net2309),
    .B(net4422));
 sg13g2_o21ai_1 _17904_ (.B1(_02129_),
    .Y(_01552_),
    .A1(net5183),
    .A2(net4422));
 sg13g2_nand2_1 _17905_ (.Y(_02130_),
    .A(net2682),
    .B(net4423));
 sg13g2_o21ai_1 _17906_ (.B1(_02130_),
    .Y(_01553_),
    .A1(net5177),
    .A2(net4423));
 sg13g2_nand2_1 _17907_ (.Y(_02131_),
    .A(net2014),
    .B(net4423));
 sg13g2_o21ai_1 _17908_ (.B1(_02131_),
    .Y(_01554_),
    .A1(net5176),
    .A2(net4424));
 sg13g2_nand2_1 _17909_ (.Y(_02132_),
    .A(net2312),
    .B(net4420));
 sg13g2_o21ai_1 _17910_ (.B1(_02132_),
    .Y(_01555_),
    .A1(net5201),
    .A2(net4420));
 sg13g2_nand2_1 _17911_ (.Y(_02133_),
    .A(net2137),
    .B(net4424));
 sg13g2_o21ai_1 _17912_ (.B1(_02133_),
    .Y(_01556_),
    .A1(net5219),
    .A2(net4424));
 sg13g2_nand2_1 _17913_ (.Y(_02134_),
    .A(net2484),
    .B(net4420));
 sg13g2_o21ai_1 _17914_ (.B1(_02134_),
    .Y(_01557_),
    .A1(net5212),
    .A2(net4420));
 sg13g2_nand2_1 _17915_ (.Y(_02135_),
    .A(net2612),
    .B(net4420));
 sg13g2_o21ai_1 _17916_ (.B1(_02135_),
    .Y(_01558_),
    .A1(net5197),
    .A2(net4420));
 sg13g2_nand2_1 _17917_ (.Y(_02136_),
    .A(net2383),
    .B(net4416));
 sg13g2_o21ai_1 _17918_ (.B1(_02136_),
    .Y(_01559_),
    .A1(net5196),
    .A2(net4416));
 sg13g2_nand2_1 _17919_ (.Y(_02137_),
    .A(net2537),
    .B(net4421));
 sg13g2_o21ai_1 _17920_ (.B1(_02137_),
    .Y(_01560_),
    .A1(net5195),
    .A2(net4421));
 sg13g2_nand2_1 _17921_ (.Y(_02138_),
    .A(net2275),
    .B(net4415));
 sg13g2_o21ai_1 _17922_ (.B1(_02138_),
    .Y(_01561_),
    .A1(net5194),
    .A2(net4415));
 sg13g2_nor2_1 _17923_ (.A(\m_sys.m_core.m_bru.io_i_s1[27] ),
    .B(net4415),
    .Y(_02139_));
 sg13g2_a21oi_1 _17924_ (.A1(_02455_),
    .A2(net4415),
    .Y(_01562_),
    .B1(_02139_));
 sg13g2_nand2_1 _17925_ (.Y(_02140_),
    .A(net2134),
    .B(net4416));
 sg13g2_o21ai_1 _17926_ (.B1(_02140_),
    .Y(_01563_),
    .A1(_02439_),
    .A2(net4416));
 sg13g2_nand2_1 _17927_ (.Y(_02141_),
    .A(net2185),
    .B(net4421));
 sg13g2_o21ai_1 _17928_ (.B1(_02141_),
    .Y(_01564_),
    .A1(net5192),
    .A2(net4421));
 sg13g2_nand2_1 _17929_ (.Y(_02142_),
    .A(net2130),
    .B(net4415));
 sg13g2_o21ai_1 _17930_ (.B1(_02142_),
    .Y(_01565_),
    .A1(_02443_),
    .A2(net4415));
 sg13g2_nand2_1 _17931_ (.Y(_02143_),
    .A(net2384),
    .B(net4415));
 sg13g2_o21ai_1 _17932_ (.B1(_02143_),
    .Y(_01566_),
    .A1(_02444_),
    .A2(net4415));
 sg13g2_nand3b_1 _17933_ (.B(_02084_),
    .C(\m_sys.m_core.m_gpr.io_b_write_addr[0] ),
    .Y(_02144_),
    .A_N(\m_sys.m_core.m_gpr.io_b_write_addr[1] ));
 sg13g2_nand2_1 _17934_ (.Y(_02145_),
    .A(net2031),
    .B(net4408));
 sg13g2_o21ai_1 _17935_ (.B1(_02145_),
    .Y(_01567_),
    .A1(_02397_),
    .A2(net4408));
 sg13g2_mux2_1 _17936_ (.A0(net5312),
    .A1(net3120),
    .S(net4408),
    .X(_01568_));
 sg13g2_nand2_1 _17937_ (.Y(_02146_),
    .A(net2425),
    .B(net4413));
 sg13g2_o21ai_1 _17938_ (.B1(_02146_),
    .Y(_01569_),
    .A1(net5231),
    .A2(net4413));
 sg13g2_mux2_1 _17939_ (.A0(net5314),
    .A1(net3097),
    .S(net4413),
    .X(_01570_));
 sg13g2_mux2_1 _17940_ (.A0(net5316),
    .A1(net3119),
    .S(net4408),
    .X(_01571_));
 sg13g2_mux2_1 _17941_ (.A0(net5319),
    .A1(net3075),
    .S(net4407),
    .X(_01572_));
 sg13g2_nand2_1 _17942_ (.Y(_02147_),
    .A(net2536),
    .B(net4408));
 sg13g2_o21ai_1 _17943_ (.B1(_02147_),
    .Y(_01573_),
    .A1(net5226),
    .A2(net4408));
 sg13g2_nand2_1 _17944_ (.Y(_02148_),
    .A(net2687),
    .B(net4408));
 sg13g2_o21ai_1 _17945_ (.B1(_02148_),
    .Y(_01574_),
    .A1(net5227),
    .A2(net4408));
 sg13g2_mux2_1 _17946_ (.A0(net5320),
    .A1(net3086),
    .S(net4413),
    .X(_01575_));
 sg13g2_nand2_1 _17947_ (.Y(_02149_),
    .A(net2307),
    .B(net4409));
 sg13g2_o21ai_1 _17948_ (.B1(_02149_),
    .Y(_01576_),
    .A1(net5228),
    .A2(net4409));
 sg13g2_nand2_1 _17949_ (.Y(_02150_),
    .A(net2486),
    .B(net4407));
 sg13g2_o21ai_1 _17950_ (.B1(_02150_),
    .Y(_01577_),
    .A1(net5229),
    .A2(net4407));
 sg13g2_nand2_1 _17951_ (.Y(_02151_),
    .A(net2664),
    .B(net4411));
 sg13g2_o21ai_1 _17952_ (.B1(_02151_),
    .Y(_01578_),
    .A1(net5230),
    .A2(net4411));
 sg13g2_nand2_1 _17953_ (.Y(_02152_),
    .A(net2401),
    .B(net4410));
 sg13g2_o21ai_1 _17954_ (.B1(_02152_),
    .Y(_01579_),
    .A1(net5223),
    .A2(net4410));
 sg13g2_nand2_1 _17955_ (.Y(_02153_),
    .A(net2514),
    .B(net4411));
 sg13g2_o21ai_1 _17956_ (.B1(_02153_),
    .Y(_01580_),
    .A1(net5224),
    .A2(net4411));
 sg13g2_nand2_1 _17957_ (.Y(_02154_),
    .A(net2807),
    .B(net4412));
 sg13g2_o21ai_1 _17958_ (.B1(_02154_),
    .Y(_01581_),
    .A1(net5222),
    .A2(net4412));
 sg13g2_nand2_1 _17959_ (.Y(_02155_),
    .A(net2830),
    .B(net4412));
 sg13g2_o21ai_1 _17960_ (.B1(_02155_),
    .Y(_01582_),
    .A1(net5191),
    .A2(net4412));
 sg13g2_nand2_1 _17961_ (.Y(_02156_),
    .A(net2792),
    .B(net4412));
 sg13g2_o21ai_1 _17962_ (.B1(_02156_),
    .Y(_01583_),
    .A1(net5187),
    .A2(net4412));
 sg13g2_nand2_1 _17963_ (.Y(_02157_),
    .A(net2801),
    .B(net4412));
 sg13g2_o21ai_1 _17964_ (.B1(_02157_),
    .Y(_01584_),
    .A1(net5183),
    .A2(net4412));
 sg13g2_nand2_1 _17965_ (.Y(_02158_),
    .A(net2348),
    .B(net4413));
 sg13g2_o21ai_1 _17966_ (.B1(_02158_),
    .Y(_01585_),
    .A1(net5177),
    .A2(net4413));
 sg13g2_nand2_1 _17967_ (.Y(_02159_),
    .A(net2352),
    .B(net4414));
 sg13g2_o21ai_1 _17968_ (.B1(_02159_),
    .Y(_01586_),
    .A1(net5176),
    .A2(net4413));
 sg13g2_nand2_1 _17969_ (.Y(_02160_),
    .A(net2573),
    .B(net4410));
 sg13g2_o21ai_1 _17970_ (.B1(_02160_),
    .Y(_01587_),
    .A1(net5201),
    .A2(net4410));
 sg13g2_nand2_1 _17971_ (.Y(_02161_),
    .A(net2630),
    .B(net4410));
 sg13g2_o21ai_1 _17972_ (.B1(_02161_),
    .Y(_01588_),
    .A1(net5219),
    .A2(net4410));
 sg13g2_nand2_1 _17973_ (.Y(_02162_),
    .A(net2460),
    .B(net4414));
 sg13g2_o21ai_1 _17974_ (.B1(_02162_),
    .Y(_01589_),
    .A1(net5212),
    .A2(net4414));
 sg13g2_nand2_1 _17975_ (.Y(_02163_),
    .A(net2416),
    .B(net4410));
 sg13g2_o21ai_1 _17976_ (.B1(_02163_),
    .Y(_01590_),
    .A1(net5197),
    .A2(net4410));
 sg13g2_nand2_1 _17977_ (.Y(_02164_),
    .A(net2475),
    .B(net4407));
 sg13g2_o21ai_1 _17978_ (.B1(_02164_),
    .Y(_01591_),
    .A1(net5196),
    .A2(net4407));
 sg13g2_nand2_1 _17979_ (.Y(_02165_),
    .A(net2466),
    .B(net4411));
 sg13g2_o21ai_1 _17980_ (.B1(_02165_),
    .Y(_01592_),
    .A1(net5195),
    .A2(net4411));
 sg13g2_nand2_1 _17981_ (.Y(_02166_),
    .A(net2598),
    .B(net4406));
 sg13g2_o21ai_1 _17982_ (.B1(_02166_),
    .Y(_01593_),
    .A1(net5194),
    .A2(net4406));
 sg13g2_nand2_1 _17983_ (.Y(_02167_),
    .A(net2441),
    .B(net4406));
 sg13g2_o21ai_1 _17984_ (.B1(_02167_),
    .Y(_01594_),
    .A1(net5193),
    .A2(net4406));
 sg13g2_nand2_1 _17985_ (.Y(_02168_),
    .A(net2684),
    .B(net4407));
 sg13g2_o21ai_1 _17986_ (.B1(_02168_),
    .Y(_01595_),
    .A1(_02439_),
    .A2(net4407));
 sg13g2_nand2_1 _17987_ (.Y(_02169_),
    .A(net2456),
    .B(net4411));
 sg13g2_o21ai_1 _17988_ (.B1(_02169_),
    .Y(_01596_),
    .A1(net5192),
    .A2(net4411));
 sg13g2_nand2_1 _17989_ (.Y(_02170_),
    .A(net2837),
    .B(net4406));
 sg13g2_o21ai_1 _17990_ (.B1(_02170_),
    .Y(_01597_),
    .A1(_02443_),
    .A2(net4406));
 sg13g2_nand2_1 _17991_ (.Y(_02171_),
    .A(net2786),
    .B(net4406));
 sg13g2_o21ai_1 _17992_ (.B1(_02171_),
    .Y(_01598_),
    .A1(_02444_),
    .A2(net4406));
 sg13g2_a21oi_1 _17993_ (.A1(_02634_),
    .A2(_02753_),
    .Y(_02172_),
    .B1(net5309));
 sg13g2_nor2_1 _17994_ (.A(_02751_),
    .B(_02172_),
    .Y(_02173_));
 sg13g2_nor3_1 _17995_ (.A(\m_sys.m_core.m_fsm.r_cstate[3] ),
    .B(\m_sys.m_core.m_fsm.r_cstate[2] ),
    .C(net3263),
    .Y(_02174_));
 sg13g2_a221oi_1 _17996_ (.B2(_02752_),
    .C1(net5375),
    .B1(net3264),
    .A1(_01938_),
    .Y(_01599_),
    .A2(_02173_));
 sg13g2_nand2_1 _17997_ (.Y(_02175_),
    .A(\m_sys.m_core.m_gpr.io_b_write_addr[0] ),
    .B(_02055_));
 sg13g2_nand2_1 _17998_ (.Y(_02176_),
    .A(net2768),
    .B(net4372));
 sg13g2_o21ai_1 _17999_ (.B1(_02176_),
    .Y(_01600_),
    .A1(_02397_),
    .A2(net4372));
 sg13g2_mux2_1 _18000_ (.A0(net5312),
    .A1(net3130),
    .S(net4371),
    .X(_01601_));
 sg13g2_nand2_1 _18001_ (.Y(_02177_),
    .A(net2784),
    .B(net4371));
 sg13g2_o21ai_1 _18002_ (.B1(_02177_),
    .Y(_01602_),
    .A1(net5231),
    .A2(net4371));
 sg13g2_mux2_1 _18003_ (.A0(net5313),
    .A1(net3089),
    .S(net4376),
    .X(_01603_));
 sg13g2_mux2_1 _18004_ (.A0(net5316),
    .A1(net3127),
    .S(net4372),
    .X(_01604_));
 sg13g2_mux2_1 _18005_ (.A0(net5319),
    .A1(net3116),
    .S(net4372),
    .X(_01605_));
 sg13g2_nand2_1 _18006_ (.Y(_02178_),
    .A(net2646),
    .B(net4372));
 sg13g2_o21ai_1 _18007_ (.B1(_02178_),
    .Y(_01606_),
    .A1(net5226),
    .A2(net4372));
 sg13g2_nand2_1 _18008_ (.Y(_02179_),
    .A(net2503),
    .B(net4372));
 sg13g2_o21ai_1 _18009_ (.B1(_02179_),
    .Y(_01607_),
    .A1(net5227),
    .A2(net4371));
 sg13g2_mux2_1 _18010_ (.A0(net5320),
    .A1(net3106),
    .S(net4376),
    .X(_01608_));
 sg13g2_nand2_1 _18011_ (.Y(_02180_),
    .A(net2551),
    .B(net4371));
 sg13g2_o21ai_1 _18012_ (.B1(_02180_),
    .Y(_01609_),
    .A1(net5228),
    .A2(net4371));
 sg13g2_nand2_1 _18013_ (.Y(_02181_),
    .A(net2725),
    .B(net4371));
 sg13g2_o21ai_1 _18014_ (.B1(_02181_),
    .Y(_01610_),
    .A1(net5229),
    .A2(net4371));
 sg13g2_nand2_1 _18015_ (.Y(_02182_),
    .A(net2648),
    .B(net4375));
 sg13g2_o21ai_1 _18016_ (.B1(_02182_),
    .Y(_01611_),
    .A1(net5230),
    .A2(net4375));
 sg13g2_nand2_1 _18017_ (.Y(_02183_),
    .A(net2635),
    .B(net4373));
 sg13g2_o21ai_1 _18018_ (.B1(_02183_),
    .Y(_01612_),
    .A1(net5223),
    .A2(net4373));
 sg13g2_nand2_1 _18019_ (.Y(_02184_),
    .A(net2701),
    .B(net4375));
 sg13g2_o21ai_1 _18020_ (.B1(_02184_),
    .Y(_01613_),
    .A1(net5224),
    .A2(net4375));
 sg13g2_nand2_1 _18021_ (.Y(_02185_),
    .A(net2588),
    .B(net4376));
 sg13g2_o21ai_1 _18022_ (.B1(_02185_),
    .Y(_01614_),
    .A1(net5222),
    .A2(net4377));
 sg13g2_nand2_1 _18023_ (.Y(_02186_),
    .A(net2585),
    .B(net4377));
 sg13g2_o21ai_1 _18024_ (.B1(_02186_),
    .Y(_01615_),
    .A1(net5191),
    .A2(net4377));
 sg13g2_nand2_1 _18025_ (.Y(_02187_),
    .A(net2277),
    .B(net4376));
 sg13g2_o21ai_1 _18026_ (.B1(_02187_),
    .Y(_01616_),
    .A1(net5187),
    .A2(net4377));
 sg13g2_nand2_1 _18027_ (.Y(_02188_),
    .A(net2822),
    .B(net4373));
 sg13g2_o21ai_1 _18028_ (.B1(_02188_),
    .Y(_01617_),
    .A1(net5180),
    .A2(net4373));
 sg13g2_nand2_1 _18029_ (.Y(_02189_),
    .A(net2257),
    .B(net4376));
 sg13g2_o21ai_1 _18030_ (.B1(_02189_),
    .Y(_01618_),
    .A1(net5177),
    .A2(net4376));
 sg13g2_nand2_1 _18031_ (.Y(_02190_),
    .A(net2774),
    .B(net4376));
 sg13g2_o21ai_1 _18032_ (.B1(_02190_),
    .Y(_01619_),
    .A1(net5176),
    .A2(net4376));
 sg13g2_nand2_1 _18033_ (.Y(_02191_),
    .A(net2850),
    .B(net4373));
 sg13g2_o21ai_1 _18034_ (.B1(_02191_),
    .Y(_01620_),
    .A1(net5201),
    .A2(net4373));
 sg13g2_nand2_1 _18035_ (.Y(_02192_),
    .A(net2297),
    .B(net4374));
 sg13g2_o21ai_1 _18036_ (.B1(_02192_),
    .Y(_01621_),
    .A1(net5219),
    .A2(net4374));
 sg13g2_nand2_1 _18037_ (.Y(_02193_),
    .A(net2429),
    .B(net4374));
 sg13g2_o21ai_1 _18038_ (.B1(_02193_),
    .Y(_01622_),
    .A1(net5212),
    .A2(net4373));
 sg13g2_nand2_1 _18039_ (.Y(_02194_),
    .A(net2394),
    .B(net4373));
 sg13g2_o21ai_1 _18040_ (.B1(_02194_),
    .Y(_01623_),
    .A1(net5197),
    .A2(net4374));
 sg13g2_nand2_1 _18041_ (.Y(_02195_),
    .A(net2631),
    .B(net4370));
 sg13g2_o21ai_1 _18042_ (.B1(_02195_),
    .Y(_01624_),
    .A1(net5196),
    .A2(net4370));
 sg13g2_nand2_1 _18043_ (.Y(_02196_),
    .A(net2633),
    .B(net4370));
 sg13g2_o21ai_1 _18044_ (.B1(_02196_),
    .Y(_01625_),
    .A1(net5195),
    .A2(net4370));
 sg13g2_nand2_1 _18045_ (.Y(_02197_),
    .A(net2653),
    .B(net4369));
 sg13g2_o21ai_1 _18046_ (.B1(_02197_),
    .Y(_01626_),
    .A1(net5194),
    .A2(net4369));
 sg13g2_nand2_1 _18047_ (.Y(_02198_),
    .A(net2224),
    .B(net4369));
 sg13g2_o21ai_1 _18048_ (.B1(_02198_),
    .Y(_01627_),
    .A1(net5193),
    .A2(net4369));
 sg13g2_nand2_1 _18049_ (.Y(_02199_),
    .A(net2871),
    .B(net4370));
 sg13g2_o21ai_1 _18050_ (.B1(_02199_),
    .Y(_01628_),
    .A1(_02439_),
    .A2(net4370));
 sg13g2_nand2_1 _18051_ (.Y(_02200_),
    .A(net2507),
    .B(net4375));
 sg13g2_o21ai_1 _18052_ (.B1(_02200_),
    .Y(_01629_),
    .A1(net5192),
    .A2(net4375));
 sg13g2_nand2_1 _18053_ (.Y(_02201_),
    .A(net2473),
    .B(net4369));
 sg13g2_o21ai_1 _18054_ (.B1(_02201_),
    .Y(_01630_),
    .A1(_02443_),
    .A2(net4369));
 sg13g2_nand2_1 _18055_ (.Y(_02202_),
    .A(net2575),
    .B(net4369));
 sg13g2_o21ai_1 _18056_ (.B1(_02202_),
    .Y(_01631_),
    .A1(_02444_),
    .A2(net4369));
 sg13g2_nand2b_1 _18057_ (.Y(_02203_),
    .B(_02113_),
    .A_N(_07465_));
 sg13g2_nor2_1 _18058_ (.A(\m_sys.m_core.m_bru.io_i_s1[0] ),
    .B(net4397),
    .Y(_02204_));
 sg13g2_a21oi_1 _18059_ (.A1(_02486_),
    .A2(net4397),
    .Y(_01632_),
    .B1(_02204_));
 sg13g2_mux2_1 _18060_ (.A0(net5312),
    .A1(net3027),
    .S(net4398),
    .X(_01633_));
 sg13g2_nand2_1 _18061_ (.Y(_02205_),
    .A(net2740),
    .B(net4403));
 sg13g2_o21ai_1 _18062_ (.B1(_02205_),
    .Y(_01634_),
    .A1(net5231),
    .A2(net4403));
 sg13g2_nor2_1 _18063_ (.A(net5313),
    .B(net4403),
    .Y(_02206_));
 sg13g2_a21oi_1 _18064_ (.A1(_02429_),
    .A2(net4403),
    .Y(_01635_),
    .B1(_02206_));
 sg13g2_mux2_1 _18065_ (.A0(net5316),
    .A1(net3020),
    .S(net4398),
    .X(_01636_));
 sg13g2_nor2_1 _18066_ (.A(net5319),
    .B(net4395),
    .Y(_02207_));
 sg13g2_a21oi_1 _18067_ (.A1(_02433_),
    .A2(net4395),
    .Y(_01637_),
    .B1(_02207_));
 sg13g2_nor2_1 _18068_ (.A(\m_sys.m_core.m_bru.io_i_s1[6] ),
    .B(net4397),
    .Y(_02208_));
 sg13g2_a21oi_1 _18069_ (.A1(_02436_),
    .A2(net4397),
    .Y(_01638_),
    .B1(_02208_));
 sg13g2_nor2_1 _18070_ (.A(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[0] ),
    .B(net4398),
    .Y(_02209_));
 sg13g2_a21oi_1 _18071_ (.A1(_02438_),
    .A2(net4398),
    .Y(_01639_),
    .B1(_02209_));
 sg13g2_mux2_1 _18072_ (.A0(net5320),
    .A1(net3026),
    .S(net4402),
    .X(_01640_));
 sg13g2_nor2_1 _18073_ (.A(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[2] ),
    .B(net4397),
    .Y(_02210_));
 sg13g2_a21oi_1 _18074_ (.A1(_02441_),
    .A2(net4397),
    .Y(_01641_),
    .B1(_02210_));
 sg13g2_nand2_1 _18075_ (.Y(_02211_),
    .A(net2321),
    .B(net4397));
 sg13g2_o21ai_1 _18076_ (.B1(_02211_),
    .Y(_01642_),
    .A1(net5229),
    .A2(net4397));
 sg13g2_nand2_1 _18077_ (.Y(_02212_),
    .A(net2524),
    .B(net4402));
 sg13g2_o21ai_1 _18078_ (.B1(_02212_),
    .Y(_01643_),
    .A1(net5230),
    .A2(net4402));
 sg13g2_nand2_1 _18079_ (.Y(_02213_),
    .A(net2412),
    .B(net4400));
 sg13g2_o21ai_1 _18080_ (.B1(_02213_),
    .Y(_01644_),
    .A1(net5223),
    .A2(net4400));
 sg13g2_nand2_1 _18081_ (.Y(_02214_),
    .A(net2520),
    .B(net4402));
 sg13g2_o21ai_1 _18082_ (.B1(_02214_),
    .Y(_01645_),
    .A1(net5224),
    .A2(net4402));
 sg13g2_nand2_1 _18083_ (.Y(_02215_),
    .A(net2771),
    .B(net4400));
 sg13g2_o21ai_1 _18084_ (.B1(_02215_),
    .Y(_01646_),
    .A1(net5222),
    .A2(net4400));
 sg13g2_nand2_1 _18085_ (.Y(_02216_),
    .A(net2843),
    .B(net4404));
 sg13g2_o21ai_1 _18086_ (.B1(_02216_),
    .Y(_01647_),
    .A1(net5191),
    .A2(net4404));
 sg13g2_nand2_1 _18087_ (.Y(_02217_),
    .A(net2563),
    .B(net4404));
 sg13g2_o21ai_1 _18088_ (.B1(_02217_),
    .Y(_01648_),
    .A1(net5187),
    .A2(net4403));
 sg13g2_nand2_1 _18089_ (.Y(_02218_),
    .A(net2899),
    .B(net4404));
 sg13g2_o21ai_1 _18090_ (.B1(_02218_),
    .Y(_01649_),
    .A1(net5182),
    .A2(net4404));
 sg13g2_nand2_1 _18091_ (.Y(_02219_),
    .A(net2867),
    .B(net4403));
 sg13g2_o21ai_1 _18092_ (.B1(_02219_),
    .Y(_01650_),
    .A1(net5177),
    .A2(net4403));
 sg13g2_nand2_1 _18093_ (.Y(_02220_),
    .A(net2007),
    .B(net4404));
 sg13g2_o21ai_1 _18094_ (.B1(_02220_),
    .Y(_01651_),
    .A1(net5176),
    .A2(net4403));
 sg13g2_nand2_1 _18095_ (.Y(_02221_),
    .A(net2109),
    .B(net4400));
 sg13g2_o21ai_1 _18096_ (.B1(_02221_),
    .Y(_01652_),
    .A1(net5202),
    .A2(net4400));
 sg13g2_nor2_1 _18097_ (.A(net5350),
    .B(net4401),
    .Y(_02222_));
 sg13g2_a21oi_1 _18098_ (.A1(_02453_),
    .A2(net4401),
    .Y(_01653_),
    .B1(_02222_));
 sg13g2_nor2_1 _18099_ (.A(net5351),
    .B(net4401),
    .Y(_02223_));
 sg13g2_a21oi_1 _18100_ (.A1(_02454_),
    .A2(net4401),
    .Y(_01654_),
    .B1(_02223_));
 sg13g2_nand2_1 _18101_ (.Y(_02224_),
    .A(net2676),
    .B(net4400));
 sg13g2_o21ai_1 _18102_ (.B1(_02224_),
    .Y(_01655_),
    .A1(net5197),
    .A2(net4400));
 sg13g2_nand2_1 _18103_ (.Y(_02225_),
    .A(net2236),
    .B(net4395));
 sg13g2_o21ai_1 _18104_ (.B1(_02225_),
    .Y(_01656_),
    .A1(net5196),
    .A2(net4395));
 sg13g2_nand2_1 _18105_ (.Y(_02226_),
    .A(net2541),
    .B(net4395));
 sg13g2_o21ai_1 _18106_ (.B1(_02226_),
    .Y(_01657_),
    .A1(net5195),
    .A2(net4395));
 sg13g2_nand2_1 _18107_ (.Y(_02227_),
    .A(net2262),
    .B(net4396));
 sg13g2_o21ai_1 _18108_ (.B1(_02227_),
    .Y(_01658_),
    .A1(net5194),
    .A2(net4396));
 sg13g2_nand2_1 _18109_ (.Y(_02228_),
    .A(net2552),
    .B(net4396));
 sg13g2_o21ai_1 _18110_ (.B1(_02228_),
    .Y(_01659_),
    .A1(net5193),
    .A2(net4399));
 sg13g2_nand2_1 _18111_ (.Y(_02229_),
    .A(net1964),
    .B(net4395));
 sg13g2_o21ai_1 _18112_ (.B1(_02229_),
    .Y(_01660_),
    .A1(_02439_),
    .A2(net4395));
 sg13g2_nand2_1 _18113_ (.Y(_02230_),
    .A(net2232),
    .B(net4402));
 sg13g2_o21ai_1 _18114_ (.B1(_02230_),
    .Y(_01661_),
    .A1(net5192),
    .A2(net4402));
 sg13g2_nor2_1 _18115_ (.A(\m_sys.m_core.m_bru.io_i_s1[30] ),
    .B(net4396),
    .Y(_02231_));
 sg13g2_a21oi_1 _18116_ (.A1(_02456_),
    .A2(net4396),
    .Y(_01662_),
    .B1(_02231_));
 sg13g2_nor2_1 _18117_ (.A(net5353),
    .B(net4396),
    .Y(_02232_));
 sg13g2_a21oi_1 _18118_ (.A1(_02457_),
    .A2(net4396),
    .Y(_01663_),
    .B1(_02232_));
 sg13g2_nor2b_1 _18119_ (.A(net4333),
    .B_N(_05848_),
    .Y(_02233_));
 sg13g2_nor2_1 _18120_ (.A(net2444),
    .B(net4059),
    .Y(_02234_));
 sg13g2_a21oi_1 _18121_ (.A1(net5136),
    .A2(net4059),
    .Y(_01664_),
    .B1(_02234_));
 sg13g2_nor2_1 _18122_ (.A(net2241),
    .B(net4060),
    .Y(_02235_));
 sg13g2_a21oi_1 _18123_ (.A1(net4997),
    .A2(net4060),
    .Y(_01665_),
    .B1(_02235_));
 sg13g2_nor2_1 _18124_ (.A(net2173),
    .B(net4059),
    .Y(_02236_));
 sg13g2_a21oi_1 _18125_ (.A1(net5133),
    .A2(net4059),
    .Y(_01666_),
    .B1(_02236_));
 sg13g2_nor2_1 _18126_ (.A(net2246),
    .B(net4060),
    .Y(_02237_));
 sg13g2_a21oi_1 _18127_ (.A1(net4990),
    .A2(net4060),
    .Y(_01667_),
    .B1(_02237_));
 sg13g2_nor2_1 _18128_ (.A(net2375),
    .B(net4059),
    .Y(_02238_));
 sg13g2_a21oi_1 _18129_ (.A1(net5129),
    .A2(net4059),
    .Y(_01668_),
    .B1(_02238_));
 sg13g2_nor2_1 _18130_ (.A(net2196),
    .B(net4059),
    .Y(_02239_));
 sg13g2_a21oi_1 _18131_ (.A1(net4984),
    .A2(net4059),
    .Y(_01669_),
    .B1(_02239_));
 sg13g2_nor2_1 _18132_ (.A(net2500),
    .B(net4060),
    .Y(_02240_));
 sg13g2_a21oi_1 _18133_ (.A1(net5123),
    .A2(net4060),
    .Y(_01670_),
    .B1(_02240_));
 sg13g2_nor2_1 _18134_ (.A(net2248),
    .B(net4060),
    .Y(_02241_));
 sg13g2_a21oi_1 _18135_ (.A1(net4981),
    .A2(net4060),
    .Y(_01671_),
    .B1(_02241_));
 sg13g2_nand2_1 _18136_ (.Y(_02242_),
    .A(net4328),
    .B(_05802_));
 sg13g2_nand2_1 _18137_ (.Y(_02243_),
    .A(net1732),
    .B(_02242_));
 sg13g2_o21ai_1 _18138_ (.B1(_02243_),
    .Y(_01672_),
    .A1(net5043),
    .A2(net4057));
 sg13g2_nand2_1 _18139_ (.Y(_02244_),
    .A(net1769),
    .B(net4058));
 sg13g2_o21ai_1 _18140_ (.B1(_02244_),
    .Y(_01673_),
    .A1(net4875),
    .A2(net4058));
 sg13g2_nand2_1 _18141_ (.Y(_02245_),
    .A(net1694),
    .B(net4057));
 sg13g2_o21ai_1 _18142_ (.B1(_02245_),
    .Y(_01674_),
    .A1(net5038),
    .A2(net4057));
 sg13g2_nand2_1 _18143_ (.Y(_02246_),
    .A(net1924),
    .B(net4057));
 sg13g2_o21ai_1 _18144_ (.B1(_02246_),
    .Y(_01675_),
    .A1(net4871),
    .A2(net4058));
 sg13g2_nand2_1 _18145_ (.Y(_02247_),
    .A(net1940),
    .B(net4057));
 sg13g2_o21ai_1 _18146_ (.B1(_02247_),
    .Y(_01676_),
    .A1(net5032),
    .A2(net4057));
 sg13g2_nand2_1 _18147_ (.Y(_02248_),
    .A(net1789),
    .B(net4057));
 sg13g2_o21ai_1 _18148_ (.B1(_02248_),
    .Y(_01677_),
    .A1(net4866),
    .A2(net4057));
 sg13g2_nand2_1 _18149_ (.Y(_02249_),
    .A(net2000),
    .B(net4058));
 sg13g2_o21ai_1 _18150_ (.B1(_02249_),
    .Y(_01678_),
    .A1(net5027),
    .A2(net4058));
 sg13g2_nand2_1 _18151_ (.Y(_02250_),
    .A(net1914),
    .B(net4058));
 sg13g2_o21ai_1 _18152_ (.B1(_02250_),
    .Y(_01679_),
    .A1(net4859),
    .A2(net4058));
 sg13g2_nand2_1 _18153_ (.Y(_02251_),
    .A(net4323),
    .B(_05848_));
 sg13g2_nand2_1 _18154_ (.Y(_02252_),
    .A(net2227),
    .B(_02251_));
 sg13g2_o21ai_1 _18155_ (.B1(_02252_),
    .Y(_01680_),
    .A1(net4856),
    .A2(net4056));
 sg13g2_nand2_1 _18156_ (.Y(_02253_),
    .A(net1713),
    .B(net4055));
 sg13g2_o21ai_1 _18157_ (.B1(_02253_),
    .Y(_01681_),
    .A1(net4849),
    .A2(net4055));
 sg13g2_nand2_1 _18158_ (.Y(_02254_),
    .A(net1978),
    .B(net4056));
 sg13g2_o21ai_1 _18159_ (.B1(_02254_),
    .Y(_01682_),
    .A1(net4846),
    .A2(net4056));
 sg13g2_nand2_1 _18160_ (.Y(_02255_),
    .A(net1715),
    .B(net4056));
 sg13g2_o21ai_1 _18161_ (.B1(_02255_),
    .Y(_01683_),
    .A1(net4840),
    .A2(net4055));
 sg13g2_nand2_1 _18162_ (.Y(_02256_),
    .A(net1664),
    .B(net4056));
 sg13g2_o21ai_1 _18163_ (.B1(_02256_),
    .Y(_01684_),
    .A1(net4834),
    .A2(net4056));
 sg13g2_nand2_1 _18164_ (.Y(_02257_),
    .A(net1976),
    .B(net4055));
 sg13g2_o21ai_1 _18165_ (.B1(_02257_),
    .Y(_01685_),
    .A1(net4827),
    .A2(net4055));
 sg13g2_nand2_1 _18166_ (.Y(_02258_),
    .A(net1922),
    .B(net4056));
 sg13g2_o21ai_1 _18167_ (.B1(_02258_),
    .Y(_01686_),
    .A1(net4823),
    .A2(net4055));
 sg13g2_nand2_1 _18168_ (.Y(_02259_),
    .A(net2222),
    .B(net4055));
 sg13g2_o21ai_1 _18169_ (.B1(_02259_),
    .Y(_01687_),
    .A1(net4818),
    .A2(net4055));
 sg13g2_nand2_1 _18170_ (.Y(_02260_),
    .A(net4323),
    .B(_05802_));
 sg13g2_nand2_1 _18171_ (.Y(_02261_),
    .A(net1771),
    .B(net4054));
 sg13g2_o21ai_1 _18172_ (.B1(_02261_),
    .Y(_01688_),
    .A1(net4856),
    .A2(net4054));
 sg13g2_nand2_1 _18173_ (.Y(_02262_),
    .A(net2019),
    .B(net4053));
 sg13g2_o21ai_1 _18174_ (.B1(_02262_),
    .Y(_01689_),
    .A1(net4849),
    .A2(net4053));
 sg13g2_nand2_1 _18175_ (.Y(_02263_),
    .A(net1974),
    .B(net4054));
 sg13g2_o21ai_1 _18176_ (.B1(_02263_),
    .Y(_01690_),
    .A1(net4846),
    .A2(net4054));
 sg13g2_nand2_1 _18177_ (.Y(_02264_),
    .A(net1916),
    .B(net4053));
 sg13g2_o21ai_1 _18178_ (.B1(_02264_),
    .Y(_01691_),
    .A1(net4840),
    .A2(net4053));
 sg13g2_nand2_1 _18179_ (.Y(_02265_),
    .A(net2001),
    .B(net4054));
 sg13g2_o21ai_1 _18180_ (.B1(_02265_),
    .Y(_01692_),
    .A1(net4834),
    .A2(net4054));
 sg13g2_nand2_1 _18181_ (.Y(_02266_),
    .A(net1970),
    .B(net4053));
 sg13g2_o21ai_1 _18182_ (.B1(_02266_),
    .Y(_01693_),
    .A1(net4827),
    .A2(net4053));
 sg13g2_nand2_1 _18183_ (.Y(_02267_),
    .A(net2133),
    .B(net4054));
 sg13g2_o21ai_1 _18184_ (.B1(_02267_),
    .Y(_01694_),
    .A1(net4823),
    .A2(net4054));
 sg13g2_nand2_1 _18185_ (.Y(_02268_),
    .A(net1763),
    .B(net4053));
 sg13g2_o21ai_1 _18186_ (.B1(_02268_),
    .Y(_01695_),
    .A1(net4818),
    .A2(net4053));
 sg13g2_nor2b_1 _18187_ (.A(net4333),
    .B_N(_05802_),
    .Y(_02269_));
 sg13g2_nor2_1 _18188_ (.A(net2186),
    .B(net4051),
    .Y(_02270_));
 sg13g2_a21oi_1 _18189_ (.A1(net5136),
    .A2(net4051),
    .Y(_01696_),
    .B1(_02270_));
 sg13g2_nor2_1 _18190_ (.A(net2234),
    .B(net4052),
    .Y(_02271_));
 sg13g2_a21oi_1 _18191_ (.A1(net4997),
    .A2(net4052),
    .Y(_01697_),
    .B1(_02271_));
 sg13g2_nor2_1 _18192_ (.A(net2482),
    .B(net4052),
    .Y(_02272_));
 sg13g2_a21oi_1 _18193_ (.A1(net5133),
    .A2(net4052),
    .Y(_01698_),
    .B1(_02272_));
 sg13g2_nor2_1 _18194_ (.A(net2735),
    .B(net4051),
    .Y(_02273_));
 sg13g2_a21oi_1 _18195_ (.A1(net4990),
    .A2(net4051),
    .Y(_01699_),
    .B1(_02273_));
 sg13g2_nor2_1 _18196_ (.A(net2733),
    .B(net4051),
    .Y(_02274_));
 sg13g2_a21oi_1 _18197_ (.A1(net5129),
    .A2(net4051),
    .Y(_01700_),
    .B1(_02274_));
 sg13g2_nor2_1 _18198_ (.A(net2181),
    .B(net4051),
    .Y(_02275_));
 sg13g2_a21oi_1 _18199_ (.A1(net4984),
    .A2(net4051),
    .Y(_01701_),
    .B1(_02275_));
 sg13g2_nor2_1 _18200_ (.A(net2420),
    .B(_02269_),
    .Y(_02276_));
 sg13g2_a21oi_1 _18201_ (.A1(net5123),
    .A2(net4052),
    .Y(_01702_),
    .B1(_02276_));
 sg13g2_nor2_1 _18202_ (.A(net2594),
    .B(net4052),
    .Y(_02277_));
 sg13g2_a21oi_1 _18203_ (.A1(net4981),
    .A2(net4052),
    .Y(_01703_),
    .B1(_02277_));
 sg13g2_nand2_1 _18204_ (.Y(_02278_),
    .A(net4328),
    .B(_07400_));
 sg13g2_nand2_1 _18205_ (.Y(_02279_),
    .A(net1957),
    .B(net4050));
 sg13g2_o21ai_1 _18206_ (.B1(_02279_),
    .Y(_01704_),
    .A1(net5043),
    .A2(net4050));
 sg13g2_nand2_1 _18207_ (.Y(_02280_),
    .A(net1968),
    .B(net4049));
 sg13g2_o21ai_1 _18208_ (.B1(_02280_),
    .Y(_01705_),
    .A1(net4875),
    .A2(net4049));
 sg13g2_nand2_1 _18209_ (.Y(_02281_),
    .A(net2245),
    .B(net4050));
 sg13g2_o21ai_1 _18210_ (.B1(_02281_),
    .Y(_01706_),
    .A1(net5038),
    .A2(net4050));
 sg13g2_nand2_1 _18211_ (.Y(_02282_),
    .A(net1835),
    .B(net4049));
 sg13g2_o21ai_1 _18212_ (.B1(_02282_),
    .Y(_01707_),
    .A1(net4871),
    .A2(net4049));
 sg13g2_nand2_1 _18213_ (.Y(_02283_),
    .A(net1850),
    .B(net4050));
 sg13g2_o21ai_1 _18214_ (.B1(_02283_),
    .Y(_01708_),
    .A1(net5032),
    .A2(net4050));
 sg13g2_nand2_1 _18215_ (.Y(_02284_),
    .A(net1822),
    .B(net4050));
 sg13g2_o21ai_1 _18216_ (.B1(_02284_),
    .Y(_01709_),
    .A1(net4866),
    .A2(net4050));
 sg13g2_nand2_1 _18217_ (.Y(_02285_),
    .A(net2039),
    .B(net4049));
 sg13g2_o21ai_1 _18218_ (.B1(_02285_),
    .Y(_01710_),
    .A1(net5026),
    .A2(net4049));
 sg13g2_nand2_1 _18219_ (.Y(_02286_),
    .A(net2281),
    .B(net4049));
 sg13g2_o21ai_1 _18220_ (.B1(_02286_),
    .Y(_01711_),
    .A1(net4859),
    .A2(net4049));
 sg13g2_nand2_1 _18221_ (.Y(_02287_),
    .A(net4323),
    .B(_07400_));
 sg13g2_nand2_1 _18222_ (.Y(_02288_),
    .A(net2207),
    .B(net4047));
 sg13g2_o21ai_1 _18223_ (.B1(_02288_),
    .Y(_01712_),
    .A1(net4856),
    .A2(net4047));
 sg13g2_nand2_1 _18224_ (.Y(_02289_),
    .A(net2178),
    .B(net4048));
 sg13g2_o21ai_1 _18225_ (.B1(_02289_),
    .Y(_01713_),
    .A1(net4849),
    .A2(net4048));
 sg13g2_nand2_1 _18226_ (.Y(_02290_),
    .A(net2070),
    .B(net4047));
 sg13g2_o21ai_1 _18227_ (.B1(_02290_),
    .Y(_01714_),
    .A1(net4846),
    .A2(net4047));
 sg13g2_nand2_1 _18228_ (.Y(_02291_),
    .A(net1876),
    .B(net4048));
 sg13g2_o21ai_1 _18229_ (.B1(_02291_),
    .Y(_01715_),
    .A1(net4840),
    .A2(net4048));
 sg13g2_nand2_1 _18230_ (.Y(_02292_),
    .A(net2324),
    .B(_02287_));
 sg13g2_o21ai_1 _18231_ (.B1(_02292_),
    .Y(_01716_),
    .A1(net4834),
    .A2(net4047));
 sg13g2_nand2_1 _18232_ (.Y(_02293_),
    .A(net2142),
    .B(net4048));
 sg13g2_o21ai_1 _18233_ (.B1(_02293_),
    .Y(_01717_),
    .A1(net4827),
    .A2(net4048));
 sg13g2_nand2_1 _18234_ (.Y(_02294_),
    .A(net2089),
    .B(net4047));
 sg13g2_o21ai_1 _18235_ (.B1(_02294_),
    .Y(_01718_),
    .A1(net4823),
    .A2(net4047));
 sg13g2_nand2_1 _18236_ (.Y(_02295_),
    .A(net2153),
    .B(net4047));
 sg13g2_o21ai_1 _18237_ (.B1(_02295_),
    .Y(_01719_),
    .A1(net4818),
    .A2(net4048));
 sg13g2_nor2b_1 _18238_ (.A(net4333),
    .B_N(_07400_),
    .Y(_02296_));
 sg13g2_nor2_1 _18239_ (.A(net2694),
    .B(net4045),
    .Y(_02297_));
 sg13g2_a21oi_1 _18240_ (.A1(net5136),
    .A2(net4045),
    .Y(_01720_),
    .B1(_02297_));
 sg13g2_nor2_1 _18241_ (.A(net2577),
    .B(net4046),
    .Y(_02298_));
 sg13g2_a21oi_1 _18242_ (.A1(net4997),
    .A2(net4046),
    .Y(_01721_),
    .B1(_02298_));
 sg13g2_nor2_1 _18243_ (.A(net2439),
    .B(net4045),
    .Y(_02299_));
 sg13g2_a21oi_1 _18244_ (.A1(net5133),
    .A2(net4045),
    .Y(_01722_),
    .B1(_02299_));
 sg13g2_nor2_1 _18245_ (.A(net2805),
    .B(net4046),
    .Y(_02300_));
 sg13g2_a21oi_1 _18246_ (.A1(net4990),
    .A2(net4046),
    .Y(_01723_),
    .B1(_02300_));
 sg13g2_nor2_1 _18247_ (.A(net2302),
    .B(net4045),
    .Y(_02301_));
 sg13g2_a21oi_1 _18248_ (.A1(net5128),
    .A2(net4045),
    .Y(_01724_),
    .B1(_02301_));
 sg13g2_nor2_1 _18249_ (.A(net2728),
    .B(net4045),
    .Y(_02302_));
 sg13g2_a21oi_1 _18250_ (.A1(net4984),
    .A2(net4045),
    .Y(_01725_),
    .B1(_02302_));
 sg13g2_nor2_1 _18251_ (.A(net2204),
    .B(net4046),
    .Y(_02303_));
 sg13g2_a21oi_1 _18252_ (.A1(net5123),
    .A2(net4046),
    .Y(_01726_),
    .B1(_02303_));
 sg13g2_nor2_1 _18253_ (.A(net2611),
    .B(net4046),
    .Y(_02304_));
 sg13g2_a21oi_1 _18254_ (.A1(net4981),
    .A2(net4046),
    .Y(_01727_),
    .B1(_02304_));
 sg13g2_nand2_1 _18255_ (.Y(_02305_),
    .A(net4327),
    .B(_05867_));
 sg13g2_nand2_1 _18256_ (.Y(_02306_),
    .A(net1748),
    .B(net4044));
 sg13g2_o21ai_1 _18257_ (.B1(_02306_),
    .Y(_01728_),
    .A1(net5041),
    .A2(net4044));
 sg13g2_nand2_1 _18258_ (.Y(_02307_),
    .A(net2115),
    .B(net4043));
 sg13g2_o21ai_1 _18259_ (.B1(_02307_),
    .Y(_01729_),
    .A1(net4876),
    .A2(net4043));
 sg13g2_nand2_1 _18260_ (.Y(_02308_),
    .A(net1745),
    .B(net4044));
 sg13g2_o21ai_1 _18261_ (.B1(_02308_),
    .Y(_01730_),
    .A1(net5037),
    .A2(net4044));
 sg13g2_nand2_1 _18262_ (.Y(_02309_),
    .A(net1818),
    .B(net4043));
 sg13g2_o21ai_1 _18263_ (.B1(_02309_),
    .Y(_01731_),
    .A1(net4873),
    .A2(net4043));
 sg13g2_nand2_1 _18264_ (.Y(_02310_),
    .A(net2041),
    .B(net4043));
 sg13g2_o21ai_1 _18265_ (.B1(_02310_),
    .Y(_01732_),
    .A1(net5034),
    .A2(net4043));
 sg13g2_nand2_1 _18266_ (.Y(_02311_),
    .A(net1668),
    .B(net4044));
 sg13g2_o21ai_1 _18267_ (.B1(_02311_),
    .Y(_01733_),
    .A1(net4865),
    .A2(net4044));
 sg13g2_nand2_1 _18268_ (.Y(_02312_),
    .A(net1661),
    .B(net4043));
 sg13g2_o21ai_1 _18269_ (.B1(_02312_),
    .Y(_01734_),
    .A1(net5028),
    .A2(net4043));
 sg13g2_nand2_1 _18270_ (.Y(_02313_),
    .A(net2064),
    .B(_02305_));
 sg13g2_o21ai_1 _18271_ (.B1(_02313_),
    .Y(_01735_),
    .A1(net4862),
    .A2(net4044));
 sg13g2_nand2_1 _18272_ (.Y(_02314_),
    .A(net4322),
    .B(_05867_));
 sg13g2_nand2_1 _18273_ (.Y(_02315_),
    .A(net1703),
    .B(net4041));
 sg13g2_o21ai_1 _18274_ (.B1(_02315_),
    .Y(_01736_),
    .A1(net4855),
    .A2(net4041));
 sg13g2_nand2_1 _18275_ (.Y(_02316_),
    .A(net1917),
    .B(net4042));
 sg13g2_o21ai_1 _18276_ (.B1(_02316_),
    .Y(_01737_),
    .A1(net4851),
    .A2(net4042));
 sg13g2_nand2_1 _18277_ (.Y(_02317_),
    .A(net2082),
    .B(net4042));
 sg13g2_o21ai_1 _18278_ (.B1(_02317_),
    .Y(_01738_),
    .A1(net4845),
    .A2(net4042));
 sg13g2_nand2_1 _18279_ (.Y(_02318_),
    .A(net1951),
    .B(net4042));
 sg13g2_o21ai_1 _18280_ (.B1(_02318_),
    .Y(_01739_),
    .A1(net4839),
    .A2(net4042));
 sg13g2_nand2_1 _18281_ (.Y(_02319_),
    .A(net1730),
    .B(net4041));
 sg13g2_o21ai_1 _18282_ (.B1(_02319_),
    .Y(_01740_),
    .A1(net4833),
    .A2(net4041));
 sg13g2_nand2_1 _18283_ (.Y(_02320_),
    .A(net1864),
    .B(net4042));
 sg13g2_o21ai_1 _18284_ (.B1(_02320_),
    .Y(_01741_),
    .A1(net4829),
    .A2(net4042));
 sg13g2_nand2_1 _18285_ (.Y(_02321_),
    .A(net1699),
    .B(net4041));
 sg13g2_o21ai_1 _18286_ (.B1(_02321_),
    .Y(_01742_),
    .A1(net4820),
    .A2(net4041));
 sg13g2_nand2_1 _18287_ (.Y(_02322_),
    .A(net1854),
    .B(net4041));
 sg13g2_o21ai_1 _18288_ (.B1(_02322_),
    .Y(_01743_),
    .A1(net4819),
    .A2(net4041));
 sg13g2_dfrbp_1 _18289_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1066),
    .D(_00147_),
    .Q_N(_09107_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[8] ));
 sg13g2_dfrbp_1 _18290_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net441),
    .D(_00148_),
    .Q_N(_09106_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[9] ));
 sg13g2_dfrbp_1 _18291_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net440),
    .D(_00149_),
    .Q_N(_09105_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[10] ));
 sg13g2_dfrbp_1 _18292_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net439),
    .D(_00150_),
    .Q_N(_09104_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[11] ));
 sg13g2_dfrbp_1 _18293_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net438),
    .D(_00151_),
    .Q_N(_00137_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[12] ));
 sg13g2_dfrbp_1 _18294_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net437),
    .D(_00152_),
    .Q_N(_00139_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[13] ));
 sg13g2_dfrbp_1 _18295_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net436),
    .D(_00153_),
    .Q_N(_00141_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[14] ));
 sg13g2_dfrbp_1 _18296_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net435),
    .D(_00154_),
    .Q_N(_00143_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[15] ));
 sg13g2_dfrbp_1 _18297_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net434),
    .D(net2459),
    .Q_N(_09103_),
    .Q(\m_sys._GEN_11[3] ));
 sg13g2_dfrbp_1 _18298_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net432),
    .D(_00156_),
    .Q_N(_00047_),
    .Q(\m_sys._GEN_11[4] ));
 sg13g2_dfrbp_1 _18299_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net430),
    .D(_00157_),
    .Q_N(_09102_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][16] ));
 sg13g2_dfrbp_1 _18300_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net429),
    .D(_00158_),
    .Q_N(_09101_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][17] ));
 sg13g2_dfrbp_1 _18301_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net428),
    .D(_00159_),
    .Q_N(_09100_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][18] ));
 sg13g2_dfrbp_1 _18302_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net427),
    .D(_00160_),
    .Q_N(_09099_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][19] ));
 sg13g2_dfrbp_1 _18303_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net426),
    .D(_00161_),
    .Q_N(_09098_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][20] ));
 sg13g2_dfrbp_1 _18304_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net425),
    .D(_00162_),
    .Q_N(_09097_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][21] ));
 sg13g2_dfrbp_1 _18305_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net424),
    .D(_00163_),
    .Q_N(_09096_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][22] ));
 sg13g2_dfrbp_1 _18306_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net423),
    .D(_00164_),
    .Q_N(_09095_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][23] ));
 sg13g2_dfrbp_1 _18307_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net422),
    .D(net3321),
    .Q_N(_00120_),
    .Q(\m_sys._m_core_io_b_mem_wdata[1] ));
 sg13g2_dfrbp_1 _18308_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net420),
    .D(net3437),
    .Q_N(_00117_),
    .Q(\m_sys._m_core_io_b_mem_wdata[2] ));
 sg13g2_dfrbp_1 _18309_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net418),
    .D(net3301),
    .Q_N(_00116_),
    .Q(\m_sys._m_core_io_b_mem_wdata[3] ));
 sg13g2_dfrbp_1 _18310_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net416),
    .D(_00168_),
    .Q_N(_00115_),
    .Q(\m_sys._m_core_io_b_mem_wdata[4] ));
 sg13g2_dfrbp_1 _18311_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net414),
    .D(net3129),
    .Q_N(_00114_),
    .Q(\m_sys._m_core_io_b_mem_wdata[5] ));
 sg13g2_dfrbp_1 _18312_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net412),
    .D(_00170_),
    .Q_N(_00112_),
    .Q(\m_sys._m_core_io_b_mem_wdata[6] ));
 sg13g2_dfrbp_1 _18313_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net410),
    .D(net3361),
    .Q_N(_09094_),
    .Q(\m_sys._m_core_io_b_mem_wdata[7] ));
 sg13g2_dfrbp_1 _18314_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net408),
    .D(net1800),
    .Q_N(_09093_),
    .Q(\m_sys._m_core_io_b_mem_wdata[8] ));
 sg13g2_dfrbp_1 _18315_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net406),
    .D(net2472),
    .Q_N(_00107_),
    .Q(\m_sys._m_core_io_b_mem_wdata[9] ));
 sg13g2_dfrbp_1 _18316_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net404),
    .D(net1656),
    .Q_N(_00104_),
    .Q(\m_sys._m_core_io_b_mem_wdata[10] ));
 sg13g2_dfrbp_1 _18317_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net402),
    .D(net3167),
    .Q_N(_00101_),
    .Q(\m_sys._m_core_io_b_mem_wdata[11] ));
 sg13g2_dfrbp_1 _18318_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net400),
    .D(net3290),
    .Q_N(_00099_),
    .Q(\m_sys._m_core_io_b_mem_wdata[12] ));
 sg13g2_dfrbp_1 _18319_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net398),
    .D(net3094),
    .Q_N(_00098_),
    .Q(\m_sys._m_core_io_b_mem_wdata[13] ));
 sg13g2_dfrbp_1 _18320_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net396),
    .D(net3157),
    .Q_N(_00097_),
    .Q(\m_sys._m_core_io_b_mem_wdata[14] ));
 sg13g2_dfrbp_1 _18321_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net394),
    .D(_00179_),
    .Q_N(_00096_),
    .Q(\m_sys._m_core_io_b_mem_wdata[15] ));
 sg13g2_dfrbp_1 _18322_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net392),
    .D(net2991),
    .Q_N(_00095_),
    .Q(\m_sys._m_core_io_b_mem_wdata[16] ));
 sg13g2_dfrbp_1 _18323_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net390),
    .D(net3378),
    .Q_N(_00094_),
    .Q(\m_sys._m_core_io_b_mem_wdata[17] ));
 sg13g2_dfrbp_1 _18324_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net388),
    .D(net3241),
    .Q_N(_00093_),
    .Q(\m_sys._m_core_io_b_mem_wdata[18] ));
 sg13g2_dfrbp_1 _18325_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net386),
    .D(net3395),
    .Q_N(_00092_),
    .Q(\m_sys._m_core_io_b_mem_wdata[19] ));
 sg13g2_dfrbp_1 _18326_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net384),
    .D(_00184_),
    .Q_N(_00091_),
    .Q(\m_sys._m_core_io_b_mem_wdata[20] ));
 sg13g2_dfrbp_1 _18327_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net382),
    .D(_00185_),
    .Q_N(_00090_),
    .Q(\m_sys._m_core_io_b_mem_wdata[21] ));
 sg13g2_dfrbp_1 _18328_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net380),
    .D(_00186_),
    .Q_N(_09092_),
    .Q(\m_sys._m_core_io_b_mem_wdata[22] ));
 sg13g2_dfrbp_1 _18329_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net378),
    .D(_00187_),
    .Q_N(_09091_),
    .Q(\m_sys._m_core_io_b_mem_wdata[23] ));
 sg13g2_dfrbp_1 _18330_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net376),
    .D(_00188_),
    .Q_N(_09090_),
    .Q(\m_sys._m_core_io_b_mem_wdata[24] ));
 sg13g2_dfrbp_1 _18331_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net374),
    .D(_00189_),
    .Q_N(_09089_),
    .Q(\m_sys._m_core_io_b_mem_wdata[25] ));
 sg13g2_dfrbp_1 _18332_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net372),
    .D(_00190_),
    .Q_N(_09088_),
    .Q(\m_sys._m_core_io_b_mem_wdata[26] ));
 sg13g2_dfrbp_1 _18333_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net370),
    .D(_00191_),
    .Q_N(_09087_),
    .Q(\m_sys._m_core_io_b_mem_wdata[27] ));
 sg13g2_dfrbp_1 _18334_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net368),
    .D(_00192_),
    .Q_N(_09086_),
    .Q(\m_sys._m_core_io_b_mem_wdata[28] ));
 sg13g2_dfrbp_1 _18335_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net366),
    .D(_00193_),
    .Q_N(_09085_),
    .Q(\m_sys._m_core_io_b_mem_wdata[29] ));
 sg13g2_dfrbp_1 _18336_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net364),
    .D(_00194_),
    .Q_N(_09084_),
    .Q(\m_sys._m_core_io_b_mem_wdata[30] ));
 sg13g2_dfrbp_1 _18337_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net362),
    .D(_00195_),
    .Q_N(_09083_),
    .Q(\m_sys._m_core_io_b_mem_wdata[31] ));
 sg13g2_dfrbp_1 _18338_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net360),
    .D(_00196_),
    .Q_N(_00080_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[31] ));
 sg13g2_dfrbp_1 _18339_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net359),
    .D(_00197_),
    .Q_N(_00077_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[30] ));
 sg13g2_dfrbp_1 _18340_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net358),
    .D(_00198_),
    .Q_N(_00076_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[29] ));
 sg13g2_dfrbp_1 _18341_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net357),
    .D(_00199_),
    .Q_N(_00075_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[28] ));
 sg13g2_dfrbp_1 _18342_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net356),
    .D(_00200_),
    .Q_N(_00074_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[27] ));
 sg13g2_dfrbp_1 _18343_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net355),
    .D(_00201_),
    .Q_N(_00073_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[26] ));
 sg13g2_dfrbp_1 _18344_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net354),
    .D(_00202_),
    .Q_N(_00072_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[25] ));
 sg13g2_dfrbp_1 _18345_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net353),
    .D(_00203_),
    .Q_N(_00071_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[24] ));
 sg13g2_dfrbp_1 _18346_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net352),
    .D(_00204_),
    .Q_N(_00069_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[23] ));
 sg13g2_dfrbp_1 _18347_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net351),
    .D(_00205_),
    .Q_N(_00067_),
    .Q(\m_sys.m_core._m_decoder_io_o_rs2[2] ));
 sg13g2_dfrbp_1 _18348_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net350),
    .D(_00206_),
    .Q_N(_00065_),
    .Q(\m_sys.m_core._m_decoder_io_o_rs2[1] ));
 sg13g2_dfrbp_1 _18349_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net349),
    .D(_00207_),
    .Q_N(_00078_),
    .Q(\m_sys.m_core._m_decoder_io_o_rs2[0] ));
 sg13g2_dfrbp_1 _18350_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net348),
    .D(_00208_),
    .Q_N(_00086_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[19] ));
 sg13g2_dfrbp_1 _18351_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net347),
    .D(_00209_),
    .Q_N(_00085_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[18] ));
 sg13g2_dfrbp_1 _18352_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net346),
    .D(_00210_),
    .Q_N(_00084_),
    .Q(\m_sys.m_core._m_decoder_io_o_rs1[2] ));
 sg13g2_dfrbp_1 _18353_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net345),
    .D(_00211_),
    .Q_N(_00083_),
    .Q(\m_sys.m_core._m_decoder_io_o_rs1[1] ));
 sg13g2_dfrbp_1 _18354_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net344),
    .D(_00212_),
    .Q_N(_00082_),
    .Q(\m_sys.m_core._m_decoder_io_o_rs1[0] ));
 sg13g2_dfrbp_1 _18355_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net343),
    .D(_00213_),
    .Q_N(_00026_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[14] ));
 sg13g2_dfrbp_1 _18356_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net342),
    .D(_00214_),
    .Q_N(_00081_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[13] ));
 sg13g2_dfrbp_1 _18357_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net341),
    .D(_00215_),
    .Q_N(_00079_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[12] ));
 sg13g2_dfrbp_1 _18358_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net340),
    .D(_00216_),
    .Q_N(_00016_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[11] ));
 sg13g2_dfrbp_1 _18359_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net339),
    .D(_00217_),
    .Q_N(_00070_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[10] ));
 sg13g2_dfrbp_1 _18360_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net338),
    .D(_00218_),
    .Q_N(_00068_),
    .Q(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[2] ));
 sg13g2_dfrbp_1 _18361_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net337),
    .D(_00219_),
    .Q_N(_00066_),
    .Q(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[1] ));
 sg13g2_dfrbp_1 _18362_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net336),
    .D(_00220_),
    .Q_N(_00018_),
    .Q(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[0] ));
 sg13g2_dfrbp_1 _18363_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net335),
    .D(_00221_),
    .Q_N(_00022_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[6] ));
 sg13g2_dfrbp_1 _18364_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net334),
    .D(_00222_),
    .Q_N(_00020_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[5] ));
 sg13g2_dfrbp_1 _18365_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net333),
    .D(_00223_),
    .Q_N(_00008_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[4] ));
 sg13g2_dfrbp_1 _18366_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net332),
    .D(_00224_),
    .Q_N(_00012_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[3] ));
 sg13g2_dfrbp_1 _18367_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net331),
    .D(_00225_),
    .Q_N(_00010_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[2] ));
 sg13g2_dfrbp_1 _18368_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net330),
    .D(_00226_),
    .Q_N(_00119_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[1] ));
 sg13g2_dfrbp_1 _18369_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net329),
    .D(net3413),
    .Q_N(_00089_),
    .Q(\m_sys.m_core.m_bru.io_i_s1[0] ));
 sg13g2_dfrbp_1 _18370_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net328),
    .D(_00228_),
    .Q_N(_09082_),
    .Q(\m_sys.m_uart.m_tx.r_cstate[1] ));
 sg13g2_dfrbp_1 _18371_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net326),
    .D(_00229_),
    .Q_N(_00014_),
    .Q(\m_sys.m_uart.m_tx.r_cstate[0] ));
 sg13g2_dfrbp_1 _18372_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net324),
    .D(_00230_),
    .Q_N(_09081_),
    .Q(\m_sys.m_uart.m_rx.r_cstate[1] ));
 sg13g2_dfrbp_1 _18373_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net322),
    .D(_00231_),
    .Q_N(_09080_),
    .Q(\m_sys.m_uart.m_rx.r_cstate[0] ));
 sg13g2_dfrbp_1 _18374_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net320),
    .D(_00232_),
    .Q_N(_09079_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][0] ));
 sg13g2_dfrbp_1 _18375_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net319),
    .D(_00233_),
    .Q_N(_09078_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][1] ));
 sg13g2_dfrbp_1 _18376_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net318),
    .D(_00234_),
    .Q_N(_09077_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][2] ));
 sg13g2_dfrbp_1 _18377_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net317),
    .D(_00235_),
    .Q_N(_09076_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][3] ));
 sg13g2_dfrbp_1 _18378_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net316),
    .D(_00236_),
    .Q_N(_09075_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][4] ));
 sg13g2_dfrbp_1 _18379_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net315),
    .D(_00237_),
    .Q_N(_09074_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][5] ));
 sg13g2_dfrbp_1 _18380_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net314),
    .D(_00238_),
    .Q_N(_09073_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][6] ));
 sg13g2_dfrbp_1 _18381_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net313),
    .D(_00239_),
    .Q_N(_09072_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][7] ));
 sg13g2_dfrbp_1 _18382_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net312),
    .D(_00240_),
    .Q_N(_09071_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][8] ));
 sg13g2_dfrbp_1 _18383_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net311),
    .D(_00241_),
    .Q_N(_09070_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][9] ));
 sg13g2_dfrbp_1 _18384_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net310),
    .D(_00242_),
    .Q_N(_09069_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][10] ));
 sg13g2_dfrbp_1 _18385_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net309),
    .D(_00243_),
    .Q_N(_09068_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][11] ));
 sg13g2_dfrbp_1 _18386_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net308),
    .D(_00244_),
    .Q_N(_09067_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][12] ));
 sg13g2_dfrbp_1 _18387_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net307),
    .D(_00245_),
    .Q_N(_09066_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][13] ));
 sg13g2_dfrbp_1 _18388_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net306),
    .D(_00246_),
    .Q_N(_09065_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][14] ));
 sg13g2_dfrbp_1 _18389_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net305),
    .D(_00247_),
    .Q_N(_09064_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][15] ));
 sg13g2_dfrbp_1 _18390_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net304),
    .D(_00248_),
    .Q_N(_09063_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][16] ));
 sg13g2_dfrbp_1 _18391_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net303),
    .D(_00249_),
    .Q_N(_09062_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][17] ));
 sg13g2_dfrbp_1 _18392_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net302),
    .D(_00250_),
    .Q_N(_09061_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][18] ));
 sg13g2_dfrbp_1 _18393_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net301),
    .D(_00251_),
    .Q_N(_09060_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][19] ));
 sg13g2_dfrbp_1 _18394_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net300),
    .D(_00252_),
    .Q_N(_09059_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][20] ));
 sg13g2_dfrbp_1 _18395_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net299),
    .D(_00253_),
    .Q_N(_09058_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][21] ));
 sg13g2_dfrbp_1 _18396_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net298),
    .D(_00254_),
    .Q_N(_09057_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][22] ));
 sg13g2_dfrbp_1 _18397_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net297),
    .D(_00255_),
    .Q_N(_09056_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][23] ));
 sg13g2_dfrbp_1 _18398_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net296),
    .D(_00256_),
    .Q_N(_09055_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][0] ));
 sg13g2_dfrbp_1 _18399_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net295),
    .D(_00257_),
    .Q_N(_09054_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][1] ));
 sg13g2_dfrbp_1 _18400_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net294),
    .D(_00258_),
    .Q_N(_09053_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][2] ));
 sg13g2_dfrbp_1 _18401_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net293),
    .D(_00259_),
    .Q_N(_09052_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][3] ));
 sg13g2_dfrbp_1 _18402_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net292),
    .D(_00260_),
    .Q_N(_09051_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][4] ));
 sg13g2_dfrbp_1 _18403_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net291),
    .D(_00261_),
    .Q_N(_09050_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][5] ));
 sg13g2_dfrbp_1 _18404_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net290),
    .D(_00262_),
    .Q_N(_09049_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][6] ));
 sg13g2_dfrbp_1 _18405_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net289),
    .D(_00263_),
    .Q_N(_09048_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][7] ));
 sg13g2_dfrbp_1 _18406_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net288),
    .D(_00264_),
    .Q_N(_09047_),
    .Q(\m_sys.m_core.m_fsm.r_cstate[2] ));
 sg13g2_dfrbp_1 _18407_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net287),
    .D(_00265_),
    .Q_N(_00027_),
    .Q(\m_sys._m_core_io_b_mem_wdata[0] ));
 sg13g2_dfrbp_1 _18408_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net286),
    .D(_00266_),
    .Q_N(_09046_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][0] ));
 sg13g2_dfrbp_1 _18409_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net285),
    .D(_00267_),
    .Q_N(_09045_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][1] ));
 sg13g2_dfrbp_1 _18410_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net284),
    .D(_00268_),
    .Q_N(_09044_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][2] ));
 sg13g2_dfrbp_1 _18411_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net283),
    .D(_00269_),
    .Q_N(_09043_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][3] ));
 sg13g2_dfrbp_1 _18412_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net282),
    .D(_00270_),
    .Q_N(_09042_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][4] ));
 sg13g2_dfrbp_1 _18413_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net281),
    .D(_00271_),
    .Q_N(_09041_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][5] ));
 sg13g2_dfrbp_1 _18414_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net280),
    .D(_00272_),
    .Q_N(_09040_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][6] ));
 sg13g2_dfrbp_1 _18415_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net279),
    .D(_00273_),
    .Q_N(_09039_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][7] ));
 sg13g2_dfrbp_1 _18416_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net278),
    .D(_00274_),
    .Q_N(_09038_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][8] ));
 sg13g2_dfrbp_1 _18417_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net277),
    .D(_00275_),
    .Q_N(_09037_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][9] ));
 sg13g2_dfrbp_1 _18418_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net276),
    .D(_00276_),
    .Q_N(_09036_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][10] ));
 sg13g2_dfrbp_1 _18419_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net275),
    .D(_00277_),
    .Q_N(_09035_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][11] ));
 sg13g2_dfrbp_1 _18420_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net274),
    .D(_00278_),
    .Q_N(_09034_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][12] ));
 sg13g2_dfrbp_1 _18421_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net273),
    .D(_00279_),
    .Q_N(_09033_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][13] ));
 sg13g2_dfrbp_1 _18422_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net272),
    .D(_00280_),
    .Q_N(_09032_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][14] ));
 sg13g2_dfrbp_1 _18423_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net271),
    .D(_00281_),
    .Q_N(_09031_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][15] ));
 sg13g2_dfrbp_1 _18424_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net270),
    .D(_00282_),
    .Q_N(_09030_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][24] ));
 sg13g2_dfrbp_1 _18425_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net269),
    .D(_00283_),
    .Q_N(_09029_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][25] ));
 sg13g2_dfrbp_1 _18426_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net268),
    .D(_00284_),
    .Q_N(_09028_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][26] ));
 sg13g2_dfrbp_1 _18427_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net267),
    .D(_00285_),
    .Q_N(_09027_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][27] ));
 sg13g2_dfrbp_1 _18428_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net266),
    .D(_00286_),
    .Q_N(_09026_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][28] ));
 sg13g2_dfrbp_1 _18429_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net265),
    .D(_00287_),
    .Q_N(_09025_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][29] ));
 sg13g2_dfrbp_1 _18430_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net264),
    .D(_00288_),
    .Q_N(_09024_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][30] ));
 sg13g2_dfrbp_1 _18431_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net263),
    .D(_00289_),
    .Q_N(_09023_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][31] ));
 sg13g2_dfrbp_1 _18432_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net262),
    .D(_00290_),
    .Q_N(_09022_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][0] ));
 sg13g2_dfrbp_1 _18433_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net261),
    .D(_00291_),
    .Q_N(_09021_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][1] ));
 sg13g2_dfrbp_1 _18434_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net260),
    .D(_00292_),
    .Q_N(_09020_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][2] ));
 sg13g2_dfrbp_1 _18435_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net259),
    .D(_00293_),
    .Q_N(_09019_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][3] ));
 sg13g2_dfrbp_1 _18436_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net258),
    .D(_00294_),
    .Q_N(_09018_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][4] ));
 sg13g2_dfrbp_1 _18437_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net257),
    .D(_00295_),
    .Q_N(_09017_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][5] ));
 sg13g2_dfrbp_1 _18438_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net256),
    .D(_00296_),
    .Q_N(_09016_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][6] ));
 sg13g2_dfrbp_1 _18439_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net255),
    .D(_00297_),
    .Q_N(_09015_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][7] ));
 sg13g2_dfrbp_1 _18440_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net254),
    .D(_00298_),
    .Q_N(_09014_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][8] ));
 sg13g2_dfrbp_1 _18441_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net253),
    .D(_00299_),
    .Q_N(_09013_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][9] ));
 sg13g2_dfrbp_1 _18442_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net252),
    .D(_00300_),
    .Q_N(_09012_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][10] ));
 sg13g2_dfrbp_1 _18443_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net251),
    .D(_00301_),
    .Q_N(_09011_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][11] ));
 sg13g2_dfrbp_1 _18444_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net250),
    .D(_00302_),
    .Q_N(_09010_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][12] ));
 sg13g2_dfrbp_1 _18445_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net249),
    .D(_00303_),
    .Q_N(_09009_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][13] ));
 sg13g2_dfrbp_1 _18446_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net248),
    .D(_00304_),
    .Q_N(_09008_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][14] ));
 sg13g2_dfrbp_1 _18447_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net247),
    .D(_00305_),
    .Q_N(_09007_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][15] ));
 sg13g2_dfrbp_1 _18448_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net246),
    .D(_00306_),
    .Q_N(_09006_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][16] ));
 sg13g2_dfrbp_1 _18449_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net245),
    .D(_00307_),
    .Q_N(_09005_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][17] ));
 sg13g2_dfrbp_1 _18450_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net244),
    .D(_00308_),
    .Q_N(_09004_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][18] ));
 sg13g2_dfrbp_1 _18451_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net243),
    .D(_00309_),
    .Q_N(_09003_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][19] ));
 sg13g2_dfrbp_1 _18452_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net242),
    .D(_00310_),
    .Q_N(_09002_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][20] ));
 sg13g2_dfrbp_1 _18453_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net241),
    .D(_00311_),
    .Q_N(_09001_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][21] ));
 sg13g2_dfrbp_1 _18454_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net240),
    .D(_00312_),
    .Q_N(_09000_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][22] ));
 sg13g2_dfrbp_1 _18455_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net239),
    .D(_00313_),
    .Q_N(_08999_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][23] ));
 sg13g2_dfrbp_1 _18456_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net238),
    .D(_00314_),
    .Q_N(_08998_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][0] ));
 sg13g2_dfrbp_1 _18457_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net237),
    .D(_00315_),
    .Q_N(_08997_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][1] ));
 sg13g2_dfrbp_1 _18458_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net236),
    .D(_00316_),
    .Q_N(_08996_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][2] ));
 sg13g2_dfrbp_1 _18459_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net235),
    .D(_00317_),
    .Q_N(_08995_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][3] ));
 sg13g2_dfrbp_1 _18460_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net234),
    .D(_00318_),
    .Q_N(_08994_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][4] ));
 sg13g2_dfrbp_1 _18461_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net233),
    .D(_00319_),
    .Q_N(_08993_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][5] ));
 sg13g2_dfrbp_1 _18462_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net232),
    .D(_00320_),
    .Q_N(_08992_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][6] ));
 sg13g2_dfrbp_1 _18463_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net231),
    .D(_00321_),
    .Q_N(_08991_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][7] ));
 sg13g2_dfrbp_1 _18464_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net230),
    .D(_00322_),
    .Q_N(_08990_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][8] ));
 sg13g2_dfrbp_1 _18465_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net229),
    .D(_00323_),
    .Q_N(_08989_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][9] ));
 sg13g2_dfrbp_1 _18466_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net228),
    .D(_00324_),
    .Q_N(_08988_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][10] ));
 sg13g2_dfrbp_1 _18467_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net227),
    .D(_00325_),
    .Q_N(_08987_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][11] ));
 sg13g2_dfrbp_1 _18468_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net226),
    .D(_00326_),
    .Q_N(_08986_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][12] ));
 sg13g2_dfrbp_1 _18469_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net225),
    .D(_00327_),
    .Q_N(_08985_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][13] ));
 sg13g2_dfrbp_1 _18470_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net224),
    .D(_00328_),
    .Q_N(_08984_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][14] ));
 sg13g2_dfrbp_1 _18471_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net223),
    .D(_00329_),
    .Q_N(_08983_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][15] ));
 sg13g2_dfrbp_1 _18472_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net222),
    .D(_00330_),
    .Q_N(_08982_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][16] ));
 sg13g2_dfrbp_1 _18473_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net221),
    .D(_00331_),
    .Q_N(_08981_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][17] ));
 sg13g2_dfrbp_1 _18474_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net220),
    .D(_00332_),
    .Q_N(_08980_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][18] ));
 sg13g2_dfrbp_1 _18475_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net219),
    .D(_00333_),
    .Q_N(_08979_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][19] ));
 sg13g2_dfrbp_1 _18476_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net218),
    .D(_00334_),
    .Q_N(_08978_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][20] ));
 sg13g2_dfrbp_1 _18477_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net217),
    .D(_00335_),
    .Q_N(_08977_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][21] ));
 sg13g2_dfrbp_1 _18478_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net216),
    .D(_00336_),
    .Q_N(_08976_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][22] ));
 sg13g2_dfrbp_1 _18479_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net215),
    .D(_00337_),
    .Q_N(_08975_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][23] ));
 sg13g2_dfrbp_1 _18480_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net214),
    .D(_00338_),
    .Q_N(_08974_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][8] ));
 sg13g2_dfrbp_1 _18481_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net213),
    .D(_00339_),
    .Q_N(_08973_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][9] ));
 sg13g2_dfrbp_1 _18482_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net212),
    .D(_00340_),
    .Q_N(_08972_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][10] ));
 sg13g2_dfrbp_1 _18483_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net211),
    .D(_00341_),
    .Q_N(_08971_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][11] ));
 sg13g2_dfrbp_1 _18484_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net210),
    .D(_00342_),
    .Q_N(_08970_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][12] ));
 sg13g2_dfrbp_1 _18485_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net209),
    .D(_00343_),
    .Q_N(_08969_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][13] ));
 sg13g2_dfrbp_1 _18486_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net208),
    .D(_00344_),
    .Q_N(_08968_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][14] ));
 sg13g2_dfrbp_1 _18487_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net207),
    .D(_00345_),
    .Q_N(_08967_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][15] ));
 sg13g2_dfrbp_1 _18488_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net206),
    .D(_00346_),
    .Q_N(_08966_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][16] ));
 sg13g2_dfrbp_1 _18489_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net205),
    .D(_00347_),
    .Q_N(_08965_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][17] ));
 sg13g2_dfrbp_1 _18490_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net204),
    .D(_00348_),
    .Q_N(_08964_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][18] ));
 sg13g2_dfrbp_1 _18491_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net203),
    .D(_00349_),
    .Q_N(_08963_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][19] ));
 sg13g2_dfrbp_1 _18492_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net202),
    .D(_00350_),
    .Q_N(_08962_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][20] ));
 sg13g2_dfrbp_1 _18493_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net201),
    .D(_00351_),
    .Q_N(_08961_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][21] ));
 sg13g2_dfrbp_1 _18494_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net200),
    .D(_00352_),
    .Q_N(_08960_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][22] ));
 sg13g2_dfrbp_1 _18495_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net199),
    .D(_00353_),
    .Q_N(_08959_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][23] ));
 sg13g2_dfrbp_1 _18496_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net198),
    .D(_00354_),
    .Q_N(_08958_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][0] ));
 sg13g2_dfrbp_1 _18497_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net197),
    .D(_00355_),
    .Q_N(_08957_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][1] ));
 sg13g2_dfrbp_1 _18498_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net196),
    .D(_00356_),
    .Q_N(_08956_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][2] ));
 sg13g2_dfrbp_1 _18499_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net195),
    .D(_00357_),
    .Q_N(_08955_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][3] ));
 sg13g2_dfrbp_1 _18500_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net194),
    .D(_00358_),
    .Q_N(_08954_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][4] ));
 sg13g2_dfrbp_1 _18501_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net193),
    .D(_00359_),
    .Q_N(_08953_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][5] ));
 sg13g2_dfrbp_1 _18502_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net192),
    .D(_00360_),
    .Q_N(_08952_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][6] ));
 sg13g2_dfrbp_1 _18503_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net191),
    .D(_00361_),
    .Q_N(_08951_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][7] ));
 sg13g2_dfrbp_1 _18504_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net190),
    .D(_00362_),
    .Q_N(_08950_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][8] ));
 sg13g2_dfrbp_1 _18505_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net189),
    .D(_00363_),
    .Q_N(_08949_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][9] ));
 sg13g2_dfrbp_1 _18506_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net188),
    .D(_00364_),
    .Q_N(_08948_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][10] ));
 sg13g2_dfrbp_1 _18507_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net187),
    .D(_00365_),
    .Q_N(_08947_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][11] ));
 sg13g2_dfrbp_1 _18508_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net186),
    .D(_00366_),
    .Q_N(_08946_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][12] ));
 sg13g2_dfrbp_1 _18509_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net185),
    .D(_00367_),
    .Q_N(_08945_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][13] ));
 sg13g2_dfrbp_1 _18510_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net184),
    .D(_00368_),
    .Q_N(_08944_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][14] ));
 sg13g2_dfrbp_1 _18511_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net183),
    .D(_00369_),
    .Q_N(_08943_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][15] ));
 sg13g2_dfrbp_1 _18512_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net182),
    .D(_00370_),
    .Q_N(_08942_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][16] ));
 sg13g2_dfrbp_1 _18513_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net181),
    .D(_00371_),
    .Q_N(_08941_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][17] ));
 sg13g2_dfrbp_1 _18514_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net180),
    .D(_00372_),
    .Q_N(_08940_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][18] ));
 sg13g2_dfrbp_1 _18515_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net179),
    .D(_00373_),
    .Q_N(_08939_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][19] ));
 sg13g2_dfrbp_1 _18516_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net178),
    .D(_00374_),
    .Q_N(_08938_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][20] ));
 sg13g2_dfrbp_1 _18517_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net177),
    .D(_00375_),
    .Q_N(_08937_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][21] ));
 sg13g2_dfrbp_1 _18518_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net176),
    .D(_00376_),
    .Q_N(_08936_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][22] ));
 sg13g2_dfrbp_1 _18519_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net175),
    .D(_00377_),
    .Q_N(_08935_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][23] ));
 sg13g2_dfrbp_1 _18520_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net174),
    .D(_00378_),
    .Q_N(_08934_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][0] ));
 sg13g2_dfrbp_1 _18521_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net173),
    .D(_00379_),
    .Q_N(_08933_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][1] ));
 sg13g2_dfrbp_1 _18522_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net172),
    .D(_00380_),
    .Q_N(_08932_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][2] ));
 sg13g2_dfrbp_1 _18523_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net171),
    .D(_00381_),
    .Q_N(_08931_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][3] ));
 sg13g2_dfrbp_1 _18524_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net170),
    .D(_00382_),
    .Q_N(_08930_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][4] ));
 sg13g2_dfrbp_1 _18525_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net169),
    .D(_00383_),
    .Q_N(_08929_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][5] ));
 sg13g2_dfrbp_1 _18526_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net168),
    .D(_00384_),
    .Q_N(_08928_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][6] ));
 sg13g2_dfrbp_1 _18527_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net167),
    .D(_00385_),
    .Q_N(_08927_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][7] ));
 sg13g2_dfrbp_1 _18528_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net166),
    .D(_00386_),
    .Q_N(_08926_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][8] ));
 sg13g2_dfrbp_1 _18529_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net165),
    .D(_00387_),
    .Q_N(_08925_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][9] ));
 sg13g2_dfrbp_1 _18530_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net164),
    .D(_00388_),
    .Q_N(_08924_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][10] ));
 sg13g2_dfrbp_1 _18531_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net163),
    .D(_00389_),
    .Q_N(_08923_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][11] ));
 sg13g2_dfrbp_1 _18532_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net162),
    .D(_00390_),
    .Q_N(_08922_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][12] ));
 sg13g2_dfrbp_1 _18533_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net161),
    .D(_00391_),
    .Q_N(_08921_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][13] ));
 sg13g2_dfrbp_1 _18534_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net160),
    .D(_00392_),
    .Q_N(_08920_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][14] ));
 sg13g2_dfrbp_1 _18535_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net159),
    .D(_00393_),
    .Q_N(_08919_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][15] ));
 sg13g2_dfrbp_1 _18536_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net158),
    .D(_00394_),
    .Q_N(_08918_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][16] ));
 sg13g2_dfrbp_1 _18537_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net157),
    .D(_00395_),
    .Q_N(_08917_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][17] ));
 sg13g2_dfrbp_1 _18538_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net156),
    .D(_00396_),
    .Q_N(_08916_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][18] ));
 sg13g2_dfrbp_1 _18539_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net155),
    .D(_00397_),
    .Q_N(_08915_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][19] ));
 sg13g2_dfrbp_1 _18540_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net154),
    .D(_00398_),
    .Q_N(_08914_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][20] ));
 sg13g2_dfrbp_1 _18541_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net153),
    .D(_00399_),
    .Q_N(_08913_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][21] ));
 sg13g2_dfrbp_1 _18542_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net152),
    .D(_00400_),
    .Q_N(_08912_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][22] ));
 sg13g2_dfrbp_1 _18543_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net151),
    .D(_00401_),
    .Q_N(_08911_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][23] ));
 sg13g2_dfrbp_1 _18544_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net150),
    .D(_00402_),
    .Q_N(_08910_),
    .Q(\m_sys.m_core.m_fsm.r_cstate[1] ));
 sg13g2_dfrbp_1 _18545_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net149),
    .D(_00403_),
    .Q_N(_00087_),
    .Q(\m_sys.m_core.m_bru.io_i_uop[0] ));
 sg13g2_dfrbp_1 _18546_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net147),
    .D(net3180),
    .Q_N(_08909_),
    .Q(\m_sys.m_core.m_bru.io_i_uop[1] ));
 sg13g2_dfrbp_1 _18547_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net145),
    .D(_00405_),
    .Q_N(_08908_),
    .Q(\m_sys.m_core.m_alu.io_i_uop[0] ));
 sg13g2_dfrbp_1 _18548_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net143),
    .D(_00406_),
    .Q_N(_00088_),
    .Q(\m_sys.m_core.m_alu.io_i_uop[1] ));
 sg13g2_dfrbp_1 _18549_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net141),
    .D(_00407_),
    .Q_N(_08907_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][24] ));
 sg13g2_dfrbp_1 _18550_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net140),
    .D(_00408_),
    .Q_N(_08906_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][25] ));
 sg13g2_dfrbp_1 _18551_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net139),
    .D(_00409_),
    .Q_N(_08905_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][26] ));
 sg13g2_dfrbp_1 _18552_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net138),
    .D(_00410_),
    .Q_N(_08904_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][27] ));
 sg13g2_dfrbp_1 _18553_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net137),
    .D(_00411_),
    .Q_N(_08903_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][28] ));
 sg13g2_dfrbp_1 _18554_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net136),
    .D(_00412_),
    .Q_N(_08902_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][29] ));
 sg13g2_dfrbp_1 _18555_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net135),
    .D(_00413_),
    .Q_N(_08901_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][30] ));
 sg13g2_dfrbp_1 _18556_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net134),
    .D(_00414_),
    .Q_N(_08900_),
    .Q(\m_sys.m_ram.m_ram.r_mem[13][31] ));
 sg13g2_dfrbp_1 _18557_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net133),
    .D(_00415_),
    .Q_N(_08899_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][0] ));
 sg13g2_dfrbp_1 _18558_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net132),
    .D(_00416_),
    .Q_N(_08898_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][1] ));
 sg13g2_dfrbp_1 _18559_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net131),
    .D(_00417_),
    .Q_N(_08897_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][2] ));
 sg13g2_dfrbp_1 _18560_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net130),
    .D(_00418_),
    .Q_N(_08896_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][3] ));
 sg13g2_dfrbp_1 _18561_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net129),
    .D(_00419_),
    .Q_N(_08895_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][4] ));
 sg13g2_dfrbp_1 _18562_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net128),
    .D(_00420_),
    .Q_N(_08894_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][5] ));
 sg13g2_dfrbp_1 _18563_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net127),
    .D(_00421_),
    .Q_N(_08893_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][6] ));
 sg13g2_dfrbp_1 _18564_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net126),
    .D(_00422_),
    .Q_N(_08892_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][7] ));
 sg13g2_dfrbp_1 _18565_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net125),
    .D(_00423_),
    .Q_N(_08891_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][24] ));
 sg13g2_dfrbp_1 _18566_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net124),
    .D(_00424_),
    .Q_N(_08890_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][25] ));
 sg13g2_dfrbp_1 _18567_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net123),
    .D(_00425_),
    .Q_N(_08889_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][26] ));
 sg13g2_dfrbp_1 _18568_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net122),
    .D(_00426_),
    .Q_N(_08888_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][27] ));
 sg13g2_dfrbp_1 _18569_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net121),
    .D(_00427_),
    .Q_N(_08887_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][28] ));
 sg13g2_dfrbp_1 _18570_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net120),
    .D(_00428_),
    .Q_N(_08886_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][29] ));
 sg13g2_dfrbp_1 _18571_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net119),
    .D(_00429_),
    .Q_N(_08885_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][30] ));
 sg13g2_dfrbp_1 _18572_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net118),
    .D(_00430_),
    .Q_N(_08884_),
    .Q(\m_sys.m_ram.m_ram.r_mem[14][31] ));
 sg13g2_dfrbp_1 _18573_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net117),
    .D(_00431_),
    .Q_N(_08883_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][8] ));
 sg13g2_dfrbp_1 _18574_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net116),
    .D(_00432_),
    .Q_N(_08882_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][9] ));
 sg13g2_dfrbp_1 _18575_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net115),
    .D(_00433_),
    .Q_N(_08881_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][10] ));
 sg13g2_dfrbp_1 _18576_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net114),
    .D(_00434_),
    .Q_N(_08880_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][11] ));
 sg13g2_dfrbp_1 _18577_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net113),
    .D(_00435_),
    .Q_N(_08879_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][12] ));
 sg13g2_dfrbp_1 _18578_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net112),
    .D(_00436_),
    .Q_N(_08878_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][13] ));
 sg13g2_dfrbp_1 _18579_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net111),
    .D(_00437_),
    .Q_N(_08877_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][14] ));
 sg13g2_dfrbp_1 _18580_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net110),
    .D(_00438_),
    .Q_N(_08876_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][15] ));
 sg13g2_dfrbp_1 _18581_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net109),
    .D(_00439_),
    .Q_N(_08875_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][24] ));
 sg13g2_dfrbp_1 _18582_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net108),
    .D(_00440_),
    .Q_N(_08874_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][25] ));
 sg13g2_dfrbp_1 _18583_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net107),
    .D(_00441_),
    .Q_N(_08873_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][26] ));
 sg13g2_dfrbp_1 _18584_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net106),
    .D(_00442_),
    .Q_N(_08872_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][27] ));
 sg13g2_dfrbp_1 _18585_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net105),
    .D(_00443_),
    .Q_N(_08871_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][28] ));
 sg13g2_dfrbp_1 _18586_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net104),
    .D(_00444_),
    .Q_N(_08870_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][29] ));
 sg13g2_dfrbp_1 _18587_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net103),
    .D(_00445_),
    .Q_N(_08869_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][30] ));
 sg13g2_dfrbp_1 _18588_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net102),
    .D(_00446_),
    .Q_N(_08868_),
    .Q(\m_sys.m_ram.m_ram.r_mem[15][31] ));
 sg13g2_dfrbp_1 _18589_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net101),
    .D(_00447_),
    .Q_N(_08867_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][16] ));
 sg13g2_dfrbp_1 _18590_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net100),
    .D(_00448_),
    .Q_N(_08866_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][17] ));
 sg13g2_dfrbp_1 _18591_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net99),
    .D(_00449_),
    .Q_N(_08865_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][18] ));
 sg13g2_dfrbp_1 _18592_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net98),
    .D(_00450_),
    .Q_N(_08864_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][19] ));
 sg13g2_dfrbp_1 _18593_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net97),
    .D(_00451_),
    .Q_N(_08863_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][20] ));
 sg13g2_dfrbp_1 _18594_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net96),
    .D(_00452_),
    .Q_N(_08862_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][21] ));
 sg13g2_dfrbp_1 _18595_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net95),
    .D(_00453_),
    .Q_N(_08861_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][22] ));
 sg13g2_dfrbp_1 _18596_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net94),
    .D(_00454_),
    .Q_N(_08860_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][23] ));
 sg13g2_dfrbp_1 _18597_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net93),
    .D(_00455_),
    .Q_N(_08859_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][24] ));
 sg13g2_dfrbp_1 _18598_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net92),
    .D(_00456_),
    .Q_N(_08858_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][25] ));
 sg13g2_dfrbp_1 _18599_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net91),
    .D(_00457_),
    .Q_N(_08857_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][26] ));
 sg13g2_dfrbp_1 _18600_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net90),
    .D(_00458_),
    .Q_N(_08856_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][27] ));
 sg13g2_dfrbp_1 _18601_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net89),
    .D(_00459_),
    .Q_N(_08855_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][28] ));
 sg13g2_dfrbp_1 _18602_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net88),
    .D(_00460_),
    .Q_N(_08854_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][29] ));
 sg13g2_dfrbp_1 _18603_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net87),
    .D(_00461_),
    .Q_N(_08853_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][30] ));
 sg13g2_dfrbp_1 _18604_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net86),
    .D(_00462_),
    .Q_N(_08852_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][31] ));
 sg13g2_dfrbp_1 _18605_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net85),
    .D(_00463_),
    .Q_N(_08851_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][0] ));
 sg13g2_dfrbp_1 _18606_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net84),
    .D(_00464_),
    .Q_N(_08850_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][1] ));
 sg13g2_dfrbp_1 _18607_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net83),
    .D(_00465_),
    .Q_N(_08849_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][2] ));
 sg13g2_dfrbp_1 _18608_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net82),
    .D(_00466_),
    .Q_N(_08848_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][3] ));
 sg13g2_dfrbp_1 _18609_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net81),
    .D(_00467_),
    .Q_N(_08847_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][4] ));
 sg13g2_dfrbp_1 _18610_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net80),
    .D(_00468_),
    .Q_N(_08846_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][5] ));
 sg13g2_dfrbp_1 _18611_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net79),
    .D(_00469_),
    .Q_N(_08845_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][6] ));
 sg13g2_dfrbp_1 _18612_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net78),
    .D(_00470_),
    .Q_N(_08844_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][7] ));
 sg13g2_dfrbp_1 _18613_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net77),
    .D(_00471_),
    .Q_N(_08843_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][24] ));
 sg13g2_dfrbp_1 _18614_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net76),
    .D(_00472_),
    .Q_N(_08842_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][25] ));
 sg13g2_dfrbp_1 _18615_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net75),
    .D(_00473_),
    .Q_N(_08841_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][26] ));
 sg13g2_dfrbp_1 _18616_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net74),
    .D(_00474_),
    .Q_N(_08840_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][27] ));
 sg13g2_dfrbp_1 _18617_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net73),
    .D(_00475_),
    .Q_N(_08839_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][28] ));
 sg13g2_dfrbp_1 _18618_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net72),
    .D(_00476_),
    .Q_N(_08838_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][29] ));
 sg13g2_dfrbp_1 _18619_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net71),
    .D(_00477_),
    .Q_N(_08837_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][30] ));
 sg13g2_dfrbp_1 _18620_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net70),
    .D(_00478_),
    .Q_N(_08836_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][31] ));
 sg13g2_dfrbp_1 _18621_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net69),
    .D(_00479_),
    .Q_N(_08835_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][8] ));
 sg13g2_dfrbp_1 _18622_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net68),
    .D(_00480_),
    .Q_N(_08834_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][9] ));
 sg13g2_dfrbp_1 _18623_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net67),
    .D(_00481_),
    .Q_N(_08833_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][10] ));
 sg13g2_dfrbp_1 _18624_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net66),
    .D(_00482_),
    .Q_N(_08832_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][11] ));
 sg13g2_dfrbp_1 _18625_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net65),
    .D(_00483_),
    .Q_N(_08831_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][12] ));
 sg13g2_dfrbp_1 _18626_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net64),
    .D(_00484_),
    .Q_N(_08830_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][13] ));
 sg13g2_dfrbp_1 _18627_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net63),
    .D(_00485_),
    .Q_N(_08829_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][14] ));
 sg13g2_dfrbp_1 _18628_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net62),
    .D(_00486_),
    .Q_N(_08828_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][15] ));
 sg13g2_dfrbp_1 _18629_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net61),
    .D(_00487_),
    .Q_N(_08827_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][16] ));
 sg13g2_dfrbp_1 _18630_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net60),
    .D(_00488_),
    .Q_N(_08826_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][17] ));
 sg13g2_dfrbp_1 _18631_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net59),
    .D(_00489_),
    .Q_N(_08825_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][18] ));
 sg13g2_dfrbp_1 _18632_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net58),
    .D(_00490_),
    .Q_N(_08824_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][19] ));
 sg13g2_dfrbp_1 _18633_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net57),
    .D(_00491_),
    .Q_N(_08823_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][20] ));
 sg13g2_dfrbp_1 _18634_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net56),
    .D(_00492_),
    .Q_N(_08822_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][21] ));
 sg13g2_dfrbp_1 _18635_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net55),
    .D(_00493_),
    .Q_N(_08821_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][22] ));
 sg13g2_dfrbp_1 _18636_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net54),
    .D(_00494_),
    .Q_N(_08820_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][23] ));
 sg13g2_dfrbp_1 _18637_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net53),
    .D(_00495_),
    .Q_N(_08819_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][24] ));
 sg13g2_dfrbp_1 _18638_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net52),
    .D(_00496_),
    .Q_N(_08818_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][25] ));
 sg13g2_dfrbp_1 _18639_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net51),
    .D(_00497_),
    .Q_N(_08817_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][26] ));
 sg13g2_dfrbp_1 _18640_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net50),
    .D(_00498_),
    .Q_N(_08816_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][27] ));
 sg13g2_dfrbp_1 _18641_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net49),
    .D(_00499_),
    .Q_N(_08815_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][28] ));
 sg13g2_dfrbp_1 _18642_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net48),
    .D(_00500_),
    .Q_N(_08814_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][29] ));
 sg13g2_dfrbp_1 _18643_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net47),
    .D(_00501_),
    .Q_N(_08813_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][30] ));
 sg13g2_dfrbp_1 _18644_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net46),
    .D(_00502_),
    .Q_N(_08812_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][31] ));
 sg13g2_dfrbp_1 _18645_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net45),
    .D(_00503_),
    .Q_N(_08811_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][16] ));
 sg13g2_dfrbp_1 _18646_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net44),
    .D(_00504_),
    .Q_N(_08810_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][17] ));
 sg13g2_dfrbp_1 _18647_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net43),
    .D(_00505_),
    .Q_N(_08809_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][18] ));
 sg13g2_dfrbp_1 _18648_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net42),
    .D(_00506_),
    .Q_N(_08808_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][19] ));
 sg13g2_dfrbp_1 _18649_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net41),
    .D(_00507_),
    .Q_N(_08807_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][20] ));
 sg13g2_dfrbp_1 _18650_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net40),
    .D(_00508_),
    .Q_N(_08806_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][21] ));
 sg13g2_dfrbp_1 _18651_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net39),
    .D(_00509_),
    .Q_N(_08805_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][22] ));
 sg13g2_dfrbp_1 _18652_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net38),
    .D(_00510_),
    .Q_N(_08804_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][23] ));
 sg13g2_dfrbp_1 _18653_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net37),
    .D(_00511_),
    .Q_N(_08803_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][24] ));
 sg13g2_dfrbp_1 _18654_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net36),
    .D(_00512_),
    .Q_N(_08802_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][25] ));
 sg13g2_dfrbp_1 _18655_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net35),
    .D(_00513_),
    .Q_N(_08801_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][26] ));
 sg13g2_dfrbp_1 _18656_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net34),
    .D(_00514_),
    .Q_N(_08800_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][27] ));
 sg13g2_dfrbp_1 _18657_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net33),
    .D(_00515_),
    .Q_N(_08799_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][28] ));
 sg13g2_dfrbp_1 _18658_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net32),
    .D(_00516_),
    .Q_N(_08798_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][29] ));
 sg13g2_dfrbp_1 _18659_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net31),
    .D(_00517_),
    .Q_N(_08797_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][30] ));
 sg13g2_dfrbp_1 _18660_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net30),
    .D(_00518_),
    .Q_N(_08796_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][31] ));
 sg13g2_dfrbp_1 _18661_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net29),
    .D(_00519_),
    .Q_N(_08795_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][0] ));
 sg13g2_dfrbp_1 _18662_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net28),
    .D(_00520_),
    .Q_N(_08794_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][1] ));
 sg13g2_dfrbp_1 _18663_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net27),
    .D(_00521_),
    .Q_N(_08793_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][2] ));
 sg13g2_dfrbp_1 _18664_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net26),
    .D(_00522_),
    .Q_N(_08792_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][3] ));
 sg13g2_dfrbp_1 _18665_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net25),
    .D(_00523_),
    .Q_N(_08791_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][4] ));
 sg13g2_dfrbp_1 _18666_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net24),
    .D(_00524_),
    .Q_N(_08790_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][5] ));
 sg13g2_dfrbp_1 _18667_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net23),
    .D(_00525_),
    .Q_N(_08789_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][6] ));
 sg13g2_dfrbp_1 _18668_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net22),
    .D(_00526_),
    .Q_N(_08788_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][7] ));
 sg13g2_dfrbp_1 _18669_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net21),
    .D(_00527_),
    .Q_N(_08787_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][24] ));
 sg13g2_dfrbp_1 _18670_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net20),
    .D(_00528_),
    .Q_N(_08786_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][25] ));
 sg13g2_dfrbp_1 _18671_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net19),
    .D(_00529_),
    .Q_N(_08785_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][26] ));
 sg13g2_dfrbp_1 _18672_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net18),
    .D(_00530_),
    .Q_N(_08784_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][27] ));
 sg13g2_dfrbp_1 _18673_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net17),
    .D(_00531_),
    .Q_N(_08783_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][28] ));
 sg13g2_dfrbp_1 _18674_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1653),
    .D(_00532_),
    .Q_N(_08782_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][29] ));
 sg13g2_dfrbp_1 _18675_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1652),
    .D(_00533_),
    .Q_N(_08781_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][30] ));
 sg13g2_dfrbp_1 _18676_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1651),
    .D(_00534_),
    .Q_N(_08780_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][31] ));
 sg13g2_dfrbp_1 _18677_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1650),
    .D(_00535_),
    .Q_N(_08779_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][8] ));
 sg13g2_dfrbp_1 _18678_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1649),
    .D(_00536_),
    .Q_N(_08778_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][9] ));
 sg13g2_dfrbp_1 _18679_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1648),
    .D(_00537_),
    .Q_N(_08777_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][10] ));
 sg13g2_dfrbp_1 _18680_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1647),
    .D(_00538_),
    .Q_N(_08776_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][11] ));
 sg13g2_dfrbp_1 _18681_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1646),
    .D(_00539_),
    .Q_N(_08775_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][12] ));
 sg13g2_dfrbp_1 _18682_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1645),
    .D(_00540_),
    .Q_N(_08774_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][13] ));
 sg13g2_dfrbp_1 _18683_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1644),
    .D(_00541_),
    .Q_N(_08773_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][14] ));
 sg13g2_dfrbp_1 _18684_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1643),
    .D(_00542_),
    .Q_N(_08772_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][15] ));
 sg13g2_dfrbp_1 _18685_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1642),
    .D(_00543_),
    .Q_N(_08771_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][24] ));
 sg13g2_dfrbp_1 _18686_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1641),
    .D(_00544_),
    .Q_N(_08770_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][25] ));
 sg13g2_dfrbp_1 _18687_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1640),
    .D(_00545_),
    .Q_N(_08769_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][26] ));
 sg13g2_dfrbp_1 _18688_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1639),
    .D(_00546_),
    .Q_N(_08768_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][27] ));
 sg13g2_dfrbp_1 _18689_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1638),
    .D(_00547_),
    .Q_N(_08767_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][28] ));
 sg13g2_dfrbp_1 _18690_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1637),
    .D(_00548_),
    .Q_N(_08766_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][29] ));
 sg13g2_dfrbp_1 _18691_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1636),
    .D(_00549_),
    .Q_N(_08765_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][30] ));
 sg13g2_dfrbp_1 _18692_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1635),
    .D(_00550_),
    .Q_N(_08764_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][31] ));
 sg13g2_dfrbp_1 _18693_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1634),
    .D(_00551_),
    .Q_N(_08763_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][16] ));
 sg13g2_dfrbp_1 _18694_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1633),
    .D(_00552_),
    .Q_N(_08762_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][17] ));
 sg13g2_dfrbp_1 _18695_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1632),
    .D(_00553_),
    .Q_N(_08761_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][18] ));
 sg13g2_dfrbp_1 _18696_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1631),
    .D(_00554_),
    .Q_N(_08760_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][19] ));
 sg13g2_dfrbp_1 _18697_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1630),
    .D(_00555_),
    .Q_N(_08759_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][20] ));
 sg13g2_dfrbp_1 _18698_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1629),
    .D(_00556_),
    .Q_N(_08758_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][21] ));
 sg13g2_dfrbp_1 _18699_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1628),
    .D(_00557_),
    .Q_N(_08757_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][22] ));
 sg13g2_dfrbp_1 _18700_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1627),
    .D(_00558_),
    .Q_N(_08756_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][23] ));
 sg13g2_dfrbp_1 _18701_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1626),
    .D(_00559_),
    .Q_N(_08755_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][24] ));
 sg13g2_dfrbp_1 _18702_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1625),
    .D(_00560_),
    .Q_N(_08754_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][25] ));
 sg13g2_dfrbp_1 _18703_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1624),
    .D(_00561_),
    .Q_N(_08753_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][26] ));
 sg13g2_dfrbp_1 _18704_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1623),
    .D(_00562_),
    .Q_N(_08752_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][27] ));
 sg13g2_dfrbp_1 _18705_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1622),
    .D(_00563_),
    .Q_N(_08751_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][28] ));
 sg13g2_dfrbp_1 _18706_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1621),
    .D(_00564_),
    .Q_N(_08750_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][29] ));
 sg13g2_dfrbp_1 _18707_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1620),
    .D(_00565_),
    .Q_N(_08749_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][30] ));
 sg13g2_dfrbp_1 _18708_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1619),
    .D(_00566_),
    .Q_N(_08748_),
    .Q(\m_sys.m_ram.m_ram.r_mem[22][31] ));
 sg13g2_dfrbp_1 _18709_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1618),
    .D(_00567_),
    .Q_N(_08747_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][0] ));
 sg13g2_dfrbp_1 _18710_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1617),
    .D(_00568_),
    .Q_N(_08746_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][1] ));
 sg13g2_dfrbp_1 _18711_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1616),
    .D(_00569_),
    .Q_N(_08745_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][2] ));
 sg13g2_dfrbp_1 _18712_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1615),
    .D(_00570_),
    .Q_N(_08744_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][3] ));
 sg13g2_dfrbp_1 _18713_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1614),
    .D(_00571_),
    .Q_N(_08743_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][4] ));
 sg13g2_dfrbp_1 _18714_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1613),
    .D(_00572_),
    .Q_N(_08742_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][5] ));
 sg13g2_dfrbp_1 _18715_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1612),
    .D(_00573_),
    .Q_N(_08741_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][6] ));
 sg13g2_dfrbp_1 _18716_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1611),
    .D(_00574_),
    .Q_N(_08740_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][7] ));
 sg13g2_dfrbp_1 _18717_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1610),
    .D(_00575_),
    .Q_N(_08739_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][24] ));
 sg13g2_dfrbp_1 _18718_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1609),
    .D(_00576_),
    .Q_N(_08738_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][25] ));
 sg13g2_dfrbp_1 _18719_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1608),
    .D(_00577_),
    .Q_N(_08737_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][26] ));
 sg13g2_dfrbp_1 _18720_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1607),
    .D(_00578_),
    .Q_N(_08736_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][27] ));
 sg13g2_dfrbp_1 _18721_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1606),
    .D(_00579_),
    .Q_N(_08735_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][28] ));
 sg13g2_dfrbp_1 _18722_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1605),
    .D(_00580_),
    .Q_N(_08734_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][29] ));
 sg13g2_dfrbp_1 _18723_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1604),
    .D(_00581_),
    .Q_N(_08733_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][30] ));
 sg13g2_dfrbp_1 _18724_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1603),
    .D(_00582_),
    .Q_N(_08732_),
    .Q(\m_sys.m_ram.m_ram.r_mem[23][31] ));
 sg13g2_dfrbp_1 _18725_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1602),
    .D(_00583_),
    .Q_N(_08731_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][8] ));
 sg13g2_dfrbp_1 _18726_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1601),
    .D(_00584_),
    .Q_N(_08730_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][9] ));
 sg13g2_dfrbp_1 _18727_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1600),
    .D(_00585_),
    .Q_N(_08729_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][10] ));
 sg13g2_dfrbp_1 _18728_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1599),
    .D(_00586_),
    .Q_N(_08728_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][11] ));
 sg13g2_dfrbp_1 _18729_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1598),
    .D(_00587_),
    .Q_N(_08727_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][12] ));
 sg13g2_dfrbp_1 _18730_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1597),
    .D(_00588_),
    .Q_N(_08726_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][13] ));
 sg13g2_dfrbp_1 _18731_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1596),
    .D(_00589_),
    .Q_N(_08725_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][14] ));
 sg13g2_dfrbp_1 _18732_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1595),
    .D(_00590_),
    .Q_N(_08724_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][15] ));
 sg13g2_dfrbp_1 _18733_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1594),
    .D(_00591_),
    .Q_N(_08723_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][24] ));
 sg13g2_dfrbp_1 _18734_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1593),
    .D(_00592_),
    .Q_N(_08722_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][25] ));
 sg13g2_dfrbp_1 _18735_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1592),
    .D(_00593_),
    .Q_N(_08721_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][26] ));
 sg13g2_dfrbp_1 _18736_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1591),
    .D(_00594_),
    .Q_N(_08720_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][27] ));
 sg13g2_dfrbp_1 _18737_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1590),
    .D(_00595_),
    .Q_N(_08719_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][28] ));
 sg13g2_dfrbp_1 _18738_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1589),
    .D(_00596_),
    .Q_N(_08718_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][29] ));
 sg13g2_dfrbp_1 _18739_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1588),
    .D(_00597_),
    .Q_N(_08717_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][30] ));
 sg13g2_dfrbp_1 _18740_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1587),
    .D(_00598_),
    .Q_N(_08716_),
    .Q(\m_sys.m_ram.m_ram.r_mem[24][31] ));
 sg13g2_dfrbp_1 _18741_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1586),
    .D(_00599_),
    .Q_N(_08715_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][16] ));
 sg13g2_dfrbp_1 _18742_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1585),
    .D(_00600_),
    .Q_N(_08714_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][17] ));
 sg13g2_dfrbp_1 _18743_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1584),
    .D(_00601_),
    .Q_N(_08713_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][18] ));
 sg13g2_dfrbp_1 _18744_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1583),
    .D(_00602_),
    .Q_N(_08712_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][19] ));
 sg13g2_dfrbp_1 _18745_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1582),
    .D(_00603_),
    .Q_N(_08711_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][20] ));
 sg13g2_dfrbp_1 _18746_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1581),
    .D(_00604_),
    .Q_N(_08710_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][21] ));
 sg13g2_dfrbp_1 _18747_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1580),
    .D(_00605_),
    .Q_N(_08709_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][22] ));
 sg13g2_dfrbp_1 _18748_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1579),
    .D(_00606_),
    .Q_N(_08708_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][23] ));
 sg13g2_dfrbp_1 _18749_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1578),
    .D(_00607_),
    .Q_N(_08707_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][16] ));
 sg13g2_dfrbp_1 _18750_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1577),
    .D(_00608_),
    .Q_N(_08706_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][17] ));
 sg13g2_dfrbp_1 _18751_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1576),
    .D(_00609_),
    .Q_N(_08705_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][18] ));
 sg13g2_dfrbp_1 _18752_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1575),
    .D(_00610_),
    .Q_N(_08704_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][19] ));
 sg13g2_dfrbp_1 _18753_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1574),
    .D(_00611_),
    .Q_N(_08703_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][20] ));
 sg13g2_dfrbp_1 _18754_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1573),
    .D(_00612_),
    .Q_N(_08702_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][21] ));
 sg13g2_dfrbp_1 _18755_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1572),
    .D(_00613_),
    .Q_N(_08701_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][22] ));
 sg13g2_dfrbp_1 _18756_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1571),
    .D(_00614_),
    .Q_N(_08700_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][23] ));
 sg13g2_dfrbp_1 _18757_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1570),
    .D(_00615_),
    .Q_N(_08699_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][24] ));
 sg13g2_dfrbp_1 _18758_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1569),
    .D(_00616_),
    .Q_N(_08698_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][25] ));
 sg13g2_dfrbp_1 _18759_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1568),
    .D(_00617_),
    .Q_N(_08697_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][26] ));
 sg13g2_dfrbp_1 _18760_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1567),
    .D(_00618_),
    .Q_N(_08696_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][27] ));
 sg13g2_dfrbp_1 _18761_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1566),
    .D(_00619_),
    .Q_N(_08695_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][28] ));
 sg13g2_dfrbp_1 _18762_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1565),
    .D(_00620_),
    .Q_N(_08694_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][29] ));
 sg13g2_dfrbp_1 _18763_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1564),
    .D(_00621_),
    .Q_N(_08693_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][30] ));
 sg13g2_dfrbp_1 _18764_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1563),
    .D(_00622_),
    .Q_N(_08692_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][31] ));
 sg13g2_dfrbp_1 _18765_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1562),
    .D(_00623_),
    .Q_N(_08691_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][24] ));
 sg13g2_dfrbp_1 _18766_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1561),
    .D(_00624_),
    .Q_N(_08690_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][25] ));
 sg13g2_dfrbp_1 _18767_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1560),
    .D(_00625_),
    .Q_N(_08689_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][26] ));
 sg13g2_dfrbp_1 _18768_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1559),
    .D(_00626_),
    .Q_N(_08688_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][27] ));
 sg13g2_dfrbp_1 _18769_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1558),
    .D(_00627_),
    .Q_N(_08687_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][28] ));
 sg13g2_dfrbp_1 _18770_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1557),
    .D(_00628_),
    .Q_N(_08686_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][29] ));
 sg13g2_dfrbp_1 _18771_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1556),
    .D(_00629_),
    .Q_N(_08685_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][30] ));
 sg13g2_dfrbp_1 _18772_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1555),
    .D(_00630_),
    .Q_N(_08684_),
    .Q(\m_sys.m_ram.m_ram.r_mem[12][31] ));
 sg13g2_dfrbp_1 _18773_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1554),
    .D(_00631_),
    .Q_N(_08683_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][24] ));
 sg13g2_dfrbp_1 _18774_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1553),
    .D(_00632_),
    .Q_N(_08682_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][25] ));
 sg13g2_dfrbp_1 _18775_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1552),
    .D(_00633_),
    .Q_N(_08681_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][26] ));
 sg13g2_dfrbp_1 _18776_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1551),
    .D(_00634_),
    .Q_N(_08680_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][27] ));
 sg13g2_dfrbp_1 _18777_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1550),
    .D(_00635_),
    .Q_N(_08679_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][28] ));
 sg13g2_dfrbp_1 _18778_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1549),
    .D(_00636_),
    .Q_N(_08678_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][29] ));
 sg13g2_dfrbp_1 _18779_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1548),
    .D(_00637_),
    .Q_N(_08677_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][30] ));
 sg13g2_dfrbp_1 _18780_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1547),
    .D(_00638_),
    .Q_N(_08676_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][31] ));
 sg13g2_dfrbp_1 _18781_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1546),
    .D(_00639_),
    .Q_N(_08675_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][0] ));
 sg13g2_dfrbp_1 _18782_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1545),
    .D(_00640_),
    .Q_N(_08674_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][1] ));
 sg13g2_dfrbp_1 _18783_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1544),
    .D(_00641_),
    .Q_N(_08673_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][2] ));
 sg13g2_dfrbp_1 _18784_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1543),
    .D(_00642_),
    .Q_N(_08672_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][3] ));
 sg13g2_dfrbp_1 _18785_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1542),
    .D(_00643_),
    .Q_N(_08671_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][4] ));
 sg13g2_dfrbp_1 _18786_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1541),
    .D(_00644_),
    .Q_N(_08670_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][5] ));
 sg13g2_dfrbp_1 _18787_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1540),
    .D(_00645_),
    .Q_N(_08669_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][6] ));
 sg13g2_dfrbp_1 _18788_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1539),
    .D(_00646_),
    .Q_N(_08668_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][7] ));
 sg13g2_dfrbp_1 _18789_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1538),
    .D(_00647_),
    .Q_N(_08667_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][0] ));
 sg13g2_dfrbp_1 _18790_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1537),
    .D(_00648_),
    .Q_N(_08666_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][1] ));
 sg13g2_dfrbp_1 _18791_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1536),
    .D(_00649_),
    .Q_N(_08665_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][2] ));
 sg13g2_dfrbp_1 _18792_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1535),
    .D(_00650_),
    .Q_N(_08664_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][3] ));
 sg13g2_dfrbp_1 _18793_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1534),
    .D(_00651_),
    .Q_N(_08663_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][4] ));
 sg13g2_dfrbp_1 _18794_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1533),
    .D(_00652_),
    .Q_N(_08662_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][5] ));
 sg13g2_dfrbp_1 _18795_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1532),
    .D(_00653_),
    .Q_N(_08661_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][6] ));
 sg13g2_dfrbp_1 _18796_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1531),
    .D(_00654_),
    .Q_N(_08660_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][7] ));
 sg13g2_dfrbp_1 _18797_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1530),
    .D(net3367),
    .Q_N(_00011_),
    .Q(\m_sys.m_core.m_bru.io_i_pc[2] ));
 sg13g2_dfrbp_1 _18798_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1528),
    .D(_00656_),
    .Q_N(_00013_),
    .Q(\m_sys.m_core.m_bru.io_i_pc[3] ));
 sg13g2_dfrbp_1 _18799_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1526),
    .D(_00657_),
    .Q_N(_00009_),
    .Q(\m_sys.m_core.m_bru.io_i_pc[4] ));
 sg13g2_dfrbp_1 _18800_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1524),
    .D(net3252),
    .Q_N(_00021_),
    .Q(\m_sys.m_core.m_bru.io_i_pc[5] ));
 sg13g2_dfrbp_1 _18801_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1522),
    .D(_00659_),
    .Q_N(_00023_),
    .Q(\m_sys.m_core.m_bru.io_i_pc[6] ));
 sg13g2_dfrbp_1 _18802_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1520),
    .D(_00660_),
    .Q_N(_00019_),
    .Q(\m_sys.m_core.m_bru.io_i_pc[7] ));
 sg13g2_dfrbp_1 _18803_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1518),
    .D(net3297),
    .Q_N(_00109_),
    .Q(\m_sys.m_core.m_bru.io_i_pc[8] ));
 sg13g2_dfrbp_1 _18804_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1516),
    .D(net3338),
    .Q_N(_00106_),
    .Q(\m_sys.m_core.m_bru.io_i_pc[9] ));
 sg13g2_dfrbp_1 _18805_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1514),
    .D(_00663_),
    .Q_N(_00103_),
    .Q(\m_sys.m_core.m_bru.io_i_pc[10] ));
 sg13g2_dfrbp_1 _18806_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1512),
    .D(_00664_),
    .Q_N(_00017_),
    .Q(\m_sys.m_core.m_bru.io_i_pc[11] ));
 sg13g2_dfrbp_1 _18807_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1510),
    .D(_00665_),
    .Q_N(_08659_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][16] ));
 sg13g2_dfrbp_1 _18808_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1509),
    .D(_00666_),
    .Q_N(_08658_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][17] ));
 sg13g2_dfrbp_1 _18809_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1508),
    .D(_00667_),
    .Q_N(_08657_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][18] ));
 sg13g2_dfrbp_1 _18810_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1507),
    .D(_00668_),
    .Q_N(_08656_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][19] ));
 sg13g2_dfrbp_1 _18811_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1506),
    .D(_00669_),
    .Q_N(_08655_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][20] ));
 sg13g2_dfrbp_1 _18812_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1505),
    .D(_00670_),
    .Q_N(_08654_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][21] ));
 sg13g2_dfrbp_1 _18813_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1504),
    .D(_00671_),
    .Q_N(_08653_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][22] ));
 sg13g2_dfrbp_1 _18814_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1503),
    .D(_00672_),
    .Q_N(_08652_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][23] ));
 sg13g2_dfrbp_1 _18815_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1502),
    .D(_00673_),
    .Q_N(_08651_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][0] ));
 sg13g2_dfrbp_1 _18816_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1501),
    .D(_00674_),
    .Q_N(_08650_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][1] ));
 sg13g2_dfrbp_1 _18817_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1500),
    .D(_00675_),
    .Q_N(_08649_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][2] ));
 sg13g2_dfrbp_1 _18818_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1499),
    .D(_00676_),
    .Q_N(_08648_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][3] ));
 sg13g2_dfrbp_1 _18819_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1498),
    .D(_00677_),
    .Q_N(_08647_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][4] ));
 sg13g2_dfrbp_1 _18820_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1497),
    .D(_00678_),
    .Q_N(_08646_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][5] ));
 sg13g2_dfrbp_1 _18821_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1496),
    .D(_00679_),
    .Q_N(_08645_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][6] ));
 sg13g2_dfrbp_1 _18822_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1495),
    .D(_00680_),
    .Q_N(_08644_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][7] ));
 sg13g2_dfrbp_1 _18823_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1494),
    .D(_00681_),
    .Q_N(_08643_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][8] ));
 sg13g2_dfrbp_1 _18824_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1493),
    .D(_00682_),
    .Q_N(_08642_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][9] ));
 sg13g2_dfrbp_1 _18825_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1492),
    .D(_00683_),
    .Q_N(_08641_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][10] ));
 sg13g2_dfrbp_1 _18826_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1491),
    .D(_00684_),
    .Q_N(_08640_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][11] ));
 sg13g2_dfrbp_1 _18827_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1490),
    .D(_00685_),
    .Q_N(_08639_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][12] ));
 sg13g2_dfrbp_1 _18828_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1489),
    .D(_00686_),
    .Q_N(_08638_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][13] ));
 sg13g2_dfrbp_1 _18829_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1488),
    .D(_00687_),
    .Q_N(_08637_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][14] ));
 sg13g2_dfrbp_1 _18830_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1487),
    .D(_00688_),
    .Q_N(_08636_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][15] ));
 sg13g2_dfrbp_1 _18831_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1486),
    .D(_00689_),
    .Q_N(_08635_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][24] ));
 sg13g2_dfrbp_1 _18832_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1485),
    .D(_00690_),
    .Q_N(_08634_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][25] ));
 sg13g2_dfrbp_1 _18833_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1484),
    .D(_00691_),
    .Q_N(_08633_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][26] ));
 sg13g2_dfrbp_1 _18834_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1483),
    .D(_00692_),
    .Q_N(_08632_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][27] ));
 sg13g2_dfrbp_1 _18835_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1482),
    .D(_00693_),
    .Q_N(_08631_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][28] ));
 sg13g2_dfrbp_1 _18836_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1481),
    .D(_00694_),
    .Q_N(_08630_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][29] ));
 sg13g2_dfrbp_1 _18837_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1480),
    .D(_00695_),
    .Q_N(_08629_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][30] ));
 sg13g2_dfrbp_1 _18838_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1479),
    .D(_00696_),
    .Q_N(_08628_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][31] ));
 sg13g2_dfrbp_1 _18839_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1478),
    .D(_00697_),
    .Q_N(_08627_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][16] ));
 sg13g2_dfrbp_1 _18840_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1477),
    .D(_00698_),
    .Q_N(_08626_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][17] ));
 sg13g2_dfrbp_1 _18841_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1476),
    .D(_00699_),
    .Q_N(_08625_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][18] ));
 sg13g2_dfrbp_1 _18842_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1475),
    .D(_00700_),
    .Q_N(_08624_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][19] ));
 sg13g2_dfrbp_1 _18843_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1474),
    .D(_00701_),
    .Q_N(_08623_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][20] ));
 sg13g2_dfrbp_1 _18844_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1473),
    .D(_00702_),
    .Q_N(_08622_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][21] ));
 sg13g2_dfrbp_1 _18845_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1472),
    .D(_00703_),
    .Q_N(_08621_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][22] ));
 sg13g2_dfrbp_1 _18846_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1471),
    .D(_00704_),
    .Q_N(_08620_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][23] ));
 sg13g2_dfrbp_1 _18847_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1470),
    .D(_00705_),
    .Q_N(_08619_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][24] ));
 sg13g2_dfrbp_1 _18848_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1469),
    .D(_00706_),
    .Q_N(_08618_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][25] ));
 sg13g2_dfrbp_1 _18849_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1468),
    .D(_00707_),
    .Q_N(_08617_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][26] ));
 sg13g2_dfrbp_1 _18850_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1467),
    .D(_00708_),
    .Q_N(_08616_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][27] ));
 sg13g2_dfrbp_1 _18851_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1466),
    .D(_00709_),
    .Q_N(_08615_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][28] ));
 sg13g2_dfrbp_1 _18852_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1465),
    .D(_00710_),
    .Q_N(_08614_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][29] ));
 sg13g2_dfrbp_1 _18853_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1464),
    .D(_00711_),
    .Q_N(_08613_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][30] ));
 sg13g2_dfrbp_1 _18854_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1463),
    .D(_00712_),
    .Q_N(_08612_),
    .Q(\m_sys.m_ram.m_ram.r_mem[27][31] ));
 sg13g2_dfrbp_1 _18855_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1462),
    .D(_00713_),
    .Q_N(_08611_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][24] ));
 sg13g2_dfrbp_1 _18856_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1461),
    .D(_00714_),
    .Q_N(_08610_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][25] ));
 sg13g2_dfrbp_1 _18857_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1460),
    .D(_00715_),
    .Q_N(_08609_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][26] ));
 sg13g2_dfrbp_1 _18858_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1459),
    .D(_00716_),
    .Q_N(_08608_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][27] ));
 sg13g2_dfrbp_1 _18859_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1458),
    .D(_00717_),
    .Q_N(_08607_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][28] ));
 sg13g2_dfrbp_1 _18860_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1457),
    .D(_00718_),
    .Q_N(_08606_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][29] ));
 sg13g2_dfrbp_1 _18861_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1456),
    .D(_00719_),
    .Q_N(_08605_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][30] ));
 sg13g2_dfrbp_1 _18862_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1455),
    .D(_00720_),
    .Q_N(_08604_),
    .Q(\m_sys.m_ram.m_ram.r_mem[11][31] ));
 sg13g2_dfrbp_1 _18863_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1454),
    .D(_00721_),
    .Q_N(_08603_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][8] ));
 sg13g2_dfrbp_1 _18864_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1453),
    .D(_00722_),
    .Q_N(_08602_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][9] ));
 sg13g2_dfrbp_1 _18865_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1452),
    .D(_00723_),
    .Q_N(_08601_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][10] ));
 sg13g2_dfrbp_1 _18866_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1451),
    .D(_00724_),
    .Q_N(_08600_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][11] ));
 sg13g2_dfrbp_1 _18867_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1450),
    .D(_00725_),
    .Q_N(_08599_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][12] ));
 sg13g2_dfrbp_1 _18868_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1449),
    .D(_00726_),
    .Q_N(_08598_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][13] ));
 sg13g2_dfrbp_1 _18869_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1448),
    .D(_00727_),
    .Q_N(_08597_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][14] ));
 sg13g2_dfrbp_1 _18870_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1447),
    .D(_00728_),
    .Q_N(_08596_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][15] ));
 sg13g2_dfrbp_1 _18871_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1446),
    .D(_00729_),
    .Q_N(_08595_),
    .Q(\m_sys.m_uart.m_tx.r_data[7] ));
 sg13g2_dfrbp_1 _18872_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1444),
    .D(_00730_),
    .Q_N(_08594_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][24] ));
 sg13g2_dfrbp_1 _18873_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1443),
    .D(_00731_),
    .Q_N(_08593_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][25] ));
 sg13g2_dfrbp_1 _18874_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1442),
    .D(_00732_),
    .Q_N(_08592_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][26] ));
 sg13g2_dfrbp_1 _18875_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1441),
    .D(_00733_),
    .Q_N(_08591_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][27] ));
 sg13g2_dfrbp_1 _18876_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1440),
    .D(_00734_),
    .Q_N(_08590_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][28] ));
 sg13g2_dfrbp_1 _18877_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1439),
    .D(_00735_),
    .Q_N(_08589_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][29] ));
 sg13g2_dfrbp_1 _18878_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1438),
    .D(_00736_),
    .Q_N(_08588_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][30] ));
 sg13g2_dfrbp_1 _18879_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1437),
    .D(_00737_),
    .Q_N(_08587_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][31] ));
 sg13g2_dfrbp_1 _18880_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1436),
    .D(_00738_),
    .Q_N(_08586_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][8] ));
 sg13g2_dfrbp_1 _18881_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1435),
    .D(_00739_),
    .Q_N(_08585_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][9] ));
 sg13g2_dfrbp_1 _18882_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1434),
    .D(_00740_),
    .Q_N(_08584_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][10] ));
 sg13g2_dfrbp_1 _18883_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1433),
    .D(_00741_),
    .Q_N(_08583_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][11] ));
 sg13g2_dfrbp_1 _18884_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1432),
    .D(_00742_),
    .Q_N(_08582_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][12] ));
 sg13g2_dfrbp_1 _18885_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1431),
    .D(_00743_),
    .Q_N(_08581_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][13] ));
 sg13g2_dfrbp_1 _18886_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1430),
    .D(_00744_),
    .Q_N(_08580_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][14] ));
 sg13g2_dfrbp_1 _18887_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1429),
    .D(_00745_),
    .Q_N(_08579_),
    .Q(\m_sys.m_ram.m_ram.r_mem[21][15] ));
 sg13g2_dfrbp_1 _18888_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1428),
    .D(_00746_),
    .Q_N(_08578_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][24] ));
 sg13g2_dfrbp_1 _18889_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1427),
    .D(_00747_),
    .Q_N(_08577_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][25] ));
 sg13g2_dfrbp_1 _18890_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1426),
    .D(_00748_),
    .Q_N(_08576_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][26] ));
 sg13g2_dfrbp_1 _18891_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1425),
    .D(_00749_),
    .Q_N(_08575_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][27] ));
 sg13g2_dfrbp_1 _18892_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1424),
    .D(_00750_),
    .Q_N(_08574_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][28] ));
 sg13g2_dfrbp_1 _18893_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1423),
    .D(_00751_),
    .Q_N(_08573_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][29] ));
 sg13g2_dfrbp_1 _18894_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1422),
    .D(_00752_),
    .Q_N(_08572_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][30] ));
 sg13g2_dfrbp_1 _18895_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1421),
    .D(_00753_),
    .Q_N(_08571_),
    .Q(\m_sys.m_ram.m_ram.r_mem[25][31] ));
 sg13g2_dfrbp_1 _18896_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1420),
    .D(_00754_),
    .Q_N(_08570_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][0] ));
 sg13g2_dfrbp_1 _18897_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1419),
    .D(_00755_),
    .Q_N(_08569_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][1] ));
 sg13g2_dfrbp_1 _18898_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1418),
    .D(_00756_),
    .Q_N(_08568_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][2] ));
 sg13g2_dfrbp_1 _18899_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1417),
    .D(_00757_),
    .Q_N(_08567_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][3] ));
 sg13g2_dfrbp_1 _18900_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1416),
    .D(_00758_),
    .Q_N(_08566_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][4] ));
 sg13g2_dfrbp_1 _18901_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1415),
    .D(_00759_),
    .Q_N(_08565_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][5] ));
 sg13g2_dfrbp_1 _18902_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1414),
    .D(_00760_),
    .Q_N(_08564_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][6] ));
 sg13g2_dfrbp_1 _18903_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1413),
    .D(_00761_),
    .Q_N(_08563_),
    .Q(\m_sys.m_ram.m_ram.r_mem[26][7] ));
 sg13g2_dfrbp_1 _18904_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1412),
    .D(_00762_),
    .Q_N(_08562_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][16] ));
 sg13g2_dfrbp_1 _18905_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1411),
    .D(_00763_),
    .Q_N(_08561_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][17] ));
 sg13g2_dfrbp_1 _18906_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1410),
    .D(_00764_),
    .Q_N(_08560_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][18] ));
 sg13g2_dfrbp_1 _18907_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1409),
    .D(_00765_),
    .Q_N(_08559_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][19] ));
 sg13g2_dfrbp_1 _18908_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1408),
    .D(_00766_),
    .Q_N(_08558_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][20] ));
 sg13g2_dfrbp_1 _18909_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1407),
    .D(_00767_),
    .Q_N(_08557_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][21] ));
 sg13g2_dfrbp_1 _18910_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1406),
    .D(_00768_),
    .Q_N(_08556_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][22] ));
 sg13g2_dfrbp_1 _18911_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1405),
    .D(_00769_),
    .Q_N(_08555_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][23] ));
 sg13g2_dfrbp_1 _18912_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1404),
    .D(_00770_),
    .Q_N(_08554_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][8] ));
 sg13g2_dfrbp_1 _18913_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1403),
    .D(_00771_),
    .Q_N(_08553_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][9] ));
 sg13g2_dfrbp_1 _18914_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1402),
    .D(_00772_),
    .Q_N(_08552_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][10] ));
 sg13g2_dfrbp_1 _18915_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1401),
    .D(_00773_),
    .Q_N(_08551_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][11] ));
 sg13g2_dfrbp_1 _18916_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1400),
    .D(_00774_),
    .Q_N(_08550_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][12] ));
 sg13g2_dfrbp_1 _18917_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1399),
    .D(_00775_),
    .Q_N(_08549_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][13] ));
 sg13g2_dfrbp_1 _18918_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1398),
    .D(_00776_),
    .Q_N(_08548_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][14] ));
 sg13g2_dfrbp_1 _18919_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1397),
    .D(_00777_),
    .Q_N(_08547_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][15] ));
 sg13g2_dfrbp_1 _18920_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1396),
    .D(_00778_),
    .Q_N(_08546_),
    .Q(\m_sys.io_b_uart_tx ));
 sg13g2_dfrbp_1 _18921_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1395),
    .D(_00779_),
    .Q_N(_08545_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][24] ));
 sg13g2_dfrbp_1 _18922_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1394),
    .D(_00780_),
    .Q_N(_08544_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][25] ));
 sg13g2_dfrbp_1 _18923_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1393),
    .D(_00781_),
    .Q_N(_08543_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][26] ));
 sg13g2_dfrbp_1 _18924_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1392),
    .D(_00782_),
    .Q_N(_08542_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][27] ));
 sg13g2_dfrbp_1 _18925_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1391),
    .D(_00783_),
    .Q_N(_08541_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][28] ));
 sg13g2_dfrbp_1 _18926_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1390),
    .D(_00784_),
    .Q_N(_08540_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][29] ));
 sg13g2_dfrbp_1 _18927_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1389),
    .D(_00785_),
    .Q_N(_08539_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][30] ));
 sg13g2_dfrbp_1 _18928_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1388),
    .D(_00786_),
    .Q_N(_08538_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][31] ));
 sg13g2_dfrbp_1 _18929_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1387),
    .D(_00787_),
    .Q_N(_08537_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][8] ));
 sg13g2_dfrbp_1 _18930_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1386),
    .D(_00788_),
    .Q_N(_08536_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][9] ));
 sg13g2_dfrbp_1 _18931_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1385),
    .D(_00789_),
    .Q_N(_08535_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][10] ));
 sg13g2_dfrbp_1 _18932_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1384),
    .D(_00790_),
    .Q_N(_08534_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][11] ));
 sg13g2_dfrbp_1 _18933_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1383),
    .D(_00791_),
    .Q_N(_08533_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][12] ));
 sg13g2_dfrbp_1 _18934_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1382),
    .D(_00792_),
    .Q_N(_08532_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][13] ));
 sg13g2_dfrbp_1 _18935_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1381),
    .D(_00793_),
    .Q_N(_08531_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][14] ));
 sg13g2_dfrbp_1 _18936_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1380),
    .D(_00794_),
    .Q_N(_08530_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][15] ));
 sg13g2_dfrbp_1 _18937_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1379),
    .D(_00795_),
    .Q_N(_08529_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][16] ));
 sg13g2_dfrbp_1 _18938_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1378),
    .D(_00796_),
    .Q_N(_08528_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][17] ));
 sg13g2_dfrbp_1 _18939_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1377),
    .D(_00797_),
    .Q_N(_08527_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][18] ));
 sg13g2_dfrbp_1 _18940_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1376),
    .D(_00798_),
    .Q_N(_08526_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][19] ));
 sg13g2_dfrbp_1 _18941_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1375),
    .D(_00799_),
    .Q_N(_08525_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][20] ));
 sg13g2_dfrbp_1 _18942_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1374),
    .D(_00800_),
    .Q_N(_08524_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][21] ));
 sg13g2_dfrbp_1 _18943_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1373),
    .D(_00801_),
    .Q_N(_08523_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][22] ));
 sg13g2_dfrbp_1 _18944_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1372),
    .D(_00802_),
    .Q_N(_08522_),
    .Q(\m_sys.m_ram.m_ram.r_mem[16][23] ));
 sg13g2_dfrbp_1 _18945_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1371),
    .D(_00803_),
    .Q_N(_08521_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][24] ));
 sg13g2_dfrbp_1 _18946_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1370),
    .D(_00804_),
    .Q_N(_08520_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][25] ));
 sg13g2_dfrbp_1 _18947_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1369),
    .D(_00805_),
    .Q_N(_08519_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][26] ));
 sg13g2_dfrbp_1 _18948_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1368),
    .D(_00806_),
    .Q_N(_08518_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][27] ));
 sg13g2_dfrbp_1 _18949_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1367),
    .D(_00807_),
    .Q_N(_08517_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][28] ));
 sg13g2_dfrbp_1 _18950_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1366),
    .D(_00808_),
    .Q_N(_08516_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][29] ));
 sg13g2_dfrbp_1 _18951_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1365),
    .D(_00809_),
    .Q_N(_08515_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][30] ));
 sg13g2_dfrbp_1 _18952_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1364),
    .D(_00810_),
    .Q_N(_08514_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][31] ));
 sg13g2_dfrbp_1 _18953_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1363),
    .D(_00811_),
    .Q_N(_08513_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][16] ));
 sg13g2_dfrbp_1 _18954_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1362),
    .D(_00812_),
    .Q_N(_08512_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][17] ));
 sg13g2_dfrbp_1 _18955_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1361),
    .D(_00813_),
    .Q_N(_08511_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][18] ));
 sg13g2_dfrbp_1 _18956_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1360),
    .D(_00814_),
    .Q_N(_08510_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][19] ));
 sg13g2_dfrbp_1 _18957_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1359),
    .D(_00815_),
    .Q_N(_08509_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][20] ));
 sg13g2_dfrbp_1 _18958_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1358),
    .D(_00816_),
    .Q_N(_08508_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][21] ));
 sg13g2_dfrbp_1 _18959_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1357),
    .D(_00817_),
    .Q_N(_08507_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][22] ));
 sg13g2_dfrbp_1 _18960_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1356),
    .D(_00818_),
    .Q_N(_08506_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][23] ));
 sg13g2_dfrbp_1 _18961_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1355),
    .D(_00819_),
    .Q_N(_08505_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][0] ));
 sg13g2_dfrbp_1 _18962_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1354),
    .D(_00820_),
    .Q_N(_08504_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][1] ));
 sg13g2_dfrbp_1 _18963_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1353),
    .D(_00821_),
    .Q_N(_08503_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][2] ));
 sg13g2_dfrbp_1 _18964_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1352),
    .D(_00822_),
    .Q_N(_08502_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][3] ));
 sg13g2_dfrbp_1 _18965_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1351),
    .D(_00823_),
    .Q_N(_08501_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][4] ));
 sg13g2_dfrbp_1 _18966_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1350),
    .D(_00824_),
    .Q_N(_08500_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][5] ));
 sg13g2_dfrbp_1 _18967_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1349),
    .D(_00825_),
    .Q_N(_08499_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][6] ));
 sg13g2_dfrbp_1 _18968_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1348),
    .D(_00826_),
    .Q_N(_08498_),
    .Q(\m_sys.m_ram.m_ram.r_mem[9][7] ));
 sg13g2_dfrbp_1 _18969_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1347),
    .D(_00827_),
    .Q_N(_08497_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][0] ));
 sg13g2_dfrbp_1 _18970_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1346),
    .D(_00828_),
    .Q_N(_08496_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][1] ));
 sg13g2_dfrbp_1 _18971_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1345),
    .D(_00829_),
    .Q_N(_08495_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][2] ));
 sg13g2_dfrbp_1 _18972_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1344),
    .D(_00830_),
    .Q_N(_08494_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][3] ));
 sg13g2_dfrbp_1 _18973_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1343),
    .D(_00831_),
    .Q_N(_08493_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][4] ));
 sg13g2_dfrbp_1 _18974_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1342),
    .D(_00832_),
    .Q_N(_08492_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][5] ));
 sg13g2_dfrbp_1 _18975_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1341),
    .D(_00833_),
    .Q_N(_08491_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][6] ));
 sg13g2_dfrbp_1 _18976_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1340),
    .D(_00834_),
    .Q_N(_08490_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][7] ));
 sg13g2_dfrbp_1 _18977_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1339),
    .D(_00835_),
    .Q_N(_08489_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][8] ));
 sg13g2_dfrbp_1 _18978_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1338),
    .D(_00836_),
    .Q_N(_08488_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][9] ));
 sg13g2_dfrbp_1 _18979_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1337),
    .D(_00837_),
    .Q_N(_08487_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][10] ));
 sg13g2_dfrbp_1 _18980_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1336),
    .D(_00838_),
    .Q_N(_08486_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][11] ));
 sg13g2_dfrbp_1 _18981_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1335),
    .D(_00839_),
    .Q_N(_08485_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][12] ));
 sg13g2_dfrbp_1 _18982_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1334),
    .D(_00840_),
    .Q_N(_08484_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][13] ));
 sg13g2_dfrbp_1 _18983_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1333),
    .D(_00841_),
    .Q_N(_08483_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][14] ));
 sg13g2_dfrbp_1 _18984_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1332),
    .D(_00842_),
    .Q_N(_08482_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][15] ));
 sg13g2_dfrbp_1 _18985_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1331),
    .D(_00843_),
    .Q_N(_08481_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][24] ));
 sg13g2_dfrbp_1 _18986_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1330),
    .D(_00844_),
    .Q_N(_08480_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][25] ));
 sg13g2_dfrbp_1 _18987_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1329),
    .D(_00845_),
    .Q_N(_08479_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][26] ));
 sg13g2_dfrbp_1 _18988_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1328),
    .D(_00846_),
    .Q_N(_08478_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][27] ));
 sg13g2_dfrbp_1 _18989_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1327),
    .D(_00847_),
    .Q_N(_08477_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][28] ));
 sg13g2_dfrbp_1 _18990_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1326),
    .D(_00848_),
    .Q_N(_08476_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][29] ));
 sg13g2_dfrbp_1 _18991_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1325),
    .D(_00849_),
    .Q_N(_08475_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][30] ));
 sg13g2_dfrbp_1 _18992_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1324),
    .D(_00850_),
    .Q_N(_08474_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][31] ));
 sg13g2_dfrbp_1 _18993_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1323),
    .D(_00851_),
    .Q_N(_08473_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][0] ));
 sg13g2_dfrbp_1 _18994_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1322),
    .D(_00852_),
    .Q_N(_08472_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][1] ));
 sg13g2_dfrbp_1 _18995_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1321),
    .D(_00853_),
    .Q_N(_08471_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][2] ));
 sg13g2_dfrbp_1 _18996_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1320),
    .D(_00854_),
    .Q_N(_08470_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][3] ));
 sg13g2_dfrbp_1 _18997_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1319),
    .D(_00855_),
    .Q_N(_08469_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][4] ));
 sg13g2_dfrbp_1 _18998_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1318),
    .D(_00856_),
    .Q_N(_08468_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][5] ));
 sg13g2_dfrbp_1 _18999_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1317),
    .D(_00857_),
    .Q_N(_08467_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][6] ));
 sg13g2_dfrbp_1 _19000_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1316),
    .D(_00858_),
    .Q_N(_08466_),
    .Q(\m_sys.m_ram.m_ram.r_mem[1][7] ));
 sg13g2_dfrbp_1 _19001_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1315),
    .D(_00859_),
    .Q_N(_08465_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][16] ));
 sg13g2_dfrbp_1 _19002_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1314),
    .D(_00860_),
    .Q_N(_08464_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][17] ));
 sg13g2_dfrbp_1 _19003_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1313),
    .D(_00861_),
    .Q_N(_08463_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][18] ));
 sg13g2_dfrbp_1 _19004_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1312),
    .D(_00862_),
    .Q_N(_08462_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][19] ));
 sg13g2_dfrbp_1 _19005_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1311),
    .D(_00863_),
    .Q_N(_08461_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][20] ));
 sg13g2_dfrbp_1 _19006_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1310),
    .D(_00864_),
    .Q_N(_08460_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][21] ));
 sg13g2_dfrbp_1 _19007_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1309),
    .D(_00865_),
    .Q_N(_08459_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][22] ));
 sg13g2_dfrbp_1 _19008_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1308),
    .D(_00866_),
    .Q_N(_08458_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][23] ));
 sg13g2_dfrbp_1 _19009_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1307),
    .D(_00867_),
    .Q_N(_08457_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][8] ));
 sg13g2_dfrbp_1 _19010_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1306),
    .D(_00868_),
    .Q_N(_08456_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][9] ));
 sg13g2_dfrbp_1 _19011_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1305),
    .D(_00869_),
    .Q_N(_08455_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][10] ));
 sg13g2_dfrbp_1 _19012_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1304),
    .D(_00870_),
    .Q_N(_08454_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][11] ));
 sg13g2_dfrbp_1 _19013_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1303),
    .D(_00871_),
    .Q_N(_08453_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][12] ));
 sg13g2_dfrbp_1 _19014_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1302),
    .D(_00872_),
    .Q_N(_08452_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][13] ));
 sg13g2_dfrbp_1 _19015_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1301),
    .D(_00873_),
    .Q_N(_08451_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][14] ));
 sg13g2_dfrbp_1 _19016_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1300),
    .D(_00874_),
    .Q_N(_08450_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][15] ));
 sg13g2_dfrbp_1 _19017_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1299),
    .D(_00875_),
    .Q_N(_08449_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][16] ));
 sg13g2_dfrbp_1 _19018_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1298),
    .D(_00876_),
    .Q_N(_08448_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][17] ));
 sg13g2_dfrbp_1 _19019_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1297),
    .D(_00877_),
    .Q_N(_08447_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][18] ));
 sg13g2_dfrbp_1 _19020_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1296),
    .D(_00878_),
    .Q_N(_08446_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][19] ));
 sg13g2_dfrbp_1 _19021_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1295),
    .D(_00879_),
    .Q_N(_08445_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][20] ));
 sg13g2_dfrbp_1 _19022_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1294),
    .D(_00880_),
    .Q_N(_08444_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][21] ));
 sg13g2_dfrbp_1 _19023_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1293),
    .D(_00881_),
    .Q_N(_08443_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][22] ));
 sg13g2_dfrbp_1 _19024_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1292),
    .D(_00882_),
    .Q_N(_08442_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][23] ));
 sg13g2_dfrbp_1 _19025_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1291),
    .D(_00883_),
    .Q_N(_08441_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][8] ));
 sg13g2_dfrbp_1 _19026_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1290),
    .D(_00884_),
    .Q_N(_08440_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][9] ));
 sg13g2_dfrbp_1 _19027_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1289),
    .D(_00885_),
    .Q_N(_08439_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][10] ));
 sg13g2_dfrbp_1 _19028_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1288),
    .D(_00886_),
    .Q_N(_08438_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][11] ));
 sg13g2_dfrbp_1 _19029_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1287),
    .D(_00887_),
    .Q_N(_08437_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][12] ));
 sg13g2_dfrbp_1 _19030_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1286),
    .D(_00888_),
    .Q_N(_08436_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][13] ));
 sg13g2_dfrbp_1 _19031_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1285),
    .D(_00889_),
    .Q_N(_08435_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][14] ));
 sg13g2_dfrbp_1 _19032_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1284),
    .D(_00890_),
    .Q_N(_08434_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][15] ));
 sg13g2_dfrbp_1 _19033_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1283),
    .D(_00891_),
    .Q_N(_08433_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][0] ));
 sg13g2_dfrbp_1 _19034_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1282),
    .D(_00892_),
    .Q_N(_08432_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][1] ));
 sg13g2_dfrbp_1 _19035_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1281),
    .D(_00893_),
    .Q_N(_08431_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][2] ));
 sg13g2_dfrbp_1 _19036_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1280),
    .D(_00894_),
    .Q_N(_08430_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][3] ));
 sg13g2_dfrbp_1 _19037_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1279),
    .D(_00895_),
    .Q_N(_08429_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][4] ));
 sg13g2_dfrbp_1 _19038_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1278),
    .D(_00896_),
    .Q_N(_08428_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][5] ));
 sg13g2_dfrbp_1 _19039_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1277),
    .D(_00897_),
    .Q_N(_08427_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][6] ));
 sg13g2_dfrbp_1 _19040_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1276),
    .D(_00898_),
    .Q_N(_08426_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][7] ));
 sg13g2_dfrbp_1 _19041_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1275),
    .D(_00899_),
    .Q_N(_08425_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][16] ));
 sg13g2_dfrbp_1 _19042_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1274),
    .D(_00900_),
    .Q_N(_08424_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][17] ));
 sg13g2_dfrbp_1 _19043_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1273),
    .D(_00901_),
    .Q_N(_08423_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][18] ));
 sg13g2_dfrbp_1 _19044_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1272),
    .D(_00902_),
    .Q_N(_08422_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][19] ));
 sg13g2_dfrbp_1 _19045_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1271),
    .D(_00903_),
    .Q_N(_08421_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][20] ));
 sg13g2_dfrbp_1 _19046_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1270),
    .D(_00904_),
    .Q_N(_08420_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][21] ));
 sg13g2_dfrbp_1 _19047_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1269),
    .D(_00905_),
    .Q_N(_08419_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][22] ));
 sg13g2_dfrbp_1 _19048_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1268),
    .D(_00906_),
    .Q_N(_08418_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][23] ));
 sg13g2_dfrbp_1 _19049_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1267),
    .D(_00907_),
    .Q_N(_08417_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][8] ));
 sg13g2_dfrbp_1 _19050_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1266),
    .D(_00908_),
    .Q_N(_08416_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][9] ));
 sg13g2_dfrbp_1 _19051_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1265),
    .D(_00909_),
    .Q_N(_08415_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][10] ));
 sg13g2_dfrbp_1 _19052_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1264),
    .D(_00910_),
    .Q_N(_08414_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][11] ));
 sg13g2_dfrbp_1 _19053_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1263),
    .D(_00911_),
    .Q_N(_08413_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][12] ));
 sg13g2_dfrbp_1 _19054_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1262),
    .D(_00912_),
    .Q_N(_08412_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][13] ));
 sg13g2_dfrbp_1 _19055_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1261),
    .D(_00913_),
    .Q_N(_08411_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][14] ));
 sg13g2_dfrbp_1 _19056_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1260),
    .D(_00914_),
    .Q_N(_08410_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][15] ));
 sg13g2_dfrbp_1 _19057_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1259),
    .D(_00915_),
    .Q_N(_08409_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][0] ));
 sg13g2_dfrbp_1 _19058_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1258),
    .D(_00916_),
    .Q_N(_08408_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][1] ));
 sg13g2_dfrbp_1 _19059_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1257),
    .D(_00917_),
    .Q_N(_08407_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][2] ));
 sg13g2_dfrbp_1 _19060_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1256),
    .D(_00918_),
    .Q_N(_08406_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][3] ));
 sg13g2_dfrbp_1 _19061_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1255),
    .D(_00919_),
    .Q_N(_08405_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][4] ));
 sg13g2_dfrbp_1 _19062_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1254),
    .D(_00920_),
    .Q_N(_08404_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][5] ));
 sg13g2_dfrbp_1 _19063_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1253),
    .D(_00921_),
    .Q_N(_08403_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][6] ));
 sg13g2_dfrbp_1 _19064_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1252),
    .D(_00922_),
    .Q_N(_08402_),
    .Q(\m_sys.m_ram.m_ram.r_mem[30][7] ));
 sg13g2_dfrbp_1 _19065_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1251),
    .D(_00923_),
    .Q_N(_08401_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][16] ));
 sg13g2_dfrbp_1 _19066_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1250),
    .D(_00924_),
    .Q_N(_08400_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][17] ));
 sg13g2_dfrbp_1 _19067_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1249),
    .D(_00925_),
    .Q_N(_08399_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][18] ));
 sg13g2_dfrbp_1 _19068_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1248),
    .D(_00926_),
    .Q_N(_08398_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][19] ));
 sg13g2_dfrbp_1 _19069_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1247),
    .D(_00927_),
    .Q_N(_08397_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][20] ));
 sg13g2_dfrbp_1 _19070_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1246),
    .D(_00928_),
    .Q_N(_08396_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][21] ));
 sg13g2_dfrbp_1 _19071_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1245),
    .D(_00929_),
    .Q_N(_08395_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][22] ));
 sg13g2_dfrbp_1 _19072_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1244),
    .D(_00930_),
    .Q_N(_08394_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][23] ));
 sg13g2_dfrbp_1 _19073_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1243),
    .D(_00931_),
    .Q_N(_08393_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][8] ));
 sg13g2_dfrbp_1 _19074_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1242),
    .D(_00932_),
    .Q_N(_08392_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][9] ));
 sg13g2_dfrbp_1 _19075_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1241),
    .D(_00933_),
    .Q_N(_08391_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][10] ));
 sg13g2_dfrbp_1 _19076_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1240),
    .D(_00934_),
    .Q_N(_08390_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][11] ));
 sg13g2_dfrbp_1 _19077_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1239),
    .D(_00935_),
    .Q_N(_08389_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][12] ));
 sg13g2_dfrbp_1 _19078_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1238),
    .D(_00936_),
    .Q_N(_08388_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][13] ));
 sg13g2_dfrbp_1 _19079_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1237),
    .D(_00937_),
    .Q_N(_08387_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][14] ));
 sg13g2_dfrbp_1 _19080_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1236),
    .D(_00938_),
    .Q_N(_08386_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][15] ));
 sg13g2_dfrbp_1 _19081_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1235),
    .D(_00939_),
    .Q_N(_08385_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][0] ));
 sg13g2_dfrbp_1 _19082_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1234),
    .D(_00940_),
    .Q_N(_08384_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][1] ));
 sg13g2_dfrbp_1 _19083_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1233),
    .D(_00941_),
    .Q_N(_08383_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][2] ));
 sg13g2_dfrbp_1 _19084_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1232),
    .D(_00942_),
    .Q_N(_08382_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][3] ));
 sg13g2_dfrbp_1 _19085_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1231),
    .D(_00943_),
    .Q_N(_08381_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][4] ));
 sg13g2_dfrbp_1 _19086_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1230),
    .D(_00944_),
    .Q_N(_08380_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][5] ));
 sg13g2_dfrbp_1 _19087_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1229),
    .D(_00945_),
    .Q_N(_08379_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][6] ));
 sg13g2_dfrbp_1 _19088_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1228),
    .D(_00946_),
    .Q_N(_08378_),
    .Q(\m_sys.m_ram.m_ram.r_mem[2][7] ));
 sg13g2_dfrbp_1 _19089_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1227),
    .D(_00947_),
    .Q_N(_08377_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][16] ));
 sg13g2_dfrbp_1 _19090_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1226),
    .D(_00948_),
    .Q_N(_08376_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][17] ));
 sg13g2_dfrbp_1 _19091_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1225),
    .D(_00949_),
    .Q_N(_08375_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][18] ));
 sg13g2_dfrbp_1 _19092_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1224),
    .D(_00950_),
    .Q_N(_08374_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][19] ));
 sg13g2_dfrbp_1 _19093_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1223),
    .D(_00951_),
    .Q_N(_08373_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][20] ));
 sg13g2_dfrbp_1 _19094_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1222),
    .D(_00952_),
    .Q_N(_08372_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][21] ));
 sg13g2_dfrbp_1 _19095_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1221),
    .D(_00953_),
    .Q_N(_08371_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][22] ));
 sg13g2_dfrbp_1 _19096_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1220),
    .D(_00954_),
    .Q_N(_08370_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][23] ));
 sg13g2_dfrbp_1 _19097_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1219),
    .D(_00955_),
    .Q_N(_08369_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][8] ));
 sg13g2_dfrbp_1 _19098_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1218),
    .D(_00956_),
    .Q_N(_08368_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][9] ));
 sg13g2_dfrbp_1 _19099_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1217),
    .D(_00957_),
    .Q_N(_08367_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][10] ));
 sg13g2_dfrbp_1 _19100_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1216),
    .D(_00958_),
    .Q_N(_08366_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][11] ));
 sg13g2_dfrbp_1 _19101_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1215),
    .D(_00959_),
    .Q_N(_08365_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][12] ));
 sg13g2_dfrbp_1 _19102_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1214),
    .D(_00960_),
    .Q_N(_08364_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][13] ));
 sg13g2_dfrbp_1 _19103_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1213),
    .D(_00961_),
    .Q_N(_08363_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][14] ));
 sg13g2_dfrbp_1 _19104_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1212),
    .D(_00962_),
    .Q_N(_08362_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][15] ));
 sg13g2_dfrbp_1 _19105_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1211),
    .D(_00963_),
    .Q_N(_08361_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][0] ));
 sg13g2_dfrbp_1 _19106_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1210),
    .D(_00964_),
    .Q_N(_08360_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][1] ));
 sg13g2_dfrbp_1 _19107_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1209),
    .D(_00965_),
    .Q_N(_08359_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][2] ));
 sg13g2_dfrbp_1 _19108_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1208),
    .D(_00966_),
    .Q_N(_08358_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][3] ));
 sg13g2_dfrbp_1 _19109_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1207),
    .D(_00967_),
    .Q_N(_08357_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][4] ));
 sg13g2_dfrbp_1 _19110_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1206),
    .D(_00968_),
    .Q_N(_08356_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][5] ));
 sg13g2_dfrbp_1 _19111_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1205),
    .D(_00969_),
    .Q_N(_08355_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][6] ));
 sg13g2_dfrbp_1 _19112_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1204),
    .D(_00970_),
    .Q_N(_08354_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][7] ));
 sg13g2_dfrbp_1 _19113_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1203),
    .D(_00971_),
    .Q_N(_08353_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][8] ));
 sg13g2_dfrbp_1 _19114_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1202),
    .D(_00972_),
    .Q_N(_08352_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][9] ));
 sg13g2_dfrbp_1 _19115_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1201),
    .D(_00973_),
    .Q_N(_08351_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][10] ));
 sg13g2_dfrbp_1 _19116_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1200),
    .D(_00974_),
    .Q_N(_08350_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][11] ));
 sg13g2_dfrbp_1 _19117_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1199),
    .D(_00975_),
    .Q_N(_08349_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][12] ));
 sg13g2_dfrbp_1 _19118_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1198),
    .D(_00976_),
    .Q_N(_08348_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][13] ));
 sg13g2_dfrbp_1 _19119_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1197),
    .D(_00977_),
    .Q_N(_08347_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][14] ));
 sg13g2_dfrbp_1 _19120_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1196),
    .D(_00978_),
    .Q_N(_08346_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][15] ));
 sg13g2_dfrbp_1 _19121_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1195),
    .D(_00979_),
    .Q_N(_08345_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][0] ));
 sg13g2_dfrbp_1 _19122_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1194),
    .D(_00980_),
    .Q_N(_08344_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][1] ));
 sg13g2_dfrbp_1 _19123_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1193),
    .D(_00981_),
    .Q_N(_08343_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][2] ));
 sg13g2_dfrbp_1 _19124_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1192),
    .D(_00982_),
    .Q_N(_08342_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][3] ));
 sg13g2_dfrbp_1 _19125_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1191),
    .D(_00983_),
    .Q_N(_08341_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][4] ));
 sg13g2_dfrbp_1 _19126_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1190),
    .D(_00984_),
    .Q_N(_08340_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][5] ));
 sg13g2_dfrbp_1 _19127_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1189),
    .D(_00985_),
    .Q_N(_08339_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][6] ));
 sg13g2_dfrbp_1 _19128_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1188),
    .D(_00986_),
    .Q_N(_08338_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][7] ));
 sg13g2_dfrbp_1 _19129_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1187),
    .D(_00987_),
    .Q_N(_08337_),
    .Q(\m_sys.m_uart.m_tx.r_data[0] ));
 sg13g2_dfrbp_1 _19130_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1186),
    .D(net2557),
    .Q_N(_08336_),
    .Q(\m_sys.m_uart.m_tx.r_data[1] ));
 sg13g2_dfrbp_1 _19131_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1185),
    .D(_00989_),
    .Q_N(_08335_),
    .Q(\m_sys.m_uart.m_tx.r_data[2] ));
 sg13g2_dfrbp_1 _19132_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1184),
    .D(_00990_),
    .Q_N(_08334_),
    .Q(\m_sys.m_uart.m_tx.r_data[3] ));
 sg13g2_dfrbp_1 _19133_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1183),
    .D(net2703),
    .Q_N(_08333_),
    .Q(\m_sys.m_uart.m_tx.r_data[4] ));
 sg13g2_dfrbp_1 _19134_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1182),
    .D(_00992_),
    .Q_N(_08332_),
    .Q(\m_sys.m_uart.m_tx.r_data[5] ));
 sg13g2_dfrbp_1 _19135_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1181),
    .D(net2285),
    .Q_N(_08331_),
    .Q(\m_sys.m_uart.m_tx.r_data[6] ));
 sg13g2_dfrbp_1 _19136_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1180),
    .D(_00994_),
    .Q_N(_08330_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][24] ));
 sg13g2_dfrbp_1 _19137_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1179),
    .D(_00995_),
    .Q_N(_08329_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][25] ));
 sg13g2_dfrbp_1 _19138_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1178),
    .D(_00996_),
    .Q_N(_08328_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][26] ));
 sg13g2_dfrbp_1 _19139_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1177),
    .D(_00997_),
    .Q_N(_08327_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][27] ));
 sg13g2_dfrbp_1 _19140_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1176),
    .D(_00998_),
    .Q_N(_08326_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][28] ));
 sg13g2_dfrbp_1 _19141_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1175),
    .D(_00999_),
    .Q_N(_08325_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][29] ));
 sg13g2_dfrbp_1 _19142_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1174),
    .D(_01000_),
    .Q_N(_08324_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][30] ));
 sg13g2_dfrbp_1 _19143_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1173),
    .D(_01001_),
    .Q_N(_08323_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][31] ));
 sg13g2_dfrbp_1 _19144_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1172),
    .D(_01002_),
    .Q_N(_08322_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][16] ));
 sg13g2_dfrbp_1 _19145_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1171),
    .D(_01003_),
    .Q_N(_08321_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][17] ));
 sg13g2_dfrbp_1 _19146_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1170),
    .D(_01004_),
    .Q_N(_08320_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][18] ));
 sg13g2_dfrbp_1 _19147_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1169),
    .D(_01005_),
    .Q_N(_08319_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][19] ));
 sg13g2_dfrbp_1 _19148_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1168),
    .D(_01006_),
    .Q_N(_08318_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][20] ));
 sg13g2_dfrbp_1 _19149_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1167),
    .D(_01007_),
    .Q_N(_08317_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][21] ));
 sg13g2_dfrbp_1 _19150_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1166),
    .D(_01008_),
    .Q_N(_08316_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][22] ));
 sg13g2_dfrbp_1 _19151_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1165),
    .D(_01009_),
    .Q_N(_08315_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][23] ));
 sg13g2_dfrbp_1 _19152_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1164),
    .D(_01010_),
    .Q_N(_08314_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][24] ));
 sg13g2_dfrbp_1 _19153_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1163),
    .D(_01011_),
    .Q_N(_08313_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][25] ));
 sg13g2_dfrbp_1 _19154_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1162),
    .D(_01012_),
    .Q_N(_08312_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][26] ));
 sg13g2_dfrbp_1 _19155_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1161),
    .D(_01013_),
    .Q_N(_08311_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][27] ));
 sg13g2_dfrbp_1 _19156_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1160),
    .D(_01014_),
    .Q_N(_08310_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][28] ));
 sg13g2_dfrbp_1 _19157_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1159),
    .D(_01015_),
    .Q_N(_08309_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][29] ));
 sg13g2_dfrbp_1 _19158_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1158),
    .D(_01016_),
    .Q_N(_08308_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][30] ));
 sg13g2_dfrbp_1 _19159_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1157),
    .D(_01017_),
    .Q_N(_08307_),
    .Q(\m_sys.m_ram.m_ram.r_mem[29][31] ));
 sg13g2_dfrbp_1 _19160_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1156),
    .D(_01018_),
    .Q_N(_08306_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][0] ));
 sg13g2_dfrbp_1 _19161_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1155),
    .D(_01019_),
    .Q_N(_08305_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][1] ));
 sg13g2_dfrbp_1 _19162_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1154),
    .D(_01020_),
    .Q_N(_08304_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][2] ));
 sg13g2_dfrbp_1 _19163_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1153),
    .D(_01021_),
    .Q_N(_08303_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][3] ));
 sg13g2_dfrbp_1 _19164_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1152),
    .D(_01022_),
    .Q_N(_08302_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][4] ));
 sg13g2_dfrbp_1 _19165_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1151),
    .D(_01023_),
    .Q_N(_08301_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][5] ));
 sg13g2_dfrbp_1 _19166_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1150),
    .D(_01024_),
    .Q_N(_08300_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][6] ));
 sg13g2_dfrbp_1 _19167_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1149),
    .D(_01025_),
    .Q_N(_08299_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][7] ));
 sg13g2_dfrbp_1 _19168_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1148),
    .D(_01026_),
    .Q_N(_08298_),
    .Q(\m_sys.m_bootloader.r_cstate[0] ));
 sg13g2_dfrbp_1 _19169_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1146),
    .D(_01027_),
    .Q_N(_08297_),
    .Q(\m_sys.m_bootloader.r_cstate[1] ));
 sg13g2_dfrbp_1 _19170_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1144),
    .D(_01028_),
    .Q_N(_08296_),
    .Q(\m_sys.m_bootloader.r_cstate[2] ));
 sg13g2_dfrbp_1 _19171_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1142),
    .D(_01029_),
    .Q_N(_08295_),
    .Q(\m_sys.m_bootloader.r_cstate[3] ));
 sg13g2_dfrbp_1 _19172_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1132),
    .D(_01030_),
    .Q_N(_00024_),
    .Q(\m_sys.m_bootloader.r_cstate[4] ));
 sg13g2_dfrbp_1 _19173_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1130),
    .D(_01031_),
    .Q_N(_00146_),
    .Q(\m_sys.m_bootloader.r_num_cnt[0] ));
 sg13g2_dfrbp_1 _19174_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1128),
    .D(net2879),
    .Q_N(_08294_),
    .Q(\m_sys.m_bootloader.r_num_cnt[1] ));
 sg13g2_dfrbp_1 _19175_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1126),
    .D(_01033_),
    .Q_N(_08293_),
    .Q(\m_sys.m_bootloader.r_num_cnt[2] ));
 sg13g2_dfrbp_1 _19176_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1108),
    .D(_01034_),
    .Q_N(_08292_),
    .Q(\m_sys.m_bootloader.r_num_cnt[3] ));
 sg13g2_dfrbp_1 _19177_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1106),
    .D(_01035_),
    .Q_N(_08291_),
    .Q(\m_sys.m_bootloader.r_num_cnt[4] ));
 sg13g2_dfrbp_1 _19178_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1104),
    .D(_01036_),
    .Q_N(_08290_),
    .Q(\m_sys.m_bootloader.r_num_cnt[5] ));
 sg13g2_dfrbp_1 _19179_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1102),
    .D(_01037_),
    .Q_N(_08289_),
    .Q(\m_sys.m_bootloader.r_num_cnt[6] ));
 sg13g2_dfrbp_1 _19180_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1100),
    .D(_01038_),
    .Q_N(_08288_),
    .Q(\m_sys.m_bootloader.r_num_cnt[7] ));
 sg13g2_dfrbp_1 _19181_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1098),
    .D(_01039_),
    .Q_N(_00046_),
    .Q(\m_sys.r_valid ));
 sg13g2_dfrbp_1 _19182_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1097),
    .D(net3327),
    .Q_N(_08287_),
    .Q(\m_sys._m_bootloader_io_b_mem_wdata[0] ));
 sg13g2_dfrbp_1 _19183_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1095),
    .D(_01041_),
    .Q_N(_08286_),
    .Q(\m_sys._m_bootloader_io_b_mem_wdata[1] ));
 sg13g2_dfrbp_1 _19184_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1093),
    .D(net3340),
    .Q_N(_08285_),
    .Q(\m_sys._m_bootloader_io_b_mem_wdata[2] ));
 sg13g2_dfrbp_1 _19185_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1091),
    .D(_01043_),
    .Q_N(_08284_),
    .Q(\m_sys._m_bootloader_io_b_mem_wdata[3] ));
 sg13g2_dfrbp_1 _19186_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1089),
    .D(_01044_),
    .Q_N(_08283_),
    .Q(\m_sys._m_bootloader_io_b_mem_wdata[4] ));
 sg13g2_dfrbp_1 _19187_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1087),
    .D(_01045_),
    .Q_N(_08282_),
    .Q(\m_sys._m_bootloader_io_b_mem_wdata[5] ));
 sg13g2_dfrbp_1 _19188_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1085),
    .D(net3287),
    .Q_N(_08281_),
    .Q(\m_sys._m_bootloader_io_b_mem_wdata[6] ));
 sg13g2_dfrbp_1 _19189_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1083),
    .D(_01047_),
    .Q_N(_08280_),
    .Q(\m_sys._m_bootloader_io_b_mem_wdata[7] ));
 sg13g2_dfrbp_1 _19190_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1065),
    .D(net2906),
    .Q_N(_08279_),
    .Q(\m_sys.m_bootloader.r_num[0] ));
 sg13g2_dfrbp_1 _19191_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1064),
    .D(_01049_),
    .Q_N(_08278_),
    .Q(\m_sys.m_bootloader.r_num[1] ));
 sg13g2_dfrbp_1 _19192_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1063),
    .D(_01050_),
    .Q_N(_08277_),
    .Q(\m_sys.m_bootloader.r_num[2] ));
 sg13g2_dfrbp_1 _19193_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1062),
    .D(_01051_),
    .Q_N(_08276_),
    .Q(\m_sys.m_bootloader.r_num[3] ));
 sg13g2_dfrbp_1 _19194_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1061),
    .D(net2800),
    .Q_N(_08275_),
    .Q(\m_sys.m_bootloader.r_num[4] ));
 sg13g2_dfrbp_1 _19195_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1060),
    .D(_01053_),
    .Q_N(_08274_),
    .Q(\m_sys.m_bootloader.r_num[5] ));
 sg13g2_dfrbp_1 _19196_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1059),
    .D(_01054_),
    .Q_N(_08273_),
    .Q(\m_sys.m_bootloader.r_num[6] ));
 sg13g2_dfrbp_1 _19197_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1058),
    .D(_01055_),
    .Q_N(_08272_),
    .Q(\m_sys.m_bootloader.r_num[7] ));
 sg13g2_dfrbp_1 _19198_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1057),
    .D(net2045),
    .Q_N(_08271_),
    .Q(\m_sys.m_bootloader._GEN_22[0] ));
 sg13g2_dfrbp_1 _19199_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1056),
    .D(net1993),
    .Q_N(_08270_),
    .Q(\m_sys.m_bootloader._GEN_22[1] ));
 sg13g2_dfrbp_1 _19200_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1055),
    .D(_01058_),
    .Q_N(_08269_),
    .Q(\m_sys.m_bootloader._GEN_22[2] ));
 sg13g2_dfrbp_1 _19201_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1054),
    .D(_01059_),
    .Q_N(_08268_),
    .Q(\m_sys.m_bootloader._GEN_22[3] ));
 sg13g2_dfrbp_1 _19202_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1053),
    .D(_01060_),
    .Q_N(_08267_),
    .Q(\m_sys.m_bootloader._GEN_22[4] ));
 sg13g2_dfrbp_1 _19203_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1052),
    .D(_01061_),
    .Q_N(_08266_),
    .Q(\m_sys.m_bootloader._GEN_22[5] ));
 sg13g2_dfrbp_1 _19204_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1051),
    .D(_01062_),
    .Q_N(_08265_),
    .Q(\m_sys.m_bootloader._GEN_22[6] ));
 sg13g2_dfrbp_1 _19205_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1050),
    .D(_01063_),
    .Q_N(_08264_),
    .Q(\m_sys.m_bootloader._GEN_22[7] ));
 sg13g2_dfrbp_1 _19206_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1049),
    .D(net2933),
    .Q_N(_08263_),
    .Q(\m_sys.m_bootloader._GEN_22[8] ));
 sg13g2_dfrbp_1 _19207_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1048),
    .D(_01065_),
    .Q_N(_08262_),
    .Q(\m_sys.m_bootloader._GEN_22[9] ));
 sg13g2_dfrbp_1 _19208_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1047),
    .D(net2614),
    .Q_N(_08261_),
    .Q(\m_sys.m_bootloader._GEN_22[10] ));
 sg13g2_dfrbp_1 _19209_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1046),
    .D(_01067_),
    .Q_N(_08260_),
    .Q(\m_sys.m_bootloader._GEN_22[11] ));
 sg13g2_dfrbp_1 _19210_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1045),
    .D(net3145),
    .Q_N(_08259_),
    .Q(\m_sys.m_bootloader.r_offset_0[0] ));
 sg13g2_dfrbp_1 _19211_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1044),
    .D(_01069_),
    .Q_N(_08258_),
    .Q(\m_sys.m_bootloader.r_offset_0[1] ));
 sg13g2_dfrbp_1 _19212_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1043),
    .D(_01070_),
    .Q_N(_08257_),
    .Q(\m_sys.m_bootloader.r_offset_0[2] ));
 sg13g2_dfrbp_1 _19213_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1042),
    .D(_01071_),
    .Q_N(_08256_),
    .Q(\m_sys.m_bootloader.r_offset_0[3] ));
 sg13g2_dfrbp_1 _19214_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1041),
    .D(_01072_),
    .Q_N(_08255_),
    .Q(\m_sys.m_bootloader.r_offset_0[4] ));
 sg13g2_dfrbp_1 _19215_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1040),
    .D(_01073_),
    .Q_N(_08254_),
    .Q(\m_sys.m_bootloader.r_offset_0[5] ));
 sg13g2_dfrbp_1 _19216_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1039),
    .D(_01074_),
    .Q_N(_00033_),
    .Q(\m_sys.m_bootloader.r_offset_0[6] ));
 sg13g2_dfrbp_1 _19217_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1038),
    .D(_01075_),
    .Q_N(_08253_),
    .Q(\m_sys.m_bootloader.r_offset_0[7] ));
 sg13g2_dfrbp_1 _19218_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1037),
    .D(net3068),
    .Q_N(_08252_),
    .Q(\m_sys.m_bootloader.r_offset_1[0] ));
 sg13g2_dfrbp_1 _19219_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1036),
    .D(_01077_),
    .Q_N(_08251_),
    .Q(\m_sys.m_bootloader.r_offset_1[1] ));
 sg13g2_dfrbp_1 _19220_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1035),
    .D(_01078_),
    .Q_N(_08250_),
    .Q(\m_sys.m_bootloader.r_offset_1[2] ));
 sg13g2_dfrbp_1 _19221_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1034),
    .D(_01079_),
    .Q_N(_08249_),
    .Q(\m_sys.m_bootloader.r_offset_1[3] ));
 sg13g2_dfrbp_1 _19222_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1033),
    .D(_01080_),
    .Q_N(_08248_),
    .Q(\m_sys.m_bootloader.r_offset_1[4] ));
 sg13g2_dfrbp_1 _19223_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1032),
    .D(_01081_),
    .Q_N(_08247_),
    .Q(\m_sys.m_bootloader.r_offset_1[5] ));
 sg13g2_dfrbp_1 _19224_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1031),
    .D(_01082_),
    .Q_N(_08246_),
    .Q(\m_sys.m_bootloader.r_offset_1[6] ));
 sg13g2_dfrbp_1 _19225_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1030),
    .D(_01083_),
    .Q_N(_08245_),
    .Q(\m_sys.m_bootloader.r_offset_1[7] ));
 sg13g2_dfrbp_1 _19226_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1029),
    .D(_01084_),
    .Q_N(_00015_),
    .Q(\m_sys._m_bootloader_io_o_bl ));
 sg13g2_dfrbp_1 _19227_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1028),
    .D(_01085_),
    .Q_N(_00025_),
    .Q(\m_sys._m_bootloader_io_b_mem_wen[0] ));
 sg13g2_dfrbp_1 _19228_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1026),
    .D(net1868),
    .Q_N(_00064_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[0] ));
 sg13g2_dfrbp_1 _19229_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1025),
    .D(net3249),
    .Q_N(_00043_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[1] ));
 sg13g2_dfrbp_1 _19230_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1024),
    .D(_01088_),
    .Q_N(_08244_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[2] ));
 sg13g2_dfrbp_1 _19231_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1023),
    .D(net3102),
    .Q_N(_08243_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[3] ));
 sg13g2_dfrbp_1 _19232_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1022),
    .D(_01090_),
    .Q_N(_08242_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[4] ));
 sg13g2_dfrbp_1 _19233_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1021),
    .D(net3134),
    .Q_N(_00044_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[5] ));
 sg13g2_dfrbp_1 _19234_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1020),
    .D(net3038),
    .Q_N(_00045_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[6] ));
 sg13g2_dfrbp_1 _19235_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1019),
    .D(net3376),
    .Q_N(_08241_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[7] ));
 sg13g2_dfrbp_1 _19236_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1018),
    .D(_01094_),
    .Q_N(_08240_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[8] ));
 sg13g2_dfrbp_1 _19237_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1017),
    .D(_01095_),
    .Q_N(_08239_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[9] ));
 sg13g2_dfrbp_1 _19238_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1016),
    .D(net3355),
    .Q_N(_08238_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[10] ));
 sg13g2_dfrbp_1 _19239_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1015),
    .D(net3246),
    .Q_N(_08237_),
    .Q(\m_sys._m_bootloader_io_b_mem_addr[11] ));
 sg13g2_dfrbp_1 _19240_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1014),
    .D(_01098_),
    .Q_N(_00048_),
    .Q(\m_sys._m_ram_io_b_port_rdata[0] ));
 sg13g2_dfrbp_1 _19241_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1012),
    .D(_01099_),
    .Q_N(_00050_),
    .Q(\m_sys._m_ram_io_b_port_rdata[1] ));
 sg13g2_dfrbp_1 _19242_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1010),
    .D(_01100_),
    .Q_N(_00052_),
    .Q(\m_sys._m_ram_io_b_port_rdata[2] ));
 sg13g2_dfrbp_1 _19243_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1008),
    .D(_01101_),
    .Q_N(_00054_),
    .Q(\m_sys._m_ram_io_b_port_rdata[3] ));
 sg13g2_dfrbp_1 _19244_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1006),
    .D(_01102_),
    .Q_N(_00056_),
    .Q(\m_sys._m_ram_io_b_port_rdata[4] ));
 sg13g2_dfrbp_1 _19245_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1004),
    .D(_01103_),
    .Q_N(_00058_),
    .Q(\m_sys._m_ram_io_b_port_rdata[5] ));
 sg13g2_dfrbp_1 _19246_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1002),
    .D(_01104_),
    .Q_N(_00060_),
    .Q(\m_sys._m_ram_io_b_port_rdata[6] ));
 sg13g2_dfrbp_1 _19247_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1000),
    .D(_01105_),
    .Q_N(_00062_),
    .Q(\m_sys._m_ram_io_b_port_rdata[7] ));
 sg13g2_dfrbp_1 _19248_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net998),
    .D(_01106_),
    .Q_N(_00049_),
    .Q(\m_sys._m_ram_io_b_port_rdata[8] ));
 sg13g2_dfrbp_1 _19249_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net996),
    .D(_01107_),
    .Q_N(_00051_),
    .Q(\m_sys._m_ram_io_b_port_rdata[9] ));
 sg13g2_dfrbp_1 _19250_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net994),
    .D(_01108_),
    .Q_N(_00053_),
    .Q(\m_sys._m_ram_io_b_port_rdata[10] ));
 sg13g2_dfrbp_1 _19251_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net992),
    .D(_01109_),
    .Q_N(_00055_),
    .Q(\m_sys._m_ram_io_b_port_rdata[11] ));
 sg13g2_dfrbp_1 _19252_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net990),
    .D(_01110_),
    .Q_N(_00057_),
    .Q(\m_sys._m_ram_io_b_port_rdata[12] ));
 sg13g2_dfrbp_1 _19253_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net988),
    .D(_01111_),
    .Q_N(_00059_),
    .Q(\m_sys._m_ram_io_b_port_rdata[13] ));
 sg13g2_dfrbp_1 _19254_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net986),
    .D(_01112_),
    .Q_N(_00061_),
    .Q(\m_sys._m_ram_io_b_port_rdata[14] ));
 sg13g2_dfrbp_1 _19255_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net984),
    .D(_01113_),
    .Q_N(_00063_),
    .Q(\m_sys._m_ram_io_b_port_rdata[15] ));
 sg13g2_dfrbp_1 _19256_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net982),
    .D(_01114_),
    .Q_N(_08236_),
    .Q(\m_sys._m_ram_io_b_port_rdata[16] ));
 sg13g2_dfrbp_1 _19257_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net980),
    .D(_01115_),
    .Q_N(_08235_),
    .Q(\m_sys._m_ram_io_b_port_rdata[17] ));
 sg13g2_dfrbp_1 _19258_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net978),
    .D(_01116_),
    .Q_N(_08234_),
    .Q(\m_sys._m_ram_io_b_port_rdata[18] ));
 sg13g2_dfrbp_1 _19259_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net976),
    .D(_01117_),
    .Q_N(_08233_),
    .Q(\m_sys._m_ram_io_b_port_rdata[19] ));
 sg13g2_dfrbp_1 _19260_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net974),
    .D(_01118_),
    .Q_N(_00138_),
    .Q(\m_sys._m_ram_io_b_port_rdata[20] ));
 sg13g2_dfrbp_1 _19261_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net972),
    .D(_01119_),
    .Q_N(_00140_),
    .Q(\m_sys._m_ram_io_b_port_rdata[21] ));
 sg13g2_dfrbp_1 _19262_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net970),
    .D(_01120_),
    .Q_N(_00142_),
    .Q(\m_sys._m_ram_io_b_port_rdata[22] ));
 sg13g2_dfrbp_1 _19263_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net968),
    .D(_01121_),
    .Q_N(_00144_),
    .Q(\m_sys._m_ram_io_b_port_rdata[23] ));
 sg13g2_dfrbp_1 _19264_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net966),
    .D(_01122_),
    .Q_N(_08232_),
    .Q(\m_sys._m_ram_io_b_port_rdata[24] ));
 sg13g2_dfrbp_1 _19265_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net964),
    .D(_01123_),
    .Q_N(_08231_),
    .Q(\m_sys._m_ram_io_b_port_rdata[25] ));
 sg13g2_dfrbp_1 _19266_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net962),
    .D(_01124_),
    .Q_N(_08230_),
    .Q(\m_sys._m_ram_io_b_port_rdata[26] ));
 sg13g2_dfrbp_1 _19267_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net960),
    .D(_01125_),
    .Q_N(_08229_),
    .Q(\m_sys._m_ram_io_b_port_rdata[27] ));
 sg13g2_dfrbp_1 _19268_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net958),
    .D(_01126_),
    .Q_N(_08228_),
    .Q(\m_sys._m_ram_io_b_port_rdata[28] ));
 sg13g2_dfrbp_1 _19269_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net956),
    .D(_01127_),
    .Q_N(_08227_),
    .Q(\m_sys._m_ram_io_b_port_rdata[29] ));
 sg13g2_dfrbp_1 _19270_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net954),
    .D(_01128_),
    .Q_N(_08226_),
    .Q(\m_sys._m_ram_io_b_port_rdata[30] ));
 sg13g2_dfrbp_1 _19271_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net952),
    .D(_01129_),
    .Q_N(_08225_),
    .Q(\m_sys._m_ram_io_b_port_rdata[31] ));
 sg13g2_dfrbp_1 _19272_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net950),
    .D(_01130_),
    .Q_N(_08224_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][24] ));
 sg13g2_dfrbp_1 _19273_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net949),
    .D(_01131_),
    .Q_N(_08223_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][25] ));
 sg13g2_dfrbp_1 _19274_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net948),
    .D(_01132_),
    .Q_N(_08222_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][26] ));
 sg13g2_dfrbp_1 _19275_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net947),
    .D(_01133_),
    .Q_N(_08221_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][27] ));
 sg13g2_dfrbp_1 _19276_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net946),
    .D(_01134_),
    .Q_N(_08220_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][28] ));
 sg13g2_dfrbp_1 _19277_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net945),
    .D(_01135_),
    .Q_N(_08219_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][29] ));
 sg13g2_dfrbp_1 _19278_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net944),
    .D(_01136_),
    .Q_N(_08218_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][30] ));
 sg13g2_dfrbp_1 _19279_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net943),
    .D(_01137_),
    .Q_N(_08217_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][31] ));
 sg13g2_dfrbp_1 _19280_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net942),
    .D(_01138_),
    .Q_N(_08216_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[0] ));
 sg13g2_dfrbp_1 _19281_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net940),
    .D(_01139_),
    .Q_N(_08215_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[1] ));
 sg13g2_dfrbp_1 _19282_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net938),
    .D(_01140_),
    .Q_N(_08214_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[2] ));
 sg13g2_dfrbp_1 _19283_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net936),
    .D(_01141_),
    .Q_N(_08213_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[3] ));
 sg13g2_dfrbp_1 _19284_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net934),
    .D(_01142_),
    .Q_N(_08212_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[4] ));
 sg13g2_dfrbp_1 _19285_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net932),
    .D(_01143_),
    .Q_N(_08211_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[5] ));
 sg13g2_dfrbp_1 _19286_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net930),
    .D(_01144_),
    .Q_N(_08210_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[6] ));
 sg13g2_dfrbp_1 _19287_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net928),
    .D(_01145_),
    .Q_N(_08209_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[7] ));
 sg13g2_dfrbp_1 _19288_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net926),
    .D(_01146_),
    .Q_N(_08208_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[8] ));
 sg13g2_dfrbp_1 _19289_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net924),
    .D(_01147_),
    .Q_N(_08207_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[9] ));
 sg13g2_dfrbp_1 _19290_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net922),
    .D(_01148_),
    .Q_N(_08206_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[10] ));
 sg13g2_dfrbp_1 _19291_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net920),
    .D(_01149_),
    .Q_N(_08205_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[11] ));
 sg13g2_dfrbp_1 _19292_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net918),
    .D(_01150_),
    .Q_N(_08204_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[12] ));
 sg13g2_dfrbp_1 _19293_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net916),
    .D(_01151_),
    .Q_N(_08203_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[13] ));
 sg13g2_dfrbp_1 _19294_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net914),
    .D(_01152_),
    .Q_N(_08202_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[14] ));
 sg13g2_dfrbp_1 _19295_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net912),
    .D(_01153_),
    .Q_N(_08201_),
    .Q(\m_sys.m_uart.m_rx.io_i_ncycle[15] ));
 sg13g2_dfrbp_1 _19296_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net910),
    .D(_01154_),
    .Q_N(_08200_),
    .Q(\m_sys.m_gpio8.r_in[0] ));
 sg13g2_dfrbp_1 _19297_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net909),
    .D(_01155_),
    .Q_N(_08199_),
    .Q(\m_sys.m_gpio8.r_in[1] ));
 sg13g2_dfrbp_1 _19298_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net908),
    .D(_01156_),
    .Q_N(_08198_),
    .Q(\m_sys.m_gpio8.r_in[2] ));
 sg13g2_dfrbp_1 _19299_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net907),
    .D(_01157_),
    .Q_N(_08197_),
    .Q(\m_sys.m_gpio8.r_in[3] ));
 sg13g2_dfrbp_1 _19300_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net906),
    .D(_01158_),
    .Q_N(_08196_),
    .Q(\m_sys.m_gpio8.r_in[4] ));
 sg13g2_dfrbp_1 _19301_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net905),
    .D(_01159_),
    .Q_N(_08195_),
    .Q(\m_sys.m_gpio8.r_in[5] ));
 sg13g2_dfrbp_1 _19302_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net904),
    .D(_01160_),
    .Q_N(_08194_),
    .Q(\m_sys.m_gpio8.r_in[6] ));
 sg13g2_dfrbp_1 _19303_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net903),
    .D(_01161_),
    .Q_N(_08193_),
    .Q(\m_sys.m_gpio8.r_in[7] ));
 sg13g2_dfrbp_1 _19304_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net902),
    .D(_01162_),
    .Q_N(_08192_),
    .Q(\m_sys.m_uart.r_rx_valid ));
 sg13g2_dfrbp_1 _19305_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net901),
    .D(_01163_),
    .Q_N(_08191_),
    .Q(\m_sys.m_uart.m_rx.r_bit_cnt[0] ));
 sg13g2_dfrbp_1 _19306_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net899),
    .D(_01164_),
    .Q_N(_08190_),
    .Q(\m_sys.m_uart.m_rx.r_bit_cnt[1] ));
 sg13g2_dfrbp_1 _19307_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net897),
    .D(net2829),
    .Q_N(_08189_),
    .Q(\m_sys.m_uart.m_rx.r_bit_cnt[2] ));
 sg13g2_dfrbp_1 _19308_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net895),
    .D(_01166_),
    .Q_N(_08188_),
    .Q(\m_sys._m_uart_io_o_bl_data[0] ));
 sg13g2_dfrbp_1 _19309_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net893),
    .D(_01167_),
    .Q_N(_08187_),
    .Q(\m_sys._m_uart_io_o_bl_data[1] ));
 sg13g2_dfrbp_1 _19310_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net891),
    .D(_01168_),
    .Q_N(_08186_),
    .Q(\m_sys._m_uart_io_o_bl_data[2] ));
 sg13g2_dfrbp_1 _19311_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net889),
    .D(_01169_),
    .Q_N(_08185_),
    .Q(\m_sys._m_uart_io_o_bl_data[3] ));
 sg13g2_dfrbp_1 _19312_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net887),
    .D(net3004),
    .Q_N(_08184_),
    .Q(\m_sys._m_uart_io_o_bl_data[4] ));
 sg13g2_dfrbp_1 _19313_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net885),
    .D(net2904),
    .Q_N(_08183_),
    .Q(\m_sys._m_uart_io_o_bl_data[5] ));
 sg13g2_dfrbp_1 _19314_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net883),
    .D(_01172_),
    .Q_N(_08182_),
    .Q(\m_sys._m_uart_io_o_bl_data[6] ));
 sg13g2_dfrbp_1 _19315_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net881),
    .D(_01173_),
    .Q_N(_08181_),
    .Q(\m_sys._m_uart_io_o_bl_data[7] ));
 sg13g2_dfrbp_1 _19316_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net879),
    .D(net2863),
    .Q_N(_08180_),
    .Q(\m_sys.m_uart.r_rx_data[0] ));
 sg13g2_dfrbp_1 _19317_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net878),
    .D(_01175_),
    .Q_N(_08179_),
    .Q(\m_sys.m_uart.r_rx_data[1] ));
 sg13g2_dfrbp_1 _19318_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net877),
    .D(_01176_),
    .Q_N(_08178_),
    .Q(\m_sys.m_uart.r_rx_data[2] ));
 sg13g2_dfrbp_1 _19319_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net876),
    .D(_01177_),
    .Q_N(_08177_),
    .Q(\m_sys.m_uart.r_rx_data[3] ));
 sg13g2_dfrbp_1 _19320_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net875),
    .D(net2446),
    .Q_N(_08176_),
    .Q(\m_sys.m_uart.r_rx_data[4] ));
 sg13g2_dfrbp_1 _19321_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net874),
    .D(_01179_),
    .Q_N(_08175_),
    .Q(\m_sys.m_uart.r_rx_data[5] ));
 sg13g2_dfrbp_1 _19322_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net873),
    .D(_01180_),
    .Q_N(_08174_),
    .Q(\m_sys.m_uart.r_rx_data[6] ));
 sg13g2_dfrbp_1 _19323_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net872),
    .D(_01181_),
    .Q_N(_08173_),
    .Q(\m_sys.m_uart.r_rx_data[7] ));
 sg13g2_dfrbp_1 _19324_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net871),
    .D(net3139),
    .Q_N(_08172_),
    .Q(\m_sys.r_addr[6] ));
 sg13g2_dfrbp_1 _19325_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net870),
    .D(net3115),
    .Q_N(_08171_),
    .Q(\m_sys.r_addr[7] ));
 sg13g2_dfrbp_1 _19326_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net869),
    .D(net3143),
    .Q_N(_08170_),
    .Q(\m_sys.r_addr[8] ));
 sg13g2_dfrbp_1 _19327_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net868),
    .D(net3165),
    .Q_N(_08169_),
    .Q(\m_sys.r_addr[9] ));
 sg13g2_dfrbp_1 _19328_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net867),
    .D(net3235),
    .Q_N(_08168_),
    .Q(\m_sys.r_addr[10] ));
 sg13g2_dfrbp_1 _19329_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net866),
    .D(net3352),
    .Q_N(_08167_),
    .Q(\m_sys.r_addr[11] ));
 sg13g2_dfrbp_1 _19330_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net865),
    .D(_01188_),
    .Q_N(_08166_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][24] ));
 sg13g2_dfrbp_1 _19331_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net864),
    .D(_01189_),
    .Q_N(_08165_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][25] ));
 sg13g2_dfrbp_1 _19332_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net863),
    .D(_01190_),
    .Q_N(_08164_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][26] ));
 sg13g2_dfrbp_1 _19333_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net862),
    .D(_01191_),
    .Q_N(_08163_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][27] ));
 sg13g2_dfrbp_1 _19334_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net861),
    .D(_01192_),
    .Q_N(_08162_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][28] ));
 sg13g2_dfrbp_1 _19335_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net860),
    .D(_01193_),
    .Q_N(_08161_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][29] ));
 sg13g2_dfrbp_1 _19336_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net859),
    .D(_01194_),
    .Q_N(_08160_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][30] ));
 sg13g2_dfrbp_1 _19337_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1067),
    .D(_01195_),
    .Q_N(_09108_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][31] ));
 sg13g2_dfrbp_1 _19338_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1068),
    .D(net3237),
    .Q_N(_09109_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[0] ));
 sg13g2_dfrbp_1 _19339_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1069),
    .D(_01751_),
    .Q_N(_09110_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[1] ));
 sg13g2_dfrbp_1 _19340_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1070),
    .D(_01752_),
    .Q_N(_09111_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[2] ));
 sg13g2_dfrbp_1 _19341_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1071),
    .D(_01753_),
    .Q_N(_09112_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[3] ));
 sg13g2_dfrbp_1 _19342_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1072),
    .D(_01754_),
    .Q_N(_09113_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[4] ));
 sg13g2_dfrbp_1 _19343_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1073),
    .D(_01755_),
    .Q_N(_09114_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[5] ));
 sg13g2_dfrbp_1 _19344_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1074),
    .D(_01756_),
    .Q_N(_09115_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[6] ));
 sg13g2_dfrbp_1 _19345_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1075),
    .D(_01757_),
    .Q_N(_09116_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[7] ));
 sg13g2_dfrbp_1 _19346_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1076),
    .D(_01758_),
    .Q_N(_09117_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[8] ));
 sg13g2_dfrbp_1 _19347_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1077),
    .D(_01759_),
    .Q_N(_09118_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[9] ));
 sg13g2_dfrbp_1 _19348_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1078),
    .D(_01745_),
    .Q_N(_09119_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[10] ));
 sg13g2_dfrbp_1 _19349_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1079),
    .D(_01746_),
    .Q_N(_09120_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[11] ));
 sg13g2_dfrbp_1 _19350_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1080),
    .D(_01747_),
    .Q_N(_09121_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[12] ));
 sg13g2_dfrbp_1 _19351_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1081),
    .D(_01748_),
    .Q_N(_09122_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[13] ));
 sg13g2_dfrbp_1 _19352_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1110),
    .D(_01749_),
    .Q_N(_09123_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[14] ));
 sg13g2_dfrbp_1 _19353_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net858),
    .D(_01750_),
    .Q_N(_08159_),
    .Q(\m_sys.m_uart.m_rx.r_cycle_cnt[15] ));
 sg13g2_dfrbp_1 _19354_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net857),
    .D(net2534),
    .Q_N(_00122_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[0] ));
 sg13g2_dfrbp_1 _19355_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net856),
    .D(_01197_),
    .Q_N(_00124_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[1] ));
 sg13g2_dfrbp_1 _19356_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net855),
    .D(_01198_),
    .Q_N(_00126_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[2] ));
 sg13g2_dfrbp_1 _19357_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net854),
    .D(_01199_),
    .Q_N(_00128_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[3] ));
 sg13g2_dfrbp_1 _19358_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net853),
    .D(_01200_),
    .Q_N(_00130_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[4] ));
 sg13g2_dfrbp_1 _19359_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net852),
    .D(_01201_),
    .Q_N(_00132_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[5] ));
 sg13g2_dfrbp_1 _19360_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net851),
    .D(_01202_),
    .Q_N(_00134_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[6] ));
 sg13g2_dfrbp_1 _19361_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net850),
    .D(_01203_),
    .Q_N(_00136_),
    .Q(\m_sys._m_uart_io_b_mem_rdata[7] ));
 sg13g2_dfrbp_1 _19362_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net849),
    .D(_01204_),
    .Q_N(_08158_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][0] ));
 sg13g2_dfrbp_1 _19363_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net848),
    .D(_01205_),
    .Q_N(_08157_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][1] ));
 sg13g2_dfrbp_1 _19364_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net847),
    .D(_01206_),
    .Q_N(_08156_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][2] ));
 sg13g2_dfrbp_1 _19365_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net846),
    .D(_01207_),
    .Q_N(_08155_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][3] ));
 sg13g2_dfrbp_1 _19366_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net845),
    .D(_01208_),
    .Q_N(_08154_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][4] ));
 sg13g2_dfrbp_1 _19367_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net844),
    .D(_01209_),
    .Q_N(_08153_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][5] ));
 sg13g2_dfrbp_1 _19368_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net843),
    .D(_01210_),
    .Q_N(_08152_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][6] ));
 sg13g2_dfrbp_1 _19369_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net842),
    .D(_01211_),
    .Q_N(_08151_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][7] ));
 sg13g2_dfrbp_1 _19370_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net841),
    .D(_01212_),
    .Q_N(_08150_),
    .Q(\m_sys.m_uart.m_tx.r_bit_cnt[0] ));
 sg13g2_dfrbp_1 _19371_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net839),
    .D(_01213_),
    .Q_N(_08149_),
    .Q(\m_sys.m_uart.m_tx.r_bit_cnt[1] ));
 sg13g2_dfrbp_1 _19372_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net837),
    .D(_01214_),
    .Q_N(_08148_),
    .Q(\m_sys.m_uart.m_tx.r_bit_cnt[2] ));
 sg13g2_dfrbp_1 _19373_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net835),
    .D(_01215_),
    .Q_N(_08147_),
    .Q(\m_sys.m_uart.m_rx.r_rx ));
 sg13g2_dfrbp_1 _19374_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net834),
    .D(_01216_),
    .Q_N(_08146_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][24] ));
 sg13g2_dfrbp_1 _19375_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net833),
    .D(_01217_),
    .Q_N(_08145_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][25] ));
 sg13g2_dfrbp_1 _19376_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net832),
    .D(_01218_),
    .Q_N(_08144_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][26] ));
 sg13g2_dfrbp_1 _19377_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net831),
    .D(_01219_),
    .Q_N(_08143_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][27] ));
 sg13g2_dfrbp_1 _19378_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net830),
    .D(_01220_),
    .Q_N(_08142_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][28] ));
 sg13g2_dfrbp_1 _19379_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net829),
    .D(_01221_),
    .Q_N(_08141_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][29] ));
 sg13g2_dfrbp_1 _19380_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net828),
    .D(_01222_),
    .Q_N(_08140_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][30] ));
 sg13g2_dfrbp_1 _19381_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1111),
    .D(_01223_),
    .Q_N(_09124_),
    .Q(\m_sys.m_ram.m_ram.r_mem[28][31] ));
 sg13g2_dfrbp_1 _19382_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1112),
    .D(_01760_),
    .Q_N(_09125_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[0] ));
 sg13g2_dfrbp_1 _19383_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1113),
    .D(_01767_),
    .Q_N(_09126_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[1] ));
 sg13g2_dfrbp_1 _19384_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1114),
    .D(net2913),
    .Q_N(_09127_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[2] ));
 sg13g2_dfrbp_1 _19385_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1115),
    .D(_01769_),
    .Q_N(_09128_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[3] ));
 sg13g2_dfrbp_1 _19386_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1116),
    .D(_01770_),
    .Q_N(_09129_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[4] ));
 sg13g2_dfrbp_1 _19387_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1117),
    .D(_01771_),
    .Q_N(_09130_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[5] ));
 sg13g2_dfrbp_1 _19388_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1118),
    .D(net3100),
    .Q_N(_09131_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[6] ));
 sg13g2_dfrbp_1 _19389_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1119),
    .D(_01773_),
    .Q_N(_09132_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[7] ));
 sg13g2_dfrbp_1 _19390_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1120),
    .D(_01774_),
    .Q_N(_09133_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[8] ));
 sg13g2_dfrbp_1 _19391_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1121),
    .D(_01775_),
    .Q_N(_09134_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[9] ));
 sg13g2_dfrbp_1 _19392_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1122),
    .D(net3033),
    .Q_N(_09135_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[10] ));
 sg13g2_dfrbp_1 _19393_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1123),
    .D(_01762_),
    .Q_N(_09136_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[11] ));
 sg13g2_dfrbp_1 _19394_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1124),
    .D(net2938),
    .Q_N(_09137_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[12] ));
 sg13g2_dfrbp_1 _19395_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1125),
    .D(_01764_),
    .Q_N(_09138_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[13] ));
 sg13g2_dfrbp_1 _19396_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1134),
    .D(_01765_),
    .Q_N(_09139_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[14] ));
 sg13g2_dfrbp_1 _19397_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net827),
    .D(_01766_),
    .Q_N(_08139_),
    .Q(\m_sys.m_uart.m_tx.r_cycle_cnt[15] ));
 sg13g2_dfrbp_1 _19398_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net826),
    .D(_01224_),
    .Q_N(_08138_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][8] ));
 sg13g2_dfrbp_1 _19399_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net825),
    .D(_01225_),
    .Q_N(_08137_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][9] ));
 sg13g2_dfrbp_1 _19400_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net824),
    .D(_01226_),
    .Q_N(_08136_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][10] ));
 sg13g2_dfrbp_1 _19401_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net823),
    .D(_01227_),
    .Q_N(_08135_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][11] ));
 sg13g2_dfrbp_1 _19402_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net822),
    .D(_01228_),
    .Q_N(_08134_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][12] ));
 sg13g2_dfrbp_1 _19403_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net821),
    .D(_01229_),
    .Q_N(_08133_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][13] ));
 sg13g2_dfrbp_1 _19404_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net820),
    .D(_01230_),
    .Q_N(_08132_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][14] ));
 sg13g2_dfrbp_1 _19405_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1135),
    .D(_01231_),
    .Q_N(_09140_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][15] ));
 sg13g2_dfrbp_1 _19406_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1136),
    .D(net3295),
    .Q_N(_00121_),
    .Q(\m_sys._m_gpio8_io_b_mem_rdata[0] ));
 sg13g2_dfrbp_1 _19407_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1137),
    .D(net3229),
    .Q_N(_00123_),
    .Q(\m_sys._m_gpio8_io_b_mem_rdata[1] ));
 sg13g2_dfrbp_1 _19408_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1138),
    .D(net3256),
    .Q_N(_00125_),
    .Q(\m_sys._m_gpio8_io_b_mem_rdata[2] ));
 sg13g2_dfrbp_1 _19409_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1139),
    .D(net3219),
    .Q_N(_00127_),
    .Q(\m_sys._m_gpio8_io_b_mem_rdata[3] ));
 sg13g2_dfrbp_1 _19410_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1140),
    .D(net3285),
    .Q_N(_00129_),
    .Q(\m_sys._m_gpio8_io_b_mem_rdata[4] ));
 sg13g2_dfrbp_1 _19411_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1141),
    .D(net3200),
    .Q_N(_00131_),
    .Q(\m_sys._m_gpio8_io_b_mem_rdata[5] ));
 sg13g2_dfrbp_1 _19412_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net645),
    .D(net3283),
    .Q_N(_00133_),
    .Q(\m_sys._m_gpio8_io_b_mem_rdata[6] ));
 sg13g2_dfrbp_1 _19413_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net819),
    .D(net3346),
    .Q_N(_00135_),
    .Q(\m_sys._m_gpio8_io_b_mem_rdata[7] ));
 sg13g2_dfrbp_1 _19414_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net818),
    .D(_01232_),
    .Q_N(_08131_),
    .Q(uio_oe[0]));
 sg13g2_dfrbp_1 _19415_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net816),
    .D(_01233_),
    .Q_N(_08130_),
    .Q(uio_oe[1]));
 sg13g2_dfrbp_1 _19416_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net814),
    .D(_01234_),
    .Q_N(_08129_),
    .Q(uio_oe[2]));
 sg13g2_dfrbp_1 _19417_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net812),
    .D(_01235_),
    .Q_N(_08128_),
    .Q(uio_oe[3]));
 sg13g2_dfrbp_1 _19418_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net810),
    .D(_01236_),
    .Q_N(_08127_),
    .Q(uio_oe[4]));
 sg13g2_dfrbp_1 _19419_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net808),
    .D(_01237_),
    .Q_N(_08126_),
    .Q(uio_oe[5]));
 sg13g2_dfrbp_1 _19420_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net806),
    .D(_01238_),
    .Q_N(_08125_),
    .Q(uio_oe[6]));
 sg13g2_dfrbp_1 _19421_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net804),
    .D(_01239_),
    .Q_N(_08124_),
    .Q(uio_oe[7]));
 sg13g2_dfrbp_1 _19422_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net802),
    .D(net2974),
    .Q_N(_08123_),
    .Q(\m_sys.m_core.m_gpr._GEN[224] ));
 sg13g2_dfrbp_1 _19423_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net801),
    .D(net3105),
    .Q_N(_08122_),
    .Q(\m_sys.m_core.m_gpr._GEN[225] ));
 sg13g2_dfrbp_1 _19424_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net800),
    .D(net3064),
    .Q_N(_08121_),
    .Q(\m_sys.m_core.m_gpr._GEN[226] ));
 sg13g2_dfrbp_1 _19425_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net799),
    .D(_01243_),
    .Q_N(_08120_),
    .Q(\m_sys.m_core.m_gpr._GEN[227] ));
 sg13g2_dfrbp_1 _19426_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net798),
    .D(net3111),
    .Q_N(_08119_),
    .Q(\m_sys.m_core.m_gpr._GEN[228] ));
 sg13g2_dfrbp_1 _19427_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net797),
    .D(_01245_),
    .Q_N(_08118_),
    .Q(\m_sys.m_core.m_gpr._GEN[229] ));
 sg13g2_dfrbp_1 _19428_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net796),
    .D(net2888),
    .Q_N(_08117_),
    .Q(\m_sys.m_core.m_gpr._GEN[230] ));
 sg13g2_dfrbp_1 _19429_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net795),
    .D(net2809),
    .Q_N(_08116_),
    .Q(\m_sys.m_core.m_gpr._GEN[231] ));
 sg13g2_dfrbp_1 _19430_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net794),
    .D(_01248_),
    .Q_N(_08115_),
    .Q(\m_sys.m_core.m_gpr._GEN[232] ));
 sg13g2_dfrbp_1 _19431_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net793),
    .D(net2997),
    .Q_N(_08114_),
    .Q(\m_sys.m_core.m_gpr._GEN[233] ));
 sg13g2_dfrbp_1 _19432_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net792),
    .D(net3078),
    .Q_N(_08113_),
    .Q(\m_sys.m_core.m_gpr._GEN[234] ));
 sg13g2_dfrbp_1 _19433_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net791),
    .D(net2957),
    .Q_N(_08112_),
    .Q(\m_sys.m_core.m_gpr._GEN[235] ));
 sg13g2_dfrbp_1 _19434_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net790),
    .D(net2836),
    .Q_N(_08111_),
    .Q(\m_sys.m_core.m_gpr._GEN[236] ));
 sg13g2_dfrbp_1 _19435_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net789),
    .D(_01253_),
    .Q_N(_08110_),
    .Q(\m_sys.m_core.m_gpr._GEN[237] ));
 sg13g2_dfrbp_1 _19436_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net788),
    .D(net2980),
    .Q_N(_08109_),
    .Q(\m_sys.m_core.m_gpr._GEN[238] ));
 sg13g2_dfrbp_1 _19437_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net787),
    .D(net2848),
    .Q_N(_08108_),
    .Q(\m_sys.m_core.m_gpr._GEN[239] ));
 sg13g2_dfrbp_1 _19438_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net786),
    .D(_01256_),
    .Q_N(_08107_),
    .Q(\m_sys.m_core.m_gpr._GEN[240] ));
 sg13g2_dfrbp_1 _19439_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net785),
    .D(_01257_),
    .Q_N(_08106_),
    .Q(\m_sys.m_core.m_gpr._GEN[241] ));
 sg13g2_dfrbp_1 _19440_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net784),
    .D(net2959),
    .Q_N(_08105_),
    .Q(\m_sys.m_core.m_gpr._GEN[242] ));
 sg13g2_dfrbp_1 _19441_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net783),
    .D(net3055),
    .Q_N(_08104_),
    .Q(\m_sys.m_core.m_gpr._GEN[243] ));
 sg13g2_dfrbp_1 _19442_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net782),
    .D(_01260_),
    .Q_N(_08103_),
    .Q(\m_sys.m_core.m_gpr._GEN[244] ));
 sg13g2_dfrbp_1 _19443_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net781),
    .D(_01261_),
    .Q_N(_08102_),
    .Q(\m_sys.m_core.m_gpr._GEN[245] ));
 sg13g2_dfrbp_1 _19444_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net780),
    .D(_01262_),
    .Q_N(_08101_),
    .Q(\m_sys.m_core.m_gpr._GEN[246] ));
 sg13g2_dfrbp_1 _19445_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net779),
    .D(net2893),
    .Q_N(_08100_),
    .Q(\m_sys.m_core.m_gpr._GEN[247] ));
 sg13g2_dfrbp_1 _19446_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net778),
    .D(net2966),
    .Q_N(_08099_),
    .Q(\m_sys.m_core.m_gpr._GEN[248] ));
 sg13g2_dfrbp_1 _19447_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net777),
    .D(net2984),
    .Q_N(_08098_),
    .Q(\m_sys.m_core.m_gpr._GEN[249] ));
 sg13g2_dfrbp_1 _19448_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net776),
    .D(net2999),
    .Q_N(_08097_),
    .Q(\m_sys.m_core.m_gpr._GEN[250] ));
 sg13g2_dfrbp_1 _19449_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net775),
    .D(net2926),
    .Q_N(_08096_),
    .Q(\m_sys.m_core.m_gpr._GEN[251] ));
 sg13g2_dfrbp_1 _19450_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net774),
    .D(net2824),
    .Q_N(_08095_),
    .Q(\m_sys.m_core.m_gpr._GEN[252] ));
 sg13g2_dfrbp_1 _19451_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net773),
    .D(net2935),
    .Q_N(_08094_),
    .Q(\m_sys.m_core.m_gpr._GEN[253] ));
 sg13g2_dfrbp_1 _19452_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net772),
    .D(net3007),
    .Q_N(_08093_),
    .Q(\m_sys.m_core.m_gpr._GEN[254] ));
 sg13g2_dfrbp_1 _19453_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net771),
    .D(net2940),
    .Q_N(_08092_),
    .Q(\m_sys.m_core.m_gpr._GEN[255] ));
 sg13g2_dfrbp_1 _19454_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net770),
    .D(_01272_),
    .Q_N(_08091_),
    .Q(uio_out[0]));
 sg13g2_dfrbp_1 _19455_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net768),
    .D(_01273_),
    .Q_N(_08090_),
    .Q(uio_out[1]));
 sg13g2_dfrbp_1 _19456_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net766),
    .D(_01274_),
    .Q_N(_08089_),
    .Q(uio_out[2]));
 sg13g2_dfrbp_1 _19457_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net764),
    .D(net3392),
    .Q_N(_08088_),
    .Q(uio_out[3]));
 sg13g2_dfrbp_1 _19458_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net762),
    .D(_01276_),
    .Q_N(_08087_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _19459_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net760),
    .D(_01277_),
    .Q_N(_08086_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _19460_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net758),
    .D(_01278_),
    .Q_N(_08085_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _19461_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net756),
    .D(_01279_),
    .Q_N(_08084_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _19462_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net754),
    .D(_01280_),
    .Q_N(_08083_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][8] ));
 sg13g2_dfrbp_1 _19463_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net753),
    .D(_01281_),
    .Q_N(_08082_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][9] ));
 sg13g2_dfrbp_1 _19464_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net752),
    .D(_01282_),
    .Q_N(_08081_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][10] ));
 sg13g2_dfrbp_1 _19465_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net751),
    .D(_01283_),
    .Q_N(_08080_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][11] ));
 sg13g2_dfrbp_1 _19466_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net750),
    .D(_01284_),
    .Q_N(_08079_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][12] ));
 sg13g2_dfrbp_1 _19467_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net749),
    .D(_01285_),
    .Q_N(_08078_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][13] ));
 sg13g2_dfrbp_1 _19468_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net748),
    .D(_01286_),
    .Q_N(_08077_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][14] ));
 sg13g2_dfrbp_1 _19469_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net747),
    .D(_01287_),
    .Q_N(_08076_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][15] ));
 sg13g2_dfrbp_1 _19470_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net746),
    .D(_01288_),
    .Q_N(_08075_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][16] ));
 sg13g2_dfrbp_1 _19471_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net745),
    .D(_01289_),
    .Q_N(_08074_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][17] ));
 sg13g2_dfrbp_1 _19472_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net744),
    .D(_01290_),
    .Q_N(_08073_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][18] ));
 sg13g2_dfrbp_1 _19473_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net743),
    .D(_01291_),
    .Q_N(_08072_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][19] ));
 sg13g2_dfrbp_1 _19474_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net742),
    .D(_01292_),
    .Q_N(_08071_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][20] ));
 sg13g2_dfrbp_1 _19475_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net741),
    .D(_01293_),
    .Q_N(_08070_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][21] ));
 sg13g2_dfrbp_1 _19476_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net740),
    .D(_01294_),
    .Q_N(_08069_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][22] ));
 sg13g2_dfrbp_1 _19477_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net739),
    .D(_01295_),
    .Q_N(_08068_),
    .Q(\m_sys.m_ram.m_ram.r_mem[0][23] ));
 sg13g2_dfrbp_1 _19478_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net738),
    .D(_01296_),
    .Q_N(_08067_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][16] ));
 sg13g2_dfrbp_1 _19479_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net737),
    .D(_01297_),
    .Q_N(_08066_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][17] ));
 sg13g2_dfrbp_1 _19480_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net736),
    .D(_01298_),
    .Q_N(_08065_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][18] ));
 sg13g2_dfrbp_1 _19481_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net735),
    .D(_01299_),
    .Q_N(_08064_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][19] ));
 sg13g2_dfrbp_1 _19482_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net734),
    .D(_01300_),
    .Q_N(_08063_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][20] ));
 sg13g2_dfrbp_1 _19483_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net733),
    .D(_01301_),
    .Q_N(_08062_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][21] ));
 sg13g2_dfrbp_1 _19484_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net732),
    .D(_01302_),
    .Q_N(_08061_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][22] ));
 sg13g2_dfrbp_1 _19485_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net731),
    .D(_01303_),
    .Q_N(_08060_),
    .Q(\m_sys.m_ram.m_ram.r_mem[20][23] ));
 sg13g2_dfrbp_1 _19486_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net730),
    .D(_01304_),
    .Q_N(_08059_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][24] ));
 sg13g2_dfrbp_1 _19487_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net729),
    .D(_01305_),
    .Q_N(_08058_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][25] ));
 sg13g2_dfrbp_1 _19488_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net728),
    .D(_01306_),
    .Q_N(_08057_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][26] ));
 sg13g2_dfrbp_1 _19489_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net727),
    .D(_01307_),
    .Q_N(_08056_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][27] ));
 sg13g2_dfrbp_1 _19490_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net726),
    .D(_01308_),
    .Q_N(_08055_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][28] ));
 sg13g2_dfrbp_1 _19491_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net725),
    .D(_01309_),
    .Q_N(_08054_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][29] ));
 sg13g2_dfrbp_1 _19492_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net724),
    .D(_01310_),
    .Q_N(_08053_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][30] ));
 sg13g2_dfrbp_1 _19493_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net723),
    .D(_01311_),
    .Q_N(_08052_),
    .Q(\m_sys.m_ram.m_ram.r_mem[10][31] ));
 sg13g2_dfrbp_1 _19494_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net722),
    .D(_01312_),
    .Q_N(_08051_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[0] ));
 sg13g2_dfrbp_1 _19495_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net720),
    .D(_01313_),
    .Q_N(_08050_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[1] ));
 sg13g2_dfrbp_1 _19496_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net718),
    .D(_01314_),
    .Q_N(_00028_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[2] ));
 sg13g2_dfrbp_1 _19497_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net716),
    .D(_01315_),
    .Q_N(_00029_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[3] ));
 sg13g2_dfrbp_1 _19498_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net714),
    .D(_01316_),
    .Q_N(_00030_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[4] ));
 sg13g2_dfrbp_1 _19499_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net712),
    .D(net3113),
    .Q_N(_00031_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[5] ));
 sg13g2_dfrbp_1 _19500_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net710),
    .D(_01318_),
    .Q_N(_00032_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[6] ));
 sg13g2_dfrbp_1 _19501_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net708),
    .D(_01319_),
    .Q_N(_00034_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[7] ));
 sg13g2_dfrbp_1 _19502_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net706),
    .D(_01320_),
    .Q_N(_00035_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[8] ));
 sg13g2_dfrbp_1 _19503_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net704),
    .D(net3023),
    .Q_N(_00036_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[9] ));
 sg13g2_dfrbp_1 _19504_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net702),
    .D(net3062),
    .Q_N(_00037_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[10] ));
 sg13g2_dfrbp_1 _19505_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net700),
    .D(net3002),
    .Q_N(_00038_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[11] ));
 sg13g2_dfrbp_1 _19506_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net698),
    .D(net2922),
    .Q_N(_00039_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[12] ));
 sg13g2_dfrbp_1 _19507_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net696),
    .D(net2834),
    .Q_N(_00040_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[13] ));
 sg13g2_dfrbp_1 _19508_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net694),
    .D(net2452),
    .Q_N(_00041_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[14] ));
 sg13g2_dfrbp_1 _19509_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net692),
    .D(net2562),
    .Q_N(_00042_),
    .Q(\m_sys.m_bootloader.r_byte_cnt[15] ));
 sg13g2_dfrbp_1 _19510_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net690),
    .D(_01328_),
    .Q_N(_08049_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[0] ));
 sg13g2_dfrbp_1 _19511_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net689),
    .D(net3203),
    .Q_N(_08048_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[1] ));
 sg13g2_dfrbp_1 _19512_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net688),
    .D(_01330_),
    .Q_N(_00118_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[2] ));
 sg13g2_dfrbp_1 _19513_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net687),
    .D(_01331_),
    .Q_N(_08047_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[3] ));
 sg13g2_dfrbp_1 _19514_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net686),
    .D(_01332_),
    .Q_N(_08046_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[4] ));
 sg13g2_dfrbp_1 _19515_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net685),
    .D(_01333_),
    .Q_N(_00113_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[5] ));
 sg13g2_dfrbp_1 _19516_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net684),
    .D(_01334_),
    .Q_N(_00111_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[6] ));
 sg13g2_dfrbp_1 _19517_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net683),
    .D(_01335_),
    .Q_N(_00110_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[7] ));
 sg13g2_dfrbp_1 _19518_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net682),
    .D(_01336_),
    .Q_N(_00108_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[8] ));
 sg13g2_dfrbp_1 _19519_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net681),
    .D(_01337_),
    .Q_N(_00105_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[9] ));
 sg13g2_dfrbp_1 _19520_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net680),
    .D(_01338_),
    .Q_N(_00102_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[10] ));
 sg13g2_dfrbp_1 _19521_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net679),
    .D(_01339_),
    .Q_N(_00100_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[11] ));
 sg13g2_dfrbp_1 _19522_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net678),
    .D(_01340_),
    .Q_N(_08045_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[12] ));
 sg13g2_dfrbp_1 _19523_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net677),
    .D(_01341_),
    .Q_N(_08044_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[13] ));
 sg13g2_dfrbp_1 _19524_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net676),
    .D(net3406),
    .Q_N(_08043_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[14] ));
 sg13g2_dfrbp_1 _19525_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net675),
    .D(_01343_),
    .Q_N(_08042_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[15] ));
 sg13g2_dfrbp_1 _19526_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net674),
    .D(_01344_),
    .Q_N(_08041_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[16] ));
 sg13g2_dfrbp_1 _19527_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net673),
    .D(_01345_),
    .Q_N(_08040_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[17] ));
 sg13g2_dfrbp_1 _19528_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net672),
    .D(_01346_),
    .Q_N(_08039_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[18] ));
 sg13g2_dfrbp_1 _19529_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net671),
    .D(net3350),
    .Q_N(_08038_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[19] ));
 sg13g2_dfrbp_1 _19530_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net670),
    .D(_01348_),
    .Q_N(_08037_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[20] ));
 sg13g2_dfrbp_1 _19531_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net669),
    .D(_01349_),
    .Q_N(_08036_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[21] ));
 sg13g2_dfrbp_1 _19532_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net668),
    .D(_01350_),
    .Q_N(_08035_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[22] ));
 sg13g2_dfrbp_1 _19533_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net667),
    .D(_01351_),
    .Q_N(_08034_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[23] ));
 sg13g2_dfrbp_1 _19534_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net666),
    .D(_01352_),
    .Q_N(_08033_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[24] ));
 sg13g2_dfrbp_1 _19535_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net665),
    .D(_01353_),
    .Q_N(_08032_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[25] ));
 sg13g2_dfrbp_1 _19536_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net664),
    .D(_01354_),
    .Q_N(_08031_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[26] ));
 sg13g2_dfrbp_1 _19537_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net663),
    .D(_01355_),
    .Q_N(_08030_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[27] ));
 sg13g2_dfrbp_1 _19538_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net662),
    .D(_01356_),
    .Q_N(_08029_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[28] ));
 sg13g2_dfrbp_1 _19539_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net661),
    .D(_01357_),
    .Q_N(_08028_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[29] ));
 sg13g2_dfrbp_1 _19540_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net660),
    .D(_01358_),
    .Q_N(_08027_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[30] ));
 sg13g2_dfrbp_1 _19541_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net659),
    .D(_01359_),
    .Q_N(_08026_),
    .Q(\m_sys.m_core.m_bru.io_i_s2[31] ));
 sg13g2_dfrbp_1 _19542_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net658),
    .D(_01360_),
    .Q_N(_08025_),
    .Q(\m_sys.m_core.m_alu.io_i_uop[2] ));
 sg13g2_dfrbp_1 _19543_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net656),
    .D(net3224),
    .Q_N(_08024_),
    .Q(\m_sys.m_core._m_bru_io_o_res[0] ));
 sg13g2_dfrbp_1 _19544_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net654),
    .D(net3175),
    .Q_N(_08023_),
    .Q(\m_sys.m_core._m_bru_io_o_res[1] ));
 sg13g2_dfrbp_1 _19545_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net652),
    .D(_01363_),
    .Q_N(_08022_),
    .Q(\m_sys.m_core.m_bru.io_i_uop[2] ));
 sg13g2_dfrbp_1 _19546_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net650),
    .D(_01364_),
    .Q_N(_08021_),
    .Q(\m_sys.m_core.m_alu.io_i_signed ));
 sg13g2_dfrbp_1 _19547_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net649),
    .D(_01365_),
    .Q_N(_08020_),
    .Q(\m_sys.m_core.r_ctrl_bru_pc_rel ));
 sg13g2_dfrbp_1 _19548_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net648),
    .D(_01366_),
    .Q_N(_08019_),
    .Q(\m_sys.m_core.r_ctrl_mem_size[0] ));
 sg13g2_dfrbp_1 _19549_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net646),
    .D(net3177),
    .Q_N(_08018_),
    .Q(\m_sys.m_core.r_ctrl_mem_size[1] ));
 sg13g2_dfrbp_1 _19550_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net644),
    .D(_01368_),
    .Q_N(_08017_),
    .Q(\m_sys.m_core.r_ctrl_mem_rw ));
 sg13g2_dfrbp_1 _19551_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net643),
    .D(_01369_),
    .Q_N(_08016_),
    .Q(\m_sys.m_core.r_ctrl_mem_signed ));
 sg13g2_dfrbp_1 _19552_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net642),
    .D(_01370_),
    .Q_N(_08015_),
    .Q(\m_sys.m_core.r_ctrl_wb_en ));
 sg13g2_dfrbp_1 _19553_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net641),
    .D(net3186),
    .Q_N(_08014_),
    .Q(\m_sys.m_core.m_gpr.io_b_write_addr[0] ));
 sg13g2_dfrbp_1 _19554_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net640),
    .D(_01372_),
    .Q_N(_08013_),
    .Q(\m_sys.m_core.m_gpr.io_b_write_addr[1] ));
 sg13g2_dfrbp_1 _19555_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net639),
    .D(_01373_),
    .Q_N(_00145_),
    .Q(\m_sys.m_core.m_gpr.io_b_write_addr[2] ));
 sg13g2_dfrbp_1 _19556_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net638),
    .D(_01374_),
    .Q_N(_08012_),
    .Q(\m_sys.m_core.m_fsm.r_cstate[3] ));
 sg13g2_dfrbp_1 _19557_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net637),
    .D(_01375_),
    .Q_N(_08011_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][24] ));
 sg13g2_dfrbp_1 _19558_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net636),
    .D(_01376_),
    .Q_N(_08010_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][25] ));
 sg13g2_dfrbp_1 _19559_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net635),
    .D(_01377_),
    .Q_N(_08009_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][26] ));
 sg13g2_dfrbp_1 _19560_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net634),
    .D(_01378_),
    .Q_N(_08008_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][27] ));
 sg13g2_dfrbp_1 _19561_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net633),
    .D(_01379_),
    .Q_N(_08007_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][28] ));
 sg13g2_dfrbp_1 _19562_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net632),
    .D(_01380_),
    .Q_N(_08006_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][29] ));
 sg13g2_dfrbp_1 _19563_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net631),
    .D(_01381_),
    .Q_N(_08005_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][30] ));
 sg13g2_dfrbp_1 _19564_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net630),
    .D(_01382_),
    .Q_N(_08004_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][31] ));
 sg13g2_dfrbp_1 _19565_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net629),
    .D(_01383_),
    .Q_N(_08003_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][16] ));
 sg13g2_dfrbp_1 _19566_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net628),
    .D(_01384_),
    .Q_N(_08002_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][17] ));
 sg13g2_dfrbp_1 _19567_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net627),
    .D(_01385_),
    .Q_N(_08001_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][18] ));
 sg13g2_dfrbp_1 _19568_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net626),
    .D(_01386_),
    .Q_N(_08000_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][19] ));
 sg13g2_dfrbp_1 _19569_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net625),
    .D(_01387_),
    .Q_N(_07999_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][20] ));
 sg13g2_dfrbp_1 _19570_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net624),
    .D(_01388_),
    .Q_N(_07998_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][21] ));
 sg13g2_dfrbp_1 _19571_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net623),
    .D(_01389_),
    .Q_N(_07997_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][22] ));
 sg13g2_dfrbp_1 _19572_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net622),
    .D(_01390_),
    .Q_N(_07996_),
    .Q(\m_sys.m_ram.m_ram.r_mem[17][23] ));
 sg13g2_dfrbp_1 _19573_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net621),
    .D(_01391_),
    .Q_N(_07995_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][0] ));
 sg13g2_dfrbp_1 _19574_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net620),
    .D(_01392_),
    .Q_N(_07994_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][1] ));
 sg13g2_dfrbp_1 _19575_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net619),
    .D(_01393_),
    .Q_N(_07993_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][2] ));
 sg13g2_dfrbp_1 _19576_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net618),
    .D(_01394_),
    .Q_N(_07992_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][3] ));
 sg13g2_dfrbp_1 _19577_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net617),
    .D(_01395_),
    .Q_N(_07991_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][4] ));
 sg13g2_dfrbp_1 _19578_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net616),
    .D(_01396_),
    .Q_N(_07990_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][5] ));
 sg13g2_dfrbp_1 _19579_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net615),
    .D(_01397_),
    .Q_N(_07989_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][6] ));
 sg13g2_dfrbp_1 _19580_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net614),
    .D(_01398_),
    .Q_N(_07988_),
    .Q(\m_sys.m_ram.m_ram.r_mem[18][7] ));
 sg13g2_dfrbp_1 _19581_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net613),
    .D(_01399_),
    .Q_N(_07987_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][8] ));
 sg13g2_dfrbp_1 _19582_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net612),
    .D(_01400_),
    .Q_N(_07986_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][9] ));
 sg13g2_dfrbp_1 _19583_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net611),
    .D(_01401_),
    .Q_N(_07985_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][10] ));
 sg13g2_dfrbp_1 _19584_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net610),
    .D(_01402_),
    .Q_N(_07984_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][11] ));
 sg13g2_dfrbp_1 _19585_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net609),
    .D(_01403_),
    .Q_N(_07983_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][12] ));
 sg13g2_dfrbp_1 _19586_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net608),
    .D(_01404_),
    .Q_N(_07982_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][13] ));
 sg13g2_dfrbp_1 _19587_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net607),
    .D(_01405_),
    .Q_N(_07981_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][14] ));
 sg13g2_dfrbp_1 _19588_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net606),
    .D(_01406_),
    .Q_N(_07980_),
    .Q(\m_sys.m_ram.m_ram.r_mem[19][15] ));
 sg13g2_dfrbp_1 _19589_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net605),
    .D(_01407_),
    .Q_N(_07979_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][24] ));
 sg13g2_dfrbp_1 _19590_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net604),
    .D(_01408_),
    .Q_N(_07978_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][25] ));
 sg13g2_dfrbp_1 _19591_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net603),
    .D(_01409_),
    .Q_N(_07977_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][26] ));
 sg13g2_dfrbp_1 _19592_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net602),
    .D(_01410_),
    .Q_N(_07976_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][27] ));
 sg13g2_dfrbp_1 _19593_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net601),
    .D(_01411_),
    .Q_N(_07975_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][28] ));
 sg13g2_dfrbp_1 _19594_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net600),
    .D(_01412_),
    .Q_N(_07974_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][29] ));
 sg13g2_dfrbp_1 _19595_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net599),
    .D(_01413_),
    .Q_N(_07973_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][30] ));
 sg13g2_dfrbp_1 _19596_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net598),
    .D(_01414_),
    .Q_N(_07972_),
    .Q(\m_sys.m_ram.m_ram.r_mem[31][31] ));
 sg13g2_dfrbp_1 _19597_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net597),
    .D(_01415_),
    .Q_N(_07971_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][0] ));
 sg13g2_dfrbp_1 _19598_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net596),
    .D(_01416_),
    .Q_N(_07970_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][1] ));
 sg13g2_dfrbp_1 _19599_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net595),
    .D(_01417_),
    .Q_N(_07969_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][2] ));
 sg13g2_dfrbp_1 _19600_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net594),
    .D(_01418_),
    .Q_N(_07968_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][3] ));
 sg13g2_dfrbp_1 _19601_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net593),
    .D(_01419_),
    .Q_N(_07967_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][4] ));
 sg13g2_dfrbp_1 _19602_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net592),
    .D(_01420_),
    .Q_N(_07966_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][5] ));
 sg13g2_dfrbp_1 _19603_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net591),
    .D(_01421_),
    .Q_N(_07965_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][6] ));
 sg13g2_dfrbp_1 _19604_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net590),
    .D(_01422_),
    .Q_N(_07964_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][7] ));
 sg13g2_dfrbp_1 _19605_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net589),
    .D(_01423_),
    .Q_N(_07963_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][8] ));
 sg13g2_dfrbp_1 _19606_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net588),
    .D(_01424_),
    .Q_N(_07962_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][9] ));
 sg13g2_dfrbp_1 _19607_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net587),
    .D(_01425_),
    .Q_N(_07961_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][10] ));
 sg13g2_dfrbp_1 _19608_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net586),
    .D(_01426_),
    .Q_N(_07960_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][11] ));
 sg13g2_dfrbp_1 _19609_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net585),
    .D(_01427_),
    .Q_N(_07959_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][12] ));
 sg13g2_dfrbp_1 _19610_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net584),
    .D(_01428_),
    .Q_N(_07958_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][13] ));
 sg13g2_dfrbp_1 _19611_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net583),
    .D(_01429_),
    .Q_N(_07957_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][14] ));
 sg13g2_dfrbp_1 _19612_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net582),
    .D(_01430_),
    .Q_N(_07956_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][15] ));
 sg13g2_dfrbp_1 _19613_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net581),
    .D(_01431_),
    .Q_N(_07955_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][16] ));
 sg13g2_dfrbp_1 _19614_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net580),
    .D(_01432_),
    .Q_N(_07954_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][17] ));
 sg13g2_dfrbp_1 _19615_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net579),
    .D(_01433_),
    .Q_N(_07953_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][18] ));
 sg13g2_dfrbp_1 _19616_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net578),
    .D(_01434_),
    .Q_N(_07952_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][19] ));
 sg13g2_dfrbp_1 _19617_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net577),
    .D(_01435_),
    .Q_N(_07951_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][20] ));
 sg13g2_dfrbp_1 _19618_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net576),
    .D(_01436_),
    .Q_N(_07950_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][21] ));
 sg13g2_dfrbp_1 _19619_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net575),
    .D(_01437_),
    .Q_N(_07949_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][22] ));
 sg13g2_dfrbp_1 _19620_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net574),
    .D(_01438_),
    .Q_N(_07948_),
    .Q(\m_sys.m_ram.m_ram.r_mem[3][23] ));
 sg13g2_dfrbp_1 _19621_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net573),
    .D(_01439_),
    .Q_N(_07947_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][0] ));
 sg13g2_dfrbp_1 _19622_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net572),
    .D(_01440_),
    .Q_N(_07946_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][1] ));
 sg13g2_dfrbp_1 _19623_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net571),
    .D(_01441_),
    .Q_N(_07945_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][2] ));
 sg13g2_dfrbp_1 _19624_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net570),
    .D(_01442_),
    .Q_N(_07944_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][3] ));
 sg13g2_dfrbp_1 _19625_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net569),
    .D(_01443_),
    .Q_N(_07943_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][4] ));
 sg13g2_dfrbp_1 _19626_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net568),
    .D(_01444_),
    .Q_N(_07942_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][5] ));
 sg13g2_dfrbp_1 _19627_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net567),
    .D(_01445_),
    .Q_N(_07941_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][6] ));
 sg13g2_dfrbp_1 _19628_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net566),
    .D(_01446_),
    .Q_N(_07940_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][7] ));
 sg13g2_dfrbp_1 _19629_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net565),
    .D(_01447_),
    .Q_N(_07939_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][8] ));
 sg13g2_dfrbp_1 _19630_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net564),
    .D(_01448_),
    .Q_N(_07938_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][9] ));
 sg13g2_dfrbp_1 _19631_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net563),
    .D(_01449_),
    .Q_N(_07937_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][10] ));
 sg13g2_dfrbp_1 _19632_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net562),
    .D(_01450_),
    .Q_N(_07936_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][11] ));
 sg13g2_dfrbp_1 _19633_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net561),
    .D(_01451_),
    .Q_N(_07935_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][12] ));
 sg13g2_dfrbp_1 _19634_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net560),
    .D(_01452_),
    .Q_N(_07934_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][13] ));
 sg13g2_dfrbp_1 _19635_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net559),
    .D(_01453_),
    .Q_N(_07933_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][14] ));
 sg13g2_dfrbp_1 _19636_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net558),
    .D(_01454_),
    .Q_N(_07932_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][15] ));
 sg13g2_dfrbp_1 _19637_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net557),
    .D(_01455_),
    .Q_N(_07931_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][16] ));
 sg13g2_dfrbp_1 _19638_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net556),
    .D(_01456_),
    .Q_N(_07930_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][17] ));
 sg13g2_dfrbp_1 _19639_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net555),
    .D(_01457_),
    .Q_N(_07929_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][18] ));
 sg13g2_dfrbp_1 _19640_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net554),
    .D(_01458_),
    .Q_N(_07928_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][19] ));
 sg13g2_dfrbp_1 _19641_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net553),
    .D(_01459_),
    .Q_N(_07927_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][20] ));
 sg13g2_dfrbp_1 _19642_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net552),
    .D(_01460_),
    .Q_N(_07926_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][21] ));
 sg13g2_dfrbp_1 _19643_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net551),
    .D(_01461_),
    .Q_N(_07925_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][22] ));
 sg13g2_dfrbp_1 _19644_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net550),
    .D(_01462_),
    .Q_N(_07924_),
    .Q(\m_sys.m_ram.m_ram.r_mem[4][23] ));
 sg13g2_dfrbp_1 _19645_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net549),
    .D(_01463_),
    .Q_N(_07923_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][0] ));
 sg13g2_dfrbp_1 _19646_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net548),
    .D(_01464_),
    .Q_N(_07922_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][1] ));
 sg13g2_dfrbp_1 _19647_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net547),
    .D(_01465_),
    .Q_N(_07921_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][2] ));
 sg13g2_dfrbp_1 _19648_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net546),
    .D(_01466_),
    .Q_N(_07920_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][3] ));
 sg13g2_dfrbp_1 _19649_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net545),
    .D(_01467_),
    .Q_N(_07919_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][4] ));
 sg13g2_dfrbp_1 _19650_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net544),
    .D(_01468_),
    .Q_N(_07918_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][5] ));
 sg13g2_dfrbp_1 _19651_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net543),
    .D(_01469_),
    .Q_N(_07917_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][6] ));
 sg13g2_dfrbp_1 _19652_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net542),
    .D(_01470_),
    .Q_N(_07916_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][7] ));
 sg13g2_dfrbp_1 _19653_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net541),
    .D(net3118),
    .Q_N(_07915_),
    .Q(\m_sys.m_core.m_gpr._GEN[128] ));
 sg13g2_dfrbp_1 _19654_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net540),
    .D(net2989),
    .Q_N(_07914_),
    .Q(\m_sys.m_core.m_gpr._GEN[129] ));
 sg13g2_dfrbp_1 _19655_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net539),
    .D(net3051),
    .Q_N(_07913_),
    .Q(\m_sys.m_core.m_gpr._GEN[130] ));
 sg13g2_dfrbp_1 _19656_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net538),
    .D(_01474_),
    .Q_N(_07912_),
    .Q(\m_sys.m_core.m_gpr._GEN[131] ));
 sg13g2_dfrbp_1 _19657_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net537),
    .D(_01475_),
    .Q_N(_07911_),
    .Q(\m_sys.m_core.m_gpr._GEN[132] ));
 sg13g2_dfrbp_1 _19658_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net536),
    .D(net2982),
    .Q_N(_07910_),
    .Q(\m_sys.m_core.m_gpr._GEN[133] ));
 sg13g2_dfrbp_1 _19659_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net535),
    .D(_01477_),
    .Q_N(_07909_),
    .Q(\m_sys.m_core.m_gpr._GEN[134] ));
 sg13g2_dfrbp_1 _19660_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net534),
    .D(_01478_),
    .Q_N(_07908_),
    .Q(\m_sys.m_core.m_gpr._GEN[135] ));
 sg13g2_dfrbp_1 _19661_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net533),
    .D(_01479_),
    .Q_N(_07907_),
    .Q(\m_sys.m_core.m_gpr._GEN[136] ));
 sg13g2_dfrbp_1 _19662_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net532),
    .D(_01480_),
    .Q_N(_07906_),
    .Q(\m_sys.m_core.m_gpr._GEN[137] ));
 sg13g2_dfrbp_1 _19663_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net531),
    .D(net2954),
    .Q_N(_07905_),
    .Q(\m_sys.m_core.m_gpr._GEN[138] ));
 sg13g2_dfrbp_1 _19664_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net530),
    .D(net2945),
    .Q_N(_07904_),
    .Q(\m_sys.m_core.m_gpr._GEN[139] ));
 sg13g2_dfrbp_1 _19665_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net529),
    .D(_01483_),
    .Q_N(_07903_),
    .Q(\m_sys.m_core.m_gpr._GEN[140] ));
 sg13g2_dfrbp_1 _19666_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net528),
    .D(_01484_),
    .Q_N(_07902_),
    .Q(\m_sys.m_core.m_gpr._GEN[141] ));
 sg13g2_dfrbp_1 _19667_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net527),
    .D(net2977),
    .Q_N(_07901_),
    .Q(\m_sys.m_core.m_gpr._GEN[142] ));
 sg13g2_dfrbp_1 _19668_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net526),
    .D(_01486_),
    .Q_N(_07900_),
    .Q(\m_sys.m_core.m_gpr._GEN[143] ));
 sg13g2_dfrbp_1 _19669_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net525),
    .D(_01487_),
    .Q_N(_07899_),
    .Q(\m_sys.m_core.m_gpr._GEN[144] ));
 sg13g2_dfrbp_1 _19670_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net524),
    .D(_01488_),
    .Q_N(_07898_),
    .Q(\m_sys.m_core.m_gpr._GEN[145] ));
 sg13g2_dfrbp_1 _19671_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net523),
    .D(net2961),
    .Q_N(_07897_),
    .Q(\m_sys.m_core.m_gpr._GEN[146] ));
 sg13g2_dfrbp_1 _19672_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net522),
    .D(net2972),
    .Q_N(_07896_),
    .Q(\m_sys.m_core.m_gpr._GEN[147] ));
 sg13g2_dfrbp_1 _19673_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net521),
    .D(_01491_),
    .Q_N(_07895_),
    .Q(\m_sys.m_core.m_gpr._GEN[148] ));
 sg13g2_dfrbp_1 _19674_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net520),
    .D(_01492_),
    .Q_N(_07894_),
    .Q(\m_sys.m_core.m_gpr._GEN[149] ));
 sg13g2_dfrbp_1 _19675_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net519),
    .D(_01493_),
    .Q_N(_07893_),
    .Q(\m_sys.m_core.m_gpr._GEN[150] ));
 sg13g2_dfrbp_1 _19676_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net518),
    .D(net3074),
    .Q_N(_07892_),
    .Q(\m_sys.m_core.m_gpr._GEN[151] ));
 sg13g2_dfrbp_1 _19677_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net517),
    .D(_01495_),
    .Q_N(_07891_),
    .Q(\m_sys.m_core.m_gpr._GEN[152] ));
 sg13g2_dfrbp_1 _19678_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net516),
    .D(net3015),
    .Q_N(_07890_),
    .Q(\m_sys.m_core.m_gpr._GEN[153] ));
 sg13g2_dfrbp_1 _19679_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net515),
    .D(_01497_),
    .Q_N(_07889_),
    .Q(\m_sys.m_core.m_gpr._GEN[154] ));
 sg13g2_dfrbp_1 _19680_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net514),
    .D(_01498_),
    .Q_N(_07888_),
    .Q(\m_sys.m_core.m_gpr._GEN[155] ));
 sg13g2_dfrbp_1 _19681_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net513),
    .D(net2950),
    .Q_N(_07887_),
    .Q(\m_sys.m_core.m_gpr._GEN[156] ));
 sg13g2_dfrbp_1 _19682_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net512),
    .D(_01500_),
    .Q_N(_07886_),
    .Q(\m_sys.m_core.m_gpr._GEN[157] ));
 sg13g2_dfrbp_1 _19683_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net511),
    .D(net2860),
    .Q_N(_07885_),
    .Q(\m_sys.m_core.m_gpr._GEN[158] ));
 sg13g2_dfrbp_1 _19684_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net510),
    .D(net3035),
    .Q_N(_07884_),
    .Q(\m_sys.m_core.m_gpr._GEN[159] ));
 sg13g2_dfrbp_1 _19685_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net509),
    .D(net3012),
    .Q_N(_07883_),
    .Q(\m_sys.m_core.m_gpr._GEN[96] ));
 sg13g2_dfrbp_1 _19686_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net508),
    .D(net3060),
    .Q_N(_07882_),
    .Q(\m_sys.m_core.m_gpr._GEN[97] ));
 sg13g2_dfrbp_1 _19687_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net507),
    .D(net2901),
    .Q_N(_07881_),
    .Q(\m_sys.m_core.m_gpr._GEN[98] ));
 sg13g2_dfrbp_1 _19688_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net506),
    .D(_01506_),
    .Q_N(_07880_),
    .Q(\m_sys.m_core.m_gpr._GEN[99] ));
 sg13g2_dfrbp_1 _19689_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net505),
    .D(_01507_),
    .Q_N(_07879_),
    .Q(\m_sys.m_core.m_gpr._GEN[100] ));
 sg13g2_dfrbp_1 _19690_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net504),
    .D(net3025),
    .Q_N(_07878_),
    .Q(\m_sys.m_core.m_gpr._GEN[101] ));
 sg13g2_dfrbp_1 _19691_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net503),
    .D(_01509_),
    .Q_N(_07877_),
    .Q(\m_sys.m_core.m_gpr._GEN[102] ));
 sg13g2_dfrbp_1 _19692_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net502),
    .D(_01510_),
    .Q_N(_07876_),
    .Q(\m_sys.m_core.m_gpr._GEN[103] ));
 sg13g2_dfrbp_1 _19693_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net501),
    .D(_01511_),
    .Q_N(_07875_),
    .Q(\m_sys.m_core.m_gpr._GEN[104] ));
 sg13g2_dfrbp_1 _19694_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net500),
    .D(_01512_),
    .Q_N(_07874_),
    .Q(\m_sys.m_core.m_gpr._GEN[105] ));
 sg13g2_dfrbp_1 _19695_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net499),
    .D(net3010),
    .Q_N(_07873_),
    .Q(\m_sys.m_core.m_gpr._GEN[106] ));
 sg13g2_dfrbp_1 _19696_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net498),
    .D(_01514_),
    .Q_N(_07872_),
    .Q(\m_sys.m_core.m_gpr._GEN[107] ));
 sg13g2_dfrbp_1 _19697_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net497),
    .D(_01515_),
    .Q_N(_07871_),
    .Q(\m_sys.m_core.m_gpr._GEN[108] ));
 sg13g2_dfrbp_1 _19698_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net496),
    .D(_01516_),
    .Q_N(_07870_),
    .Q(\m_sys.m_core.m_gpr._GEN[109] ));
 sg13g2_dfrbp_1 _19699_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net495),
    .D(_01517_),
    .Q_N(_07869_),
    .Q(\m_sys.m_core.m_gpr._GEN[110] ));
 sg13g2_dfrbp_1 _19700_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net494),
    .D(_01518_),
    .Q_N(_07868_),
    .Q(\m_sys.m_core.m_gpr._GEN[111] ));
 sg13g2_dfrbp_1 _19701_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net493),
    .D(_01519_),
    .Q_N(_07867_),
    .Q(\m_sys.m_core.m_gpr._GEN[112] ));
 sg13g2_dfrbp_1 _19702_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net492),
    .D(_01520_),
    .Q_N(_07866_),
    .Q(\m_sys.m_core.m_gpr._GEN[113] ));
 sg13g2_dfrbp_1 _19703_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net491),
    .D(_01521_),
    .Q_N(_07865_),
    .Q(\m_sys.m_core.m_gpr._GEN[114] ));
 sg13g2_dfrbp_1 _19704_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net490),
    .D(_01522_),
    .Q_N(_07864_),
    .Q(\m_sys.m_core.m_gpr._GEN[115] ));
 sg13g2_dfrbp_1 _19705_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net489),
    .D(_01523_),
    .Q_N(_07863_),
    .Q(\m_sys.m_core.m_gpr._GEN[116] ));
 sg13g2_dfrbp_1 _19706_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net488),
    .D(_01524_),
    .Q_N(_07862_),
    .Q(\m_sys.m_core.m_gpr._GEN[117] ));
 sg13g2_dfrbp_1 _19707_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net487),
    .D(_01525_),
    .Q_N(_07861_),
    .Q(\m_sys.m_core.m_gpr._GEN[118] ));
 sg13g2_dfrbp_1 _19708_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net486),
    .D(_01526_),
    .Q_N(_07860_),
    .Q(\m_sys.m_core.m_gpr._GEN[119] ));
 sg13g2_dfrbp_1 _19709_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net485),
    .D(_01527_),
    .Q_N(_07859_),
    .Q(\m_sys.m_core.m_gpr._GEN[120] ));
 sg13g2_dfrbp_1 _19710_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net484),
    .D(_01528_),
    .Q_N(_07858_),
    .Q(\m_sys.m_core.m_gpr._GEN[121] ));
 sg13g2_dfrbp_1 _19711_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net483),
    .D(_01529_),
    .Q_N(_07857_),
    .Q(\m_sys.m_core.m_gpr._GEN[122] ));
 sg13g2_dfrbp_1 _19712_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net482),
    .D(_01530_),
    .Q_N(_07856_),
    .Q(\m_sys.m_core.m_gpr._GEN[123] ));
 sg13g2_dfrbp_1 _19713_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net481),
    .D(net3030),
    .Q_N(_07855_),
    .Q(\m_sys.m_core.m_gpr._GEN[124] ));
 sg13g2_dfrbp_1 _19714_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net480),
    .D(_01532_),
    .Q_N(_07854_),
    .Q(\m_sys.m_core.m_gpr._GEN[125] ));
 sg13g2_dfrbp_1 _19715_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net479),
    .D(net2969),
    .Q_N(_07853_),
    .Q(\m_sys.m_core.m_gpr._GEN[126] ));
 sg13g2_dfrbp_1 _19716_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net478),
    .D(net2995),
    .Q_N(_07852_),
    .Q(\m_sys.m_core.m_gpr._GEN[127] ));
 sg13g2_dfrbp_1 _19717_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net477),
    .D(net1981),
    .Q_N(_07851_),
    .Q(\m_sys.m_core.m_gpr._GEN[64] ));
 sg13g2_dfrbp_1 _19718_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net476),
    .D(_01536_),
    .Q_N(_07850_),
    .Q(\m_sys.m_core.m_gpr._GEN[65] ));
 sg13g2_dfrbp_1 _19719_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net475),
    .D(_01537_),
    .Q_N(_07849_),
    .Q(\m_sys.m_core.m_gpr._GEN[66] ));
 sg13g2_dfrbp_1 _19720_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net474),
    .D(_01538_),
    .Q_N(_07848_),
    .Q(\m_sys.m_core.m_gpr._GEN[67] ));
 sg13g2_dfrbp_1 _19721_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net473),
    .D(_01539_),
    .Q_N(_07847_),
    .Q(\m_sys.m_core.m_gpr._GEN[68] ));
 sg13g2_dfrbp_1 _19722_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net472),
    .D(_01540_),
    .Q_N(_07846_),
    .Q(\m_sys.m_core.m_gpr._GEN[69] ));
 sg13g2_dfrbp_1 _19723_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net471),
    .D(_01541_),
    .Q_N(_07845_),
    .Q(\m_sys.m_core.m_gpr._GEN[70] ));
 sg13g2_dfrbp_1 _19724_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net470),
    .D(_01542_),
    .Q_N(_07844_),
    .Q(\m_sys.m_core.m_gpr._GEN[71] ));
 sg13g2_dfrbp_1 _19725_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net469),
    .D(_01543_),
    .Q_N(_07843_),
    .Q(\m_sys.m_core.m_gpr._GEN[72] ));
 sg13g2_dfrbp_1 _19726_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net468),
    .D(_01544_),
    .Q_N(_07842_),
    .Q(\m_sys.m_core.m_gpr._GEN[73] ));
 sg13g2_dfrbp_1 _19727_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net467),
    .D(net2332),
    .Q_N(_07841_),
    .Q(\m_sys.m_core.m_gpr._GEN[74] ));
 sg13g2_dfrbp_1 _19728_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net466),
    .D(_01546_),
    .Q_N(_07840_),
    .Q(\m_sys.m_core.m_gpr._GEN[75] ));
 sg13g2_dfrbp_1 _19729_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net465),
    .D(_01547_),
    .Q_N(_07839_),
    .Q(\m_sys.m_core.m_gpr._GEN[76] ));
 sg13g2_dfrbp_1 _19730_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net464),
    .D(_01548_),
    .Q_N(_07838_),
    .Q(\m_sys.m_core.m_gpr._GEN[77] ));
 sg13g2_dfrbp_1 _19731_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net463),
    .D(_01549_),
    .Q_N(_07837_),
    .Q(\m_sys.m_core.m_gpr._GEN[78] ));
 sg13g2_dfrbp_1 _19732_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net462),
    .D(_01550_),
    .Q_N(_07836_),
    .Q(\m_sys.m_core.m_gpr._GEN[79] ));
 sg13g2_dfrbp_1 _19733_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net461),
    .D(_01551_),
    .Q_N(_07835_),
    .Q(\m_sys.m_core.m_gpr._GEN[80] ));
 sg13g2_dfrbp_1 _19734_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net460),
    .D(_01552_),
    .Q_N(_07834_),
    .Q(\m_sys.m_core.m_gpr._GEN[81] ));
 sg13g2_dfrbp_1 _19735_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net459),
    .D(_01553_),
    .Q_N(_07833_),
    .Q(\m_sys.m_core.m_gpr._GEN[82] ));
 sg13g2_dfrbp_1 _19736_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net458),
    .D(_01554_),
    .Q_N(_07832_),
    .Q(\m_sys.m_core.m_gpr._GEN[83] ));
 sg13g2_dfrbp_1 _19737_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net457),
    .D(_01555_),
    .Q_N(_07831_),
    .Q(\m_sys.m_core.m_gpr._GEN[84] ));
 sg13g2_dfrbp_1 _19738_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net456),
    .D(_01556_),
    .Q_N(_07830_),
    .Q(\m_sys.m_core.m_gpr._GEN[85] ));
 sg13g2_dfrbp_1 _19739_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net455),
    .D(_01557_),
    .Q_N(_07829_),
    .Q(\m_sys.m_core.m_gpr._GEN[86] ));
 sg13g2_dfrbp_1 _19740_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net454),
    .D(_01558_),
    .Q_N(_07828_),
    .Q(\m_sys.m_core.m_gpr._GEN[87] ));
 sg13g2_dfrbp_1 _19741_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net453),
    .D(_01559_),
    .Q_N(_07827_),
    .Q(\m_sys.m_core.m_gpr._GEN[88] ));
 sg13g2_dfrbp_1 _19742_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net452),
    .D(_01560_),
    .Q_N(_07826_),
    .Q(\m_sys.m_core.m_gpr._GEN[89] ));
 sg13g2_dfrbp_1 _19743_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net451),
    .D(_01561_),
    .Q_N(_07825_),
    .Q(\m_sys.m_core.m_gpr._GEN[90] ));
 sg13g2_dfrbp_1 _19744_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net450),
    .D(net2826),
    .Q_N(_07824_),
    .Q(\m_sys.m_core.m_gpr._GEN[91] ));
 sg13g2_dfrbp_1 _19745_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net449),
    .D(net2135),
    .Q_N(_07823_),
    .Q(\m_sys.m_core.m_gpr._GEN[92] ));
 sg13g2_dfrbp_1 _19746_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net448),
    .D(_01564_),
    .Q_N(_07822_),
    .Q(\m_sys.m_core.m_gpr._GEN[93] ));
 sg13g2_dfrbp_1 _19747_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net447),
    .D(net2131),
    .Q_N(_07821_),
    .Q(\m_sys.m_core.m_gpr._GEN[94] ));
 sg13g2_dfrbp_1 _19748_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net446),
    .D(net2385),
    .Q_N(_07820_),
    .Q(\m_sys.m_core.m_gpr._GEN[95] ));
 sg13g2_dfrbp_1 _19749_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net445),
    .D(net2032),
    .Q_N(_07819_),
    .Q(\m_sys.m_core.m_gpr._GEN[32] ));
 sg13g2_dfrbp_1 _19750_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net444),
    .D(_01568_),
    .Q_N(_07818_),
    .Q(\m_sys.m_core.m_gpr._GEN[33] ));
 sg13g2_dfrbp_1 _19751_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net443),
    .D(_01569_),
    .Q_N(_07817_),
    .Q(\m_sys.m_core.m_gpr._GEN[34] ));
 sg13g2_dfrbp_1 _19752_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net442),
    .D(_01570_),
    .Q_N(_07816_),
    .Q(\m_sys.m_core.m_gpr._GEN[35] ));
 sg13g2_dfrbp_1 _19753_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net433),
    .D(_01571_),
    .Q_N(_07815_),
    .Q(\m_sys.m_core.m_gpr._GEN[36] ));
 sg13g2_dfrbp_1 _19754_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net431),
    .D(_01572_),
    .Q_N(_07814_),
    .Q(\m_sys.m_core.m_gpr._GEN[37] ));
 sg13g2_dfrbp_1 _19755_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net421),
    .D(_01573_),
    .Q_N(_07813_),
    .Q(\m_sys.m_core.m_gpr._GEN[38] ));
 sg13g2_dfrbp_1 _19756_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net419),
    .D(_01574_),
    .Q_N(_07812_),
    .Q(\m_sys.m_core.m_gpr._GEN[39] ));
 sg13g2_dfrbp_1 _19757_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net417),
    .D(_01575_),
    .Q_N(_07811_),
    .Q(\m_sys.m_core.m_gpr._GEN[40] ));
 sg13g2_dfrbp_1 _19758_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net415),
    .D(_01576_),
    .Q_N(_07810_),
    .Q(\m_sys.m_core.m_gpr._GEN[41] ));
 sg13g2_dfrbp_1 _19759_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net413),
    .D(net2487),
    .Q_N(_07809_),
    .Q(\m_sys.m_core.m_gpr._GEN[42] ));
 sg13g2_dfrbp_1 _19760_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net411),
    .D(_01578_),
    .Q_N(_07808_),
    .Q(\m_sys.m_core.m_gpr._GEN[43] ));
 sg13g2_dfrbp_1 _19761_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net409),
    .D(_01579_),
    .Q_N(_07807_),
    .Q(\m_sys.m_core.m_gpr._GEN[44] ));
 sg13g2_dfrbp_1 _19762_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net407),
    .D(_01580_),
    .Q_N(_07806_),
    .Q(\m_sys.m_core.m_gpr._GEN[45] ));
 sg13g2_dfrbp_1 _19763_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net405),
    .D(_01581_),
    .Q_N(_07805_),
    .Q(\m_sys.m_core.m_gpr._GEN[46] ));
 sg13g2_dfrbp_1 _19764_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net403),
    .D(_01582_),
    .Q_N(_07804_),
    .Q(\m_sys.m_core.m_gpr._GEN[47] ));
 sg13g2_dfrbp_1 _19765_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net401),
    .D(_01583_),
    .Q_N(_07803_),
    .Q(\m_sys.m_core.m_gpr._GEN[48] ));
 sg13g2_dfrbp_1 _19766_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net399),
    .D(_01584_),
    .Q_N(_07802_),
    .Q(\m_sys.m_core.m_gpr._GEN[49] ));
 sg13g2_dfrbp_1 _19767_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net397),
    .D(_01585_),
    .Q_N(_07801_),
    .Q(\m_sys.m_core.m_gpr._GEN[50] ));
 sg13g2_dfrbp_1 _19768_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net395),
    .D(_01586_),
    .Q_N(_07800_),
    .Q(\m_sys.m_core.m_gpr._GEN[51] ));
 sg13g2_dfrbp_1 _19769_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net393),
    .D(_01587_),
    .Q_N(_07799_),
    .Q(\m_sys.m_core.m_gpr._GEN[52] ));
 sg13g2_dfrbp_1 _19770_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net391),
    .D(_01588_),
    .Q_N(_07798_),
    .Q(\m_sys.m_core.m_gpr._GEN[53] ));
 sg13g2_dfrbp_1 _19771_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net389),
    .D(_01589_),
    .Q_N(_07797_),
    .Q(\m_sys.m_core.m_gpr._GEN[54] ));
 sg13g2_dfrbp_1 _19772_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net387),
    .D(_01590_),
    .Q_N(_07796_),
    .Q(\m_sys.m_core.m_gpr._GEN[55] ));
 sg13g2_dfrbp_1 _19773_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net385),
    .D(_01591_),
    .Q_N(_07795_),
    .Q(\m_sys.m_core.m_gpr._GEN[56] ));
 sg13g2_dfrbp_1 _19774_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net383),
    .D(_01592_),
    .Q_N(_07794_),
    .Q(\m_sys.m_core.m_gpr._GEN[57] ));
 sg13g2_dfrbp_1 _19775_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net381),
    .D(_01593_),
    .Q_N(_07793_),
    .Q(\m_sys.m_core.m_gpr._GEN[58] ));
 sg13g2_dfrbp_1 _19776_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net379),
    .D(_01594_),
    .Q_N(_07792_),
    .Q(\m_sys.m_core.m_gpr._GEN[59] ));
 sg13g2_dfrbp_1 _19777_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net377),
    .D(net2685),
    .Q_N(_07791_),
    .Q(\m_sys.m_core.m_gpr._GEN[60] ));
 sg13g2_dfrbp_1 _19778_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net375),
    .D(_01596_),
    .Q_N(_07790_),
    .Q(\m_sys.m_core.m_gpr._GEN[61] ));
 sg13g2_dfrbp_1 _19779_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net373),
    .D(net2838),
    .Q_N(_07789_),
    .Q(\m_sys.m_core.m_gpr._GEN[62] ));
 sg13g2_dfrbp_1 _19780_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net371),
    .D(net2787),
    .Q_N(_07788_),
    .Q(\m_sys.m_core.m_gpr._GEN[63] ));
 sg13g2_dfrbp_1 _19781_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net369),
    .D(net3265),
    .Q_N(_07787_),
    .Q(\m_sys.m_core.m_fsm.r_cstate[0] ));
 sg13g2_dfrbp_1 _19782_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net367),
    .D(net2769),
    .Q_N(_07786_),
    .Q(\m_sys.m_core.m_gpr._GEN[160] ));
 sg13g2_dfrbp_1 _19783_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net365),
    .D(_01601_),
    .Q_N(_07785_),
    .Q(\m_sys.m_core.m_gpr._GEN[161] ));
 sg13g2_dfrbp_1 _19784_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net363),
    .D(_01602_),
    .Q_N(_07784_),
    .Q(\m_sys.m_core.m_gpr._GEN[162] ));
 sg13g2_dfrbp_1 _19785_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net361),
    .D(_01603_),
    .Q_N(_07783_),
    .Q(\m_sys.m_core.m_gpr._GEN[163] ));
 sg13g2_dfrbp_1 _19786_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net327),
    .D(_01604_),
    .Q_N(_07782_),
    .Q(\m_sys.m_core.m_gpr._GEN[164] ));
 sg13g2_dfrbp_1 _19787_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net325),
    .D(_01605_),
    .Q_N(_07781_),
    .Q(\m_sys.m_core.m_gpr._GEN[165] ));
 sg13g2_dfrbp_1 _19788_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net323),
    .D(_01606_),
    .Q_N(_07780_),
    .Q(\m_sys.m_core.m_gpr._GEN[166] ));
 sg13g2_dfrbp_1 _19789_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net321),
    .D(_01607_),
    .Q_N(_07779_),
    .Q(\m_sys.m_core.m_gpr._GEN[167] ));
 sg13g2_dfrbp_1 _19790_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net148),
    .D(_01608_),
    .Q_N(_07778_),
    .Q(\m_sys.m_core.m_gpr._GEN[168] ));
 sg13g2_dfrbp_1 _19791_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net146),
    .D(_01609_),
    .Q_N(_07777_),
    .Q(\m_sys.m_core.m_gpr._GEN[169] ));
 sg13g2_dfrbp_1 _19792_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net144),
    .D(net2726),
    .Q_N(_07776_),
    .Q(\m_sys.m_core.m_gpr._GEN[170] ));
 sg13g2_dfrbp_1 _19793_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net142),
    .D(_01611_),
    .Q_N(_07775_),
    .Q(\m_sys.m_core.m_gpr._GEN[171] ));
 sg13g2_dfrbp_1 _19794_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1529),
    .D(_01612_),
    .Q_N(_07774_),
    .Q(\m_sys.m_core.m_gpr._GEN[172] ));
 sg13g2_dfrbp_1 _19795_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1527),
    .D(_01613_),
    .Q_N(_07773_),
    .Q(\m_sys.m_core.m_gpr._GEN[173] ));
 sg13g2_dfrbp_1 _19796_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1525),
    .D(_01614_),
    .Q_N(_07772_),
    .Q(\m_sys.m_core.m_gpr._GEN[174] ));
 sg13g2_dfrbp_1 _19797_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1523),
    .D(_01615_),
    .Q_N(_07771_),
    .Q(\m_sys.m_core.m_gpr._GEN[175] ));
 sg13g2_dfrbp_1 _19798_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1521),
    .D(_01616_),
    .Q_N(_07770_),
    .Q(\m_sys.m_core.m_gpr._GEN[176] ));
 sg13g2_dfrbp_1 _19799_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1519),
    .D(_01617_),
    .Q_N(_07769_),
    .Q(\m_sys.m_core.m_gpr._GEN[177] ));
 sg13g2_dfrbp_1 _19800_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1517),
    .D(_01618_),
    .Q_N(_07768_),
    .Q(\m_sys.m_core.m_gpr._GEN[178] ));
 sg13g2_dfrbp_1 _19801_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1515),
    .D(_01619_),
    .Q_N(_07767_),
    .Q(\m_sys.m_core.m_gpr._GEN[179] ));
 sg13g2_dfrbp_1 _19802_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1513),
    .D(_01620_),
    .Q_N(_07766_),
    .Q(\m_sys.m_core.m_gpr._GEN[180] ));
 sg13g2_dfrbp_1 _19803_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1511),
    .D(_01621_),
    .Q_N(_07765_),
    .Q(\m_sys.m_core.m_gpr._GEN[181] ));
 sg13g2_dfrbp_1 _19804_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1445),
    .D(_01622_),
    .Q_N(_07764_),
    .Q(\m_sys.m_core.m_gpr._GEN[182] ));
 sg13g2_dfrbp_1 _19805_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1147),
    .D(_01623_),
    .Q_N(_07763_),
    .Q(\m_sys.m_core.m_gpr._GEN[183] ));
 sg13g2_dfrbp_1 _19806_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1145),
    .D(_01624_),
    .Q_N(_07762_),
    .Q(\m_sys.m_core.m_gpr._GEN[184] ));
 sg13g2_dfrbp_1 _19807_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1143),
    .D(_01625_),
    .Q_N(_07761_),
    .Q(\m_sys.m_core.m_gpr._GEN[185] ));
 sg13g2_dfrbp_1 _19808_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1133),
    .D(_01626_),
    .Q_N(_07760_),
    .Q(\m_sys.m_core.m_gpr._GEN[186] ));
 sg13g2_dfrbp_1 _19809_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1131),
    .D(_01627_),
    .Q_N(_07759_),
    .Q(\m_sys.m_core.m_gpr._GEN[187] ));
 sg13g2_dfrbp_1 _19810_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1129),
    .D(net2872),
    .Q_N(_07758_),
    .Q(\m_sys.m_core.m_gpr._GEN[188] ));
 sg13g2_dfrbp_1 _19811_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1127),
    .D(_01629_),
    .Q_N(_07757_),
    .Q(\m_sys.m_core.m_gpr._GEN[189] ));
 sg13g2_dfrbp_1 _19812_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1109),
    .D(net2474),
    .Q_N(_07756_),
    .Q(\m_sys.m_core.m_gpr._GEN[190] ));
 sg13g2_dfrbp_1 _19813_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1107),
    .D(net2576),
    .Q_N(_07755_),
    .Q(\m_sys.m_core.m_gpr._GEN[191] ));
 sg13g2_dfrbp_1 _19814_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1105),
    .D(net3132),
    .Q_N(_07754_),
    .Q(\m_sys.m_core.m_gpr._GEN[192] ));
 sg13g2_dfrbp_1 _19815_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1103),
    .D(_01633_),
    .Q_N(_07753_),
    .Q(\m_sys.m_core.m_gpr._GEN[193] ));
 sg13g2_dfrbp_1 _19816_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1101),
    .D(_01634_),
    .Q_N(_07752_),
    .Q(\m_sys.m_core.m_gpr._GEN[194] ));
 sg13g2_dfrbp_1 _19817_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1099),
    .D(_01635_),
    .Q_N(_07751_),
    .Q(\m_sys.m_core.m_gpr._GEN[195] ));
 sg13g2_dfrbp_1 _19818_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1096),
    .D(_01636_),
    .Q_N(_07750_),
    .Q(\m_sys.m_core.m_gpr._GEN[196] ));
 sg13g2_dfrbp_1 _19819_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1094),
    .D(_01637_),
    .Q_N(_07749_),
    .Q(\m_sys.m_core.m_gpr._GEN[197] ));
 sg13g2_dfrbp_1 _19820_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1092),
    .D(net2796),
    .Q_N(_07748_),
    .Q(\m_sys.m_core.m_gpr._GEN[198] ));
 sg13g2_dfrbp_1 _19821_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1090),
    .D(net2869),
    .Q_N(_07747_),
    .Q(\m_sys.m_core.m_gpr._GEN[199] ));
 sg13g2_dfrbp_1 _19822_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1088),
    .D(_01640_),
    .Q_N(_07746_),
    .Q(\m_sys.m_core.m_gpr._GEN[200] ));
 sg13g2_dfrbp_1 _19823_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1086),
    .D(net2919),
    .Q_N(_07745_),
    .Q(\m_sys.m_core.m_gpr._GEN[201] ));
 sg13g2_dfrbp_1 _19824_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1084),
    .D(net2322),
    .Q_N(_07744_),
    .Q(\m_sys.m_core.m_gpr._GEN[202] ));
 sg13g2_dfrbp_1 _19825_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1082),
    .D(_01643_),
    .Q_N(_07743_),
    .Q(\m_sys.m_core.m_gpr._GEN[203] ));
 sg13g2_dfrbp_1 _19826_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1027),
    .D(_01644_),
    .Q_N(_07742_),
    .Q(\m_sys.m_core.m_gpr._GEN[204] ));
 sg13g2_dfrbp_1 _19827_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1013),
    .D(_01645_),
    .Q_N(_07741_),
    .Q(\m_sys.m_core.m_gpr._GEN[205] ));
 sg13g2_dfrbp_1 _19828_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1011),
    .D(_01646_),
    .Q_N(_07740_),
    .Q(\m_sys.m_core.m_gpr._GEN[206] ));
 sg13g2_dfrbp_1 _19829_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1009),
    .D(_01647_),
    .Q_N(_07739_),
    .Q(\m_sys.m_core.m_gpr._GEN[207] ));
 sg13g2_dfrbp_1 _19830_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1007),
    .D(_01648_),
    .Q_N(_07738_),
    .Q(\m_sys.m_core.m_gpr._GEN[208] ));
 sg13g2_dfrbp_1 _19831_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1005),
    .D(_01649_),
    .Q_N(_07737_),
    .Q(\m_sys.m_core.m_gpr._GEN[209] ));
 sg13g2_dfrbp_1 _19832_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1003),
    .D(_01650_),
    .Q_N(_07736_),
    .Q(\m_sys.m_core.m_gpr._GEN[210] ));
 sg13g2_dfrbp_1 _19833_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1001),
    .D(_01651_),
    .Q_N(_07735_),
    .Q(\m_sys.m_core.m_gpr._GEN[211] ));
 sg13g2_dfrbp_1 _19834_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net999),
    .D(_01652_),
    .Q_N(_07734_),
    .Q(\m_sys.m_core.m_gpr._GEN[212] ));
 sg13g2_dfrbp_1 _19835_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net997),
    .D(net2845),
    .Q_N(_07733_),
    .Q(\m_sys.m_core.m_gpr._GEN[213] ));
 sg13g2_dfrbp_1 _19836_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net995),
    .D(_01654_),
    .Q_N(_07732_),
    .Q(\m_sys.m_core.m_gpr._GEN[214] ));
 sg13g2_dfrbp_1 _19837_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net993),
    .D(_01655_),
    .Q_N(_07731_),
    .Q(\m_sys.m_core.m_gpr._GEN[215] ));
 sg13g2_dfrbp_1 _19838_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net991),
    .D(_01656_),
    .Q_N(_07730_),
    .Q(\m_sys.m_core.m_gpr._GEN[216] ));
 sg13g2_dfrbp_1 _19839_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net989),
    .D(_01657_),
    .Q_N(_07729_),
    .Q(\m_sys.m_core.m_gpr._GEN[217] ));
 sg13g2_dfrbp_1 _19840_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net987),
    .D(_01658_),
    .Q_N(_07728_),
    .Q(\m_sys.m_core.m_gpr._GEN[218] ));
 sg13g2_dfrbp_1 _19841_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net985),
    .D(_01659_),
    .Q_N(_07727_),
    .Q(\m_sys.m_core.m_gpr._GEN[219] ));
 sg13g2_dfrbp_1 _19842_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net983),
    .D(net1965),
    .Q_N(_07726_),
    .Q(\m_sys.m_core.m_gpr._GEN[220] ));
 sg13g2_dfrbp_1 _19843_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net981),
    .D(_01661_),
    .Q_N(_07725_),
    .Q(\m_sys.m_core.m_gpr._GEN[221] ));
 sg13g2_dfrbp_1 _19844_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net979),
    .D(net2750),
    .Q_N(_07724_),
    .Q(\m_sys.m_core.m_gpr._GEN[222] ));
 sg13g2_dfrbp_1 _19845_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net977),
    .D(net2722),
    .Q_N(_07723_),
    .Q(\m_sys.m_core.m_gpr._GEN[223] ));
 sg13g2_dfrbp_1 _19846_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net975),
    .D(_01664_),
    .Q_N(_07722_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][16] ));
 sg13g2_dfrbp_1 _19847_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net973),
    .D(_01665_),
    .Q_N(_07721_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][17] ));
 sg13g2_dfrbp_1 _19848_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net971),
    .D(_01666_),
    .Q_N(_07720_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][18] ));
 sg13g2_dfrbp_1 _19849_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net969),
    .D(_01667_),
    .Q_N(_07719_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][19] ));
 sg13g2_dfrbp_1 _19850_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net967),
    .D(_01668_),
    .Q_N(_07718_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][20] ));
 sg13g2_dfrbp_1 _19851_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net965),
    .D(_01669_),
    .Q_N(_07717_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][21] ));
 sg13g2_dfrbp_1 _19852_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net963),
    .D(_01670_),
    .Q_N(_07716_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][22] ));
 sg13g2_dfrbp_1 _19853_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net961),
    .D(_01671_),
    .Q_N(_07715_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][23] ));
 sg13g2_dfrbp_1 _19854_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net959),
    .D(_01672_),
    .Q_N(_07714_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][0] ));
 sg13g2_dfrbp_1 _19855_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net957),
    .D(_01673_),
    .Q_N(_07713_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][1] ));
 sg13g2_dfrbp_1 _19856_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net955),
    .D(_01674_),
    .Q_N(_07712_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][2] ));
 sg13g2_dfrbp_1 _19857_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net953),
    .D(_01675_),
    .Q_N(_07711_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][3] ));
 sg13g2_dfrbp_1 _19858_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net951),
    .D(_01676_),
    .Q_N(_07710_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][4] ));
 sg13g2_dfrbp_1 _19859_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net941),
    .D(_01677_),
    .Q_N(_07709_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][5] ));
 sg13g2_dfrbp_1 _19860_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net939),
    .D(_01678_),
    .Q_N(_07708_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][6] ));
 sg13g2_dfrbp_1 _19861_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net937),
    .D(_01679_),
    .Q_N(_07707_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][7] ));
 sg13g2_dfrbp_1 _19862_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net935),
    .D(_01680_),
    .Q_N(_07706_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][8] ));
 sg13g2_dfrbp_1 _19863_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net933),
    .D(_01681_),
    .Q_N(_07705_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][9] ));
 sg13g2_dfrbp_1 _19864_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net931),
    .D(_01682_),
    .Q_N(_07704_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][10] ));
 sg13g2_dfrbp_1 _19865_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net929),
    .D(_01683_),
    .Q_N(_07703_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][11] ));
 sg13g2_dfrbp_1 _19866_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net927),
    .D(_01684_),
    .Q_N(_07702_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][12] ));
 sg13g2_dfrbp_1 _19867_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net925),
    .D(_01685_),
    .Q_N(_07701_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][13] ));
 sg13g2_dfrbp_1 _19868_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net923),
    .D(_01686_),
    .Q_N(_07700_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][14] ));
 sg13g2_dfrbp_1 _19869_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net921),
    .D(_01687_),
    .Q_N(_07699_),
    .Q(\m_sys.m_ram.m_ram.r_mem[5][15] ));
 sg13g2_dfrbp_1 _19870_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net919),
    .D(_01688_),
    .Q_N(_07698_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][8] ));
 sg13g2_dfrbp_1 _19871_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net917),
    .D(_01689_),
    .Q_N(_07697_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][9] ));
 sg13g2_dfrbp_1 _19872_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net915),
    .D(_01690_),
    .Q_N(_07696_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][10] ));
 sg13g2_dfrbp_1 _19873_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net913),
    .D(_01691_),
    .Q_N(_07695_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][11] ));
 sg13g2_dfrbp_1 _19874_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net911),
    .D(_01692_),
    .Q_N(_07694_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][12] ));
 sg13g2_dfrbp_1 _19875_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net900),
    .D(_01693_),
    .Q_N(_07693_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][13] ));
 sg13g2_dfrbp_1 _19876_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net898),
    .D(_01694_),
    .Q_N(_07692_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][14] ));
 sg13g2_dfrbp_1 _19877_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net896),
    .D(_01695_),
    .Q_N(_07691_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][15] ));
 sg13g2_dfrbp_1 _19878_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net894),
    .D(_01696_),
    .Q_N(_07690_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][16] ));
 sg13g2_dfrbp_1 _19879_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net892),
    .D(_01697_),
    .Q_N(_07689_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][17] ));
 sg13g2_dfrbp_1 _19880_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net890),
    .D(_01698_),
    .Q_N(_07688_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][18] ));
 sg13g2_dfrbp_1 _19881_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net888),
    .D(_01699_),
    .Q_N(_07687_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][19] ));
 sg13g2_dfrbp_1 _19882_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net886),
    .D(_01700_),
    .Q_N(_07686_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][20] ));
 sg13g2_dfrbp_1 _19883_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net884),
    .D(_01701_),
    .Q_N(_07685_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][21] ));
 sg13g2_dfrbp_1 _19884_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net882),
    .D(_01702_),
    .Q_N(_07684_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][22] ));
 sg13g2_dfrbp_1 _19885_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net880),
    .D(_01703_),
    .Q_N(_07683_),
    .Q(\m_sys.m_ram.m_ram.r_mem[6][23] ));
 sg13g2_dfrbp_1 _19886_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net840),
    .D(_01704_),
    .Q_N(_07682_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][0] ));
 sg13g2_dfrbp_1 _19887_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net838),
    .D(_01705_),
    .Q_N(_07681_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][1] ));
 sg13g2_dfrbp_1 _19888_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net836),
    .D(_01706_),
    .Q_N(_07680_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][2] ));
 sg13g2_dfrbp_1 _19889_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net817),
    .D(_01707_),
    .Q_N(_07679_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][3] ));
 sg13g2_dfrbp_1 _19890_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net815),
    .D(_01708_),
    .Q_N(_07678_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][4] ));
 sg13g2_dfrbp_1 _19891_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net813),
    .D(_01709_),
    .Q_N(_07677_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][5] ));
 sg13g2_dfrbp_1 _19892_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net811),
    .D(_01710_),
    .Q_N(_07676_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][6] ));
 sg13g2_dfrbp_1 _19893_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net809),
    .D(_01711_),
    .Q_N(_07675_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][7] ));
 sg13g2_dfrbp_1 _19894_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net807),
    .D(_01712_),
    .Q_N(_07674_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][8] ));
 sg13g2_dfrbp_1 _19895_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net805),
    .D(_01713_),
    .Q_N(_07673_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][9] ));
 sg13g2_dfrbp_1 _19896_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net803),
    .D(_01714_),
    .Q_N(_07672_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][10] ));
 sg13g2_dfrbp_1 _19897_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net769),
    .D(_01715_),
    .Q_N(_07671_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][11] ));
 sg13g2_dfrbp_1 _19898_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net767),
    .D(_01716_),
    .Q_N(_07670_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][12] ));
 sg13g2_dfrbp_1 _19899_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net765),
    .D(_01717_),
    .Q_N(_07669_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][13] ));
 sg13g2_dfrbp_1 _19900_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net763),
    .D(_01718_),
    .Q_N(_07668_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][14] ));
 sg13g2_dfrbp_1 _19901_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net761),
    .D(_01719_),
    .Q_N(_07667_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][15] ));
 sg13g2_dfrbp_1 _19902_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net759),
    .D(_01720_),
    .Q_N(_07666_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][16] ));
 sg13g2_dfrbp_1 _19903_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net757),
    .D(_01721_),
    .Q_N(_07665_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][17] ));
 sg13g2_dfrbp_1 _19904_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net755),
    .D(_01722_),
    .Q_N(_07664_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][18] ));
 sg13g2_dfrbp_1 _19905_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net721),
    .D(_01723_),
    .Q_N(_07663_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][19] ));
 sg13g2_dfrbp_1 _19906_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net719),
    .D(_01724_),
    .Q_N(_07662_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][20] ));
 sg13g2_dfrbp_1 _19907_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net717),
    .D(_01725_),
    .Q_N(_07661_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][21] ));
 sg13g2_dfrbp_1 _19908_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net715),
    .D(_01726_),
    .Q_N(_07660_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][22] ));
 sg13g2_dfrbp_1 _19909_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net713),
    .D(_01727_),
    .Q_N(_07659_),
    .Q(\m_sys.m_ram.m_ram.r_mem[7][23] ));
 sg13g2_dfrbp_1 _19910_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net711),
    .D(_01728_),
    .Q_N(_07658_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][0] ));
 sg13g2_dfrbp_1 _19911_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net709),
    .D(_01729_),
    .Q_N(_07657_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][1] ));
 sg13g2_dfrbp_1 _19912_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net707),
    .D(_01730_),
    .Q_N(_07656_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][2] ));
 sg13g2_dfrbp_1 _19913_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net705),
    .D(_01731_),
    .Q_N(_07655_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][3] ));
 sg13g2_dfrbp_1 _19914_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net703),
    .D(_01732_),
    .Q_N(_07654_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][4] ));
 sg13g2_dfrbp_1 _19915_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net701),
    .D(_01733_),
    .Q_N(_07653_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][5] ));
 sg13g2_dfrbp_1 _19916_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net699),
    .D(_01734_),
    .Q_N(_07652_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][6] ));
 sg13g2_dfrbp_1 _19917_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net697),
    .D(_01735_),
    .Q_N(_07651_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][7] ));
 sg13g2_dfrbp_1 _19918_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net695),
    .D(_01736_),
    .Q_N(_07650_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][8] ));
 sg13g2_dfrbp_1 _19919_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net693),
    .D(_01737_),
    .Q_N(_07649_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][9] ));
 sg13g2_dfrbp_1 _19920_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net691),
    .D(_01738_),
    .Q_N(_07648_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][10] ));
 sg13g2_dfrbp_1 _19921_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net657),
    .D(_01739_),
    .Q_N(_07647_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][11] ));
 sg13g2_dfrbp_1 _19922_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net655),
    .D(_01740_),
    .Q_N(_07646_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][12] ));
 sg13g2_dfrbp_1 _19923_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net653),
    .D(_01741_),
    .Q_N(_07645_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][13] ));
 sg13g2_dfrbp_1 _19924_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net651),
    .D(_01742_),
    .Q_N(_07644_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][14] ));
 sg13g2_dfrbp_1 _19925_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net647),
    .D(_01743_),
    .Q_N(_07643_),
    .Q(\m_sys.m_ram.m_ram.r_mem[8][15] ));
 sg13g2_tiehi _18672__18 (.L_HI(net18));
 sg13g2_tiehi _18671__19 (.L_HI(net19));
 sg13g2_tiehi _18670__20 (.L_HI(net20));
 sg13g2_tiehi _18669__21 (.L_HI(net21));
 sg13g2_tiehi _18668__22 (.L_HI(net22));
 sg13g2_tiehi _18667__23 (.L_HI(net23));
 sg13g2_tiehi _18666__24 (.L_HI(net24));
 sg13g2_tiehi _18665__25 (.L_HI(net25));
 sg13g2_tiehi _18664__26 (.L_HI(net26));
 sg13g2_tiehi _18663__27 (.L_HI(net27));
 sg13g2_tiehi _18662__28 (.L_HI(net28));
 sg13g2_tiehi _18661__29 (.L_HI(net29));
 sg13g2_tiehi _18660__30 (.L_HI(net30));
 sg13g2_tiehi _18659__31 (.L_HI(net31));
 sg13g2_tiehi _18658__32 (.L_HI(net32));
 sg13g2_tiehi _18657__33 (.L_HI(net33));
 sg13g2_tiehi _18656__34 (.L_HI(net34));
 sg13g2_tiehi _18655__35 (.L_HI(net35));
 sg13g2_tiehi _18654__36 (.L_HI(net36));
 sg13g2_tiehi _18653__37 (.L_HI(net37));
 sg13g2_tiehi _18652__38 (.L_HI(net38));
 sg13g2_tiehi _18651__39 (.L_HI(net39));
 sg13g2_tiehi _18650__40 (.L_HI(net40));
 sg13g2_tiehi _18649__41 (.L_HI(net41));
 sg13g2_tiehi _18648__42 (.L_HI(net42));
 sg13g2_tiehi _18647__43 (.L_HI(net43));
 sg13g2_tiehi _18646__44 (.L_HI(net44));
 sg13g2_tiehi _18645__45 (.L_HI(net45));
 sg13g2_tiehi _18644__46 (.L_HI(net46));
 sg13g2_tiehi _18643__47 (.L_HI(net47));
 sg13g2_tiehi _18642__48 (.L_HI(net48));
 sg13g2_tiehi _18641__49 (.L_HI(net49));
 sg13g2_tiehi _18640__50 (.L_HI(net50));
 sg13g2_tiehi _18639__51 (.L_HI(net51));
 sg13g2_tiehi _18638__52 (.L_HI(net52));
 sg13g2_tiehi _18637__53 (.L_HI(net53));
 sg13g2_tiehi _18636__54 (.L_HI(net54));
 sg13g2_tiehi _18635__55 (.L_HI(net55));
 sg13g2_tiehi _18634__56 (.L_HI(net56));
 sg13g2_tiehi _18633__57 (.L_HI(net57));
 sg13g2_tiehi _18632__58 (.L_HI(net58));
 sg13g2_tiehi _18631__59 (.L_HI(net59));
 sg13g2_tiehi _18630__60 (.L_HI(net60));
 sg13g2_tiehi _18629__61 (.L_HI(net61));
 sg13g2_tiehi _18628__62 (.L_HI(net62));
 sg13g2_tiehi _18627__63 (.L_HI(net63));
 sg13g2_tiehi _18626__64 (.L_HI(net64));
 sg13g2_tiehi _18625__65 (.L_HI(net65));
 sg13g2_tiehi _18624__66 (.L_HI(net66));
 sg13g2_tiehi _18623__67 (.L_HI(net67));
 sg13g2_tiehi _18622__68 (.L_HI(net68));
 sg13g2_tiehi _18621__69 (.L_HI(net69));
 sg13g2_tiehi _18620__70 (.L_HI(net70));
 sg13g2_tiehi _18619__71 (.L_HI(net71));
 sg13g2_tiehi _18618__72 (.L_HI(net72));
 sg13g2_tiehi _18617__73 (.L_HI(net73));
 sg13g2_tiehi _18616__74 (.L_HI(net74));
 sg13g2_tiehi _18615__75 (.L_HI(net75));
 sg13g2_tiehi _18614__76 (.L_HI(net76));
 sg13g2_tiehi _18613__77 (.L_HI(net77));
 sg13g2_tiehi _18612__78 (.L_HI(net78));
 sg13g2_tiehi _18611__79 (.L_HI(net79));
 sg13g2_tiehi _18610__80 (.L_HI(net80));
 sg13g2_tiehi _18609__81 (.L_HI(net81));
 sg13g2_tiehi _18608__82 (.L_HI(net82));
 sg13g2_tiehi _18607__83 (.L_HI(net83));
 sg13g2_tiehi _18606__84 (.L_HI(net84));
 sg13g2_tiehi _18605__85 (.L_HI(net85));
 sg13g2_tiehi _18604__86 (.L_HI(net86));
 sg13g2_tiehi _18603__87 (.L_HI(net87));
 sg13g2_tiehi _18602__88 (.L_HI(net88));
 sg13g2_tiehi _18601__89 (.L_HI(net89));
 sg13g2_tiehi _18600__90 (.L_HI(net90));
 sg13g2_tiehi _18599__91 (.L_HI(net91));
 sg13g2_tiehi _18598__92 (.L_HI(net92));
 sg13g2_tiehi _18597__93 (.L_HI(net93));
 sg13g2_tiehi _18596__94 (.L_HI(net94));
 sg13g2_tiehi _18595__95 (.L_HI(net95));
 sg13g2_tiehi _18594__96 (.L_HI(net96));
 sg13g2_tiehi _18593__97 (.L_HI(net97));
 sg13g2_tiehi _18592__98 (.L_HI(net98));
 sg13g2_tiehi _18591__99 (.L_HI(net99));
 sg13g2_tiehi _18590__100 (.L_HI(net100));
 sg13g2_tiehi _18589__101 (.L_HI(net101));
 sg13g2_tiehi _18588__102 (.L_HI(net102));
 sg13g2_tiehi _18587__103 (.L_HI(net103));
 sg13g2_tiehi _18586__104 (.L_HI(net104));
 sg13g2_tiehi _18585__105 (.L_HI(net105));
 sg13g2_tiehi _18584__106 (.L_HI(net106));
 sg13g2_tiehi _18583__107 (.L_HI(net107));
 sg13g2_tiehi _18582__108 (.L_HI(net108));
 sg13g2_tiehi _18581__109 (.L_HI(net109));
 sg13g2_tiehi _18580__110 (.L_HI(net110));
 sg13g2_tiehi _18579__111 (.L_HI(net111));
 sg13g2_tiehi _18578__112 (.L_HI(net112));
 sg13g2_tiehi _18577__113 (.L_HI(net113));
 sg13g2_tiehi _18576__114 (.L_HI(net114));
 sg13g2_tiehi _18575__115 (.L_HI(net115));
 sg13g2_tiehi _18574__116 (.L_HI(net116));
 sg13g2_tiehi _18573__117 (.L_HI(net117));
 sg13g2_tiehi _18572__118 (.L_HI(net118));
 sg13g2_tiehi _18571__119 (.L_HI(net119));
 sg13g2_tiehi _18570__120 (.L_HI(net120));
 sg13g2_tiehi _18569__121 (.L_HI(net121));
 sg13g2_tiehi _18568__122 (.L_HI(net122));
 sg13g2_tiehi _18567__123 (.L_HI(net123));
 sg13g2_tiehi _18566__124 (.L_HI(net124));
 sg13g2_tiehi _18565__125 (.L_HI(net125));
 sg13g2_tiehi _18564__126 (.L_HI(net126));
 sg13g2_tiehi _18563__127 (.L_HI(net127));
 sg13g2_tiehi _18562__128 (.L_HI(net128));
 sg13g2_tiehi _18561__129 (.L_HI(net129));
 sg13g2_tiehi _18560__130 (.L_HI(net130));
 sg13g2_tiehi _18559__131 (.L_HI(net131));
 sg13g2_tiehi _18558__132 (.L_HI(net132));
 sg13g2_tiehi _18557__133 (.L_HI(net133));
 sg13g2_tiehi _18556__134 (.L_HI(net134));
 sg13g2_tiehi _18555__135 (.L_HI(net135));
 sg13g2_tiehi _18554__136 (.L_HI(net136));
 sg13g2_tiehi _18553__137 (.L_HI(net137));
 sg13g2_tiehi _18552__138 (.L_HI(net138));
 sg13g2_tiehi _18551__139 (.L_HI(net139));
 sg13g2_tiehi _18550__140 (.L_HI(net140));
 sg13g2_tiehi _18549__141 (.L_HI(net141));
 sg13g2_tiehi _19793__142 (.L_HI(net142));
 sg13g2_tiehi _18548__143 (.L_HI(net143));
 sg13g2_tiehi _19792__144 (.L_HI(net144));
 sg13g2_tiehi _18547__145 (.L_HI(net145));
 sg13g2_tiehi _19791__146 (.L_HI(net146));
 sg13g2_tiehi _18546__147 (.L_HI(net147));
 sg13g2_tiehi _19790__148 (.L_HI(net148));
 sg13g2_tiehi _18545__149 (.L_HI(net149));
 sg13g2_tiehi _18544__150 (.L_HI(net150));
 sg13g2_tiehi _18543__151 (.L_HI(net151));
 sg13g2_tiehi _18542__152 (.L_HI(net152));
 sg13g2_tiehi _18541__153 (.L_HI(net153));
 sg13g2_tiehi _18540__154 (.L_HI(net154));
 sg13g2_tiehi _18539__155 (.L_HI(net155));
 sg13g2_tiehi _18538__156 (.L_HI(net156));
 sg13g2_tiehi _18537__157 (.L_HI(net157));
 sg13g2_tiehi _18536__158 (.L_HI(net158));
 sg13g2_tiehi _18535__159 (.L_HI(net159));
 sg13g2_tiehi _18534__160 (.L_HI(net160));
 sg13g2_tiehi _18533__161 (.L_HI(net161));
 sg13g2_tiehi _18532__162 (.L_HI(net162));
 sg13g2_tiehi _18531__163 (.L_HI(net163));
 sg13g2_tiehi _18530__164 (.L_HI(net164));
 sg13g2_tiehi _18529__165 (.L_HI(net165));
 sg13g2_tiehi _18528__166 (.L_HI(net166));
 sg13g2_tiehi _18527__167 (.L_HI(net167));
 sg13g2_tiehi _18526__168 (.L_HI(net168));
 sg13g2_tiehi _18525__169 (.L_HI(net169));
 sg13g2_tiehi _18524__170 (.L_HI(net170));
 sg13g2_tiehi _18523__171 (.L_HI(net171));
 sg13g2_tiehi _18522__172 (.L_HI(net172));
 sg13g2_tiehi _18521__173 (.L_HI(net173));
 sg13g2_tiehi _18520__174 (.L_HI(net174));
 sg13g2_tiehi _18519__175 (.L_HI(net175));
 sg13g2_tiehi _18518__176 (.L_HI(net176));
 sg13g2_tiehi _18517__177 (.L_HI(net177));
 sg13g2_tiehi _18516__178 (.L_HI(net178));
 sg13g2_tiehi _18515__179 (.L_HI(net179));
 sg13g2_tiehi _18514__180 (.L_HI(net180));
 sg13g2_tiehi _18513__181 (.L_HI(net181));
 sg13g2_tiehi _18512__182 (.L_HI(net182));
 sg13g2_tiehi _18511__183 (.L_HI(net183));
 sg13g2_tiehi _18510__184 (.L_HI(net184));
 sg13g2_tiehi _18509__185 (.L_HI(net185));
 sg13g2_tiehi _18508__186 (.L_HI(net186));
 sg13g2_tiehi _18507__187 (.L_HI(net187));
 sg13g2_tiehi _18506__188 (.L_HI(net188));
 sg13g2_tiehi _18505__189 (.L_HI(net189));
 sg13g2_tiehi _18504__190 (.L_HI(net190));
 sg13g2_tiehi _18503__191 (.L_HI(net191));
 sg13g2_tiehi _18502__192 (.L_HI(net192));
 sg13g2_tiehi _18501__193 (.L_HI(net193));
 sg13g2_tiehi _18500__194 (.L_HI(net194));
 sg13g2_tiehi _18499__195 (.L_HI(net195));
 sg13g2_tiehi _18498__196 (.L_HI(net196));
 sg13g2_tiehi _18497__197 (.L_HI(net197));
 sg13g2_tiehi _18496__198 (.L_HI(net198));
 sg13g2_tiehi _18495__199 (.L_HI(net199));
 sg13g2_tiehi _18494__200 (.L_HI(net200));
 sg13g2_tiehi _18493__201 (.L_HI(net201));
 sg13g2_tiehi _18492__202 (.L_HI(net202));
 sg13g2_tiehi _18491__203 (.L_HI(net203));
 sg13g2_tiehi _18490__204 (.L_HI(net204));
 sg13g2_tiehi _18489__205 (.L_HI(net205));
 sg13g2_tiehi _18488__206 (.L_HI(net206));
 sg13g2_tiehi _18487__207 (.L_HI(net207));
 sg13g2_tiehi _18486__208 (.L_HI(net208));
 sg13g2_tiehi _18485__209 (.L_HI(net209));
 sg13g2_tiehi _18484__210 (.L_HI(net210));
 sg13g2_tiehi _18483__211 (.L_HI(net211));
 sg13g2_tiehi _18482__212 (.L_HI(net212));
 sg13g2_tiehi _18481__213 (.L_HI(net213));
 sg13g2_tiehi _18480__214 (.L_HI(net214));
 sg13g2_tiehi _18479__215 (.L_HI(net215));
 sg13g2_tiehi _18478__216 (.L_HI(net216));
 sg13g2_tiehi _18477__217 (.L_HI(net217));
 sg13g2_tiehi _18476__218 (.L_HI(net218));
 sg13g2_tiehi _18475__219 (.L_HI(net219));
 sg13g2_tiehi _18474__220 (.L_HI(net220));
 sg13g2_tiehi _18473__221 (.L_HI(net221));
 sg13g2_tiehi _18472__222 (.L_HI(net222));
 sg13g2_tiehi _18471__223 (.L_HI(net223));
 sg13g2_tiehi _18470__224 (.L_HI(net224));
 sg13g2_tiehi _18469__225 (.L_HI(net225));
 sg13g2_tiehi _18468__226 (.L_HI(net226));
 sg13g2_tiehi _18467__227 (.L_HI(net227));
 sg13g2_tiehi _18466__228 (.L_HI(net228));
 sg13g2_tiehi _18465__229 (.L_HI(net229));
 sg13g2_tiehi _18464__230 (.L_HI(net230));
 sg13g2_tiehi _18463__231 (.L_HI(net231));
 sg13g2_tiehi _18462__232 (.L_HI(net232));
 sg13g2_tiehi _18461__233 (.L_HI(net233));
 sg13g2_tiehi _18460__234 (.L_HI(net234));
 sg13g2_tiehi _18459__235 (.L_HI(net235));
 sg13g2_tiehi _18458__236 (.L_HI(net236));
 sg13g2_tiehi _18457__237 (.L_HI(net237));
 sg13g2_tiehi _18456__238 (.L_HI(net238));
 sg13g2_tiehi _18455__239 (.L_HI(net239));
 sg13g2_tiehi _18454__240 (.L_HI(net240));
 sg13g2_tiehi _18453__241 (.L_HI(net241));
 sg13g2_tiehi _18452__242 (.L_HI(net242));
 sg13g2_tiehi _18451__243 (.L_HI(net243));
 sg13g2_tiehi _18450__244 (.L_HI(net244));
 sg13g2_tiehi _18449__245 (.L_HI(net245));
 sg13g2_tiehi _18448__246 (.L_HI(net246));
 sg13g2_tiehi _18447__247 (.L_HI(net247));
 sg13g2_tiehi _18446__248 (.L_HI(net248));
 sg13g2_tiehi _18445__249 (.L_HI(net249));
 sg13g2_tiehi _18444__250 (.L_HI(net250));
 sg13g2_tiehi _18443__251 (.L_HI(net251));
 sg13g2_tiehi _18442__252 (.L_HI(net252));
 sg13g2_tiehi _18441__253 (.L_HI(net253));
 sg13g2_tiehi _18440__254 (.L_HI(net254));
 sg13g2_tiehi _18439__255 (.L_HI(net255));
 sg13g2_tiehi _18438__256 (.L_HI(net256));
 sg13g2_tiehi _18437__257 (.L_HI(net257));
 sg13g2_tiehi _18436__258 (.L_HI(net258));
 sg13g2_tiehi _18435__259 (.L_HI(net259));
 sg13g2_tiehi _18434__260 (.L_HI(net260));
 sg13g2_tiehi _18433__261 (.L_HI(net261));
 sg13g2_tiehi _18432__262 (.L_HI(net262));
 sg13g2_tiehi _18431__263 (.L_HI(net263));
 sg13g2_tiehi _18430__264 (.L_HI(net264));
 sg13g2_tiehi _18429__265 (.L_HI(net265));
 sg13g2_tiehi _18428__266 (.L_HI(net266));
 sg13g2_tiehi _18427__267 (.L_HI(net267));
 sg13g2_tiehi _18426__268 (.L_HI(net268));
 sg13g2_tiehi _18425__269 (.L_HI(net269));
 sg13g2_tiehi _18424__270 (.L_HI(net270));
 sg13g2_tiehi _18423__271 (.L_HI(net271));
 sg13g2_tiehi _18422__272 (.L_HI(net272));
 sg13g2_tiehi _18421__273 (.L_HI(net273));
 sg13g2_tiehi _18420__274 (.L_HI(net274));
 sg13g2_tiehi _18419__275 (.L_HI(net275));
 sg13g2_tiehi _18418__276 (.L_HI(net276));
 sg13g2_tiehi _18417__277 (.L_HI(net277));
 sg13g2_tiehi _18416__278 (.L_HI(net278));
 sg13g2_tiehi _18415__279 (.L_HI(net279));
 sg13g2_tiehi _18414__280 (.L_HI(net280));
 sg13g2_tiehi _18413__281 (.L_HI(net281));
 sg13g2_tiehi _18412__282 (.L_HI(net282));
 sg13g2_tiehi _18411__283 (.L_HI(net283));
 sg13g2_tiehi _18410__284 (.L_HI(net284));
 sg13g2_tiehi _18409__285 (.L_HI(net285));
 sg13g2_tiehi _18408__286 (.L_HI(net286));
 sg13g2_tiehi _18407__287 (.L_HI(net287));
 sg13g2_tiehi _18406__288 (.L_HI(net288));
 sg13g2_tiehi _18405__289 (.L_HI(net289));
 sg13g2_tiehi _18404__290 (.L_HI(net290));
 sg13g2_tiehi _18403__291 (.L_HI(net291));
 sg13g2_tiehi _18402__292 (.L_HI(net292));
 sg13g2_tiehi _18401__293 (.L_HI(net293));
 sg13g2_tiehi _18400__294 (.L_HI(net294));
 sg13g2_tiehi _18399__295 (.L_HI(net295));
 sg13g2_tiehi _18398__296 (.L_HI(net296));
 sg13g2_tiehi _18397__297 (.L_HI(net297));
 sg13g2_tiehi _18396__298 (.L_HI(net298));
 sg13g2_tiehi _18395__299 (.L_HI(net299));
 sg13g2_tiehi _18394__300 (.L_HI(net300));
 sg13g2_tiehi _18393__301 (.L_HI(net301));
 sg13g2_tiehi _18392__302 (.L_HI(net302));
 sg13g2_tiehi _18391__303 (.L_HI(net303));
 sg13g2_tiehi _18390__304 (.L_HI(net304));
 sg13g2_tiehi _18389__305 (.L_HI(net305));
 sg13g2_tiehi _18388__306 (.L_HI(net306));
 sg13g2_tiehi _18387__307 (.L_HI(net307));
 sg13g2_tiehi _18386__308 (.L_HI(net308));
 sg13g2_tiehi _18385__309 (.L_HI(net309));
 sg13g2_tiehi _18384__310 (.L_HI(net310));
 sg13g2_tiehi _18383__311 (.L_HI(net311));
 sg13g2_tiehi _18382__312 (.L_HI(net312));
 sg13g2_tiehi _18381__313 (.L_HI(net313));
 sg13g2_tiehi _18380__314 (.L_HI(net314));
 sg13g2_tiehi _18379__315 (.L_HI(net315));
 sg13g2_tiehi _18378__316 (.L_HI(net316));
 sg13g2_tiehi _18377__317 (.L_HI(net317));
 sg13g2_tiehi _18376__318 (.L_HI(net318));
 sg13g2_tiehi _18375__319 (.L_HI(net319));
 sg13g2_tiehi _18374__320 (.L_HI(net320));
 sg13g2_tiehi _19789__321 (.L_HI(net321));
 sg13g2_tiehi _18373__322 (.L_HI(net322));
 sg13g2_tiehi _19788__323 (.L_HI(net323));
 sg13g2_tiehi _18372__324 (.L_HI(net324));
 sg13g2_tiehi _19787__325 (.L_HI(net325));
 sg13g2_tiehi _18371__326 (.L_HI(net326));
 sg13g2_tiehi _19786__327 (.L_HI(net327));
 sg13g2_tiehi _18370__328 (.L_HI(net328));
 sg13g2_tiehi _18369__329 (.L_HI(net329));
 sg13g2_tiehi _18368__330 (.L_HI(net330));
 sg13g2_tiehi _18367__331 (.L_HI(net331));
 sg13g2_tiehi _18366__332 (.L_HI(net332));
 sg13g2_tiehi _18365__333 (.L_HI(net333));
 sg13g2_tiehi _18364__334 (.L_HI(net334));
 sg13g2_tiehi _18363__335 (.L_HI(net335));
 sg13g2_tiehi _18362__336 (.L_HI(net336));
 sg13g2_tiehi _18361__337 (.L_HI(net337));
 sg13g2_tiehi _18360__338 (.L_HI(net338));
 sg13g2_tiehi _18359__339 (.L_HI(net339));
 sg13g2_tiehi _18358__340 (.L_HI(net340));
 sg13g2_tiehi _18357__341 (.L_HI(net341));
 sg13g2_tiehi _18356__342 (.L_HI(net342));
 sg13g2_tiehi _18355__343 (.L_HI(net343));
 sg13g2_tiehi _18354__344 (.L_HI(net344));
 sg13g2_tiehi _18353__345 (.L_HI(net345));
 sg13g2_tiehi _18352__346 (.L_HI(net346));
 sg13g2_tiehi _18351__347 (.L_HI(net347));
 sg13g2_tiehi _18350__348 (.L_HI(net348));
 sg13g2_tiehi _18349__349 (.L_HI(net349));
 sg13g2_tiehi _18348__350 (.L_HI(net350));
 sg13g2_tiehi _18347__351 (.L_HI(net351));
 sg13g2_tiehi _18346__352 (.L_HI(net352));
 sg13g2_tiehi _18345__353 (.L_HI(net353));
 sg13g2_tiehi _18344__354 (.L_HI(net354));
 sg13g2_tiehi _18343__355 (.L_HI(net355));
 sg13g2_tiehi _18342__356 (.L_HI(net356));
 sg13g2_tiehi _18341__357 (.L_HI(net357));
 sg13g2_tiehi _18340__358 (.L_HI(net358));
 sg13g2_tiehi _18339__359 (.L_HI(net359));
 sg13g2_tiehi _18338__360 (.L_HI(net360));
 sg13g2_tiehi _19785__361 (.L_HI(net361));
 sg13g2_tiehi _18337__362 (.L_HI(net362));
 sg13g2_tiehi _19784__363 (.L_HI(net363));
 sg13g2_tiehi _18336__364 (.L_HI(net364));
 sg13g2_tiehi _19783__365 (.L_HI(net365));
 sg13g2_tiehi _18335__366 (.L_HI(net366));
 sg13g2_tiehi _19782__367 (.L_HI(net367));
 sg13g2_tiehi _18334__368 (.L_HI(net368));
 sg13g2_tiehi _19781__369 (.L_HI(net369));
 sg13g2_tiehi _18333__370 (.L_HI(net370));
 sg13g2_tiehi _19780__371 (.L_HI(net371));
 sg13g2_tiehi _18332__372 (.L_HI(net372));
 sg13g2_tiehi _19779__373 (.L_HI(net373));
 sg13g2_tiehi _18331__374 (.L_HI(net374));
 sg13g2_tiehi _19778__375 (.L_HI(net375));
 sg13g2_tiehi _18330__376 (.L_HI(net376));
 sg13g2_tiehi _19777__377 (.L_HI(net377));
 sg13g2_tiehi _18329__378 (.L_HI(net378));
 sg13g2_tiehi _19776__379 (.L_HI(net379));
 sg13g2_tiehi _18328__380 (.L_HI(net380));
 sg13g2_tiehi _19775__381 (.L_HI(net381));
 sg13g2_tiehi _18327__382 (.L_HI(net382));
 sg13g2_tiehi _19774__383 (.L_HI(net383));
 sg13g2_tiehi _18326__384 (.L_HI(net384));
 sg13g2_tiehi _19773__385 (.L_HI(net385));
 sg13g2_tiehi _18325__386 (.L_HI(net386));
 sg13g2_tiehi _19772__387 (.L_HI(net387));
 sg13g2_tiehi _18324__388 (.L_HI(net388));
 sg13g2_tiehi _19771__389 (.L_HI(net389));
 sg13g2_tiehi _18323__390 (.L_HI(net390));
 sg13g2_tiehi _19770__391 (.L_HI(net391));
 sg13g2_tiehi _18322__392 (.L_HI(net392));
 sg13g2_tiehi _19769__393 (.L_HI(net393));
 sg13g2_tiehi _18321__394 (.L_HI(net394));
 sg13g2_tiehi _19768__395 (.L_HI(net395));
 sg13g2_tiehi _18320__396 (.L_HI(net396));
 sg13g2_tiehi _19767__397 (.L_HI(net397));
 sg13g2_tiehi _18319__398 (.L_HI(net398));
 sg13g2_tiehi _19766__399 (.L_HI(net399));
 sg13g2_tiehi _18318__400 (.L_HI(net400));
 sg13g2_tiehi _19765__401 (.L_HI(net401));
 sg13g2_tiehi _18317__402 (.L_HI(net402));
 sg13g2_tiehi _19764__403 (.L_HI(net403));
 sg13g2_tiehi _18316__404 (.L_HI(net404));
 sg13g2_tiehi _19763__405 (.L_HI(net405));
 sg13g2_tiehi _18315__406 (.L_HI(net406));
 sg13g2_tiehi _19762__407 (.L_HI(net407));
 sg13g2_tiehi _18314__408 (.L_HI(net408));
 sg13g2_tiehi _19761__409 (.L_HI(net409));
 sg13g2_tiehi _18313__410 (.L_HI(net410));
 sg13g2_tiehi _19760__411 (.L_HI(net411));
 sg13g2_tiehi _18312__412 (.L_HI(net412));
 sg13g2_tiehi _19759__413 (.L_HI(net413));
 sg13g2_tiehi _18311__414 (.L_HI(net414));
 sg13g2_tiehi _19758__415 (.L_HI(net415));
 sg13g2_tiehi _18310__416 (.L_HI(net416));
 sg13g2_tiehi _19757__417 (.L_HI(net417));
 sg13g2_tiehi _18309__418 (.L_HI(net418));
 sg13g2_tiehi _19756__419 (.L_HI(net419));
 sg13g2_tiehi _18308__420 (.L_HI(net420));
 sg13g2_tiehi _19755__421 (.L_HI(net421));
 sg13g2_tiehi _18307__422 (.L_HI(net422));
 sg13g2_tiehi _18306__423 (.L_HI(net423));
 sg13g2_tiehi _18305__424 (.L_HI(net424));
 sg13g2_tiehi _18304__425 (.L_HI(net425));
 sg13g2_tiehi _18303__426 (.L_HI(net426));
 sg13g2_tiehi _18302__427 (.L_HI(net427));
 sg13g2_tiehi _18301__428 (.L_HI(net428));
 sg13g2_tiehi _18300__429 (.L_HI(net429));
 sg13g2_tiehi _18299__430 (.L_HI(net430));
 sg13g2_tiehi _19754__431 (.L_HI(net431));
 sg13g2_tiehi _18298__432 (.L_HI(net432));
 sg13g2_tiehi _19753__433 (.L_HI(net433));
 sg13g2_tiehi _18297__434 (.L_HI(net434));
 sg13g2_tiehi _18296__435 (.L_HI(net435));
 sg13g2_tiehi _18295__436 (.L_HI(net436));
 sg13g2_tiehi _18294__437 (.L_HI(net437));
 sg13g2_tiehi _18293__438 (.L_HI(net438));
 sg13g2_tiehi _18292__439 (.L_HI(net439));
 sg13g2_tiehi _18291__440 (.L_HI(net440));
 sg13g2_tiehi _18290__441 (.L_HI(net441));
 sg13g2_tiehi _19752__442 (.L_HI(net442));
 sg13g2_tiehi _19751__443 (.L_HI(net443));
 sg13g2_tiehi _19750__444 (.L_HI(net444));
 sg13g2_tiehi _19749__445 (.L_HI(net445));
 sg13g2_tiehi _19748__446 (.L_HI(net446));
 sg13g2_tiehi _19747__447 (.L_HI(net447));
 sg13g2_tiehi _19746__448 (.L_HI(net448));
 sg13g2_tiehi _19745__449 (.L_HI(net449));
 sg13g2_tiehi _19744__450 (.L_HI(net450));
 sg13g2_tiehi _19743__451 (.L_HI(net451));
 sg13g2_tiehi _19742__452 (.L_HI(net452));
 sg13g2_tiehi _19741__453 (.L_HI(net453));
 sg13g2_tiehi _19740__454 (.L_HI(net454));
 sg13g2_tiehi _19739__455 (.L_HI(net455));
 sg13g2_tiehi _19738__456 (.L_HI(net456));
 sg13g2_tiehi _19737__457 (.L_HI(net457));
 sg13g2_tiehi _19736__458 (.L_HI(net458));
 sg13g2_tiehi _19735__459 (.L_HI(net459));
 sg13g2_tiehi _19734__460 (.L_HI(net460));
 sg13g2_tiehi _19733__461 (.L_HI(net461));
 sg13g2_tiehi _19732__462 (.L_HI(net462));
 sg13g2_tiehi _19731__463 (.L_HI(net463));
 sg13g2_tiehi _19730__464 (.L_HI(net464));
 sg13g2_tiehi _19729__465 (.L_HI(net465));
 sg13g2_tiehi _19728__466 (.L_HI(net466));
 sg13g2_tiehi _19727__467 (.L_HI(net467));
 sg13g2_tiehi _19726__468 (.L_HI(net468));
 sg13g2_tiehi _19725__469 (.L_HI(net469));
 sg13g2_tiehi _19724__470 (.L_HI(net470));
 sg13g2_tiehi _19723__471 (.L_HI(net471));
 sg13g2_tiehi _19722__472 (.L_HI(net472));
 sg13g2_tiehi _19721__473 (.L_HI(net473));
 sg13g2_tiehi _19720__474 (.L_HI(net474));
 sg13g2_tiehi _19719__475 (.L_HI(net475));
 sg13g2_tiehi _19718__476 (.L_HI(net476));
 sg13g2_tiehi _19717__477 (.L_HI(net477));
 sg13g2_tiehi _19716__478 (.L_HI(net478));
 sg13g2_tiehi _19715__479 (.L_HI(net479));
 sg13g2_tiehi _19714__480 (.L_HI(net480));
 sg13g2_tiehi _19713__481 (.L_HI(net481));
 sg13g2_tiehi _19712__482 (.L_HI(net482));
 sg13g2_tiehi _19711__483 (.L_HI(net483));
 sg13g2_tiehi _19710__484 (.L_HI(net484));
 sg13g2_tiehi _19709__485 (.L_HI(net485));
 sg13g2_tiehi _19708__486 (.L_HI(net486));
 sg13g2_tiehi _19707__487 (.L_HI(net487));
 sg13g2_tiehi _19706__488 (.L_HI(net488));
 sg13g2_tiehi _19705__489 (.L_HI(net489));
 sg13g2_tiehi _19704__490 (.L_HI(net490));
 sg13g2_tiehi _19703__491 (.L_HI(net491));
 sg13g2_tiehi _19702__492 (.L_HI(net492));
 sg13g2_tiehi _19701__493 (.L_HI(net493));
 sg13g2_tiehi _19700__494 (.L_HI(net494));
 sg13g2_tiehi _19699__495 (.L_HI(net495));
 sg13g2_tiehi _19698__496 (.L_HI(net496));
 sg13g2_tiehi _19697__497 (.L_HI(net497));
 sg13g2_tiehi _19696__498 (.L_HI(net498));
 sg13g2_tiehi _19695__499 (.L_HI(net499));
 sg13g2_tiehi _19694__500 (.L_HI(net500));
 sg13g2_tiehi _19693__501 (.L_HI(net501));
 sg13g2_tiehi _19692__502 (.L_HI(net502));
 sg13g2_tiehi _19691__503 (.L_HI(net503));
 sg13g2_tiehi _19690__504 (.L_HI(net504));
 sg13g2_tiehi _19689__505 (.L_HI(net505));
 sg13g2_tiehi _19688__506 (.L_HI(net506));
 sg13g2_tiehi _19687__507 (.L_HI(net507));
 sg13g2_tiehi _19686__508 (.L_HI(net508));
 sg13g2_tiehi _19685__509 (.L_HI(net509));
 sg13g2_tiehi _19684__510 (.L_HI(net510));
 sg13g2_tiehi _19683__511 (.L_HI(net511));
 sg13g2_tiehi _19682__512 (.L_HI(net512));
 sg13g2_tiehi _19681__513 (.L_HI(net513));
 sg13g2_tiehi _19680__514 (.L_HI(net514));
 sg13g2_tiehi _19679__515 (.L_HI(net515));
 sg13g2_tiehi _19678__516 (.L_HI(net516));
 sg13g2_tiehi _19677__517 (.L_HI(net517));
 sg13g2_tiehi _19676__518 (.L_HI(net518));
 sg13g2_tiehi _19675__519 (.L_HI(net519));
 sg13g2_tiehi _19674__520 (.L_HI(net520));
 sg13g2_tiehi _19673__521 (.L_HI(net521));
 sg13g2_tiehi _19672__522 (.L_HI(net522));
 sg13g2_tiehi _19671__523 (.L_HI(net523));
 sg13g2_tiehi _19670__524 (.L_HI(net524));
 sg13g2_tiehi _19669__525 (.L_HI(net525));
 sg13g2_tiehi _19668__526 (.L_HI(net526));
 sg13g2_tiehi _19667__527 (.L_HI(net527));
 sg13g2_tiehi _19666__528 (.L_HI(net528));
 sg13g2_tiehi _19665__529 (.L_HI(net529));
 sg13g2_tiehi _19664__530 (.L_HI(net530));
 sg13g2_tiehi _19663__531 (.L_HI(net531));
 sg13g2_tiehi _19662__532 (.L_HI(net532));
 sg13g2_tiehi _19661__533 (.L_HI(net533));
 sg13g2_tiehi _19660__534 (.L_HI(net534));
 sg13g2_tiehi _19659__535 (.L_HI(net535));
 sg13g2_tiehi _19658__536 (.L_HI(net536));
 sg13g2_tiehi _19657__537 (.L_HI(net537));
 sg13g2_tiehi _19656__538 (.L_HI(net538));
 sg13g2_tiehi _19655__539 (.L_HI(net539));
 sg13g2_tiehi _19654__540 (.L_HI(net540));
 sg13g2_tiehi _19653__541 (.L_HI(net541));
 sg13g2_tiehi _19652__542 (.L_HI(net542));
 sg13g2_tiehi _19651__543 (.L_HI(net543));
 sg13g2_tiehi _19650__544 (.L_HI(net544));
 sg13g2_tiehi _19649__545 (.L_HI(net545));
 sg13g2_tiehi _19648__546 (.L_HI(net546));
 sg13g2_tiehi _19647__547 (.L_HI(net547));
 sg13g2_tiehi _19646__548 (.L_HI(net548));
 sg13g2_tiehi _19645__549 (.L_HI(net549));
 sg13g2_tiehi _19644__550 (.L_HI(net550));
 sg13g2_tiehi _19643__551 (.L_HI(net551));
 sg13g2_tiehi _19642__552 (.L_HI(net552));
 sg13g2_tiehi _19641__553 (.L_HI(net553));
 sg13g2_tiehi _19640__554 (.L_HI(net554));
 sg13g2_tiehi _19639__555 (.L_HI(net555));
 sg13g2_tiehi _19638__556 (.L_HI(net556));
 sg13g2_tiehi _19637__557 (.L_HI(net557));
 sg13g2_tiehi _19636__558 (.L_HI(net558));
 sg13g2_tiehi _19635__559 (.L_HI(net559));
 sg13g2_tiehi _19634__560 (.L_HI(net560));
 sg13g2_tiehi _19633__561 (.L_HI(net561));
 sg13g2_tiehi _19632__562 (.L_HI(net562));
 sg13g2_tiehi _19631__563 (.L_HI(net563));
 sg13g2_tiehi _19630__564 (.L_HI(net564));
 sg13g2_tiehi _19629__565 (.L_HI(net565));
 sg13g2_tiehi _19628__566 (.L_HI(net566));
 sg13g2_tiehi _19627__567 (.L_HI(net567));
 sg13g2_tiehi _19626__568 (.L_HI(net568));
 sg13g2_tiehi _19625__569 (.L_HI(net569));
 sg13g2_tiehi _19624__570 (.L_HI(net570));
 sg13g2_tiehi _19623__571 (.L_HI(net571));
 sg13g2_tiehi _19622__572 (.L_HI(net572));
 sg13g2_tiehi _19621__573 (.L_HI(net573));
 sg13g2_tiehi _19620__574 (.L_HI(net574));
 sg13g2_tiehi _19619__575 (.L_HI(net575));
 sg13g2_tiehi _19618__576 (.L_HI(net576));
 sg13g2_tiehi _19617__577 (.L_HI(net577));
 sg13g2_tiehi _19616__578 (.L_HI(net578));
 sg13g2_tiehi _19615__579 (.L_HI(net579));
 sg13g2_tiehi _19614__580 (.L_HI(net580));
 sg13g2_tiehi _19613__581 (.L_HI(net581));
 sg13g2_tiehi _19612__582 (.L_HI(net582));
 sg13g2_tiehi _19611__583 (.L_HI(net583));
 sg13g2_tiehi _19610__584 (.L_HI(net584));
 sg13g2_tiehi _19609__585 (.L_HI(net585));
 sg13g2_tiehi _19608__586 (.L_HI(net586));
 sg13g2_tiehi _19607__587 (.L_HI(net587));
 sg13g2_tiehi _19606__588 (.L_HI(net588));
 sg13g2_tiehi _19605__589 (.L_HI(net589));
 sg13g2_tiehi _19604__590 (.L_HI(net590));
 sg13g2_tiehi _19603__591 (.L_HI(net591));
 sg13g2_tiehi _19602__592 (.L_HI(net592));
 sg13g2_tiehi _19601__593 (.L_HI(net593));
 sg13g2_tiehi _19600__594 (.L_HI(net594));
 sg13g2_tiehi _19599__595 (.L_HI(net595));
 sg13g2_tiehi _19598__596 (.L_HI(net596));
 sg13g2_tiehi _19597__597 (.L_HI(net597));
 sg13g2_tiehi _19596__598 (.L_HI(net598));
 sg13g2_tiehi _19595__599 (.L_HI(net599));
 sg13g2_tiehi _19594__600 (.L_HI(net600));
 sg13g2_tiehi _19593__601 (.L_HI(net601));
 sg13g2_tiehi _19592__602 (.L_HI(net602));
 sg13g2_tiehi _19591__603 (.L_HI(net603));
 sg13g2_tiehi _19590__604 (.L_HI(net604));
 sg13g2_tiehi _19589__605 (.L_HI(net605));
 sg13g2_tiehi _19588__606 (.L_HI(net606));
 sg13g2_tiehi _19587__607 (.L_HI(net607));
 sg13g2_tiehi _19586__608 (.L_HI(net608));
 sg13g2_tiehi _19585__609 (.L_HI(net609));
 sg13g2_tiehi _19584__610 (.L_HI(net610));
 sg13g2_tiehi _19583__611 (.L_HI(net611));
 sg13g2_tiehi _19582__612 (.L_HI(net612));
 sg13g2_tiehi _19581__613 (.L_HI(net613));
 sg13g2_tiehi _19580__614 (.L_HI(net614));
 sg13g2_tiehi _19579__615 (.L_HI(net615));
 sg13g2_tiehi _19578__616 (.L_HI(net616));
 sg13g2_tiehi _19577__617 (.L_HI(net617));
 sg13g2_tiehi _19576__618 (.L_HI(net618));
 sg13g2_tiehi _19575__619 (.L_HI(net619));
 sg13g2_tiehi _19574__620 (.L_HI(net620));
 sg13g2_tiehi _19573__621 (.L_HI(net621));
 sg13g2_tiehi _19572__622 (.L_HI(net622));
 sg13g2_tiehi _19571__623 (.L_HI(net623));
 sg13g2_tiehi _19570__624 (.L_HI(net624));
 sg13g2_tiehi _19569__625 (.L_HI(net625));
 sg13g2_tiehi _19568__626 (.L_HI(net626));
 sg13g2_tiehi _19567__627 (.L_HI(net627));
 sg13g2_tiehi _19566__628 (.L_HI(net628));
 sg13g2_tiehi _19565__629 (.L_HI(net629));
 sg13g2_tiehi _19564__630 (.L_HI(net630));
 sg13g2_tiehi _19563__631 (.L_HI(net631));
 sg13g2_tiehi _19562__632 (.L_HI(net632));
 sg13g2_tiehi _19561__633 (.L_HI(net633));
 sg13g2_tiehi _19560__634 (.L_HI(net634));
 sg13g2_tiehi _19559__635 (.L_HI(net635));
 sg13g2_tiehi _19558__636 (.L_HI(net636));
 sg13g2_tiehi _19557__637 (.L_HI(net637));
 sg13g2_tiehi _19556__638 (.L_HI(net638));
 sg13g2_tiehi _19555__639 (.L_HI(net639));
 sg13g2_tiehi _19554__640 (.L_HI(net640));
 sg13g2_tiehi _19553__641 (.L_HI(net641));
 sg13g2_tiehi _19552__642 (.L_HI(net642));
 sg13g2_tiehi _19551__643 (.L_HI(net643));
 sg13g2_tiehi _19550__644 (.L_HI(net644));
 sg13g2_tiehi _19412__645 (.L_HI(net645));
 sg13g2_tiehi _19549__646 (.L_HI(net646));
 sg13g2_tiehi _19925__647 (.L_HI(net647));
 sg13g2_tiehi _19548__648 (.L_HI(net648));
 sg13g2_tiehi _19547__649 (.L_HI(net649));
 sg13g2_tiehi _19546__650 (.L_HI(net650));
 sg13g2_tiehi _19924__651 (.L_HI(net651));
 sg13g2_tiehi _19545__652 (.L_HI(net652));
 sg13g2_tiehi _19923__653 (.L_HI(net653));
 sg13g2_tiehi _19544__654 (.L_HI(net654));
 sg13g2_tiehi _19922__655 (.L_HI(net655));
 sg13g2_tiehi _19543__656 (.L_HI(net656));
 sg13g2_tiehi _19921__657 (.L_HI(net657));
 sg13g2_tiehi _19542__658 (.L_HI(net658));
 sg13g2_tiehi _19541__659 (.L_HI(net659));
 sg13g2_tiehi _19540__660 (.L_HI(net660));
 sg13g2_tiehi _19539__661 (.L_HI(net661));
 sg13g2_tiehi _19538__662 (.L_HI(net662));
 sg13g2_tiehi _19537__663 (.L_HI(net663));
 sg13g2_tiehi _19536__664 (.L_HI(net664));
 sg13g2_tiehi _19535__665 (.L_HI(net665));
 sg13g2_tiehi _19534__666 (.L_HI(net666));
 sg13g2_tiehi _19533__667 (.L_HI(net667));
 sg13g2_tiehi _19532__668 (.L_HI(net668));
 sg13g2_tiehi _19531__669 (.L_HI(net669));
 sg13g2_tiehi _19530__670 (.L_HI(net670));
 sg13g2_tiehi _19529__671 (.L_HI(net671));
 sg13g2_tiehi _19528__672 (.L_HI(net672));
 sg13g2_tiehi _19527__673 (.L_HI(net673));
 sg13g2_tiehi _19526__674 (.L_HI(net674));
 sg13g2_tiehi _19525__675 (.L_HI(net675));
 sg13g2_tiehi _19524__676 (.L_HI(net676));
 sg13g2_tiehi _19523__677 (.L_HI(net677));
 sg13g2_tiehi _19522__678 (.L_HI(net678));
 sg13g2_tiehi _19521__679 (.L_HI(net679));
 sg13g2_tiehi _19520__680 (.L_HI(net680));
 sg13g2_tiehi _19519__681 (.L_HI(net681));
 sg13g2_tiehi _19518__682 (.L_HI(net682));
 sg13g2_tiehi _19517__683 (.L_HI(net683));
 sg13g2_tiehi _19516__684 (.L_HI(net684));
 sg13g2_tiehi _19515__685 (.L_HI(net685));
 sg13g2_tiehi _19514__686 (.L_HI(net686));
 sg13g2_tiehi _19513__687 (.L_HI(net687));
 sg13g2_tiehi _19512__688 (.L_HI(net688));
 sg13g2_tiehi _19511__689 (.L_HI(net689));
 sg13g2_tiehi _19510__690 (.L_HI(net690));
 sg13g2_tiehi _19920__691 (.L_HI(net691));
 sg13g2_tiehi _19509__692 (.L_HI(net692));
 sg13g2_tiehi _19919__693 (.L_HI(net693));
 sg13g2_tiehi _19508__694 (.L_HI(net694));
 sg13g2_tiehi _19918__695 (.L_HI(net695));
 sg13g2_tiehi _19507__696 (.L_HI(net696));
 sg13g2_tiehi _19917__697 (.L_HI(net697));
 sg13g2_tiehi _19506__698 (.L_HI(net698));
 sg13g2_tiehi _19916__699 (.L_HI(net699));
 sg13g2_tiehi _19505__700 (.L_HI(net700));
 sg13g2_tiehi _19915__701 (.L_HI(net701));
 sg13g2_tiehi _19504__702 (.L_HI(net702));
 sg13g2_tiehi _19914__703 (.L_HI(net703));
 sg13g2_tiehi _19503__704 (.L_HI(net704));
 sg13g2_tiehi _19913__705 (.L_HI(net705));
 sg13g2_tiehi _19502__706 (.L_HI(net706));
 sg13g2_tiehi _19912__707 (.L_HI(net707));
 sg13g2_tiehi _19501__708 (.L_HI(net708));
 sg13g2_tiehi _19911__709 (.L_HI(net709));
 sg13g2_tiehi _19500__710 (.L_HI(net710));
 sg13g2_tiehi _19910__711 (.L_HI(net711));
 sg13g2_tiehi _19499__712 (.L_HI(net712));
 sg13g2_tiehi _19909__713 (.L_HI(net713));
 sg13g2_tiehi _19498__714 (.L_HI(net714));
 sg13g2_tiehi _19908__715 (.L_HI(net715));
 sg13g2_tiehi _19497__716 (.L_HI(net716));
 sg13g2_tiehi _19907__717 (.L_HI(net717));
 sg13g2_tiehi _19496__718 (.L_HI(net718));
 sg13g2_tiehi _19906__719 (.L_HI(net719));
 sg13g2_tiehi _19495__720 (.L_HI(net720));
 sg13g2_tiehi _19905__721 (.L_HI(net721));
 sg13g2_tiehi _19494__722 (.L_HI(net722));
 sg13g2_tiehi _19493__723 (.L_HI(net723));
 sg13g2_tiehi _19492__724 (.L_HI(net724));
 sg13g2_tiehi _19491__725 (.L_HI(net725));
 sg13g2_tiehi _19490__726 (.L_HI(net726));
 sg13g2_tiehi _19489__727 (.L_HI(net727));
 sg13g2_tiehi _19488__728 (.L_HI(net728));
 sg13g2_tiehi _19487__729 (.L_HI(net729));
 sg13g2_tiehi _19486__730 (.L_HI(net730));
 sg13g2_tiehi _19485__731 (.L_HI(net731));
 sg13g2_tiehi _19484__732 (.L_HI(net732));
 sg13g2_tiehi _19483__733 (.L_HI(net733));
 sg13g2_tiehi _19482__734 (.L_HI(net734));
 sg13g2_tiehi _19481__735 (.L_HI(net735));
 sg13g2_tiehi _19480__736 (.L_HI(net736));
 sg13g2_tiehi _19479__737 (.L_HI(net737));
 sg13g2_tiehi _19478__738 (.L_HI(net738));
 sg13g2_tiehi _19477__739 (.L_HI(net739));
 sg13g2_tiehi _19476__740 (.L_HI(net740));
 sg13g2_tiehi _19475__741 (.L_HI(net741));
 sg13g2_tiehi _19474__742 (.L_HI(net742));
 sg13g2_tiehi _19473__743 (.L_HI(net743));
 sg13g2_tiehi _19472__744 (.L_HI(net744));
 sg13g2_tiehi _19471__745 (.L_HI(net745));
 sg13g2_tiehi _19470__746 (.L_HI(net746));
 sg13g2_tiehi _19469__747 (.L_HI(net747));
 sg13g2_tiehi _19468__748 (.L_HI(net748));
 sg13g2_tiehi _19467__749 (.L_HI(net749));
 sg13g2_tiehi _19466__750 (.L_HI(net750));
 sg13g2_tiehi _19465__751 (.L_HI(net751));
 sg13g2_tiehi _19464__752 (.L_HI(net752));
 sg13g2_tiehi _19463__753 (.L_HI(net753));
 sg13g2_tiehi _19462__754 (.L_HI(net754));
 sg13g2_tiehi _19904__755 (.L_HI(net755));
 sg13g2_tiehi _19461__756 (.L_HI(net756));
 sg13g2_tiehi _19903__757 (.L_HI(net757));
 sg13g2_tiehi _19460__758 (.L_HI(net758));
 sg13g2_tiehi _19902__759 (.L_HI(net759));
 sg13g2_tiehi _19459__760 (.L_HI(net760));
 sg13g2_tiehi _19901__761 (.L_HI(net761));
 sg13g2_tiehi _19458__762 (.L_HI(net762));
 sg13g2_tiehi _19900__763 (.L_HI(net763));
 sg13g2_tiehi _19457__764 (.L_HI(net764));
 sg13g2_tiehi _19899__765 (.L_HI(net765));
 sg13g2_tiehi _19456__766 (.L_HI(net766));
 sg13g2_tiehi _19898__767 (.L_HI(net767));
 sg13g2_tiehi _19455__768 (.L_HI(net768));
 sg13g2_tiehi _19897__769 (.L_HI(net769));
 sg13g2_tiehi _19454__770 (.L_HI(net770));
 sg13g2_tiehi _19453__771 (.L_HI(net771));
 sg13g2_tiehi _19452__772 (.L_HI(net772));
 sg13g2_tiehi _19451__773 (.L_HI(net773));
 sg13g2_tiehi _19450__774 (.L_HI(net774));
 sg13g2_tiehi _19449__775 (.L_HI(net775));
 sg13g2_tiehi _19448__776 (.L_HI(net776));
 sg13g2_tiehi _19447__777 (.L_HI(net777));
 sg13g2_tiehi _19446__778 (.L_HI(net778));
 sg13g2_tiehi _19445__779 (.L_HI(net779));
 sg13g2_tiehi _19444__780 (.L_HI(net780));
 sg13g2_tiehi _19443__781 (.L_HI(net781));
 sg13g2_tiehi _19442__782 (.L_HI(net782));
 sg13g2_tiehi _19441__783 (.L_HI(net783));
 sg13g2_tiehi _19440__784 (.L_HI(net784));
 sg13g2_tiehi _19439__785 (.L_HI(net785));
 sg13g2_tiehi _19438__786 (.L_HI(net786));
 sg13g2_tiehi _19437__787 (.L_HI(net787));
 sg13g2_tiehi _19436__788 (.L_HI(net788));
 sg13g2_tiehi _19435__789 (.L_HI(net789));
 sg13g2_tiehi _19434__790 (.L_HI(net790));
 sg13g2_tiehi _19433__791 (.L_HI(net791));
 sg13g2_tiehi _19432__792 (.L_HI(net792));
 sg13g2_tiehi _19431__793 (.L_HI(net793));
 sg13g2_tiehi _19430__794 (.L_HI(net794));
 sg13g2_tiehi _19429__795 (.L_HI(net795));
 sg13g2_tiehi _19428__796 (.L_HI(net796));
 sg13g2_tiehi _19427__797 (.L_HI(net797));
 sg13g2_tiehi _19426__798 (.L_HI(net798));
 sg13g2_tiehi _19425__799 (.L_HI(net799));
 sg13g2_tiehi _19424__800 (.L_HI(net800));
 sg13g2_tiehi _19423__801 (.L_HI(net801));
 sg13g2_tiehi _19422__802 (.L_HI(net802));
 sg13g2_tiehi _19896__803 (.L_HI(net803));
 sg13g2_tiehi _19421__804 (.L_HI(net804));
 sg13g2_tiehi _19895__805 (.L_HI(net805));
 sg13g2_tiehi _19420__806 (.L_HI(net806));
 sg13g2_tiehi _19894__807 (.L_HI(net807));
 sg13g2_tiehi _19419__808 (.L_HI(net808));
 sg13g2_tiehi _19893__809 (.L_HI(net809));
 sg13g2_tiehi _19418__810 (.L_HI(net810));
 sg13g2_tiehi _19892__811 (.L_HI(net811));
 sg13g2_tiehi _19417__812 (.L_HI(net812));
 sg13g2_tiehi _19891__813 (.L_HI(net813));
 sg13g2_tiehi _19416__814 (.L_HI(net814));
 sg13g2_tiehi _19890__815 (.L_HI(net815));
 sg13g2_tiehi _19415__816 (.L_HI(net816));
 sg13g2_tiehi _19889__817 (.L_HI(net817));
 sg13g2_tiehi _19414__818 (.L_HI(net818));
 sg13g2_tiehi _19413__819 (.L_HI(net819));
 sg13g2_tiehi _19404__820 (.L_HI(net820));
 sg13g2_tiehi _19403__821 (.L_HI(net821));
 sg13g2_tiehi _19402__822 (.L_HI(net822));
 sg13g2_tiehi _19401__823 (.L_HI(net823));
 sg13g2_tiehi _19400__824 (.L_HI(net824));
 sg13g2_tiehi _19399__825 (.L_HI(net825));
 sg13g2_tiehi _19398__826 (.L_HI(net826));
 sg13g2_tiehi _19397__827 (.L_HI(net827));
 sg13g2_tiehi _19380__828 (.L_HI(net828));
 sg13g2_tiehi _19379__829 (.L_HI(net829));
 sg13g2_tiehi _19378__830 (.L_HI(net830));
 sg13g2_tiehi _19377__831 (.L_HI(net831));
 sg13g2_tiehi _19376__832 (.L_HI(net832));
 sg13g2_tiehi _19375__833 (.L_HI(net833));
 sg13g2_tiehi _19374__834 (.L_HI(net834));
 sg13g2_tiehi _19373__835 (.L_HI(net835));
 sg13g2_tiehi _19888__836 (.L_HI(net836));
 sg13g2_tiehi _19372__837 (.L_HI(net837));
 sg13g2_tiehi _19887__838 (.L_HI(net838));
 sg13g2_tiehi _19371__839 (.L_HI(net839));
 sg13g2_tiehi _19886__840 (.L_HI(net840));
 sg13g2_tiehi _19370__841 (.L_HI(net841));
 sg13g2_tiehi _19369__842 (.L_HI(net842));
 sg13g2_tiehi _19368__843 (.L_HI(net843));
 sg13g2_tiehi _19367__844 (.L_HI(net844));
 sg13g2_tiehi _19366__845 (.L_HI(net845));
 sg13g2_tiehi _19365__846 (.L_HI(net846));
 sg13g2_tiehi _19364__847 (.L_HI(net847));
 sg13g2_tiehi _19363__848 (.L_HI(net848));
 sg13g2_tiehi _19362__849 (.L_HI(net849));
 sg13g2_tiehi _19361__850 (.L_HI(net850));
 sg13g2_tiehi _19360__851 (.L_HI(net851));
 sg13g2_tiehi _19359__852 (.L_HI(net852));
 sg13g2_tiehi _19358__853 (.L_HI(net853));
 sg13g2_tiehi _19357__854 (.L_HI(net854));
 sg13g2_tiehi _19356__855 (.L_HI(net855));
 sg13g2_tiehi _19355__856 (.L_HI(net856));
 sg13g2_tiehi _19354__857 (.L_HI(net857));
 sg13g2_tiehi _19353__858 (.L_HI(net858));
 sg13g2_tiehi _19336__859 (.L_HI(net859));
 sg13g2_tiehi _19335__860 (.L_HI(net860));
 sg13g2_tiehi _19334__861 (.L_HI(net861));
 sg13g2_tiehi _19333__862 (.L_HI(net862));
 sg13g2_tiehi _19332__863 (.L_HI(net863));
 sg13g2_tiehi _19331__864 (.L_HI(net864));
 sg13g2_tiehi _19330__865 (.L_HI(net865));
 sg13g2_tiehi _19329__866 (.L_HI(net866));
 sg13g2_tiehi _19328__867 (.L_HI(net867));
 sg13g2_tiehi _19327__868 (.L_HI(net868));
 sg13g2_tiehi _19326__869 (.L_HI(net869));
 sg13g2_tiehi _19325__870 (.L_HI(net870));
 sg13g2_tiehi _19324__871 (.L_HI(net871));
 sg13g2_tiehi _19323__872 (.L_HI(net872));
 sg13g2_tiehi _19322__873 (.L_HI(net873));
 sg13g2_tiehi _19321__874 (.L_HI(net874));
 sg13g2_tiehi _19320__875 (.L_HI(net875));
 sg13g2_tiehi _19319__876 (.L_HI(net876));
 sg13g2_tiehi _19318__877 (.L_HI(net877));
 sg13g2_tiehi _19317__878 (.L_HI(net878));
 sg13g2_tiehi _19316__879 (.L_HI(net879));
 sg13g2_tiehi _19885__880 (.L_HI(net880));
 sg13g2_tiehi _19315__881 (.L_HI(net881));
 sg13g2_tiehi _19884__882 (.L_HI(net882));
 sg13g2_tiehi _19314__883 (.L_HI(net883));
 sg13g2_tiehi _19883__884 (.L_HI(net884));
 sg13g2_tiehi _19313__885 (.L_HI(net885));
 sg13g2_tiehi _19882__886 (.L_HI(net886));
 sg13g2_tiehi _19312__887 (.L_HI(net887));
 sg13g2_tiehi _19881__888 (.L_HI(net888));
 sg13g2_tiehi _19311__889 (.L_HI(net889));
 sg13g2_tiehi _19880__890 (.L_HI(net890));
 sg13g2_tiehi _19310__891 (.L_HI(net891));
 sg13g2_tiehi _19879__892 (.L_HI(net892));
 sg13g2_tiehi _19309__893 (.L_HI(net893));
 sg13g2_tiehi _19878__894 (.L_HI(net894));
 sg13g2_tiehi _19308__895 (.L_HI(net895));
 sg13g2_tiehi _19877__896 (.L_HI(net896));
 sg13g2_tiehi _19307__897 (.L_HI(net897));
 sg13g2_tiehi _19876__898 (.L_HI(net898));
 sg13g2_tiehi _19306__899 (.L_HI(net899));
 sg13g2_tiehi _19875__900 (.L_HI(net900));
 sg13g2_tiehi _19305__901 (.L_HI(net901));
 sg13g2_tiehi _19304__902 (.L_HI(net902));
 sg13g2_tiehi _19303__903 (.L_HI(net903));
 sg13g2_tiehi _19302__904 (.L_HI(net904));
 sg13g2_tiehi _19301__905 (.L_HI(net905));
 sg13g2_tiehi _19300__906 (.L_HI(net906));
 sg13g2_tiehi _19299__907 (.L_HI(net907));
 sg13g2_tiehi _19298__908 (.L_HI(net908));
 sg13g2_tiehi _19297__909 (.L_HI(net909));
 sg13g2_tiehi _19296__910 (.L_HI(net910));
 sg13g2_tiehi _19874__911 (.L_HI(net911));
 sg13g2_tiehi _19295__912 (.L_HI(net912));
 sg13g2_tiehi _19873__913 (.L_HI(net913));
 sg13g2_tiehi _19294__914 (.L_HI(net914));
 sg13g2_tiehi _19872__915 (.L_HI(net915));
 sg13g2_tiehi _19293__916 (.L_HI(net916));
 sg13g2_tiehi _19871__917 (.L_HI(net917));
 sg13g2_tiehi _19292__918 (.L_HI(net918));
 sg13g2_tiehi _19870__919 (.L_HI(net919));
 sg13g2_tiehi _19291__920 (.L_HI(net920));
 sg13g2_tiehi _19869__921 (.L_HI(net921));
 sg13g2_tiehi _19290__922 (.L_HI(net922));
 sg13g2_tiehi _19868__923 (.L_HI(net923));
 sg13g2_tiehi _19289__924 (.L_HI(net924));
 sg13g2_tiehi _19867__925 (.L_HI(net925));
 sg13g2_tiehi _19288__926 (.L_HI(net926));
 sg13g2_tiehi _19866__927 (.L_HI(net927));
 sg13g2_tiehi _19287__928 (.L_HI(net928));
 sg13g2_tiehi _19865__929 (.L_HI(net929));
 sg13g2_tiehi _19286__930 (.L_HI(net930));
 sg13g2_tiehi _19864__931 (.L_HI(net931));
 sg13g2_tiehi _19285__932 (.L_HI(net932));
 sg13g2_tiehi _19863__933 (.L_HI(net933));
 sg13g2_tiehi _19284__934 (.L_HI(net934));
 sg13g2_tiehi _19862__935 (.L_HI(net935));
 sg13g2_tiehi _19283__936 (.L_HI(net936));
 sg13g2_tiehi _19861__937 (.L_HI(net937));
 sg13g2_tiehi _19282__938 (.L_HI(net938));
 sg13g2_tiehi _19860__939 (.L_HI(net939));
 sg13g2_tiehi _19281__940 (.L_HI(net940));
 sg13g2_tiehi _19859__941 (.L_HI(net941));
 sg13g2_tiehi _19280__942 (.L_HI(net942));
 sg13g2_tiehi _19279__943 (.L_HI(net943));
 sg13g2_tiehi _19278__944 (.L_HI(net944));
 sg13g2_tiehi _19277__945 (.L_HI(net945));
 sg13g2_tiehi _19276__946 (.L_HI(net946));
 sg13g2_tiehi _19275__947 (.L_HI(net947));
 sg13g2_tiehi _19274__948 (.L_HI(net948));
 sg13g2_tiehi _19273__949 (.L_HI(net949));
 sg13g2_tiehi _19272__950 (.L_HI(net950));
 sg13g2_tiehi _19858__951 (.L_HI(net951));
 sg13g2_tiehi _19271__952 (.L_HI(net952));
 sg13g2_tiehi _19857__953 (.L_HI(net953));
 sg13g2_tiehi _19270__954 (.L_HI(net954));
 sg13g2_tiehi _19856__955 (.L_HI(net955));
 sg13g2_tiehi _19269__956 (.L_HI(net956));
 sg13g2_tiehi _19855__957 (.L_HI(net957));
 sg13g2_tiehi _19268__958 (.L_HI(net958));
 sg13g2_tiehi _19854__959 (.L_HI(net959));
 sg13g2_tiehi _19267__960 (.L_HI(net960));
 sg13g2_tiehi _19853__961 (.L_HI(net961));
 sg13g2_tiehi _19266__962 (.L_HI(net962));
 sg13g2_tiehi _19852__963 (.L_HI(net963));
 sg13g2_tiehi _19265__964 (.L_HI(net964));
 sg13g2_tiehi _19851__965 (.L_HI(net965));
 sg13g2_tiehi _19264__966 (.L_HI(net966));
 sg13g2_tiehi _19850__967 (.L_HI(net967));
 sg13g2_tiehi _19263__968 (.L_HI(net968));
 sg13g2_tiehi _19849__969 (.L_HI(net969));
 sg13g2_tiehi _19262__970 (.L_HI(net970));
 sg13g2_tiehi _19848__971 (.L_HI(net971));
 sg13g2_tiehi _19261__972 (.L_HI(net972));
 sg13g2_tiehi _19847__973 (.L_HI(net973));
 sg13g2_tiehi _19260__974 (.L_HI(net974));
 sg13g2_tiehi _19846__975 (.L_HI(net975));
 sg13g2_tiehi _19259__976 (.L_HI(net976));
 sg13g2_tiehi _19845__977 (.L_HI(net977));
 sg13g2_tiehi _19258__978 (.L_HI(net978));
 sg13g2_tiehi _19844__979 (.L_HI(net979));
 sg13g2_tiehi _19257__980 (.L_HI(net980));
 sg13g2_tiehi _19843__981 (.L_HI(net981));
 sg13g2_tiehi _19256__982 (.L_HI(net982));
 sg13g2_tiehi _19842__983 (.L_HI(net983));
 sg13g2_tiehi _19255__984 (.L_HI(net984));
 sg13g2_tiehi _19841__985 (.L_HI(net985));
 sg13g2_tiehi _19254__986 (.L_HI(net986));
 sg13g2_tiehi _19840__987 (.L_HI(net987));
 sg13g2_tiehi _19253__988 (.L_HI(net988));
 sg13g2_tiehi _19839__989 (.L_HI(net989));
 sg13g2_tiehi _19252__990 (.L_HI(net990));
 sg13g2_tiehi _19838__991 (.L_HI(net991));
 sg13g2_tiehi _19251__992 (.L_HI(net992));
 sg13g2_tiehi _19837__993 (.L_HI(net993));
 sg13g2_tiehi _19250__994 (.L_HI(net994));
 sg13g2_tiehi _19836__995 (.L_HI(net995));
 sg13g2_tiehi _19249__996 (.L_HI(net996));
 sg13g2_tiehi _19835__997 (.L_HI(net997));
 sg13g2_tiehi _19248__998 (.L_HI(net998));
 sg13g2_tiehi _19834__999 (.L_HI(net999));
 sg13g2_tiehi _19247__1000 (.L_HI(net1000));
 sg13g2_tiehi _19833__1001 (.L_HI(net1001));
 sg13g2_tiehi _19246__1002 (.L_HI(net1002));
 sg13g2_tiehi _19832__1003 (.L_HI(net1003));
 sg13g2_tiehi _19245__1004 (.L_HI(net1004));
 sg13g2_tiehi _19831__1005 (.L_HI(net1005));
 sg13g2_tiehi _19244__1006 (.L_HI(net1006));
 sg13g2_tiehi _19830__1007 (.L_HI(net1007));
 sg13g2_tiehi _19243__1008 (.L_HI(net1008));
 sg13g2_tiehi _19829__1009 (.L_HI(net1009));
 sg13g2_tiehi _19242__1010 (.L_HI(net1010));
 sg13g2_tiehi _19828__1011 (.L_HI(net1011));
 sg13g2_tiehi _19241__1012 (.L_HI(net1012));
 sg13g2_tiehi _19827__1013 (.L_HI(net1013));
 sg13g2_tiehi _19240__1014 (.L_HI(net1014));
 sg13g2_tiehi _19239__1015 (.L_HI(net1015));
 sg13g2_tiehi _19238__1016 (.L_HI(net1016));
 sg13g2_tiehi _19237__1017 (.L_HI(net1017));
 sg13g2_tiehi _19236__1018 (.L_HI(net1018));
 sg13g2_tiehi _19235__1019 (.L_HI(net1019));
 sg13g2_tiehi _19234__1020 (.L_HI(net1020));
 sg13g2_tiehi _19233__1021 (.L_HI(net1021));
 sg13g2_tiehi _19232__1022 (.L_HI(net1022));
 sg13g2_tiehi _19231__1023 (.L_HI(net1023));
 sg13g2_tiehi _19230__1024 (.L_HI(net1024));
 sg13g2_tiehi _19229__1025 (.L_HI(net1025));
 sg13g2_tiehi _19228__1026 (.L_HI(net1026));
 sg13g2_tiehi _19826__1027 (.L_HI(net1027));
 sg13g2_tiehi _19227__1028 (.L_HI(net1028));
 sg13g2_tiehi _19226__1029 (.L_HI(net1029));
 sg13g2_tiehi _19225__1030 (.L_HI(net1030));
 sg13g2_tiehi _19224__1031 (.L_HI(net1031));
 sg13g2_tiehi _19223__1032 (.L_HI(net1032));
 sg13g2_tiehi _19222__1033 (.L_HI(net1033));
 sg13g2_tiehi _19221__1034 (.L_HI(net1034));
 sg13g2_tiehi _19220__1035 (.L_HI(net1035));
 sg13g2_tiehi _19219__1036 (.L_HI(net1036));
 sg13g2_tiehi _19218__1037 (.L_HI(net1037));
 sg13g2_tiehi _19217__1038 (.L_HI(net1038));
 sg13g2_tiehi _19216__1039 (.L_HI(net1039));
 sg13g2_tiehi _19215__1040 (.L_HI(net1040));
 sg13g2_tiehi _19214__1041 (.L_HI(net1041));
 sg13g2_tiehi _19213__1042 (.L_HI(net1042));
 sg13g2_tiehi _19212__1043 (.L_HI(net1043));
 sg13g2_tiehi _19211__1044 (.L_HI(net1044));
 sg13g2_tiehi _19210__1045 (.L_HI(net1045));
 sg13g2_tiehi _19209__1046 (.L_HI(net1046));
 sg13g2_tiehi _19208__1047 (.L_HI(net1047));
 sg13g2_tiehi _19207__1048 (.L_HI(net1048));
 sg13g2_tiehi _19206__1049 (.L_HI(net1049));
 sg13g2_tiehi _19205__1050 (.L_HI(net1050));
 sg13g2_tiehi _19204__1051 (.L_HI(net1051));
 sg13g2_tiehi _19203__1052 (.L_HI(net1052));
 sg13g2_tiehi _19202__1053 (.L_HI(net1053));
 sg13g2_tiehi _19201__1054 (.L_HI(net1054));
 sg13g2_tiehi _19200__1055 (.L_HI(net1055));
 sg13g2_tiehi _19199__1056 (.L_HI(net1056));
 sg13g2_tiehi _19198__1057 (.L_HI(net1057));
 sg13g2_tiehi _19197__1058 (.L_HI(net1058));
 sg13g2_tiehi _19196__1059 (.L_HI(net1059));
 sg13g2_tiehi _19195__1060 (.L_HI(net1060));
 sg13g2_tiehi _19194__1061 (.L_HI(net1061));
 sg13g2_tiehi _19193__1062 (.L_HI(net1062));
 sg13g2_tiehi _19192__1063 (.L_HI(net1063));
 sg13g2_tiehi _19191__1064 (.L_HI(net1064));
 sg13g2_tiehi _19190__1065 (.L_HI(net1065));
 sg13g2_tiehi _18289__1066 (.L_HI(net1066));
 sg13g2_tiehi _19337__1067 (.L_HI(net1067));
 sg13g2_tiehi _19338__1068 (.L_HI(net1068));
 sg13g2_tiehi _19339__1069 (.L_HI(net1069));
 sg13g2_tiehi _19340__1070 (.L_HI(net1070));
 sg13g2_tiehi _19341__1071 (.L_HI(net1071));
 sg13g2_tiehi _19342__1072 (.L_HI(net1072));
 sg13g2_tiehi _19343__1073 (.L_HI(net1073));
 sg13g2_tiehi _19344__1074 (.L_HI(net1074));
 sg13g2_tiehi _19345__1075 (.L_HI(net1075));
 sg13g2_tiehi _19346__1076 (.L_HI(net1076));
 sg13g2_tiehi _19347__1077 (.L_HI(net1077));
 sg13g2_tiehi _19348__1078 (.L_HI(net1078));
 sg13g2_tiehi _19349__1079 (.L_HI(net1079));
 sg13g2_tiehi _19350__1080 (.L_HI(net1080));
 sg13g2_tiehi _19351__1081 (.L_HI(net1081));
 sg13g2_tiehi _19825__1082 (.L_HI(net1082));
 sg13g2_tiehi _19189__1083 (.L_HI(net1083));
 sg13g2_tiehi _19824__1084 (.L_HI(net1084));
 sg13g2_tiehi _19188__1085 (.L_HI(net1085));
 sg13g2_tiehi _19823__1086 (.L_HI(net1086));
 sg13g2_tiehi _19187__1087 (.L_HI(net1087));
 sg13g2_tiehi _19822__1088 (.L_HI(net1088));
 sg13g2_tiehi _19186__1089 (.L_HI(net1089));
 sg13g2_tiehi _19821__1090 (.L_HI(net1090));
 sg13g2_tiehi _19185__1091 (.L_HI(net1091));
 sg13g2_tiehi _19820__1092 (.L_HI(net1092));
 sg13g2_tiehi _19184__1093 (.L_HI(net1093));
 sg13g2_tiehi _19819__1094 (.L_HI(net1094));
 sg13g2_tiehi _19183__1095 (.L_HI(net1095));
 sg13g2_tiehi _19818__1096 (.L_HI(net1096));
 sg13g2_tiehi _19182__1097 (.L_HI(net1097));
 sg13g2_tiehi _19181__1098 (.L_HI(net1098));
 sg13g2_tiehi _19817__1099 (.L_HI(net1099));
 sg13g2_tiehi _19180__1100 (.L_HI(net1100));
 sg13g2_tiehi _19816__1101 (.L_HI(net1101));
 sg13g2_tiehi _19179__1102 (.L_HI(net1102));
 sg13g2_tiehi _19815__1103 (.L_HI(net1103));
 sg13g2_tiehi _19178__1104 (.L_HI(net1104));
 sg13g2_tiehi _19814__1105 (.L_HI(net1105));
 sg13g2_tiehi _19177__1106 (.L_HI(net1106));
 sg13g2_tiehi _19813__1107 (.L_HI(net1107));
 sg13g2_tiehi _19176__1108 (.L_HI(net1108));
 sg13g2_tiehi _19812__1109 (.L_HI(net1109));
 sg13g2_tiehi _19352__1110 (.L_HI(net1110));
 sg13g2_tiehi _19381__1111 (.L_HI(net1111));
 sg13g2_tiehi _19382__1112 (.L_HI(net1112));
 sg13g2_tiehi _19383__1113 (.L_HI(net1113));
 sg13g2_tiehi _19384__1114 (.L_HI(net1114));
 sg13g2_tiehi _19385__1115 (.L_HI(net1115));
 sg13g2_tiehi _19386__1116 (.L_HI(net1116));
 sg13g2_tiehi _19387__1117 (.L_HI(net1117));
 sg13g2_tiehi _19388__1118 (.L_HI(net1118));
 sg13g2_tiehi _19389__1119 (.L_HI(net1119));
 sg13g2_tiehi _19390__1120 (.L_HI(net1120));
 sg13g2_tiehi _19391__1121 (.L_HI(net1121));
 sg13g2_tiehi _19392__1122 (.L_HI(net1122));
 sg13g2_tiehi _19393__1123 (.L_HI(net1123));
 sg13g2_tiehi _19394__1124 (.L_HI(net1124));
 sg13g2_tiehi _19395__1125 (.L_HI(net1125));
 sg13g2_tiehi _19175__1126 (.L_HI(net1126));
 sg13g2_tiehi _19811__1127 (.L_HI(net1127));
 sg13g2_tiehi _19174__1128 (.L_HI(net1128));
 sg13g2_tiehi _19810__1129 (.L_HI(net1129));
 sg13g2_tiehi _19173__1130 (.L_HI(net1130));
 sg13g2_tiehi _19809__1131 (.L_HI(net1131));
 sg13g2_tiehi _19172__1132 (.L_HI(net1132));
 sg13g2_tiehi _19808__1133 (.L_HI(net1133));
 sg13g2_tiehi _19396__1134 (.L_HI(net1134));
 sg13g2_tiehi _19405__1135 (.L_HI(net1135));
 sg13g2_tiehi _19406__1136 (.L_HI(net1136));
 sg13g2_tiehi _19407__1137 (.L_HI(net1137));
 sg13g2_tiehi _19408__1138 (.L_HI(net1138));
 sg13g2_tiehi _19409__1139 (.L_HI(net1139));
 sg13g2_tiehi _19410__1140 (.L_HI(net1140));
 sg13g2_tiehi _19411__1141 (.L_HI(net1141));
 sg13g2_tiehi _19171__1142 (.L_HI(net1142));
 sg13g2_tiehi _19807__1143 (.L_HI(net1143));
 sg13g2_tiehi _19170__1144 (.L_HI(net1144));
 sg13g2_tiehi _19806__1145 (.L_HI(net1145));
 sg13g2_tiehi _19169__1146 (.L_HI(net1146));
 sg13g2_tiehi _19805__1147 (.L_HI(net1147));
 sg13g2_tiehi _19168__1148 (.L_HI(net1148));
 sg13g2_tiehi _19167__1149 (.L_HI(net1149));
 sg13g2_tiehi _19166__1150 (.L_HI(net1150));
 sg13g2_tiehi _19165__1151 (.L_HI(net1151));
 sg13g2_tiehi _19164__1152 (.L_HI(net1152));
 sg13g2_tiehi _19163__1153 (.L_HI(net1153));
 sg13g2_tiehi _19162__1154 (.L_HI(net1154));
 sg13g2_tiehi _19161__1155 (.L_HI(net1155));
 sg13g2_tiehi _19160__1156 (.L_HI(net1156));
 sg13g2_tiehi _19159__1157 (.L_HI(net1157));
 sg13g2_tiehi _19158__1158 (.L_HI(net1158));
 sg13g2_tiehi _19157__1159 (.L_HI(net1159));
 sg13g2_tiehi _19156__1160 (.L_HI(net1160));
 sg13g2_tiehi _19155__1161 (.L_HI(net1161));
 sg13g2_tiehi _19154__1162 (.L_HI(net1162));
 sg13g2_tiehi _19153__1163 (.L_HI(net1163));
 sg13g2_tiehi _19152__1164 (.L_HI(net1164));
 sg13g2_tiehi _19151__1165 (.L_HI(net1165));
 sg13g2_tiehi _19150__1166 (.L_HI(net1166));
 sg13g2_tiehi _19149__1167 (.L_HI(net1167));
 sg13g2_tiehi _19148__1168 (.L_HI(net1168));
 sg13g2_tiehi _19147__1169 (.L_HI(net1169));
 sg13g2_tiehi _19146__1170 (.L_HI(net1170));
 sg13g2_tiehi _19145__1171 (.L_HI(net1171));
 sg13g2_tiehi _19144__1172 (.L_HI(net1172));
 sg13g2_tiehi _19143__1173 (.L_HI(net1173));
 sg13g2_tiehi _19142__1174 (.L_HI(net1174));
 sg13g2_tiehi _19141__1175 (.L_HI(net1175));
 sg13g2_tiehi _19140__1176 (.L_HI(net1176));
 sg13g2_tiehi _19139__1177 (.L_HI(net1177));
 sg13g2_tiehi _19138__1178 (.L_HI(net1178));
 sg13g2_tiehi _19137__1179 (.L_HI(net1179));
 sg13g2_tiehi _19136__1180 (.L_HI(net1180));
 sg13g2_tiehi _19135__1181 (.L_HI(net1181));
 sg13g2_tiehi _19134__1182 (.L_HI(net1182));
 sg13g2_tiehi _19133__1183 (.L_HI(net1183));
 sg13g2_tiehi _19132__1184 (.L_HI(net1184));
 sg13g2_tiehi _19131__1185 (.L_HI(net1185));
 sg13g2_tiehi _19130__1186 (.L_HI(net1186));
 sg13g2_tiehi _19129__1187 (.L_HI(net1187));
 sg13g2_tiehi _19128__1188 (.L_HI(net1188));
 sg13g2_tiehi _19127__1189 (.L_HI(net1189));
 sg13g2_tiehi _19126__1190 (.L_HI(net1190));
 sg13g2_tiehi _19125__1191 (.L_HI(net1191));
 sg13g2_tiehi _19124__1192 (.L_HI(net1192));
 sg13g2_tiehi _19123__1193 (.L_HI(net1193));
 sg13g2_tiehi _19122__1194 (.L_HI(net1194));
 sg13g2_tiehi _19121__1195 (.L_HI(net1195));
 sg13g2_tiehi _19120__1196 (.L_HI(net1196));
 sg13g2_tiehi _19119__1197 (.L_HI(net1197));
 sg13g2_tiehi _19118__1198 (.L_HI(net1198));
 sg13g2_tiehi _19117__1199 (.L_HI(net1199));
 sg13g2_tiehi _19116__1200 (.L_HI(net1200));
 sg13g2_tiehi _19115__1201 (.L_HI(net1201));
 sg13g2_tiehi _19114__1202 (.L_HI(net1202));
 sg13g2_tiehi _19113__1203 (.L_HI(net1203));
 sg13g2_tiehi _19112__1204 (.L_HI(net1204));
 sg13g2_tiehi _19111__1205 (.L_HI(net1205));
 sg13g2_tiehi _19110__1206 (.L_HI(net1206));
 sg13g2_tiehi _19109__1207 (.L_HI(net1207));
 sg13g2_tiehi _19108__1208 (.L_HI(net1208));
 sg13g2_tiehi _19107__1209 (.L_HI(net1209));
 sg13g2_tiehi _19106__1210 (.L_HI(net1210));
 sg13g2_tiehi _19105__1211 (.L_HI(net1211));
 sg13g2_tiehi _19104__1212 (.L_HI(net1212));
 sg13g2_tiehi _19103__1213 (.L_HI(net1213));
 sg13g2_tiehi _19102__1214 (.L_HI(net1214));
 sg13g2_tiehi _19101__1215 (.L_HI(net1215));
 sg13g2_tiehi _19100__1216 (.L_HI(net1216));
 sg13g2_tiehi _19099__1217 (.L_HI(net1217));
 sg13g2_tiehi _19098__1218 (.L_HI(net1218));
 sg13g2_tiehi _19097__1219 (.L_HI(net1219));
 sg13g2_tiehi _19096__1220 (.L_HI(net1220));
 sg13g2_tiehi _19095__1221 (.L_HI(net1221));
 sg13g2_tiehi _19094__1222 (.L_HI(net1222));
 sg13g2_tiehi _19093__1223 (.L_HI(net1223));
 sg13g2_tiehi _19092__1224 (.L_HI(net1224));
 sg13g2_tiehi _19091__1225 (.L_HI(net1225));
 sg13g2_tiehi _19090__1226 (.L_HI(net1226));
 sg13g2_tiehi _19089__1227 (.L_HI(net1227));
 sg13g2_tiehi _19088__1228 (.L_HI(net1228));
 sg13g2_tiehi _19087__1229 (.L_HI(net1229));
 sg13g2_tiehi _19086__1230 (.L_HI(net1230));
 sg13g2_tiehi _19085__1231 (.L_HI(net1231));
 sg13g2_tiehi _19084__1232 (.L_HI(net1232));
 sg13g2_tiehi _19083__1233 (.L_HI(net1233));
 sg13g2_tiehi _19082__1234 (.L_HI(net1234));
 sg13g2_tiehi _19081__1235 (.L_HI(net1235));
 sg13g2_tiehi _19080__1236 (.L_HI(net1236));
 sg13g2_tiehi _19079__1237 (.L_HI(net1237));
 sg13g2_tiehi _19078__1238 (.L_HI(net1238));
 sg13g2_tiehi _19077__1239 (.L_HI(net1239));
 sg13g2_tiehi _19076__1240 (.L_HI(net1240));
 sg13g2_tiehi _19075__1241 (.L_HI(net1241));
 sg13g2_tiehi _19074__1242 (.L_HI(net1242));
 sg13g2_tiehi _19073__1243 (.L_HI(net1243));
 sg13g2_tiehi _19072__1244 (.L_HI(net1244));
 sg13g2_tiehi _19071__1245 (.L_HI(net1245));
 sg13g2_tiehi _19070__1246 (.L_HI(net1246));
 sg13g2_tiehi _19069__1247 (.L_HI(net1247));
 sg13g2_tiehi _19068__1248 (.L_HI(net1248));
 sg13g2_tiehi _19067__1249 (.L_HI(net1249));
 sg13g2_tiehi _19066__1250 (.L_HI(net1250));
 sg13g2_tiehi _19065__1251 (.L_HI(net1251));
 sg13g2_tiehi _19064__1252 (.L_HI(net1252));
 sg13g2_tiehi _19063__1253 (.L_HI(net1253));
 sg13g2_tiehi _19062__1254 (.L_HI(net1254));
 sg13g2_tiehi _19061__1255 (.L_HI(net1255));
 sg13g2_tiehi _19060__1256 (.L_HI(net1256));
 sg13g2_tiehi _19059__1257 (.L_HI(net1257));
 sg13g2_tiehi _19058__1258 (.L_HI(net1258));
 sg13g2_tiehi _19057__1259 (.L_HI(net1259));
 sg13g2_tiehi _19056__1260 (.L_HI(net1260));
 sg13g2_tiehi _19055__1261 (.L_HI(net1261));
 sg13g2_tiehi _19054__1262 (.L_HI(net1262));
 sg13g2_tiehi _19053__1263 (.L_HI(net1263));
 sg13g2_tiehi _19052__1264 (.L_HI(net1264));
 sg13g2_tiehi _19051__1265 (.L_HI(net1265));
 sg13g2_tiehi _19050__1266 (.L_HI(net1266));
 sg13g2_tiehi _19049__1267 (.L_HI(net1267));
 sg13g2_tiehi _19048__1268 (.L_HI(net1268));
 sg13g2_tiehi _19047__1269 (.L_HI(net1269));
 sg13g2_tiehi _19046__1270 (.L_HI(net1270));
 sg13g2_tiehi _19045__1271 (.L_HI(net1271));
 sg13g2_tiehi _19044__1272 (.L_HI(net1272));
 sg13g2_tiehi _19043__1273 (.L_HI(net1273));
 sg13g2_tiehi _19042__1274 (.L_HI(net1274));
 sg13g2_tiehi _19041__1275 (.L_HI(net1275));
 sg13g2_tiehi _19040__1276 (.L_HI(net1276));
 sg13g2_tiehi _19039__1277 (.L_HI(net1277));
 sg13g2_tiehi _19038__1278 (.L_HI(net1278));
 sg13g2_tiehi _19037__1279 (.L_HI(net1279));
 sg13g2_tiehi _19036__1280 (.L_HI(net1280));
 sg13g2_tiehi _19035__1281 (.L_HI(net1281));
 sg13g2_tiehi _19034__1282 (.L_HI(net1282));
 sg13g2_tiehi _19033__1283 (.L_HI(net1283));
 sg13g2_tiehi _19032__1284 (.L_HI(net1284));
 sg13g2_tiehi _19031__1285 (.L_HI(net1285));
 sg13g2_tiehi _19030__1286 (.L_HI(net1286));
 sg13g2_tiehi _19029__1287 (.L_HI(net1287));
 sg13g2_tiehi _19028__1288 (.L_HI(net1288));
 sg13g2_tiehi _19027__1289 (.L_HI(net1289));
 sg13g2_tiehi _19026__1290 (.L_HI(net1290));
 sg13g2_tiehi _19025__1291 (.L_HI(net1291));
 sg13g2_tiehi _19024__1292 (.L_HI(net1292));
 sg13g2_tiehi _19023__1293 (.L_HI(net1293));
 sg13g2_tiehi _19022__1294 (.L_HI(net1294));
 sg13g2_tiehi _19021__1295 (.L_HI(net1295));
 sg13g2_tiehi _19020__1296 (.L_HI(net1296));
 sg13g2_tiehi _19019__1297 (.L_HI(net1297));
 sg13g2_tiehi _19018__1298 (.L_HI(net1298));
 sg13g2_tiehi _19017__1299 (.L_HI(net1299));
 sg13g2_tiehi _19016__1300 (.L_HI(net1300));
 sg13g2_tiehi _19015__1301 (.L_HI(net1301));
 sg13g2_tiehi _19014__1302 (.L_HI(net1302));
 sg13g2_tiehi _19013__1303 (.L_HI(net1303));
 sg13g2_tiehi _19012__1304 (.L_HI(net1304));
 sg13g2_tiehi _19011__1305 (.L_HI(net1305));
 sg13g2_tiehi _19010__1306 (.L_HI(net1306));
 sg13g2_tiehi _19009__1307 (.L_HI(net1307));
 sg13g2_tiehi _19008__1308 (.L_HI(net1308));
 sg13g2_tiehi _19007__1309 (.L_HI(net1309));
 sg13g2_tiehi _19006__1310 (.L_HI(net1310));
 sg13g2_tiehi _19005__1311 (.L_HI(net1311));
 sg13g2_tiehi _19004__1312 (.L_HI(net1312));
 sg13g2_tiehi _19003__1313 (.L_HI(net1313));
 sg13g2_tiehi _19002__1314 (.L_HI(net1314));
 sg13g2_tiehi _19001__1315 (.L_HI(net1315));
 sg13g2_tiehi _19000__1316 (.L_HI(net1316));
 sg13g2_tiehi _18999__1317 (.L_HI(net1317));
 sg13g2_tiehi _18998__1318 (.L_HI(net1318));
 sg13g2_tiehi _18997__1319 (.L_HI(net1319));
 sg13g2_tiehi _18996__1320 (.L_HI(net1320));
 sg13g2_tiehi _18995__1321 (.L_HI(net1321));
 sg13g2_tiehi _18994__1322 (.L_HI(net1322));
 sg13g2_tiehi _18993__1323 (.L_HI(net1323));
 sg13g2_tiehi _18992__1324 (.L_HI(net1324));
 sg13g2_tiehi _18991__1325 (.L_HI(net1325));
 sg13g2_tiehi _18990__1326 (.L_HI(net1326));
 sg13g2_tiehi _18989__1327 (.L_HI(net1327));
 sg13g2_tiehi _18988__1328 (.L_HI(net1328));
 sg13g2_tiehi _18987__1329 (.L_HI(net1329));
 sg13g2_tiehi _18986__1330 (.L_HI(net1330));
 sg13g2_tiehi _18985__1331 (.L_HI(net1331));
 sg13g2_tiehi _18984__1332 (.L_HI(net1332));
 sg13g2_tiehi _18983__1333 (.L_HI(net1333));
 sg13g2_tiehi _18982__1334 (.L_HI(net1334));
 sg13g2_tiehi _18981__1335 (.L_HI(net1335));
 sg13g2_tiehi _18980__1336 (.L_HI(net1336));
 sg13g2_tiehi _18979__1337 (.L_HI(net1337));
 sg13g2_tiehi _18978__1338 (.L_HI(net1338));
 sg13g2_tiehi _18977__1339 (.L_HI(net1339));
 sg13g2_tiehi _18976__1340 (.L_HI(net1340));
 sg13g2_tiehi _18975__1341 (.L_HI(net1341));
 sg13g2_tiehi _18974__1342 (.L_HI(net1342));
 sg13g2_tiehi _18973__1343 (.L_HI(net1343));
 sg13g2_tiehi _18972__1344 (.L_HI(net1344));
 sg13g2_tiehi _18971__1345 (.L_HI(net1345));
 sg13g2_tiehi _18970__1346 (.L_HI(net1346));
 sg13g2_tiehi _18969__1347 (.L_HI(net1347));
 sg13g2_tiehi _18968__1348 (.L_HI(net1348));
 sg13g2_tiehi _18967__1349 (.L_HI(net1349));
 sg13g2_tiehi _18966__1350 (.L_HI(net1350));
 sg13g2_tiehi _18965__1351 (.L_HI(net1351));
 sg13g2_tiehi _18964__1352 (.L_HI(net1352));
 sg13g2_tiehi _18963__1353 (.L_HI(net1353));
 sg13g2_tiehi _18962__1354 (.L_HI(net1354));
 sg13g2_tiehi _18961__1355 (.L_HI(net1355));
 sg13g2_tiehi _18960__1356 (.L_HI(net1356));
 sg13g2_tiehi _18959__1357 (.L_HI(net1357));
 sg13g2_tiehi _18958__1358 (.L_HI(net1358));
 sg13g2_tiehi _18957__1359 (.L_HI(net1359));
 sg13g2_tiehi _18956__1360 (.L_HI(net1360));
 sg13g2_tiehi _18955__1361 (.L_HI(net1361));
 sg13g2_tiehi _18954__1362 (.L_HI(net1362));
 sg13g2_tiehi _18953__1363 (.L_HI(net1363));
 sg13g2_tiehi _18952__1364 (.L_HI(net1364));
 sg13g2_tiehi _18951__1365 (.L_HI(net1365));
 sg13g2_tiehi _18950__1366 (.L_HI(net1366));
 sg13g2_tiehi _18949__1367 (.L_HI(net1367));
 sg13g2_tiehi _18948__1368 (.L_HI(net1368));
 sg13g2_tiehi _18947__1369 (.L_HI(net1369));
 sg13g2_tiehi _18946__1370 (.L_HI(net1370));
 sg13g2_tiehi _18945__1371 (.L_HI(net1371));
 sg13g2_tiehi _18944__1372 (.L_HI(net1372));
 sg13g2_tiehi _18943__1373 (.L_HI(net1373));
 sg13g2_tiehi _18942__1374 (.L_HI(net1374));
 sg13g2_tiehi _18941__1375 (.L_HI(net1375));
 sg13g2_tiehi _18940__1376 (.L_HI(net1376));
 sg13g2_tiehi _18939__1377 (.L_HI(net1377));
 sg13g2_tiehi _18938__1378 (.L_HI(net1378));
 sg13g2_tiehi _18937__1379 (.L_HI(net1379));
 sg13g2_tiehi _18936__1380 (.L_HI(net1380));
 sg13g2_tiehi _18935__1381 (.L_HI(net1381));
 sg13g2_tiehi _18934__1382 (.L_HI(net1382));
 sg13g2_tiehi _18933__1383 (.L_HI(net1383));
 sg13g2_tiehi _18932__1384 (.L_HI(net1384));
 sg13g2_tiehi _18931__1385 (.L_HI(net1385));
 sg13g2_tiehi _18930__1386 (.L_HI(net1386));
 sg13g2_tiehi _18929__1387 (.L_HI(net1387));
 sg13g2_tiehi _18928__1388 (.L_HI(net1388));
 sg13g2_tiehi _18927__1389 (.L_HI(net1389));
 sg13g2_tiehi _18926__1390 (.L_HI(net1390));
 sg13g2_tiehi _18925__1391 (.L_HI(net1391));
 sg13g2_tiehi _18924__1392 (.L_HI(net1392));
 sg13g2_tiehi _18923__1393 (.L_HI(net1393));
 sg13g2_tiehi _18922__1394 (.L_HI(net1394));
 sg13g2_tiehi _18921__1395 (.L_HI(net1395));
 sg13g2_tiehi _18920__1396 (.L_HI(net1396));
 sg13g2_tiehi _18919__1397 (.L_HI(net1397));
 sg13g2_tiehi _18918__1398 (.L_HI(net1398));
 sg13g2_tiehi _18917__1399 (.L_HI(net1399));
 sg13g2_tiehi _18916__1400 (.L_HI(net1400));
 sg13g2_tiehi _18915__1401 (.L_HI(net1401));
 sg13g2_tiehi _18914__1402 (.L_HI(net1402));
 sg13g2_tiehi _18913__1403 (.L_HI(net1403));
 sg13g2_tiehi _18912__1404 (.L_HI(net1404));
 sg13g2_tiehi _18911__1405 (.L_HI(net1405));
 sg13g2_tiehi _18910__1406 (.L_HI(net1406));
 sg13g2_tiehi _18909__1407 (.L_HI(net1407));
 sg13g2_tiehi _18908__1408 (.L_HI(net1408));
 sg13g2_tiehi _18907__1409 (.L_HI(net1409));
 sg13g2_tiehi _18906__1410 (.L_HI(net1410));
 sg13g2_tiehi _18905__1411 (.L_HI(net1411));
 sg13g2_tiehi _18904__1412 (.L_HI(net1412));
 sg13g2_tiehi _18903__1413 (.L_HI(net1413));
 sg13g2_tiehi _18902__1414 (.L_HI(net1414));
 sg13g2_tiehi _18901__1415 (.L_HI(net1415));
 sg13g2_tiehi _18900__1416 (.L_HI(net1416));
 sg13g2_tiehi _18899__1417 (.L_HI(net1417));
 sg13g2_tiehi _18898__1418 (.L_HI(net1418));
 sg13g2_tiehi _18897__1419 (.L_HI(net1419));
 sg13g2_tiehi _18896__1420 (.L_HI(net1420));
 sg13g2_tiehi _18895__1421 (.L_HI(net1421));
 sg13g2_tiehi _18894__1422 (.L_HI(net1422));
 sg13g2_tiehi _18893__1423 (.L_HI(net1423));
 sg13g2_tiehi _18892__1424 (.L_HI(net1424));
 sg13g2_tiehi _18891__1425 (.L_HI(net1425));
 sg13g2_tiehi _18890__1426 (.L_HI(net1426));
 sg13g2_tiehi _18889__1427 (.L_HI(net1427));
 sg13g2_tiehi _18888__1428 (.L_HI(net1428));
 sg13g2_tiehi _18887__1429 (.L_HI(net1429));
 sg13g2_tiehi _18886__1430 (.L_HI(net1430));
 sg13g2_tiehi _18885__1431 (.L_HI(net1431));
 sg13g2_tiehi _18884__1432 (.L_HI(net1432));
 sg13g2_tiehi _18883__1433 (.L_HI(net1433));
 sg13g2_tiehi _18882__1434 (.L_HI(net1434));
 sg13g2_tiehi _18881__1435 (.L_HI(net1435));
 sg13g2_tiehi _18880__1436 (.L_HI(net1436));
 sg13g2_tiehi _18879__1437 (.L_HI(net1437));
 sg13g2_tiehi _18878__1438 (.L_HI(net1438));
 sg13g2_tiehi _18877__1439 (.L_HI(net1439));
 sg13g2_tiehi _18876__1440 (.L_HI(net1440));
 sg13g2_tiehi _18875__1441 (.L_HI(net1441));
 sg13g2_tiehi _18874__1442 (.L_HI(net1442));
 sg13g2_tiehi _18873__1443 (.L_HI(net1443));
 sg13g2_tiehi _18872__1444 (.L_HI(net1444));
 sg13g2_tiehi _19804__1445 (.L_HI(net1445));
 sg13g2_tiehi _18871__1446 (.L_HI(net1446));
 sg13g2_tiehi _18870__1447 (.L_HI(net1447));
 sg13g2_tiehi _18869__1448 (.L_HI(net1448));
 sg13g2_tiehi _18868__1449 (.L_HI(net1449));
 sg13g2_tiehi _18867__1450 (.L_HI(net1450));
 sg13g2_tiehi _18866__1451 (.L_HI(net1451));
 sg13g2_tiehi _18865__1452 (.L_HI(net1452));
 sg13g2_tiehi _18864__1453 (.L_HI(net1453));
 sg13g2_tiehi _18863__1454 (.L_HI(net1454));
 sg13g2_tiehi _18862__1455 (.L_HI(net1455));
 sg13g2_tiehi _18861__1456 (.L_HI(net1456));
 sg13g2_tiehi _18860__1457 (.L_HI(net1457));
 sg13g2_tiehi _18859__1458 (.L_HI(net1458));
 sg13g2_tiehi _18858__1459 (.L_HI(net1459));
 sg13g2_tiehi _18857__1460 (.L_HI(net1460));
 sg13g2_tiehi _18856__1461 (.L_HI(net1461));
 sg13g2_tiehi _18855__1462 (.L_HI(net1462));
 sg13g2_tiehi _18854__1463 (.L_HI(net1463));
 sg13g2_tiehi _18853__1464 (.L_HI(net1464));
 sg13g2_tiehi _18852__1465 (.L_HI(net1465));
 sg13g2_tiehi _18851__1466 (.L_HI(net1466));
 sg13g2_tiehi _18850__1467 (.L_HI(net1467));
 sg13g2_tiehi _18849__1468 (.L_HI(net1468));
 sg13g2_tiehi _18848__1469 (.L_HI(net1469));
 sg13g2_tiehi _18847__1470 (.L_HI(net1470));
 sg13g2_tiehi _18846__1471 (.L_HI(net1471));
 sg13g2_tiehi _18845__1472 (.L_HI(net1472));
 sg13g2_tiehi _18844__1473 (.L_HI(net1473));
 sg13g2_tiehi _18843__1474 (.L_HI(net1474));
 sg13g2_tiehi _18842__1475 (.L_HI(net1475));
 sg13g2_tiehi _18841__1476 (.L_HI(net1476));
 sg13g2_tiehi _18840__1477 (.L_HI(net1477));
 sg13g2_tiehi _18839__1478 (.L_HI(net1478));
 sg13g2_tiehi _18838__1479 (.L_HI(net1479));
 sg13g2_tiehi _18837__1480 (.L_HI(net1480));
 sg13g2_tiehi _18836__1481 (.L_HI(net1481));
 sg13g2_tiehi _18835__1482 (.L_HI(net1482));
 sg13g2_tiehi _18834__1483 (.L_HI(net1483));
 sg13g2_tiehi _18833__1484 (.L_HI(net1484));
 sg13g2_tiehi _18832__1485 (.L_HI(net1485));
 sg13g2_tiehi _18831__1486 (.L_HI(net1486));
 sg13g2_tiehi _18830__1487 (.L_HI(net1487));
 sg13g2_tiehi _18829__1488 (.L_HI(net1488));
 sg13g2_tiehi _18828__1489 (.L_HI(net1489));
 sg13g2_tiehi _18827__1490 (.L_HI(net1490));
 sg13g2_tiehi _18826__1491 (.L_HI(net1491));
 sg13g2_tiehi _18825__1492 (.L_HI(net1492));
 sg13g2_tiehi _18824__1493 (.L_HI(net1493));
 sg13g2_tiehi _18823__1494 (.L_HI(net1494));
 sg13g2_tiehi _18822__1495 (.L_HI(net1495));
 sg13g2_tiehi _18821__1496 (.L_HI(net1496));
 sg13g2_tiehi _18820__1497 (.L_HI(net1497));
 sg13g2_tiehi _18819__1498 (.L_HI(net1498));
 sg13g2_tiehi _18818__1499 (.L_HI(net1499));
 sg13g2_tiehi _18817__1500 (.L_HI(net1500));
 sg13g2_tiehi _18816__1501 (.L_HI(net1501));
 sg13g2_tiehi _18815__1502 (.L_HI(net1502));
 sg13g2_tiehi _18814__1503 (.L_HI(net1503));
 sg13g2_tiehi _18813__1504 (.L_HI(net1504));
 sg13g2_tiehi _18812__1505 (.L_HI(net1505));
 sg13g2_tiehi _18811__1506 (.L_HI(net1506));
 sg13g2_tiehi _18810__1507 (.L_HI(net1507));
 sg13g2_tiehi _18809__1508 (.L_HI(net1508));
 sg13g2_tiehi _18808__1509 (.L_HI(net1509));
 sg13g2_tiehi _18807__1510 (.L_HI(net1510));
 sg13g2_tiehi _19803__1511 (.L_HI(net1511));
 sg13g2_tiehi _18806__1512 (.L_HI(net1512));
 sg13g2_tiehi _19802__1513 (.L_HI(net1513));
 sg13g2_tiehi _18805__1514 (.L_HI(net1514));
 sg13g2_tiehi _19801__1515 (.L_HI(net1515));
 sg13g2_tiehi _18804__1516 (.L_HI(net1516));
 sg13g2_tiehi _19800__1517 (.L_HI(net1517));
 sg13g2_tiehi _18803__1518 (.L_HI(net1518));
 sg13g2_tiehi _19799__1519 (.L_HI(net1519));
 sg13g2_tiehi _18802__1520 (.L_HI(net1520));
 sg13g2_tiehi _19798__1521 (.L_HI(net1521));
 sg13g2_tiehi _18801__1522 (.L_HI(net1522));
 sg13g2_tiehi _19797__1523 (.L_HI(net1523));
 sg13g2_tiehi _18800__1524 (.L_HI(net1524));
 sg13g2_tiehi _19796__1525 (.L_HI(net1525));
 sg13g2_tiehi _18799__1526 (.L_HI(net1526));
 sg13g2_tiehi _19795__1527 (.L_HI(net1527));
 sg13g2_tiehi _18798__1528 (.L_HI(net1528));
 sg13g2_tiehi _19794__1529 (.L_HI(net1529));
 sg13g2_tiehi _18797__1530 (.L_HI(net1530));
 sg13g2_tiehi _18796__1531 (.L_HI(net1531));
 sg13g2_tiehi _18795__1532 (.L_HI(net1532));
 sg13g2_tiehi _18794__1533 (.L_HI(net1533));
 sg13g2_tiehi _18793__1534 (.L_HI(net1534));
 sg13g2_tiehi _18792__1535 (.L_HI(net1535));
 sg13g2_tiehi _18791__1536 (.L_HI(net1536));
 sg13g2_tiehi _18790__1537 (.L_HI(net1537));
 sg13g2_tiehi _18789__1538 (.L_HI(net1538));
 sg13g2_tiehi _18788__1539 (.L_HI(net1539));
 sg13g2_tiehi _18787__1540 (.L_HI(net1540));
 sg13g2_tiehi _18786__1541 (.L_HI(net1541));
 sg13g2_tiehi _18785__1542 (.L_HI(net1542));
 sg13g2_tiehi _18784__1543 (.L_HI(net1543));
 sg13g2_tiehi _18783__1544 (.L_HI(net1544));
 sg13g2_tiehi _18782__1545 (.L_HI(net1545));
 sg13g2_tiehi _18781__1546 (.L_HI(net1546));
 sg13g2_tiehi _18780__1547 (.L_HI(net1547));
 sg13g2_tiehi _18779__1548 (.L_HI(net1548));
 sg13g2_tiehi _18778__1549 (.L_HI(net1549));
 sg13g2_tiehi _18777__1550 (.L_HI(net1550));
 sg13g2_tiehi _18776__1551 (.L_HI(net1551));
 sg13g2_tiehi _18775__1552 (.L_HI(net1552));
 sg13g2_tiehi _18774__1553 (.L_HI(net1553));
 sg13g2_tiehi _18773__1554 (.L_HI(net1554));
 sg13g2_tiehi _18772__1555 (.L_HI(net1555));
 sg13g2_tiehi _18771__1556 (.L_HI(net1556));
 sg13g2_tiehi _18770__1557 (.L_HI(net1557));
 sg13g2_tiehi _18769__1558 (.L_HI(net1558));
 sg13g2_tiehi _18768__1559 (.L_HI(net1559));
 sg13g2_tiehi _18767__1560 (.L_HI(net1560));
 sg13g2_tiehi _18766__1561 (.L_HI(net1561));
 sg13g2_tiehi _18765__1562 (.L_HI(net1562));
 sg13g2_tiehi _18764__1563 (.L_HI(net1563));
 sg13g2_tiehi _18763__1564 (.L_HI(net1564));
 sg13g2_tiehi _18762__1565 (.L_HI(net1565));
 sg13g2_tiehi _18761__1566 (.L_HI(net1566));
 sg13g2_tiehi _18760__1567 (.L_HI(net1567));
 sg13g2_tiehi _18759__1568 (.L_HI(net1568));
 sg13g2_tiehi _18758__1569 (.L_HI(net1569));
 sg13g2_tiehi _18757__1570 (.L_HI(net1570));
 sg13g2_tiehi _18756__1571 (.L_HI(net1571));
 sg13g2_tiehi _18755__1572 (.L_HI(net1572));
 sg13g2_tiehi _18754__1573 (.L_HI(net1573));
 sg13g2_tiehi _18753__1574 (.L_HI(net1574));
 sg13g2_tiehi _18752__1575 (.L_HI(net1575));
 sg13g2_tiehi _18751__1576 (.L_HI(net1576));
 sg13g2_tiehi _18750__1577 (.L_HI(net1577));
 sg13g2_tiehi _18749__1578 (.L_HI(net1578));
 sg13g2_tiehi _18748__1579 (.L_HI(net1579));
 sg13g2_tiehi _18747__1580 (.L_HI(net1580));
 sg13g2_tiehi _18746__1581 (.L_HI(net1581));
 sg13g2_tiehi _18745__1582 (.L_HI(net1582));
 sg13g2_tiehi _18744__1583 (.L_HI(net1583));
 sg13g2_tiehi _18743__1584 (.L_HI(net1584));
 sg13g2_tiehi _18742__1585 (.L_HI(net1585));
 sg13g2_tiehi _18741__1586 (.L_HI(net1586));
 sg13g2_tiehi _18740__1587 (.L_HI(net1587));
 sg13g2_tiehi _18739__1588 (.L_HI(net1588));
 sg13g2_tiehi _18738__1589 (.L_HI(net1589));
 sg13g2_tiehi _18737__1590 (.L_HI(net1590));
 sg13g2_tiehi _18736__1591 (.L_HI(net1591));
 sg13g2_tiehi _18735__1592 (.L_HI(net1592));
 sg13g2_tiehi _18734__1593 (.L_HI(net1593));
 sg13g2_tiehi _18733__1594 (.L_HI(net1594));
 sg13g2_tiehi _18732__1595 (.L_HI(net1595));
 sg13g2_tiehi _18731__1596 (.L_HI(net1596));
 sg13g2_tiehi _18730__1597 (.L_HI(net1597));
 sg13g2_tiehi _18729__1598 (.L_HI(net1598));
 sg13g2_tiehi _18728__1599 (.L_HI(net1599));
 sg13g2_tiehi _18727__1600 (.L_HI(net1600));
 sg13g2_tiehi _18726__1601 (.L_HI(net1601));
 sg13g2_tiehi _18725__1602 (.L_HI(net1602));
 sg13g2_tiehi _18724__1603 (.L_HI(net1603));
 sg13g2_tiehi _18723__1604 (.L_HI(net1604));
 sg13g2_tiehi _18722__1605 (.L_HI(net1605));
 sg13g2_tiehi _18721__1606 (.L_HI(net1606));
 sg13g2_tiehi _18720__1607 (.L_HI(net1607));
 sg13g2_tiehi _18719__1608 (.L_HI(net1608));
 sg13g2_tiehi _18718__1609 (.L_HI(net1609));
 sg13g2_tiehi _18717__1610 (.L_HI(net1610));
 sg13g2_tiehi _18716__1611 (.L_HI(net1611));
 sg13g2_tiehi _18715__1612 (.L_HI(net1612));
 sg13g2_tiehi _18714__1613 (.L_HI(net1613));
 sg13g2_tiehi _18713__1614 (.L_HI(net1614));
 sg13g2_tiehi _18712__1615 (.L_HI(net1615));
 sg13g2_tiehi _18711__1616 (.L_HI(net1616));
 sg13g2_tiehi _18710__1617 (.L_HI(net1617));
 sg13g2_tiehi _18709__1618 (.L_HI(net1618));
 sg13g2_tiehi _18708__1619 (.L_HI(net1619));
 sg13g2_tiehi _18707__1620 (.L_HI(net1620));
 sg13g2_tiehi _18706__1621 (.L_HI(net1621));
 sg13g2_tiehi _18705__1622 (.L_HI(net1622));
 sg13g2_tiehi _18704__1623 (.L_HI(net1623));
 sg13g2_tiehi _18703__1624 (.L_HI(net1624));
 sg13g2_tiehi _18702__1625 (.L_HI(net1625));
 sg13g2_tiehi _18701__1626 (.L_HI(net1626));
 sg13g2_tiehi _18700__1627 (.L_HI(net1627));
 sg13g2_tiehi _18699__1628 (.L_HI(net1628));
 sg13g2_tiehi _18698__1629 (.L_HI(net1629));
 sg13g2_tiehi _18697__1630 (.L_HI(net1630));
 sg13g2_tiehi _18696__1631 (.L_HI(net1631));
 sg13g2_tiehi _18695__1632 (.L_HI(net1632));
 sg13g2_tiehi _18694__1633 (.L_HI(net1633));
 sg13g2_tiehi _18693__1634 (.L_HI(net1634));
 sg13g2_tiehi _18692__1635 (.L_HI(net1635));
 sg13g2_tiehi _18691__1636 (.L_HI(net1636));
 sg13g2_tiehi _18690__1637 (.L_HI(net1637));
 sg13g2_tiehi _18689__1638 (.L_HI(net1638));
 sg13g2_tiehi _18688__1639 (.L_HI(net1639));
 sg13g2_tiehi _18687__1640 (.L_HI(net1640));
 sg13g2_tiehi _18686__1641 (.L_HI(net1641));
 sg13g2_tiehi _18685__1642 (.L_HI(net1642));
 sg13g2_tiehi _18684__1643 (.L_HI(net1643));
 sg13g2_tiehi _18683__1644 (.L_HI(net1644));
 sg13g2_tiehi _18682__1645 (.L_HI(net1645));
 sg13g2_tiehi _18681__1646 (.L_HI(net1646));
 sg13g2_tiehi _18680__1647 (.L_HI(net1647));
 sg13g2_tiehi _18679__1648 (.L_HI(net1648));
 sg13g2_tiehi _18678__1649 (.L_HI(net1649));
 sg13g2_tiehi _18677__1650 (.L_HI(net1650));
 sg13g2_tiehi _18676__1651 (.L_HI(net1651));
 sg13g2_tiehi _18675__1652 (.L_HI(net1652));
 sg13g2_tiehi _18674__1653 (.L_HI(net1653));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_2 _21563_ (.A(\m_sys.io_b_uart_tx ),
    .X(uo_out[4]));
 sg13g2_buf_2 fanout4038 (.A(net4039),
    .X(net4038));
 sg13g2_buf_2 fanout4039 (.A(net4040),
    .X(net4039));
 sg13g2_buf_2 fanout4040 (.A(_03540_),
    .X(net4040));
 sg13g2_buf_2 fanout4041 (.A(_02314_),
    .X(net4041));
 sg13g2_buf_4 fanout4042 (.X(net4042),
    .A(_02314_));
 sg13g2_buf_2 fanout4043 (.A(net4044),
    .X(net4043));
 sg13g2_buf_2 fanout4044 (.A(_02305_),
    .X(net4044));
 sg13g2_buf_2 fanout4045 (.A(_02296_),
    .X(net4045));
 sg13g2_buf_2 fanout4046 (.A(_02296_),
    .X(net4046));
 sg13g2_buf_2 fanout4047 (.A(net4048),
    .X(net4047));
 sg13g2_buf_2 fanout4048 (.A(_02287_),
    .X(net4048));
 sg13g2_buf_2 fanout4049 (.A(_02278_),
    .X(net4049));
 sg13g2_buf_2 fanout4050 (.A(_02278_),
    .X(net4050));
 sg13g2_buf_2 fanout4051 (.A(net4052),
    .X(net4051));
 sg13g2_buf_2 fanout4052 (.A(_02269_),
    .X(net4052));
 sg13g2_buf_2 fanout4053 (.A(_02260_),
    .X(net4053));
 sg13g2_buf_2 fanout4054 (.A(_02260_),
    .X(net4054));
 sg13g2_buf_2 fanout4055 (.A(net4056),
    .X(net4055));
 sg13g2_buf_2 fanout4056 (.A(_02251_),
    .X(net4056));
 sg13g2_buf_2 fanout4057 (.A(net4058),
    .X(net4057));
 sg13g2_buf_2 fanout4058 (.A(_02242_),
    .X(net4058));
 sg13g2_buf_2 fanout4059 (.A(_02233_),
    .X(net4059));
 sg13g2_buf_2 fanout4060 (.A(_02233_),
    .X(net4060));
 sg13g2_buf_2 fanout4061 (.A(net4062),
    .X(net4061));
 sg13g2_buf_2 fanout4062 (.A(_02046_),
    .X(net4062));
 sg13g2_buf_2 fanout4063 (.A(_02037_),
    .X(net4063));
 sg13g2_buf_2 fanout4064 (.A(_02037_),
    .X(net4064));
 sg13g2_buf_2 fanout4065 (.A(net4066),
    .X(net4065));
 sg13g2_buf_2 fanout4066 (.A(_02028_),
    .X(net4066));
 sg13g2_buf_2 fanout4067 (.A(net4068),
    .X(net4067));
 sg13g2_buf_2 fanout4068 (.A(_02019_),
    .X(net4068));
 sg13g2_buf_2 fanout4069 (.A(net4070),
    .X(net4069));
 sg13g2_buf_2 fanout4070 (.A(_02010_),
    .X(net4070));
 sg13g2_buf_2 fanout4071 (.A(net4072),
    .X(net4071));
 sg13g2_buf_1 fanout4072 (.A(net4073),
    .X(net4072));
 sg13g2_buf_2 fanout4073 (.A(_02001_),
    .X(net4073));
 sg13g2_buf_2 fanout4074 (.A(_01992_),
    .X(net4074));
 sg13g2_buf_2 fanout4075 (.A(_01992_),
    .X(net4075));
 sg13g2_buf_2 fanout4076 (.A(net4077),
    .X(net4076));
 sg13g2_buf_2 fanout4077 (.A(_01983_),
    .X(net4077));
 sg13g2_buf_2 fanout4078 (.A(_01974_),
    .X(net4078));
 sg13g2_buf_2 fanout4079 (.A(_01974_),
    .X(net4079));
 sg13g2_buf_2 fanout4080 (.A(net4082),
    .X(net4080));
 sg13g2_buf_1 fanout4081 (.A(net4082),
    .X(net4081));
 sg13g2_buf_2 fanout4082 (.A(_01965_),
    .X(net4082));
 sg13g2_buf_2 fanout4083 (.A(_01956_),
    .X(net4083));
 sg13g2_buf_2 fanout4084 (.A(_01956_),
    .X(net4084));
 sg13g2_buf_2 fanout4085 (.A(net4087),
    .X(net4085));
 sg13g2_buf_1 fanout4086 (.A(net4087),
    .X(net4086));
 sg13g2_buf_2 fanout4087 (.A(_01947_),
    .X(net4087));
 sg13g2_buf_2 fanout4088 (.A(net4090),
    .X(net4088));
 sg13g2_buf_1 fanout4089 (.A(net4090),
    .X(net4089));
 sg13g2_buf_2 fanout4090 (.A(_07531_),
    .X(net4090));
 sg13g2_buf_2 fanout4091 (.A(_07522_),
    .X(net4091));
 sg13g2_buf_2 fanout4092 (.A(_07522_),
    .X(net4092));
 sg13g2_buf_2 fanout4093 (.A(net4094),
    .X(net4093));
 sg13g2_buf_2 fanout4094 (.A(_07513_),
    .X(net4094));
 sg13g2_buf_2 fanout4095 (.A(net4096),
    .X(net4095));
 sg13g2_buf_2 fanout4096 (.A(_07504_),
    .X(net4096));
 sg13g2_buf_2 fanout4097 (.A(net4098),
    .X(net4097));
 sg13g2_buf_2 fanout4098 (.A(_07443_),
    .X(net4098));
 sg13g2_buf_2 fanout4099 (.A(_07434_),
    .X(net4099));
 sg13g2_buf_2 fanout4100 (.A(_07434_),
    .X(net4100));
 sg13g2_buf_2 fanout4101 (.A(net4102),
    .X(net4101));
 sg13g2_buf_2 fanout4102 (.A(_07420_),
    .X(net4102));
 sg13g2_buf_2 fanout4103 (.A(_07401_),
    .X(net4103));
 sg13g2_buf_2 fanout4104 (.A(_07401_),
    .X(net4104));
 sg13g2_buf_2 fanout4105 (.A(_07322_),
    .X(net4105));
 sg13g2_buf_2 fanout4106 (.A(_07322_),
    .X(net4106));
 sg13g2_buf_2 fanout4107 (.A(net4109),
    .X(net4107));
 sg13g2_buf_1 fanout4108 (.A(net4109),
    .X(net4108));
 sg13g2_buf_2 fanout4109 (.A(_06069_),
    .X(net4109));
 sg13g2_buf_2 fanout4110 (.A(net4111),
    .X(net4110));
 sg13g2_buf_4 fanout4111 (.X(net4111),
    .A(_06060_));
 sg13g2_buf_2 fanout4112 (.A(net4113),
    .X(net4112));
 sg13g2_buf_2 fanout4113 (.A(_06051_),
    .X(net4113));
 sg13g2_buf_2 fanout4114 (.A(net4116),
    .X(net4114));
 sg13g2_buf_1 fanout4115 (.A(net4116),
    .X(net4115));
 sg13g2_buf_2 fanout4116 (.A(_06042_),
    .X(net4116));
 sg13g2_buf_2 fanout4117 (.A(_06005_),
    .X(net4117));
 sg13g2_buf_2 fanout4118 (.A(_06005_),
    .X(net4118));
 sg13g2_buf_2 fanout4119 (.A(_05996_),
    .X(net4119));
 sg13g2_buf_2 fanout4120 (.A(_05996_),
    .X(net4120));
 sg13g2_buf_2 fanout4121 (.A(_05987_),
    .X(net4121));
 sg13g2_buf_2 fanout4122 (.A(_05987_),
    .X(net4122));
 sg13g2_buf_2 fanout4123 (.A(_05978_),
    .X(net4123));
 sg13g2_buf_2 fanout4124 (.A(_05978_),
    .X(net4124));
 sg13g2_buf_2 fanout4125 (.A(net4126),
    .X(net4125));
 sg13g2_buf_2 fanout4126 (.A(_05969_),
    .X(net4126));
 sg13g2_buf_2 fanout4127 (.A(net4128),
    .X(net4127));
 sg13g2_buf_2 fanout4128 (.A(_05959_),
    .X(net4128));
 sg13g2_buf_2 fanout4129 (.A(net4130),
    .X(net4129));
 sg13g2_buf_2 fanout4130 (.A(_05950_),
    .X(net4130));
 sg13g2_buf_2 fanout4131 (.A(net4132),
    .X(net4131));
 sg13g2_buf_2 fanout4132 (.A(_05941_),
    .X(net4132));
 sg13g2_buf_2 fanout4133 (.A(net4134),
    .X(net4133));
 sg13g2_buf_2 fanout4134 (.A(_05932_),
    .X(net4134));
 sg13g2_buf_2 fanout4135 (.A(_05923_),
    .X(net4135));
 sg13g2_buf_2 fanout4136 (.A(_05923_),
    .X(net4136));
 sg13g2_buf_2 fanout4137 (.A(net4138),
    .X(net4137));
 sg13g2_buf_2 fanout4138 (.A(_05914_),
    .X(net4138));
 sg13g2_buf_2 fanout4139 (.A(net4140),
    .X(net4139));
 sg13g2_buf_2 fanout4140 (.A(_05905_),
    .X(net4140));
 sg13g2_buf_2 fanout4141 (.A(_05896_),
    .X(net4141));
 sg13g2_buf_2 fanout4142 (.A(_05896_),
    .X(net4142));
 sg13g2_buf_2 fanout4143 (.A(_05887_),
    .X(net4143));
 sg13g2_buf_2 fanout4144 (.A(_05887_),
    .X(net4144));
 sg13g2_buf_2 fanout4145 (.A(net4146),
    .X(net4145));
 sg13g2_buf_2 fanout4146 (.A(_05877_),
    .X(net4146));
 sg13g2_buf_2 fanout4147 (.A(_05868_),
    .X(net4147));
 sg13g2_buf_2 fanout4148 (.A(_05868_),
    .X(net4148));
 sg13g2_buf_2 fanout4149 (.A(net4150),
    .X(net4149));
 sg13g2_buf_2 fanout4150 (.A(_05858_),
    .X(net4150));
 sg13g2_buf_2 fanout4151 (.A(net4152),
    .X(net4151));
 sg13g2_buf_4 fanout4152 (.X(net4152),
    .A(_05849_));
 sg13g2_buf_2 fanout4153 (.A(_05839_),
    .X(net4153));
 sg13g2_buf_2 fanout4154 (.A(_05839_),
    .X(net4154));
 sg13g2_buf_2 fanout4155 (.A(net4156),
    .X(net4155));
 sg13g2_buf_2 fanout4156 (.A(net4157),
    .X(net4156));
 sg13g2_buf_2 fanout4157 (.A(_05830_),
    .X(net4157));
 sg13g2_buf_2 fanout4158 (.A(_05821_),
    .X(net4158));
 sg13g2_buf_2 fanout4159 (.A(_05821_),
    .X(net4159));
 sg13g2_buf_2 fanout4160 (.A(net4161),
    .X(net4160));
 sg13g2_buf_2 fanout4161 (.A(_05812_),
    .X(net4161));
 sg13g2_buf_2 fanout4162 (.A(_05803_),
    .X(net4162));
 sg13g2_buf_2 fanout4163 (.A(_05803_),
    .X(net4163));
 sg13g2_buf_2 fanout4164 (.A(_05793_),
    .X(net4164));
 sg13g2_buf_2 fanout4165 (.A(_05793_),
    .X(net4165));
 sg13g2_buf_2 fanout4166 (.A(net4167),
    .X(net4166));
 sg13g2_buf_2 fanout4167 (.A(_05784_),
    .X(net4167));
 sg13g2_buf_2 fanout4168 (.A(_05775_),
    .X(net4168));
 sg13g2_buf_2 fanout4169 (.A(_05775_),
    .X(net4169));
 sg13g2_buf_2 fanout4170 (.A(_05763_),
    .X(net4170));
 sg13g2_buf_2 fanout4171 (.A(_05763_),
    .X(net4171));
 sg13g2_buf_2 fanout4172 (.A(_05754_),
    .X(net4172));
 sg13g2_buf_2 fanout4173 (.A(_05754_),
    .X(net4173));
 sg13g2_buf_2 fanout4174 (.A(net4175),
    .X(net4174));
 sg13g2_buf_2 fanout4175 (.A(_05745_),
    .X(net4175));
 sg13g2_buf_2 fanout4176 (.A(net4177),
    .X(net4176));
 sg13g2_buf_2 fanout4177 (.A(_05736_),
    .X(net4177));
 sg13g2_buf_2 fanout4178 (.A(net4179),
    .X(net4178));
 sg13g2_buf_2 fanout4179 (.A(_05727_),
    .X(net4179));
 sg13g2_buf_2 fanout4180 (.A(_05718_),
    .X(net4180));
 sg13g2_buf_2 fanout4181 (.A(_05718_),
    .X(net4181));
 sg13g2_buf_2 fanout4182 (.A(_05706_),
    .X(net4182));
 sg13g2_buf_2 fanout4183 (.A(_05706_),
    .X(net4183));
 sg13g2_buf_2 fanout4184 (.A(net4186),
    .X(net4184));
 sg13g2_buf_1 fanout4185 (.A(net4186),
    .X(net4185));
 sg13g2_buf_2 fanout4186 (.A(_05697_),
    .X(net4186));
 sg13g2_buf_2 fanout4187 (.A(net4188),
    .X(net4187));
 sg13g2_buf_2 fanout4188 (.A(_05688_),
    .X(net4188));
 sg13g2_buf_2 fanout4189 (.A(_05679_),
    .X(net4189));
 sg13g2_buf_2 fanout4190 (.A(_05679_),
    .X(net4190));
 sg13g2_buf_2 fanout4191 (.A(net4192),
    .X(net4191));
 sg13g2_buf_2 fanout4192 (.A(_05669_),
    .X(net4192));
 sg13g2_buf_2 fanout4193 (.A(_05659_),
    .X(net4193));
 sg13g2_buf_2 fanout4194 (.A(_05659_),
    .X(net4194));
 sg13g2_buf_2 fanout4195 (.A(net4196),
    .X(net4195));
 sg13g2_buf_2 fanout4196 (.A(_05650_),
    .X(net4196));
 sg13g2_buf_2 fanout4197 (.A(net4198),
    .X(net4197));
 sg13g2_buf_2 fanout4198 (.A(_05641_),
    .X(net4198));
 sg13g2_buf_2 fanout4199 (.A(net4200),
    .X(net4199));
 sg13g2_buf_2 fanout4200 (.A(_05600_),
    .X(net4200));
 sg13g2_buf_4 fanout4201 (.X(net4201),
    .A(net4202));
 sg13g2_buf_2 fanout4202 (.A(_05591_),
    .X(net4202));
 sg13g2_buf_2 fanout4203 (.A(net4205),
    .X(net4203));
 sg13g2_buf_1 fanout4204 (.A(net4205),
    .X(net4204));
 sg13g2_buf_2 fanout4205 (.A(_05582_),
    .X(net4205));
 sg13g2_buf_2 fanout4206 (.A(net4207),
    .X(net4206));
 sg13g2_buf_2 fanout4207 (.A(_05572_),
    .X(net4207));
 sg13g2_buf_2 fanout4208 (.A(net4209),
    .X(net4208));
 sg13g2_buf_2 fanout4209 (.A(_05563_),
    .X(net4209));
 sg13g2_buf_2 fanout4210 (.A(net4211),
    .X(net4210));
 sg13g2_buf_2 fanout4211 (.A(_05552_),
    .X(net4211));
 sg13g2_buf_2 fanout4212 (.A(_05542_),
    .X(net4212));
 sg13g2_buf_2 fanout4213 (.A(_05542_),
    .X(net4213));
 sg13g2_buf_2 fanout4214 (.A(net4216),
    .X(net4214));
 sg13g2_buf_1 fanout4215 (.A(net4216),
    .X(net4215));
 sg13g2_buf_2 fanout4216 (.A(_05533_),
    .X(net4216));
 sg13g2_buf_2 fanout4217 (.A(_05524_),
    .X(net4217));
 sg13g2_buf_2 fanout4218 (.A(_05524_),
    .X(net4218));
 sg13g2_buf_2 fanout4219 (.A(net4220),
    .X(net4219));
 sg13g2_buf_2 fanout4220 (.A(net4221),
    .X(net4220));
 sg13g2_buf_2 fanout4221 (.A(_05515_),
    .X(net4221));
 sg13g2_buf_2 fanout4222 (.A(net4223),
    .X(net4222));
 sg13g2_buf_2 fanout4223 (.A(_05506_),
    .X(net4223));
 sg13g2_buf_2 fanout4224 (.A(net4225),
    .X(net4224));
 sg13g2_buf_2 fanout4225 (.A(_05496_),
    .X(net4225));
 sg13g2_buf_2 fanout4226 (.A(_05487_),
    .X(net4226));
 sg13g2_buf_2 fanout4227 (.A(_05487_),
    .X(net4227));
 sg13g2_buf_2 fanout4228 (.A(net4229),
    .X(net4228));
 sg13g2_buf_2 fanout4229 (.A(_05478_),
    .X(net4229));
 sg13g2_buf_2 fanout4230 (.A(_05469_),
    .X(net4230));
 sg13g2_buf_2 fanout4231 (.A(_05469_),
    .X(net4231));
 sg13g2_buf_2 fanout4232 (.A(net4233),
    .X(net4232));
 sg13g2_buf_2 fanout4233 (.A(_05460_),
    .X(net4233));
 sg13g2_buf_2 fanout4234 (.A(net4235),
    .X(net4234));
 sg13g2_buf_2 fanout4235 (.A(_05450_),
    .X(net4235));
 sg13g2_buf_2 fanout4236 (.A(_05440_),
    .X(net4236));
 sg13g2_buf_2 fanout4237 (.A(_05440_),
    .X(net4237));
 sg13g2_buf_2 fanout4238 (.A(_05430_),
    .X(net4238));
 sg13g2_buf_2 fanout4239 (.A(_05430_),
    .X(net4239));
 sg13g2_buf_2 fanout4240 (.A(net4241),
    .X(net4240));
 sg13g2_buf_2 fanout4241 (.A(_05421_),
    .X(net4241));
 sg13g2_buf_2 fanout4242 (.A(_05411_),
    .X(net4242));
 sg13g2_buf_2 fanout4243 (.A(_05411_),
    .X(net4243));
 sg13g2_buf_2 fanout4244 (.A(net4245),
    .X(net4244));
 sg13g2_buf_2 fanout4245 (.A(_05401_),
    .X(net4245));
 sg13g2_buf_2 fanout4246 (.A(net4248),
    .X(net4246));
 sg13g2_buf_1 fanout4247 (.A(net4248),
    .X(net4247));
 sg13g2_buf_2 fanout4248 (.A(_05392_),
    .X(net4248));
 sg13g2_buf_4 fanout4249 (.X(net4249),
    .A(_05382_));
 sg13g2_buf_2 fanout4250 (.A(_05382_),
    .X(net4250));
 sg13g2_buf_2 fanout4251 (.A(net4252),
    .X(net4251));
 sg13g2_buf_2 fanout4252 (.A(_05372_),
    .X(net4252));
 sg13g2_buf_2 fanout4253 (.A(_05361_),
    .X(net4253));
 sg13g2_buf_2 fanout4254 (.A(_05361_),
    .X(net4254));
 sg13g2_buf_2 fanout4255 (.A(net4256),
    .X(net4255));
 sg13g2_buf_2 fanout4256 (.A(_05352_),
    .X(net4256));
 sg13g2_buf_2 fanout4257 (.A(net4258),
    .X(net4257));
 sg13g2_buf_2 fanout4258 (.A(_05343_),
    .X(net4258));
 sg13g2_buf_2 fanout4259 (.A(net4260),
    .X(net4259));
 sg13g2_buf_2 fanout4260 (.A(_05334_),
    .X(net4260));
 sg13g2_buf_2 fanout4261 (.A(net4262),
    .X(net4261));
 sg13g2_buf_2 fanout4262 (.A(_05325_),
    .X(net4262));
 sg13g2_buf_2 fanout4263 (.A(net4264),
    .X(net4263));
 sg13g2_buf_2 fanout4264 (.A(_05313_),
    .X(net4264));
 sg13g2_buf_2 fanout4265 (.A(_05276_),
    .X(net4265));
 sg13g2_buf_2 fanout4266 (.A(_05276_),
    .X(net4266));
 sg13g2_buf_2 fanout4267 (.A(_05267_),
    .X(net4267));
 sg13g2_buf_2 fanout4268 (.A(_05267_),
    .X(net4268));
 sg13g2_buf_2 fanout4269 (.A(_05258_),
    .X(net4269));
 sg13g2_buf_2 fanout4270 (.A(_05258_),
    .X(net4270));
 sg13g2_buf_2 fanout4271 (.A(_05248_),
    .X(net4271));
 sg13g2_buf_2 fanout4272 (.A(_05248_),
    .X(net4272));
 sg13g2_buf_2 fanout4273 (.A(_05239_),
    .X(net4273));
 sg13g2_buf_2 fanout4274 (.A(_05239_),
    .X(net4274));
 sg13g2_buf_2 fanout4275 (.A(net4276),
    .X(net4275));
 sg13g2_buf_2 fanout4276 (.A(_05230_),
    .X(net4276));
 sg13g2_buf_2 fanout4277 (.A(net4278),
    .X(net4277));
 sg13g2_buf_2 fanout4278 (.A(_05220_),
    .X(net4278));
 sg13g2_buf_2 fanout4279 (.A(_05211_),
    .X(net4279));
 sg13g2_buf_2 fanout4280 (.A(_05211_),
    .X(net4280));
 sg13g2_buf_2 fanout4281 (.A(_05202_),
    .X(net4281));
 sg13g2_buf_2 fanout4282 (.A(_05202_),
    .X(net4282));
 sg13g2_buf_2 fanout4283 (.A(net4284),
    .X(net4283));
 sg13g2_buf_2 fanout4284 (.A(_05193_),
    .X(net4284));
 sg13g2_buf_2 fanout4285 (.A(net4286),
    .X(net4285));
 sg13g2_buf_2 fanout4286 (.A(_05184_),
    .X(net4286));
 sg13g2_buf_2 fanout4287 (.A(_05174_),
    .X(net4287));
 sg13g2_buf_2 fanout4288 (.A(_05174_),
    .X(net4288));
 sg13g2_buf_2 fanout4289 (.A(net4290),
    .X(net4289));
 sg13g2_buf_2 fanout4290 (.A(_05165_),
    .X(net4290));
 sg13g2_buf_2 fanout4291 (.A(_05156_),
    .X(net4291));
 sg13g2_buf_2 fanout4292 (.A(_05156_),
    .X(net4292));
 sg13g2_buf_2 fanout4293 (.A(net4295),
    .X(net4293));
 sg13g2_buf_1 fanout4294 (.A(net4295),
    .X(net4294));
 sg13g2_buf_2 fanout4295 (.A(_05128_),
    .X(net4295));
 sg13g2_buf_2 fanout4296 (.A(net4297),
    .X(net4296));
 sg13g2_buf_2 fanout4297 (.A(_05118_),
    .X(net4297));
 sg13g2_buf_2 fanout4298 (.A(_05109_),
    .X(net4298));
 sg13g2_buf_2 fanout4299 (.A(_05109_),
    .X(net4299));
 sg13g2_buf_2 fanout4300 (.A(net4301),
    .X(net4300));
 sg13g2_buf_2 fanout4301 (.A(_04990_),
    .X(net4301));
 sg13g2_buf_2 fanout4302 (.A(net4303),
    .X(net4302));
 sg13g2_buf_2 fanout4303 (.A(_04980_),
    .X(net4303));
 sg13g2_buf_4 fanout4304 (.X(net4304),
    .A(_04957_));
 sg13g2_buf_2 fanout4305 (.A(_04957_),
    .X(net4305));
 sg13g2_buf_2 fanout4306 (.A(net4307),
    .X(net4306));
 sg13g2_buf_2 fanout4307 (.A(_04934_),
    .X(net4307));
 sg13g2_buf_2 fanout4308 (.A(_02726_),
    .X(net4308));
 sg13g2_buf_2 fanout4309 (.A(_02726_),
    .X(net4309));
 sg13g2_buf_2 fanout4310 (.A(net4313),
    .X(net4310));
 sg13g2_buf_2 fanout4311 (.A(net4313),
    .X(net4311));
 sg13g2_buf_1 fanout4312 (.A(net4313),
    .X(net4312));
 sg13g2_buf_1 fanout4313 (.A(_06362_),
    .X(net4313));
 sg13g2_buf_2 fanout4314 (.A(net4319),
    .X(net4314));
 sg13g2_buf_2 fanout4315 (.A(net4319),
    .X(net4315));
 sg13g2_buf_2 fanout4316 (.A(net4319),
    .X(net4316));
 sg13g2_buf_2 fanout4317 (.A(net4319),
    .X(net4317));
 sg13g2_buf_1 fanout4318 (.A(net4319),
    .X(net4318));
 sg13g2_buf_4 fanout4319 (.X(net4319),
    .A(_05127_));
 sg13g2_buf_4 fanout4320 (.X(net4320),
    .A(net4322));
 sg13g2_buf_1 fanout4321 (.A(net4322),
    .X(net4321));
 sg13g2_buf_4 fanout4322 (.X(net4322),
    .A(net4325));
 sg13g2_buf_2 fanout4323 (.A(net4325),
    .X(net4323));
 sg13g2_buf_1 fanout4324 (.A(net4325),
    .X(net4324));
 sg13g2_buf_8 fanout4325 (.A(_04956_),
    .X(net4325));
 sg13g2_buf_2 fanout4326 (.A(net4327),
    .X(net4326));
 sg13g2_buf_4 fanout4327 (.X(net4327),
    .A(_04933_));
 sg13g2_buf_2 fanout4328 (.A(net4330),
    .X(net4328));
 sg13g2_buf_2 fanout4329 (.A(net4330),
    .X(net4329));
 sg13g2_buf_4 fanout4330 (.X(net4330),
    .A(_04933_));
 sg13g2_buf_2 fanout4331 (.A(net4332),
    .X(net4331));
 sg13g2_buf_4 fanout4332 (.X(net4332),
    .A(net4335));
 sg13g2_buf_4 fanout4333 (.X(net4333),
    .A(net4335));
 sg13g2_buf_2 fanout4334 (.A(net4335),
    .X(net4334));
 sg13g2_buf_2 fanout4335 (.A(_02725_),
    .X(net4335));
 sg13g2_buf_2 fanout4336 (.A(_06198_),
    .X(net4336));
 sg13g2_buf_2 fanout4337 (.A(net4338),
    .X(net4337));
 sg13g2_buf_2 fanout4338 (.A(_07495_),
    .X(net4338));
 sg13g2_buf_2 fanout4339 (.A(_07455_),
    .X(net4339));
 sg13g2_buf_2 fanout4340 (.A(_07455_),
    .X(net4340));
 sg13g2_buf_2 fanout4341 (.A(net4345),
    .X(net4341));
 sg13g2_buf_1 fanout4342 (.A(net4345),
    .X(net4342));
 sg13g2_buf_2 fanout4343 (.A(net4345),
    .X(net4343));
 sg13g2_buf_1 fanout4344 (.A(net4345),
    .X(net4344));
 sg13g2_buf_1 fanout4345 (.A(net4346),
    .X(net4345));
 sg13g2_buf_2 fanout4346 (.A(_07334_),
    .X(net4346));
 sg13g2_buf_2 fanout4347 (.A(_06126_),
    .X(net4347));
 sg13g2_buf_4 fanout4348 (.X(net4348),
    .A(_01843_));
 sg13g2_buf_2 fanout4349 (.A(net4350),
    .X(net4349));
 sg13g2_buf_2 fanout4350 (.A(_07545_),
    .X(net4350));
 sg13g2_buf_2 fanout4351 (.A(net4352),
    .X(net4351));
 sg13g2_buf_2 fanout4352 (.A(_07543_),
    .X(net4352));
 sg13g2_buf_2 fanout4353 (.A(_07363_),
    .X(net4353));
 sg13g2_buf_4 fanout4354 (.X(net4354),
    .A(_06354_));
 sg13g2_buf_4 fanout4355 (.X(net4355),
    .A(net4357));
 sg13g2_buf_2 fanout4356 (.A(net4357),
    .X(net4356));
 sg13g2_buf_2 fanout4357 (.A(net4366),
    .X(net4357));
 sg13g2_buf_2 fanout4358 (.A(net4359),
    .X(net4358));
 sg13g2_buf_2 fanout4359 (.A(net4361),
    .X(net4359));
 sg13g2_buf_2 fanout4360 (.A(net4361),
    .X(net4360));
 sg13g2_buf_2 fanout4361 (.A(net4366),
    .X(net4361));
 sg13g2_buf_4 fanout4362 (.X(net4362),
    .A(net4366));
 sg13g2_buf_4 fanout4363 (.X(net4363),
    .A(net4366));
 sg13g2_buf_2 fanout4364 (.A(net4365),
    .X(net4364));
 sg13g2_buf_4 fanout4365 (.X(net4365),
    .A(net4366));
 sg13g2_buf_8 fanout4366 (.A(_02718_),
    .X(net4366));
 sg13g2_buf_2 fanout4367 (.A(net4368),
    .X(net4367));
 sg13g2_buf_2 fanout4368 (.A(_02601_),
    .X(net4368));
 sg13g2_buf_2 fanout4369 (.A(net4378),
    .X(net4369));
 sg13g2_buf_2 fanout4370 (.A(net4378),
    .X(net4370));
 sg13g2_buf_4 fanout4371 (.X(net4371),
    .A(net4372));
 sg13g2_buf_4 fanout4372 (.X(net4372),
    .A(net4378));
 sg13g2_buf_2 fanout4373 (.A(net4375),
    .X(net4373));
 sg13g2_buf_1 fanout4374 (.A(net4375),
    .X(net4374));
 sg13g2_buf_4 fanout4375 (.X(net4375),
    .A(net4378));
 sg13g2_buf_4 fanout4376 (.X(net4376),
    .A(net4378));
 sg13g2_buf_2 fanout4377 (.A(net4378),
    .X(net4377));
 sg13g2_buf_4 fanout4378 (.X(net4378),
    .A(_02175_));
 sg13g2_buf_4 fanout4379 (.X(net4379),
    .A(_01842_));
 sg13g2_buf_4 fanout4380 (.X(net4380),
    .A(_06351_));
 sg13g2_buf_4 fanout4381 (.X(net4381),
    .A(_06342_));
 sg13g2_buf_4 fanout4382 (.X(net4382),
    .A(_06262_));
 sg13g2_buf_2 fanout4383 (.A(_06097_),
    .X(net4383));
 sg13g2_buf_2 fanout4384 (.A(_06097_),
    .X(net4384));
 sg13g2_buf_4 fanout4385 (.X(net4385),
    .A(net4386));
 sg13g2_buf_4 fanout4386 (.X(net4386),
    .A(_03559_));
 sg13g2_buf_4 fanout4387 (.X(net4387),
    .A(_03523_));
 sg13g2_buf_2 fanout4388 (.A(net4389),
    .X(net4388));
 sg13g2_buf_2 fanout4389 (.A(net4390),
    .X(net4389));
 sg13g2_buf_2 fanout4390 (.A(_02672_),
    .X(net4390));
 sg13g2_buf_4 fanout4391 (.X(net4391),
    .A(net4392));
 sg13g2_buf_2 fanout4392 (.A(_02651_),
    .X(net4392));
 sg13g2_buf_2 fanout4393 (.A(_02648_),
    .X(net4393));
 sg13g2_buf_4 fanout4394 (.X(net4394),
    .A(_02648_));
 sg13g2_buf_2 fanout4395 (.A(net4396),
    .X(net4395));
 sg13g2_buf_2 fanout4396 (.A(net4399),
    .X(net4396));
 sg13g2_buf_4 fanout4397 (.X(net4397),
    .A(net4399));
 sg13g2_buf_2 fanout4398 (.A(net4399),
    .X(net4398));
 sg13g2_buf_2 fanout4399 (.A(_02203_),
    .X(net4399));
 sg13g2_buf_4 fanout4400 (.X(net4400),
    .A(net4405));
 sg13g2_buf_1 fanout4401 (.A(net4402),
    .X(net4401));
 sg13g2_buf_4 fanout4402 (.X(net4402),
    .A(net4405));
 sg13g2_buf_2 fanout4403 (.A(net4405),
    .X(net4403));
 sg13g2_buf_2 fanout4404 (.A(net4405),
    .X(net4404));
 sg13g2_buf_2 fanout4405 (.A(_02203_),
    .X(net4405));
 sg13g2_buf_4 fanout4406 (.X(net4406),
    .A(net4409));
 sg13g2_buf_2 fanout4407 (.A(net4409),
    .X(net4407));
 sg13g2_buf_4 fanout4408 (.X(net4408),
    .A(net4409));
 sg13g2_buf_2 fanout4409 (.A(_02144_),
    .X(net4409));
 sg13g2_buf_2 fanout4410 (.A(net4414),
    .X(net4410));
 sg13g2_buf_2 fanout4411 (.A(net4414),
    .X(net4411));
 sg13g2_buf_2 fanout4412 (.A(net4413),
    .X(net4412));
 sg13g2_buf_4 fanout4413 (.X(net4413),
    .A(net4414));
 sg13g2_buf_4 fanout4414 (.X(net4414),
    .A(_02144_));
 sg13g2_buf_4 fanout4415 (.X(net4415),
    .A(net4419));
 sg13g2_buf_2 fanout4416 (.A(net4419),
    .X(net4416));
 sg13g2_buf_2 fanout4417 (.A(net4419),
    .X(net4417));
 sg13g2_buf_1 fanout4418 (.A(net4419),
    .X(net4418));
 sg13g2_buf_2 fanout4419 (.A(_02114_),
    .X(net4419));
 sg13g2_buf_4 fanout4420 (.X(net4420),
    .A(net4424));
 sg13g2_buf_2 fanout4421 (.A(net4424),
    .X(net4421));
 sg13g2_buf_2 fanout4422 (.A(net4423),
    .X(net4422));
 sg13g2_buf_4 fanout4423 (.X(net4423),
    .A(net4424));
 sg13g2_buf_4 fanout4424 (.X(net4424),
    .A(_02114_));
 sg13g2_buf_4 fanout4425 (.X(net4425),
    .A(net4434));
 sg13g2_buf_1 fanout4426 (.A(net4434),
    .X(net4426));
 sg13g2_buf_2 fanout4427 (.A(net4428),
    .X(net4427));
 sg13g2_buf_4 fanout4428 (.X(net4428),
    .A(net4434));
 sg13g2_buf_4 fanout4429 (.X(net4429),
    .A(net4434));
 sg13g2_buf_2 fanout4430 (.A(net4434),
    .X(net4430));
 sg13g2_buf_2 fanout4431 (.A(net4433),
    .X(net4431));
 sg13g2_buf_2 fanout4432 (.A(net4433),
    .X(net4432));
 sg13g2_buf_2 fanout4433 (.A(net4434),
    .X(net4433));
 sg13g2_buf_4 fanout4434 (.X(net4434),
    .A(_02056_));
 sg13g2_buf_4 fanout4435 (.X(net4435),
    .A(net4439));
 sg13g2_buf_2 fanout4436 (.A(net4439),
    .X(net4436));
 sg13g2_buf_2 fanout4437 (.A(net4439),
    .X(net4437));
 sg13g2_buf_2 fanout4438 (.A(net4439),
    .X(net4438));
 sg13g2_buf_1 fanout4439 (.A(_07467_),
    .X(net4439));
 sg13g2_buf_2 fanout4440 (.A(net4441),
    .X(net4440));
 sg13g2_buf_4 fanout4441 (.X(net4441),
    .A(net4444));
 sg13g2_buf_2 fanout4442 (.A(net4443),
    .X(net4442));
 sg13g2_buf_4 fanout4443 (.X(net4443),
    .A(net4444));
 sg13g2_buf_2 fanout4444 (.A(_07467_),
    .X(net4444));
 sg13g2_buf_2 fanout4445 (.A(_07367_),
    .X(net4445));
 sg13g2_buf_2 fanout4446 (.A(_07362_),
    .X(net4446));
 sg13g2_buf_4 fanout4447 (.X(net4447),
    .A(_06338_));
 sg13g2_buf_4 fanout4448 (.X(net4448),
    .A(net4449));
 sg13g2_buf_2 fanout4449 (.A(net4450),
    .X(net4449));
 sg13g2_buf_4 fanout4450 (.X(net4450),
    .A(net4453));
 sg13g2_buf_4 fanout4451 (.X(net4451),
    .A(net4452));
 sg13g2_buf_4 fanout4452 (.X(net4452),
    .A(net4453));
 sg13g2_buf_8 fanout4453 (.A(_05773_),
    .X(net4453));
 sg13g2_buf_2 fanout4454 (.A(_05715_),
    .X(net4454));
 sg13g2_buf_2 fanout4455 (.A(_05715_),
    .X(net4455));
 sg13g2_buf_4 fanout4456 (.X(net4456),
    .A(net4458));
 sg13g2_buf_2 fanout4457 (.A(net4458),
    .X(net4457));
 sg13g2_buf_4 fanout4458 (.X(net4458),
    .A(net4461));
 sg13g2_buf_4 fanout4459 (.X(net4459),
    .A(net4461));
 sg13g2_buf_4 fanout4460 (.X(net4460),
    .A(net4461));
 sg13g2_buf_4 fanout4461 (.X(net4461),
    .A(_05561_));
 sg13g2_buf_4 fanout4462 (.X(net4462),
    .A(net4464));
 sg13g2_buf_2 fanout4463 (.A(net4464),
    .X(net4463));
 sg13g2_buf_4 fanout4464 (.X(net4464),
    .A(_05370_));
 sg13g2_buf_4 fanout4465 (.X(net4465),
    .A(net4467));
 sg13g2_buf_2 fanout4466 (.A(net4467),
    .X(net4466));
 sg13g2_buf_4 fanout4467 (.X(net4467),
    .A(_05370_));
 sg13g2_buf_4 fanout4468 (.X(net4468),
    .A(net4470));
 sg13g2_buf_4 fanout4469 (.X(net4469),
    .A(net4470));
 sg13g2_buf_4 fanout4470 (.X(net4470),
    .A(net4473));
 sg13g2_buf_4 fanout4471 (.X(net4471),
    .A(net4472));
 sg13g2_buf_4 fanout4472 (.X(net4472),
    .A(net4473));
 sg13g2_buf_4 fanout4473 (.X(net4473),
    .A(_05323_));
 sg13g2_buf_4 fanout4474 (.X(net4474),
    .A(net4476));
 sg13g2_buf_4 fanout4475 (.X(net4475),
    .A(net4476));
 sg13g2_buf_4 fanout4476 (.X(net4476),
    .A(net4479));
 sg13g2_buf_4 fanout4477 (.X(net4477),
    .A(net4478));
 sg13g2_buf_4 fanout4478 (.X(net4478),
    .A(net4479));
 sg13g2_buf_4 fanout4479 (.X(net4479),
    .A(_05154_));
 sg13g2_buf_4 fanout4480 (.X(net4480),
    .A(net4481));
 sg13g2_buf_2 fanout4481 (.A(_05107_),
    .X(net4481));
 sg13g2_buf_4 fanout4482 (.X(net4482),
    .A(net4485));
 sg13g2_buf_2 fanout4483 (.A(net4484),
    .X(net4483));
 sg13g2_buf_4 fanout4484 (.X(net4484),
    .A(net4485));
 sg13g2_buf_4 fanout4485 (.X(net4485),
    .A(_05107_));
 sg13g2_buf_4 fanout4486 (.X(net4486),
    .A(net4488));
 sg13g2_buf_2 fanout4487 (.A(net4488),
    .X(net4487));
 sg13g2_buf_4 fanout4488 (.X(net4488),
    .A(net4491));
 sg13g2_buf_4 fanout4489 (.X(net4489),
    .A(net4491));
 sg13g2_buf_4 fanout4490 (.X(net4490),
    .A(net4491));
 sg13g2_buf_4 fanout4491 (.X(net4491),
    .A(_04930_));
 sg13g2_buf_4 fanout4492 (.X(net4492),
    .A(_03558_));
 sg13g2_buf_4 fanout4493 (.X(net4493),
    .A(net4498));
 sg13g2_buf_1 fanout4494 (.A(net4498),
    .X(net4494));
 sg13g2_buf_2 fanout4495 (.A(net4497),
    .X(net4495));
 sg13g2_buf_1 fanout4496 (.A(net4498),
    .X(net4496));
 sg13g2_buf_2 fanout4497 (.A(net4498),
    .X(net4497));
 sg13g2_buf_2 fanout4498 (.A(_02697_),
    .X(net4498));
 sg13g2_buf_4 fanout4499 (.X(net4499),
    .A(net4502));
 sg13g2_buf_2 fanout4500 (.A(net4502),
    .X(net4500));
 sg13g2_buf_4 fanout4501 (.X(net4501),
    .A(net4502));
 sg13g2_buf_2 fanout4502 (.A(_02683_),
    .X(net4502));
 sg13g2_buf_4 fanout4503 (.X(net4503),
    .A(net4505));
 sg13g2_buf_2 fanout4504 (.A(net4505),
    .X(net4504));
 sg13g2_buf_4 fanout4505 (.X(net4505),
    .A(_02683_));
 sg13g2_buf_8 fanout4506 (.A(_02675_),
    .X(net4506));
 sg13g2_buf_4 fanout4507 (.X(net4507),
    .A(net4508));
 sg13g2_buf_4 fanout4508 (.X(net4508),
    .A(net4512));
 sg13g2_buf_4 fanout4509 (.X(net4509),
    .A(net4511));
 sg13g2_buf_2 fanout4510 (.A(net4511),
    .X(net4510));
 sg13g2_buf_4 fanout4511 (.X(net4511),
    .A(net4512));
 sg13g2_buf_2 fanout4512 (.A(net4550),
    .X(net4512));
 sg13g2_buf_4 fanout4513 (.X(net4513),
    .A(net4517));
 sg13g2_buf_4 fanout4514 (.X(net4514),
    .A(net4517));
 sg13g2_buf_4 fanout4515 (.X(net4515),
    .A(net4517));
 sg13g2_buf_2 fanout4516 (.A(net4517),
    .X(net4516));
 sg13g2_buf_2 fanout4517 (.A(net4550),
    .X(net4517));
 sg13g2_buf_4 fanout4518 (.X(net4518),
    .A(net4522));
 sg13g2_buf_4 fanout4519 (.X(net4519),
    .A(net4522));
 sg13g2_buf_4 fanout4520 (.X(net4520),
    .A(net4522));
 sg13g2_buf_2 fanout4521 (.A(net4522),
    .X(net4521));
 sg13g2_buf_2 fanout4522 (.A(net4528),
    .X(net4522));
 sg13g2_buf_4 fanout4523 (.X(net4523),
    .A(net4525));
 sg13g2_buf_4 fanout4524 (.X(net4524),
    .A(net4525));
 sg13g2_buf_4 fanout4525 (.X(net4525),
    .A(net4528));
 sg13g2_buf_4 fanout4526 (.X(net4526),
    .A(net4527));
 sg13g2_buf_4 fanout4527 (.X(net4527),
    .A(net4528));
 sg13g2_buf_2 fanout4528 (.A(net4550),
    .X(net4528));
 sg13g2_buf_4 fanout4529 (.X(net4529),
    .A(net4530));
 sg13g2_buf_4 fanout4530 (.X(net4530),
    .A(net4537));
 sg13g2_buf_4 fanout4531 (.X(net4531),
    .A(net4537));
 sg13g2_buf_4 fanout4532 (.X(net4532),
    .A(net4537));
 sg13g2_buf_4 fanout4533 (.X(net4533),
    .A(net4534));
 sg13g2_buf_4 fanout4534 (.X(net4534),
    .A(net4537));
 sg13g2_buf_4 fanout4535 (.X(net4535),
    .A(net4536));
 sg13g2_buf_4 fanout4536 (.X(net4536),
    .A(net4537));
 sg13g2_buf_2 fanout4537 (.A(net4550),
    .X(net4537));
 sg13g2_buf_4 fanout4538 (.X(net4538),
    .A(net4540));
 sg13g2_buf_4 fanout4539 (.X(net4539),
    .A(net4543));
 sg13g2_buf_2 fanout4540 (.A(net4543),
    .X(net4540));
 sg13g2_buf_4 fanout4541 (.X(net4541),
    .A(net4543));
 sg13g2_buf_4 fanout4542 (.X(net4542),
    .A(net4543));
 sg13g2_buf_2 fanout4543 (.A(net4550),
    .X(net4543));
 sg13g2_buf_4 fanout4544 (.X(net4544),
    .A(net4549));
 sg13g2_buf_4 fanout4545 (.X(net4545),
    .A(net4549));
 sg13g2_buf_4 fanout4546 (.X(net4546),
    .A(net4549));
 sg13g2_buf_2 fanout4547 (.A(net4548),
    .X(net4547));
 sg13g2_buf_4 fanout4548 (.X(net4548),
    .A(net4549));
 sg13g2_buf_2 fanout4549 (.A(net4550),
    .X(net4549));
 sg13g2_buf_8 fanout4550 (.A(_02674_),
    .X(net4550));
 sg13g2_buf_4 fanout4551 (.X(net4551),
    .A(_02650_));
 sg13g2_buf_4 fanout4552 (.X(net4552),
    .A(net4554));
 sg13g2_buf_4 fanout4553 (.X(net4553),
    .A(net4554));
 sg13g2_buf_2 fanout4554 (.A(net4557),
    .X(net4554));
 sg13g2_buf_4 fanout4555 (.X(net4555),
    .A(net4556));
 sg13g2_buf_4 fanout4556 (.X(net4556),
    .A(net4557));
 sg13g2_buf_2 fanout4557 (.A(net4596),
    .X(net4557));
 sg13g2_buf_4 fanout4558 (.X(net4558),
    .A(net4562));
 sg13g2_buf_2 fanout4559 (.A(net4562),
    .X(net4559));
 sg13g2_buf_4 fanout4560 (.X(net4560),
    .A(net4562));
 sg13g2_buf_2 fanout4561 (.A(net4562),
    .X(net4561));
 sg13g2_buf_2 fanout4562 (.A(net4596),
    .X(net4562));
 sg13g2_buf_4 fanout4563 (.X(net4563),
    .A(net4564));
 sg13g2_buf_4 fanout4564 (.X(net4564),
    .A(net4567));
 sg13g2_buf_4 fanout4565 (.X(net4565),
    .A(net4567));
 sg13g2_buf_2 fanout4566 (.A(net4567),
    .X(net4566));
 sg13g2_buf_2 fanout4567 (.A(net4573),
    .X(net4567));
 sg13g2_buf_4 fanout4568 (.X(net4568),
    .A(net4570));
 sg13g2_buf_4 fanout4569 (.X(net4569),
    .A(net4570));
 sg13g2_buf_2 fanout4570 (.A(net4573),
    .X(net4570));
 sg13g2_buf_4 fanout4571 (.X(net4571),
    .A(net4572));
 sg13g2_buf_4 fanout4572 (.X(net4572),
    .A(net4573));
 sg13g2_buf_2 fanout4573 (.A(net4596),
    .X(net4573));
 sg13g2_buf_4 fanout4574 (.X(net4574),
    .A(net4575));
 sg13g2_buf_4 fanout4575 (.X(net4575),
    .A(net4595));
 sg13g2_buf_4 fanout4576 (.X(net4576),
    .A(net4577));
 sg13g2_buf_4 fanout4577 (.X(net4577),
    .A(net4595));
 sg13g2_buf_4 fanout4578 (.X(net4578),
    .A(net4582));
 sg13g2_buf_4 fanout4579 (.X(net4579),
    .A(net4582));
 sg13g2_buf_4 fanout4580 (.X(net4580),
    .A(net4582));
 sg13g2_buf_4 fanout4581 (.X(net4581),
    .A(net4582));
 sg13g2_buf_2 fanout4582 (.A(net4595),
    .X(net4582));
 sg13g2_buf_4 fanout4583 (.X(net4583),
    .A(net4585));
 sg13g2_buf_4 fanout4584 (.X(net4584),
    .A(net4588));
 sg13g2_buf_2 fanout4585 (.A(net4588),
    .X(net4585));
 sg13g2_buf_4 fanout4586 (.X(net4586),
    .A(net4587));
 sg13g2_buf_4 fanout4587 (.X(net4587),
    .A(net4588));
 sg13g2_buf_2 fanout4588 (.A(net4595),
    .X(net4588));
 sg13g2_buf_4 fanout4589 (.X(net4589),
    .A(net4594));
 sg13g2_buf_2 fanout4590 (.A(net4594),
    .X(net4590));
 sg13g2_buf_4 fanout4591 (.X(net4591),
    .A(net4594));
 sg13g2_buf_2 fanout4592 (.A(net4593),
    .X(net4592));
 sg13g2_buf_4 fanout4593 (.X(net4593),
    .A(net4594));
 sg13g2_buf_2 fanout4594 (.A(net4595),
    .X(net4594));
 sg13g2_buf_4 fanout4595 (.X(net4595),
    .A(net4596));
 sg13g2_buf_4 fanout4596 (.X(net4596),
    .A(_02649_));
 sg13g2_buf_4 fanout4597 (.X(net4597),
    .A(_02647_));
 sg13g2_buf_4 fanout4598 (.X(net4598),
    .A(net4599));
 sg13g2_buf_4 fanout4599 (.X(net4599),
    .A(net4608));
 sg13g2_buf_4 fanout4600 (.X(net4600),
    .A(net4602));
 sg13g2_buf_1 fanout4601 (.A(net4602),
    .X(net4601));
 sg13g2_buf_4 fanout4602 (.X(net4602),
    .A(net4608));
 sg13g2_buf_4 fanout4603 (.X(net4603),
    .A(net4604));
 sg13g2_buf_4 fanout4604 (.X(net4604),
    .A(net4607));
 sg13g2_buf_4 fanout4605 (.X(net4605),
    .A(net4607));
 sg13g2_buf_4 fanout4606 (.X(net4606),
    .A(net4607));
 sg13g2_buf_2 fanout4607 (.A(net4608),
    .X(net4607));
 sg13g2_buf_2 fanout4608 (.A(_02646_),
    .X(net4608));
 sg13g2_buf_4 fanout4609 (.X(net4609),
    .A(net4610));
 sg13g2_buf_4 fanout4610 (.X(net4610),
    .A(net4613));
 sg13g2_buf_4 fanout4611 (.X(net4611),
    .A(net4613));
 sg13g2_buf_2 fanout4612 (.A(net4613),
    .X(net4612));
 sg13g2_buf_2 fanout4613 (.A(net4620),
    .X(net4613));
 sg13g2_buf_4 fanout4614 (.X(net4614),
    .A(net4617));
 sg13g2_buf_2 fanout4615 (.A(net4617),
    .X(net4615));
 sg13g2_buf_4 fanout4616 (.X(net4616),
    .A(net4617));
 sg13g2_buf_2 fanout4617 (.A(net4620),
    .X(net4617));
 sg13g2_buf_4 fanout4618 (.X(net4618),
    .A(net4620));
 sg13g2_buf_4 fanout4619 (.X(net4619),
    .A(net4620));
 sg13g2_buf_2 fanout4620 (.A(_02646_),
    .X(net4620));
 sg13g2_buf_4 fanout4621 (.X(net4621),
    .A(net4625));
 sg13g2_buf_4 fanout4622 (.X(net4622),
    .A(net4625));
 sg13g2_buf_4 fanout4623 (.X(net4623),
    .A(net4625));
 sg13g2_buf_2 fanout4624 (.A(net4625),
    .X(net4624));
 sg13g2_buf_2 fanout4625 (.A(net4642),
    .X(net4625));
 sg13g2_buf_4 fanout4626 (.X(net4626),
    .A(net4627));
 sg13g2_buf_4 fanout4627 (.X(net4627),
    .A(net4630));
 sg13g2_buf_4 fanout4628 (.X(net4628),
    .A(net4630));
 sg13g2_buf_4 fanout4629 (.X(net4629),
    .A(net4630));
 sg13g2_buf_2 fanout4630 (.A(net4642),
    .X(net4630));
 sg13g2_buf_4 fanout4631 (.X(net4631),
    .A(net4632));
 sg13g2_buf_4 fanout4632 (.X(net4632),
    .A(net4635));
 sg13g2_buf_4 fanout4633 (.X(net4633),
    .A(net4635));
 sg13g2_buf_4 fanout4634 (.X(net4634),
    .A(net4635));
 sg13g2_buf_2 fanout4635 (.A(net4642),
    .X(net4635));
 sg13g2_buf_4 fanout4636 (.X(net4636),
    .A(net4641));
 sg13g2_buf_2 fanout4637 (.A(net4641),
    .X(net4637));
 sg13g2_buf_4 fanout4638 (.X(net4638),
    .A(net4641));
 sg13g2_buf_2 fanout4639 (.A(net4640),
    .X(net4639));
 sg13g2_buf_4 fanout4640 (.X(net4640),
    .A(net4641));
 sg13g2_buf_2 fanout4641 (.A(net4642),
    .X(net4641));
 sg13g2_buf_2 fanout4642 (.A(_02646_),
    .X(net4642));
 sg13g2_buf_8 fanout4643 (.A(_02644_),
    .X(net4643));
 sg13g2_buf_4 fanout4644 (.X(net4644),
    .A(net4648));
 sg13g2_buf_2 fanout4645 (.A(net4648),
    .X(net4645));
 sg13g2_buf_4 fanout4646 (.X(net4646),
    .A(net4648));
 sg13g2_buf_2 fanout4647 (.A(net4648),
    .X(net4647));
 sg13g2_buf_2 fanout4648 (.A(net4666),
    .X(net4648));
 sg13g2_buf_2 fanout4649 (.A(net4651),
    .X(net4649));
 sg13g2_buf_4 fanout4650 (.X(net4650),
    .A(net4651));
 sg13g2_buf_2 fanout4651 (.A(net4666),
    .X(net4651));
 sg13g2_buf_4 fanout4652 (.X(net4652),
    .A(net4653));
 sg13g2_buf_4 fanout4653 (.X(net4653),
    .A(net4666));
 sg13g2_buf_4 fanout4654 (.X(net4654),
    .A(net4658));
 sg13g2_buf_1 fanout4655 (.A(net4658),
    .X(net4655));
 sg13g2_buf_4 fanout4656 (.X(net4656),
    .A(net4658));
 sg13g2_buf_4 fanout4657 (.X(net4657),
    .A(net4658));
 sg13g2_buf_2 fanout4658 (.A(net4665),
    .X(net4658));
 sg13g2_buf_4 fanout4659 (.X(net4659),
    .A(net4662));
 sg13g2_buf_2 fanout4660 (.A(net4662),
    .X(net4660));
 sg13g2_buf_4 fanout4661 (.X(net4661),
    .A(net4662));
 sg13g2_buf_2 fanout4662 (.A(net4665),
    .X(net4662));
 sg13g2_buf_4 fanout4663 (.X(net4663),
    .A(net4665));
 sg13g2_buf_1 fanout4664 (.A(net4665),
    .X(net4664));
 sg13g2_buf_2 fanout4665 (.A(net4666),
    .X(net4665));
 sg13g2_buf_2 fanout4666 (.A(_02643_),
    .X(net4666));
 sg13g2_buf_4 fanout4667 (.X(net4667),
    .A(net4670));
 sg13g2_buf_1 fanout4668 (.A(net4670),
    .X(net4668));
 sg13g2_buf_4 fanout4669 (.X(net4669),
    .A(net4670));
 sg13g2_buf_2 fanout4670 (.A(net4678),
    .X(net4670));
 sg13g2_buf_2 fanout4671 (.A(net4675),
    .X(net4671));
 sg13g2_buf_2 fanout4672 (.A(net4675),
    .X(net4672));
 sg13g2_buf_4 fanout4673 (.X(net4673),
    .A(net4675));
 sg13g2_buf_2 fanout4674 (.A(net4675),
    .X(net4674));
 sg13g2_buf_2 fanout4675 (.A(net4678),
    .X(net4675));
 sg13g2_buf_2 fanout4676 (.A(net4677),
    .X(net4676));
 sg13g2_buf_4 fanout4677 (.X(net4677),
    .A(net4678));
 sg13g2_buf_2 fanout4678 (.A(_02643_),
    .X(net4678));
 sg13g2_buf_2 fanout4679 (.A(net4683),
    .X(net4679));
 sg13g2_buf_2 fanout4680 (.A(net4683),
    .X(net4680));
 sg13g2_buf_4 fanout4681 (.X(net4681),
    .A(net4683));
 sg13g2_buf_2 fanout4682 (.A(net4683),
    .X(net4682));
 sg13g2_buf_2 fanout4683 (.A(net4690),
    .X(net4683));
 sg13g2_buf_4 fanout4684 (.X(net4684),
    .A(net4687));
 sg13g2_buf_4 fanout4685 (.X(net4685),
    .A(net4687));
 sg13g2_buf_2 fanout4686 (.A(net4687),
    .X(net4686));
 sg13g2_buf_2 fanout4687 (.A(net4690),
    .X(net4687));
 sg13g2_buf_4 fanout4688 (.X(net4688),
    .A(net4690));
 sg13g2_buf_2 fanout4689 (.A(net4690),
    .X(net4689));
 sg13g2_buf_4 fanout4690 (.X(net4690),
    .A(_02643_));
 sg13g2_buf_2 fanout4691 (.A(_02528_),
    .X(net4691));
 sg13g2_buf_2 fanout4692 (.A(_02528_),
    .X(net4692));
 sg13g2_buf_4 fanout4693 (.X(net4693),
    .A(net4694));
 sg13g2_buf_4 fanout4694 (.X(net4694),
    .A(net4702));
 sg13g2_buf_4 fanout4695 (.X(net4695),
    .A(net4702));
 sg13g2_buf_1 fanout4696 (.A(net4702),
    .X(net4696));
 sg13g2_buf_2 fanout4697 (.A(net4698),
    .X(net4697));
 sg13g2_buf_4 fanout4698 (.X(net4698),
    .A(net4701));
 sg13g2_buf_2 fanout4699 (.A(net4700),
    .X(net4699));
 sg13g2_buf_4 fanout4700 (.X(net4700),
    .A(net4701));
 sg13g2_buf_2 fanout4701 (.A(net4702),
    .X(net4701));
 sg13g2_buf_2 fanout4702 (.A(_02085_),
    .X(net4702));
 sg13g2_buf_4 fanout4703 (.X(net4703),
    .A(net4704));
 sg13g2_buf_4 fanout4704 (.X(net4704),
    .A(_01781_));
 sg13g2_buf_2 fanout4705 (.A(_01781_),
    .X(net4705));
 sg13g2_buf_4 fanout4706 (.X(net4706),
    .A(net4707));
 sg13g2_buf_4 fanout4707 (.X(net4707),
    .A(_01780_));
 sg13g2_buf_2 fanout4708 (.A(_07366_),
    .X(net4708));
 sg13g2_buf_2 fanout4709 (.A(net4710),
    .X(net4709));
 sg13g2_buf_2 fanout4710 (.A(_06350_),
    .X(net4710));
 sg13g2_buf_2 fanout4711 (.A(net4712),
    .X(net4711));
 sg13g2_buf_1 fanout4712 (.A(_06349_),
    .X(net4712));
 sg13g2_buf_2 fanout4713 (.A(net4714),
    .X(net4713));
 sg13g2_buf_2 fanout4714 (.A(net4715),
    .X(net4714));
 sg13g2_buf_4 fanout4715 (.X(net4715),
    .A(_06084_));
 sg13g2_buf_2 fanout4716 (.A(_03969_),
    .X(net4716));
 sg13g2_buf_1 fanout4717 (.A(_03969_),
    .X(net4717));
 sg13g2_buf_2 fanout4718 (.A(net4720),
    .X(net4718));
 sg13g2_buf_2 fanout4719 (.A(net4720),
    .X(net4719));
 sg13g2_buf_2 fanout4720 (.A(net4721),
    .X(net4720));
 sg13g2_buf_2 fanout4721 (.A(net4722),
    .X(net4721));
 sg13g2_buf_2 fanout4722 (.A(_03550_),
    .X(net4722));
 sg13g2_buf_2 fanout4723 (.A(net4728),
    .X(net4723));
 sg13g2_buf_2 fanout4724 (.A(net4726),
    .X(net4724));
 sg13g2_buf_2 fanout4725 (.A(net4726),
    .X(net4725));
 sg13g2_buf_2 fanout4726 (.A(net4727),
    .X(net4726));
 sg13g2_buf_2 fanout4727 (.A(net4728),
    .X(net4727));
 sg13g2_buf_2 fanout4728 (.A(_03550_),
    .X(net4728));
 sg13g2_buf_2 fanout4729 (.A(_02883_),
    .X(net4729));
 sg13g2_buf_1 fanout4730 (.A(_02883_),
    .X(net4730));
 sg13g2_buf_4 fanout4731 (.X(net4731),
    .A(net4732));
 sg13g2_buf_4 fanout4732 (.X(net4732),
    .A(_02777_));
 sg13g2_buf_4 fanout4733 (.X(net4733),
    .A(net4734));
 sg13g2_buf_4 fanout4734 (.X(net4734),
    .A(_02776_));
 sg13g2_buf_2 fanout4735 (.A(net4737),
    .X(net4735));
 sg13g2_buf_2 fanout4736 (.A(net4737),
    .X(net4736));
 sg13g2_buf_2 fanout4737 (.A(_02759_),
    .X(net4737));
 sg13g2_buf_4 fanout4738 (.X(net4738),
    .A(net4739));
 sg13g2_buf_2 fanout4739 (.A(_02759_),
    .X(net4739));
 sg13g2_buf_2 fanout4740 (.A(_03819_),
    .X(net4740));
 sg13g2_buf_2 fanout4741 (.A(net4744),
    .X(net4741));
 sg13g2_buf_2 fanout4742 (.A(net4744),
    .X(net4742));
 sg13g2_buf_1 fanout4743 (.A(net4744),
    .X(net4743));
 sg13g2_buf_4 fanout4744 (.X(net4744),
    .A(_03553_));
 sg13g2_buf_2 fanout4745 (.A(net4746),
    .X(net4745));
 sg13g2_buf_1 fanout4746 (.A(net4747),
    .X(net4746));
 sg13g2_buf_1 fanout4747 (.A(_03541_),
    .X(net4747));
 sg13g2_buf_4 fanout4748 (.X(net4748),
    .A(net4750));
 sg13g2_buf_2 fanout4749 (.A(net4750),
    .X(net4749));
 sg13g2_buf_4 fanout4750 (.X(net4750),
    .A(net4754));
 sg13g2_buf_2 fanout4751 (.A(net4752),
    .X(net4751));
 sg13g2_buf_2 fanout4752 (.A(net4753),
    .X(net4752));
 sg13g2_buf_1 fanout4753 (.A(net4754),
    .X(net4753));
 sg13g2_buf_2 fanout4754 (.A(_03497_),
    .X(net4754));
 sg13g2_buf_2 fanout4755 (.A(net4756),
    .X(net4755));
 sg13g2_buf_4 fanout4756 (.X(net4756),
    .A(net4760));
 sg13g2_buf_2 fanout4757 (.A(net4760),
    .X(net4757));
 sg13g2_buf_2 fanout4758 (.A(net4759),
    .X(net4758));
 sg13g2_buf_2 fanout4759 (.A(net4760),
    .X(net4759));
 sg13g2_buf_2 fanout4760 (.A(_03496_),
    .X(net4760));
 sg13g2_buf_2 fanout4761 (.A(net4764),
    .X(net4761));
 sg13g2_buf_2 fanout4762 (.A(net4763),
    .X(net4762));
 sg13g2_buf_2 fanout4763 (.A(net4764),
    .X(net4763));
 sg13g2_buf_4 fanout4764 (.X(net4764),
    .A(_03460_));
 sg13g2_buf_2 fanout4765 (.A(net4766),
    .X(net4765));
 sg13g2_buf_2 fanout4766 (.A(_03459_),
    .X(net4766));
 sg13g2_buf_4 fanout4767 (.X(net4767),
    .A(net4768));
 sg13g2_buf_4 fanout4768 (.X(net4768),
    .A(_03410_));
 sg13g2_buf_2 fanout4769 (.A(net4770),
    .X(net4769));
 sg13g2_buf_2 fanout4770 (.A(_03409_),
    .X(net4770));
 sg13g2_buf_4 fanout4771 (.X(net4771),
    .A(net4773));
 sg13g2_buf_1 fanout4772 (.A(net4773),
    .X(net4772));
 sg13g2_buf_1 fanout4773 (.A(net4774),
    .X(net4773));
 sg13g2_buf_2 fanout4774 (.A(_03319_),
    .X(net4774));
 sg13g2_buf_2 fanout4775 (.A(net4777),
    .X(net4775));
 sg13g2_buf_1 fanout4776 (.A(net4777),
    .X(net4776));
 sg13g2_buf_2 fanout4777 (.A(net4778),
    .X(net4777));
 sg13g2_buf_2 fanout4778 (.A(net4785),
    .X(net4778));
 sg13g2_buf_2 fanout4779 (.A(net4780),
    .X(net4779));
 sg13g2_buf_2 fanout4780 (.A(net4785),
    .X(net4780));
 sg13g2_buf_2 fanout4781 (.A(net4783),
    .X(net4781));
 sg13g2_buf_2 fanout4782 (.A(net4783),
    .X(net4782));
 sg13g2_buf_2 fanout4783 (.A(net4784),
    .X(net4783));
 sg13g2_buf_2 fanout4784 (.A(net4785),
    .X(net4784));
 sg13g2_buf_4 fanout4785 (.X(net4785),
    .A(_03123_));
 sg13g2_buf_4 fanout4786 (.X(net4786),
    .A(net4788));
 sg13g2_buf_2 fanout4787 (.A(net4788),
    .X(net4787));
 sg13g2_buf_2 fanout4788 (.A(_02783_),
    .X(net4788));
 sg13g2_buf_2 fanout4789 (.A(_06111_),
    .X(net4789));
 sg13g2_buf_2 fanout4790 (.A(_06107_),
    .X(net4790));
 sg13g2_buf_2 fanout4791 (.A(net4792),
    .X(net4791));
 sg13g2_buf_2 fanout4792 (.A(_06080_),
    .X(net4792));
 sg13g2_buf_2 fanout4793 (.A(_05610_),
    .X(net4793));
 sg13g2_buf_4 fanout4794 (.X(net4794),
    .A(_05610_));
 sg13g2_buf_2 fanout4795 (.A(net4797),
    .X(net4795));
 sg13g2_buf_4 fanout4796 (.X(net4796),
    .A(net4797));
 sg13g2_buf_2 fanout4797 (.A(_05153_),
    .X(net4797));
 sg13g2_buf_2 fanout4798 (.A(_05153_),
    .X(net4798));
 sg13g2_buf_1 fanout4799 (.A(_05153_),
    .X(net4799));
 sg13g2_buf_2 fanout4800 (.A(net4804),
    .X(net4800));
 sg13g2_buf_2 fanout4801 (.A(net4804),
    .X(net4801));
 sg13g2_buf_2 fanout4802 (.A(net4804),
    .X(net4802));
 sg13g2_buf_2 fanout4803 (.A(net4804),
    .X(net4803));
 sg13g2_buf_4 fanout4804 (.X(net4804),
    .A(_05147_));
 sg13g2_buf_4 fanout4805 (.X(net4805),
    .A(net4807));
 sg13g2_buf_2 fanout4806 (.A(net4807),
    .X(net4806));
 sg13g2_buf_2 fanout4807 (.A(_05141_),
    .X(net4807));
 sg13g2_buf_2 fanout4808 (.A(net4809),
    .X(net4808));
 sg13g2_buf_2 fanout4809 (.A(_05141_),
    .X(net4809));
 sg13g2_buf_2 fanout4810 (.A(_05135_),
    .X(net4810));
 sg13g2_buf_2 fanout4811 (.A(_05135_),
    .X(net4811));
 sg13g2_buf_2 fanout4812 (.A(net4813),
    .X(net4812));
 sg13g2_buf_1 fanout4813 (.A(net4814),
    .X(net4813));
 sg13g2_buf_2 fanout4814 (.A(_05135_),
    .X(net4814));
 sg13g2_buf_2 fanout4815 (.A(net4816),
    .X(net4815));
 sg13g2_buf_4 fanout4816 (.X(net4816),
    .A(_04978_));
 sg13g2_buf_4 fanout4817 (.X(net4817),
    .A(net4819));
 sg13g2_buf_1 fanout4818 (.A(net4819),
    .X(net4818));
 sg13g2_buf_2 fanout4819 (.A(_04978_),
    .X(net4819));
 sg13g2_buf_4 fanout4820 (.X(net4820),
    .A(net4821));
 sg13g2_buf_4 fanout4821 (.X(net4821),
    .A(net4824));
 sg13g2_buf_4 fanout4822 (.X(net4822),
    .A(net4824));
 sg13g2_buf_4 fanout4823 (.X(net4823),
    .A(net4824));
 sg13g2_buf_4 fanout4824 (.X(net4824),
    .A(_04975_));
 sg13g2_buf_4 fanout4825 (.X(net4825),
    .A(net4830));
 sg13g2_buf_2 fanout4826 (.A(net4830),
    .X(net4826));
 sg13g2_buf_4 fanout4827 (.X(net4827),
    .A(net4828));
 sg13g2_buf_2 fanout4828 (.A(net4830),
    .X(net4828));
 sg13g2_buf_2 fanout4829 (.A(net4830),
    .X(net4829));
 sg13g2_buf_2 fanout4830 (.A(_04972_),
    .X(net4830));
 sg13g2_buf_4 fanout4831 (.X(net4831),
    .A(net4833));
 sg13g2_buf_2 fanout4832 (.A(net4833),
    .X(net4832));
 sg13g2_buf_4 fanout4833 (.X(net4833),
    .A(net4836));
 sg13g2_buf_2 fanout4834 (.A(net4836),
    .X(net4834));
 sg13g2_buf_1 fanout4835 (.A(net4836),
    .X(net4835));
 sg13g2_buf_8 fanout4836 (.A(_04969_),
    .X(net4836));
 sg13g2_buf_4 fanout4837 (.X(net4837),
    .A(_04966_));
 sg13g2_buf_1 fanout4838 (.A(_04966_),
    .X(net4838));
 sg13g2_buf_2 fanout4839 (.A(net4841),
    .X(net4839));
 sg13g2_buf_4 fanout4840 (.X(net4840),
    .A(net4841));
 sg13g2_buf_2 fanout4841 (.A(_04966_),
    .X(net4841));
 sg13g2_buf_4 fanout4842 (.X(net4842),
    .A(net4844));
 sg13g2_buf_1 fanout4843 (.A(net4844),
    .X(net4843));
 sg13g2_buf_2 fanout4844 (.A(_04963_),
    .X(net4844));
 sg13g2_buf_4 fanout4845 (.X(net4845),
    .A(_04963_));
 sg13g2_buf_4 fanout4846 (.X(net4846),
    .A(_04963_));
 sg13g2_buf_4 fanout4847 (.X(net4847),
    .A(net4852));
 sg13g2_buf_1 fanout4848 (.A(net4852),
    .X(net4848));
 sg13g2_buf_4 fanout4849 (.X(net4849),
    .A(net4852));
 sg13g2_buf_2 fanout4850 (.A(net4852),
    .X(net4850));
 sg13g2_buf_4 fanout4851 (.X(net4851),
    .A(net4852));
 sg13g2_buf_8 fanout4852 (.A(_04960_),
    .X(net4852));
 sg13g2_buf_4 fanout4853 (.X(net4853),
    .A(net4855));
 sg13g2_buf_1 fanout4854 (.A(net4855),
    .X(net4854));
 sg13g2_buf_4 fanout4855 (.X(net4855),
    .A(net4858));
 sg13g2_buf_4 fanout4856 (.X(net4856),
    .A(net4858));
 sg13g2_buf_1 fanout4857 (.A(net4858),
    .X(net4857));
 sg13g2_buf_4 fanout4858 (.X(net4858),
    .A(_04952_));
 sg13g2_buf_2 fanout4859 (.A(net4861),
    .X(net4859));
 sg13g2_buf_1 fanout4860 (.A(net4861),
    .X(net4860));
 sg13g2_buf_2 fanout4861 (.A(_04948_),
    .X(net4861));
 sg13g2_buf_4 fanout4862 (.X(net4862),
    .A(_04948_));
 sg13g2_buf_4 fanout4863 (.X(net4863),
    .A(_04948_));
 sg13g2_buf_4 fanout4864 (.X(net4864),
    .A(net4865));
 sg13g2_buf_4 fanout4865 (.X(net4865),
    .A(_04944_));
 sg13g2_buf_2 fanout4866 (.A(net4868),
    .X(net4866));
 sg13g2_buf_1 fanout4867 (.A(net4868),
    .X(net4867));
 sg13g2_buf_4 fanout4868 (.X(net4868),
    .A(_04944_));
 sg13g2_buf_4 fanout4869 (.X(net4869),
    .A(_04940_));
 sg13g2_buf_2 fanout4870 (.A(_04940_),
    .X(net4870));
 sg13g2_buf_2 fanout4871 (.A(net4873),
    .X(net4871));
 sg13g2_buf_1 fanout4872 (.A(net4873),
    .X(net4872));
 sg13g2_buf_4 fanout4873 (.X(net4873),
    .A(_04940_));
 sg13g2_buf_2 fanout4874 (.A(net4875),
    .X(net4874));
 sg13g2_buf_4 fanout4875 (.X(net4875),
    .A(_04936_));
 sg13g2_buf_4 fanout4876 (.X(net4876),
    .A(_04936_));
 sg13g2_buf_4 fanout4877 (.X(net4877),
    .A(_04936_));
 sg13g2_buf_2 fanout4878 (.A(net4879),
    .X(net4878));
 sg13g2_buf_2 fanout4879 (.A(_03532_),
    .X(net4879));
 sg13g2_buf_4 fanout4880 (.X(net4880),
    .A(_03515_));
 sg13g2_buf_1 fanout4881 (.A(_03515_),
    .X(net4881));
 sg13g2_buf_2 fanout4882 (.A(_03514_),
    .X(net4882));
 sg13g2_buf_2 fanout4883 (.A(_03506_),
    .X(net4883));
 sg13g2_buf_4 fanout4884 (.X(net4884),
    .A(_03402_));
 sg13g2_buf_2 fanout4885 (.A(net4887),
    .X(net4885));
 sg13g2_buf_1 fanout4886 (.A(net4887),
    .X(net4886));
 sg13g2_buf_1 fanout4887 (.A(_03318_),
    .X(net4887));
 sg13g2_buf_2 fanout4888 (.A(net4889),
    .X(net4888));
 sg13g2_buf_1 fanout4889 (.A(net4890),
    .X(net4889));
 sg13g2_buf_2 fanout4890 (.A(net4891),
    .X(net4890));
 sg13g2_buf_2 fanout4891 (.A(_03318_),
    .X(net4891));
 sg13g2_buf_2 fanout4892 (.A(net4893),
    .X(net4892));
 sg13g2_buf_2 fanout4893 (.A(net4894),
    .X(net4893));
 sg13g2_buf_2 fanout4894 (.A(_03152_),
    .X(net4894));
 sg13g2_buf_4 fanout4895 (.X(net4895),
    .A(_03151_));
 sg13g2_buf_2 fanout4896 (.A(net4897),
    .X(net4896));
 sg13g2_buf_2 fanout4897 (.A(net4898),
    .X(net4897));
 sg13g2_buf_2 fanout4898 (.A(net4900),
    .X(net4898));
 sg13g2_buf_2 fanout4899 (.A(net4900),
    .X(net4899));
 sg13g2_buf_1 fanout4900 (.A(_03137_),
    .X(net4900));
 sg13g2_buf_2 fanout4901 (.A(net4903),
    .X(net4901));
 sg13g2_buf_1 fanout4902 (.A(net4903),
    .X(net4902));
 sg13g2_buf_2 fanout4903 (.A(_03137_),
    .X(net4903));
 sg13g2_buf_2 fanout4904 (.A(net4905),
    .X(net4904));
 sg13g2_buf_2 fanout4905 (.A(net4911),
    .X(net4905));
 sg13g2_buf_2 fanout4906 (.A(net4907),
    .X(net4906));
 sg13g2_buf_2 fanout4907 (.A(net4910),
    .X(net4907));
 sg13g2_buf_2 fanout4908 (.A(net4909),
    .X(net4908));
 sg13g2_buf_1 fanout4909 (.A(net4910),
    .X(net4909));
 sg13g2_buf_2 fanout4910 (.A(net4911),
    .X(net4910));
 sg13g2_buf_2 fanout4911 (.A(_03136_),
    .X(net4911));
 sg13g2_buf_2 fanout4912 (.A(net4913),
    .X(net4912));
 sg13g2_buf_1 fanout4913 (.A(net4923),
    .X(net4913));
 sg13g2_buf_2 fanout4914 (.A(net4923),
    .X(net4914));
 sg13g2_buf_2 fanout4915 (.A(net4923),
    .X(net4915));
 sg13g2_buf_2 fanout4916 (.A(net4922),
    .X(net4916));
 sg13g2_buf_1 fanout4917 (.A(net4922),
    .X(net4917));
 sg13g2_buf_2 fanout4918 (.A(net4922),
    .X(net4918));
 sg13g2_buf_1 fanout4919 (.A(net4922),
    .X(net4919));
 sg13g2_buf_2 fanout4920 (.A(net4921),
    .X(net4920));
 sg13g2_buf_2 fanout4921 (.A(net4922),
    .X(net4921));
 sg13g2_buf_2 fanout4922 (.A(net4923),
    .X(net4922));
 sg13g2_buf_2 fanout4923 (.A(_03132_),
    .X(net4923));
 sg13g2_buf_2 fanout4924 (.A(net4926),
    .X(net4924));
 sg13g2_buf_1 fanout4925 (.A(net4926),
    .X(net4925));
 sg13g2_buf_2 fanout4926 (.A(net4927),
    .X(net4926));
 sg13g2_buf_2 fanout4927 (.A(net4934),
    .X(net4927));
 sg13g2_buf_2 fanout4928 (.A(net4929),
    .X(net4928));
 sg13g2_buf_2 fanout4929 (.A(net4933),
    .X(net4929));
 sg13g2_buf_2 fanout4930 (.A(net4931),
    .X(net4930));
 sg13g2_buf_1 fanout4931 (.A(net4932),
    .X(net4931));
 sg13g2_buf_2 fanout4932 (.A(net4933),
    .X(net4932));
 sg13g2_buf_2 fanout4933 (.A(net4934),
    .X(net4933));
 sg13g2_buf_2 fanout4934 (.A(_03131_),
    .X(net4934));
 sg13g2_buf_2 fanout4935 (.A(net4936),
    .X(net4935));
 sg13g2_buf_2 fanout4936 (.A(net4939),
    .X(net4936));
 sg13g2_buf_2 fanout4937 (.A(net4939),
    .X(net4937));
 sg13g2_buf_2 fanout4938 (.A(net4939),
    .X(net4938));
 sg13g2_buf_2 fanout4939 (.A(_03128_),
    .X(net4939));
 sg13g2_buf_2 fanout4940 (.A(net4944),
    .X(net4940));
 sg13g2_buf_2 fanout4941 (.A(net4942),
    .X(net4941));
 sg13g2_buf_2 fanout4942 (.A(net4943),
    .X(net4942));
 sg13g2_buf_2 fanout4943 (.A(net4944),
    .X(net4943));
 sg13g2_buf_2 fanout4944 (.A(_03127_),
    .X(net4944));
 sg13g2_buf_2 fanout4945 (.A(_03127_),
    .X(net4945));
 sg13g2_buf_2 fanout4946 (.A(net4947),
    .X(net4946));
 sg13g2_buf_2 fanout4947 (.A(net4948),
    .X(net4947));
 sg13g2_buf_2 fanout4948 (.A(_03122_),
    .X(net4948));
 sg13g2_buf_2 fanout4949 (.A(net4951),
    .X(net4949));
 sg13g2_buf_2 fanout4950 (.A(net4951),
    .X(net4950));
 sg13g2_buf_2 fanout4951 (.A(_03122_),
    .X(net4951));
 sg13g2_buf_2 fanout4952 (.A(net4956),
    .X(net4952));
 sg13g2_buf_2 fanout4953 (.A(net4956),
    .X(net4953));
 sg13g2_buf_2 fanout4954 (.A(net4955),
    .X(net4954));
 sg13g2_buf_1 fanout4955 (.A(net4956),
    .X(net4955));
 sg13g2_buf_2 fanout4956 (.A(_03122_),
    .X(net4956));
 sg13g2_buf_2 fanout4957 (.A(_02782_),
    .X(net4957));
 sg13g2_buf_4 fanout4958 (.X(net4958),
    .A(net4961));
 sg13g2_buf_2 fanout4959 (.A(net4960),
    .X(net4959));
 sg13g2_buf_2 fanout4960 (.A(net4961),
    .X(net4960));
 sg13g2_buf_2 fanout4961 (.A(net4970),
    .X(net4961));
 sg13g2_buf_2 fanout4962 (.A(net4964),
    .X(net4962));
 sg13g2_buf_1 fanout4963 (.A(net4964),
    .X(net4963));
 sg13g2_buf_2 fanout4964 (.A(net4965),
    .X(net4964));
 sg13g2_buf_2 fanout4965 (.A(net4970),
    .X(net4965));
 sg13g2_buf_2 fanout4966 (.A(net4967),
    .X(net4966));
 sg13g2_buf_2 fanout4967 (.A(net4970),
    .X(net4967));
 sg13g2_buf_2 fanout4968 (.A(net4970),
    .X(net4968));
 sg13g2_buf_1 fanout4969 (.A(net4970),
    .X(net4969));
 sg13g2_buf_4 fanout4970 (.X(net4970),
    .A(_02757_));
 sg13g2_buf_2 fanout4971 (.A(net4973),
    .X(net4971));
 sg13g2_buf_2 fanout4972 (.A(net4973),
    .X(net4972));
 sg13g2_buf_2 fanout4973 (.A(net4974),
    .X(net4973));
 sg13g2_buf_2 fanout4974 (.A(_02756_),
    .X(net4974));
 sg13g2_buf_2 fanout4975 (.A(net4977),
    .X(net4975));
 sg13g2_buf_2 fanout4976 (.A(net4977),
    .X(net4976));
 sg13g2_buf_4 fanout4977 (.X(net4977),
    .A(_02756_));
 sg13g2_buf_2 fanout4978 (.A(net4980),
    .X(net4978));
 sg13g2_buf_1 fanout4979 (.A(net4980),
    .X(net4979));
 sg13g2_buf_2 fanout4980 (.A(_02750_),
    .X(net4980));
 sg13g2_buf_4 fanout4981 (.X(net4981),
    .A(_02750_));
 sg13g2_buf_4 fanout4982 (.X(net4982),
    .A(_02750_));
 sg13g2_buf_4 fanout4983 (.X(net4983),
    .A(net4984));
 sg13g2_buf_4 fanout4984 (.X(net4984),
    .A(net4987));
 sg13g2_buf_2 fanout4985 (.A(net4986),
    .X(net4985));
 sg13g2_buf_2 fanout4986 (.A(net4987),
    .X(net4986));
 sg13g2_buf_4 fanout4987 (.X(net4987),
    .A(_02744_));
 sg13g2_buf_2 fanout4988 (.A(net4989),
    .X(net4988));
 sg13g2_buf_2 fanout4989 (.A(net4990),
    .X(net4989));
 sg13g2_buf_2 fanout4990 (.A(_02738_),
    .X(net4990));
 sg13g2_buf_2 fanout4991 (.A(_02738_),
    .X(net4991));
 sg13g2_buf_1 fanout4992 (.A(_02738_),
    .X(net4992));
 sg13g2_buf_2 fanout4993 (.A(net4994),
    .X(net4993));
 sg13g2_buf_4 fanout4994 (.X(net4994),
    .A(_02732_));
 sg13g2_buf_2 fanout4995 (.A(net4996),
    .X(net4995));
 sg13g2_buf_2 fanout4996 (.A(net4997),
    .X(net4996));
 sg13g2_buf_4 fanout4997 (.X(net4997),
    .A(_02732_));
 sg13g2_buf_2 fanout4998 (.A(net4999),
    .X(net4998));
 sg13g2_buf_2 fanout4999 (.A(_06268_),
    .X(net4999));
 sg13g2_buf_2 fanout5000 (.A(net5001),
    .X(net5000));
 sg13g2_buf_2 fanout5001 (.A(_06112_),
    .X(net5001));
 sg13g2_buf_2 fanout5002 (.A(net5004),
    .X(net5002));
 sg13g2_buf_1 fanout5003 (.A(net5004),
    .X(net5003));
 sg13g2_buf_2 fanout5004 (.A(_06078_),
    .X(net5004));
 sg13g2_buf_4 fanout5005 (.X(net5005),
    .A(net5009));
 sg13g2_buf_4 fanout5006 (.X(net5006),
    .A(net5009));
 sg13g2_buf_4 fanout5007 (.X(net5007),
    .A(net5008));
 sg13g2_buf_4 fanout5008 (.X(net5008),
    .A(net5009));
 sg13g2_buf_2 fanout5009 (.A(_05150_),
    .X(net5009));
 sg13g2_buf_2 fanout5010 (.A(_05144_),
    .X(net5010));
 sg13g2_buf_2 fanout5011 (.A(_05144_),
    .X(net5011));
 sg13g2_buf_2 fanout5012 (.A(net5013),
    .X(net5012));
 sg13g2_buf_2 fanout5013 (.A(net5014),
    .X(net5013));
 sg13g2_buf_2 fanout5014 (.A(_05144_),
    .X(net5014));
 sg13g2_buf_4 fanout5015 (.X(net5015),
    .A(net5017));
 sg13g2_buf_2 fanout5016 (.A(net5017),
    .X(net5016));
 sg13g2_buf_2 fanout5017 (.A(_05138_),
    .X(net5017));
 sg13g2_buf_4 fanout5018 (.X(net5018),
    .A(net5019));
 sg13g2_buf_4 fanout5019 (.X(net5019),
    .A(_05138_));
 sg13g2_buf_2 fanout5020 (.A(net5022),
    .X(net5020));
 sg13g2_buf_1 fanout5021 (.A(net5022),
    .X(net5021));
 sg13g2_buf_4 fanout5022 (.X(net5022),
    .A(net5025));
 sg13g2_buf_4 fanout5023 (.X(net5023),
    .A(net5025));
 sg13g2_buf_1 fanout5024 (.A(net5025),
    .X(net5024));
 sg13g2_buf_4 fanout5025 (.X(net5025),
    .A(_05132_));
 sg13g2_buf_4 fanout5026 (.X(net5026),
    .A(net5027));
 sg13g2_buf_4 fanout5027 (.X(net5027),
    .A(_04946_));
 sg13g2_buf_4 fanout5028 (.X(net5028),
    .A(_04946_));
 sg13g2_buf_4 fanout5029 (.X(net5029),
    .A(_04946_));
 sg13g2_buf_4 fanout5030 (.X(net5030),
    .A(net5031));
 sg13g2_buf_4 fanout5031 (.X(net5031),
    .A(_04942_));
 sg13g2_buf_4 fanout5032 (.X(net5032),
    .A(net5034));
 sg13g2_buf_1 fanout5033 (.A(net5034),
    .X(net5033));
 sg13g2_buf_4 fanout5034 (.X(net5034),
    .A(_04942_));
 sg13g2_buf_4 fanout5035 (.X(net5035),
    .A(net5037));
 sg13g2_buf_1 fanout5036 (.A(net5037),
    .X(net5036));
 sg13g2_buf_2 fanout5037 (.A(_04938_),
    .X(net5037));
 sg13g2_buf_4 fanout5038 (.X(net5038),
    .A(net5040));
 sg13g2_buf_1 fanout5039 (.A(net5040),
    .X(net5039));
 sg13g2_buf_4 fanout5040 (.X(net5040),
    .A(_04938_));
 sg13g2_buf_4 fanout5041 (.X(net5041),
    .A(net5042));
 sg13g2_buf_4 fanout5042 (.X(net5042),
    .A(_04928_));
 sg13g2_buf_2 fanout5043 (.A(net5045),
    .X(net5043));
 sg13g2_buf_1 fanout5044 (.A(net5045),
    .X(net5044));
 sg13g2_buf_4 fanout5045 (.X(net5045),
    .A(_04928_));
 sg13g2_buf_4 fanout5046 (.X(net5046),
    .A(net5049));
 sg13g2_buf_4 fanout5047 (.X(net5047),
    .A(net5049));
 sg13g2_buf_4 fanout5048 (.X(net5048),
    .A(net5049));
 sg13g2_buf_4 fanout5049 (.X(net5049),
    .A(_03565_));
 sg13g2_buf_4 fanout5050 (.X(net5050),
    .A(net5051));
 sg13g2_buf_2 fanout5051 (.A(net5053),
    .X(net5051));
 sg13g2_buf_4 fanout5052 (.X(net5052),
    .A(net5053));
 sg13g2_buf_2 fanout5053 (.A(_03563_),
    .X(net5053));
 sg13g2_buf_2 fanout5054 (.A(net5055),
    .X(net5054));
 sg13g2_buf_2 fanout5055 (.A(net5058),
    .X(net5055));
 sg13g2_buf_2 fanout5056 (.A(net5058),
    .X(net5056));
 sg13g2_buf_2 fanout5057 (.A(net5058),
    .X(net5057));
 sg13g2_buf_2 fanout5058 (.A(_03563_),
    .X(net5058));
 sg13g2_buf_2 fanout5059 (.A(net5060),
    .X(net5059));
 sg13g2_buf_2 fanout5060 (.A(net5062),
    .X(net5060));
 sg13g2_buf_2 fanout5061 (.A(net5062),
    .X(net5061));
 sg13g2_buf_2 fanout5062 (.A(net5068),
    .X(net5062));
 sg13g2_buf_2 fanout5063 (.A(net5065),
    .X(net5063));
 sg13g2_buf_1 fanout5064 (.A(net5065),
    .X(net5064));
 sg13g2_buf_4 fanout5065 (.X(net5065),
    .A(net5068));
 sg13g2_buf_2 fanout5066 (.A(net5068),
    .X(net5066));
 sg13g2_buf_2 fanout5067 (.A(net5068),
    .X(net5067));
 sg13g2_buf_2 fanout5068 (.A(_03561_),
    .X(net5068));
 sg13g2_buf_2 fanout5069 (.A(_03533_),
    .X(net5069));
 sg13g2_buf_2 fanout5070 (.A(net5071),
    .X(net5070));
 sg13g2_buf_2 fanout5071 (.A(_03533_),
    .X(net5071));
 sg13g2_buf_2 fanout5072 (.A(net5073),
    .X(net5072));
 sg13g2_buf_2 fanout5073 (.A(_03507_),
    .X(net5073));
 sg13g2_buf_4 fanout5074 (.X(net5074),
    .A(net5075));
 sg13g2_buf_4 fanout5075 (.X(net5075),
    .A(net5076));
 sg13g2_buf_4 fanout5076 (.X(net5076),
    .A(net5081));
 sg13g2_buf_2 fanout5077 (.A(net5080),
    .X(net5077));
 sg13g2_buf_2 fanout5078 (.A(net5080),
    .X(net5078));
 sg13g2_buf_4 fanout5079 (.X(net5079),
    .A(net5080));
 sg13g2_buf_2 fanout5080 (.A(net5081),
    .X(net5080));
 sg13g2_buf_2 fanout5081 (.A(_03069_),
    .X(net5081));
 sg13g2_buf_2 fanout5082 (.A(net5092),
    .X(net5082));
 sg13g2_buf_2 fanout5083 (.A(net5084),
    .X(net5083));
 sg13g2_buf_2 fanout5084 (.A(net5092),
    .X(net5084));
 sg13g2_buf_2 fanout5085 (.A(net5086),
    .X(net5085));
 sg13g2_buf_2 fanout5086 (.A(net5091),
    .X(net5086));
 sg13g2_buf_2 fanout5087 (.A(net5088),
    .X(net5087));
 sg13g2_buf_2 fanout5088 (.A(net5091),
    .X(net5088));
 sg13g2_buf_2 fanout5089 (.A(net5091),
    .X(net5089));
 sg13g2_buf_2 fanout5090 (.A(net5091),
    .X(net5090));
 sg13g2_buf_2 fanout5091 (.A(net5092),
    .X(net5091));
 sg13g2_buf_2 fanout5092 (.A(_03069_),
    .X(net5092));
 sg13g2_buf_4 fanout5093 (.X(net5093),
    .A(_03067_));
 sg13g2_buf_4 fanout5094 (.X(net5094),
    .A(net5096));
 sg13g2_buf_1 fanout5095 (.A(net5096),
    .X(net5095));
 sg13g2_buf_4 fanout5096 (.X(net5096),
    .A(_03066_));
 sg13g2_buf_4 fanout5097 (.X(net5097),
    .A(net5098));
 sg13g2_buf_4 fanout5098 (.X(net5098),
    .A(_03065_));
 sg13g2_buf_4 fanout5099 (.X(net5099),
    .A(_03064_));
 sg13g2_buf_2 fanout5100 (.A(_03064_),
    .X(net5100));
 sg13g2_buf_4 fanout5101 (.X(net5101),
    .A(_03064_));
 sg13g2_buf_4 fanout5102 (.X(net5102),
    .A(net5103));
 sg13g2_buf_4 fanout5103 (.X(net5103),
    .A(net5104));
 sg13g2_buf_4 fanout5104 (.X(net5104),
    .A(_02781_));
 sg13g2_buf_4 fanout5105 (.X(net5105),
    .A(net5106));
 sg13g2_buf_4 fanout5106 (.X(net5106),
    .A(_02766_));
 sg13g2_buf_4 fanout5107 (.X(net5107),
    .A(net5109));
 sg13g2_buf_2 fanout5108 (.A(net5109),
    .X(net5108));
 sg13g2_buf_4 fanout5109 (.X(net5109),
    .A(_02765_));
 sg13g2_buf_2 fanout5110 (.A(net5119),
    .X(net5110));
 sg13g2_buf_2 fanout5111 (.A(net5119),
    .X(net5111));
 sg13g2_buf_2 fanout5112 (.A(net5113),
    .X(net5112));
 sg13g2_buf_2 fanout5113 (.A(net5119),
    .X(net5113));
 sg13g2_buf_2 fanout5114 (.A(net5115),
    .X(net5114));
 sg13g2_buf_2 fanout5115 (.A(net5118),
    .X(net5115));
 sg13g2_buf_2 fanout5116 (.A(net5118),
    .X(net5116));
 sg13g2_buf_2 fanout5117 (.A(net5118),
    .X(net5117));
 sg13g2_buf_2 fanout5118 (.A(net5119),
    .X(net5118));
 sg13g2_buf_2 fanout5119 (.A(_02763_),
    .X(net5119));
 sg13g2_buf_2 fanout5120 (.A(net5124),
    .X(net5120));
 sg13g2_buf_4 fanout5121 (.X(net5121),
    .A(net5124));
 sg13g2_buf_2 fanout5122 (.A(net5124),
    .X(net5122));
 sg13g2_buf_2 fanout5123 (.A(net5124),
    .X(net5123));
 sg13g2_buf_4 fanout5124 (.X(net5124),
    .A(_02747_));
 sg13g2_buf_4 fanout5125 (.X(net5125),
    .A(net5127));
 sg13g2_buf_1 fanout5126 (.A(net5127),
    .X(net5126));
 sg13g2_buf_4 fanout5127 (.X(net5127),
    .A(_02741_));
 sg13g2_buf_4 fanout5128 (.X(net5128),
    .A(net5129));
 sg13g2_buf_4 fanout5129 (.X(net5129),
    .A(_02741_));
 sg13g2_buf_2 fanout5130 (.A(net5132),
    .X(net5130));
 sg13g2_buf_1 fanout5131 (.A(net5132),
    .X(net5131));
 sg13g2_buf_2 fanout5132 (.A(_02735_),
    .X(net5132));
 sg13g2_buf_2 fanout5133 (.A(net5134),
    .X(net5133));
 sg13g2_buf_4 fanout5134 (.X(net5134),
    .A(_02735_));
 sg13g2_buf_4 fanout5135 (.X(net5135),
    .A(_02729_));
 sg13g2_buf_2 fanout5136 (.A(_02729_),
    .X(net5136));
 sg13g2_buf_2 fanout5137 (.A(net5139),
    .X(net5137));
 sg13g2_buf_2 fanout5138 (.A(net5139),
    .X(net5138));
 sg13g2_buf_4 fanout5139 (.X(net5139),
    .A(_02729_));
 sg13g2_buf_2 fanout5140 (.A(_02716_),
    .X(net5140));
 sg13g2_buf_2 fanout5141 (.A(_02636_),
    .X(net5141));
 sg13g2_buf_2 fanout5142 (.A(_02636_),
    .X(net5142));
 sg13g2_buf_4 fanout5143 (.X(net5143),
    .A(_05131_));
 sg13g2_buf_2 fanout5144 (.A(_05131_),
    .X(net5144));
 sg13g2_buf_2 fanout5145 (.A(net5147),
    .X(net5145));
 sg13g2_buf_2 fanout5146 (.A(net5147),
    .X(net5146));
 sg13g2_buf_4 fanout5147 (.X(net5147),
    .A(_04892_));
 sg13g2_buf_4 fanout5148 (.X(net5148),
    .A(net5152));
 sg13g2_buf_2 fanout5149 (.A(net5152),
    .X(net5149));
 sg13g2_buf_4 fanout5150 (.X(net5150),
    .A(net5151));
 sg13g2_buf_4 fanout5151 (.X(net5151),
    .A(net5152));
 sg13g2_buf_2 fanout5152 (.A(_03554_),
    .X(net5152));
 sg13g2_buf_4 fanout5153 (.X(net5153),
    .A(net5157));
 sg13g2_buf_4 fanout5154 (.X(net5154),
    .A(net5157));
 sg13g2_buf_4 fanout5155 (.X(net5155),
    .A(net5156));
 sg13g2_buf_4 fanout5156 (.X(net5156),
    .A(net5157));
 sg13g2_buf_4 fanout5157 (.X(net5157),
    .A(_02761_));
 sg13g2_buf_2 fanout5158 (.A(_02723_),
    .X(net5158));
 sg13g2_buf_4 fanout5159 (.X(net5159),
    .A(_02631_));
 sg13g2_buf_4 fanout5160 (.X(net5160),
    .A(_02496_));
 sg13g2_buf_2 fanout5161 (.A(net5162),
    .X(net5161));
 sg13g2_buf_2 fanout5162 (.A(_02490_),
    .X(net5162));
 sg13g2_buf_2 fanout5163 (.A(net5166),
    .X(net5163));
 sg13g2_buf_2 fanout5164 (.A(net5166),
    .X(net5164));
 sg13g2_buf_2 fanout5165 (.A(net5166),
    .X(net5165));
 sg13g2_buf_2 fanout5166 (.A(_02490_),
    .X(net5166));
 sg13g2_buf_4 fanout5167 (.X(net5167),
    .A(_02489_));
 sg13g2_buf_2 fanout5168 (.A(_02489_),
    .X(net5168));
 sg13g2_buf_4 fanout5169 (.X(net5169),
    .A(_02489_));
 sg13g2_buf_2 fanout5170 (.A(net5171),
    .X(net5170));
 sg13g2_buf_1 fanout5171 (.A(net5175),
    .X(net5171));
 sg13g2_buf_2 fanout5172 (.A(net5175),
    .X(net5172));
 sg13g2_buf_2 fanout5173 (.A(net5174),
    .X(net5173));
 sg13g2_buf_4 fanout5174 (.X(net5174),
    .A(net5175));
 sg13g2_buf_2 fanout5175 (.A(_02487_),
    .X(net5175));
 sg13g2_buf_4 fanout5176 (.X(net5176),
    .A(_02452_));
 sg13g2_buf_4 fanout5177 (.X(net5177),
    .A(_02450_));
 sg13g2_buf_4 fanout5178 (.X(net5178),
    .A(net5179));
 sg13g2_buf_4 fanout5179 (.X(net5179),
    .A(_02448_));
 sg13g2_buf_2 fanout5180 (.A(net5181),
    .X(net5180));
 sg13g2_buf_2 fanout5181 (.A(net5183),
    .X(net5181));
 sg13g2_buf_4 fanout5182 (.X(net5182),
    .A(net5183));
 sg13g2_buf_2 fanout5183 (.A(_02448_),
    .X(net5183));
 sg13g2_buf_4 fanout5184 (.X(net5184),
    .A(net5185));
 sg13g2_buf_4 fanout5185 (.X(net5185),
    .A(net5190));
 sg13g2_buf_4 fanout5186 (.X(net5186),
    .A(net5190));
 sg13g2_buf_2 fanout5187 (.A(net5188),
    .X(net5187));
 sg13g2_buf_2 fanout5188 (.A(net5189),
    .X(net5188));
 sg13g2_buf_2 fanout5189 (.A(net5190),
    .X(net5189));
 sg13g2_buf_2 fanout5190 (.A(_02447_),
    .X(net5190));
 sg13g2_buf_4 fanout5191 (.X(net5191),
    .A(_02445_));
 sg13g2_buf_4 fanout5192 (.X(net5192),
    .A(_02440_));
 sg13g2_buf_2 fanout5193 (.A(_02437_),
    .X(net5193));
 sg13g2_buf_4 fanout5194 (.X(net5194),
    .A(_02434_));
 sg13g2_buf_4 fanout5195 (.X(net5195),
    .A(_02432_));
 sg13g2_buf_4 fanout5196 (.X(net5196),
    .A(_02430_));
 sg13g2_buf_4 fanout5197 (.X(net5197),
    .A(_02427_));
 sg13g2_buf_2 fanout5198 (.A(net5200),
    .X(net5198));
 sg13g2_buf_4 fanout5199 (.X(net5199),
    .A(net5200));
 sg13g2_buf_2 fanout5200 (.A(net5207),
    .X(net5200));
 sg13g2_buf_2 fanout5201 (.A(net5202),
    .X(net5201));
 sg13g2_buf_1 fanout5202 (.A(net5203),
    .X(net5202));
 sg13g2_buf_2 fanout5203 (.A(net5204),
    .X(net5203));
 sg13g2_buf_2 fanout5204 (.A(net5207),
    .X(net5204));
 sg13g2_buf_4 fanout5205 (.X(net5205),
    .A(net5207));
 sg13g2_buf_2 fanout5206 (.A(net5207),
    .X(net5206));
 sg13g2_buf_2 fanout5207 (.A(_02424_),
    .X(net5207));
 sg13g2_buf_2 fanout5208 (.A(net5217),
    .X(net5208));
 sg13g2_buf_2 fanout5209 (.A(net5217),
    .X(net5209));
 sg13g2_buf_2 fanout5210 (.A(net5211),
    .X(net5210));
 sg13g2_buf_2 fanout5211 (.A(net5217),
    .X(net5211));
 sg13g2_buf_2 fanout5212 (.A(net5213),
    .X(net5212));
 sg13g2_buf_2 fanout5213 (.A(net5214),
    .X(net5213));
 sg13g2_buf_2 fanout5214 (.A(net5217),
    .X(net5214));
 sg13g2_buf_2 fanout5215 (.A(net5217),
    .X(net5215));
 sg13g2_buf_2 fanout5216 (.A(net5217),
    .X(net5216));
 sg13g2_buf_4 fanout5217 (.X(net5217),
    .A(_02423_));
 sg13g2_buf_4 fanout5218 (.X(net5218),
    .A(net5220));
 sg13g2_buf_2 fanout5219 (.A(net5220),
    .X(net5219));
 sg13g2_buf_2 fanout5220 (.A(_02422_),
    .X(net5220));
 sg13g2_buf_4 fanout5221 (.X(net5221),
    .A(_02402_));
 sg13g2_buf_4 fanout5222 (.X(net5222),
    .A(_02400_));
 sg13g2_buf_4 fanout5223 (.X(net5223),
    .A(_02399_));
 sg13g2_buf_4 fanout5224 (.X(net5224),
    .A(_02398_));
 sg13g2_buf_1 fanout5225 (.A(_02398_),
    .X(net5225));
 sg13g2_buf_4 fanout5226 (.X(net5226),
    .A(_02386_));
 sg13g2_buf_4 fanout5227 (.X(net5227),
    .A(_02385_));
 sg13g2_buf_4 fanout5228 (.X(net5228),
    .A(_02384_));
 sg13g2_buf_8 fanout5229 (.A(_02383_),
    .X(net5229));
 sg13g2_buf_4 fanout5230 (.X(net5230),
    .A(_02381_));
 sg13g2_buf_8 fanout5231 (.A(_02371_),
    .X(net5231));
 sg13g2_buf_4 fanout5232 (.X(net5232),
    .A(_02369_));
 sg13g2_buf_2 fanout5233 (.A(net5236),
    .X(net5233));
 sg13g2_buf_4 fanout5234 (.X(net5234),
    .A(net5236));
 sg13g2_buf_2 fanout5235 (.A(net5236),
    .X(net5235));
 sg13g2_buf_2 fanout5236 (.A(_02366_),
    .X(net5236));
 sg13g2_buf_2 fanout5237 (.A(net5238),
    .X(net5237));
 sg13g2_buf_1 fanout5238 (.A(_02366_),
    .X(net5238));
 sg13g2_buf_2 fanout5239 (.A(net5241),
    .X(net5239));
 sg13g2_buf_1 fanout5240 (.A(net5241),
    .X(net5240));
 sg13g2_buf_2 fanout5241 (.A(_02366_),
    .X(net5241));
 sg13g2_buf_2 fanout5242 (.A(\m_sys.m_core.m_fsm.r_cstate[0] ),
    .X(net5242));
 sg13g2_buf_2 fanout5243 (.A(net5244),
    .X(net5243));
 sg13g2_buf_2 fanout5244 (.A(net5254),
    .X(net5244));
 sg13g2_buf_2 fanout5245 (.A(net5246),
    .X(net5245));
 sg13g2_buf_2 fanout5246 (.A(net5254),
    .X(net5246));
 sg13g2_buf_2 fanout5247 (.A(net5249),
    .X(net5247));
 sg13g2_buf_2 fanout5248 (.A(net5249),
    .X(net5248));
 sg13g2_buf_2 fanout5249 (.A(net5254),
    .X(net5249));
 sg13g2_buf_2 fanout5250 (.A(net5252),
    .X(net5250));
 sg13g2_buf_1 fanout5251 (.A(net5252),
    .X(net5251));
 sg13g2_buf_2 fanout5252 (.A(net5254),
    .X(net5252));
 sg13g2_buf_2 fanout5253 (.A(net5254),
    .X(net5253));
 sg13g2_buf_2 fanout5254 (.A(\m_sys.m_core.m_alu.io_i_signed ),
    .X(net5254));
 sg13g2_buf_4 fanout5255 (.X(net5255),
    .A(net5256));
 sg13g2_buf_4 fanout5256 (.X(net5256),
    .A(net5259));
 sg13g2_buf_2 fanout5257 (.A(net5259),
    .X(net5257));
 sg13g2_buf_2 fanout5258 (.A(net5259),
    .X(net5258));
 sg13g2_buf_2 fanout5259 (.A(\m_sys.m_core.m_alu.io_i_uop[2] ),
    .X(net5259));
 sg13g2_buf_4 fanout5260 (.X(net5260),
    .A(net2811));
 sg13g2_buf_4 fanout5261 (.X(net5261),
    .A(net2663));
 sg13g2_buf_4 fanout5262 (.X(net5262),
    .A(net2759));
 sg13g2_buf_4 fanout5263 (.X(net5263),
    .A(net3003));
 sg13g2_buf_4 fanout5264 (.X(net5264),
    .A(net2846));
 sg13g2_buf_4 fanout5265 (.X(net5265),
    .A(net2752));
 sg13g2_buf_2 fanout5266 (.A(net5267),
    .X(net5266));
 sg13g2_buf_4 fanout5267 (.X(net5267),
    .A(\m_sys._m_bootloader_io_b_mem_addr[0] ));
 sg13g2_buf_2 fanout5268 (.A(net5270),
    .X(net5268));
 sg13g2_buf_1 fanout5269 (.A(net5270),
    .X(net5269));
 sg13g2_buf_4 fanout5270 (.X(net5270),
    .A(net5271));
 sg13g2_buf_4 fanout5271 (.X(net5271),
    .A(net5273));
 sg13g2_buf_4 fanout5272 (.X(net5272),
    .A(net5273));
 sg13g2_buf_2 fanout5273 (.A(\m_sys._m_bootloader_io_o_bl ),
    .X(net5273));
 sg13g2_buf_2 fanout5274 (.A(net5277),
    .X(net5274));
 sg13g2_buf_2 fanout5275 (.A(net5277),
    .X(net5275));
 sg13g2_buf_1 fanout5276 (.A(net5277),
    .X(net5276));
 sg13g2_buf_2 fanout5277 (.A(net5279),
    .X(net5277));
 sg13g2_buf_2 fanout5278 (.A(net5279),
    .X(net5278));
 sg13g2_buf_2 fanout5279 (.A(\m_sys.r_valid ),
    .X(net5279));
 sg13g2_buf_2 fanout5280 (.A(net5281),
    .X(net5280));
 sg13g2_buf_2 fanout5281 (.A(\m_sys.r_valid ),
    .X(net5281));
 sg13g2_buf_2 fanout5282 (.A(\m_sys.m_bootloader.r_cstate[3] ),
    .X(net5282));
 sg13g2_buf_4 fanout5283 (.X(net5283),
    .A(net3425));
 sg13g2_buf_2 fanout5284 (.A(net5285),
    .X(net5284));
 sg13g2_buf_2 fanout5285 (.A(net5286),
    .X(net5285));
 sg13g2_buf_2 fanout5286 (.A(\m_sys.m_bootloader.r_cstate[0] ),
    .X(net5286));
 sg13g2_buf_2 fanout5287 (.A(net3396),
    .X(net5287));
 sg13g2_buf_4 fanout5288 (.X(net5288),
    .A(\m_sys.m_core.m_alu.io_i_uop[1] ));
 sg13g2_buf_2 fanout5289 (.A(net5292),
    .X(net5289));
 sg13g2_buf_1 fanout5290 (.A(net5292),
    .X(net5290));
 sg13g2_buf_2 fanout5291 (.A(net5292),
    .X(net5291));
 sg13g2_buf_2 fanout5292 (.A(\m_sys.m_core.m_alu.io_i_uop[1] ),
    .X(net5292));
 sg13g2_buf_2 fanout5293 (.A(net5294),
    .X(net5293));
 sg13g2_buf_1 fanout5294 (.A(net5302),
    .X(net5294));
 sg13g2_buf_2 fanout5295 (.A(net5301),
    .X(net5295));
 sg13g2_buf_1 fanout5296 (.A(net5301),
    .X(net5296));
 sg13g2_buf_2 fanout5297 (.A(net5301),
    .X(net5297));
 sg13g2_buf_2 fanout5298 (.A(net5299),
    .X(net5298));
 sg13g2_buf_1 fanout5299 (.A(net5300),
    .X(net5299));
 sg13g2_buf_1 fanout5300 (.A(net5301),
    .X(net5300));
 sg13g2_buf_2 fanout5301 (.A(net5302),
    .X(net5301));
 sg13g2_buf_2 fanout5302 (.A(net3428),
    .X(net5302));
 sg13g2_buf_2 fanout5303 (.A(net5306),
    .X(net5303));
 sg13g2_buf_2 fanout5304 (.A(net5306),
    .X(net5304));
 sg13g2_buf_2 fanout5305 (.A(net5306),
    .X(net5305));
 sg13g2_buf_2 fanout5306 (.A(net5308),
    .X(net5306));
 sg13g2_buf_4 fanout5307 (.X(net5307),
    .A(net5308));
 sg13g2_buf_2 fanout5308 (.A(\m_sys.m_core.m_alu.io_i_uop[0] ),
    .X(net5308));
 sg13g2_buf_2 fanout5309 (.A(\m_sys.m_core.m_fsm.r_cstate[1] ),
    .X(net5309));
 sg13g2_buf_4 fanout5310 (.X(net5310),
    .A(net5311));
 sg13g2_buf_4 fanout5311 (.X(net5311),
    .A(\m_sys._m_core_io_b_mem_wdata[0] ));
 sg13g2_buf_4 fanout5312 (.X(net5312),
    .A(\m_sys.m_core.m_bru.io_i_s1[1] ));
 sg13g2_buf_4 fanout5313 (.X(net5313),
    .A(\m_sys.m_core.m_bru.io_i_s1[3] ));
 sg13g2_buf_1 fanout5314 (.A(\m_sys.m_core.m_bru.io_i_s1[3] ),
    .X(net5314));
 sg13g2_buf_4 fanout5315 (.X(net5315),
    .A(net5316));
 sg13g2_buf_4 fanout5316 (.X(net5316),
    .A(\m_sys.m_core.m_bru.io_i_s1[4] ));
 sg13g2_buf_4 fanout5317 (.X(net5317),
    .A(net5318));
 sg13g2_buf_2 fanout5318 (.A(net5319),
    .X(net5318));
 sg13g2_buf_4 fanout5319 (.X(net5319),
    .A(\m_sys.m_core.m_bru.io_i_s1[5] ));
 sg13g2_buf_4 fanout5320 (.X(net5320),
    .A(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[1] ));
 sg13g2_buf_2 fanout5321 (.A(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[1] ),
    .X(net5321));
 sg13g2_buf_2 fanout5322 (.A(\m_sys.m_core.m_bru.io_i_s1[12] ),
    .X(net5322));
 sg13g2_buf_2 fanout5323 (.A(\m_sys.m_core.m_bru.io_i_s1[13] ),
    .X(net5323));
 sg13g2_buf_8 fanout5324 (.A(\m_sys.m_core._m_decoder_io_o_rs1[0] ),
    .X(net5324));
 sg13g2_buf_4 fanout5325 (.X(net5325),
    .A(net5326));
 sg13g2_buf_4 fanout5326 (.X(net5326),
    .A(\m_sys.m_core._m_decoder_io_o_rs1[1] ));
 sg13g2_buf_4 fanout5327 (.X(net5327),
    .A(net5328));
 sg13g2_buf_4 fanout5328 (.X(net5328),
    .A(\m_sys.m_core._m_decoder_io_o_rs1[2] ));
 sg13g2_buf_2 fanout5329 (.A(net5331),
    .X(net5329));
 sg13g2_buf_4 fanout5330 (.X(net5330),
    .A(net5331));
 sg13g2_buf_2 fanout5331 (.A(\m_sys.m_core._m_decoder_io_o_rs1[2] ),
    .X(net5331));
 sg13g2_buf_4 fanout5332 (.X(net5332),
    .A(net5335));
 sg13g2_buf_2 fanout5333 (.A(net5335),
    .X(net5333));
 sg13g2_buf_4 fanout5334 (.X(net5334),
    .A(net5335));
 sg13g2_buf_2 fanout5335 (.A(\m_sys.m_core._m_decoder_io_o_rs2[0] ),
    .X(net5335));
 sg13g2_buf_4 fanout5336 (.X(net5336),
    .A(net5340));
 sg13g2_buf_4 fanout5337 (.X(net5337),
    .A(net5340));
 sg13g2_buf_4 fanout5338 (.X(net5338),
    .A(net5339));
 sg13g2_buf_4 fanout5339 (.X(net5339),
    .A(net5340));
 sg13g2_buf_4 fanout5340 (.X(net5340),
    .A(\m_sys.m_core._m_decoder_io_o_rs2[0] ));
 sg13g2_buf_4 fanout5341 (.X(net5341),
    .A(net5344));
 sg13g2_buf_2 fanout5342 (.A(net5344),
    .X(net5342));
 sg13g2_buf_4 fanout5343 (.X(net5343),
    .A(net5344));
 sg13g2_buf_2 fanout5344 (.A(net5350),
    .X(net5344));
 sg13g2_buf_4 fanout5345 (.X(net5345),
    .A(net5346));
 sg13g2_buf_2 fanout5346 (.A(net5350),
    .X(net5346));
 sg13g2_buf_2 fanout5347 (.A(net5349),
    .X(net5347));
 sg13g2_buf_2 fanout5348 (.A(net5349),
    .X(net5348));
 sg13g2_buf_2 fanout5349 (.A(net5350),
    .X(net5349));
 sg13g2_buf_2 fanout5350 (.A(\m_sys.m_core._m_decoder_io_o_rs2[1] ),
    .X(net5350));
 sg13g2_buf_4 fanout5351 (.X(net5351),
    .A(net5352));
 sg13g2_buf_4 fanout5352 (.X(net5352),
    .A(\m_sys.m_core._m_decoder_io_o_rs2[2] ));
 sg13g2_buf_4 fanout5353 (.X(net5353),
    .A(\m_sys.m_core.m_bru.io_i_s1[31] ));
 sg13g2_buf_2 fanout5354 (.A(net5355),
    .X(net5354));
 sg13g2_buf_2 fanout5355 (.A(net5359),
    .X(net5355));
 sg13g2_buf_1 fanout5356 (.A(net5359),
    .X(net5356));
 sg13g2_buf_2 fanout5357 (.A(net5359),
    .X(net5357));
 sg13g2_buf_2 fanout5358 (.A(net5359),
    .X(net5358));
 sg13g2_buf_1 fanout5359 (.A(\m_sys._GEN_11[4] ),
    .X(net5359));
 sg13g2_buf_4 fanout5360 (.X(net5360),
    .A(net5361));
 sg13g2_buf_2 fanout5361 (.A(\m_sys._GEN_11[3] ),
    .X(net5361));
 sg13g2_buf_2 fanout5362 (.A(net5366),
    .X(net5362));
 sg13g2_buf_2 fanout5363 (.A(net5365),
    .X(net5363));
 sg13g2_buf_2 fanout5364 (.A(net5366),
    .X(net5364));
 sg13g2_buf_1 fanout5365 (.A(net5366),
    .X(net5365));
 sg13g2_buf_2 fanout5366 (.A(\m_sys._GEN_11[3] ),
    .X(net5366));
 sg13g2_buf_2 fanout5367 (.A(net5368),
    .X(net5367));
 sg13g2_buf_4 fanout5368 (.X(net5368),
    .A(net5378));
 sg13g2_buf_4 fanout5369 (.X(net5369),
    .A(net5370));
 sg13g2_buf_1 fanout5370 (.A(net5378),
    .X(net5370));
 sg13g2_buf_2 fanout5371 (.A(net5375),
    .X(net5371));
 sg13g2_buf_1 fanout5372 (.A(net5375),
    .X(net5372));
 sg13g2_buf_2 fanout5373 (.A(net5375),
    .X(net5373));
 sg13g2_buf_1 fanout5374 (.A(net5375),
    .X(net5374));
 sg13g2_buf_2 fanout5375 (.A(net5378),
    .X(net5375));
 sg13g2_buf_4 fanout5376 (.X(net5376),
    .A(net5378));
 sg13g2_buf_2 fanout5377 (.A(net5378),
    .X(net5377));
 sg13g2_buf_4 fanout5378 (.X(net5378),
    .A(_02396_));
 sg13g2_buf_4 fanout5379 (.X(net5379),
    .A(net5385));
 sg13g2_buf_1 fanout5380 (.A(net5385),
    .X(net5380));
 sg13g2_buf_2 fanout5381 (.A(net5383),
    .X(net5381));
 sg13g2_buf_1 fanout5382 (.A(net5383),
    .X(net5382));
 sg13g2_buf_2 fanout5383 (.A(net5385),
    .X(net5383));
 sg13g2_buf_4 fanout5384 (.X(net5384),
    .A(net5385));
 sg13g2_buf_4 fanout5385 (.X(net5385),
    .A(rst_n));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tiehi _18673__17 (.L_HI(net17));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_leaf_85_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_2 clkbuf_leaf_86_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_2 clkbuf_leaf_87_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_2 clkbuf_leaf_88_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_2 clkbuf_leaf_89_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_2 clkbuf_leaf_90_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_2 clkbuf_leaf_91_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_2 clkbuf_leaf_92_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_2 clkbuf_leaf_93_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_2 clkbuf_leaf_94_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_2 clkbuf_leaf_95_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_2 clkbuf_leaf_96_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_2 clkbuf_leaf_97_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_2 clkbuf_leaf_98_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_2 clkbuf_leaf_99_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_2 clkbuf_leaf_100_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_2 clkbuf_leaf_101_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_2 clkbuf_leaf_102_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_2 clkbuf_leaf_103_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_2 clkbuf_leaf_104_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_2 clkbuf_leaf_105_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_2 clkbuf_leaf_106_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_2 clkbuf_leaf_107_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_2 clkbuf_leaf_108_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_2 clkbuf_leaf_109_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_2 clkbuf_leaf_110_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_2 clkbuf_leaf_111_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_2 clkbuf_leaf_112_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_2 clkbuf_leaf_113_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_2 clkbuf_leaf_114_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_2 clkbuf_leaf_115_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_2 clkbuf_leaf_116_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_2 clkbuf_leaf_117_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_2 clkbuf_leaf_118_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_2 clkbuf_leaf_119_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_2 clkbuf_leaf_120_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_2 clkbuf_leaf_121_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_2 clkbuf_leaf_122_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_2 clkbuf_leaf_123_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_2 clkbuf_leaf_124_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_2 clkbuf_leaf_125_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_2 clkbuf_leaf_126_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_2 clkbuf_leaf_127_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_2 clkbuf_leaf_128_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_2 clkbuf_leaf_129_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_2 clkbuf_leaf_130_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_2 clkbuf_leaf_131_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_2 clkbuf_leaf_132_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_2 clkbuf_leaf_133_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_2 clkbuf_leaf_134_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_2 clkbuf_leaf_135_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_2 clkbuf_leaf_136_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_2 clkbuf_leaf_137_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_2 clkbuf_leaf_138_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_2 clkbuf_leaf_139_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_2 clkbuf_leaf_140_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_2 clkbuf_leaf_141_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_2 clkbuf_leaf_142_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_2 clkbuf_leaf_143_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_2 clkbuf_leaf_144_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_2 clkbuf_leaf_145_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_2 clkbuf_leaf_146_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_2 clkbuf_leaf_147_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_2 clkbuf_leaf_148_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_2 clkbuf_leaf_149_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_2 clkbuf_leaf_150_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_2 clkbuf_leaf_151_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_2 clkbuf_leaf_152_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_2 clkbuf_leaf_153_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_2 clkbuf_leaf_154_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_2 clkbuf_leaf_155_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_2 clkbuf_leaf_156_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_2 clkbuf_leaf_157_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_2 clkbuf_leaf_158_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_2 clkbuf_leaf_159_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_2 clkbuf_leaf_160_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_2 clkbuf_leaf_161_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_2 clkbuf_leaf_162_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_2 clkbuf_leaf_163_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_2 clkbuf_leaf_164_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_2 clkbuf_leaf_165_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_2 clkbuf_leaf_166_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_2 clkbuf_leaf_167_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_2 clkbuf_leaf_168_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_2 clkbuf_leaf_169_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_2 clkbuf_leaf_170_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_2 clkbuf_leaf_171_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_2 clkbuf_leaf_172_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_2 clkbuf_leaf_173_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_2 clkbuf_leaf_174_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_2 clkbuf_leaf_175_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_2 clkbuf_leaf_176_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_2 clkbuf_leaf_177_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_2 clkbuf_leaf_178_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_2 clkbuf_leaf_179_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_2 clkbuf_leaf_180_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_2 clkbuf_leaf_181_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_2 clkbuf_leaf_182_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_2 clkbuf_leaf_183_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_2 clkbuf_leaf_184_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_2 clkbuf_leaf_185_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_2 clkbuf_leaf_186_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_2 clkbuf_leaf_187_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_2 clkbuf_leaf_188_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_2 clkbuf_leaf_189_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_2 clkbuf_leaf_190_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_2 clkbuf_leaf_191_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_2 clkbuf_leaf_192_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_2 clkbuf_leaf_193_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_2 clkbuf_leaf_194_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_2 clkbuf_leaf_195_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_2 clkbuf_leaf_196_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_2 clkbuf_leaf_197_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_2 clkbuf_leaf_198_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_2 clkbuf_leaf_199_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_2 clkbuf_leaf_200_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_2 clkbuf_leaf_201_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_2 clkbuf_leaf_202_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_2 clkbuf_leaf_203_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_2 clkbuf_leaf_204_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_2 clkbuf_leaf_205_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_2 clkbuf_leaf_206_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_2 clkbuf_leaf_207_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_2 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_2 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_2 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_2 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_2 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_2 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_2 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkload7 (.A(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkload8 (.A(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkload9 (.A(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkload10 (.A(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkload11 (.A(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkload12 (.A(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkload13 (.A(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkload14 (.A(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkload15 (.A(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_207_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_59_clk));
 sg13g2_inv_4 clkload18 (.A(clknet_leaf_35_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_34_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_70_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_144_clk));
 sg13g2_inv_4 clkload22 (.A(clknet_leaf_83_clk));
 sg13g2_inv_8 clkload23 (.A(clknet_leaf_84_clk));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_87_clk));
 sg13g2_inv_1 clkload25 (.A(clknet_leaf_89_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_00046_),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold2 (.A(_00077_),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold3 (.A(_00174_),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold4 (.A(\m_sys.m_uart.r_rx_data[6] ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold5 (.A(_07418_),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold6 (.A(\m_sys.m_uart.r_rx_data[5] ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold7 (.A(_07417_),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold8 (.A(\m_sys.m_ram.m_ram.r_mem[8][6] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold9 (.A(\m_sys.m_ram.m_ram.r_mem[17][7] ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold10 (.A(\m_sys.m_ram.m_ram.r_mem[21][1] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold11 (.A(\m_sys.m_ram.m_ram.r_mem[5][12] ),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold12 (.A(\m_sys.m_ram.m_ram.r_mem[4][5] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold13 (.A(\m_sys.m_ram.m_ram.r_mem[29][4] ),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold14 (.A(\m_sys.m_ram.m_ram.r_mem[20][5] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold15 (.A(\m_sys.m_ram.m_ram.r_mem[8][5] ),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold16 (.A(\m_sys.m_ram.m_ram.r_mem[5][0] ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold17 (.A(\m_sys.m_ram.m_ram.r_mem[1][11] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold18 (.A(\m_sys.m_ram.m_ram.r_mem[20][3] ),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold19 (.A(\m_sys.m_ram.m_ram.r_mem[9][9] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold20 (.A(\m_sys.m_ram.m_ram.r_mem[25][2] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold21 (.A(\m_sys.m_ram.m_ram.r_mem[1][13] ),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold22 (.A(\m_sys.m_ram.m_ram.r_mem[1][15] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold23 (.A(\m_sys.m_ram.m_ram.r_mem[18][6] ),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold24 (.A(\m_sys.m_ram.m_ram.r_mem[1][10] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold25 (.A(\m_sys.m_ram.m_ram.r_mem[21][3] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold26 (.A(\m_sys.m_ram.m_ram.r_mem[18][7] ),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold27 (.A(\m_sys.m_ram.m_ram.r_mem[29][1] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold28 (.A(\m_sys.m_ram.m_ram.r_mem[18][10] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold29 (.A(\m_sys.m_ram.m_ram.r_mem[30][14] ),
    .X(net1682));
 sg13g2_dlygate4sd3_1 hold30 (.A(\m_sys.m_ram.m_ram.r_mem[5][2] ),
    .X(net1683));
 sg13g2_dlygate4sd3_1 hold31 (.A(\m_sys.m_ram.m_ram.r_mem[29][0] ),
    .X(net1684));
 sg13g2_dlygate4sd3_1 hold32 (.A(\m_sys.m_ram.m_ram.r_mem[24][8] ),
    .X(net1685));
 sg13g2_dlygate4sd3_1 hold33 (.A(\m_sys.m_ram.m_ram.r_mem[28][2] ),
    .X(net1686));
 sg13g2_dlygate4sd3_1 hold34 (.A(\m_sys.m_ram.m_ram.r_mem[0][0] ),
    .X(net1687));
 sg13g2_dlygate4sd3_1 hold35 (.A(\m_sys.m_ram.m_ram.r_mem[2][13] ),
    .X(net1688));
 sg13g2_dlygate4sd3_1 hold36 (.A(\m_sys.m_ram.m_ram.r_mem[20][6] ),
    .X(net1689));
 sg13g2_dlygate4sd3_1 hold37 (.A(\m_sys.m_ram.m_ram.r_mem[21][14] ),
    .X(net1690));
 sg13g2_dlygate4sd3_1 hold38 (.A(\m_sys.m_ram.m_ram.r_mem[29][15] ),
    .X(net1691));
 sg13g2_dlygate4sd3_1 hold39 (.A(\m_sys.m_ram.m_ram.r_mem[1][1] ),
    .X(net1692));
 sg13g2_dlygate4sd3_1 hold40 (.A(\m_sys.m_ram.m_ram.r_mem[16][11] ),
    .X(net1693));
 sg13g2_dlygate4sd3_1 hold41 (.A(\m_sys.m_ram.m_ram.r_mem[6][2] ),
    .X(net1694));
 sg13g2_dlygate4sd3_1 hold42 (.A(\m_sys.m_ram.m_ram.r_mem[21][4] ),
    .X(net1695));
 sg13g2_dlygate4sd3_1 hold43 (.A(\m_sys.m_ram.m_ram.r_mem[0][14] ),
    .X(net1696));
 sg13g2_dlygate4sd3_1 hold44 (.A(\m_sys.m_ram.m_ram.r_mem[25][10] ),
    .X(net1697));
 sg13g2_dlygate4sd3_1 hold45 (.A(\m_sys.m_ram.m_ram.r_mem[12][14] ),
    .X(net1698));
 sg13g2_dlygate4sd3_1 hold46 (.A(\m_sys.m_ram.m_ram.r_mem[8][14] ),
    .X(net1699));
 sg13g2_dlygate4sd3_1 hold47 (.A(\m_sys.m_ram.m_ram.r_mem[1][6] ),
    .X(net1700));
 sg13g2_dlygate4sd3_1 hold48 (.A(\m_sys.m_ram.m_ram.r_mem[20][15] ),
    .X(net1701));
 sg13g2_dlygate4sd3_1 hold49 (.A(\m_sys.m_ram.m_ram.r_mem[21][8] ),
    .X(net1702));
 sg13g2_dlygate4sd3_1 hold50 (.A(\m_sys.m_ram.m_ram.r_mem[8][8] ),
    .X(net1703));
 sg13g2_dlygate4sd3_1 hold51 (.A(\m_sys.m_ram.m_ram.r_mem[12][15] ),
    .X(net1704));
 sg13g2_dlygate4sd3_1 hold52 (.A(\m_sys.m_ram.m_ram.r_mem[9][7] ),
    .X(net1705));
 sg13g2_dlygate4sd3_1 hold53 (.A(\m_sys.m_ram.m_ram.r_mem[21][6] ),
    .X(net1706));
 sg13g2_dlygate4sd3_1 hold54 (.A(\m_sys.m_ram.m_ram.r_mem[26][11] ),
    .X(net1707));
 sg13g2_dlygate4sd3_1 hold55 (.A(\m_sys.m_ram.m_ram.r_mem[1][9] ),
    .X(net1708));
 sg13g2_dlygate4sd3_1 hold56 (.A(\m_sys.m_ram.m_ram.r_mem[31][8] ),
    .X(net1709));
 sg13g2_dlygate4sd3_1 hold57 (.A(\m_sys.m_ram.m_ram.r_mem[25][3] ),
    .X(net1710));
 sg13g2_dlygate4sd3_1 hold58 (.A(\m_sys.m_ram.m_ram.r_mem[14][13] ),
    .X(net1711));
 sg13g2_dlygate4sd3_1 hold59 (.A(\m_sys.m_ram.m_ram.r_mem[2][9] ),
    .X(net1712));
 sg13g2_dlygate4sd3_1 hold60 (.A(\m_sys.m_ram.m_ram.r_mem[5][9] ),
    .X(net1713));
 sg13g2_dlygate4sd3_1 hold61 (.A(\m_sys.m_ram.m_ram.r_mem[17][6] ),
    .X(net1714));
 sg13g2_dlygate4sd3_1 hold62 (.A(\m_sys.m_ram.m_ram.r_mem[5][11] ),
    .X(net1715));
 sg13g2_dlygate4sd3_1 hold63 (.A(\m_sys.m_ram.m_ram.r_mem[29][8] ),
    .X(net1716));
 sg13g2_dlygate4sd3_1 hold64 (.A(\m_sys.m_ram.m_ram.r_mem[26][13] ),
    .X(net1717));
 sg13g2_dlygate4sd3_1 hold65 (.A(\m_sys.m_ram.m_ram.r_mem[28][4] ),
    .X(net1718));
 sg13g2_dlygate4sd3_1 hold66 (.A(\m_sys.m_ram.m_ram.r_mem[12][9] ),
    .X(net1719));
 sg13g2_dlygate4sd3_1 hold67 (.A(\m_sys.m_ram.m_ram.r_mem[20][14] ),
    .X(net1720));
 sg13g2_dlygate4sd3_1 hold68 (.A(\m_sys.m_ram.m_ram.r_mem[21][15] ),
    .X(net1721));
 sg13g2_dlygate4sd3_1 hold69 (.A(\m_sys.m_ram.m_ram.r_mem[9][3] ),
    .X(net1722));
 sg13g2_dlygate4sd3_1 hold70 (.A(\m_sys.m_ram.m_ram.r_mem[9][5] ),
    .X(net1723));
 sg13g2_dlygate4sd3_1 hold71 (.A(\m_sys.m_ram.m_ram.r_mem[0][6] ),
    .X(net1724));
 sg13g2_dlygate4sd3_1 hold72 (.A(\m_sys.m_ram.m_ram.r_mem[28][14] ),
    .X(net1725));
 sg13g2_dlygate4sd3_1 hold73 (.A(\m_sys.m_ram.m_ram.r_mem[14][11] ),
    .X(net1726));
 sg13g2_dlygate4sd3_1 hold74 (.A(\m_sys.m_ram.m_ram.r_mem[21][9] ),
    .X(net1727));
 sg13g2_dlygate4sd3_1 hold75 (.A(\m_sys.m_ram.m_ram.r_mem[25][13] ),
    .X(net1728));
 sg13g2_dlygate4sd3_1 hold76 (.A(\m_sys.m_ram.m_ram.r_mem[4][15] ),
    .X(net1729));
 sg13g2_dlygate4sd3_1 hold77 (.A(\m_sys.m_ram.m_ram.r_mem[8][12] ),
    .X(net1730));
 sg13g2_dlygate4sd3_1 hold78 (.A(\m_sys.m_ram.m_ram.r_mem[1][12] ),
    .X(net1731));
 sg13g2_dlygate4sd3_1 hold79 (.A(\m_sys.m_ram.m_ram.r_mem[6][0] ),
    .X(net1732));
 sg13g2_dlygate4sd3_1 hold80 (.A(\m_sys.m_ram.m_ram.r_mem[21][12] ),
    .X(net1733));
 sg13g2_dlygate4sd3_1 hold81 (.A(\m_sys.m_ram.m_ram.r_mem[25][15] ),
    .X(net1734));
 sg13g2_dlygate4sd3_1 hold82 (.A(\m_sys.m_ram.m_ram.r_mem[18][2] ),
    .X(net1735));
 sg13g2_dlygate4sd3_1 hold83 (.A(\m_sys.m_ram.m_ram.r_mem[16][5] ),
    .X(net1736));
 sg13g2_dlygate4sd3_1 hold84 (.A(\m_sys.m_ram.m_ram.r_mem[12][12] ),
    .X(net1737));
 sg13g2_dlygate4sd3_1 hold85 (.A(\m_sys.m_ram.m_ram.r_mem[26][2] ),
    .X(net1738));
 sg13g2_dlygate4sd3_1 hold86 (.A(\m_sys.m_ram.m_ram.r_mem[29][12] ),
    .X(net1739));
 sg13g2_dlygate4sd3_1 hold87 (.A(\m_sys.m_ram.m_ram.r_mem[16][14] ),
    .X(net1740));
 sg13g2_dlygate4sd3_1 hold88 (.A(\m_sys.m_ram.m_ram.r_mem[1][5] ),
    .X(net1741));
 sg13g2_dlygate4sd3_1 hold89 (.A(\m_sys.m_ram.m_ram.r_mem[30][10] ),
    .X(net1742));
 sg13g2_dlygate4sd3_1 hold90 (.A(\m_sys.m_ram.m_ram.r_mem[25][7] ),
    .X(net1743));
 sg13g2_dlygate4sd3_1 hold91 (.A(\m_sys.m_ram.m_ram.r_mem[9][1] ),
    .X(net1744));
 sg13g2_dlygate4sd3_1 hold92 (.A(\m_sys.m_ram.m_ram.r_mem[8][2] ),
    .X(net1745));
 sg13g2_dlygate4sd3_1 hold93 (.A(\m_sys.m_ram.m_ram.r_mem[17][11] ),
    .X(net1746));
 sg13g2_dlygate4sd3_1 hold94 (.A(\m_sys.m_ram.m_ram.r_mem[0][2] ),
    .X(net1747));
 sg13g2_dlygate4sd3_1 hold95 (.A(\m_sys.m_ram.m_ram.r_mem[8][0] ),
    .X(net1748));
 sg13g2_dlygate4sd3_1 hold96 (.A(\m_sys.m_ram.m_ram.r_mem[3][9] ),
    .X(net1749));
 sg13g2_dlygate4sd3_1 hold97 (.A(\m_sys.m_ram.m_ram.r_mem[16][1] ),
    .X(net1750));
 sg13g2_dlygate4sd3_1 hold98 (.A(\m_sys.m_ram.m_ram.r_mem[19][2] ),
    .X(net1751));
 sg13g2_dlygate4sd3_1 hold99 (.A(\m_sys.m_ram.m_ram.r_mem[24][15] ),
    .X(net1752));
 sg13g2_dlygate4sd3_1 hold100 (.A(\m_sys.m_ram.m_ram.r_mem[27][12] ),
    .X(net1753));
 sg13g2_dlygate4sd3_1 hold101 (.A(\m_sys.m_ram.m_ram.r_mem[24][11] ),
    .X(net1754));
 sg13g2_dlygate4sd3_1 hold102 (.A(\m_sys.m_ram.m_ram.r_mem[17][4] ),
    .X(net1755));
 sg13g2_dlygate4sd3_1 hold103 (.A(\m_sys.m_ram.m_ram.r_mem[16][13] ),
    .X(net1756));
 sg13g2_dlygate4sd3_1 hold104 (.A(\m_sys.m_ram.m_ram.r_mem[25][11] ),
    .X(net1757));
 sg13g2_dlygate4sd3_1 hold105 (.A(\m_sys.m_ram.m_ram.r_mem[28][3] ),
    .X(net1758));
 sg13g2_dlygate4sd3_1 hold106 (.A(\m_sys.m_ram.m_ram.r_mem[2][15] ),
    .X(net1759));
 sg13g2_dlygate4sd3_1 hold107 (.A(\m_sys.m_ram.m_ram.r_mem[30][8] ),
    .X(net1760));
 sg13g2_dlygate4sd3_1 hold108 (.A(\m_sys.m_ram.m_ram.r_mem[9][0] ),
    .X(net1761));
 sg13g2_dlygate4sd3_1 hold109 (.A(\m_sys.m_ram.m_ram.r_mem[13][4] ),
    .X(net1762));
 sg13g2_dlygate4sd3_1 hold110 (.A(\m_sys.m_ram.m_ram.r_mem[6][15] ),
    .X(net1763));
 sg13g2_dlygate4sd3_1 hold111 (.A(\m_sys.m_ram.m_ram.r_mem[14][14] ),
    .X(net1764));
 sg13g2_dlygate4sd3_1 hold112 (.A(\m_sys.m_ram.m_ram.r_mem[23][6] ),
    .X(net1765));
 sg13g2_dlygate4sd3_1 hold113 (.A(\m_sys.m_ram.m_ram.r_mem[3][15] ),
    .X(net1766));
 sg13g2_dlygate4sd3_1 hold114 (.A(\m_sys.m_ram.m_ram.r_mem[4][8] ),
    .X(net1767));
 sg13g2_dlygate4sd3_1 hold115 (.A(\m_sys.m_ram.m_ram.r_mem[21][2] ),
    .X(net1768));
 sg13g2_dlygate4sd3_1 hold116 (.A(\m_sys.m_ram.m_ram.r_mem[6][1] ),
    .X(net1769));
 sg13g2_dlygate4sd3_1 hold117 (.A(\m_sys.m_ram.m_ram.r_mem[28][6] ),
    .X(net1770));
 sg13g2_dlygate4sd3_1 hold118 (.A(\m_sys.m_ram.m_ram.r_mem[6][8] ),
    .X(net1771));
 sg13g2_dlygate4sd3_1 hold119 (.A(\m_sys.m_ram.m_ram.r_mem[17][9] ),
    .X(net1772));
 sg13g2_dlygate4sd3_1 hold120 (.A(\m_sys.m_ram.m_ram.r_mem[21][11] ),
    .X(net1773));
 sg13g2_dlygate4sd3_1 hold121 (.A(\m_sys.m_ram.m_ram.r_mem[19][9] ),
    .X(net1774));
 sg13g2_dlygate4sd3_1 hold122 (.A(\m_sys.m_ram.m_ram.r_mem[27][15] ),
    .X(net1775));
 sg13g2_dlygate4sd3_1 hold123 (.A(\m_sys.m_ram.m_ram.r_mem[9][8] ),
    .X(net1776));
 sg13g2_dlygate4sd3_1 hold124 (.A(\m_sys.m_ram.m_ram.r_mem[15][7] ),
    .X(net1777));
 sg13g2_dlygate4sd3_1 hold125 (.A(\m_sys.m_ram.m_ram.r_mem[10][3] ),
    .X(net1778));
 sg13g2_dlygate4sd3_1 hold126 (.A(\m_sys.m_ram.m_ram.r_mem[27][8] ),
    .X(net1779));
 sg13g2_dlygate4sd3_1 hold127 (.A(\m_sys.m_ram.m_ram.r_mem[5][7] ),
    .X(net1780));
 sg13g2_dlygate4sd3_1 hold128 (.A(\m_sys.m_ram.m_ram.r_mem[2][12] ),
    .X(net1781));
 sg13g2_dlygate4sd3_1 hold129 (.A(\m_sys.m_ram.m_ram.r_mem[4][12] ),
    .X(net1782));
 sg13g2_dlygate4sd3_1 hold130 (.A(\m_sys.m_ram.m_ram.r_mem[16][0] ),
    .X(net1783));
 sg13g2_dlygate4sd3_1 hold131 (.A(\m_sys.m_ram.m_ram.r_mem[26][0] ),
    .X(net1784));
 sg13g2_dlygate4sd3_1 hold132 (.A(\m_sys.m_ram.m_ram.r_mem[29][3] ),
    .X(net1785));
 sg13g2_dlygate4sd3_1 hold133 (.A(\m_sys.m_ram.m_ram.r_mem[30][11] ),
    .X(net1786));
 sg13g2_dlygate4sd3_1 hold134 (.A(\m_sys.m_ram.m_ram.r_mem[13][2] ),
    .X(net1787));
 sg13g2_dlygate4sd3_1 hold135 (.A(\m_sys.m_ram.m_ram.r_mem[11][0] ),
    .X(net1788));
 sg13g2_dlygate4sd3_1 hold136 (.A(\m_sys.m_ram.m_ram.r_mem[6][5] ),
    .X(net1789));
 sg13g2_dlygate4sd3_1 hold137 (.A(\m_sys.m_ram.m_ram.r_mem[23][4] ),
    .X(net1790));
 sg13g2_dlygate4sd3_1 hold138 (.A(\m_sys.m_ram.m_ram.r_mem[31][7] ),
    .X(net1791));
 sg13g2_dlygate4sd3_1 hold139 (.A(\m_sys.m_ram.m_ram.r_mem[19][12] ),
    .X(net1792));
 sg13g2_dlygate4sd3_1 hold140 (.A(\m_sys.m_ram.m_ram.r_mem[26][15] ),
    .X(net1793));
 sg13g2_dlygate4sd3_1 hold141 (.A(\m_sys.m_ram.m_ram.r_mem[1][2] ),
    .X(net1794));
 sg13g2_dlygate4sd3_1 hold142 (.A(\m_sys.m_ram.m_ram.r_mem[23][14] ),
    .X(net1795));
 sg13g2_dlygate4sd3_1 hold143 (.A(\m_sys.m_ram.m_ram.r_mem[10][5] ),
    .X(net1796));
 sg13g2_dlygate4sd3_1 hold144 (.A(\m_sys.m_ram.m_ram.r_mem[23][8] ),
    .X(net1797));
 sg13g2_dlygate4sd3_1 hold145 (.A(\m_sys.m_ram.m_ram.r_mem[22][4] ),
    .X(net1798));
 sg13g2_dlygate4sd3_1 hold146 (.A(_00075_),
    .X(net1799));
 sg13g2_dlygate4sd3_1 hold147 (.A(_00172_),
    .X(net1800));
 sg13g2_dlygate4sd3_1 hold148 (.A(\m_sys.m_ram.m_ram.r_mem[20][10] ),
    .X(net1801));
 sg13g2_dlygate4sd3_1 hold149 (.A(\m_sys.m_ram.m_ram.r_mem[29][9] ),
    .X(net1802));
 sg13g2_dlygate4sd3_1 hold150 (.A(\m_sys.m_ram.m_ram.r_mem[19][5] ),
    .X(net1803));
 sg13g2_dlygate4sd3_1 hold151 (.A(\m_sys.m_ram.m_ram.r_mem[25][1] ),
    .X(net1804));
 sg13g2_dlygate4sd3_1 hold152 (.A(\m_sys.m_ram.m_ram.r_mem[9][2] ),
    .X(net1805));
 sg13g2_dlygate4sd3_1 hold153 (.A(\m_sys.m_ram.m_ram.r_mem[26][6] ),
    .X(net1806));
 sg13g2_dlygate4sd3_1 hold154 (.A(\m_sys.m_ram.m_ram.r_mem[28][9] ),
    .X(net1807));
 sg13g2_dlygate4sd3_1 hold155 (.A(\m_sys.m_ram.m_ram.r_mem[5][1] ),
    .X(net1808));
 sg13g2_dlygate4sd3_1 hold156 (.A(\m_sys.m_ram.m_ram.r_mem[16][8] ),
    .X(net1809));
 sg13g2_dlygate4sd3_1 hold157 (.A(\m_sys.m_ram.m_ram.r_mem[31][15] ),
    .X(net1810));
 sg13g2_dlygate4sd3_1 hold158 (.A(\m_sys.m_ram.m_ram.r_mem[10][4] ),
    .X(net1811));
 sg13g2_dlygate4sd3_1 hold159 (.A(\m_sys.m_ram.m_ram.r_mem[10][8] ),
    .X(net1812));
 sg13g2_dlygate4sd3_1 hold160 (.A(\m_sys.m_ram.m_ram.r_mem[19][7] ),
    .X(net1813));
 sg13g2_dlygate4sd3_1 hold161 (.A(\m_sys.m_ram.m_ram.r_mem[16][12] ),
    .X(net1814));
 sg13g2_dlygate4sd3_1 hold162 (.A(\m_sys.m_ram.m_ram.r_mem[1][3] ),
    .X(net1815));
 sg13g2_dlygate4sd3_1 hold163 (.A(\m_sys.m_ram.m_ram.r_mem[28][8] ),
    .X(net1816));
 sg13g2_dlygate4sd3_1 hold164 (.A(\m_sys.m_ram.m_ram.r_mem[12][13] ),
    .X(net1817));
 sg13g2_dlygate4sd3_1 hold165 (.A(\m_sys.m_ram.m_ram.r_mem[8][3] ),
    .X(net1818));
 sg13g2_dlygate4sd3_1 hold166 (.A(\m_sys.m_ram.m_ram.r_mem[27][6] ),
    .X(net1819));
 sg13g2_dlygate4sd3_1 hold167 (.A(\m_sys.m_ram.m_ram.r_mem[14][9] ),
    .X(net1820));
 sg13g2_dlygate4sd3_1 hold168 (.A(\m_sys.m_ram.m_ram.r_mem[15][8] ),
    .X(net1821));
 sg13g2_dlygate4sd3_1 hold169 (.A(\m_sys.m_ram.m_ram.r_mem[7][5] ),
    .X(net1822));
 sg13g2_dlygate4sd3_1 hold170 (.A(\m_sys.m_ram.m_ram.r_mem[20][7] ),
    .X(net1823));
 sg13g2_dlygate4sd3_1 hold171 (.A(\m_sys.m_ram.m_ram.r_mem[17][15] ),
    .X(net1824));
 sg13g2_dlygate4sd3_1 hold172 (.A(\m_sys.m_ram.m_ram.r_mem[14][8] ),
    .X(net1825));
 sg13g2_dlygate4sd3_1 hold173 (.A(\m_sys.m_ram.m_ram.r_mem[15][9] ),
    .X(net1826));
 sg13g2_dlygate4sd3_1 hold174 (.A(\m_sys.m_ram.m_ram.r_mem[19][6] ),
    .X(net1827));
 sg13g2_dlygate4sd3_1 hold175 (.A(\m_sys.m_ram.m_ram.r_mem[29][14] ),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold176 (.A(\m_sys.m_ram.m_ram.r_mem[11][1] ),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold177 (.A(\m_sys.m_ram.m_ram.r_mem[4][4] ),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold178 (.A(\m_sys.m_ram.m_ram.r_mem[31][10] ),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold179 (.A(\m_sys.m_ram.m_ram.r_mem[18][11] ),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold180 (.A(\m_sys.m_ram.m_ram.r_mem[29][6] ),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold181 (.A(\m_sys.m_ram.m_ram.r_mem[14][0] ),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold182 (.A(\m_sys.m_ram.m_ram.r_mem[7][3] ),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold183 (.A(\m_sys.m_ram.m_ram.r_mem[0][13] ),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold184 (.A(\m_sys.m_ram.m_ram.r_mem[24][10] ),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold185 (.A(\m_sys.m_ram.m_ram.r_mem[23][0] ),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold186 (.A(\m_sys.m_ram.m_ram.r_mem[10][13] ),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold187 (.A(\m_sys.m_ram.m_ram.r_mem[25][9] ),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold188 (.A(\m_sys.m_ram.m_ram.r_mem[30][13] ),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold189 (.A(\m_sys.m_ram.m_ram.r_mem[24][6] ),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold190 (.A(\m_sys.m_ram.m_ram.r_mem[24][7] ),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold191 (.A(\m_sys.m_ram.m_ram.r_mem[12][1] ),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold192 (.A(\m_sys.m_ram.m_ram.r_mem[28][1] ),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold193 (.A(\m_sys.m_ram.m_ram.r_mem[2][6] ),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold194 (.A(\m_sys.m_ram.m_ram.r_mem[3][13] ),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold195 (.A(\m_sys.m_ram.m_ram.r_mem[28][7] ),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold196 (.A(\m_sys.m_ram.m_ram.r_mem[2][11] ),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold197 (.A(\m_sys.m_ram.m_ram.r_mem[7][4] ),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold198 (.A(\m_sys.m_ram.m_ram.r_mem[31][14] ),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold199 (.A(\m_sys.m_ram.m_ram.r_mem[0][11] ),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold200 (.A(\m_sys.m_ram.m_ram.r_mem[31][1] ),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold201 (.A(\m_sys.m_ram.m_ram.r_mem[8][15] ),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold202 (.A(\m_sys.m_ram.m_ram.r_mem[29][7] ),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold203 (.A(\m_sys.m_ram.m_ram.r_mem[1][8] ),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold204 (.A(\m_sys.m_ram.m_ram.r_mem[5][5] ),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold205 (.A(\m_sys.m_ram.m_ram.r_mem[27][13] ),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold206 (.A(\m_sys.m_ram.m_ram.r_mem[13][9] ),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold207 (.A(\m_sys.m_ram.m_ram.r_mem[30][1] ),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold208 (.A(\m_sys.m_ram.m_ram.r_mem[17][2] ),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold209 (.A(\m_sys.m_ram.m_ram.r_mem[23][15] ),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold210 (.A(\m_sys.m_ram.m_ram.r_mem[16][2] ),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold211 (.A(\m_sys.m_ram.m_ram.r_mem[8][13] ),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold212 (.A(\m_sys.m_ram.m_ram.r_mem[20][0] ),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold213 (.A(_00064_),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold214 (.A(_06366_),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold215 (.A(_01086_),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold216 (.A(\m_sys.m_ram.m_ram.r_mem[2][7] ),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold217 (.A(\m_sys.m_ram.m_ram.r_mem[22][5] ),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold218 (.A(\m_sys.m_ram.m_ram.r_mem[18][1] ),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold219 (.A(\m_sys.m_ram.m_ram.r_mem[23][11] ),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold220 (.A(\m_sys.m_ram.m_ram.r_mem[1][0] ),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold221 (.A(\m_sys.m_ram.m_ram.r_mem[22][2] ),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold222 (.A(\m_sys.m_ram.m_ram.r_mem[30][12] ),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold223 (.A(\m_sys.m_ram.m_ram.r_mem[7][11] ),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold224 (.A(\m_sys.m_ram.m_ram.r_mem[15][15] ),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold225 (.A(\m_sys.m_ram.m_ram.r_mem[25][0] ),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold226 (.A(\m_sys.m_ram.m_ram.r_mem[30][2] ),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold227 (.A(\m_sys.m_ram.m_ram.r_mem[21][10] ),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold228 (.A(\m_sys.m_ram.m_ram.r_mem[2][8] ),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold229 (.A(\m_sys.m_ram.m_ram.r_mem[4][10] ),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold230 (.A(\m_sys.m_ram.m_ram.r_mem[24][1] ),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold231 (.A(\m_sys.m_ram.m_ram.r_mem[2][4] ),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold232 (.A(\m_sys.m_ram.m_ram.r_mem[17][1] ),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold233 (.A(\m_sys.m_ram.m_ram.r_mem[22][0] ),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold234 (.A(\m_sys.m_ram.m_ram.r_mem[23][13] ),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold235 (.A(\m_sys.m_ram.m_ram.r_mem[9][15] ),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold236 (.A(\m_sys.m_ram.m_ram.r_mem[12][4] ),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold237 (.A(\m_sys.m_ram.m_ram.r_mem[21][5] ),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold238 (.A(\m_sys.m_ram.m_ram.r_mem[13][5] ),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold239 (.A(\m_sys.m_ram.m_ram.r_mem[24][4] ),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold240 (.A(\m_sys.m_ram.m_ram.r_mem[16][15] ),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold241 (.A(\m_sys.m_ram.m_ram.r_mem[29][10] ),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold242 (.A(\m_sys.m_ram.m_ram.r_mem[25][12] ),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold243 (.A(\m_sys.m_ram.m_ram.r_mem[22][11] ),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold244 (.A(\m_sys.m_ram.m_ram.r_mem[12][6] ),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold245 (.A(\m_sys.m_ram.m_ram.r_mem[13][1] ),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold246 (.A(\m_sys.m_ram.m_ram.r_mem[16][9] ),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold247 (.A(\m_sys.m_ram.m_ram.r_mem[26][4] ),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold248 (.A(\m_sys.m_ram.m_ram.r_mem[14][6] ),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold249 (.A(\m_sys.m_ram.m_ram.r_mem[12][10] ),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold250 (.A(\m_sys.m_ram.m_ram.r_mem[18][14] ),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold251 (.A(\m_sys.m_ram.m_ram.r_mem[30][0] ),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold252 (.A(\m_sys.m_ram.m_ram.r_mem[11][15] ),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold253 (.A(\m_sys.m_ram.m_ram.r_mem[23][10] ),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold254 (.A(\m_sys.m_ram.m_ram.r_mem[4][14] ),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold255 (.A(\m_sys.m_ram.m_ram.r_mem[20][11] ),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold256 (.A(\m_sys.m_ram.m_ram.r_mem[9][4] ),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold257 (.A(\m_sys.m_ram.m_ram.r_mem[13][10] ),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold258 (.A(\m_sys.m_ram.m_ram.r_mem[17][13] ),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold259 (.A(\m_sys.m_ram.m_ram.r_mem[17][5] ),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold260 (.A(\m_sys.m_ram.m_ram.r_mem[20][8] ),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold261 (.A(\m_sys.m_ram.m_ram.r_mem[6][7] ),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold262 (.A(\m_sys.m_ram.m_ram.r_mem[0][5] ),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold263 (.A(\m_sys.m_ram.m_ram.r_mem[6][11] ),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold264 (.A(\m_sys.m_ram.m_ram.r_mem[8][9] ),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold265 (.A(\m_sys.m_ram.m_ram.r_mem[10][7] ),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold266 (.A(\m_sys.m_ram.m_ram.r_mem[30][3] ),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold267 (.A(\m_sys.m_ram.m_ram.r_mem[1][14] ),
    .X(net1920));
 sg13g2_dlygate4sd3_1 hold268 (.A(\m_sys.m_ram.m_ram.r_mem[21][0] ),
    .X(net1921));
 sg13g2_dlygate4sd3_1 hold269 (.A(\m_sys.m_ram.m_ram.r_mem[5][14] ),
    .X(net1922));
 sg13g2_dlygate4sd3_1 hold270 (.A(\m_sys.m_ram.m_ram.r_mem[21][7] ),
    .X(net1923));
 sg13g2_dlygate4sd3_1 hold271 (.A(\m_sys.m_ram.m_ram.r_mem[6][3] ),
    .X(net1924));
 sg13g2_dlygate4sd3_1 hold272 (.A(\m_sys.m_ram.m_ram.r_mem[24][13] ),
    .X(net1925));
 sg13g2_dlygate4sd3_1 hold273 (.A(\m_sys.m_ram.m_ram.r_mem[31][11] ),
    .X(net1926));
 sg13g2_dlygate4sd3_1 hold274 (.A(\m_sys.m_ram.m_ram.r_mem[30][5] ),
    .X(net1927));
 sg13g2_dlygate4sd3_1 hold275 (.A(\m_sys.m_ram.m_ram.r_mem[13][6] ),
    .X(net1928));
 sg13g2_dlygate4sd3_1 hold276 (.A(\m_sys.m_ram.m_ram.r_mem[20][4] ),
    .X(net1929));
 sg13g2_dlygate4sd3_1 hold277 (.A(\m_sys.m_ram.m_ram.r_mem[31][3] ),
    .X(net1930));
 sg13g2_dlygate4sd3_1 hold278 (.A(\m_sys.m_ram.m_ram.r_mem[15][13] ),
    .X(net1931));
 sg13g2_dlygate4sd3_1 hold279 (.A(\m_sys.m_ram.m_ram.r_mem[19][3] ),
    .X(net1932));
 sg13g2_dlygate4sd3_1 hold280 (.A(\m_sys.m_ram.m_ram.r_mem[26][5] ),
    .X(net1933));
 sg13g2_dlygate4sd3_1 hold281 (.A(\m_sys.m_ram.m_ram.r_mem[5][4] ),
    .X(net1934));
 sg13g2_dlygate4sd3_1 hold282 (.A(\m_sys.m_ram.m_ram.r_mem[27][1] ),
    .X(net1935));
 sg13g2_dlygate4sd3_1 hold283 (.A(\m_sys.m_ram.m_ram.r_mem[9][6] ),
    .X(net1936));
 sg13g2_dlygate4sd3_1 hold284 (.A(\m_sys.m_ram.m_ram.r_mem[9][10] ),
    .X(net1937));
 sg13g2_dlygate4sd3_1 hold285 (.A(\m_sys.m_ram.m_ram.r_mem[22][9] ),
    .X(net1938));
 sg13g2_dlygate4sd3_1 hold286 (.A(\m_sys.m_ram.m_ram.r_mem[3][8] ),
    .X(net1939));
 sg13g2_dlygate4sd3_1 hold287 (.A(\m_sys.m_ram.m_ram.r_mem[6][4] ),
    .X(net1940));
 sg13g2_dlygate4sd3_1 hold288 (.A(\m_sys.m_ram.m_ram.r_mem[24][12] ),
    .X(net1941));
 sg13g2_dlygate4sd3_1 hold289 (.A(\m_sys.m_ram.m_ram.r_mem[28][15] ),
    .X(net1942));
 sg13g2_dlygate4sd3_1 hold290 (.A(\m_sys.m_ram.m_ram.r_mem[0][9] ),
    .X(net1943));
 sg13g2_dlygate4sd3_1 hold291 (.A(\m_sys.m_ram.m_ram.r_mem[4][13] ),
    .X(net1944));
 sg13g2_dlygate4sd3_1 hold292 (.A(\m_sys.m_ram.m_ram.r_mem[4][3] ),
    .X(net1945));
 sg13g2_dlygate4sd3_1 hold293 (.A(\m_sys.m_ram.m_ram.r_mem[27][10] ),
    .X(net1946));
 sg13g2_dlygate4sd3_1 hold294 (.A(\m_sys.m_ram.m_ram.r_mem[31][2] ),
    .X(net1947));
 sg13g2_dlygate4sd3_1 hold295 (.A(\m_sys.m_ram.m_ram.r_mem[27][9] ),
    .X(net1948));
 sg13g2_dlygate4sd3_1 hold296 (.A(\m_sys.m_ram.m_ram.r_mem[4][11] ),
    .X(net1949));
 sg13g2_dlygate4sd3_1 hold297 (.A(\m_sys.m_ram.m_ram.r_mem[27][7] ),
    .X(net1950));
 sg13g2_dlygate4sd3_1 hold298 (.A(\m_sys.m_ram.m_ram.r_mem[8][11] ),
    .X(net1951));
 sg13g2_dlygate4sd3_1 hold299 (.A(\m_sys.m_ram.m_ram.r_mem[19][8] ),
    .X(net1952));
 sg13g2_dlygate4sd3_1 hold300 (.A(\m_sys.m_ram.m_ram.r_mem[10][12] ),
    .X(net1953));
 sg13g2_dlygate4sd3_1 hold301 (.A(\m_sys.m_ram.m_ram.r_mem[18][5] ),
    .X(net1954));
 sg13g2_dlygate4sd3_1 hold302 (.A(\m_sys.m_ram.m_ram.r_mem[19][1] ),
    .X(net1955));
 sg13g2_dlygate4sd3_1 hold303 (.A(\m_sys.m_ram.m_ram.r_mem[26][12] ),
    .X(net1956));
 sg13g2_dlygate4sd3_1 hold304 (.A(\m_sys.m_ram.m_ram.r_mem[7][0] ),
    .X(net1957));
 sg13g2_dlygate4sd3_1 hold305 (.A(\m_sys.m_ram.m_ram.r_mem[28][5] ),
    .X(net1958));
 sg13g2_dlygate4sd3_1 hold306 (.A(\m_sys.m_ram.m_ram.r_mem[3][12] ),
    .X(net1959));
 sg13g2_dlygate4sd3_1 hold307 (.A(\m_sys.m_ram.m_ram.r_mem[29][5] ),
    .X(net1960));
 sg13g2_dlygate4sd3_1 hold308 (.A(\m_sys.m_ram.m_ram.r_mem[9][11] ),
    .X(net1961));
 sg13g2_dlygate4sd3_1 hold309 (.A(\m_sys.m_ram.m_ram.r_mem[26][10] ),
    .X(net1962));
 sg13g2_dlygate4sd3_1 hold310 (.A(\m_sys.m_ram.m_ram.r_mem[15][2] ),
    .X(net1963));
 sg13g2_dlygate4sd3_1 hold311 (.A(\m_sys.m_core.m_gpr._GEN[220] ),
    .X(net1964));
 sg13g2_dlygate4sd3_1 hold312 (.A(_01660_),
    .X(net1965));
 sg13g2_dlygate4sd3_1 hold313 (.A(\m_sys.m_ram.m_ram.r_mem[15][3] ),
    .X(net1966));
 sg13g2_dlygate4sd3_1 hold314 (.A(\m_sys.m_ram.m_ram.r_mem[26][3] ),
    .X(net1967));
 sg13g2_dlygate4sd3_1 hold315 (.A(\m_sys.m_ram.m_ram.r_mem[7][1] ),
    .X(net1968));
 sg13g2_dlygate4sd3_1 hold316 (.A(\m_sys.m_ram.m_ram.r_mem[26][14] ),
    .X(net1969));
 sg13g2_dlygate4sd3_1 hold317 (.A(\m_sys.m_ram.m_ram.r_mem[6][13] ),
    .X(net1970));
 sg13g2_dlygate4sd3_1 hold318 (.A(\m_sys.m_ram.m_ram.r_mem[25][6] ),
    .X(net1971));
 sg13g2_dlygate4sd3_1 hold319 (.A(\m_sys.m_ram.m_ram.r_mem[26][1] ),
    .X(net1972));
 sg13g2_dlygate4sd3_1 hold320 (.A(\m_sys.m_ram.m_ram.r_mem[3][6] ),
    .X(net1973));
 sg13g2_dlygate4sd3_1 hold321 (.A(\m_sys.m_ram.m_ram.r_mem[6][10] ),
    .X(net1974));
 sg13g2_dlygate4sd3_1 hold322 (.A(\m_sys.m_ram.m_ram.r_mem[17][3] ),
    .X(net1975));
 sg13g2_dlygate4sd3_1 hold323 (.A(\m_sys.m_ram.m_ram.r_mem[5][13] ),
    .X(net1976));
 sg13g2_dlygate4sd3_1 hold324 (.A(\m_sys.m_ram.m_ram.r_mem[31][6] ),
    .X(net1977));
 sg13g2_dlygate4sd3_1 hold325 (.A(\m_sys.m_ram.m_ram.r_mem[5][10] ),
    .X(net1978));
 sg13g2_dlygate4sd3_1 hold326 (.A(\m_sys.m_ram.m_ram.r_mem[23][2] ),
    .X(net1979));
 sg13g2_dlygate4sd3_1 hold327 (.A(\m_sys.m_core.m_gpr._GEN[64] ),
    .X(net1980));
 sg13g2_dlygate4sd3_1 hold328 (.A(_01535_),
    .X(net1981));
 sg13g2_dlygate4sd3_1 hold329 (.A(\m_sys.m_ram.m_ram.r_mem[16][6] ),
    .X(net1982));
 sg13g2_dlygate4sd3_1 hold330 (.A(\m_sys.m_ram.m_ram.r_mem[19][13] ),
    .X(net1983));
 sg13g2_dlygate4sd3_1 hold331 (.A(\m_sys.m_ram.m_ram.r_mem[13][12] ),
    .X(net1984));
 sg13g2_dlygate4sd3_1 hold332 (.A(\m_sys.m_ram.m_ram.r_mem[10][15] ),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold333 (.A(\m_sys.m_ram.m_ram.r_mem[1][4] ),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold334 (.A(\m_sys.m_ram.m_ram.r_mem[15][1] ),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold335 (.A(\m_sys.m_ram.m_ram.r_mem[20][13] ),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold336 (.A(\m_sys.m_ram.m_ram.r_mem[27][14] ),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold337 (.A(\m_sys.m_ram.m_ram.r_mem[18][4] ),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold338 (.A(\m_sys.m_ram.m_ram.r_mem[27][3] ),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold339 (.A(\m_sys.m_bootloader._GEN_22[1] ),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold340 (.A(_01057_),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold341 (.A(\m_sys.m_ram.m_ram.r_mem[14][15] ),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold342 (.A(\m_sys.m_ram.m_ram.r_mem[28][10] ),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold343 (.A(\m_sys.m_ram.m_ram.r_mem[20][9] ),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold344 (.A(\m_sys.m_ram.m_ram.r_mem[31][12] ),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold345 (.A(\m_sys.m_ram.m_ram.r_mem[10][0] ),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold346 (.A(\m_sys.m_ram.m_ram.r_mem[25][4] ),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold347 (.A(\m_sys.m_ram.m_ram.r_mem[6][6] ),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold348 (.A(\m_sys.m_ram.m_ram.r_mem[6][12] ),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold349 (.A(\m_sys.m_ram.m_ram.r_mem[3][7] ),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold350 (.A(\m_sys.m_ram.m_ram.r_mem[2][10] ),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold351 (.A(\m_sys.m_ram.m_ram.r_mem[0][12] ),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold352 (.A(\m_sys.m_ram.m_ram.r_mem[9][13] ),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold353 (.A(\m_sys.m_ram.m_ram.r_mem[14][10] ),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold354 (.A(\m_sys.m_core.m_gpr._GEN[211] ),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold355 (.A(\m_sys.m_ram.m_ram.r_mem[22][3] ),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold356 (.A(\m_sys.m_ram.m_ram.r_mem[31][9] ),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold357 (.A(\m_sys.m_uart.r_rx_data[1] ),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold358 (.A(_07412_),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold359 (.A(\m_sys.m_ram.m_ram.r_mem[18][13] ),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold360 (.A(\m_sys.m_ram.m_ram.r_mem[4][2] ),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold361 (.A(\m_sys.m_core.m_gpr._GEN[83] ),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold362 (.A(\m_sys.m_ram.m_ram.r_mem[14][12] ),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold363 (.A(\m_sys.m_ram.m_ram.r_mem[9][12] ),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold364 (.A(\m_sys.m_ram.m_ram.r_mem[2][1] ),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold365 (.A(\m_sys.m_ram.m_ram.r_mem[23][1] ),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold366 (.A(\m_sys.m_ram.m_ram.r_mem[6][9] ),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold367 (.A(\m_sys.m_ram.m_ram.r_mem[23][9] ),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold368 (.A(\m_sys.m_ram.m_ram.r_mem[24][9] ),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold369 (.A(\m_sys.m_ram.m_ram.r_mem[25][8] ),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold370 (.A(\m_sys.m_ram.m_ram.r_mem[4][7] ),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold371 (.A(\m_sys.m_ram.m_ram.r_mem[0][8] ),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold372 (.A(\m_sys.m_ram.m_ram.r_mem[19][10] ),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold373 (.A(\m_sys.m_ram.m_ram.r_mem[10][11] ),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold374 (.A(\m_sys.m_ram.m_ram.r_mem[27][11] ),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold375 (.A(\m_sys.m_ram.m_ram.r_mem[22][12] ),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold376 (.A(\m_sys.m_ram.m_ram.r_mem[31][4] ),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold377 (.A(\m_sys.m_ram.m_ram.r_mem[2][2] ),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold378 (.A(\m_sys.m_core.m_gpr._GEN[32] ),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold379 (.A(_01567_),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold380 (.A(\m_sys.m_ram.m_ram.r_mem[18][12] ),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold381 (.A(\m_sys.m_ram.m_ram.r_mem[2][5] ),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold382 (.A(\m_sys.m_ram.m_ram.r_mem[4][1] ),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold383 (.A(\m_sys.m_ram.m_ram.r_mem[11][13] ),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold384 (.A(\m_sys.m_ram.m_ram.r_mem[17][8] ),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold385 (.A(\m_sys.m_ram.m_ram.r_mem[28][13] ),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold386 (.A(\m_sys.m_ram.m_ram.r_mem[7][6] ),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold387 (.A(\m_sys.m_ram.m_ram.r_mem[13][8] ),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold388 (.A(\m_sys.m_ram.m_ram.r_mem[8][4] ),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold389 (.A(\m_sys.m_ram.m_ram.r_mem[13][14] ),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold390 (.A(\m_sys.m_ram.m_ram.r_mem[2][14] ),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold391 (.A(\m_sys.m_bootloader._GEN_22[0] ),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold392 (.A(_01056_),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold393 (.A(\m_sys.m_ram.m_ram.r_mem[1][7] ),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold394 (.A(\m_sys.m_ram.m_ram.r_mem[11][6] ),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold395 (.A(\m_sys.m_ram.m_ram.r_mem[28][0] ),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold396 (.A(\m_sys.m_ram.m_ram.r_mem[12][2] ),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold397 (.A(\m_sys.m_ram.m_ram.r_mem[20][12] ),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold398 (.A(\m_sys.m_ram.m_ram.r_mem[13][3] ),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold399 (.A(\m_sys.m_ram.m_ram.r_mem[12][8] ),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold400 (.A(\m_sys.m_ram.m_ram.r_mem[13][13] ),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold401 (.A(\m_sys.m_ram.m_ram.r_mem[14][7] ),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold402 (.A(\m_sys.m_ram.m_ram.r_mem[31][5] ),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold403 (.A(\m_sys.m_ram.m_ram.r_mem[24][3] ),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold404 (.A(\m_sys.m_ram.m_ram.r_mem[3][14] ),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold405 (.A(\m_sys.m_ram.m_ram.r_mem[30][7] ),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold406 (.A(\m_sys.m_ram.m_ram.r_mem[15][12] ),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold407 (.A(\m_sys.m_ram.m_ram.r_mem[23][12] ),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold408 (.A(\m_sys.m_ram.m_ram.r_mem[17][12] ),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold409 (.A(\m_sys.m_ram.m_ram.r_mem[15][11] ),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold410 (.A(\m_sys.m_ram.m_ram.r_mem[15][4] ),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold411 (.A(\m_sys.m_ram.m_ram.r_mem[8][7] ),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold412 (.A(\m_sys.m_ram.m_ram.r_mem[10][6] ),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold413 (.A(\m_sys.m_ram.m_ram.r_mem[3][5] ),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold414 (.A(\m_sys.m_ram.m_ram.r_mem[10][14] ),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold415 (.A(\m_sys.m_ram.m_ram.r_mem[22][15] ),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold416 (.A(\m_sys.m_ram.m_ram.r_mem[18][8] ),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold417 (.A(\m_sys.m_ram.m_ram.r_mem[7][10] ),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold418 (.A(\m_sys.m_ram.m_ram.r_mem[17][14] ),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold419 (.A(\m_sys.m_ram.m_ram.r_mem[15][10] ),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold420 (.A(\m_sys.m_ram.m_ram.r_mem[22][14] ),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold421 (.A(\m_sys.m_ram.m_ram.r_mem[13][11] ),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold422 (.A(\m_sys.m_ram.m_ram.r_mem[5][6] ),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold423 (.A(\m_sys.m_ram.m_ram.r_mem[10][1] ),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold424 (.A(\m_sys.m_ram.m_ram.r_mem[4][0] ),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold425 (.A(\m_sys.m_ram.m_ram.r_mem[18][0] ),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold426 (.A(\m_sys.m_ram.m_ram.r_mem[16][7] ),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold427 (.A(\m_sys.m_ram.m_ram.r_mem[19][0] ),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold428 (.A(\m_sys.m_ram.m_ram.r_mem[11][8] ),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold429 (.A(\m_sys.m_ram.m_ram.r_mem[8][10] ),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold430 (.A(\m_sys.m_core.m_gpr._GEN[71] ),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold431 (.A(\m_sys.m_ram.m_ram.r_mem[0][10] ),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold432 (.A(\m_sys.m_ram.m_ram.r_mem[2][0] ),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold433 (.A(\m_sys.m_ram.m_ram.r_mem[16][3] ),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold434 (.A(\m_sys.m_ram.m_ram.r_mem[17][0] ),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold435 (.A(\m_sys.m_ram.m_ram.r_mem[14][2] ),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold436 (.A(\m_sys.m_ram.m_ram.r_mem[7][14] ),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold437 (.A(\m_sys.m_ram.m_ram.r_mem[20][1] ),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold438 (.A(\m_sys.m_ram.m_ram.r_mem[30][6] ),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold439 (.A(\m_sys.m_ram.m_ram.r_mem[11][11] ),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold440 (.A(\m_sys.m_ram.m_ram.r_mem[3][10] ),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold441 (.A(\m_sys.m_ram.m_ram.r_mem[30][4] ),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold442 (.A(\m_sys.m_ram.m_ram.r_mem[21][13] ),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold443 (.A(\m_sys.m_ram.m_ram.r_mem[24][5] ),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold444 (.A(\m_sys.m_ram.m_ram.r_mem[12][11] ),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold445 (.A(\m_sys.m_ram.m_ram.r_mem[27][2] ),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold446 (.A(\m_sys.m_ram.m_ram.r_mem[27][5] ),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold447 (.A(\m_sys.m_ram.m_ram.r_mem[14][1] ),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold448 (.A(\m_sys.m_ram.m_ram.r_mem[26][9] ),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold449 (.A(\m_sys.m_ram.m_ram.r_mem[22][8] ),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold450 (.A(\m_sys.m_ram.m_ram.r_mem[13][15] ),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold451 (.A(\m_sys.m_ram.m_ram.r_mem[15][6] ),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold452 (.A(\m_sys.m_ram.m_ram.r_mem[31][0] ),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold453 (.A(\m_sys.m_ram.m_ram.r_mem[11][14] ),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold454 (.A(\m_sys.m_ram.m_ram.r_mem[11][9] ),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold455 (.A(\m_sys.m_ram.m_ram.r_mem[16][10] ),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold456 (.A(\m_sys.m_core.m_gpr._GEN[212] ),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold457 (.A(\m_sys.m_ram.m_ram.r_mem[19][4] ),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold458 (.A(\m_sys.m_ram.m_ram.r_mem[30][9] ),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold459 (.A(\m_sys.m_ram.m_ram.r_mem[30][15] ),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold460 (.A(\m_sys.m_ram.m_ram.r_mem[11][4] ),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold461 (.A(\m_sys.m_ram.m_ram.r_mem[19][11] ),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold462 (.A(\m_sys.m_ram.m_ram.r_mem[8][1] ),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold463 (.A(\m_sys.m_ram.m_ram.r_mem[18][15] ),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold464 (.A(\m_sys.m_ram.m_ram.r_mem[31][13] ),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold465 (.A(\m_sys.m_ram.m_ram.r_mem[11][2] ),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold466 (.A(\m_sys.m_ram.m_ram.r_mem[11][10] ),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold467 (.A(\m_sys.m_uart.r_rx_data[7] ),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold468 (.A(_07419_),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold469 (.A(\m_sys.m_ram.m_ram.r_mem[15][14] ),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold470 (.A(\m_sys.m_uart.r_rx_data[3] ),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold471 (.A(_07414_),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold472 (.A(\m_sys.m_ram.m_ram.r_mem[9][14] ),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold473 (.A(\m_sys.m_ram.m_ram.r_mem[11][3] ),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold474 (.A(\m_sys.m_ram.m_ram.r_mem[9][28] ),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold475 (.A(\m_sys.m_ram.m_ram.r_mem[18][9] ),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold476 (.A(\m_sys.m_ram.m_ram.r_mem[11][5] ),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold477 (.A(\m_sys.m_core.m_gpr._GEN[94] ),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold478 (.A(_01565_),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold479 (.A(\m_sys.m_ram.m_ram.r_mem[22][13] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold480 (.A(\m_sys.m_ram.m_ram.r_mem[6][14] ),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold481 (.A(\m_sys.m_core.m_gpr._GEN[92] ),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold482 (.A(_01563_),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold483 (.A(\m_sys.m_ram.m_ram.r_mem[15][5] ),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold484 (.A(\m_sys.m_core.m_gpr._GEN[85] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold485 (.A(\m_sys.m_ram.m_ram.r_mem[0][15] ),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold486 (.A(\m_sys.m_ram.m_ram.r_mem[28][11] ),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold487 (.A(\m_sys.m_ram.m_ram.r_mem[14][5] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold488 (.A(\m_sys.m_ram.m_ram.r_mem[22][10] ),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold489 (.A(\m_sys.m_ram.m_ram.r_mem[7][13] ),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold490 (.A(\m_sys.m_ram.m_ram.r_mem[5][3] ),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold491 (.A(\m_sys.m_ram.m_ram.r_mem[3][4] ),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold492 (.A(\m_sys.m_ram.m_ram.r_mem[18][3] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold493 (.A(\m_sys.m_ram.m_ram.r_mem[21][25] ),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold494 (.A(\m_sys.m_ram.m_ram.r_mem[25][28] ),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold495 (.A(\m_sys.m_ram.m_ram.r_mem[0][7] ),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold496 (.A(\m_sys.m_ram.m_ram.r_mem[13][16] ),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold497 (.A(\m_sys.m_ram.m_ram.r_mem[17][10] ),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold498 (.A(\m_sys.m_ram.m_ram.r_mem[12][5] ),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold499 (.A(\m_sys.m_ram.m_ram.r_mem[26][7] ),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold500 (.A(\m_sys.m_ram.m_ram.r_mem[7][15] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold501 (.A(\m_sys.m_ram.m_ram.r_mem[6][28] ),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold502 (.A(\m_sys.m_ram.m_ram.r_mem[3][11] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold503 (.A(\m_sys.m_ram.m_ram.r_mem[25][27] ),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold504 (.A(\m_sys.m_ram.m_ram.r_mem[24][2] ),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold505 (.A(\m_sys.m_ram.m_ram.r_mem[1][19] ),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold506 (.A(\m_sys.m_ram.m_ram.r_mem[15][0] ),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold507 (.A(\m_sys.m_ram.m_ram.r_mem[10][28] ),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold508 (.A(\m_sys.m_ram.m_ram.r_mem[13][7] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold509 (.A(\m_sys.m_ram.m_ram.r_mem[20][2] ),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold510 (.A(\m_sys.m_ram.m_ram.r_mem[27][4] ),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold511 (.A(\m_sys.m_ram.m_ram.r_mem[26][8] ),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold512 (.A(\m_sys.m_ram.m_ram.r_mem[18][24] ),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold513 (.A(\m_sys.m_ram.m_ram.r_mem[8][22] ),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold514 (.A(\m_sys.m_ram.m_ram.r_mem[30][22] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold515 (.A(\m_sys.m_ram.m_ram.r_mem[11][12] ),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold516 (.A(\m_sys.m_ram.m_ram.r_mem[4][9] ),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold517 (.A(\m_sys.m_ram.m_ram.r_mem[24][14] ),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold518 (.A(\m_sys.m_ram.m_ram.r_mem[12][3] ),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold519 (.A(\m_sys.m_ram.m_ram.r_mem[26][26] ),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold520 (.A(\m_sys.m_ram.m_ram.r_mem[5][18] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold521 (.A(\m_sys.m_ram.m_ram.r_mem[21][21] ),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold522 (.A(\m_sys.m_ram.m_ram.r_mem[14][3] ),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold523 (.A(\m_sys.m_ram.m_ram.r_mem[19][15] ),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold524 (.A(\m_sys.m_ram.m_ram.r_mem[6][25] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold525 (.A(\m_sys.m_ram.m_ram.r_mem[7][9] ),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold526 (.A(\m_sys.m_ram.m_ram.r_mem[2][3] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold527 (.A(\m_sys.m_ram.m_ram.r_mem[24][0] ),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold528 (.A(\m_sys.m_ram.m_ram.r_mem[6][21] ),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold529 (.A(\m_sys.m_ram.m_ram.r_mem[26][23] ),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold530 (.A(\m_sys.m_ram.m_ram.r_mem[3][1] ),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold531 (.A(\m_sys.m_ram.m_ram.r_mem[24][20] ),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold532 (.A(\m_sys.m_core.m_gpr._GEN[93] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold533 (.A(\m_sys.m_ram.m_ram.r_mem[6][16] ),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold534 (.A(\m_sys.m_ram.m_ram.r_mem[4][31] ),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold535 (.A(\m_sys.m_ram.m_ram.r_mem[27][0] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold536 (.A(\m_sys.m_ram.m_ram.r_mem[25][26] ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold537 (.A(\m_sys.m_ram.m_ram.r_mem[29][13] ),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold538 (.A(\m_sys.m_ram.m_ram.r_mem[29][27] ),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold539 (.A(\m_sys.m_ram.m_ram.r_mem[10][10] ),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold540 (.A(\m_sys.m_ram.m_ram.r_mem[23][7] ),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold541 (.A(\m_sys.m_ram.m_ram.r_mem[17][29] ),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold542 (.A(\m_sys.m_ram.m_ram.r_mem[24][30] ),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold543 (.A(\m_sys.m_ram.m_ram.r_mem[5][21] ),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold544 (.A(\m_sys.m_ram.m_ram.r_mem[1][20] ),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold545 (.A(\m_sys.m_ram.m_ram.r_mem[12][28] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold546 (.A(\m_sys.m_ram.m_ram.r_mem[0][4] ),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold547 (.A(\m_sys.m_ram.m_ram.r_mem[17][16] ),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold548 (.A(\m_sys.m_ram.m_ram.r_mem[4][29] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold549 (.A(\m_sys.m_ram.m_ram.r_mem[6][30] ),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold550 (.A(\m_sys.m_ram.m_ram.r_mem[16][4] ),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold551 (.A(\m_sys.m_ram.m_ram.r_mem[7][22] ),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold552 (.A(\m_sys.m_ram.m_ram.r_mem[25][29] ),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold553 (.A(\m_sys.m_ram.m_ram.r_mem[24][21] ),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold554 (.A(\m_sys.m_ram.m_ram.r_mem[7][8] ),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold555 (.A(\m_sys.m_ram.m_ram.r_mem[8][26] ),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold556 (.A(\m_sys.m_ram.m_ram.r_mem[26][18] ),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold557 (.A(\m_sys.m_ram.m_ram.r_mem[28][25] ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold558 (.A(\m_sys.m_ram.m_ram.r_mem[12][27] ),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold559 (.A(\m_sys.m_ram.m_ram.r_mem[0][20] ),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold560 (.A(\m_sys.m_ram.m_ram.r_mem[28][12] ),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold561 (.A(\m_sys.m_ram.m_ram.r_mem[14][4] ),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold562 (.A(\m_sys.m_ram.m_ram.r_mem[0][1] ),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold563 (.A(\m_sys.m_ram.m_ram.r_mem[21][27] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold564 (.A(\m_sys.m_ram.m_ram.r_mem[17][24] ),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold565 (.A(\m_sys.m_ram.m_ram.r_mem[11][18] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold566 (.A(\m_sys.m_ram.m_ram.r_mem[25][21] ),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold567 (.A(\m_sys.m_ram.m_ram.r_mem[10][9] ),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold568 (.A(\m_sys.m_ram.m_ram.r_mem[12][20] ),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold569 (.A(\m_sys.m_ram.m_ram.r_mem[5][15] ),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold570 (.A(\m_sys.m_ram.m_ram.r_mem[21][26] ),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold571 (.A(\m_sys.m_core.m_gpr._GEN[187] ),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold572 (.A(\m_sys.m_ram.m_ram.r_mem[4][6] ),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold573 (.A(\m_sys.m_ram.m_ram.r_mem[28][28] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold574 (.A(\m_sys.m_ram.m_ram.r_mem[5][8] ),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold575 (.A(\m_sys.m_ram.m_ram.r_mem[13][24] ),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold576 (.A(\m_sys.m_ram.m_ram.r_mem[22][31] ),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold577 (.A(\m_sys.m_ram.m_ram.r_mem[20][26] ),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold578 (.A(\m_sys.m_ram.m_ram.r_mem[11][7] ),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold579 (.A(\m_sys.m_core.m_gpr._GEN[221] ),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold580 (.A(\m_sys.m_ram.m_ram.r_mem[2][24] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold581 (.A(\m_sys.m_ram.m_ram.r_mem[6][17] ),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold582 (.A(\m_sys.m_ram.m_ram.r_mem[2][29] ),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold583 (.A(\m_sys.m_core.m_gpr._GEN[216] ),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold584 (.A(\m_sys.m_ram.m_ram.r_mem[25][14] ),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold585 (.A(\m_sys.m_ram.m_ram.r_mem[3][16] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold586 (.A(\m_sys.m_ram.m_ram.r_mem[29][11] ),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold587 (.A(\m_sys.m_ram.m_ram.r_mem[20][28] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold588 (.A(\m_sys.m_ram.m_ram.r_mem[5][17] ),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold589 (.A(\m_sys.m_ram.m_ram.r_mem[13][28] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold590 (.A(\m_sys.m_ram.m_ram.r_mem[19][14] ),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold591 (.A(\m_sys.m_ram.m_ram.r_mem[30][18] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold592 (.A(\m_sys.m_ram.m_ram.r_mem[7][2] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold593 (.A(\m_sys.m_ram.m_ram.r_mem[5][19] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold594 (.A(\m_sys.m_ram.m_ram.r_mem[0][19] ),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold595 (.A(\m_sys.m_ram.m_ram.r_mem[5][23] ),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold596 (.A(\m_sys.m_ram.m_ram.r_mem[23][3] ),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold597 (.A(\m_sys.m_ram.m_ram.r_mem[29][23] ),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold598 (.A(\m_sys.m_ram.m_ram.r_mem[23][19] ),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold599 (.A(\m_sys.m_ram.m_ram.r_mem[29][2] ),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold600 (.A(\m_sys.m_ram.m_ram.r_mem[2][21] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold601 (.A(\m_sys.m_ram.m_ram.r_mem[29][28] ),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold602 (.A(\m_sys.m_ram.m_ram.r_mem[29][18] ),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold603 (.A(\m_sys.m_ram.m_ram.r_mem[28][20] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold604 (.A(\m_sys.m_core.m_gpr._GEN[178] ),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold605 (.A(\m_sys.m_ram.m_ram.r_mem[21][28] ),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold606 (.A(\m_sys.m_ram.m_ram.r_mem[21][29] ),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold607 (.A(\m_sys.m_ram.m_ram.r_mem[29][24] ),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold608 (.A(\m_sys.m_ram.m_ram.r_mem[20][24] ),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold609 (.A(\m_sys.m_core.m_gpr._GEN[218] ),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold610 (.A(\m_sys.m_ram.m_ram.r_mem[18][26] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold611 (.A(\m_sys.m_ram.m_ram.r_mem[19][29] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold612 (.A(\m_sys.m_ram.m_ram.r_mem[3][2] ),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold613 (.A(\m_sys.m_ram.m_ram.r_mem[9][25] ),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold614 (.A(\m_sys.m_ram.m_ram.r_mem[30][28] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold615 (.A(\m_sys.m_ram.m_ram.r_mem[0][3] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold616 (.A(\m_sys.m_ram.m_ram.r_mem[21][22] ),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold617 (.A(\m_sys.m_ram.m_ram.r_mem[0][16] ),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold618 (.A(\m_sys.m_ram.m_ram.r_mem[12][30] ),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold619 (.A(\m_sys.m_ram.m_ram.r_mem[5][27] ),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold620 (.A(\m_sys.m_ram.m_ram.r_mem[7][29] ),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold621 (.A(\m_sys.m_ram.m_ram.r_mem[22][25] ),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold622 (.A(\m_sys.m_core.m_gpr._GEN[90] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold623 (.A(\m_sys.m_ram.m_ram.r_mem[0][21] ),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold624 (.A(\m_sys.m_core.m_gpr._GEN[176] ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold625 (.A(\m_sys.m_ram.m_ram.r_mem[3][0] ),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold626 (.A(\m_sys.m_ram.m_ram.r_mem[16][21] ),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold627 (.A(\m_sys.m_ram.m_ram.r_mem[30][16] ),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold628 (.A(\m_sys.m_ram.m_ram.r_mem[7][7] ),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold629 (.A(\m_sys.m_ram.m_ram.r_mem[13][27] ),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold630 (.A(\m_sys.m_ram.m_ram.r_mem[10][30] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold631 (.A(\m_sys.m_uart.m_tx.r_data[6] ),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold632 (.A(_00993_),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold633 (.A(\m_sys.m_ram.m_ram.r_mem[21][18] ),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold634 (.A(\m_sys.m_ram.m_ram.r_mem[2][20] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold635 (.A(\m_sys.m_ram.m_ram.r_mem[24][22] ),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold636 (.A(\m_sys.m_ram.m_ram.r_mem[13][20] ),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold637 (.A(\m_sys.m_ram.m_ram.r_mem[5][31] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold638 (.A(\m_sys.m_ram.m_ram.r_mem[14][17] ),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold639 (.A(\m_sys.m_ram.m_ram.r_mem[1][30] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold640 (.A(\m_sys.m_ram.m_ram.r_mem[1][29] ),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold641 (.A(\m_sys.m_ram.m_ram.r_mem[3][17] ),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold642 (.A(\m_sys.m_ram.m_ram.r_mem[15][17] ),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold643 (.A(\m_sys.m_ram.m_ram.r_mem[21][31] ),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold644 (.A(\m_sys.m_core.m_gpr._GEN[181] ),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold645 (.A(\m_sys.m_ram.m_ram.r_mem[15][31] ),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold646 (.A(\m_sys.m_ram.m_ram.r_mem[13][30] ),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold647 (.A(\m_sys.m_ram.m_ram.r_mem[9][19] ),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold648 (.A(\m_sys.m_ram.m_ram.r_mem[27][25] ),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold649 (.A(\m_sys.m_ram.m_ram.r_mem[7][20] ),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold650 (.A(\m_sys.m_ram.m_ram.r_mem[14][31] ),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold651 (.A(\m_sys.m_ram.m_ram.r_mem[9][24] ),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold652 (.A(\m_sys.m_ram.m_ram.r_mem[9][21] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold653 (.A(\m_sys.m_ram.m_ram.r_mem[5][24] ),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold654 (.A(\m_sys.m_core.m_gpr._GEN[41] ),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold655 (.A(\m_sys.m_ram.m_ram.r_mem[10][25] ),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold656 (.A(\m_sys.m_core.m_gpr._GEN[81] ),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold657 (.A(\m_sys.m_ram.m_ram.r_mem[3][24] ),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold658 (.A(\m_sys.m_ram.m_ram.r_mem[26][24] ),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold659 (.A(\m_sys.m_core.m_gpr._GEN[84] ),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold660 (.A(\m_sys.m_ram.m_ram.r_mem[4][17] ),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold661 (.A(\m_sys.m_ram.m_ram.r_mem[29][21] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold662 (.A(\m_sys.m_ram.m_ram.r_mem[31][31] ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold663 (.A(\m_sys.m_ram.m_ram.r_mem[17][21] ),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold664 (.A(\m_sys.m_ram.m_ram.r_mem[1][27] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold665 (.A(\m_sys.m_ram.m_ram.r_mem[31][30] ),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold666 (.A(\m_sys.m_ram.m_ram.r_mem[23][27] ),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold667 (.A(\m_sys.m_ram.m_ram.r_mem[31][18] ),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold668 (.A(\m_sys.m_core.m_gpr._GEN[202] ),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold669 (.A(_01642_),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold670 (.A(\m_sys.m_ram.m_ram.r_mem[25][22] ),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold671 (.A(\m_sys.m_ram.m_ram.r_mem[7][12] ),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold672 (.A(\m_sys.m_ram.m_ram.r_mem[10][21] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold673 (.A(\m_sys.m_ram.m_ram.r_mem[12][18] ),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold674 (.A(\m_sys.m_ram.m_ram.r_mem[18][23] ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold675 (.A(\m_sys.m_ram.m_ram.r_mem[25][18] ),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold676 (.A(\m_sys.m_core.m_gpr._GEN[78] ),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold677 (.A(\m_sys.m_ram.m_ram.r_mem[25][20] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold678 (.A(\m_sys.m_core.m_gpr._GEN[74] ),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold679 (.A(_01545_),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold680 (.A(\m_sys.m_ram.m_ram.r_mem[12][26] ),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold681 (.A(\m_sys.m_ram.m_ram.r_mem[9][26] ),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold682 (.A(\m_sys.m_ram.m_ram.r_mem[12][16] ),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold683 (.A(\m_sys.m_ram.m_ram.r_mem[1][21] ),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold684 (.A(\m_sys.m_ram.m_ram.r_mem[24][26] ),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold685 (.A(\m_sys.m_ram.m_ram.r_mem[2][26] ),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold686 (.A(\m_sys.m_ram.m_ram.r_mem[16][31] ),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold687 (.A(\m_sys.m_ram.m_ram.r_mem[2][30] ),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold688 (.A(\m_sys.m_ram.m_ram.r_mem[14][23] ),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold689 (.A(\m_sys.m_ram.m_ram.r_mem[20][27] ),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold690 (.A(\m_sys.m_ram.m_ram.r_mem[8][20] ),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold691 (.A(\m_sys.m_ram.m_ram.r_mem[31][28] ),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold692 (.A(\m_sys.m_ram.m_ram.r_mem[10][19] ),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold693 (.A(\m_sys.m_ram.m_ram.r_mem[13][18] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold694 (.A(\m_sys.m_ram.m_ram.r_mem[18][31] ),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold695 (.A(\m_sys.m_core.m_gpr._GEN[50] ),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold696 (.A(\m_sys.m_ram.m_ram.r_mem[13][23] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold697 (.A(\m_sys.m_core.m_gpr._GEN[76] ),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold698 (.A(\m_sys.m_ram.m_ram.r_mem[18][19] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold699 (.A(\m_sys.m_core.m_gpr._GEN[51] ),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold700 (.A(\m_sys.m_ram.m_ram.r_mem[23][5] ),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold701 (.A(\m_sys.m_ram.m_ram.r_mem[16][23] ),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold702 (.A(\m_sys.m_ram.m_ram.r_mem[8][16] ),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold703 (.A(\m_sys.m_ram.m_ram.r_mem[27][31] ),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold704 (.A(\m_sys.m_ram.m_ram.r_mem[13][0] ),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold705 (.A(\m_sys.m_ram.m_ram.r_mem[0][30] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold706 (.A(\m_sys.m_core.m_gpr._GEN[70] ),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold707 (.A(\m_sys.m_ram.m_ram.r_mem[22][21] ),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold708 (.A(\m_sys.m_ram.m_ram.r_mem[8][23] ),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold709 (.A(\m_sys.m_ram.m_ram.r_mem[21][20] ),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold710 (.A(\m_sys.m_ram.m_ram.r_mem[24][19] ),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold711 (.A(\m_sys.m_ram.m_ram.r_mem[22][6] ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold712 (.A(\m_sys.m_ram.m_ram.r_mem[11][31] ),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold713 (.A(\m_sys.m_ram.m_ram.r_mem[7][26] ),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold714 (.A(\m_sys.m_ram.m_ram.r_mem[8][21] ),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold715 (.A(\m_sys.m_ram.m_ram.r_mem[11][16] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold716 (.A(\m_sys.m_ram.m_ram.r_mem[13][17] ),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold717 (.A(\m_sys.m_ram.m_ram.r_mem[18][20] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold718 (.A(\m_sys.m_ram.m_ram.r_mem[25][17] ),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold719 (.A(\m_sys.m_ram.m_ram.r_mem[8][18] ),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold720 (.A(\m_sys.m_ram.m_ram.r_mem[8][19] ),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold721 (.A(\m_sys.m_ram.m_ram.r_mem[13][31] ),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold722 (.A(\m_sys.m_ram.m_ram.r_mem[5][20] ),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold723 (.A(\m_sys.m_ram.m_ram.r_mem[11][20] ),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold724 (.A(\m_sys.m_ram.m_ram.r_mem[3][25] ),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold725 (.A(\m_sys.m_uart.r_rx_data[2] ),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold726 (.A(_07413_),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold727 (.A(\m_sys.m_ram.m_ram.r_mem[27][29] ),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold728 (.A(\m_sys.m_ram.m_ram.r_mem[28][17] ),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold729 (.A(\m_sys.m_ram.m_ram.r_mem[25][23] ),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold730 (.A(\m_sys.m_core.m_gpr._GEN[88] ),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold731 (.A(\m_sys.m_core.m_gpr._GEN[95] ),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold732 (.A(_01566_),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold733 (.A(\m_sys.m_ram.m_ram.r_mem[13][26] ),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold734 (.A(\m_sys.m_ram.m_ram.r_mem[14][25] ),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold735 (.A(\m_sys.m_ram.m_ram.r_mem[14][19] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold736 (.A(\m_sys.m_ram.m_ram.r_mem[19][30] ),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold737 (.A(\m_sys.m_ram.m_ram.r_mem[17][25] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold738 (.A(\m_sys.m_ram.m_ram.r_mem[26][19] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold739 (.A(\m_sys.m_ram.m_ram.r_mem[13][25] ),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold740 (.A(\m_sys.m_ram.m_ram.r_mem[3][26] ),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold741 (.A(\m_sys.m_core.m_gpr._GEN[183] ),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold742 (.A(\m_sys.m_ram.m_ram.r_mem[23][18] ),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold743 (.A(\m_sys.m_ram.m_ram.r_mem[5][29] ),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold744 (.A(\m_sys.m_ram.m_ram.r_mem[28][24] ),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold745 (.A(\m_sys.m_ram.m_ram.r_mem[5][28] ),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold746 (.A(\m_sys.m_ram.m_ram.r_mem[24][29] ),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold747 (.A(\m_sys.m_ram.m_ram.r_mem[12][0] ),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold748 (.A(\m_sys.m_core.m_gpr._GEN[44] ),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold749 (.A(\m_sys.m_ram.m_ram.r_mem[12][22] ),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold750 (.A(\m_sys.m_ram.m_ram.r_mem[20][16] ),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold751 (.A(\m_sys.m_ram.m_ram.r_mem[16][20] ),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold752 (.A(\m_sys.m_ram.m_ram.r_mem[10][20] ),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold753 (.A(\m_sys.m_ram.m_ram.r_mem[27][23] ),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold754 (.A(\m_sys.m_ram.m_ram.r_mem[26][27] ),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold755 (.A(\m_sys.m_ram.m_ram.r_mem[17][28] ),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold756 (.A(\m_sys.m_ram.m_ram.r_mem[30][21] ),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold757 (.A(\m_sys.m_ram.m_ram.r_mem[22][1] ),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold758 (.A(\m_sys.m_ram.m_ram.r_mem[5][25] ),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold759 (.A(\m_sys.m_core.m_gpr._GEN[204] ),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold760 (.A(\m_sys.m_ram.m_ram.r_mem[3][21] ),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold761 (.A(\m_sys.m_ram.m_ram.r_mem[22][19] ),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold762 (.A(\m_sys.m_ram.m_ram.r_mem[7][28] ),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold763 (.A(\m_sys.m_core.m_gpr._GEN[55] ),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold764 (.A(\m_sys.m_ram.m_ram.r_mem[15][26] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold765 (.A(\m_sys.m_ram.m_ram.r_mem[28][23] ),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold766 (.A(\m_sys.m_ram.m_ram.r_mem[29][30] ),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold767 (.A(\m_sys.m_ram.m_ram.r_mem[6][22] ),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold768 (.A(\m_sys.m_core.m_gpr._GEN[77] ),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold769 (.A(\m_sys.m_ram.m_ram.r_mem[21][23] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold770 (.A(\m_sys.m_ram.m_ram.r_mem[27][26] ),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold771 (.A(\m_sys.m_ram.m_ram.r_mem[12][19] ),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold772 (.A(\m_sys.m_core.m_gpr._GEN[34] ),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold773 (.A(\m_sys.m_ram.m_ram.r_mem[21][16] ),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold774 (.A(\m_sys.m_ram.m_ram.r_mem[28][19] ),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold775 (.A(\m_sys.m_ram.m_ram.r_mem[14][21] ),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold776 (.A(\m_sys.m_core.m_gpr._GEN[182] ),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold777 (.A(\m_sys.m_ram.m_ram.r_mem[10][2] ),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold778 (.A(\m_sys.m_ram.m_ram.r_mem[5][26] ),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold779 (.A(\m_sys.m_ram.m_ram.r_mem[19][26] ),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold780 (.A(\m_sys.m_ram.m_ram.r_mem[14][16] ),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold781 (.A(\m_sys.m_ram.m_ram.r_mem[22][20] ),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold782 (.A(\m_sys.m_ram.m_ram.r_mem[6][24] ),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold783 (.A(\m_sys.m_ram.m_ram.r_mem[16][19] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold784 (.A(\m_sys.m_ram.m_ram.r_mem[4][23] ),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold785 (.A(\m_sys.m_ram.m_ram.r_mem[6][31] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold786 (.A(\m_sys.m_ram.m_ram.r_mem[7][18] ),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold787 (.A(\m_sys.m_ram.m_ram.r_mem[25][25] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold788 (.A(\m_sys.m_core.m_gpr._GEN[59] ),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold789 (.A(\m_sys.m_ram.m_ram.r_mem[26][30] ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold790 (.A(\m_sys.m_ram.m_ram.r_mem[3][30] ),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold791 (.A(\m_sys.m_ram.m_ram.r_mem[5][16] ),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold792 (.A(\m_sys.m_uart.r_rx_data[4] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold793 (.A(_01178_),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold794 (.A(\m_sys.m_core.m_gpr._GEN[75] ),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold795 (.A(\m_sys.m_ram.m_ram.r_mem[28][27] ),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold796 (.A(\m_sys.m_core.m_gpr._GEN[102] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold797 (.A(\m_sys.m_ram.m_ram.r_mem[15][29] ),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold798 (.A(\m_sys.m_bootloader.r_byte_cnt[14] ),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold799 (.A(_01326_),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold800 (.A(\m_sys.m_ram.m_ram.r_mem[7][25] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold801 (.A(\m_sys.m_ram.m_ram.r_mem[16][27] ),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold802 (.A(\m_sys.m_ram.m_ram.r_mem[26][17] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold803 (.A(\m_sys.m_core.m_gpr._GEN[61] ),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold804 (.A(\m_sys.m_ram.m_ram.r_mem[25][16] ),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold805 (.A(\m_sys._GEN_11[3] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold806 (.A(_00155_),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold807 (.A(\m_sys.m_core.m_gpr._GEN[54] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold808 (.A(\m_sys.m_ram.m_ram.r_mem[9][27] ),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold809 (.A(\m_sys.m_ram.m_ram.r_mem[3][22] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold810 (.A(\m_sys.m_ram.m_ram.r_mem[14][28] ),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold811 (.A(\m_sys.m_ram.m_ram.r_mem[19][24] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold812 (.A(\m_sys.m_ram.m_ram.r_mem[28][29] ),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold813 (.A(\m_sys.m_core.m_gpr._GEN[57] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold814 (.A(\m_sys.m_ram.m_ram.r_mem[26][28] ),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold815 (.A(\m_sys.m_ram.m_ram.r_mem[23][17] ),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold816 (.A(\m_sys.m_ram.m_ram.r_mem[25][5] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold817 (.A(\m_sys.m_ram.m_ram.r_mem[1][26] ),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold818 (.A(_00076_),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold819 (.A(_00173_),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold820 (.A(\m_sys.m_core.m_gpr._GEN[190] ),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold821 (.A(_01630_),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold822 (.A(\m_sys.m_core.m_gpr._GEN[56] ),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold823 (.A(\m_sys.m_ram.m_ram.r_mem[10][18] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold824 (.A(\m_sys.m_ram.m_ram.r_mem[9][30] ),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold825 (.A(\m_sys.m_ram.m_ram.r_mem[9][18] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold826 (.A(\m_sys.m_ram.m_ram.r_mem[29][17] ),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold827 (.A(\m_sys.m_ram.m_ram.r_mem[17][22] ),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold828 (.A(\m_sys.m_ram.m_ram.r_mem[11][23] ),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold829 (.A(\m_sys.m_ram.m_ram.r_mem[6][18] ),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold830 (.A(\m_sys.m_ram.m_ram.r_mem[19][25] ),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold831 (.A(\m_sys.m_core.m_gpr._GEN[86] ),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold832 (.A(\m_sys.m_ram.m_ram.r_mem[11][19] ),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold833 (.A(\m_sys.m_core.m_gpr._GEN[42] ),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold834 (.A(_01577_),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold835 (.A(\m_sys.m_ram.m_ram.r_mem[18][21] ),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold836 (.A(\m_sys.m_ram.m_ram.r_mem[25][31] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold837 (.A(\m_sys.m_ram.m_ram.r_mem[31][24] ),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold838 (.A(\m_sys.m_ram.m_ram.r_mem[3][20] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold839 (.A(\m_sys.m_ram.m_ram.r_mem[27][30] ),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold840 (.A(\m_sys.m_ram.m_ram.r_mem[5][30] ),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold841 (.A(\m_sys.m_ram.m_ram.r_mem[19][20] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold842 (.A(\m_sys.m_ram.m_ram.r_mem[2][22] ),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold843 (.A(\m_sys.m_ram.m_ram.r_mem[3][23] ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold844 (.A(\m_sys.m_ram.m_ram.r_mem[30][29] ),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold845 (.A(\m_sys.m_ram.m_ram.r_mem[22][7] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold846 (.A(\m_sys.m_ram.m_ram.r_mem[20][25] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold847 (.A(\m_sys.m_ram.m_ram.r_mem[5][22] ),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold848 (.A(\m_sys.m_ram.m_ram.r_mem[10][31] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold849 (.A(\m_sys.m_ram.m_ram.r_mem[4][16] ),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold850 (.A(\m_sys.m_core.m_gpr._GEN[167] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold851 (.A(\m_sys.m_ram.m_ram.r_mem[19][31] ),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold852 (.A(\m_sys.m_ram.m_ram.r_mem[16][16] ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold853 (.A(\m_sys.m_ram.m_ram.r_mem[17][20] ),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold854 (.A(\m_sys.m_core.m_gpr._GEN[189] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold855 (.A(\m_sys.m_ram.m_ram.r_mem[28][26] ),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold856 (.A(\m_sys.m_ram.m_ram.r_mem[9][17] ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold857 (.A(\m_sys.m_core.m_gpr._GEN[68] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold858 (.A(\m_sys.m_core.m_gpr._GEN[65] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold859 (.A(\m_sys.m_ram.m_ram.r_mem[20][22] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold860 (.A(\m_sys.m_ram.m_ram.r_mem[16][29] ),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold861 (.A(\m_sys.m_core.m_gpr._GEN[45] ),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold862 (.A(\m_sys.m_ram.m_ram.r_mem[8][30] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold863 (.A(\m_sys.m_ram.m_ram.r_mem[30][17] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold864 (.A(\m_sys.m_ram.m_ram.r_mem[18][16] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold865 (.A(\m_sys.m_ram.m_ram.r_mem[18][29] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold866 (.A(\m_sys.m_ram.m_ram.r_mem[15][18] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold867 (.A(\m_sys.m_core.m_gpr._GEN[205] ),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold868 (.A(\m_sys.m_ram.m_ram.r_mem[4][20] ),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold869 (.A(\m_sys._m_uart_io_o_bl_data[1] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold870 (.A(\m_sys.m_ram.m_ram.r_mem[15][28] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold871 (.A(\m_sys.m_core.m_gpr._GEN[203] ),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold872 (.A(\m_sys.m_ram.m_ram.r_mem[4][18] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold873 (.A(\m_sys.m_ram.m_ram.r_mem[2][17] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold874 (.A(\m_sys.m_ram.m_ram.r_mem[31][29] ),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold875 (.A(\m_sys.m_ram.m_ram.r_mem[14][27] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold876 (.A(\m_sys.m_ram.m_ram.r_mem[9][31] ),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold877 (.A(\m_sys.m_ram.m_ram.r_mem[25][19] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold878 (.A(\m_sys.m_ram.m_ram.r_mem[22][18] ),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold879 (.A(\m_sys.m_ram.m_ram.r_mem[11][22] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold880 (.A(\m_sys.m_uart.r_rx_valid ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold881 (.A(_01196_),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold882 (.A(\m_sys.m_ram.m_ram.r_mem[21][30] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold883 (.A(\m_sys.m_core.m_gpr._GEN[38] ),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold884 (.A(\m_sys.m_core.m_gpr._GEN[89] ),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold885 (.A(\m_sys.m_ram.m_ram.r_mem[4][27] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold886 (.A(\m_sys.m_ram.m_ram.r_mem[17][17] ),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold887 (.A(\m_sys.m_ram.m_ram.r_mem[14][29] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold888 (.A(\m_sys.m_core.m_gpr._GEN[217] ),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold889 (.A(\m_sys.m_core.m_gpr._GEN[73] ),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold890 (.A(\m_sys.m_ram.m_ram.r_mem[0][23] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold891 (.A(\m_sys.m_ram.m_ram.r_mem[15][24] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold892 (.A(\m_sys.m_ram.m_ram.r_mem[21][24] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold893 (.A(\m_sys.m_ram.m_ram.r_mem[17][19] ),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold894 (.A(\m_sys.m_ram.m_ram.r_mem[26][29] ),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold895 (.A(\m_sys.m_ram.m_ram.r_mem[28][21] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold896 (.A(\m_sys.m_ram.m_ram.r_mem[9][16] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold897 (.A(\m_sys.m_ram.m_ram.r_mem[15][21] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold898 (.A(\m_sys.m_core.m_gpr._GEN[169] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold899 (.A(\m_sys.m_core.m_gpr._GEN[219] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold900 (.A(\m_sys.m_ram.m_ram.r_mem[31][16] ),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold901 (.A(\m_sys.m_ram.m_ram.r_mem[8][27] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold902 (.A(\m_sys.m_ram.m_ram.r_mem[12][7] ),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold903 (.A(\m_sys.m_uart.m_tx.r_data[1] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold904 (.A(_00988_),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold905 (.A(\m_sys.m_ram.m_ram.r_mem[4][26] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold906 (.A(\m_sys.m_ram.m_ram.r_mem[0][18] ),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold907 (.A(\m_sys.m_ram.m_ram.r_mem[22][26] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold908 (.A(\m_sys.m_bootloader.r_byte_cnt[15] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold909 (.A(_01327_),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold910 (.A(\m_sys.m_core.m_gpr._GEN[208] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold911 (.A(\m_sys.m_ram.m_ram.r_mem[17][27] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold912 (.A(\m_sys.m_ram.m_ram.r_mem[31][27] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold913 (.A(\m_sys.m_ram.m_ram.r_mem[11][17] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold914 (.A(\m_sys.m_uart.m_tx.r_data[0] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold915 (.A(\m_sys.m_ram.m_ram.r_mem[19][23] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold916 (.A(\m_sys.m_ram.m_ram.r_mem[20][31] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold917 (.A(\m_sys.m_ram.m_ram.r_mem[27][27] ),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold918 (.A(\m_sys.m_ram.m_ram.r_mem[31][17] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold919 (.A(\m_sys.m_ram.m_ram.r_mem[24][24] ),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold920 (.A(\m_sys.m_core.m_gpr._GEN[52] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold921 (.A(\m_sys.m_ram.m_ram.r_mem[10][17] ),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold922 (.A(\m_sys.m_core.m_gpr._GEN[191] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold923 (.A(_01631_),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold924 (.A(\m_sys.m_ram.m_ram.r_mem[7][17] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold925 (.A(\m_sys.m_bootloader._GEN_22[9] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold926 (.A(\m_sys.m_ram.m_ram.r_mem[10][23] ),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold927 (.A(\m_sys.m_ram.m_ram.r_mem[28][22] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold928 (.A(\m_sys.m_ram.m_ram.r_mem[2][19] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold929 (.A(\m_sys.m_ram.m_ram.r_mem[24][27] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold930 (.A(\m_sys.m_ram.m_ram.r_mem[1][31] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold931 (.A(\m_sys.m_ram.m_ram.r_mem[4][24] ),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold932 (.A(\m_sys.m_core.m_gpr._GEN[175] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold933 (.A(\m_sys.m_ram.m_ram.r_mem[16][30] ),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold934 (.A(\m_sys.m_ram.m_ram.r_mem[11][25] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold935 (.A(\m_sys.m_core.m_gpr._GEN[174] ),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold936 (.A(\m_sys.m_ram.m_ram.r_mem[3][3] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold937 (.A(\m_sys.m_uart.m_tx.r_data[7] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold938 (.A(\m_sys.m_ram.m_ram.r_mem[4][28] ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold939 (.A(\m_sys.m_ram.m_ram.r_mem[15][25] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold940 (.A(\m_sys.m_ram.m_ram.r_mem[17][18] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold941 (.A(\m_sys.m_ram.m_ram.r_mem[6][23] ),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold942 (.A(\m_sys.m_ram.m_ram.r_mem[29][29] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold943 (.A(\m_sys.m_ram.m_ram.r_mem[1][24] ),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold944 (.A(\m_sys.m_ram.m_ram.r_mem[1][22] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold945 (.A(\m_sys.m_core.m_gpr._GEN[58] ),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold946 (.A(\m_sys.m_ram.m_ram.r_mem[9][20] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold947 (.A(\m_sys.m_ram.m_ram.r_mem[10][27] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold948 (.A(\m_sys.m_ram.m_ram.r_mem[31][21] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold949 (.A(\m_sys.m_ram.m_ram.r_mem[0][17] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold950 (.A(\m_sys.m_ram.m_ram.r_mem[0][22] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold951 (.A(\m_sys.m_ram.m_ram.r_mem[23][29] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold952 (.A(\m_sys.m_ram.m_ram.r_mem[8][17] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold953 (.A(\m_sys.m_ram.m_ram.r_mem[30][26] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold954 (.A(\m_sys.m_ram.m_ram.r_mem[20][30] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold955 (.A(\m_sys.m_ram.m_ram.r_mem[29][20] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold956 (.A(\m_sys.m_ram.m_ram.r_mem[11][27] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold957 (.A(\m_sys.m_ram.m_ram.r_mem[6][26] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold958 (.A(\m_sys.m_ram.m_ram.r_mem[7][23] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold959 (.A(\m_sys.m_core.m_gpr._GEN[87] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold960 (.A(\m_sys.m_bootloader._GEN_22[10] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold961 (.A(_01066_),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold962 (.A(\m_sys.m_ram.m_ram.r_mem[31][22] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold963 (.A(\m_sys.m_ram.m_ram.r_mem[30][27] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold964 (.A(\m_sys.m_ram.m_ram.r_mem[18][22] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold965 (.A(\m_sys.m_ram.m_ram.r_mem[0][26] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold966 (.A(\m_sys.m_ram.m_ram.r_mem[10][29] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold967 (.A(\m_sys.m_ram.m_ram.r_mem[23][25] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold968 (.A(\m_sys.m_ram.m_ram.r_mem[20][19] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold969 (.A(\m_sys.m_ram.m_ram.r_mem[21][17] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold970 (.A(\m_sys.m_ram.m_ram.r_mem[18][18] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold971 (.A(\m_sys.m_ram.m_ram.r_mem[17][30] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold972 (.A(\m_sys.m_ram.m_ram.r_mem[13][22] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold973 (.A(\m_sys.m_ram.m_ram.r_mem[9][23] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold974 (.A(\m_sys.m_ram.m_ram.r_mem[13][29] ),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold975 (.A(\m_sys.m_ram.m_ram.r_mem[22][23] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold976 (.A(\m_sys.m_ram.m_ram.r_mem[7][24] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold977 (.A(\m_sys.m_core.m_gpr._GEN[53] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold978 (.A(\m_sys.m_core.m_gpr._GEN[184] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold979 (.A(\m_sys.m_ram.m_ram.r_mem[29][19] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold980 (.A(\m_sys.m_core.m_gpr._GEN[185] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold981 (.A(\m_sys.m_ram.m_ram.r_mem[23][16] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold982 (.A(\m_sys.m_core.m_gpr._GEN[172] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold983 (.A(\m_sys.m_ram.m_ram.r_mem[22][24] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold984 (.A(\m_sys.m_ram.m_ram.r_mem[21][19] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold985 (.A(\m_sys.m_ram.m_ram.r_mem[0][31] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold986 (.A(\m_sys.m_ram.m_ram.r_mem[12][17] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold987 (.A(\m_sys.m_ram.m_ram.r_mem[28][31] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold988 (.A(\m_sys.m_ram.m_ram.r_mem[26][22] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold989 (.A(\m_sys.m_ram.m_ram.r_mem[1][28] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold990 (.A(\m_sys.m_ram.m_ram.r_mem[16][28] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold991 (.A(\m_sys.m_ram.m_ram.r_mem[2][18] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold992 (.A(\m_sys.m_ram.m_ram.r_mem[27][20] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold993 (.A(\m_sys.m_core.m_gpr._GEN[166] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold994 (.A(\m_sys.m_ram.m_ram.r_mem[26][20] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold995 (.A(\m_sys.m_core.m_gpr._GEN[171] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold996 (.A(\m_sys.m_ram.m_ram.r_mem[1][23] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold997 (.A(\m_sys.m_ram.m_ram.r_mem[6][29] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold998 (.A(\m_sys.m_ram.m_ram.r_mem[2][23] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold999 (.A(\m_sys.m_ram.m_ram.r_mem[3][27] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\m_sys.m_core.m_gpr._GEN[186] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\m_sys.m_ram.m_ram.r_mem[23][30] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\m_sys.m_ram.m_ram.r_mem[11][28] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\m_sys.m_ram.m_ram.r_mem[29][31] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\m_sys.m_ram.m_ram.r_mem[11][21] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\m_sys.m_ram.m_ram.r_mem[30][24] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\m_sys.m_ram.m_ram.r_mem[12][21] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\m_sys.m_ram.m_ram.r_mem[24][17] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\m_sys.m_ram.m_ram.r_mem[0][27] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\m_sys.m_ram.m_ram.r_mem[1][18] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\m_sys._m_uart_io_o_bl_data[6] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\m_sys.m_core.m_gpr._GEN[43] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\m_sys.m_ram.m_ram.r_mem[20][18] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\m_sys.m_ram.m_ram.r_mem[6][27] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\m_sys.m_ram.m_ram.r_mem[16][26] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\m_sys.m_ram.m_ram.r_mem[8][28] ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\m_sys.m_ram.m_ram.r_mem[30][23] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\m_sys.m_core.m_gpr._GEN[80] ),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\m_sys.m_ram.m_ram.r_mem[0][28] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\m_sys.m_ram.m_ram.r_mem[2][25] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\m_sys.m_ram.m_ram.r_mem[1][17] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\m_sys.m_ram.m_ram.r_mem[17][23] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\m_sys.m_ram.m_ram.r_mem[3][31] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\m_sys.m_core.m_gpr._GEN[215] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\m_sys.m_ram.m_ram.r_mem[4][19] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\m_sys.m_ram.m_ram.r_mem[13][21] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\m_sys.m_ram.m_ram.r_mem[28][30] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\m_sys.m_ram.m_ram.r_mem[30][19] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\m_sys.m_ram.m_ram.r_mem[29][16] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\m_sys.m_core.m_gpr._GEN[82] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\m_sys.m_ram.m_ram.r_mem[3][18] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\m_sys.m_core.m_gpr._GEN[60] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold1032 (.A(_01595_),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\m_sys.m_ram.m_ram.r_mem[2][27] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\m_sys.m_core.m_gpr._GEN[39] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\m_sys.m_ram.m_ram.r_mem[19][16] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\m_sys.m_ram.m_ram.r_mem[31][19] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\m_sys.m_ram.m_ram.r_mem[16][22] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\m_sys.m_ram.m_ram.r_mem[25][24] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\m_sys.m_ram.m_ram.r_mem[22][17] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\m_sys.m_ram.m_ram.r_mem[20][20] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\m_sys.m_ram.m_ram.r_mem[7][16] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\m_sys.m_ram.m_ram.r_mem[30][20] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\m_sys.m_ram.m_ram.r_mem[27][21] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\m_sys.m_ram.m_ram.r_mem[27][17] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\m_sys.m_ram.m_ram.r_mem[29][25] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\m_sys.m_ram.m_ram.r_mem[8][29] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\m_sys.m_ram.m_ram.r_mem[12][24] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\m_sys.m_core.m_gpr._GEN[173] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\m_sys.m_uart.m_tx.r_data[4] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold1050 (.A(_00991_),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\m_sys.m_ram.m_ram.r_mem[23][23] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\m_sys.m_ram.m_ram.r_mem[27][28] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\m_sys.m_ram.m_ram.r_mem[28][18] ),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\m_sys.m_ram.m_ram.r_mem[27][22] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\m_sys.m_core.m_gpr._GEN[79] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\m_sys.m_ram.m_ram.r_mem[10][26] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\m_sys.m_ram.m_ram.r_mem[24][18] ),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\m_sys.m_ram.m_ram.r_mem[27][19] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\m_sys.m_ram.m_ram.r_mem[15][23] ),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\m_sys.m_ram.m_ram.r_mem[26][31] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\m_sys.m_ram.m_ram.r_mem[31][26] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\m_sys.m_uart.m_tx.r_data[5] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\m_sys.m_ram.m_ram.r_mem[27][16] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\m_sys.m_ram.m_ram.r_mem[18][17] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\m_sys.m_ram.m_ram.r_mem[29][26] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\m_sys.m_ram.m_ram.r_mem[12][31] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\m_sys.m_ram.m_ram.r_mem[22][16] ),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\m_sys.m_core.m_gpr._GEN[223] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold1069 (.A(_01663_),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\m_sys.m_ram.m_ram.r_mem[14][22] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\m_sys.m_ram.m_ram.r_mem[27][18] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\m_sys.m_core.m_gpr._GEN[170] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold1073 (.A(_01610_),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\m_sys.m_ram.m_ram.r_mem[4][22] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\m_sys.m_ram.m_ram.r_mem[7][21] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\m_sys.m_ram.m_ram.r_mem[20][23] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\m_sys.m_ram.m_ram.r_mem[1][16] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\m_sys.m_ram.m_ram.r_mem[10][22] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\m_sys.m_ram.m_ram.r_mem[9][22] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\m_sys.m_ram.m_ram.r_mem[6][20] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\m_sys.m_ram.m_ram.r_mem[31][25] ),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\m_sys.m_ram.m_ram.r_mem[6][19] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\m_sys.m_ram.m_ram.r_mem[2][31] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\m_sys.m_uart.m_tx.r_data[3] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\m_sys.m_ram.m_ram.r_mem[12][29] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\m_sys.m_ram.m_ram.r_mem[26][16] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\m_sys.m_core.m_gpr._GEN[194] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\m_sys.m_ram.m_ram.r_mem[15][27] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\m_sys.m_ram.m_ram.r_mem[11][24] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\m_sys.m_ram.m_ram.r_mem[14][30] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\m_sys.m_ram.m_ram.r_mem[19][22] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\m_sys.m_ram.m_ram.r_mem[24][16] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\m_sys.m_ram.m_ram.r_mem[23][21] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\m_sys.m_ram.m_ram.r_mem[12][25] ),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\m_sys.m_core.m_gpr._GEN[66] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\m_sys.m_core.m_gpr._GEN[222] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold1097 (.A(_01662_),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\m_sys.m_ram.m_ram.r_mem[19][17] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\m_sys._m_uart_io_o_bl_data[2] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\m_sys.m_ram.m_ram.r_mem[3][29] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\m_sys.m_ram.m_ram.r_mem[17][26] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\m_sys.m_ram.m_ram.r_mem[19][28] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\m_sys.m_ram.m_ram.r_mem[11][26] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\m_sys.m_ram.m_ram.r_mem[4][25] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\m_sys.m_ram.m_ram.r_mem[13][19] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\m_sys._m_uart_io_o_bl_data[5] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\m_sys.m_ram.m_ram.r_mem[16][25] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\m_sys.m_ram.m_ram.r_mem[24][28] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\m_sys.m_ram.m_ram.r_mem[8][25] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\m_sys.m_ram.m_ram.r_mem[28][16] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\m_sys.m_ram.m_ram.r_mem[29][22] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\m_sys.m_ram.m_ram.r_mem[30][25] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\m_sys.m_ram.m_ram.r_mem[1][25] ),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\m_sys.m_ram.m_ram.r_mem[31][20] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\m_sys.m_core.m_gpr._GEN[160] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold1116 (.A(_01600_),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\m_sys.m_ram.m_ram.r_mem[20][21] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\m_sys.m_core.m_gpr._GEN[206] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\m_sys.m_ram.m_ram.r_mem[30][30] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\m_sys.m_ram.m_ram.r_mem[19][18] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\m_sys.m_core.m_gpr._GEN[179] ),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\m_sys.m_ram.m_ram.r_mem[15][16] ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\m_sys.m_ram.m_ram.r_mem[31][23] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\m_sys.m_ram.m_ram.r_mem[7][27] ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\m_sys.m_ram.m_ram.r_mem[20][17] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\m_sys.m_ram.m_ram.r_mem[22][29] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\m_sys.m_ram.m_ram.r_mem[26][21] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\m_sys.m_ram.m_ram.r_mem[14][24] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\m_sys.m_ram.m_ram.r_mem[22][28] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\m_sys.m_ram.m_ram.r_mem[18][25] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\m_sys.m_core.m_gpr._GEN[162] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\m_sys.m_ram.m_ram.r_mem[17][31] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\m_sys.m_core.m_gpr._GEN[63] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold1134 (.A(_01598_),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\m_sys.m_ram.m_ram.r_mem[16][18] ),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\m_sys.m_ram.m_ram.r_mem[11][29] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\m_sys.m_ram.m_ram.r_mem[22][30] ),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\m_sys.m_ram.m_ram.r_mem[8][24] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\m_sys.m_core.m_gpr._GEN[48] ),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\m_sys.m_ram.m_ram.r_mem[25][30] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\m_sys.m_ram.m_ram.r_mem[23][22] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\m_sys.m_core.m_gpr._GEN[198] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold1143 (.A(_01638_),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\m_sys.m_ram.m_ram.r_mem[23][20] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\m_sys.m_ram.m_ram.r_mem[23][31] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\m_sys.m_bootloader.r_num[4] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold1147 (.A(_01052_),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\m_sys.m_core.m_gpr._GEN[49] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\m_sys.m_core.m_gpr._GEN[197] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\m_sys.m_ram.m_ram.r_mem[19][19] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\m_sys.m_ram.m_ram.r_mem[30][31] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\m_sys.m_ram.m_ram.r_mem[7][19] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\m_sys.m_ram.m_ram.r_mem[3][19] ),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\m_sys.m_core.m_gpr._GEN[46] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\m_sys.m_core.m_gpr._GEN[231] ),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold1156 (.A(_01247_),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\m_sys.m_ram.m_ram.r_mem[24][25] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\m_sys._m_uart_io_o_bl_data[7] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\m_sys.m_ram.m_ram.r_mem[27][24] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\m_sys.m_ram.m_ram.r_mem[24][31] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\m_sys.m_ram.m_ram.r_mem[4][21] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\m_sys.m_ram.m_ram.r_mem[16][17] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\m_sys.m_ram.m_ram.r_mem[16][24] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\m_sys.m_ram.m_ram.r_mem[11][30] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\m_sys.m_ram.m_ram.r_mem[19][27] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\m_sys.m_ram.m_ram.r_mem[14][18] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\m_sys.m_ram.m_ram.r_mem[22][27] ),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\m_sys.m_ram.m_ram.r_mem[15][20] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\m_sys.m_core.m_gpr._GEN[177] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\m_sys.m_core.m_gpr._GEN[252] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold1171 (.A(_01268_),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\m_sys.m_core.m_gpr._GEN[91] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold1173 (.A(_01562_),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\m_sys.m_core.m_gpr._GEN[214] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\m_sys.m_uart.m_rx.r_bit_cnt[2] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold1176 (.A(_01165_),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\m_sys.m_core.m_gpr._GEN[47] ),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\m_sys.m_ram.m_ram.r_mem[26][25] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\m_sys.m_ram.m_ram.r_mem[18][30] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\m_sys.m_bootloader.r_byte_cnt[13] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold1181 (.A(_01325_),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\m_sys.m_core.m_gpr._GEN[236] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold1183 (.A(_01252_),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\m_sys.m_core.m_gpr._GEN[62] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold1185 (.A(_01597_),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\m_sys.m_ram.m_ram.r_mem[23][28] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\m_sys.m_ram.m_ram.r_mem[0][25] ),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\m_sys.m_ram.m_ram.r_mem[14][20] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\m_sys.m_ram.m_ram.r_mem[2][16] ),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\m_sys.m_core.m_gpr._GEN[207] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\m_sys.m_core.m_gpr._GEN[213] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold1192 (.A(_01653_),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\m_sys._m_uart_io_o_bl_data[3] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\m_sys.m_core.m_gpr._GEN[239] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold1195 (.A(_01255_),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\m_sys.m_ram.m_ram.r_mem[10][24] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\m_sys.m_core.m_gpr._GEN[180] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\m_sys.m_ram.m_ram.r_mem[3][28] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\m_sys.m_ram.m_ram.r_mem[15][30] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\m_sys.m_ram.m_ram.r_mem[4][30] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\m_sys.m_bootloader.r_num[3] ),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\m_sys.m_ram.m_ram.r_mem[8][31] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\m_sys.m_ram.m_ram.r_mem[14][26] ),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\m_sys.m_ram.m_ram.r_mem[24][23] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\m_sys.m_ram.m_ram.r_mem[7][30] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\m_sys.m_core.m_gpr._GEN[158] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold1207 (.A(_01501_),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\m_sys.m_ram.m_ram.r_mem[7][31] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\m_sys.m_uart.r_rx_data[0] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold1210 (.A(_01174_),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\m_sys.m_ram.m_ram.r_mem[18][27] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\m_sys.m_ram.m_ram.r_mem[0][29] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\m_sys.m_ram.m_ram.r_mem[15][19] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\m_sys.m_core.m_gpr._GEN[210] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\m_sys.m_core.m_gpr._GEN[199] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold1216 (.A(_01639_),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\m_sys.m_core.m_gpr._GEN[157] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\m_sys.m_core.m_gpr._GEN[188] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold1219 (.A(_01628_),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\m_sys.m_ram.m_ram.r_mem[22][22] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\m_sys.m_ram.m_ram.r_mem[19][21] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\m_sys.m_ram.m_ram.r_mem[18][28] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\m_sys.m_ram.m_ram.r_mem[10][16] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\m_sys.m_bootloader.r_num_cnt[1] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold1225 (.A(_06246_),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold1226 (.A(_01032_),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\m_sys.m_bootloader.r_byte_cnt[6] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\m_sys.m_ram.m_ram.r_mem[12][23] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\m_sys.m_bootloader.r_num[2] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\m_sys.m_core.m_gpr._GEN[140] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\m_sys.m_uart.m_tx.r_cstate[0] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold1232 (.A(_04919_),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\m_sys.m_ram.m_ram.r_mem[15][22] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\m_sys.m_core.m_gpr._GEN[230] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold1235 (.A(_01246_),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\m_sys.m_core.m_gpr._GEN[115] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\m_sys.m_bootloader.r_num[5] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\m_sys.m_bootloader.r_num[6] ),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\m_sys.m_core.m_gpr._GEN[247] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold1240 (.A(_01263_),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\m_sys.m_core.m_gpr._GEN[112] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\m_sys.m_core.m_gpr._GEN[229] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\m_sys.m_bootloader._GEN_22[11] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\m_sys.m_bootloader.r_num[7] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\m_sys.m_core.m_gpr._GEN[141] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\m_sys.m_core.m_gpr._GEN[209] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\m_sys.m_core.m_gpr._GEN[98] ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold1248 (.A(_01505_),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\m_sys.m_core.m_gpr._GEN[246] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\m_sys.m_uart.m_rx.r_cstate[0] ),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold1251 (.A(_01171_),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\m_sys.m_bootloader.r_num[0] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold1253 (.A(_01048_),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\m_sys.m_ram.m_ram.r_mem[23][26] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\m_sys.m_core.m_gpr._GEN[241] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\m_sys.m_ram.m_ram.r_mem[23][24] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\m_sys.m_core.m_gpr._GEN[105] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[2] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold1259 (.A(_02531_),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold1260 (.A(_01768_),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\m_sys.m_core.m_gpr._GEN[149] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\m_sys.m_ram.m_ram.r_mem[0][24] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\m_sys.m_uart.m_tx.r_data[2] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\m_sys.m_bootloader._GEN_22[2] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\m_sys.m_core.m_gpr._GEN[201] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold1266 (.A(_01641_),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\m_sys.m_ram.m_ram.r_mem[2][28] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\m_sys.m_bootloader.r_byte_cnt[12] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold1269 (.A(_01324_),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\m_sys.m_core.m_gpr._GEN[114] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\m_sys.m_core.m_gpr._GEN[111] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\m_sys.m_core.m_gpr._GEN[251] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold1273 (.A(_01267_),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\m_sys.m_bootloader.r_offset_1[7] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\m_sys.m_core.m_gpr._GEN[244] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\m_sys.m_core.m_gpr._GEN[107] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\m_sys.m_core.m_gpr._GEN[152] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\m_sys.m_core.m_gpr.io_b_write_addr[2] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\m_sys.m_bootloader._GEN_22[8] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold1280 (.A(_01064_),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\m_sys.m_core.m_gpr._GEN[253] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold1282 (.A(_01269_),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[12] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold1284 (.A(_02547_),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold1285 (.A(_01763_),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\m_sys.m_core.m_gpr._GEN[255] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold1287 (.A(_01271_),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\m_sys.m_core.m_gpr._GEN[240] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\m_sys.m_core.m_gpr._GEN[155] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\m_sys.m_core.m_gpr._GEN[237] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\m_sys.m_core.m_gpr._GEN[139] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold1292 (.A(_01482_),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\m_sys.m_core.r_ctrl_mem_rw ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\m_sys.m_core.m_gpr._GEN[117] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\m_sys.m_bootloader.r_offset_0[6] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\m_sys.m_core.m_gpr._GEN[156] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold1297 (.A(_01499_),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\m_sys.m_core.m_gpr._GEN[110] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[8] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\m_sys.m_core.m_gpr._GEN[138] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold1301 (.A(_01481_),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\m_sys.m_ram.m_ram.r_mem[20][29] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\m_sys.m_core.m_gpr._GEN[235] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold1304 (.A(_01251_),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\m_sys.m_core.m_gpr._GEN[242] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold1306 (.A(_01258_),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\m_sys.m_core.m_gpr._GEN[146] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold1308 (.A(_01489_),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\m_sys.m_core.m_gpr._GEN[232] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\m_sys.m_core.m_gpr._GEN[119] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\m_sys.m_core.r_ctrl_wb_en ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\m_sys.m_core.m_gpr._GEN[248] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold1313 (.A(_01264_),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\m_sys.m_core.m_gpr._GEN[103] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\m_sys.m_core.m_gpr._GEN[126] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold1316 (.A(_01533_),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\m_sys.m_bootloader.r_num[1] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\m_sys.m_core.m_gpr._GEN[147] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold1319 (.A(_01490_),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\m_sys.m_core.m_gpr._GEN[224] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold1321 (.A(_01240_),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\m_sys.m_core.m_gpr._GEN[245] ),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\m_sys.m_core.m_gpr._GEN[142] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold1324 (.A(_01485_),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\m_sys.m_core.m_gpr._GEN[67] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\m_sys.m_core.m_gpr._GEN[238] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold1327 (.A(_01254_),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\m_sys.m_core.m_gpr._GEN[133] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold1329 (.A(_01476_),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\m_sys.m_core.m_gpr._GEN[249] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold1331 (.A(_01265_),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\m_sys.m_bootloader.r_cstate[4] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\m_sys.m_core.m_gpr._GEN[195] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\m_sys.m_core.m_gpr._GEN[132] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\m_sys.m_core.m_gpr._GEN[129] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold1336 (.A(_01472_),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold1337 (.A(_00083_),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold1338 (.A(_00180_),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\m_sys.m_core.m_gpr._GEN[120] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\m_sys.m_core.m_gpr._GEN[109] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\m_sys.m_core.m_gpr._GEN[127] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold1342 (.A(_01534_),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\m_sys.m_core.m_gpr._GEN[233] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold1344 (.A(_01249_),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\m_sys.m_core.m_gpr._GEN[250] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold1346 (.A(_01266_),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\m_sys.m_core.m_gpr._GEN[118] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\m_sys.m_bootloader.r_byte_cnt[11] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold1349 (.A(_01323_),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\m_sys._m_uart_io_o_bl_data[4] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold1351 (.A(_01170_),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\m_sys.m_core.m_gpr._GEN[150] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\m_sys.m_core.m_gpr._GEN[254] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold1354 (.A(_01270_),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\m_sys.m_core.m_gpr._GEN[136] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\m_sys.m_core.m_gpr._GEN[106] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold1357 (.A(_01513_),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\m_sys.m_core.m_gpr._GEN[96] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold1359 (.A(_01503_),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\m_sys.m_core.m_gpr._GEN[108] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\m_sys.m_core.m_gpr._GEN[153] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold1362 (.A(_01496_),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\m_sys.m_core.m_gpr._GEN[123] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\m_sys.m_core.m_gpr._GEN[125] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\m_sys.m_core.m_gpr._GEN[72] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\m_sys.m_core.m_bru.io_i_s2[10] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\m_sys.m_core.m_gpr._GEN[196] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\m_sys.m_core.m_gpr._GEN[69] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\m_sys.m_bootloader.r_byte_cnt[9] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold1370 (.A(_01321_),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\m_sys.m_core.m_gpr._GEN[101] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold1372 (.A(_01508_),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\m_sys.m_core.m_gpr._GEN[200] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\m_sys.m_core.m_gpr._GEN[193] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\m_sys.m_core.m_bru.io_i_s2[9] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\m_sys.m_core.m_gpr._GEN[124] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold1377 (.A(_01531_),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[10] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold1379 (.A(_02544_),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold1380 (.A(_01761_),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\m_sys.m_core.m_gpr._GEN[159] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold1382 (.A(_01502_),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\m_sys.m_core.m_gpr._GEN[145] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\m_sys._m_bootloader_io_b_mem_addr[6] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold1385 (.A(_01092_),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\m_sys.m_ram.m_ram.r_mem[9][29] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\m_sys.m_core.m_gpr._GEN[121] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\m_sys.m_bootloader._GEN_22[3] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\m_sys.m_core.m_gpr._GEN[104] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\m_sys.m_core.m_bru.io_i_s2[26] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\m_sys.m_core.m_gpr._GEN[116] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\m_sys.m_bootloader._GEN_22[7] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\m_sys.m_bootloader.r_byte_cnt[8] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\m_sys.m_core.m_gpr._GEN[144] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\m_sys.m_core.m_gpr._GEN[134] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\m_sys.m_bootloader._GEN_22[4] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\m_sys.m_core.m_gpr._GEN[130] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold1398 (.A(_01473_),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\m_sys.m_core.m_gpr._GEN[137] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[15] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\m_sys.m_core.m_gpr._GEN[243] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold1402 (.A(_01259_),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\m_sys.m_bootloader._GEN_22[6] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\m_sys.m_core.m_gpr._GEN[122] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\m_sys.m_core.m_gpr._GEN[154] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\m_sys.m_core.m_gpr._GEN[97] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold1407 (.A(_01504_),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\m_sys.m_bootloader.r_byte_cnt[10] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold1409 (.A(_01322_),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\m_sys.m_core.m_gpr._GEN[226] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold1411 (.A(_01242_),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\m_sys.m_core.m_gpr._GEN[100] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\m_sys.m_core.m_bru.io_i_uop[2] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\m_sys.m_bootloader.r_offset_1[0] ),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold1415 (.A(_01076_),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\m_sys.m_core.m_gpr._GEN[131] ),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\m_sys.m_core.m_gpr._GEN[99] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\m_sys.m_core.r_ctrl_mem_signed ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\m_sys.m_bootloader._GEN_22[5] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\m_sys.m_core.m_gpr._GEN[151] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold1421 (.A(_01494_),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\m_sys.m_core.m_gpr._GEN[37] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[10] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\m_sys.m_core.m_gpr._GEN[234] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold1425 (.A(_01250_),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\m_sys.m_bootloader.r_byte_cnt[4] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\m_sys.m_core.r_ctrl_bru_pc_rel ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\m_sys.m_core.m_gpr._GEN[148] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\m_sys.m_core.m_gpr._GEN[135] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\m_sys.m_core.m_bru.io_i_pc[11] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold1431 (.A(_05639_),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\m_sys.m_core.m_bru.io_i_uop[0] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\m_sys.m_core.m_gpr._GEN[40] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\m_sys.m_bootloader.r_offset_1[1] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\m_sys.m_bootloader.r_offset_1[5] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\m_sys.m_core.m_gpr._GEN[163] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[13] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\m_sys.m_bootloader.r_offset_1[6] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\m_sys.m_core.m_gpr._GEN[227] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\m_sys._m_core_io_b_mem_wdata[13] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold1441 (.A(_00177_),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[0] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\m_sys._m_ram_io_b_port_rdata[13] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\m_sys.m_core.m_gpr._GEN[35] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[6] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold1446 (.A(_02537_),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold1447 (.A(_01772_),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\m_sys._m_bootloader_io_b_mem_addr[3] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold1449 (.A(_01089_),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\m_sys.m_core.m_gpr._GEN[113] ),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\m_sys.m_core.m_gpr._GEN[225] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold1452 (.A(_01241_),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\m_sys.m_core.m_gpr._GEN[168] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\m_sys.m_bootloader.r_num_cnt[2] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold1455 (.A(_06248_),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[9] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\m_sys.m_core.m_gpr._GEN[228] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold1458 (.A(_01244_),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\m_sys.m_bootloader.r_byte_cnt[5] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold1460 (.A(_01317_),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\m_sys.r_addr[7] ),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold1462 (.A(_01183_),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\m_sys.m_core.m_gpr._GEN[165] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\m_sys.m_core.m_gpr._GEN[128] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold1465 (.A(_01471_),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\m_sys.m_core.m_gpr._GEN[36] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\m_sys.m_core.m_gpr._GEN[33] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\m_sys.m_bootloader.r_num_cnt[6] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold1469 (.A(_06256_),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\m_sys.m_bootloader.r_num_cnt[5] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold1471 (.A(_06254_),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\m_sys.m_uart.m_rx.r_cstate[1] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold1473 (.A(_04923_),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\m_sys.m_core.m_gpr._GEN[164] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold1475 (.A(_00072_),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold1476 (.A(_00169_),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\m_sys.m_core.m_gpr._GEN[161] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\m_sys.m_core.m_gpr._GEN[192] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold1479 (.A(_01632_),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\m_sys._m_bootloader_io_b_mem_addr[5] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold1481 (.A(_01091_),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\m_sys.m_bootloader.r_byte_cnt[7] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\m_sys._m_ram_io_b_port_rdata[15] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\m_sys.m_bootloader.r_num_cnt[3] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\m_sys.r_addr[6] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold1486 (.A(_01182_),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[9] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold1488 (.A(_02543_),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\m_sys.r_addr[8] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold1490 (.A(_01184_),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\m_sys.m_bootloader.r_offset_0[0] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold1492 (.A(_01068_),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[13] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold1494 (.A(_02549_),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\m_sys.m_uart.m_rx.r_rx ),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[10] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold1497 (.A(_02619_),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\m_sys.m_bootloader.r_offset_0[1] ),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[4] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\m_sys.m_core.m_bru.io_i_s1[10] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\m_sys.m_bootloader.r_offset_1[4] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\m_sys._m_ram_io_b_port_rdata[20] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\m_sys._m_core_io_b_mem_wdata[14] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold1504 (.A(_00178_),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\m_sys._m_ram_io_b_port_rdata[14] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\m_sys._m_ram_io_b_port_rdata[23] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\m_sys.m_bootloader.r_offset_1[3] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\m_sys.m_uart.m_tx.r_bit_cnt[2] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold1509 (.A(_07432_),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[14] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\m_sys.r_addr[9] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold1512 (.A(_01185_),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\m_sys._m_core_io_b_mem_wdata[11] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold1514 (.A(_00175_),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[4] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold1516 (.A(_02534_),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\m_sys.m_bootloader.r_byte_cnt[2] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\m_sys.m_bootloader.r_num_cnt[7] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\m_sys.m_bootloader.r_byte_cnt[3] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\m_sys.m_core._m_bru_io_o_res[1] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold1521 (.A(_01928_),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold1522 (.A(_01362_),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\m_sys.m_core.r_ctrl_mem_size[1] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold1524 (.A(_01367_),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\m_sys.m_core.m_bru.io_i_s2[7] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\m_sys.m_core.m_bru.io_i_uop[1] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold1527 (.A(_00404_),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\m_sys.m_bootloader.r_num_cnt[4] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[2] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold1530 (.A(_02604_),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\m_sys.m_bootloader.r_offset_0[2] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\m_sys.m_core.m_gpr.io_b_write_addr[0] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold1533 (.A(_01371_),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\m_sys.m_core.m_gpr._GEN[143] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\m_sys.m_bootloader.r_offset_0[7] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\m_sys._m_bootloader_io_b_mem_wdata[7] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\m_sys._m_ram_io_b_port_rdata[21] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\m_sys._m_ram_io_b_port_rdata[12] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\m_sys.m_core.m_bru.io_i_s2[28] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[11] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold1541 (.A(_02621_),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\m_sys._m_bootloader_io_b_mem_wen[0] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold1543 (.A(_06358_),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold1544 (.A(\m_sys._m_bootloader_io_b_mem_addr[8] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\m_sys.m_gpio8.r_in[5] ),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold1546 (.A(_02662_),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold1547 (.A(_00005_),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[11] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\m_sys.m_core.m_bru.io_i_s2[1] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold1550 (.A(_01329_),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[3] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold1552 (.A(_02532_),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold1553 (.A(_00014_),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold1554 (.A(_04910_),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\m_sys.m_uart.m_tx.r_bit_cnt[1] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold1556 (.A(_07431_),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold1557 (.A(_00146_),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold1558 (.A(_06245_),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\m_sys.m_bootloader.r_offset_0[3] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[7] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold1561 (.A(_02540_),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\m_sys.m_core.m_bru.io_i_s2[30] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[14] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\m_sys.m_gpio8.r_in[3] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold1565 (.A(_02658_),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold1566 (.A(_00003_),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\m_sys._m_ram_io_b_port_rdata[18] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[8] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\m_sys.m_core._m_bru_io_o_res[0] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold1570 (.A(_01926_),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold1571 (.A(_01361_),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold1572 (.A(uio_out[4]),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\m_sys._m_core_io_b_mem_wdata[15] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\m_sys.m_gpio8.r_in[1] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold1575 (.A(_02654_),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold1576 (.A(_00001_),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[1] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\m_sys.m_core.m_bru.io_i_s2[29] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold1579 (.A(_00073_),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\m_sys.m_core.m_bru.io_i_s2[6] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\m_sys.r_addr[10] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold1582 (.A(_01186_),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[0] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold1584 (.A(_01744_),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\m_sys._m_ram_io_b_port_rdata[11] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\m_sys.m_bootloader.r_offset_0[5] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold1587 (.A(_00085_),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold1588 (.A(_00182_),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\m_sys._m_ram_io_b_port_rdata[8] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\m_sys.m_core.m_bru.io_i_s2[0] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\m_sys._m_bootloader_io_b_mem_wdata[4] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\m_sys._m_bootloader_io_b_mem_addr[11] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold1593 (.A(_01097_),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[11] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\m_sys._m_bootloader_io_b_mem_addr[1] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold1596 (.A(_01087_),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\m_sys.m_core.m_bru.io_i_pc[6] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\m_sys.m_core.m_bru.io_i_s2[5] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_00658_),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\m_sys.m_core.m_bru.io_i_s2[13] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\m_sys.m_gpio8.r_in[2] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold1602 (.A(_02656_),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold1603 (.A(_00002_),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\m_sys.m_core.m_bru.io_i_pc[10] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\m_sys._m_ram_io_b_port_rdata[4] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[6] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold1607 (.A(_02613_),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\m_sys.m_core.m_bru.io_i_s2[11] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\m_sys.m_core.m_bru.io_i_s2[22] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold1610 (.A(_00015_),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold1611 (.A(_02174_),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold1612 (.A(_01599_),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[8] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold1614 (.A(_02617_),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[3] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold1616 (.A(_02607_),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\m_sys._m_ram_io_b_port_rdata[22] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\m_sys._m_ram_io_b_port_rdata[10] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\m_sys._m_bootloader_io_b_mem_wdata[3] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[5] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold1621 (.A(_02611_),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\m_sys.m_core.m_bru.io_i_s2[25] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\m_sys._m_core_io_b_mem_wdata[20] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[7] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[15] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\m_sys.m_core.m_bru.io_i_s2[31] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\m_sys.m_bootloader.r_offset_1[2] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\m_sys.m_gpio8.r_in[6] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold1629 (.A(_02664_),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold1630 (.A(_00006_),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\m_sys.m_gpio8.r_in[4] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold1632 (.A(_00004_),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\m_sys._m_bootloader_io_b_mem_wdata[6] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold1634 (.A(_01046_),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[1] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold1636 (.A(_00079_),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold1637 (.A(_00176_),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold1638 (.A(\m_sys.m_uart.m_rx.r_bit_cnt[1] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold1639 (.A(_04921_),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\m_sys.m_gpio8.r_in[0] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold1641 (.A(_02652_),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold1642 (.A(_00000_),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\m_sys.m_core.m_bru.io_i_s2[8] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold1644 (.A(_00661_),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\m_sys.m_core.m_bru.io_i_s2[4] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold1646 (.A(_00070_),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold1647 (.A(_02804_),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold1648 (.A(_00167_),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\m_sys.m_uart.m_tx.r_bit_cnt[0] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold1650 (.A(_07429_),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\m_sys.m_core.m_bru.io_i_s2[21] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\m_sys._m_ram_io_b_port_rdata[9] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold1653 (.A(uio_out[7]),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\m_sys.m_uart.m_tx.r_cycle_cnt[5] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\m_sys._m_ram_io_b_port_rdata[0] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\m_sys._m_ram_io_b_port_rdata[7] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\m_sys.m_core.m_bru.io_i_s2[23] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\m_sys._m_ram_io_b_port_rdata[19] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\m_sys.m_core.r_ctrl_mem_size[0] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\m_sys.m_core.m_bru.io_i_pc[7] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\m_sys._m_ram_io_b_port_rdata[17] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\m_sys._m_bootloader_io_b_mem_wdata[1] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\m_sys.m_core.m_bru.io_i_s2[18] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[4] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\m_sys._m_ram_io_b_port_rdata[3] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[12] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold1667 (.A(_00066_),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold1668 (.A(_00165_),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\m_sys._m_core_io_b_mem_wdata[21] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\m_sys._m_bootloader_io_b_mem_wdata[5] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\m_sys._m_ram_io_b_port_rdata[2] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\m_sys._m_ram_io_b_port_rdata[6] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\m_sys._m_bootloader_io_b_mem_wdata[0] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold1674 (.A(_01040_),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\m_sys.m_core.m_bru.io_i_s2[17] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\m_sys.m_core.m_gpr.io_b_write_addr[1] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\m_sys._m_core_io_b_mem_wdata[31] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\m_sys._m_core_io_b_mem_wdata[29] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[13] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold1680 (.A(_02626_),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[15] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold1682 (.A(_02630_),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\m_sys._m_ram_io_b_port_rdata[16] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\m_sys.m_core.m_bru.io_i_pc[9] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold1685 (.A(_00662_),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold1686 (.A(\m_sys._m_bootloader_io_b_mem_wdata[2] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold1687 (.A(_01042_),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[12] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\m_sys._m_ram_io_b_port_rdata[1] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\m_sys.m_core.m_bru.io_i_pc[3] ),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold1691 (.A(_05616_),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\m_sys.m_gpio8.r_in[7] ),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold1693 (.A(_00007_),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\m_sys.m_core.m_bru.io_i_s2[15] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\m_sys.m_core.m_bru.io_i_s2[2] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\m_sys.m_core.m_bru.io_i_s2[19] ),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold1697 (.A(_01347_),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\m_sys.r_addr[11] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold1699 (.A(_01187_),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\m_sys.m_uart.m_tx.r_cstate[1] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\m_sys._m_bootloader_io_b_mem_addr[10] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold1702 (.A(_01096_),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[1] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\m_sys.m_uart.m_rx.r_bit_cnt[0] ),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[5] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\m_sys.m_core.m_bru.io_i_s2[20] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold1707 (.A(_00074_),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold1708 (.A(_00171_),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\m_sys._m_ram_io_b_port_rdata[5] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\m_sys.m_core.m_bru.io_i_s1[31] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\m_sys.m_bootloader.r_byte_cnt[0] ),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\m_sys.m_core.m_fsm.r_cstate[1] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\m_sys.m_core.m_bru.io_i_pc[2] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold1714 (.A(_00655_),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[7] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\m_sys.m_bootloader.r_offset_0[4] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\m_sys._m_bootloader_io_b_mem_addr[4] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\m_sys._m_core_io_b_mem_wdata[25] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\m_sys.m_core.m_bru.io_i_s2[27] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold1720 (.A(uio_oe[4]),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold1721 (.A(uio_out[6]),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\m_sys._m_bootloader_io_b_mem_addr[7] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold1723 (.A(_01093_),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold1724 (.A(_00084_),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold1725 (.A(_00181_),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[9] ),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\m_sys.m_uart.m_rx.r_cstate[0] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[6] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\m_sys.m_core.m_bru.io_i_s2[3] ),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold1730 (.A(uio_out[2]),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\m_sys._m_core_io_b_mem_wdata[23] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\m_sys.m_core.m_bru.io_i_pc[4] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold1733 (.A(uio_oe[7]),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\m_sys._m_bootloader_io_b_mem_addr[2] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\m_sys.m_core.m_bru.io_i_s2[12] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\m_sys._m_core_io_b_mem_wdata[27] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold1737 (.A(uio_out[5]),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold1738 (.A(uio_out[3]),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold1739 (.A(_01275_),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\m_sys.m_core.m_bru.io_i_s2[24] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold1741 (.A(_00086_),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold1742 (.A(_00183_),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\m_sys.m_core.m_alu.io_i_uop[1] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold1744 (.A(uio_out[0]),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\m_sys._m_ram_io_b_port_rdata[25] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\m_sys._m_core_io_b_mem_wdata[22] ),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[14] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\m_sys._m_core_io_b_mem_wdata[12] ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\m_sys._m_core_io_b_mem_wdata[4] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold1750 (.A(\m_sys._m_ram_io_b_port_rdata[30] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\m_sys._m_ram_io_b_port_rdata[24] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold1752 (.A(\m_sys.m_core.m_bru.io_i_s2[14] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold1753 (.A(_01342_),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\m_sys._m_core_io_b_mem_wdata[10] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\m_sys.m_uart.m_rx.r_cstate[1] ),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold1756 (.A(uio_out[1]),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\m_sys.m_bootloader.r_cstate[1] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\m_sys._m_core_io_b_mem_wdata[30] ),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\m_sys.m_core.m_bru.io_i_s1[0] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold1760 (.A(_00227_),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[3] ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold1762 (.A(_00011_),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold1763 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[0] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\m_sys.m_bootloader.r_byte_cnt[1] ),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\m_sys.m_core.m_bru.io_i_s2[16] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold1766 (.A(uio_oe[6]),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\m_sys._m_ram_io_b_port_rdata[27] ),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\m_sys._m_bootloader_io_b_mem_addr[9] ),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\m_sys.m_uart.m_rx.io_i_ncycle[2] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold1770 (.A(_00071_),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold1771 (.A(_02816_),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\m_sys.m_bootloader.r_cstate[2] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold1773 (.A(uio_oe[5]),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\m_sys._m_ram_io_b_port_rdata[28] ),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\m_sys.m_core.m_alu.io_i_uop[0] ),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\m_sys._m_core_io_b_mem_wdata[28] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\m_sys._m_ram_io_b_port_rdata[31] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\m_sys._m_ram_io_b_port_rdata[26] ),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\m_sys._m_ram_io_b_port_rdata[29] ),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\m_sys.m_core.m_bru.io_i_s1[6] ),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold1781 (.A(uio_oe[0]),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold1782 (.A(uio_oe[2]),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold1783 (.A(_00068_),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold1784 (.A(_00166_),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold1785 (.A(uio_oe[1]),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold1786 (.A(uio_oe[3]),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\m_sys._m_core_io_b_mem_wdata[26] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\m_sys.m_core.m_bru.io_i_s1[28] ),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\m_sys._m_core_io_b_mem_wdata[24] ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\m_sys._m_uart_io_o_bl_data[0] ),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold1791 (.A(_00026_),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\m_sys.m_core._m_decoder_io_o_ctrl_wb_addr[2] ),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\m_sys.m_core.m_bru.io_i_pc[5] ),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\m_sys.m_core.m_bru.io_i_pc[8] ),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\m_sys.m_core.m_fsm.r_cstate[3] ),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\m_sys.m_core.m_gpr._GEN[187] ),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[9] ),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\m_sys.m_uart.m_rx.r_cycle_cnt[0] ),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\m_sys._m_bootloader_io_b_mem_addr[7] ),
    .X(net3452));
 sg13g2_antennanp ANTENNA_1 (.A(_04247_));
 sg13g2_antennanp ANTENNA_2 (.A(_04334_));
 sg13g2_antennanp ANTENNA_3 (.A(_04371_));
 sg13g2_antennanp ANTENNA_4 (.A(_04455_));
 sg13g2_antennanp ANTENNA_5 (.A(_04497_));
 sg13g2_antennanp ANTENNA_6 (.A(_04541_));
 sg13g2_antennanp ANTENNA_7 (.A(_04579_));
 sg13g2_antennanp ANTENNA_8 (.A(_04615_));
 sg13g2_antennanp ANTENNA_9 (.A(_04650_));
 sg13g2_antennanp ANTENNA_10 (.A(_04733_));
 sg13g2_antennanp ANTENNA_11 (.A(_04774_));
 sg13g2_antennanp ANTENNA_12 (.A(_04810_));
 sg13g2_antennanp ANTENNA_13 (.A(_04843_));
 sg13g2_antennanp ANTENNA_14 (.A(_04883_));
 sg13g2_antennanp ANTENNA_15 (.A(_05153_));
 sg13g2_antennanp ANTENNA_16 (.A(_05153_));
 sg13g2_antennanp ANTENNA_17 (.A(_05153_));
 sg13g2_antennanp ANTENNA_18 (.A(_05153_));
 sg13g2_antennanp ANTENNA_19 (.A(_05153_));
 sg13g2_antennanp ANTENNA_20 (.A(_05155_));
 sg13g2_antennanp ANTENNA_21 (.A(_05155_));
 sg13g2_antennanp ANTENNA_22 (.A(_05155_));
 sg13g2_antennanp ANTENNA_23 (.A(_05155_));
 sg13g2_antennanp ANTENNA_24 (.A(_05183_));
 sg13g2_antennanp ANTENNA_25 (.A(_05183_));
 sg13g2_antennanp ANTENNA_26 (.A(_05183_));
 sg13g2_antennanp ANTENNA_27 (.A(_05183_));
 sg13g2_antennanp ANTENNA_28 (.A(_05183_));
 sg13g2_antennanp ANTENNA_29 (.A(_05183_));
 sg13g2_antennanp ANTENNA_30 (.A(_05183_));
 sg13g2_antennanp ANTENNA_31 (.A(_05183_));
 sg13g2_antennanp ANTENNA_32 (.A(_05371_));
 sg13g2_antennanp ANTENNA_33 (.A(_05371_));
 sg13g2_antennanp ANTENNA_34 (.A(_05371_));
 sg13g2_antennanp ANTENNA_35 (.A(_05371_));
 sg13g2_antennanp ANTENNA_36 (.A(_05371_));
 sg13g2_antennanp ANTENNA_37 (.A(_05371_));
 sg13g2_antennanp ANTENNA_38 (.A(_05391_));
 sg13g2_antennanp ANTENNA_39 (.A(_05391_));
 sg13g2_antennanp ANTENNA_40 (.A(_05391_));
 sg13g2_antennanp ANTENNA_41 (.A(_05391_));
 sg13g2_antennanp ANTENNA_42 (.A(_05391_));
 sg13g2_antennanp ANTENNA_43 (.A(_05391_));
 sg13g2_antennanp ANTENNA_44 (.A(_05391_));
 sg13g2_antennanp ANTENNA_45 (.A(_05459_));
 sg13g2_antennanp ANTENNA_46 (.A(_05459_));
 sg13g2_antennanp ANTENNA_47 (.A(_05459_));
 sg13g2_antennanp ANTENNA_48 (.A(_05459_));
 sg13g2_antennanp ANTENNA_49 (.A(_05459_));
 sg13g2_antennanp ANTENNA_50 (.A(_05459_));
 sg13g2_antennanp ANTENNA_51 (.A(_05459_));
 sg13g2_antennanp ANTENNA_52 (.A(_05459_));
 sg13g2_antennanp ANTENNA_53 (.A(_05459_));
 sg13g2_antennanp ANTENNA_54 (.A(_05459_));
 sg13g2_antennanp ANTENNA_55 (.A(_05459_));
 sg13g2_antennanp ANTENNA_56 (.A(_05459_));
 sg13g2_antennanp ANTENNA_57 (.A(_05459_));
 sg13g2_antennanp ANTENNA_58 (.A(_05459_));
 sg13g2_antennanp ANTENNA_59 (.A(_05459_));
 sg13g2_antennanp ANTENNA_60 (.A(_05459_));
 sg13g2_antennanp ANTENNA_61 (.A(_05459_));
 sg13g2_antennanp ANTENNA_62 (.A(_05459_));
 sg13g2_antennanp ANTENNA_63 (.A(_05459_));
 sg13g2_antennanp ANTENNA_64 (.A(_05459_));
 sg13g2_antennanp ANTENNA_65 (.A(_05459_));
 sg13g2_antennanp ANTENNA_66 (.A(_05459_));
 sg13g2_antennanp ANTENNA_67 (.A(_05459_));
 sg13g2_antennanp ANTENNA_68 (.A(_05459_));
 sg13g2_antennanp ANTENNA_69 (.A(_05551_));
 sg13g2_antennanp ANTENNA_70 (.A(_05551_));
 sg13g2_antennanp ANTENNA_71 (.A(_05551_));
 sg13g2_antennanp ANTENNA_72 (.A(_05551_));
 sg13g2_antennanp ANTENNA_73 (.A(_05562_));
 sg13g2_antennanp ANTENNA_74 (.A(_05562_));
 sg13g2_antennanp ANTENNA_75 (.A(_05562_));
 sg13g2_antennanp ANTENNA_76 (.A(_05562_));
 sg13g2_antennanp ANTENNA_77 (.A(_05678_));
 sg13g2_antennanp ANTENNA_78 (.A(_05678_));
 sg13g2_antennanp ANTENNA_79 (.A(_05678_));
 sg13g2_antennanp ANTENNA_80 (.A(_05678_));
 sg13g2_antennanp ANTENNA_81 (.A(_05774_));
 sg13g2_antennanp ANTENNA_82 (.A(_05774_));
 sg13g2_antennanp ANTENNA_83 (.A(_05774_));
 sg13g2_antennanp ANTENNA_84 (.A(_05774_));
 sg13g2_antennanp ANTENNA_85 (.A(_05774_));
 sg13g2_antennanp ANTENNA_86 (.A(_05774_));
 sg13g2_antennanp ANTENNA_87 (.A(_05774_));
 sg13g2_antennanp ANTENNA_88 (.A(_05774_));
 sg13g2_antennanp ANTENNA_89 (.A(_05774_));
 sg13g2_antennanp ANTENNA_90 (.A(_05774_));
 sg13g2_antennanp ANTENNA_91 (.A(_06479_));
 sg13g2_antennanp ANTENNA_92 (.A(_06507_));
 sg13g2_antennanp ANTENNA_93 (.A(_06619_));
 sg13g2_antennanp ANTENNA_94 (.A(_06703_));
 sg13g2_antennanp ANTENNA_95 (.A(_06815_));
 sg13g2_antennanp ANTENNA_96 (.A(_06843_));
 sg13g2_antennanp ANTENNA_97 (.A(_07400_));
 sg13g2_antennanp ANTENNA_98 (.A(_07400_));
 sg13g2_antennanp ANTENNA_99 (.A(_07400_));
 sg13g2_antennanp ANTENNA_100 (.A(_07400_));
 sg13g2_antennanp ANTENNA_101 (.A(_07400_));
 sg13g2_antennanp ANTENNA_102 (.A(_07400_));
 sg13g2_antennanp ANTENNA_103 (.A(_07400_));
 sg13g2_antennanp ANTENNA_104 (.A(_07400_));
 sg13g2_antennanp ANTENNA_105 (.A(clk));
 sg13g2_antennanp ANTENNA_106 (.A(clk));
 sg13g2_antennanp ANTENNA_107 (.A(uio_out[4]));
 sg13g2_antennanp ANTENNA_108 (.A(_00074_));
 sg13g2_antennanp ANTENNA_109 (.A(_00074_));
 sg13g2_antennanp ANTENNA_110 (.A(_00074_));
 sg13g2_antennanp ANTENNA_111 (.A(_00074_));
 sg13g2_antennanp ANTENNA_112 (.A(_00074_));
 sg13g2_antennanp ANTENNA_113 (.A(_04334_));
 sg13g2_antennanp ANTENNA_114 (.A(_04371_));
 sg13g2_antennanp ANTENNA_115 (.A(_04455_));
 sg13g2_antennanp ANTENNA_116 (.A(_04497_));
 sg13g2_antennanp ANTENNA_117 (.A(_04541_));
 sg13g2_antennanp ANTENNA_118 (.A(_04579_));
 sg13g2_antennanp ANTENNA_119 (.A(_04615_));
 sg13g2_antennanp ANTENNA_120 (.A(_04733_));
 sg13g2_antennanp ANTENNA_121 (.A(_04774_));
 sg13g2_antennanp ANTENNA_122 (.A(_04810_));
 sg13g2_antennanp ANTENNA_123 (.A(_04843_));
 sg13g2_antennanp ANTENNA_124 (.A(_04883_));
 sg13g2_antennanp ANTENNA_125 (.A(_05155_));
 sg13g2_antennanp ANTENNA_126 (.A(_05155_));
 sg13g2_antennanp ANTENNA_127 (.A(_05155_));
 sg13g2_antennanp ANTENNA_128 (.A(_05155_));
 sg13g2_antennanp ANTENNA_129 (.A(_05155_));
 sg13g2_antennanp ANTENNA_130 (.A(_05155_));
 sg13g2_antennanp ANTENNA_131 (.A(_05155_));
 sg13g2_antennanp ANTENNA_132 (.A(_05155_));
 sg13g2_antennanp ANTENNA_133 (.A(_05155_));
 sg13g2_antennanp ANTENNA_134 (.A(_05155_));
 sg13g2_antennanp ANTENNA_135 (.A(_05155_));
 sg13g2_antennanp ANTENNA_136 (.A(_05155_));
 sg13g2_antennanp ANTENNA_137 (.A(_05155_));
 sg13g2_antennanp ANTENNA_138 (.A(_05155_));
 sg13g2_antennanp ANTENNA_139 (.A(_05155_));
 sg13g2_antennanp ANTENNA_140 (.A(_05155_));
 sg13g2_antennanp ANTENNA_141 (.A(_05155_));
 sg13g2_antennanp ANTENNA_142 (.A(_05155_));
 sg13g2_antennanp ANTENNA_143 (.A(_05155_));
 sg13g2_antennanp ANTENNA_144 (.A(_05155_));
 sg13g2_antennanp ANTENNA_145 (.A(_05257_));
 sg13g2_antennanp ANTENNA_146 (.A(_05257_));
 sg13g2_antennanp ANTENNA_147 (.A(_05257_));
 sg13g2_antennanp ANTENNA_148 (.A(_05257_));
 sg13g2_antennanp ANTENNA_149 (.A(_05371_));
 sg13g2_antennanp ANTENNA_150 (.A(_05371_));
 sg13g2_antennanp ANTENNA_151 (.A(_05371_));
 sg13g2_antennanp ANTENNA_152 (.A(_05371_));
 sg13g2_antennanp ANTENNA_153 (.A(_05371_));
 sg13g2_antennanp ANTENNA_154 (.A(_05371_));
 sg13g2_antennanp ANTENNA_155 (.A(_05391_));
 sg13g2_antennanp ANTENNA_156 (.A(_05391_));
 sg13g2_antennanp ANTENNA_157 (.A(_05391_));
 sg13g2_antennanp ANTENNA_158 (.A(_05391_));
 sg13g2_antennanp ANTENNA_159 (.A(_05391_));
 sg13g2_antennanp ANTENNA_160 (.A(_05391_));
 sg13g2_antennanp ANTENNA_161 (.A(_05391_));
 sg13g2_antennanp ANTENNA_162 (.A(_05391_));
 sg13g2_antennanp ANTENNA_163 (.A(_05391_));
 sg13g2_antennanp ANTENNA_164 (.A(_05505_));
 sg13g2_antennanp ANTENNA_165 (.A(_05505_));
 sg13g2_antennanp ANTENNA_166 (.A(_05505_));
 sg13g2_antennanp ANTENNA_167 (.A(_05505_));
 sg13g2_antennanp ANTENNA_168 (.A(_05551_));
 sg13g2_antennanp ANTENNA_169 (.A(_05551_));
 sg13g2_antennanp ANTENNA_170 (.A(_05551_));
 sg13g2_antennanp ANTENNA_171 (.A(_05551_));
 sg13g2_antennanp ANTENNA_172 (.A(_05551_));
 sg13g2_antennanp ANTENNA_173 (.A(_05551_));
 sg13g2_antennanp ANTENNA_174 (.A(_05551_));
 sg13g2_antennanp ANTENNA_175 (.A(_05562_));
 sg13g2_antennanp ANTENNA_176 (.A(_05562_));
 sg13g2_antennanp ANTENNA_177 (.A(_05562_));
 sg13g2_antennanp ANTENNA_178 (.A(_05562_));
 sg13g2_antennanp ANTENNA_179 (.A(_05802_));
 sg13g2_antennanp ANTENNA_180 (.A(_05802_));
 sg13g2_antennanp ANTENNA_181 (.A(_05802_));
 sg13g2_antennanp ANTENNA_182 (.A(_05802_));
 sg13g2_antennanp ANTENNA_183 (.A(_05802_));
 sg13g2_antennanp ANTENNA_184 (.A(_05802_));
 sg13g2_antennanp ANTENNA_185 (.A(_05802_));
 sg13g2_antennanp ANTENNA_186 (.A(_05848_));
 sg13g2_antennanp ANTENNA_187 (.A(_05848_));
 sg13g2_antennanp ANTENNA_188 (.A(_05848_));
 sg13g2_antennanp ANTENNA_189 (.A(_05848_));
 sg13g2_antennanp ANTENNA_190 (.A(_05848_));
 sg13g2_antennanp ANTENNA_191 (.A(_05886_));
 sg13g2_antennanp ANTENNA_192 (.A(_05886_));
 sg13g2_antennanp ANTENNA_193 (.A(_05886_));
 sg13g2_antennanp ANTENNA_194 (.A(_05886_));
 sg13g2_antennanp ANTENNA_195 (.A(_05886_));
 sg13g2_antennanp ANTENNA_196 (.A(_05886_));
 sg13g2_antennanp ANTENNA_197 (.A(_05886_));
 sg13g2_antennanp ANTENNA_198 (.A(_06507_));
 sg13g2_antennanp ANTENNA_199 (.A(_06619_));
 sg13g2_antennanp ANTENNA_200 (.A(_06815_));
 sg13g2_antennanp ANTENNA_201 (.A(clk));
 sg13g2_antennanp ANTENNA_202 (.A(clk));
 sg13g2_antennanp ANTENNA_203 (.A(uio_out[4]));
 sg13g2_antennanp ANTENNA_204 (.A(_00074_));
 sg13g2_antennanp ANTENNA_205 (.A(_00074_));
 sg13g2_antennanp ANTENNA_206 (.A(_04334_));
 sg13g2_antennanp ANTENNA_207 (.A(_04371_));
 sg13g2_antennanp ANTENNA_208 (.A(_04455_));
 sg13g2_antennanp ANTENNA_209 (.A(_04497_));
 sg13g2_antennanp ANTENNA_210 (.A(_04541_));
 sg13g2_antennanp ANTENNA_211 (.A(_04579_));
 sg13g2_antennanp ANTENNA_212 (.A(_04615_));
 sg13g2_antennanp ANTENNA_213 (.A(_04650_));
 sg13g2_antennanp ANTENNA_214 (.A(_04733_));
 sg13g2_antennanp ANTENNA_215 (.A(_04774_));
 sg13g2_antennanp ANTENNA_216 (.A(_04843_));
 sg13g2_antennanp ANTENNA_217 (.A(_04883_));
 sg13g2_antennanp ANTENNA_218 (.A(_05155_));
 sg13g2_antennanp ANTENNA_219 (.A(_05155_));
 sg13g2_antennanp ANTENNA_220 (.A(_05155_));
 sg13g2_antennanp ANTENNA_221 (.A(_05155_));
 sg13g2_antennanp ANTENNA_222 (.A(_05155_));
 sg13g2_antennanp ANTENNA_223 (.A(_05155_));
 sg13g2_antennanp ANTENNA_224 (.A(_05155_));
 sg13g2_antennanp ANTENNA_225 (.A(_05155_));
 sg13g2_antennanp ANTENNA_226 (.A(_05155_));
 sg13g2_antennanp ANTENNA_227 (.A(_05155_));
 sg13g2_antennanp ANTENNA_228 (.A(_05155_));
 sg13g2_antennanp ANTENNA_229 (.A(_05155_));
 sg13g2_antennanp ANTENNA_230 (.A(_05155_));
 sg13g2_antennanp ANTENNA_231 (.A(_05155_));
 sg13g2_antennanp ANTENNA_232 (.A(_05155_));
 sg13g2_antennanp ANTENNA_233 (.A(_05155_));
 sg13g2_antennanp ANTENNA_234 (.A(_05155_));
 sg13g2_antennanp ANTENNA_235 (.A(_05155_));
 sg13g2_antennanp ANTENNA_236 (.A(_05257_));
 sg13g2_antennanp ANTENNA_237 (.A(_05257_));
 sg13g2_antennanp ANTENNA_238 (.A(_05257_));
 sg13g2_antennanp ANTENNA_239 (.A(_05257_));
 sg13g2_antennanp ANTENNA_240 (.A(_05371_));
 sg13g2_antennanp ANTENNA_241 (.A(_05371_));
 sg13g2_antennanp ANTENNA_242 (.A(_05371_));
 sg13g2_antennanp ANTENNA_243 (.A(_05371_));
 sg13g2_antennanp ANTENNA_244 (.A(_05371_));
 sg13g2_antennanp ANTENNA_245 (.A(_05371_));
 sg13g2_antennanp ANTENNA_246 (.A(_05371_));
 sg13g2_antennanp ANTENNA_247 (.A(_05371_));
 sg13g2_antennanp ANTENNA_248 (.A(_05505_));
 sg13g2_antennanp ANTENNA_249 (.A(_05505_));
 sg13g2_antennanp ANTENNA_250 (.A(_05505_));
 sg13g2_antennanp ANTENNA_251 (.A(_05505_));
 sg13g2_antennanp ANTENNA_252 (.A(_05551_));
 sg13g2_antennanp ANTENNA_253 (.A(_05551_));
 sg13g2_antennanp ANTENNA_254 (.A(_05551_));
 sg13g2_antennanp ANTENNA_255 (.A(_05551_));
 sg13g2_antennanp ANTENNA_256 (.A(_05562_));
 sg13g2_antennanp ANTENNA_257 (.A(_05562_));
 sg13g2_antennanp ANTENNA_258 (.A(_05562_));
 sg13g2_antennanp ANTENNA_259 (.A(_05562_));
 sg13g2_antennanp ANTENNA_260 (.A(_05774_));
 sg13g2_antennanp ANTENNA_261 (.A(_05774_));
 sg13g2_antennanp ANTENNA_262 (.A(_05774_));
 sg13g2_antennanp ANTENNA_263 (.A(_05774_));
 sg13g2_antennanp ANTENNA_264 (.A(_05774_));
 sg13g2_antennanp ANTENNA_265 (.A(_05774_));
 sg13g2_antennanp ANTENNA_266 (.A(_05774_));
 sg13g2_antennanp ANTENNA_267 (.A(_05774_));
 sg13g2_antennanp ANTENNA_268 (.A(_05886_));
 sg13g2_antennanp ANTENNA_269 (.A(_05886_));
 sg13g2_antennanp ANTENNA_270 (.A(_05886_));
 sg13g2_antennanp ANTENNA_271 (.A(_05886_));
 sg13g2_antennanp ANTENNA_272 (.A(_05886_));
 sg13g2_antennanp ANTENNA_273 (.A(_05886_));
 sg13g2_antennanp ANTENNA_274 (.A(_05886_));
 sg13g2_antennanp ANTENNA_275 (.A(_06507_));
 sg13g2_antennanp ANTENNA_276 (.A(_06815_));
 sg13g2_antennanp ANTENNA_277 (.A(_07400_));
 sg13g2_antennanp ANTENNA_278 (.A(_07400_));
 sg13g2_antennanp ANTENNA_279 (.A(_07400_));
 sg13g2_antennanp ANTENNA_280 (.A(_07400_));
 sg13g2_antennanp ANTENNA_281 (.A(_07400_));
 sg13g2_antennanp ANTENNA_282 (.A(_07400_));
 sg13g2_antennanp ANTENNA_283 (.A(_07400_));
 sg13g2_antennanp ANTENNA_284 (.A(clk));
 sg13g2_antennanp ANTENNA_285 (.A(clk));
 sg13g2_antennanp ANTENNA_286 (.A(uio_out[4]));
 sg13g2_antennanp ANTENNA_287 (.A(uio_out[4]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_4 FILLER_0_273 ();
 sg13g2_fill_1 FILLER_0_277 ();
 sg13g2_decap_4 FILLER_0_282 ();
 sg13g2_fill_1 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_fill_2 FILLER_0_517 ();
 sg13g2_fill_1 FILLER_0_519 ();
 sg13g2_fill_1 FILLER_0_589 ();
 sg13g2_fill_2 FILLER_0_599 ();
 sg13g2_fill_1 FILLER_0_601 ();
 sg13g2_fill_1 FILLER_0_667 ();
 sg13g2_fill_2 FILLER_0_677 ();
 sg13g2_fill_1 FILLER_0_679 ();
 sg13g2_fill_1 FILLER_0_684 ();
 sg13g2_fill_1 FILLER_0_729 ();
 sg13g2_fill_2 FILLER_0_746 ();
 sg13g2_fill_1 FILLER_0_748 ();
 sg13g2_fill_1 FILLER_0_754 ();
 sg13g2_fill_1 FILLER_0_767 ();
 sg13g2_fill_2 FILLER_0_782 ();
 sg13g2_decap_8 FILLER_0_796 ();
 sg13g2_decap_4 FILLER_0_803 ();
 sg13g2_fill_2 FILLER_0_807 ();
 sg13g2_fill_1 FILLER_0_835 ();
 sg13g2_fill_1 FILLER_0_864 ();
 sg13g2_fill_1 FILLER_0_903 ();
 sg13g2_fill_2 FILLER_0_908 ();
 sg13g2_fill_1 FILLER_0_910 ();
 sg13g2_fill_1 FILLER_0_916 ();
 sg13g2_fill_1 FILLER_0_952 ();
 sg13g2_fill_2 FILLER_0_967 ();
 sg13g2_fill_1 FILLER_0_969 ();
 sg13g2_fill_2 FILLER_0_983 ();
 sg13g2_fill_1 FILLER_0_1025 ();
 sg13g2_fill_2 FILLER_0_1092 ();
 sg13g2_fill_1 FILLER_0_1132 ();
 sg13g2_fill_2 FILLER_0_1159 ();
 sg13g2_fill_1 FILLER_0_1161 ();
 sg13g2_decap_8 FILLER_0_1244 ();
 sg13g2_decap_8 FILLER_0_1251 ();
 sg13g2_decap_8 FILLER_0_1258 ();
 sg13g2_decap_8 FILLER_0_1265 ();
 sg13g2_decap_8 FILLER_0_1272 ();
 sg13g2_decap_8 FILLER_0_1279 ();
 sg13g2_decap_8 FILLER_0_1286 ();
 sg13g2_decap_8 FILLER_0_1293 ();
 sg13g2_decap_8 FILLER_0_1300 ();
 sg13g2_decap_8 FILLER_0_1307 ();
 sg13g2_decap_8 FILLER_0_1314 ();
 sg13g2_decap_8 FILLER_0_1321 ();
 sg13g2_decap_8 FILLER_0_1328 ();
 sg13g2_decap_8 FILLER_0_1335 ();
 sg13g2_decap_8 FILLER_0_1342 ();
 sg13g2_decap_8 FILLER_0_1349 ();
 sg13g2_decap_8 FILLER_0_1356 ();
 sg13g2_decap_8 FILLER_0_1363 ();
 sg13g2_decap_8 FILLER_0_1370 ();
 sg13g2_decap_8 FILLER_0_1377 ();
 sg13g2_decap_8 FILLER_0_1384 ();
 sg13g2_decap_8 FILLER_0_1391 ();
 sg13g2_decap_8 FILLER_0_1398 ();
 sg13g2_decap_8 FILLER_0_1405 ();
 sg13g2_decap_8 FILLER_0_1412 ();
 sg13g2_decap_8 FILLER_0_1419 ();
 sg13g2_decap_8 FILLER_0_1426 ();
 sg13g2_decap_8 FILLER_0_1433 ();
 sg13g2_decap_8 FILLER_0_1440 ();
 sg13g2_decap_8 FILLER_0_1447 ();
 sg13g2_decap_8 FILLER_0_1454 ();
 sg13g2_decap_8 FILLER_0_1461 ();
 sg13g2_decap_8 FILLER_0_1468 ();
 sg13g2_decap_8 FILLER_0_1475 ();
 sg13g2_decap_8 FILLER_0_1482 ();
 sg13g2_decap_8 FILLER_0_1489 ();
 sg13g2_decap_8 FILLER_0_1496 ();
 sg13g2_decap_8 FILLER_0_1503 ();
 sg13g2_decap_8 FILLER_0_1510 ();
 sg13g2_decap_8 FILLER_0_1517 ();
 sg13g2_decap_8 FILLER_0_1524 ();
 sg13g2_decap_8 FILLER_0_1531 ();
 sg13g2_decap_8 FILLER_0_1538 ();
 sg13g2_decap_8 FILLER_0_1545 ();
 sg13g2_decap_8 FILLER_0_1552 ();
 sg13g2_decap_8 FILLER_0_1559 ();
 sg13g2_decap_8 FILLER_0_1566 ();
 sg13g2_decap_8 FILLER_0_1573 ();
 sg13g2_decap_8 FILLER_0_1580 ();
 sg13g2_decap_8 FILLER_0_1587 ();
 sg13g2_decap_8 FILLER_0_1594 ();
 sg13g2_decap_8 FILLER_0_1601 ();
 sg13g2_decap_8 FILLER_0_1608 ();
 sg13g2_decap_8 FILLER_0_1615 ();
 sg13g2_decap_8 FILLER_0_1622 ();
 sg13g2_decap_8 FILLER_0_1629 ();
 sg13g2_decap_8 FILLER_0_1636 ();
 sg13g2_decap_8 FILLER_0_1643 ();
 sg13g2_decap_8 FILLER_0_1650 ();
 sg13g2_decap_8 FILLER_0_1657 ();
 sg13g2_decap_8 FILLER_0_1664 ();
 sg13g2_decap_8 FILLER_0_1671 ();
 sg13g2_decap_8 FILLER_0_1678 ();
 sg13g2_decap_8 FILLER_0_1685 ();
 sg13g2_decap_8 FILLER_0_1692 ();
 sg13g2_decap_8 FILLER_0_1699 ();
 sg13g2_decap_8 FILLER_0_1706 ();
 sg13g2_decap_8 FILLER_0_1713 ();
 sg13g2_decap_8 FILLER_0_1720 ();
 sg13g2_decap_8 FILLER_0_1727 ();
 sg13g2_decap_8 FILLER_0_1734 ();
 sg13g2_decap_8 FILLER_0_1741 ();
 sg13g2_decap_8 FILLER_0_1748 ();
 sg13g2_decap_8 FILLER_0_1755 ();
 sg13g2_decap_4 FILLER_0_1762 ();
 sg13g2_fill_2 FILLER_0_1766 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_fill_2 FILLER_1_154 ();
 sg13g2_fill_1 FILLER_1_156 ();
 sg13g2_fill_2 FILLER_1_177 ();
 sg13g2_fill_1 FILLER_1_179 ();
 sg13g2_decap_4 FILLER_1_210 ();
 sg13g2_fill_1 FILLER_1_218 ();
 sg13g2_decap_4 FILLER_1_231 ();
 sg13g2_fill_1 FILLER_1_235 ();
 sg13g2_fill_2 FILLER_1_240 ();
 sg13g2_fill_1 FILLER_1_242 ();
 sg13g2_decap_4 FILLER_1_261 ();
 sg13g2_fill_2 FILLER_1_265 ();
 sg13g2_fill_1 FILLER_1_276 ();
 sg13g2_fill_2 FILLER_1_290 ();
 sg13g2_fill_1 FILLER_1_292 ();
 sg13g2_fill_2 FILLER_1_306 ();
 sg13g2_fill_1 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_321 ();
 sg13g2_decap_8 FILLER_1_328 ();
 sg13g2_decap_4 FILLER_1_335 ();
 sg13g2_fill_1 FILLER_1_339 ();
 sg13g2_fill_2 FILLER_1_349 ();
 sg13g2_fill_2 FILLER_1_458 ();
 sg13g2_fill_1 FILLER_1_460 ();
 sg13g2_fill_2 FILLER_1_496 ();
 sg13g2_fill_2 FILLER_1_530 ();
 sg13g2_fill_1 FILLER_1_532 ();
 sg13g2_fill_2 FILLER_1_542 ();
 sg13g2_fill_2 FILLER_1_554 ();
 sg13g2_fill_1 FILLER_1_556 ();
 sg13g2_fill_2 FILLER_1_640 ();
 sg13g2_fill_1 FILLER_1_642 ();
 sg13g2_fill_2 FILLER_1_713 ();
 sg13g2_fill_1 FILLER_1_715 ();
 sg13g2_decap_4 FILLER_1_799 ();
 sg13g2_fill_1 FILLER_1_803 ();
 sg13g2_decap_4 FILLER_1_880 ();
 sg13g2_fill_1 FILLER_1_884 ();
 sg13g2_fill_2 FILLER_1_943 ();
 sg13g2_fill_2 FILLER_1_1115 ();
 sg13g2_fill_2 FILLER_1_1161 ();
 sg13g2_fill_1 FILLER_1_1163 ();
 sg13g2_fill_2 FILLER_1_1173 ();
 sg13g2_fill_2 FILLER_1_1188 ();
 sg13g2_fill_1 FILLER_1_1190 ();
 sg13g2_fill_2 FILLER_1_1247 ();
 sg13g2_decap_8 FILLER_1_1253 ();
 sg13g2_decap_8 FILLER_1_1260 ();
 sg13g2_decap_8 FILLER_1_1267 ();
 sg13g2_decap_8 FILLER_1_1274 ();
 sg13g2_decap_8 FILLER_1_1281 ();
 sg13g2_decap_8 FILLER_1_1288 ();
 sg13g2_decap_8 FILLER_1_1295 ();
 sg13g2_decap_8 FILLER_1_1302 ();
 sg13g2_decap_8 FILLER_1_1309 ();
 sg13g2_decap_8 FILLER_1_1316 ();
 sg13g2_decap_8 FILLER_1_1323 ();
 sg13g2_decap_8 FILLER_1_1330 ();
 sg13g2_decap_8 FILLER_1_1337 ();
 sg13g2_decap_8 FILLER_1_1344 ();
 sg13g2_decap_8 FILLER_1_1351 ();
 sg13g2_decap_8 FILLER_1_1358 ();
 sg13g2_decap_8 FILLER_1_1365 ();
 sg13g2_decap_8 FILLER_1_1372 ();
 sg13g2_decap_8 FILLER_1_1379 ();
 sg13g2_decap_8 FILLER_1_1386 ();
 sg13g2_decap_8 FILLER_1_1393 ();
 sg13g2_decap_8 FILLER_1_1400 ();
 sg13g2_decap_8 FILLER_1_1407 ();
 sg13g2_decap_8 FILLER_1_1414 ();
 sg13g2_decap_8 FILLER_1_1421 ();
 sg13g2_decap_8 FILLER_1_1428 ();
 sg13g2_decap_8 FILLER_1_1435 ();
 sg13g2_decap_8 FILLER_1_1442 ();
 sg13g2_decap_8 FILLER_1_1449 ();
 sg13g2_decap_8 FILLER_1_1456 ();
 sg13g2_decap_8 FILLER_1_1463 ();
 sg13g2_decap_8 FILLER_1_1470 ();
 sg13g2_decap_8 FILLER_1_1477 ();
 sg13g2_decap_8 FILLER_1_1484 ();
 sg13g2_decap_8 FILLER_1_1491 ();
 sg13g2_decap_8 FILLER_1_1498 ();
 sg13g2_decap_8 FILLER_1_1505 ();
 sg13g2_decap_8 FILLER_1_1512 ();
 sg13g2_decap_8 FILLER_1_1519 ();
 sg13g2_decap_8 FILLER_1_1526 ();
 sg13g2_decap_8 FILLER_1_1533 ();
 sg13g2_decap_8 FILLER_1_1540 ();
 sg13g2_decap_8 FILLER_1_1547 ();
 sg13g2_decap_8 FILLER_1_1554 ();
 sg13g2_decap_8 FILLER_1_1561 ();
 sg13g2_decap_8 FILLER_1_1568 ();
 sg13g2_decap_8 FILLER_1_1575 ();
 sg13g2_decap_8 FILLER_1_1582 ();
 sg13g2_decap_8 FILLER_1_1589 ();
 sg13g2_decap_8 FILLER_1_1596 ();
 sg13g2_decap_8 FILLER_1_1603 ();
 sg13g2_decap_8 FILLER_1_1610 ();
 sg13g2_decap_8 FILLER_1_1617 ();
 sg13g2_decap_8 FILLER_1_1624 ();
 sg13g2_decap_8 FILLER_1_1631 ();
 sg13g2_decap_8 FILLER_1_1638 ();
 sg13g2_decap_8 FILLER_1_1645 ();
 sg13g2_decap_8 FILLER_1_1652 ();
 sg13g2_decap_8 FILLER_1_1659 ();
 sg13g2_decap_8 FILLER_1_1666 ();
 sg13g2_decap_8 FILLER_1_1673 ();
 sg13g2_decap_8 FILLER_1_1680 ();
 sg13g2_decap_8 FILLER_1_1687 ();
 sg13g2_decap_8 FILLER_1_1694 ();
 sg13g2_decap_8 FILLER_1_1701 ();
 sg13g2_decap_8 FILLER_1_1708 ();
 sg13g2_decap_8 FILLER_1_1715 ();
 sg13g2_decap_8 FILLER_1_1722 ();
 sg13g2_decap_8 FILLER_1_1729 ();
 sg13g2_decap_8 FILLER_1_1736 ();
 sg13g2_decap_8 FILLER_1_1743 ();
 sg13g2_decap_8 FILLER_1_1750 ();
 sg13g2_decap_8 FILLER_1_1757 ();
 sg13g2_decap_4 FILLER_1_1764 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_fill_1 FILLER_2_186 ();
 sg13g2_fill_2 FILLER_2_195 ();
 sg13g2_fill_1 FILLER_2_231 ();
 sg13g2_fill_1 FILLER_2_266 ();
 sg13g2_fill_1 FILLER_2_297 ();
 sg13g2_decap_8 FILLER_2_324 ();
 sg13g2_fill_1 FILLER_2_484 ();
 sg13g2_fill_1 FILLER_2_515 ();
 sg13g2_fill_1 FILLER_2_529 ();
 sg13g2_fill_1 FILLER_2_561 ();
 sg13g2_fill_2 FILLER_2_660 ();
 sg13g2_fill_2 FILLER_2_686 ();
 sg13g2_fill_1 FILLER_2_688 ();
 sg13g2_fill_1 FILLER_2_694 ();
 sg13g2_fill_1 FILLER_2_701 ();
 sg13g2_fill_2 FILLER_2_708 ();
 sg13g2_fill_1 FILLER_2_710 ();
 sg13g2_fill_1 FILLER_2_730 ();
 sg13g2_fill_2 FILLER_2_740 ();
 sg13g2_fill_2 FILLER_2_751 ();
 sg13g2_fill_1 FILLER_2_798 ();
 sg13g2_decap_4 FILLER_2_915 ();
 sg13g2_fill_2 FILLER_2_932 ();
 sg13g2_fill_1 FILLER_2_984 ();
 sg13g2_fill_2 FILLER_2_1004 ();
 sg13g2_fill_2 FILLER_2_1041 ();
 sg13g2_fill_1 FILLER_2_1043 ();
 sg13g2_fill_2 FILLER_2_1084 ();
 sg13g2_fill_1 FILLER_2_1086 ();
 sg13g2_fill_1 FILLER_2_1149 ();
 sg13g2_fill_1 FILLER_2_1202 ();
 sg13g2_fill_1 FILLER_2_1212 ();
 sg13g2_fill_2 FILLER_2_1222 ();
 sg13g2_decap_8 FILLER_2_1276 ();
 sg13g2_decap_8 FILLER_2_1283 ();
 sg13g2_decap_8 FILLER_2_1290 ();
 sg13g2_decap_8 FILLER_2_1297 ();
 sg13g2_decap_8 FILLER_2_1304 ();
 sg13g2_decap_8 FILLER_2_1311 ();
 sg13g2_decap_4 FILLER_2_1318 ();
 sg13g2_decap_8 FILLER_2_1326 ();
 sg13g2_decap_8 FILLER_2_1333 ();
 sg13g2_decap_8 FILLER_2_1340 ();
 sg13g2_decap_8 FILLER_2_1351 ();
 sg13g2_fill_1 FILLER_2_1358 ();
 sg13g2_decap_8 FILLER_2_1363 ();
 sg13g2_fill_1 FILLER_2_1370 ();
 sg13g2_decap_8 FILLER_2_1379 ();
 sg13g2_decap_8 FILLER_2_1386 ();
 sg13g2_decap_8 FILLER_2_1393 ();
 sg13g2_decap_8 FILLER_2_1400 ();
 sg13g2_decap_8 FILLER_2_1407 ();
 sg13g2_decap_8 FILLER_2_1414 ();
 sg13g2_decap_8 FILLER_2_1421 ();
 sg13g2_decap_8 FILLER_2_1428 ();
 sg13g2_decap_8 FILLER_2_1435 ();
 sg13g2_decap_8 FILLER_2_1442 ();
 sg13g2_decap_8 FILLER_2_1449 ();
 sg13g2_decap_8 FILLER_2_1456 ();
 sg13g2_decap_8 FILLER_2_1463 ();
 sg13g2_decap_8 FILLER_2_1470 ();
 sg13g2_decap_8 FILLER_2_1477 ();
 sg13g2_decap_8 FILLER_2_1484 ();
 sg13g2_decap_8 FILLER_2_1491 ();
 sg13g2_decap_8 FILLER_2_1498 ();
 sg13g2_decap_8 FILLER_2_1505 ();
 sg13g2_decap_8 FILLER_2_1512 ();
 sg13g2_decap_8 FILLER_2_1519 ();
 sg13g2_decap_8 FILLER_2_1526 ();
 sg13g2_decap_8 FILLER_2_1533 ();
 sg13g2_decap_8 FILLER_2_1540 ();
 sg13g2_decap_8 FILLER_2_1547 ();
 sg13g2_decap_8 FILLER_2_1554 ();
 sg13g2_decap_8 FILLER_2_1561 ();
 sg13g2_decap_8 FILLER_2_1568 ();
 sg13g2_decap_8 FILLER_2_1575 ();
 sg13g2_decap_8 FILLER_2_1582 ();
 sg13g2_decap_8 FILLER_2_1589 ();
 sg13g2_decap_8 FILLER_2_1596 ();
 sg13g2_decap_8 FILLER_2_1603 ();
 sg13g2_decap_8 FILLER_2_1610 ();
 sg13g2_decap_8 FILLER_2_1617 ();
 sg13g2_decap_8 FILLER_2_1624 ();
 sg13g2_decap_8 FILLER_2_1631 ();
 sg13g2_decap_8 FILLER_2_1638 ();
 sg13g2_decap_8 FILLER_2_1645 ();
 sg13g2_decap_8 FILLER_2_1652 ();
 sg13g2_decap_8 FILLER_2_1659 ();
 sg13g2_decap_8 FILLER_2_1666 ();
 sg13g2_decap_8 FILLER_2_1673 ();
 sg13g2_decap_8 FILLER_2_1680 ();
 sg13g2_decap_8 FILLER_2_1687 ();
 sg13g2_decap_8 FILLER_2_1694 ();
 sg13g2_decap_8 FILLER_2_1701 ();
 sg13g2_decap_8 FILLER_2_1708 ();
 sg13g2_decap_8 FILLER_2_1715 ();
 sg13g2_decap_8 FILLER_2_1722 ();
 sg13g2_decap_8 FILLER_2_1729 ();
 sg13g2_decap_8 FILLER_2_1736 ();
 sg13g2_decap_8 FILLER_2_1743 ();
 sg13g2_decap_8 FILLER_2_1750 ();
 sg13g2_decap_8 FILLER_2_1757 ();
 sg13g2_decap_4 FILLER_2_1764 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_fill_2 FILLER_3_105 ();
 sg13g2_decap_4 FILLER_3_115 ();
 sg13g2_decap_4 FILLER_3_123 ();
 sg13g2_fill_2 FILLER_3_167 ();
 sg13g2_fill_1 FILLER_3_169 ();
 sg13g2_fill_1 FILLER_3_190 ();
 sg13g2_fill_2 FILLER_3_223 ();
 sg13g2_fill_1 FILLER_3_225 ();
 sg13g2_fill_2 FILLER_3_252 ();
 sg13g2_fill_1 FILLER_3_254 ();
 sg13g2_fill_2 FILLER_3_280 ();
 sg13g2_fill_2 FILLER_3_344 ();
 sg13g2_fill_1 FILLER_3_424 ();
 sg13g2_fill_1 FILLER_3_480 ();
 sg13g2_fill_2 FILLER_3_525 ();
 sg13g2_fill_1 FILLER_3_527 ();
 sg13g2_fill_2 FILLER_3_546 ();
 sg13g2_fill_1 FILLER_3_582 ();
 sg13g2_fill_1 FILLER_3_592 ();
 sg13g2_fill_2 FILLER_3_610 ();
 sg13g2_fill_1 FILLER_3_626 ();
 sg13g2_fill_1 FILLER_3_705 ();
 sg13g2_fill_1 FILLER_3_732 ();
 sg13g2_decap_8 FILLER_3_800 ();
 sg13g2_fill_2 FILLER_3_807 ();
 sg13g2_fill_1 FILLER_3_809 ();
 sg13g2_fill_2 FILLER_3_848 ();
 sg13g2_fill_1 FILLER_3_892 ();
 sg13g2_fill_1 FILLER_3_936 ();
 sg13g2_fill_1 FILLER_3_974 ();
 sg13g2_fill_2 FILLER_3_1030 ();
 sg13g2_fill_1 FILLER_3_1041 ();
 sg13g2_fill_2 FILLER_3_1066 ();
 sg13g2_fill_2 FILLER_3_1086 ();
 sg13g2_fill_1 FILLER_3_1088 ();
 sg13g2_fill_1 FILLER_3_1112 ();
 sg13g2_fill_1 FILLER_3_1122 ();
 sg13g2_fill_2 FILLER_3_1136 ();
 sg13g2_fill_1 FILLER_3_1143 ();
 sg13g2_fill_1 FILLER_3_1179 ();
 sg13g2_fill_1 FILLER_3_1189 ();
 sg13g2_fill_2 FILLER_3_1224 ();
 sg13g2_fill_1 FILLER_3_1226 ();
 sg13g2_fill_2 FILLER_3_1261 ();
 sg13g2_fill_2 FILLER_3_1288 ();
 sg13g2_fill_1 FILLER_3_1290 ();
 sg13g2_decap_8 FILLER_3_1303 ();
 sg13g2_decap_4 FILLER_3_1310 ();
 sg13g2_fill_1 FILLER_3_1314 ();
 sg13g2_decap_4 FILLER_3_1337 ();
 sg13g2_fill_2 FILLER_3_1341 ();
 sg13g2_fill_2 FILLER_3_1347 ();
 sg13g2_fill_1 FILLER_3_1353 ();
 sg13g2_decap_8 FILLER_3_1397 ();
 sg13g2_decap_8 FILLER_3_1404 ();
 sg13g2_decap_8 FILLER_3_1411 ();
 sg13g2_decap_8 FILLER_3_1418 ();
 sg13g2_decap_8 FILLER_3_1425 ();
 sg13g2_fill_2 FILLER_3_1432 ();
 sg13g2_decap_8 FILLER_3_1446 ();
 sg13g2_decap_8 FILLER_3_1453 ();
 sg13g2_decap_8 FILLER_3_1460 ();
 sg13g2_decap_8 FILLER_3_1467 ();
 sg13g2_decap_8 FILLER_3_1474 ();
 sg13g2_decap_8 FILLER_3_1481 ();
 sg13g2_decap_8 FILLER_3_1488 ();
 sg13g2_decap_8 FILLER_3_1495 ();
 sg13g2_decap_8 FILLER_3_1502 ();
 sg13g2_decap_8 FILLER_3_1509 ();
 sg13g2_decap_8 FILLER_3_1516 ();
 sg13g2_decap_8 FILLER_3_1523 ();
 sg13g2_decap_8 FILLER_3_1530 ();
 sg13g2_decap_8 FILLER_3_1537 ();
 sg13g2_decap_8 FILLER_3_1544 ();
 sg13g2_decap_8 FILLER_3_1551 ();
 sg13g2_decap_8 FILLER_3_1558 ();
 sg13g2_decap_8 FILLER_3_1565 ();
 sg13g2_decap_8 FILLER_3_1572 ();
 sg13g2_decap_8 FILLER_3_1579 ();
 sg13g2_decap_8 FILLER_3_1586 ();
 sg13g2_decap_8 FILLER_3_1593 ();
 sg13g2_decap_8 FILLER_3_1600 ();
 sg13g2_decap_8 FILLER_3_1607 ();
 sg13g2_decap_8 FILLER_3_1614 ();
 sg13g2_decap_8 FILLER_3_1621 ();
 sg13g2_decap_8 FILLER_3_1628 ();
 sg13g2_decap_8 FILLER_3_1635 ();
 sg13g2_decap_8 FILLER_3_1642 ();
 sg13g2_decap_8 FILLER_3_1649 ();
 sg13g2_decap_8 FILLER_3_1656 ();
 sg13g2_decap_8 FILLER_3_1663 ();
 sg13g2_decap_8 FILLER_3_1670 ();
 sg13g2_decap_8 FILLER_3_1677 ();
 sg13g2_decap_8 FILLER_3_1684 ();
 sg13g2_decap_8 FILLER_3_1691 ();
 sg13g2_decap_8 FILLER_3_1698 ();
 sg13g2_decap_8 FILLER_3_1705 ();
 sg13g2_decap_8 FILLER_3_1712 ();
 sg13g2_decap_8 FILLER_3_1719 ();
 sg13g2_decap_8 FILLER_3_1726 ();
 sg13g2_decap_8 FILLER_3_1733 ();
 sg13g2_decap_8 FILLER_3_1740 ();
 sg13g2_decap_8 FILLER_3_1747 ();
 sg13g2_decap_8 FILLER_3_1754 ();
 sg13g2_decap_8 FILLER_3_1761 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_4 FILLER_4_84 ();
 sg13g2_fill_1 FILLER_4_88 ();
 sg13g2_fill_2 FILLER_4_109 ();
 sg13g2_fill_1 FILLER_4_111 ();
 sg13g2_fill_1 FILLER_4_146 ();
 sg13g2_fill_2 FILLER_4_202 ();
 sg13g2_fill_2 FILLER_4_214 ();
 sg13g2_fill_1 FILLER_4_240 ();
 sg13g2_fill_2 FILLER_4_251 ();
 sg13g2_fill_1 FILLER_4_253 ();
 sg13g2_fill_2 FILLER_4_307 ();
 sg13g2_fill_1 FILLER_4_330 ();
 sg13g2_fill_1 FILLER_4_353 ();
 sg13g2_fill_1 FILLER_4_363 ();
 sg13g2_fill_2 FILLER_4_373 ();
 sg13g2_fill_2 FILLER_4_384 ();
 sg13g2_fill_1 FILLER_4_403 ();
 sg13g2_fill_1 FILLER_4_425 ();
 sg13g2_fill_1 FILLER_4_460 ();
 sg13g2_fill_2 FILLER_4_501 ();
 sg13g2_fill_1 FILLER_4_604 ();
 sg13g2_fill_2 FILLER_4_646 ();
 sg13g2_fill_2 FILLER_4_657 ();
 sg13g2_fill_2 FILLER_4_668 ();
 sg13g2_fill_2 FILLER_4_689 ();
 sg13g2_fill_1 FILLER_4_700 ();
 sg13g2_fill_2 FILLER_4_714 ();
 sg13g2_fill_1 FILLER_4_716 ();
 sg13g2_fill_2 FILLER_4_735 ();
 sg13g2_fill_1 FILLER_4_769 ();
 sg13g2_fill_2 FILLER_4_827 ();
 sg13g2_fill_1 FILLER_4_829 ();
 sg13g2_fill_2 FILLER_4_843 ();
 sg13g2_fill_2 FILLER_4_849 ();
 sg13g2_fill_2 FILLER_4_868 ();
 sg13g2_fill_1 FILLER_4_922 ();
 sg13g2_fill_2 FILLER_4_941 ();
 sg13g2_fill_1 FILLER_4_943 ();
 sg13g2_fill_2 FILLER_4_956 ();
 sg13g2_fill_1 FILLER_4_1011 ();
 sg13g2_fill_1 FILLER_4_1038 ();
 sg13g2_fill_2 FILLER_4_1065 ();
 sg13g2_fill_2 FILLER_4_1158 ();
 sg13g2_fill_2 FILLER_4_1170 ();
 sg13g2_fill_1 FILLER_4_1172 ();
 sg13g2_fill_2 FILLER_4_1187 ();
 sg13g2_fill_1 FILLER_4_1189 ();
 sg13g2_fill_2 FILLER_4_1256 ();
 sg13g2_fill_1 FILLER_4_1258 ();
 sg13g2_fill_1 FILLER_4_1418 ();
 sg13g2_fill_2 FILLER_4_1439 ();
 sg13g2_decap_8 FILLER_4_1461 ();
 sg13g2_decap_8 FILLER_4_1468 ();
 sg13g2_decap_8 FILLER_4_1475 ();
 sg13g2_decap_8 FILLER_4_1482 ();
 sg13g2_decap_8 FILLER_4_1489 ();
 sg13g2_decap_8 FILLER_4_1496 ();
 sg13g2_decap_8 FILLER_4_1503 ();
 sg13g2_decap_8 FILLER_4_1510 ();
 sg13g2_decap_8 FILLER_4_1517 ();
 sg13g2_decap_8 FILLER_4_1524 ();
 sg13g2_decap_8 FILLER_4_1531 ();
 sg13g2_decap_8 FILLER_4_1538 ();
 sg13g2_decap_8 FILLER_4_1545 ();
 sg13g2_decap_8 FILLER_4_1552 ();
 sg13g2_decap_8 FILLER_4_1559 ();
 sg13g2_decap_8 FILLER_4_1566 ();
 sg13g2_decap_8 FILLER_4_1573 ();
 sg13g2_decap_8 FILLER_4_1580 ();
 sg13g2_decap_8 FILLER_4_1587 ();
 sg13g2_decap_8 FILLER_4_1594 ();
 sg13g2_decap_8 FILLER_4_1601 ();
 sg13g2_decap_8 FILLER_4_1608 ();
 sg13g2_decap_8 FILLER_4_1615 ();
 sg13g2_decap_8 FILLER_4_1622 ();
 sg13g2_decap_8 FILLER_4_1629 ();
 sg13g2_decap_8 FILLER_4_1636 ();
 sg13g2_decap_8 FILLER_4_1643 ();
 sg13g2_decap_8 FILLER_4_1650 ();
 sg13g2_decap_8 FILLER_4_1657 ();
 sg13g2_decap_8 FILLER_4_1664 ();
 sg13g2_decap_8 FILLER_4_1671 ();
 sg13g2_decap_8 FILLER_4_1678 ();
 sg13g2_decap_8 FILLER_4_1685 ();
 sg13g2_decap_8 FILLER_4_1692 ();
 sg13g2_decap_8 FILLER_4_1699 ();
 sg13g2_decap_8 FILLER_4_1706 ();
 sg13g2_decap_8 FILLER_4_1713 ();
 sg13g2_decap_8 FILLER_4_1720 ();
 sg13g2_decap_8 FILLER_4_1727 ();
 sg13g2_decap_8 FILLER_4_1734 ();
 sg13g2_decap_8 FILLER_4_1741 ();
 sg13g2_decap_8 FILLER_4_1748 ();
 sg13g2_decap_8 FILLER_4_1755 ();
 sg13g2_decap_4 FILLER_4_1762 ();
 sg13g2_fill_2 FILLER_4_1766 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_fill_1 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_47 ();
 sg13g2_decap_8 FILLER_5_54 ();
 sg13g2_decap_8 FILLER_5_61 ();
 sg13g2_decap_8 FILLER_5_68 ();
 sg13g2_decap_4 FILLER_5_75 ();
 sg13g2_decap_4 FILLER_5_83 ();
 sg13g2_fill_1 FILLER_5_181 ();
 sg13g2_fill_2 FILLER_5_199 ();
 sg13g2_fill_2 FILLER_5_257 ();
 sg13g2_fill_1 FILLER_5_297 ();
 sg13g2_fill_1 FILLER_5_307 ();
 sg13g2_fill_1 FILLER_5_312 ();
 sg13g2_fill_2 FILLER_5_322 ();
 sg13g2_fill_1 FILLER_5_324 ();
 sg13g2_fill_2 FILLER_5_334 ();
 sg13g2_fill_2 FILLER_5_434 ();
 sg13g2_fill_2 FILLER_5_507 ();
 sg13g2_fill_1 FILLER_5_549 ();
 sg13g2_fill_2 FILLER_5_558 ();
 sg13g2_fill_1 FILLER_5_571 ();
 sg13g2_fill_1 FILLER_5_585 ();
 sg13g2_fill_2 FILLER_5_630 ();
 sg13g2_fill_1 FILLER_5_632 ();
 sg13g2_fill_2 FILLER_5_674 ();
 sg13g2_fill_1 FILLER_5_735 ();
 sg13g2_fill_2 FILLER_5_745 ();
 sg13g2_fill_1 FILLER_5_747 ();
 sg13g2_fill_2 FILLER_5_763 ();
 sg13g2_fill_1 FILLER_5_765 ();
 sg13g2_fill_2 FILLER_5_805 ();
 sg13g2_fill_1 FILLER_5_807 ();
 sg13g2_fill_2 FILLER_5_887 ();
 sg13g2_fill_1 FILLER_5_889 ();
 sg13g2_fill_2 FILLER_5_904 ();
 sg13g2_fill_2 FILLER_5_1003 ();
 sg13g2_fill_1 FILLER_5_1005 ();
 sg13g2_fill_2 FILLER_5_1019 ();
 sg13g2_fill_1 FILLER_5_1032 ();
 sg13g2_fill_1 FILLER_5_1046 ();
 sg13g2_fill_2 FILLER_5_1051 ();
 sg13g2_fill_1 FILLER_5_1053 ();
 sg13g2_fill_1 FILLER_5_1097 ();
 sg13g2_fill_2 FILLER_5_1111 ();
 sg13g2_fill_1 FILLER_5_1113 ();
 sg13g2_fill_1 FILLER_5_1146 ();
 sg13g2_fill_1 FILLER_5_1203 ();
 sg13g2_fill_1 FILLER_5_1273 ();
 sg13g2_fill_1 FILLER_5_1323 ();
 sg13g2_fill_2 FILLER_5_1328 ();
 sg13g2_fill_1 FILLER_5_1330 ();
 sg13g2_fill_2 FILLER_5_1351 ();
 sg13g2_fill_1 FILLER_5_1383 ();
 sg13g2_fill_1 FILLER_5_1397 ();
 sg13g2_fill_2 FILLER_5_1402 ();
 sg13g2_fill_1 FILLER_5_1404 ();
 sg13g2_fill_2 FILLER_5_1431 ();
 sg13g2_decap_8 FILLER_5_1458 ();
 sg13g2_decap_8 FILLER_5_1465 ();
 sg13g2_decap_8 FILLER_5_1472 ();
 sg13g2_decap_8 FILLER_5_1479 ();
 sg13g2_decap_8 FILLER_5_1486 ();
 sg13g2_decap_8 FILLER_5_1493 ();
 sg13g2_decap_8 FILLER_5_1500 ();
 sg13g2_decap_8 FILLER_5_1507 ();
 sg13g2_decap_8 FILLER_5_1514 ();
 sg13g2_decap_8 FILLER_5_1521 ();
 sg13g2_decap_8 FILLER_5_1528 ();
 sg13g2_decap_8 FILLER_5_1535 ();
 sg13g2_decap_8 FILLER_5_1542 ();
 sg13g2_decap_8 FILLER_5_1549 ();
 sg13g2_decap_8 FILLER_5_1556 ();
 sg13g2_decap_8 FILLER_5_1563 ();
 sg13g2_decap_8 FILLER_5_1570 ();
 sg13g2_decap_8 FILLER_5_1577 ();
 sg13g2_decap_8 FILLER_5_1584 ();
 sg13g2_decap_8 FILLER_5_1591 ();
 sg13g2_decap_8 FILLER_5_1598 ();
 sg13g2_decap_8 FILLER_5_1605 ();
 sg13g2_decap_8 FILLER_5_1612 ();
 sg13g2_decap_8 FILLER_5_1619 ();
 sg13g2_decap_8 FILLER_5_1626 ();
 sg13g2_decap_8 FILLER_5_1633 ();
 sg13g2_decap_8 FILLER_5_1640 ();
 sg13g2_decap_8 FILLER_5_1647 ();
 sg13g2_decap_8 FILLER_5_1654 ();
 sg13g2_decap_8 FILLER_5_1661 ();
 sg13g2_decap_8 FILLER_5_1668 ();
 sg13g2_decap_8 FILLER_5_1675 ();
 sg13g2_decap_8 FILLER_5_1682 ();
 sg13g2_decap_8 FILLER_5_1689 ();
 sg13g2_decap_8 FILLER_5_1696 ();
 sg13g2_decap_8 FILLER_5_1703 ();
 sg13g2_decap_8 FILLER_5_1710 ();
 sg13g2_decap_8 FILLER_5_1717 ();
 sg13g2_decap_8 FILLER_5_1724 ();
 sg13g2_decap_8 FILLER_5_1731 ();
 sg13g2_decap_8 FILLER_5_1738 ();
 sg13g2_decap_8 FILLER_5_1745 ();
 sg13g2_decap_8 FILLER_5_1752 ();
 sg13g2_decap_8 FILLER_5_1759 ();
 sg13g2_fill_2 FILLER_5_1766 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_21 ();
 sg13g2_fill_2 FILLER_6_46 ();
 sg13g2_fill_1 FILLER_6_48 ();
 sg13g2_decap_4 FILLER_6_66 ();
 sg13g2_fill_1 FILLER_6_70 ();
 sg13g2_fill_2 FILLER_6_75 ();
 sg13g2_fill_1 FILLER_6_103 ();
 sg13g2_fill_2 FILLER_6_116 ();
 sg13g2_fill_1 FILLER_6_118 ();
 sg13g2_fill_1 FILLER_6_123 ();
 sg13g2_fill_2 FILLER_6_205 ();
 sg13g2_fill_2 FILLER_6_213 ();
 sg13g2_fill_2 FILLER_6_224 ();
 sg13g2_fill_2 FILLER_6_381 ();
 sg13g2_fill_2 FILLER_6_392 ();
 sg13g2_fill_2 FILLER_6_498 ();
 sg13g2_fill_2 FILLER_6_509 ();
 sg13g2_fill_1 FILLER_6_584 ();
 sg13g2_fill_2 FILLER_6_599 ();
 sg13g2_fill_2 FILLER_6_607 ();
 sg13g2_fill_1 FILLER_6_641 ();
 sg13g2_fill_1 FILLER_6_707 ();
 sg13g2_fill_1 FILLER_6_760 ();
 sg13g2_fill_2 FILLER_6_792 ();
 sg13g2_fill_1 FILLER_6_794 ();
 sg13g2_fill_2 FILLER_6_807 ();
 sg13g2_fill_1 FILLER_6_822 ();
 sg13g2_fill_1 FILLER_6_837 ();
 sg13g2_fill_2 FILLER_6_843 ();
 sg13g2_fill_1 FILLER_6_845 ();
 sg13g2_fill_2 FILLER_6_954 ();
 sg13g2_fill_1 FILLER_6_956 ();
 sg13g2_fill_1 FILLER_6_995 ();
 sg13g2_fill_2 FILLER_6_1031 ();
 sg13g2_fill_1 FILLER_6_1033 ();
 sg13g2_fill_2 FILLER_6_1047 ();
 sg13g2_fill_1 FILLER_6_1049 ();
 sg13g2_fill_2 FILLER_6_1054 ();
 sg13g2_fill_1 FILLER_6_1056 ();
 sg13g2_fill_2 FILLER_6_1081 ();
 sg13g2_fill_1 FILLER_6_1087 ();
 sg13g2_fill_2 FILLER_6_1093 ();
 sg13g2_fill_1 FILLER_6_1095 ();
 sg13g2_fill_1 FILLER_6_1112 ();
 sg13g2_fill_2 FILLER_6_1127 ();
 sg13g2_fill_1 FILLER_6_1129 ();
 sg13g2_fill_1 FILLER_6_1169 ();
 sg13g2_fill_2 FILLER_6_1195 ();
 sg13g2_fill_1 FILLER_6_1197 ();
 sg13g2_fill_2 FILLER_6_1272 ();
 sg13g2_fill_1 FILLER_6_1274 ();
 sg13g2_fill_2 FILLER_6_1327 ();
 sg13g2_fill_1 FILLER_6_1329 ();
 sg13g2_fill_2 FILLER_6_1370 ();
 sg13g2_fill_1 FILLER_6_1428 ();
 sg13g2_decap_8 FILLER_6_1481 ();
 sg13g2_decap_8 FILLER_6_1488 ();
 sg13g2_decap_8 FILLER_6_1495 ();
 sg13g2_decap_8 FILLER_6_1502 ();
 sg13g2_decap_8 FILLER_6_1509 ();
 sg13g2_decap_8 FILLER_6_1516 ();
 sg13g2_decap_8 FILLER_6_1523 ();
 sg13g2_decap_8 FILLER_6_1530 ();
 sg13g2_decap_8 FILLER_6_1537 ();
 sg13g2_decap_8 FILLER_6_1544 ();
 sg13g2_decap_8 FILLER_6_1551 ();
 sg13g2_decap_8 FILLER_6_1558 ();
 sg13g2_decap_8 FILLER_6_1565 ();
 sg13g2_decap_8 FILLER_6_1572 ();
 sg13g2_decap_8 FILLER_6_1579 ();
 sg13g2_decap_8 FILLER_6_1586 ();
 sg13g2_decap_8 FILLER_6_1593 ();
 sg13g2_decap_8 FILLER_6_1600 ();
 sg13g2_decap_8 FILLER_6_1607 ();
 sg13g2_decap_8 FILLER_6_1614 ();
 sg13g2_decap_8 FILLER_6_1621 ();
 sg13g2_decap_8 FILLER_6_1628 ();
 sg13g2_decap_8 FILLER_6_1635 ();
 sg13g2_decap_8 FILLER_6_1642 ();
 sg13g2_decap_8 FILLER_6_1649 ();
 sg13g2_decap_8 FILLER_6_1656 ();
 sg13g2_decap_8 FILLER_6_1663 ();
 sg13g2_decap_8 FILLER_6_1670 ();
 sg13g2_decap_8 FILLER_6_1677 ();
 sg13g2_decap_8 FILLER_6_1684 ();
 sg13g2_decap_8 FILLER_6_1691 ();
 sg13g2_decap_8 FILLER_6_1698 ();
 sg13g2_decap_8 FILLER_6_1705 ();
 sg13g2_decap_8 FILLER_6_1712 ();
 sg13g2_decap_8 FILLER_6_1719 ();
 sg13g2_decap_8 FILLER_6_1726 ();
 sg13g2_decap_8 FILLER_6_1733 ();
 sg13g2_decap_8 FILLER_6_1740 ();
 sg13g2_decap_8 FILLER_6_1747 ();
 sg13g2_decap_8 FILLER_6_1754 ();
 sg13g2_decap_8 FILLER_6_1761 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_22 ();
 sg13g2_fill_1 FILLER_7_24 ();
 sg13g2_fill_1 FILLER_7_34 ();
 sg13g2_fill_2 FILLER_7_44 ();
 sg13g2_fill_1 FILLER_7_46 ();
 sg13g2_fill_1 FILLER_7_81 ();
 sg13g2_fill_1 FILLER_7_173 ();
 sg13g2_fill_2 FILLER_7_183 ();
 sg13g2_fill_1 FILLER_7_185 ();
 sg13g2_fill_2 FILLER_7_204 ();
 sg13g2_fill_1 FILLER_7_275 ();
 sg13g2_fill_1 FILLER_7_290 ();
 sg13g2_fill_1 FILLER_7_311 ();
 sg13g2_fill_1 FILLER_7_321 ();
 sg13g2_fill_2 FILLER_7_342 ();
 sg13g2_fill_1 FILLER_7_344 ();
 sg13g2_fill_2 FILLER_7_351 ();
 sg13g2_fill_1 FILLER_7_353 ();
 sg13g2_fill_1 FILLER_7_366 ();
 sg13g2_fill_2 FILLER_7_398 ();
 sg13g2_fill_2 FILLER_7_435 ();
 sg13g2_fill_2 FILLER_7_496 ();
 sg13g2_fill_2 FILLER_7_529 ();
 sg13g2_fill_1 FILLER_7_576 ();
 sg13g2_fill_2 FILLER_7_607 ();
 sg13g2_fill_1 FILLER_7_677 ();
 sg13g2_fill_2 FILLER_7_728 ();
 sg13g2_fill_1 FILLER_7_857 ();
 sg13g2_fill_1 FILLER_7_897 ();
 sg13g2_fill_1 FILLER_7_933 ();
 sg13g2_fill_2 FILLER_7_986 ();
 sg13g2_fill_2 FILLER_7_1006 ();
 sg13g2_fill_2 FILLER_7_1022 ();
 sg13g2_fill_1 FILLER_7_1024 ();
 sg13g2_fill_1 FILLER_7_1039 ();
 sg13g2_fill_2 FILLER_7_1092 ();
 sg13g2_fill_1 FILLER_7_1176 ();
 sg13g2_fill_1 FILLER_7_1322 ();
 sg13g2_fill_2 FILLER_7_1349 ();
 sg13g2_fill_2 FILLER_7_1382 ();
 sg13g2_fill_1 FILLER_7_1384 ();
 sg13g2_fill_2 FILLER_7_1433 ();
 sg13g2_fill_2 FILLER_7_1439 ();
 sg13g2_fill_1 FILLER_7_1441 ();
 sg13g2_fill_1 FILLER_7_1447 ();
 sg13g2_decap_8 FILLER_7_1494 ();
 sg13g2_decap_8 FILLER_7_1501 ();
 sg13g2_decap_8 FILLER_7_1508 ();
 sg13g2_decap_8 FILLER_7_1515 ();
 sg13g2_decap_8 FILLER_7_1522 ();
 sg13g2_decap_8 FILLER_7_1529 ();
 sg13g2_decap_8 FILLER_7_1536 ();
 sg13g2_decap_8 FILLER_7_1543 ();
 sg13g2_decap_8 FILLER_7_1550 ();
 sg13g2_decap_8 FILLER_7_1557 ();
 sg13g2_decap_8 FILLER_7_1564 ();
 sg13g2_decap_8 FILLER_7_1571 ();
 sg13g2_decap_8 FILLER_7_1578 ();
 sg13g2_decap_8 FILLER_7_1585 ();
 sg13g2_decap_8 FILLER_7_1592 ();
 sg13g2_decap_8 FILLER_7_1599 ();
 sg13g2_decap_8 FILLER_7_1606 ();
 sg13g2_decap_8 FILLER_7_1613 ();
 sg13g2_decap_8 FILLER_7_1620 ();
 sg13g2_decap_8 FILLER_7_1627 ();
 sg13g2_decap_8 FILLER_7_1634 ();
 sg13g2_decap_8 FILLER_7_1641 ();
 sg13g2_decap_8 FILLER_7_1648 ();
 sg13g2_decap_8 FILLER_7_1655 ();
 sg13g2_decap_8 FILLER_7_1662 ();
 sg13g2_decap_8 FILLER_7_1669 ();
 sg13g2_decap_8 FILLER_7_1676 ();
 sg13g2_decap_8 FILLER_7_1683 ();
 sg13g2_decap_8 FILLER_7_1690 ();
 sg13g2_decap_8 FILLER_7_1697 ();
 sg13g2_decap_8 FILLER_7_1704 ();
 sg13g2_decap_8 FILLER_7_1711 ();
 sg13g2_decap_8 FILLER_7_1718 ();
 sg13g2_decap_8 FILLER_7_1725 ();
 sg13g2_decap_8 FILLER_7_1732 ();
 sg13g2_decap_8 FILLER_7_1739 ();
 sg13g2_decap_8 FILLER_7_1746 ();
 sg13g2_decap_8 FILLER_7_1753 ();
 sg13g2_decap_8 FILLER_7_1760 ();
 sg13g2_fill_1 FILLER_7_1767 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_15 ();
 sg13g2_fill_2 FILLER_8_21 ();
 sg13g2_fill_1 FILLER_8_49 ();
 sg13g2_fill_2 FILLER_8_95 ();
 sg13g2_fill_1 FILLER_8_97 ();
 sg13g2_fill_2 FILLER_8_112 ();
 sg13g2_fill_2 FILLER_8_158 ();
 sg13g2_fill_2 FILLER_8_191 ();
 sg13g2_fill_1 FILLER_8_207 ();
 sg13g2_fill_2 FILLER_8_218 ();
 sg13g2_fill_1 FILLER_8_233 ();
 sg13g2_fill_1 FILLER_8_242 ();
 sg13g2_fill_2 FILLER_8_255 ();
 sg13g2_fill_1 FILLER_8_257 ();
 sg13g2_fill_2 FILLER_8_337 ();
 sg13g2_fill_1 FILLER_8_339 ();
 sg13g2_fill_2 FILLER_8_439 ();
 sg13g2_fill_2 FILLER_8_476 ();
 sg13g2_fill_2 FILLER_8_495 ();
 sg13g2_fill_2 FILLER_8_581 ();
 sg13g2_fill_1 FILLER_8_583 ();
 sg13g2_fill_2 FILLER_8_614 ();
 sg13g2_fill_1 FILLER_8_616 ();
 sg13g2_fill_2 FILLER_8_806 ();
 sg13g2_fill_1 FILLER_8_840 ();
 sg13g2_fill_2 FILLER_8_850 ();
 sg13g2_fill_2 FILLER_8_862 ();
 sg13g2_fill_1 FILLER_8_868 ();
 sg13g2_fill_2 FILLER_8_882 ();
 sg13g2_decap_8 FILLER_8_892 ();
 sg13g2_decap_4 FILLER_8_899 ();
 sg13g2_fill_2 FILLER_8_903 ();
 sg13g2_fill_1 FILLER_8_913 ();
 sg13g2_fill_2 FILLER_8_918 ();
 sg13g2_fill_2 FILLER_8_937 ();
 sg13g2_fill_2 FILLER_8_965 ();
 sg13g2_fill_2 FILLER_8_990 ();
 sg13g2_fill_1 FILLER_8_992 ();
 sg13g2_fill_1 FILLER_8_1054 ();
 sg13g2_fill_2 FILLER_8_1097 ();
 sg13g2_fill_1 FILLER_8_1099 ();
 sg13g2_fill_1 FILLER_8_1109 ();
 sg13g2_fill_2 FILLER_8_1114 ();
 sg13g2_fill_2 FILLER_8_1146 ();
 sg13g2_fill_1 FILLER_8_1148 ();
 sg13g2_fill_2 FILLER_8_1170 ();
 sg13g2_fill_1 FILLER_8_1172 ();
 sg13g2_fill_2 FILLER_8_1177 ();
 sg13g2_fill_1 FILLER_8_1281 ();
 sg13g2_fill_1 FILLER_8_1301 ();
 sg13g2_fill_2 FILLER_8_1312 ();
 sg13g2_fill_2 FILLER_8_1337 ();
 sg13g2_fill_2 FILLER_8_1358 ();
 sg13g2_fill_2 FILLER_8_1386 ();
 sg13g2_fill_1 FILLER_8_1388 ();
 sg13g2_fill_2 FILLER_8_1437 ();
 sg13g2_fill_2 FILLER_8_1454 ();
 sg13g2_fill_2 FILLER_8_1465 ();
 sg13g2_fill_1 FILLER_8_1467 ();
 sg13g2_decap_8 FILLER_8_1520 ();
 sg13g2_decap_8 FILLER_8_1527 ();
 sg13g2_decap_8 FILLER_8_1534 ();
 sg13g2_decap_8 FILLER_8_1541 ();
 sg13g2_decap_8 FILLER_8_1548 ();
 sg13g2_decap_8 FILLER_8_1555 ();
 sg13g2_decap_8 FILLER_8_1562 ();
 sg13g2_decap_8 FILLER_8_1569 ();
 sg13g2_decap_8 FILLER_8_1576 ();
 sg13g2_decap_8 FILLER_8_1583 ();
 sg13g2_decap_8 FILLER_8_1590 ();
 sg13g2_decap_8 FILLER_8_1597 ();
 sg13g2_decap_8 FILLER_8_1604 ();
 sg13g2_decap_8 FILLER_8_1611 ();
 sg13g2_decap_8 FILLER_8_1618 ();
 sg13g2_decap_8 FILLER_8_1625 ();
 sg13g2_decap_8 FILLER_8_1632 ();
 sg13g2_decap_8 FILLER_8_1639 ();
 sg13g2_decap_8 FILLER_8_1646 ();
 sg13g2_decap_8 FILLER_8_1653 ();
 sg13g2_decap_8 FILLER_8_1660 ();
 sg13g2_decap_8 FILLER_8_1667 ();
 sg13g2_decap_8 FILLER_8_1674 ();
 sg13g2_decap_8 FILLER_8_1681 ();
 sg13g2_decap_8 FILLER_8_1688 ();
 sg13g2_decap_8 FILLER_8_1695 ();
 sg13g2_decap_8 FILLER_8_1702 ();
 sg13g2_decap_8 FILLER_8_1709 ();
 sg13g2_decap_8 FILLER_8_1716 ();
 sg13g2_decap_8 FILLER_8_1723 ();
 sg13g2_decap_8 FILLER_8_1730 ();
 sg13g2_decap_8 FILLER_8_1737 ();
 sg13g2_decap_8 FILLER_8_1744 ();
 sg13g2_decap_8 FILLER_8_1751 ();
 sg13g2_decap_8 FILLER_8_1758 ();
 sg13g2_fill_2 FILLER_8_1765 ();
 sg13g2_fill_1 FILLER_8_1767 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_fill_1 FILLER_9_65 ();
 sg13g2_fill_2 FILLER_9_110 ();
 sg13g2_fill_2 FILLER_9_188 ();
 sg13g2_fill_2 FILLER_9_196 ();
 sg13g2_fill_2 FILLER_9_224 ();
 sg13g2_fill_1 FILLER_9_234 ();
 sg13g2_fill_1 FILLER_9_284 ();
 sg13g2_fill_1 FILLER_9_307 ();
 sg13g2_fill_2 FILLER_9_335 ();
 sg13g2_fill_1 FILLER_9_337 ();
 sg13g2_fill_2 FILLER_9_405 ();
 sg13g2_fill_2 FILLER_9_439 ();
 sg13g2_fill_2 FILLER_9_486 ();
 sg13g2_fill_1 FILLER_9_508 ();
 sg13g2_fill_1 FILLER_9_534 ();
 sg13g2_fill_2 FILLER_9_544 ();
 sg13g2_fill_1 FILLER_9_602 ();
 sg13g2_fill_2 FILLER_9_634 ();
 sg13g2_fill_1 FILLER_9_646 ();
 sg13g2_fill_1 FILLER_9_656 ();
 sg13g2_fill_1 FILLER_9_662 ();
 sg13g2_fill_2 FILLER_9_671 ();
 sg13g2_fill_2 FILLER_9_678 ();
 sg13g2_fill_1 FILLER_9_729 ();
 sg13g2_fill_1 FILLER_9_735 ();
 sg13g2_fill_2 FILLER_9_769 ();
 sg13g2_fill_1 FILLER_9_771 ();
 sg13g2_fill_1 FILLER_9_796 ();
 sg13g2_decap_4 FILLER_9_888 ();
 sg13g2_fill_2 FILLER_9_892 ();
 sg13g2_fill_2 FILLER_9_926 ();
 sg13g2_fill_1 FILLER_9_928 ();
 sg13g2_fill_1 FILLER_9_960 ();
 sg13g2_decap_8 FILLER_9_972 ();
 sg13g2_fill_2 FILLER_9_1012 ();
 sg13g2_fill_2 FILLER_9_1026 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_fill_2 FILLER_9_1060 ();
 sg13g2_fill_1 FILLER_9_1062 ();
 sg13g2_fill_1 FILLER_9_1137 ();
 sg13g2_fill_2 FILLER_9_1145 ();
 sg13g2_fill_2 FILLER_9_1157 ();
 sg13g2_fill_2 FILLER_9_1226 ();
 sg13g2_fill_1 FILLER_9_1274 ();
 sg13g2_fill_2 FILLER_9_1315 ();
 sg13g2_fill_1 FILLER_9_1317 ();
 sg13g2_fill_1 FILLER_9_1344 ();
 sg13g2_fill_2 FILLER_9_1362 ();
 sg13g2_fill_2 FILLER_9_1439 ();
 sg13g2_fill_1 FILLER_9_1482 ();
 sg13g2_fill_2 FILLER_9_1501 ();
 sg13g2_fill_1 FILLER_9_1503 ();
 sg13g2_decap_8 FILLER_9_1529 ();
 sg13g2_decap_8 FILLER_9_1536 ();
 sg13g2_decap_8 FILLER_9_1543 ();
 sg13g2_decap_8 FILLER_9_1550 ();
 sg13g2_decap_8 FILLER_9_1557 ();
 sg13g2_decap_8 FILLER_9_1564 ();
 sg13g2_decap_8 FILLER_9_1571 ();
 sg13g2_decap_8 FILLER_9_1578 ();
 sg13g2_decap_8 FILLER_9_1585 ();
 sg13g2_decap_8 FILLER_9_1592 ();
 sg13g2_decap_8 FILLER_9_1599 ();
 sg13g2_decap_8 FILLER_9_1606 ();
 sg13g2_decap_8 FILLER_9_1613 ();
 sg13g2_decap_8 FILLER_9_1620 ();
 sg13g2_decap_8 FILLER_9_1627 ();
 sg13g2_decap_8 FILLER_9_1634 ();
 sg13g2_decap_8 FILLER_9_1641 ();
 sg13g2_decap_8 FILLER_9_1648 ();
 sg13g2_decap_8 FILLER_9_1655 ();
 sg13g2_decap_8 FILLER_9_1662 ();
 sg13g2_decap_8 FILLER_9_1669 ();
 sg13g2_decap_8 FILLER_9_1676 ();
 sg13g2_decap_8 FILLER_9_1683 ();
 sg13g2_decap_8 FILLER_9_1690 ();
 sg13g2_decap_8 FILLER_9_1697 ();
 sg13g2_decap_8 FILLER_9_1704 ();
 sg13g2_decap_8 FILLER_9_1711 ();
 sg13g2_decap_8 FILLER_9_1718 ();
 sg13g2_decap_8 FILLER_9_1725 ();
 sg13g2_decap_8 FILLER_9_1732 ();
 sg13g2_decap_8 FILLER_9_1739 ();
 sg13g2_decap_8 FILLER_9_1746 ();
 sg13g2_decap_8 FILLER_9_1753 ();
 sg13g2_decap_8 FILLER_9_1760 ();
 sg13g2_fill_1 FILLER_9_1767 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_fill_2 FILLER_10_53 ();
 sg13g2_fill_2 FILLER_10_75 ();
 sg13g2_fill_1 FILLER_10_142 ();
 sg13g2_fill_2 FILLER_10_153 ();
 sg13g2_fill_1 FILLER_10_169 ();
 sg13g2_fill_2 FILLER_10_202 ();
 sg13g2_fill_2 FILLER_10_367 ();
 sg13g2_fill_1 FILLER_10_369 ();
 sg13g2_fill_1 FILLER_10_375 ();
 sg13g2_fill_1 FILLER_10_394 ();
 sg13g2_fill_2 FILLER_10_442 ();
 sg13g2_fill_2 FILLER_10_478 ();
 sg13g2_fill_2 FILLER_10_499 ();
 sg13g2_fill_1 FILLER_10_579 ();
 sg13g2_fill_2 FILLER_10_589 ();
 sg13g2_fill_1 FILLER_10_595 ();
 sg13g2_fill_2 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_799 ();
 sg13g2_decap_4 FILLER_10_806 ();
 sg13g2_decap_4 FILLER_10_814 ();
 sg13g2_fill_1 FILLER_10_818 ();
 sg13g2_decap_4 FILLER_10_824 ();
 sg13g2_fill_2 FILLER_10_828 ();
 sg13g2_fill_2 FILLER_10_848 ();
 sg13g2_fill_1 FILLER_10_850 ();
 sg13g2_fill_1 FILLER_10_914 ();
 sg13g2_fill_1 FILLER_10_972 ();
 sg13g2_fill_1 FILLER_10_982 ();
 sg13g2_fill_1 FILLER_10_995 ();
 sg13g2_fill_2 FILLER_10_1052 ();
 sg13g2_fill_1 FILLER_10_1054 ();
 sg13g2_fill_1 FILLER_10_1078 ();
 sg13g2_fill_2 FILLER_10_1089 ();
 sg13g2_fill_1 FILLER_10_1091 ();
 sg13g2_fill_2 FILLER_10_1112 ();
 sg13g2_fill_1 FILLER_10_1122 ();
 sg13g2_fill_2 FILLER_10_1154 ();
 sg13g2_fill_2 FILLER_10_1168 ();
 sg13g2_fill_1 FILLER_10_1179 ();
 sg13g2_fill_1 FILLER_10_1240 ();
 sg13g2_fill_2 FILLER_10_1295 ();
 sg13g2_fill_2 FILLER_10_1310 ();
 sg13g2_fill_2 FILLER_10_1360 ();
 sg13g2_fill_1 FILLER_10_1397 ();
 sg13g2_fill_1 FILLER_10_1456 ();
 sg13g2_fill_1 FILLER_10_1476 ();
 sg13g2_fill_1 FILLER_10_1488 ();
 sg13g2_decap_8 FILLER_10_1528 ();
 sg13g2_decap_8 FILLER_10_1535 ();
 sg13g2_decap_8 FILLER_10_1542 ();
 sg13g2_decap_8 FILLER_10_1549 ();
 sg13g2_decap_8 FILLER_10_1556 ();
 sg13g2_decap_8 FILLER_10_1563 ();
 sg13g2_decap_8 FILLER_10_1570 ();
 sg13g2_decap_8 FILLER_10_1577 ();
 sg13g2_decap_8 FILLER_10_1584 ();
 sg13g2_decap_8 FILLER_10_1591 ();
 sg13g2_decap_8 FILLER_10_1598 ();
 sg13g2_decap_8 FILLER_10_1605 ();
 sg13g2_decap_8 FILLER_10_1612 ();
 sg13g2_decap_8 FILLER_10_1619 ();
 sg13g2_decap_8 FILLER_10_1626 ();
 sg13g2_decap_8 FILLER_10_1633 ();
 sg13g2_decap_8 FILLER_10_1640 ();
 sg13g2_decap_8 FILLER_10_1647 ();
 sg13g2_decap_8 FILLER_10_1654 ();
 sg13g2_decap_8 FILLER_10_1661 ();
 sg13g2_decap_8 FILLER_10_1668 ();
 sg13g2_decap_8 FILLER_10_1675 ();
 sg13g2_decap_8 FILLER_10_1682 ();
 sg13g2_decap_8 FILLER_10_1689 ();
 sg13g2_decap_8 FILLER_10_1696 ();
 sg13g2_decap_8 FILLER_10_1703 ();
 sg13g2_decap_8 FILLER_10_1710 ();
 sg13g2_decap_8 FILLER_10_1717 ();
 sg13g2_decap_8 FILLER_10_1724 ();
 sg13g2_decap_8 FILLER_10_1731 ();
 sg13g2_decap_8 FILLER_10_1738 ();
 sg13g2_decap_8 FILLER_10_1745 ();
 sg13g2_decap_8 FILLER_10_1752 ();
 sg13g2_decap_8 FILLER_10_1759 ();
 sg13g2_fill_2 FILLER_10_1766 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_fill_1 FILLER_11_52 ();
 sg13g2_fill_2 FILLER_11_79 ();
 sg13g2_fill_1 FILLER_11_81 ();
 sg13g2_fill_1 FILLER_11_102 ();
 sg13g2_fill_1 FILLER_11_118 ();
 sg13g2_fill_2 FILLER_11_128 ();
 sg13g2_fill_1 FILLER_11_130 ();
 sg13g2_fill_2 FILLER_11_137 ();
 sg13g2_fill_1 FILLER_11_139 ();
 sg13g2_fill_2 FILLER_11_175 ();
 sg13g2_fill_2 FILLER_11_208 ();
 sg13g2_fill_2 FILLER_11_255 ();
 sg13g2_fill_1 FILLER_11_283 ();
 sg13g2_fill_2 FILLER_11_289 ();
 sg13g2_fill_1 FILLER_11_291 ();
 sg13g2_fill_2 FILLER_11_310 ();
 sg13g2_fill_2 FILLER_11_317 ();
 sg13g2_fill_1 FILLER_11_319 ();
 sg13g2_fill_2 FILLER_11_372 ();
 sg13g2_fill_1 FILLER_11_374 ();
 sg13g2_fill_1 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_464 ();
 sg13g2_fill_1 FILLER_11_512 ();
 sg13g2_fill_1 FILLER_11_517 ();
 sg13g2_fill_1 FILLER_11_551 ();
 sg13g2_fill_2 FILLER_11_572 ();
 sg13g2_fill_1 FILLER_11_574 ();
 sg13g2_fill_2 FILLER_11_610 ();
 sg13g2_fill_1 FILLER_11_636 ();
 sg13g2_fill_1 FILLER_11_646 ();
 sg13g2_fill_2 FILLER_11_669 ();
 sg13g2_fill_2 FILLER_11_712 ();
 sg13g2_fill_1 FILLER_11_731 ();
 sg13g2_fill_1 FILLER_11_763 ();
 sg13g2_fill_2 FILLER_11_778 ();
 sg13g2_decap_4 FILLER_11_806 ();
 sg13g2_fill_2 FILLER_11_844 ();
 sg13g2_fill_1 FILLER_11_918 ();
 sg13g2_fill_2 FILLER_11_933 ();
 sg13g2_fill_1 FILLER_11_940 ();
 sg13g2_fill_2 FILLER_11_1021 ();
 sg13g2_fill_1 FILLER_11_1034 ();
 sg13g2_fill_2 FILLER_11_1049 ();
 sg13g2_fill_1 FILLER_11_1051 ();
 sg13g2_fill_2 FILLER_11_1106 ();
 sg13g2_fill_1 FILLER_11_1108 ();
 sg13g2_fill_2 FILLER_11_1138 ();
 sg13g2_fill_2 FILLER_11_1153 ();
 sg13g2_fill_2 FILLER_11_1160 ();
 sg13g2_fill_2 FILLER_11_1190 ();
 sg13g2_fill_2 FILLER_11_1222 ();
 sg13g2_fill_1 FILLER_11_1256 ();
 sg13g2_fill_2 FILLER_11_1374 ();
 sg13g2_fill_2 FILLER_11_1389 ();
 sg13g2_fill_2 FILLER_11_1448 ();
 sg13g2_fill_1 FILLER_11_1473 ();
 sg13g2_fill_2 FILLER_11_1500 ();
 sg13g2_fill_1 FILLER_11_1502 ();
 sg13g2_decap_8 FILLER_11_1538 ();
 sg13g2_decap_8 FILLER_11_1545 ();
 sg13g2_decap_8 FILLER_11_1552 ();
 sg13g2_decap_8 FILLER_11_1559 ();
 sg13g2_decap_8 FILLER_11_1566 ();
 sg13g2_decap_8 FILLER_11_1573 ();
 sg13g2_decap_8 FILLER_11_1580 ();
 sg13g2_decap_8 FILLER_11_1587 ();
 sg13g2_decap_8 FILLER_11_1594 ();
 sg13g2_decap_8 FILLER_11_1601 ();
 sg13g2_decap_8 FILLER_11_1608 ();
 sg13g2_decap_8 FILLER_11_1615 ();
 sg13g2_decap_8 FILLER_11_1622 ();
 sg13g2_decap_8 FILLER_11_1629 ();
 sg13g2_decap_8 FILLER_11_1636 ();
 sg13g2_decap_8 FILLER_11_1643 ();
 sg13g2_decap_8 FILLER_11_1650 ();
 sg13g2_decap_8 FILLER_11_1657 ();
 sg13g2_decap_8 FILLER_11_1664 ();
 sg13g2_decap_8 FILLER_11_1671 ();
 sg13g2_decap_8 FILLER_11_1678 ();
 sg13g2_decap_8 FILLER_11_1685 ();
 sg13g2_decap_8 FILLER_11_1692 ();
 sg13g2_decap_8 FILLER_11_1699 ();
 sg13g2_decap_8 FILLER_11_1706 ();
 sg13g2_decap_8 FILLER_11_1713 ();
 sg13g2_decap_8 FILLER_11_1720 ();
 sg13g2_decap_8 FILLER_11_1727 ();
 sg13g2_decap_8 FILLER_11_1734 ();
 sg13g2_decap_8 FILLER_11_1741 ();
 sg13g2_decap_8 FILLER_11_1748 ();
 sg13g2_decap_8 FILLER_11_1755 ();
 sg13g2_decap_4 FILLER_11_1762 ();
 sg13g2_fill_2 FILLER_11_1766 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_69 ();
 sg13g2_fill_1 FILLER_12_71 ();
 sg13g2_fill_1 FILLER_12_194 ();
 sg13g2_fill_1 FILLER_12_254 ();
 sg13g2_fill_2 FILLER_12_263 ();
 sg13g2_fill_1 FILLER_12_273 ();
 sg13g2_fill_1 FILLER_12_309 ();
 sg13g2_fill_2 FILLER_12_344 ();
 sg13g2_fill_2 FILLER_12_376 ();
 sg13g2_fill_2 FILLER_12_391 ();
 sg13g2_fill_2 FILLER_12_432 ();
 sg13g2_fill_2 FILLER_12_495 ();
 sg13g2_fill_2 FILLER_12_511 ();
 sg13g2_fill_1 FILLER_12_548 ();
 sg13g2_fill_2 FILLER_12_583 ();
 sg13g2_fill_1 FILLER_12_585 ();
 sg13g2_fill_1 FILLER_12_590 ();
 sg13g2_fill_1 FILLER_12_596 ();
 sg13g2_fill_2 FILLER_12_602 ();
 sg13g2_fill_1 FILLER_12_604 ();
 sg13g2_fill_2 FILLER_12_611 ();
 sg13g2_fill_1 FILLER_12_613 ();
 sg13g2_fill_2 FILLER_12_714 ();
 sg13g2_fill_2 FILLER_12_725 ();
 sg13g2_fill_1 FILLER_12_727 ();
 sg13g2_fill_1 FILLER_12_760 ();
 sg13g2_fill_2 FILLER_12_795 ();
 sg13g2_decap_8 FILLER_12_814 ();
 sg13g2_fill_1 FILLER_12_845 ();
 sg13g2_decap_4 FILLER_12_884 ();
 sg13g2_fill_2 FILLER_12_928 ();
 sg13g2_fill_1 FILLER_12_930 ();
 sg13g2_fill_2 FILLER_12_957 ();
 sg13g2_fill_2 FILLER_12_980 ();
 sg13g2_fill_1 FILLER_12_982 ();
 sg13g2_fill_1 FILLER_12_1015 ();
 sg13g2_fill_2 FILLER_12_1022 ();
 sg13g2_fill_1 FILLER_12_1024 ();
 sg13g2_fill_1 FILLER_12_1055 ();
 sg13g2_fill_1 FILLER_12_1065 ();
 sg13g2_fill_2 FILLER_12_1075 ();
 sg13g2_fill_1 FILLER_12_1191 ();
 sg13g2_fill_1 FILLER_12_1231 ();
 sg13g2_fill_2 FILLER_12_1237 ();
 sg13g2_fill_2 FILLER_12_1265 ();
 sg13g2_fill_1 FILLER_12_1267 ();
 sg13g2_fill_1 FILLER_12_1300 ();
 sg13g2_fill_1 FILLER_12_1321 ();
 sg13g2_fill_1 FILLER_12_1334 ();
 sg13g2_fill_1 FILLER_12_1406 ();
 sg13g2_fill_2 FILLER_12_1430 ();
 sg13g2_fill_1 FILLER_12_1432 ();
 sg13g2_fill_1 FILLER_12_1506 ();
 sg13g2_decap_8 FILLER_12_1561 ();
 sg13g2_decap_8 FILLER_12_1568 ();
 sg13g2_decap_8 FILLER_12_1575 ();
 sg13g2_decap_8 FILLER_12_1582 ();
 sg13g2_decap_8 FILLER_12_1589 ();
 sg13g2_decap_8 FILLER_12_1596 ();
 sg13g2_decap_8 FILLER_12_1603 ();
 sg13g2_decap_8 FILLER_12_1610 ();
 sg13g2_decap_8 FILLER_12_1617 ();
 sg13g2_decap_8 FILLER_12_1624 ();
 sg13g2_decap_8 FILLER_12_1631 ();
 sg13g2_decap_8 FILLER_12_1638 ();
 sg13g2_decap_8 FILLER_12_1645 ();
 sg13g2_decap_8 FILLER_12_1652 ();
 sg13g2_decap_8 FILLER_12_1659 ();
 sg13g2_decap_8 FILLER_12_1666 ();
 sg13g2_decap_8 FILLER_12_1673 ();
 sg13g2_decap_8 FILLER_12_1680 ();
 sg13g2_decap_8 FILLER_12_1687 ();
 sg13g2_decap_8 FILLER_12_1694 ();
 sg13g2_decap_8 FILLER_12_1701 ();
 sg13g2_decap_8 FILLER_12_1708 ();
 sg13g2_decap_8 FILLER_12_1715 ();
 sg13g2_decap_8 FILLER_12_1722 ();
 sg13g2_decap_8 FILLER_12_1729 ();
 sg13g2_decap_8 FILLER_12_1736 ();
 sg13g2_decap_8 FILLER_12_1743 ();
 sg13g2_decap_8 FILLER_12_1750 ();
 sg13g2_decap_8 FILLER_12_1757 ();
 sg13g2_decap_4 FILLER_12_1764 ();
 sg13g2_fill_2 FILLER_13_26 ();
 sg13g2_fill_1 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_64 ();
 sg13g2_fill_2 FILLER_13_92 ();
 sg13g2_fill_1 FILLER_13_94 ();
 sg13g2_fill_2 FILLER_13_101 ();
 sg13g2_fill_2 FILLER_13_134 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_fill_1 FILLER_13_163 ();
 sg13g2_fill_1 FILLER_13_181 ();
 sg13g2_fill_1 FILLER_13_200 ();
 sg13g2_fill_1 FILLER_13_209 ();
 sg13g2_fill_1 FILLER_13_218 ();
 sg13g2_fill_2 FILLER_13_233 ();
 sg13g2_fill_2 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_fill_2 FILLER_13_300 ();
 sg13g2_fill_1 FILLER_13_302 ();
 sg13g2_fill_2 FILLER_13_317 ();
 sg13g2_fill_1 FILLER_13_319 ();
 sg13g2_fill_2 FILLER_13_334 ();
 sg13g2_fill_1 FILLER_13_377 ();
 sg13g2_fill_2 FILLER_13_410 ();
 sg13g2_fill_2 FILLER_13_446 ();
 sg13g2_fill_2 FILLER_13_481 ();
 sg13g2_fill_1 FILLER_13_540 ();
 sg13g2_fill_1 FILLER_13_550 ();
 sg13g2_fill_2 FILLER_13_566 ();
 sg13g2_fill_2 FILLER_13_633 ();
 sg13g2_fill_2 FILLER_13_648 ();
 sg13g2_fill_2 FILLER_13_654 ();
 sg13g2_fill_1 FILLER_13_656 ();
 sg13g2_fill_1 FILLER_13_700 ();
 sg13g2_fill_2 FILLER_13_731 ();
 sg13g2_fill_2 FILLER_13_759 ();
 sg13g2_fill_1 FILLER_13_779 ();
 sg13g2_fill_1 FILLER_13_785 ();
 sg13g2_fill_2 FILLER_13_812 ();
 sg13g2_decap_4 FILLER_13_840 ();
 sg13g2_fill_2 FILLER_13_849 ();
 sg13g2_decap_4 FILLER_13_859 ();
 sg13g2_decap_8 FILLER_13_890 ();
 sg13g2_fill_1 FILLER_13_897 ();
 sg13g2_fill_1 FILLER_13_906 ();
 sg13g2_fill_1 FILLER_13_939 ();
 sg13g2_fill_1 FILLER_13_992 ();
 sg13g2_fill_2 FILLER_13_1071 ();
 sg13g2_fill_1 FILLER_13_1073 ();
 sg13g2_fill_1 FILLER_13_1111 ();
 sg13g2_fill_2 FILLER_13_1190 ();
 sg13g2_fill_2 FILLER_13_1202 ();
 sg13g2_fill_1 FILLER_13_1204 ();
 sg13g2_fill_2 FILLER_13_1240 ();
 sg13g2_fill_2 FILLER_13_1277 ();
 sg13g2_fill_1 FILLER_13_1288 ();
 sg13g2_fill_2 FILLER_13_1326 ();
 sg13g2_fill_1 FILLER_13_1328 ();
 sg13g2_fill_2 FILLER_13_1375 ();
 sg13g2_fill_1 FILLER_13_1391 ();
 sg13g2_fill_2 FILLER_13_1400 ();
 sg13g2_fill_2 FILLER_13_1444 ();
 sg13g2_decap_8 FILLER_13_1540 ();
 sg13g2_decap_8 FILLER_13_1547 ();
 sg13g2_decap_8 FILLER_13_1554 ();
 sg13g2_decap_8 FILLER_13_1561 ();
 sg13g2_decap_8 FILLER_13_1568 ();
 sg13g2_decap_8 FILLER_13_1575 ();
 sg13g2_decap_8 FILLER_13_1582 ();
 sg13g2_decap_8 FILLER_13_1589 ();
 sg13g2_decap_8 FILLER_13_1596 ();
 sg13g2_decap_8 FILLER_13_1603 ();
 sg13g2_decap_8 FILLER_13_1610 ();
 sg13g2_decap_8 FILLER_13_1617 ();
 sg13g2_decap_8 FILLER_13_1624 ();
 sg13g2_decap_8 FILLER_13_1631 ();
 sg13g2_decap_8 FILLER_13_1638 ();
 sg13g2_decap_8 FILLER_13_1645 ();
 sg13g2_decap_8 FILLER_13_1652 ();
 sg13g2_decap_8 FILLER_13_1659 ();
 sg13g2_decap_8 FILLER_13_1666 ();
 sg13g2_decap_8 FILLER_13_1673 ();
 sg13g2_decap_8 FILLER_13_1680 ();
 sg13g2_decap_8 FILLER_13_1687 ();
 sg13g2_decap_8 FILLER_13_1694 ();
 sg13g2_decap_8 FILLER_13_1701 ();
 sg13g2_decap_8 FILLER_13_1708 ();
 sg13g2_decap_8 FILLER_13_1715 ();
 sg13g2_decap_8 FILLER_13_1722 ();
 sg13g2_decap_8 FILLER_13_1729 ();
 sg13g2_decap_8 FILLER_13_1736 ();
 sg13g2_decap_8 FILLER_13_1743 ();
 sg13g2_decap_8 FILLER_13_1750 ();
 sg13g2_decap_8 FILLER_13_1757 ();
 sg13g2_decap_4 FILLER_13_1764 ();
 sg13g2_fill_2 FILLER_14_26 ();
 sg13g2_fill_1 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_34 ();
 sg13g2_fill_1 FILLER_14_36 ();
 sg13g2_fill_1 FILLER_14_67 ();
 sg13g2_fill_1 FILLER_14_99 ();
 sg13g2_fill_2 FILLER_14_106 ();
 sg13g2_fill_1 FILLER_14_108 ();
 sg13g2_fill_2 FILLER_14_123 ();
 sg13g2_fill_1 FILLER_14_133 ();
 sg13g2_fill_2 FILLER_14_139 ();
 sg13g2_fill_1 FILLER_14_141 ();
 sg13g2_fill_1 FILLER_14_218 ();
 sg13g2_fill_2 FILLER_14_258 ();
 sg13g2_fill_2 FILLER_14_301 ();
 sg13g2_fill_1 FILLER_14_303 ();
 sg13g2_fill_1 FILLER_14_312 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_fill_2 FILLER_14_354 ();
 sg13g2_fill_1 FILLER_14_356 ();
 sg13g2_fill_1 FILLER_14_389 ();
 sg13g2_fill_1 FILLER_14_431 ();
 sg13g2_fill_2 FILLER_14_463 ();
 sg13g2_fill_2 FILLER_14_471 ();
 sg13g2_fill_2 FILLER_14_497 ();
 sg13g2_fill_1 FILLER_14_504 ();
 sg13g2_fill_2 FILLER_14_514 ();
 sg13g2_fill_1 FILLER_14_516 ();
 sg13g2_fill_2 FILLER_14_563 ();
 sg13g2_decap_4 FILLER_14_600 ();
 sg13g2_fill_2 FILLER_14_635 ();
 sg13g2_fill_1 FILLER_14_667 ();
 sg13g2_fill_1 FILLER_14_673 ();
 sg13g2_fill_1 FILLER_14_689 ();
 sg13g2_fill_2 FILLER_14_715 ();
 sg13g2_fill_2 FILLER_14_767 ();
 sg13g2_decap_8 FILLER_14_801 ();
 sg13g2_decap_4 FILLER_14_808 ();
 sg13g2_fill_1 FILLER_14_812 ();
 sg13g2_decap_4 FILLER_14_880 ();
 sg13g2_fill_1 FILLER_14_915 ();
 sg13g2_fill_2 FILLER_14_925 ();
 sg13g2_fill_1 FILLER_14_927 ();
 sg13g2_fill_1 FILLER_14_937 ();
 sg13g2_fill_1 FILLER_14_969 ();
 sg13g2_fill_2 FILLER_14_989 ();
 sg13g2_fill_1 FILLER_14_991 ();
 sg13g2_fill_1 FILLER_14_996 ();
 sg13g2_fill_2 FILLER_14_1051 ();
 sg13g2_fill_2 FILLER_14_1110 ();
 sg13g2_fill_1 FILLER_14_1112 ();
 sg13g2_fill_2 FILLER_14_1139 ();
 sg13g2_fill_1 FILLER_14_1141 ();
 sg13g2_fill_2 FILLER_14_1162 ();
 sg13g2_fill_1 FILLER_14_1164 ();
 sg13g2_fill_2 FILLER_14_1196 ();
 sg13g2_fill_1 FILLER_14_1198 ();
 sg13g2_fill_2 FILLER_14_1226 ();
 sg13g2_fill_2 FILLER_14_1262 ();
 sg13g2_fill_1 FILLER_14_1277 ();
 sg13g2_fill_2 FILLER_14_1283 ();
 sg13g2_fill_1 FILLER_14_1285 ();
 sg13g2_fill_2 FILLER_14_1345 ();
 sg13g2_fill_2 FILLER_14_1356 ();
 sg13g2_fill_1 FILLER_14_1358 ();
 sg13g2_fill_2 FILLER_14_1371 ();
 sg13g2_fill_2 FILLER_14_1415 ();
 sg13g2_fill_1 FILLER_14_1468 ();
 sg13g2_fill_1 FILLER_14_1495 ();
 sg13g2_decap_8 FILLER_14_1554 ();
 sg13g2_decap_8 FILLER_14_1561 ();
 sg13g2_decap_8 FILLER_14_1568 ();
 sg13g2_decap_8 FILLER_14_1575 ();
 sg13g2_decap_8 FILLER_14_1582 ();
 sg13g2_decap_8 FILLER_14_1589 ();
 sg13g2_decap_8 FILLER_14_1596 ();
 sg13g2_decap_8 FILLER_14_1603 ();
 sg13g2_decap_8 FILLER_14_1610 ();
 sg13g2_decap_8 FILLER_14_1617 ();
 sg13g2_decap_8 FILLER_14_1624 ();
 sg13g2_decap_8 FILLER_14_1631 ();
 sg13g2_decap_8 FILLER_14_1638 ();
 sg13g2_decap_8 FILLER_14_1645 ();
 sg13g2_decap_8 FILLER_14_1652 ();
 sg13g2_decap_8 FILLER_14_1659 ();
 sg13g2_decap_8 FILLER_14_1666 ();
 sg13g2_decap_8 FILLER_14_1673 ();
 sg13g2_decap_8 FILLER_14_1680 ();
 sg13g2_decap_8 FILLER_14_1687 ();
 sg13g2_decap_8 FILLER_14_1694 ();
 sg13g2_decap_8 FILLER_14_1701 ();
 sg13g2_decap_8 FILLER_14_1708 ();
 sg13g2_decap_8 FILLER_14_1715 ();
 sg13g2_decap_8 FILLER_14_1722 ();
 sg13g2_decap_8 FILLER_14_1729 ();
 sg13g2_decap_8 FILLER_14_1736 ();
 sg13g2_decap_8 FILLER_14_1743 ();
 sg13g2_decap_8 FILLER_14_1750 ();
 sg13g2_decap_8 FILLER_14_1757 ();
 sg13g2_decap_4 FILLER_14_1764 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_19 ();
 sg13g2_fill_2 FILLER_15_56 ();
 sg13g2_fill_2 FILLER_15_117 ();
 sg13g2_fill_1 FILLER_15_119 ();
 sg13g2_fill_2 FILLER_15_151 ();
 sg13g2_fill_1 FILLER_15_153 ();
 sg13g2_fill_1 FILLER_15_222 ();
 sg13g2_fill_1 FILLER_15_247 ();
 sg13g2_fill_2 FILLER_15_258 ();
 sg13g2_fill_2 FILLER_15_265 ();
 sg13g2_fill_1 FILLER_15_299 ();
 sg13g2_fill_2 FILLER_15_309 ();
 sg13g2_fill_1 FILLER_15_311 ();
 sg13g2_fill_2 FILLER_15_325 ();
 sg13g2_fill_1 FILLER_15_327 ();
 sg13g2_fill_2 FILLER_15_332 ();
 sg13g2_fill_1 FILLER_15_334 ();
 sg13g2_fill_2 FILLER_15_397 ();
 sg13g2_fill_1 FILLER_15_454 ();
 sg13g2_fill_2 FILLER_15_520 ();
 sg13g2_fill_2 FILLER_15_528 ();
 sg13g2_fill_2 FILLER_15_558 ();
 sg13g2_fill_1 FILLER_15_560 ();
 sg13g2_fill_1 FILLER_15_575 ();
 sg13g2_fill_1 FILLER_15_717 ();
 sg13g2_fill_2 FILLER_15_850 ();
 sg13g2_decap_4 FILLER_15_883 ();
 sg13g2_fill_2 FILLER_15_887 ();
 sg13g2_fill_1 FILLER_15_912 ();
 sg13g2_fill_2 FILLER_15_918 ();
 sg13g2_decap_4 FILLER_15_955 ();
 sg13g2_fill_2 FILLER_15_998 ();
 sg13g2_fill_1 FILLER_15_1000 ();
 sg13g2_fill_2 FILLER_15_1063 ();
 sg13g2_fill_2 FILLER_15_1071 ();
 sg13g2_fill_1 FILLER_15_1073 ();
 sg13g2_fill_2 FILLER_15_1089 ();
 sg13g2_fill_2 FILLER_15_1100 ();
 sg13g2_fill_1 FILLER_15_1134 ();
 sg13g2_fill_2 FILLER_15_1171 ();
 sg13g2_fill_2 FILLER_15_1203 ();
 sg13g2_fill_1 FILLER_15_1205 ();
 sg13g2_fill_1 FILLER_15_1236 ();
 sg13g2_fill_2 FILLER_15_1250 ();
 sg13g2_fill_2 FILLER_15_1266 ();
 sg13g2_fill_1 FILLER_15_1268 ();
 sg13g2_fill_1 FILLER_15_1323 ();
 sg13g2_fill_1 FILLER_15_1356 ();
 sg13g2_fill_2 FILLER_15_1396 ();
 sg13g2_fill_2 FILLER_15_1419 ();
 sg13g2_fill_2 FILLER_15_1447 ();
 sg13g2_fill_1 FILLER_15_1479 ();
 sg13g2_fill_2 FILLER_15_1499 ();
 sg13g2_fill_1 FILLER_15_1501 ();
 sg13g2_fill_1 FILLER_15_1518 ();
 sg13g2_decap_8 FILLER_15_1552 ();
 sg13g2_decap_8 FILLER_15_1559 ();
 sg13g2_decap_8 FILLER_15_1566 ();
 sg13g2_decap_8 FILLER_15_1573 ();
 sg13g2_decap_8 FILLER_15_1580 ();
 sg13g2_decap_8 FILLER_15_1587 ();
 sg13g2_decap_8 FILLER_15_1594 ();
 sg13g2_decap_8 FILLER_15_1601 ();
 sg13g2_decap_8 FILLER_15_1608 ();
 sg13g2_decap_8 FILLER_15_1615 ();
 sg13g2_decap_8 FILLER_15_1622 ();
 sg13g2_decap_8 FILLER_15_1629 ();
 sg13g2_decap_8 FILLER_15_1636 ();
 sg13g2_decap_8 FILLER_15_1643 ();
 sg13g2_decap_8 FILLER_15_1650 ();
 sg13g2_decap_8 FILLER_15_1657 ();
 sg13g2_decap_8 FILLER_15_1664 ();
 sg13g2_decap_8 FILLER_15_1671 ();
 sg13g2_decap_8 FILLER_15_1678 ();
 sg13g2_decap_8 FILLER_15_1685 ();
 sg13g2_decap_8 FILLER_15_1692 ();
 sg13g2_decap_8 FILLER_15_1699 ();
 sg13g2_decap_8 FILLER_15_1706 ();
 sg13g2_decap_8 FILLER_15_1713 ();
 sg13g2_decap_8 FILLER_15_1720 ();
 sg13g2_decap_8 FILLER_15_1727 ();
 sg13g2_decap_8 FILLER_15_1734 ();
 sg13g2_decap_8 FILLER_15_1741 ();
 sg13g2_decap_8 FILLER_15_1748 ();
 sg13g2_decap_8 FILLER_15_1755 ();
 sg13g2_decap_4 FILLER_15_1762 ();
 sg13g2_fill_2 FILLER_15_1766 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_6 ();
 sg13g2_fill_1 FILLER_16_16 ();
 sg13g2_fill_2 FILLER_16_39 ();
 sg13g2_fill_1 FILLER_16_55 ();
 sg13g2_fill_2 FILLER_16_81 ();
 sg13g2_fill_1 FILLER_16_88 ();
 sg13g2_fill_2 FILLER_16_106 ();
 sg13g2_fill_2 FILLER_16_134 ();
 sg13g2_fill_1 FILLER_16_136 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_fill_2 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_208 ();
 sg13g2_fill_2 FILLER_16_278 ();
 sg13g2_fill_1 FILLER_16_280 ();
 sg13g2_fill_2 FILLER_16_313 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_fill_2 FILLER_16_395 ();
 sg13g2_fill_2 FILLER_16_405 ();
 sg13g2_fill_2 FILLER_16_412 ();
 sg13g2_fill_1 FILLER_16_431 ();
 sg13g2_fill_2 FILLER_16_497 ();
 sg13g2_fill_1 FILLER_16_499 ();
 sg13g2_fill_2 FILLER_16_550 ();
 sg13g2_fill_1 FILLER_16_552 ();
 sg13g2_fill_2 FILLER_16_566 ();
 sg13g2_fill_1 FILLER_16_568 ();
 sg13g2_fill_1 FILLER_16_626 ();
 sg13g2_fill_2 FILLER_16_704 ();
 sg13g2_fill_1 FILLER_16_706 ();
 sg13g2_fill_1 FILLER_16_735 ();
 sg13g2_fill_2 FILLER_16_776 ();
 sg13g2_fill_1 FILLER_16_778 ();
 sg13g2_fill_2 FILLER_16_818 ();
 sg13g2_fill_1 FILLER_16_833 ();
 sg13g2_fill_1 FILLER_16_844 ();
 sg13g2_fill_2 FILLER_16_926 ();
 sg13g2_fill_1 FILLER_16_928 ();
 sg13g2_fill_1 FILLER_16_941 ();
 sg13g2_fill_1 FILLER_16_995 ();
 sg13g2_fill_1 FILLER_16_1039 ();
 sg13g2_fill_2 FILLER_16_1073 ();
 sg13g2_fill_1 FILLER_16_1075 ();
 sg13g2_fill_2 FILLER_16_1102 ();
 sg13g2_fill_2 FILLER_16_1148 ();
 sg13g2_fill_1 FILLER_16_1159 ();
 sg13g2_fill_2 FILLER_16_1200 ();
 sg13g2_fill_1 FILLER_16_1202 ();
 sg13g2_fill_2 FILLER_16_1218 ();
 sg13g2_fill_1 FILLER_16_1220 ();
 sg13g2_fill_1 FILLER_16_1336 ();
 sg13g2_fill_2 FILLER_16_1348 ();
 sg13g2_fill_2 FILLER_16_1360 ();
 sg13g2_fill_1 FILLER_16_1362 ();
 sg13g2_fill_2 FILLER_16_1381 ();
 sg13g2_fill_2 FILLER_16_1435 ();
 sg13g2_fill_1 FILLER_16_1437 ();
 sg13g2_fill_2 FILLER_16_1444 ();
 sg13g2_fill_1 FILLER_16_1446 ();
 sg13g2_fill_2 FILLER_16_1475 ();
 sg13g2_fill_2 FILLER_16_1482 ();
 sg13g2_fill_1 FILLER_16_1484 ();
 sg13g2_decap_8 FILLER_16_1567 ();
 sg13g2_decap_8 FILLER_16_1574 ();
 sg13g2_decap_8 FILLER_16_1581 ();
 sg13g2_decap_8 FILLER_16_1588 ();
 sg13g2_decap_8 FILLER_16_1595 ();
 sg13g2_decap_8 FILLER_16_1602 ();
 sg13g2_decap_8 FILLER_16_1609 ();
 sg13g2_decap_8 FILLER_16_1616 ();
 sg13g2_decap_8 FILLER_16_1623 ();
 sg13g2_decap_8 FILLER_16_1630 ();
 sg13g2_decap_8 FILLER_16_1637 ();
 sg13g2_decap_8 FILLER_16_1644 ();
 sg13g2_decap_8 FILLER_16_1651 ();
 sg13g2_decap_8 FILLER_16_1658 ();
 sg13g2_decap_8 FILLER_16_1665 ();
 sg13g2_decap_8 FILLER_16_1672 ();
 sg13g2_decap_8 FILLER_16_1679 ();
 sg13g2_decap_8 FILLER_16_1686 ();
 sg13g2_decap_8 FILLER_16_1693 ();
 sg13g2_decap_8 FILLER_16_1700 ();
 sg13g2_decap_8 FILLER_16_1707 ();
 sg13g2_decap_8 FILLER_16_1714 ();
 sg13g2_decap_8 FILLER_16_1721 ();
 sg13g2_decap_8 FILLER_16_1728 ();
 sg13g2_decap_8 FILLER_16_1735 ();
 sg13g2_decap_8 FILLER_16_1742 ();
 sg13g2_decap_8 FILLER_16_1749 ();
 sg13g2_decap_8 FILLER_16_1756 ();
 sg13g2_decap_4 FILLER_16_1763 ();
 sg13g2_fill_1 FILLER_16_1767 ();
 sg13g2_fill_1 FILLER_17_40 ();
 sg13g2_fill_1 FILLER_17_54 ();
 sg13g2_fill_2 FILLER_17_72 ();
 sg13g2_fill_2 FILLER_17_118 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_fill_1 FILLER_17_257 ();
 sg13g2_fill_1 FILLER_17_314 ();
 sg13g2_fill_2 FILLER_17_335 ();
 sg13g2_fill_1 FILLER_17_337 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_381 ();
 sg13g2_fill_1 FILLER_17_423 ();
 sg13g2_fill_2 FILLER_17_439 ();
 sg13g2_fill_1 FILLER_17_450 ();
 sg13g2_fill_2 FILLER_17_460 ();
 sg13g2_fill_2 FILLER_17_476 ();
 sg13g2_fill_1 FILLER_17_478 ();
 sg13g2_fill_1 FILLER_17_488 ();
 sg13g2_fill_2 FILLER_17_532 ();
 sg13g2_fill_1 FILLER_17_534 ();
 sg13g2_fill_2 FILLER_17_593 ();
 sg13g2_decap_8 FILLER_17_599 ();
 sg13g2_fill_1 FILLER_17_606 ();
 sg13g2_fill_1 FILLER_17_615 ();
 sg13g2_fill_1 FILLER_17_642 ();
 sg13g2_fill_1 FILLER_17_699 ();
 sg13g2_fill_1 FILLER_17_748 ();
 sg13g2_fill_1 FILLER_17_811 ();
 sg13g2_decap_8 FILLER_17_877 ();
 sg13g2_decap_4 FILLER_17_892 ();
 sg13g2_fill_2 FILLER_17_896 ();
 sg13g2_fill_1 FILLER_17_902 ();
 sg13g2_fill_2 FILLER_17_908 ();
 sg13g2_fill_1 FILLER_17_910 ();
 sg13g2_fill_1 FILLER_17_957 ();
 sg13g2_fill_2 FILLER_17_977 ();
 sg13g2_fill_1 FILLER_17_979 ();
 sg13g2_fill_1 FILLER_17_1007 ();
 sg13g2_fill_2 FILLER_17_1048 ();
 sg13g2_fill_2 FILLER_17_1068 ();
 sg13g2_fill_1 FILLER_17_1117 ();
 sg13g2_fill_2 FILLER_17_1183 ();
 sg13g2_fill_2 FILLER_17_1237 ();
 sg13g2_fill_1 FILLER_17_1239 ();
 sg13g2_fill_2 FILLER_17_1253 ();
 sg13g2_fill_1 FILLER_17_1255 ();
 sg13g2_fill_2 FILLER_17_1305 ();
 sg13g2_fill_1 FILLER_17_1307 ();
 sg13g2_fill_1 FILLER_17_1339 ();
 sg13g2_fill_2 FILLER_17_1459 ();
 sg13g2_fill_1 FILLER_17_1461 ();
 sg13g2_fill_1 FILLER_17_1468 ();
 sg13g2_fill_2 FILLER_17_1502 ();
 sg13g2_fill_1 FILLER_17_1504 ();
 sg13g2_fill_1 FILLER_17_1520 ();
 sg13g2_decap_8 FILLER_17_1559 ();
 sg13g2_decap_8 FILLER_17_1566 ();
 sg13g2_decap_8 FILLER_17_1573 ();
 sg13g2_decap_8 FILLER_17_1580 ();
 sg13g2_decap_8 FILLER_17_1587 ();
 sg13g2_decap_8 FILLER_17_1594 ();
 sg13g2_decap_8 FILLER_17_1601 ();
 sg13g2_decap_8 FILLER_17_1608 ();
 sg13g2_decap_8 FILLER_17_1615 ();
 sg13g2_decap_8 FILLER_17_1622 ();
 sg13g2_decap_8 FILLER_17_1629 ();
 sg13g2_decap_8 FILLER_17_1636 ();
 sg13g2_decap_8 FILLER_17_1643 ();
 sg13g2_decap_8 FILLER_17_1650 ();
 sg13g2_decap_8 FILLER_17_1657 ();
 sg13g2_decap_8 FILLER_17_1664 ();
 sg13g2_decap_8 FILLER_17_1671 ();
 sg13g2_decap_8 FILLER_17_1678 ();
 sg13g2_decap_8 FILLER_17_1685 ();
 sg13g2_decap_8 FILLER_17_1692 ();
 sg13g2_decap_8 FILLER_17_1699 ();
 sg13g2_decap_8 FILLER_17_1706 ();
 sg13g2_decap_8 FILLER_17_1713 ();
 sg13g2_decap_8 FILLER_17_1720 ();
 sg13g2_decap_8 FILLER_17_1727 ();
 sg13g2_decap_8 FILLER_17_1734 ();
 sg13g2_decap_8 FILLER_17_1741 ();
 sg13g2_decap_8 FILLER_17_1748 ();
 sg13g2_decap_8 FILLER_17_1755 ();
 sg13g2_decap_4 FILLER_17_1762 ();
 sg13g2_fill_2 FILLER_17_1766 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_1 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_139 ();
 sg13g2_fill_2 FILLER_18_149 ();
 sg13g2_fill_2 FILLER_18_202 ();
 sg13g2_fill_1 FILLER_18_204 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_fill_2 FILLER_18_274 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_fill_2 FILLER_18_289 ();
 sg13g2_fill_1 FILLER_18_300 ();
 sg13g2_fill_2 FILLER_18_323 ();
 sg13g2_fill_1 FILLER_18_325 ();
 sg13g2_fill_2 FILLER_18_343 ();
 sg13g2_fill_2 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_356 ();
 sg13g2_fill_2 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_470 ();
 sg13g2_fill_1 FILLER_18_489 ();
 sg13g2_fill_2 FILLER_18_498 ();
 sg13g2_fill_2 FILLER_18_529 ();
 sg13g2_fill_1 FILLER_18_531 ();
 sg13g2_fill_2 FILLER_18_558 ();
 sg13g2_fill_1 FILLER_18_569 ();
 sg13g2_fill_1 FILLER_18_610 ();
 sg13g2_fill_2 FILLER_18_634 ();
 sg13g2_fill_2 FILLER_18_728 ();
 sg13g2_fill_1 FILLER_18_730 ();
 sg13g2_fill_2 FILLER_18_762 ();
 sg13g2_fill_2 FILLER_18_803 ();
 sg13g2_fill_2 FILLER_18_821 ();
 sg13g2_fill_1 FILLER_18_837 ();
 sg13g2_fill_2 FILLER_18_852 ();
 sg13g2_fill_1 FILLER_18_905 ();
 sg13g2_decap_4 FILLER_18_922 ();
 sg13g2_fill_2 FILLER_18_926 ();
 sg13g2_fill_2 FILLER_18_957 ();
 sg13g2_fill_2 FILLER_18_1026 ();
 sg13g2_fill_1 FILLER_18_1028 ();
 sg13g2_fill_2 FILLER_18_1063 ();
 sg13g2_fill_1 FILLER_18_1065 ();
 sg13g2_fill_2 FILLER_18_1157 ();
 sg13g2_fill_1 FILLER_18_1159 ();
 sg13g2_fill_1 FILLER_18_1182 ();
 sg13g2_fill_2 FILLER_18_1187 ();
 sg13g2_fill_2 FILLER_18_1193 ();
 sg13g2_fill_1 FILLER_18_1195 ();
 sg13g2_fill_2 FILLER_18_1220 ();
 sg13g2_fill_1 FILLER_18_1222 ();
 sg13g2_fill_2 FILLER_18_1258 ();
 sg13g2_fill_2 FILLER_18_1336 ();
 sg13g2_fill_2 FILLER_18_1364 ();
 sg13g2_fill_1 FILLER_18_1366 ();
 sg13g2_fill_2 FILLER_18_1421 ();
 sg13g2_fill_1 FILLER_18_1423 ();
 sg13g2_fill_2 FILLER_18_1448 ();
 sg13g2_fill_1 FILLER_18_1458 ();
 sg13g2_fill_2 FILLER_18_1485 ();
 sg13g2_fill_1 FILLER_18_1487 ();
 sg13g2_fill_1 FILLER_18_1528 ();
 sg13g2_decap_8 FILLER_18_1563 ();
 sg13g2_decap_8 FILLER_18_1570 ();
 sg13g2_decap_8 FILLER_18_1577 ();
 sg13g2_decap_8 FILLER_18_1584 ();
 sg13g2_decap_8 FILLER_18_1591 ();
 sg13g2_decap_8 FILLER_18_1598 ();
 sg13g2_decap_8 FILLER_18_1605 ();
 sg13g2_decap_8 FILLER_18_1612 ();
 sg13g2_decap_8 FILLER_18_1619 ();
 sg13g2_decap_8 FILLER_18_1626 ();
 sg13g2_decap_8 FILLER_18_1633 ();
 sg13g2_decap_8 FILLER_18_1640 ();
 sg13g2_decap_8 FILLER_18_1647 ();
 sg13g2_decap_8 FILLER_18_1654 ();
 sg13g2_decap_8 FILLER_18_1661 ();
 sg13g2_decap_8 FILLER_18_1668 ();
 sg13g2_decap_8 FILLER_18_1675 ();
 sg13g2_decap_8 FILLER_18_1682 ();
 sg13g2_decap_8 FILLER_18_1689 ();
 sg13g2_decap_8 FILLER_18_1696 ();
 sg13g2_decap_8 FILLER_18_1703 ();
 sg13g2_decap_8 FILLER_18_1710 ();
 sg13g2_decap_8 FILLER_18_1717 ();
 sg13g2_decap_8 FILLER_18_1724 ();
 sg13g2_decap_8 FILLER_18_1731 ();
 sg13g2_decap_8 FILLER_18_1738 ();
 sg13g2_decap_8 FILLER_18_1745 ();
 sg13g2_decap_8 FILLER_18_1752 ();
 sg13g2_decap_8 FILLER_18_1759 ();
 sg13g2_fill_2 FILLER_18_1766 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_83 ();
 sg13g2_fill_2 FILLER_19_115 ();
 sg13g2_fill_2 FILLER_19_143 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_fill_2 FILLER_19_284 ();
 sg13g2_fill_1 FILLER_19_286 ();
 sg13g2_fill_2 FILLER_19_365 ();
 sg13g2_fill_1 FILLER_19_367 ();
 sg13g2_decap_4 FILLER_19_407 ();
 sg13g2_fill_1 FILLER_19_433 ();
 sg13g2_fill_2 FILLER_19_439 ();
 sg13g2_fill_1 FILLER_19_441 ();
 sg13g2_fill_2 FILLER_19_454 ();
 sg13g2_fill_1 FILLER_19_456 ();
 sg13g2_fill_1 FILLER_19_498 ();
 sg13g2_fill_2 FILLER_19_503 ();
 sg13g2_fill_1 FILLER_19_505 ();
 sg13g2_fill_2 FILLER_19_514 ();
 sg13g2_fill_1 FILLER_19_530 ();
 sg13g2_fill_1 FILLER_19_566 ();
 sg13g2_fill_1 FILLER_19_577 ();
 sg13g2_fill_2 FILLER_19_649 ();
 sg13g2_fill_1 FILLER_19_677 ();
 sg13g2_fill_2 FILLER_19_704 ();
 sg13g2_fill_1 FILLER_19_706 ();
 sg13g2_fill_2 FILLER_19_766 ();
 sg13g2_fill_1 FILLER_19_768 ();
 sg13g2_fill_2 FILLER_19_804 ();
 sg13g2_fill_1 FILLER_19_806 ();
 sg13g2_fill_2 FILLER_19_884 ();
 sg13g2_fill_1 FILLER_19_886 ();
 sg13g2_fill_1 FILLER_19_953 ();
 sg13g2_fill_2 FILLER_19_1003 ();
 sg13g2_fill_1 FILLER_19_1011 ();
 sg13g2_fill_2 FILLER_19_1029 ();
 sg13g2_fill_2 FILLER_19_1036 ();
 sg13g2_fill_2 FILLER_19_1090 ();
 sg13g2_fill_1 FILLER_19_1092 ();
 sg13g2_fill_1 FILLER_19_1163 ();
 sg13g2_fill_2 FILLER_19_1191 ();
 sg13g2_fill_2 FILLER_19_1223 ();
 sg13g2_fill_1 FILLER_19_1267 ();
 sg13g2_fill_2 FILLER_19_1341 ();
 sg13g2_fill_1 FILLER_19_1348 ();
 sg13g2_fill_1 FILLER_19_1378 ();
 sg13g2_fill_1 FILLER_19_1388 ();
 sg13g2_fill_1 FILLER_19_1394 ();
 sg13g2_fill_1 FILLER_19_1407 ();
 sg13g2_fill_2 FILLER_19_1418 ();
 sg13g2_fill_2 FILLER_19_1434 ();
 sg13g2_fill_2 FILLER_19_1475 ();
 sg13g2_fill_1 FILLER_19_1477 ();
 sg13g2_fill_2 FILLER_19_1487 ();
 sg13g2_fill_1 FILLER_19_1489 ();
 sg13g2_fill_1 FILLER_19_1550 ();
 sg13g2_decap_8 FILLER_19_1572 ();
 sg13g2_decap_8 FILLER_19_1579 ();
 sg13g2_decap_8 FILLER_19_1586 ();
 sg13g2_decap_8 FILLER_19_1593 ();
 sg13g2_decap_8 FILLER_19_1600 ();
 sg13g2_decap_8 FILLER_19_1607 ();
 sg13g2_decap_8 FILLER_19_1614 ();
 sg13g2_decap_8 FILLER_19_1621 ();
 sg13g2_decap_8 FILLER_19_1628 ();
 sg13g2_decap_8 FILLER_19_1635 ();
 sg13g2_decap_8 FILLER_19_1642 ();
 sg13g2_decap_8 FILLER_19_1649 ();
 sg13g2_decap_8 FILLER_19_1656 ();
 sg13g2_decap_8 FILLER_19_1663 ();
 sg13g2_decap_8 FILLER_19_1670 ();
 sg13g2_decap_8 FILLER_19_1677 ();
 sg13g2_decap_8 FILLER_19_1684 ();
 sg13g2_decap_8 FILLER_19_1691 ();
 sg13g2_decap_8 FILLER_19_1698 ();
 sg13g2_decap_8 FILLER_19_1705 ();
 sg13g2_decap_8 FILLER_19_1712 ();
 sg13g2_decap_8 FILLER_19_1719 ();
 sg13g2_decap_8 FILLER_19_1726 ();
 sg13g2_decap_8 FILLER_19_1733 ();
 sg13g2_decap_8 FILLER_19_1740 ();
 sg13g2_decap_8 FILLER_19_1747 ();
 sg13g2_decap_8 FILLER_19_1754 ();
 sg13g2_decap_8 FILLER_19_1761 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_27 ();
 sg13g2_fill_2 FILLER_20_53 ();
 sg13g2_fill_1 FILLER_20_55 ();
 sg13g2_fill_2 FILLER_20_62 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_fill_1 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_186 ();
 sg13g2_fill_1 FILLER_20_222 ();
 sg13g2_fill_1 FILLER_20_249 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_fill_1 FILLER_20_308 ();
 sg13g2_fill_2 FILLER_20_332 ();
 sg13g2_fill_1 FILLER_20_339 ();
 sg13g2_fill_1 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_fill_1 FILLER_20_450 ();
 sg13g2_fill_2 FILLER_20_515 ();
 sg13g2_fill_1 FILLER_20_517 ();
 sg13g2_fill_2 FILLER_20_558 ();
 sg13g2_fill_1 FILLER_20_560 ();
 sg13g2_fill_1 FILLER_20_576 ();
 sg13g2_fill_1 FILLER_20_582 ();
 sg13g2_fill_2 FILLER_20_601 ();
 sg13g2_fill_1 FILLER_20_670 ();
 sg13g2_fill_1 FILLER_20_702 ();
 sg13g2_fill_1 FILLER_20_708 ();
 sg13g2_fill_2 FILLER_20_725 ();
 sg13g2_fill_1 FILLER_20_805 ();
 sg13g2_fill_1 FILLER_20_822 ();
 sg13g2_fill_2 FILLER_20_914 ();
 sg13g2_fill_1 FILLER_20_916 ();
 sg13g2_fill_2 FILLER_20_929 ();
 sg13g2_fill_1 FILLER_20_931 ();
 sg13g2_fill_1 FILLER_20_970 ();
 sg13g2_fill_2 FILLER_20_1035 ();
 sg13g2_fill_1 FILLER_20_1037 ();
 sg13g2_decap_8 FILLER_20_1051 ();
 sg13g2_fill_1 FILLER_20_1072 ();
 sg13g2_fill_2 FILLER_20_1079 ();
 sg13g2_fill_1 FILLER_20_1143 ();
 sg13g2_fill_2 FILLER_20_1205 ();
 sg13g2_fill_1 FILLER_20_1207 ();
 sg13g2_fill_1 FILLER_20_1223 ();
 sg13g2_fill_1 FILLER_20_1240 ();
 sg13g2_fill_1 FILLER_20_1256 ();
 sg13g2_fill_2 FILLER_20_1303 ();
 sg13g2_fill_1 FILLER_20_1305 ();
 sg13g2_fill_2 FILLER_20_1398 ();
 sg13g2_fill_2 FILLER_20_1431 ();
 sg13g2_fill_1 FILLER_20_1433 ();
 sg13g2_fill_2 FILLER_20_1460 ();
 sg13g2_fill_1 FILLER_20_1462 ();
 sg13g2_fill_2 FILLER_20_1495 ();
 sg13g2_fill_1 FILLER_20_1497 ();
 sg13g2_fill_2 FILLER_20_1515 ();
 sg13g2_fill_1 FILLER_20_1540 ();
 sg13g2_decap_8 FILLER_20_1583 ();
 sg13g2_decap_8 FILLER_20_1590 ();
 sg13g2_decap_8 FILLER_20_1597 ();
 sg13g2_decap_8 FILLER_20_1604 ();
 sg13g2_decap_8 FILLER_20_1611 ();
 sg13g2_decap_8 FILLER_20_1618 ();
 sg13g2_decap_8 FILLER_20_1625 ();
 sg13g2_decap_8 FILLER_20_1632 ();
 sg13g2_decap_8 FILLER_20_1639 ();
 sg13g2_decap_8 FILLER_20_1646 ();
 sg13g2_decap_8 FILLER_20_1653 ();
 sg13g2_decap_8 FILLER_20_1660 ();
 sg13g2_decap_8 FILLER_20_1667 ();
 sg13g2_decap_8 FILLER_20_1674 ();
 sg13g2_decap_8 FILLER_20_1681 ();
 sg13g2_decap_8 FILLER_20_1688 ();
 sg13g2_decap_8 FILLER_20_1695 ();
 sg13g2_decap_8 FILLER_20_1702 ();
 sg13g2_decap_8 FILLER_20_1709 ();
 sg13g2_decap_8 FILLER_20_1716 ();
 sg13g2_decap_8 FILLER_20_1723 ();
 sg13g2_decap_8 FILLER_20_1730 ();
 sg13g2_decap_8 FILLER_20_1737 ();
 sg13g2_decap_8 FILLER_20_1744 ();
 sg13g2_decap_8 FILLER_20_1751 ();
 sg13g2_decap_8 FILLER_20_1758 ();
 sg13g2_fill_2 FILLER_20_1765 ();
 sg13g2_fill_1 FILLER_20_1767 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_32 ();
 sg13g2_fill_1 FILLER_21_34 ();
 sg13g2_fill_1 FILLER_21_87 ();
 sg13g2_fill_1 FILLER_21_116 ();
 sg13g2_decap_4 FILLER_21_148 ();
 sg13g2_fill_1 FILLER_21_152 ();
 sg13g2_fill_1 FILLER_21_183 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_244 ();
 sg13g2_fill_2 FILLER_21_258 ();
 sg13g2_fill_2 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_331 ();
 sg13g2_fill_2 FILLER_21_359 ();
 sg13g2_fill_1 FILLER_21_381 ();
 sg13g2_fill_2 FILLER_21_394 ();
 sg13g2_fill_2 FILLER_21_414 ();
 sg13g2_fill_1 FILLER_21_416 ();
 sg13g2_fill_2 FILLER_21_434 ();
 sg13g2_fill_2 FILLER_21_457 ();
 sg13g2_fill_1 FILLER_21_459 ();
 sg13g2_fill_2 FILLER_21_495 ();
 sg13g2_fill_2 FILLER_21_525 ();
 sg13g2_fill_2 FILLER_21_541 ();
 sg13g2_fill_1 FILLER_21_543 ();
 sg13g2_decap_4 FILLER_21_612 ();
 sg13g2_fill_2 FILLER_21_616 ();
 sg13g2_decap_4 FILLER_21_626 ();
 sg13g2_fill_2 FILLER_21_635 ();
 sg13g2_fill_1 FILLER_21_651 ();
 sg13g2_fill_2 FILLER_21_662 ();
 sg13g2_fill_1 FILLER_21_694 ();
 sg13g2_fill_1 FILLER_21_703 ();
 sg13g2_fill_2 FILLER_21_730 ();
 sg13g2_fill_1 FILLER_21_759 ();
 sg13g2_fill_2 FILLER_21_769 ();
 sg13g2_fill_1 FILLER_21_771 ();
 sg13g2_fill_1 FILLER_21_786 ();
 sg13g2_fill_1 FILLER_21_791 ();
 sg13g2_fill_2 FILLER_21_818 ();
 sg13g2_fill_2 FILLER_21_835 ();
 sg13g2_fill_1 FILLER_21_837 ();
 sg13g2_fill_1 FILLER_21_906 ();
 sg13g2_fill_1 FILLER_21_964 ();
 sg13g2_fill_1 FILLER_21_970 ();
 sg13g2_decap_4 FILLER_21_1050 ();
 sg13g2_fill_1 FILLER_21_1106 ();
 sg13g2_fill_2 FILLER_21_1118 ();
 sg13g2_fill_1 FILLER_21_1125 ();
 sg13g2_fill_2 FILLER_21_1133 ();
 sg13g2_fill_1 FILLER_21_1148 ();
 sg13g2_fill_1 FILLER_21_1158 ();
 sg13g2_fill_2 FILLER_21_1212 ();
 sg13g2_fill_1 FILLER_21_1235 ();
 sg13g2_fill_2 FILLER_21_1245 ();
 sg13g2_fill_2 FILLER_21_1292 ();
 sg13g2_fill_2 FILLER_21_1339 ();
 sg13g2_fill_1 FILLER_21_1369 ();
 sg13g2_fill_2 FILLER_21_1426 ();
 sg13g2_fill_1 FILLER_21_1455 ();
 sg13g2_fill_1 FILLER_21_1479 ();
 sg13g2_fill_2 FILLER_21_1520 ();
 sg13g2_fill_1 FILLER_21_1522 ();
 sg13g2_fill_2 FILLER_21_1528 ();
 sg13g2_fill_1 FILLER_21_1530 ();
 sg13g2_decap_8 FILLER_21_1566 ();
 sg13g2_decap_8 FILLER_21_1573 ();
 sg13g2_decap_8 FILLER_21_1580 ();
 sg13g2_decap_8 FILLER_21_1587 ();
 sg13g2_decap_8 FILLER_21_1594 ();
 sg13g2_decap_8 FILLER_21_1601 ();
 sg13g2_decap_8 FILLER_21_1608 ();
 sg13g2_decap_8 FILLER_21_1615 ();
 sg13g2_decap_8 FILLER_21_1622 ();
 sg13g2_decap_8 FILLER_21_1629 ();
 sg13g2_decap_8 FILLER_21_1636 ();
 sg13g2_decap_8 FILLER_21_1643 ();
 sg13g2_decap_8 FILLER_21_1650 ();
 sg13g2_decap_8 FILLER_21_1657 ();
 sg13g2_decap_8 FILLER_21_1664 ();
 sg13g2_decap_8 FILLER_21_1671 ();
 sg13g2_decap_8 FILLER_21_1678 ();
 sg13g2_decap_8 FILLER_21_1685 ();
 sg13g2_decap_8 FILLER_21_1692 ();
 sg13g2_decap_8 FILLER_21_1699 ();
 sg13g2_decap_8 FILLER_21_1706 ();
 sg13g2_decap_8 FILLER_21_1713 ();
 sg13g2_decap_8 FILLER_21_1720 ();
 sg13g2_decap_8 FILLER_21_1727 ();
 sg13g2_decap_8 FILLER_21_1734 ();
 sg13g2_decap_8 FILLER_21_1741 ();
 sg13g2_decap_8 FILLER_21_1748 ();
 sg13g2_decap_8 FILLER_21_1755 ();
 sg13g2_decap_4 FILLER_21_1762 ();
 sg13g2_fill_2 FILLER_21_1766 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_36 ();
 sg13g2_fill_1 FILLER_22_38 ();
 sg13g2_fill_2 FILLER_22_67 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_fill_2 FILLER_22_80 ();
 sg13g2_fill_1 FILLER_22_170 ();
 sg13g2_fill_1 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_199 ();
 sg13g2_fill_1 FILLER_22_201 ();
 sg13g2_fill_2 FILLER_22_257 ();
 sg13g2_fill_2 FILLER_22_272 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_355 ();
 sg13g2_fill_1 FILLER_22_374 ();
 sg13g2_fill_2 FILLER_22_399 ();
 sg13g2_decap_4 FILLER_22_409 ();
 sg13g2_fill_1 FILLER_22_439 ();
 sg13g2_fill_1 FILLER_22_462 ();
 sg13g2_fill_1 FILLER_22_476 ();
 sg13g2_fill_2 FILLER_22_483 ();
 sg13g2_fill_1 FILLER_22_485 ();
 sg13g2_fill_1 FILLER_22_491 ();
 sg13g2_fill_2 FILLER_22_556 ();
 sg13g2_decap_4 FILLER_22_590 ();
 sg13g2_fill_1 FILLER_22_638 ();
 sg13g2_fill_1 FILLER_22_675 ();
 sg13g2_fill_2 FILLER_22_689 ();
 sg13g2_fill_2 FILLER_22_695 ();
 sg13g2_fill_1 FILLER_22_697 ();
 sg13g2_fill_2 FILLER_22_727 ();
 sg13g2_fill_1 FILLER_22_729 ();
 sg13g2_fill_2 FILLER_22_736 ();
 sg13g2_fill_1 FILLER_22_805 ();
 sg13g2_fill_1 FILLER_22_848 ();
 sg13g2_fill_2 FILLER_22_918 ();
 sg13g2_fill_2 FILLER_22_953 ();
 sg13g2_fill_2 FILLER_22_994 ();
 sg13g2_fill_1 FILLER_22_996 ();
 sg13g2_fill_1 FILLER_22_1065 ();
 sg13g2_fill_1 FILLER_22_1128 ();
 sg13g2_fill_2 FILLER_22_1136 ();
 sg13g2_fill_2 FILLER_22_1203 ();
 sg13g2_fill_1 FILLER_22_1205 ();
 sg13g2_fill_2 FILLER_22_1328 ();
 sg13g2_fill_2 FILLER_22_1345 ();
 sg13g2_fill_1 FILLER_22_1377 ();
 sg13g2_fill_1 FILLER_22_1383 ();
 sg13g2_fill_2 FILLER_22_1396 ();
 sg13g2_decap_4 FILLER_22_1431 ();
 sg13g2_decap_8 FILLER_22_1571 ();
 sg13g2_decap_8 FILLER_22_1578 ();
 sg13g2_decap_8 FILLER_22_1585 ();
 sg13g2_decap_8 FILLER_22_1592 ();
 sg13g2_decap_8 FILLER_22_1599 ();
 sg13g2_decap_8 FILLER_22_1606 ();
 sg13g2_decap_8 FILLER_22_1613 ();
 sg13g2_decap_8 FILLER_22_1620 ();
 sg13g2_decap_8 FILLER_22_1627 ();
 sg13g2_decap_8 FILLER_22_1634 ();
 sg13g2_decap_8 FILLER_22_1641 ();
 sg13g2_decap_8 FILLER_22_1648 ();
 sg13g2_decap_8 FILLER_22_1655 ();
 sg13g2_decap_8 FILLER_22_1662 ();
 sg13g2_decap_8 FILLER_22_1669 ();
 sg13g2_decap_8 FILLER_22_1676 ();
 sg13g2_decap_8 FILLER_22_1683 ();
 sg13g2_decap_8 FILLER_22_1690 ();
 sg13g2_decap_8 FILLER_22_1697 ();
 sg13g2_decap_8 FILLER_22_1704 ();
 sg13g2_decap_8 FILLER_22_1711 ();
 sg13g2_decap_8 FILLER_22_1718 ();
 sg13g2_decap_8 FILLER_22_1725 ();
 sg13g2_decap_8 FILLER_22_1732 ();
 sg13g2_decap_8 FILLER_22_1739 ();
 sg13g2_decap_8 FILLER_22_1746 ();
 sg13g2_decap_8 FILLER_22_1753 ();
 sg13g2_decap_8 FILLER_22_1760 ();
 sg13g2_fill_1 FILLER_22_1767 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_37 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_80 ();
 sg13g2_fill_1 FILLER_23_87 ();
 sg13g2_fill_1 FILLER_23_118 ();
 sg13g2_fill_2 FILLER_23_129 ();
 sg13g2_fill_1 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_fill_2 FILLER_23_203 ();
 sg13g2_fill_2 FILLER_23_218 ();
 sg13g2_fill_2 FILLER_23_230 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_260 ();
 sg13g2_fill_2 FILLER_23_313 ();
 sg13g2_fill_1 FILLER_23_325 ();
 sg13g2_fill_1 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_388 ();
 sg13g2_fill_2 FILLER_23_392 ();
 sg13g2_fill_1 FILLER_23_400 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_fill_2 FILLER_23_446 ();
 sg13g2_fill_1 FILLER_23_448 ();
 sg13g2_fill_2 FILLER_23_454 ();
 sg13g2_fill_1 FILLER_23_456 ();
 sg13g2_fill_2 FILLER_23_535 ();
 sg13g2_fill_1 FILLER_23_537 ();
 sg13g2_fill_1 FILLER_23_562 ();
 sg13g2_decap_4 FILLER_23_593 ();
 sg13g2_fill_1 FILLER_23_602 ();
 sg13g2_fill_2 FILLER_23_620 ();
 sg13g2_fill_2 FILLER_23_647 ();
 sg13g2_fill_1 FILLER_23_662 ();
 sg13g2_fill_1 FILLER_23_672 ();
 sg13g2_fill_2 FILLER_23_688 ();
 sg13g2_fill_1 FILLER_23_690 ();
 sg13g2_fill_1 FILLER_23_794 ();
 sg13g2_fill_2 FILLER_23_800 ();
 sg13g2_fill_1 FILLER_23_802 ();
 sg13g2_fill_1 FILLER_23_808 ();
 sg13g2_fill_1 FILLER_23_821 ();
 sg13g2_fill_2 FILLER_23_841 ();
 sg13g2_fill_2 FILLER_23_852 ();
 sg13g2_fill_1 FILLER_23_863 ();
 sg13g2_fill_2 FILLER_23_868 ();
 sg13g2_decap_4 FILLER_23_898 ();
 sg13g2_fill_1 FILLER_23_902 ();
 sg13g2_fill_1 FILLER_23_907 ();
 sg13g2_fill_2 FILLER_23_918 ();
 sg13g2_fill_1 FILLER_23_920 ();
 sg13g2_fill_2 FILLER_23_958 ();
 sg13g2_fill_1 FILLER_23_965 ();
 sg13g2_fill_2 FILLER_23_981 ();
 sg13g2_fill_1 FILLER_23_1009 ();
 sg13g2_fill_2 FILLER_23_1166 ();
 sg13g2_fill_2 FILLER_23_1187 ();
 sg13g2_fill_2 FILLER_23_1224 ();
 sg13g2_fill_1 FILLER_23_1226 ();
 sg13g2_fill_2 FILLER_23_1235 ();
 sg13g2_fill_2 FILLER_23_1324 ();
 sg13g2_fill_1 FILLER_23_1326 ();
 sg13g2_fill_1 FILLER_23_1392 ();
 sg13g2_fill_2 FILLER_23_1415 ();
 sg13g2_fill_2 FILLER_23_1439 ();
 sg13g2_fill_1 FILLER_23_1441 ();
 sg13g2_fill_2 FILLER_23_1478 ();
 sg13g2_fill_1 FILLER_23_1480 ();
 sg13g2_fill_2 FILLER_23_1486 ();
 sg13g2_fill_2 FILLER_23_1528 ();
 sg13g2_decap_8 FILLER_23_1556 ();
 sg13g2_decap_8 FILLER_23_1563 ();
 sg13g2_decap_8 FILLER_23_1570 ();
 sg13g2_decap_8 FILLER_23_1577 ();
 sg13g2_decap_8 FILLER_23_1584 ();
 sg13g2_decap_8 FILLER_23_1591 ();
 sg13g2_decap_8 FILLER_23_1598 ();
 sg13g2_decap_8 FILLER_23_1605 ();
 sg13g2_decap_8 FILLER_23_1612 ();
 sg13g2_decap_8 FILLER_23_1619 ();
 sg13g2_decap_8 FILLER_23_1626 ();
 sg13g2_decap_8 FILLER_23_1633 ();
 sg13g2_decap_8 FILLER_23_1640 ();
 sg13g2_decap_8 FILLER_23_1647 ();
 sg13g2_decap_8 FILLER_23_1654 ();
 sg13g2_decap_8 FILLER_23_1661 ();
 sg13g2_decap_8 FILLER_23_1668 ();
 sg13g2_decap_8 FILLER_23_1675 ();
 sg13g2_decap_8 FILLER_23_1682 ();
 sg13g2_decap_8 FILLER_23_1689 ();
 sg13g2_decap_8 FILLER_23_1696 ();
 sg13g2_decap_8 FILLER_23_1703 ();
 sg13g2_decap_8 FILLER_23_1710 ();
 sg13g2_decap_8 FILLER_23_1717 ();
 sg13g2_decap_8 FILLER_23_1724 ();
 sg13g2_decap_8 FILLER_23_1731 ();
 sg13g2_decap_8 FILLER_23_1738 ();
 sg13g2_decap_8 FILLER_23_1745 ();
 sg13g2_decap_8 FILLER_23_1752 ();
 sg13g2_decap_8 FILLER_23_1759 ();
 sg13g2_fill_2 FILLER_23_1766 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_fill_2 FILLER_24_61 ();
 sg13g2_fill_1 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_155 ();
 sg13g2_fill_1 FILLER_24_157 ();
 sg13g2_fill_2 FILLER_24_169 ();
 sg13g2_fill_2 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_324 ();
 sg13g2_fill_1 FILLER_24_330 ();
 sg13g2_fill_1 FILLER_24_339 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_1 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_371 ();
 sg13g2_decap_4 FILLER_24_402 ();
 sg13g2_fill_2 FILLER_24_414 ();
 sg13g2_fill_1 FILLER_24_416 ();
 sg13g2_fill_1 FILLER_24_438 ();
 sg13g2_fill_2 FILLER_24_448 ();
 sg13g2_fill_1 FILLER_24_450 ();
 sg13g2_fill_2 FILLER_24_464 ();
 sg13g2_fill_1 FILLER_24_510 ();
 sg13g2_fill_1 FILLER_24_546 ();
 sg13g2_decap_4 FILLER_24_587 ();
 sg13g2_fill_2 FILLER_24_591 ();
 sg13g2_fill_1 FILLER_24_619 ();
 sg13g2_fill_2 FILLER_24_689 ();
 sg13g2_fill_2 FILLER_24_716 ();
 sg13g2_fill_1 FILLER_24_731 ();
 sg13g2_fill_1 FILLER_24_763 ();
 sg13g2_fill_1 FILLER_24_852 ();
 sg13g2_fill_2 FILLER_24_888 ();
 sg13g2_fill_1 FILLER_24_911 ();
 sg13g2_fill_2 FILLER_24_920 ();
 sg13g2_fill_1 FILLER_24_922 ();
 sg13g2_fill_1 FILLER_24_936 ();
 sg13g2_fill_1 FILLER_24_993 ();
 sg13g2_fill_2 FILLER_24_1005 ();
 sg13g2_fill_1 FILLER_24_1007 ();
 sg13g2_fill_2 FILLER_24_1057 ();
 sg13g2_fill_1 FILLER_24_1086 ();
 sg13g2_fill_1 FILLER_24_1105 ();
 sg13g2_fill_1 FILLER_24_1136 ();
 sg13g2_fill_2 FILLER_24_1191 ();
 sg13g2_fill_1 FILLER_24_1224 ();
 sg13g2_fill_1 FILLER_24_1233 ();
 sg13g2_fill_1 FILLER_24_1247 ();
 sg13g2_fill_1 FILLER_24_1256 ();
 sg13g2_fill_2 FILLER_24_1262 ();
 sg13g2_fill_2 FILLER_24_1287 ();
 sg13g2_fill_1 FILLER_24_1289 ();
 sg13g2_fill_1 FILLER_24_1307 ();
 sg13g2_fill_2 FILLER_24_1321 ();
 sg13g2_fill_1 FILLER_24_1364 ();
 sg13g2_fill_1 FILLER_24_1384 ();
 sg13g2_fill_2 FILLER_24_1403 ();
 sg13g2_fill_1 FILLER_24_1448 ();
 sg13g2_fill_2 FILLER_24_1461 ();
 sg13g2_fill_1 FILLER_24_1476 ();
 sg13g2_fill_2 FILLER_24_1486 ();
 sg13g2_fill_2 FILLER_24_1494 ();
 sg13g2_fill_1 FILLER_24_1496 ();
 sg13g2_fill_2 FILLER_24_1513 ();
 sg13g2_fill_1 FILLER_24_1515 ();
 sg13g2_decap_8 FILLER_24_1554 ();
 sg13g2_decap_8 FILLER_24_1561 ();
 sg13g2_decap_8 FILLER_24_1568 ();
 sg13g2_decap_8 FILLER_24_1575 ();
 sg13g2_decap_8 FILLER_24_1582 ();
 sg13g2_decap_8 FILLER_24_1589 ();
 sg13g2_decap_8 FILLER_24_1596 ();
 sg13g2_decap_8 FILLER_24_1603 ();
 sg13g2_decap_8 FILLER_24_1610 ();
 sg13g2_decap_8 FILLER_24_1617 ();
 sg13g2_decap_8 FILLER_24_1624 ();
 sg13g2_decap_8 FILLER_24_1631 ();
 sg13g2_decap_8 FILLER_24_1638 ();
 sg13g2_decap_8 FILLER_24_1645 ();
 sg13g2_decap_8 FILLER_24_1652 ();
 sg13g2_decap_8 FILLER_24_1659 ();
 sg13g2_decap_8 FILLER_24_1666 ();
 sg13g2_decap_8 FILLER_24_1673 ();
 sg13g2_decap_8 FILLER_24_1680 ();
 sg13g2_decap_8 FILLER_24_1687 ();
 sg13g2_decap_8 FILLER_24_1694 ();
 sg13g2_decap_8 FILLER_24_1701 ();
 sg13g2_decap_8 FILLER_24_1708 ();
 sg13g2_decap_8 FILLER_24_1715 ();
 sg13g2_decap_8 FILLER_24_1722 ();
 sg13g2_decap_8 FILLER_24_1729 ();
 sg13g2_decap_8 FILLER_24_1736 ();
 sg13g2_decap_8 FILLER_24_1743 ();
 sg13g2_decap_8 FILLER_24_1750 ();
 sg13g2_decap_8 FILLER_24_1757 ();
 sg13g2_decap_4 FILLER_24_1764 ();
 sg13g2_fill_1 FILLER_25_35 ();
 sg13g2_fill_1 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_66 ();
 sg13g2_fill_1 FILLER_25_161 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_215 ();
 sg13g2_fill_2 FILLER_25_242 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_281 ();
 sg13g2_fill_2 FILLER_25_304 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_fill_2 FILLER_25_410 ();
 sg13g2_fill_1 FILLER_25_474 ();
 sg13g2_fill_2 FILLER_25_480 ();
 sg13g2_fill_1 FILLER_25_482 ();
 sg13g2_fill_2 FILLER_25_494 ();
 sg13g2_fill_1 FILLER_25_496 ();
 sg13g2_fill_2 FILLER_25_523 ();
 sg13g2_fill_1 FILLER_25_525 ();
 sg13g2_fill_1 FILLER_25_535 ();
 sg13g2_decap_8 FILLER_25_587 ();
 sg13g2_fill_2 FILLER_25_599 ();
 sg13g2_fill_1 FILLER_25_605 ();
 sg13g2_fill_1 FILLER_25_638 ();
 sg13g2_fill_1 FILLER_25_656 ();
 sg13g2_fill_1 FILLER_25_663 ();
 sg13g2_fill_2 FILLER_25_759 ();
 sg13g2_fill_2 FILLER_25_800 ();
 sg13g2_fill_1 FILLER_25_802 ();
 sg13g2_fill_2 FILLER_25_849 ();
 sg13g2_fill_2 FILLER_25_863 ();
 sg13g2_fill_1 FILLER_25_878 ();
 sg13g2_decap_8 FILLER_25_887 ();
 sg13g2_fill_2 FILLER_25_894 ();
 sg13g2_fill_1 FILLER_25_896 ();
 sg13g2_fill_2 FILLER_25_927 ();
 sg13g2_decap_4 FILLER_25_942 ();
 sg13g2_fill_2 FILLER_25_954 ();
 sg13g2_fill_1 FILLER_25_956 ();
 sg13g2_fill_2 FILLER_25_967 ();
 sg13g2_fill_1 FILLER_25_995 ();
 sg13g2_fill_2 FILLER_25_1004 ();
 sg13g2_fill_2 FILLER_25_1035 ();
 sg13g2_fill_2 FILLER_25_1076 ();
 sg13g2_fill_2 FILLER_25_1112 ();
 sg13g2_fill_2 FILLER_25_1119 ();
 sg13g2_fill_2 FILLER_25_1130 ();
 sg13g2_fill_1 FILLER_25_1132 ();
 sg13g2_fill_2 FILLER_25_1138 ();
 sg13g2_fill_1 FILLER_25_1155 ();
 sg13g2_fill_2 FILLER_25_1210 ();
 sg13g2_fill_1 FILLER_25_1212 ();
 sg13g2_fill_1 FILLER_25_1222 ();
 sg13g2_fill_2 FILLER_25_1352 ();
 sg13g2_fill_1 FILLER_25_1354 ();
 sg13g2_fill_1 FILLER_25_1431 ();
 sg13g2_fill_2 FILLER_25_1473 ();
 sg13g2_fill_2 FILLER_25_1515 ();
 sg13g2_fill_1 FILLER_25_1517 ();
 sg13g2_decap_8 FILLER_25_1549 ();
 sg13g2_decap_8 FILLER_25_1556 ();
 sg13g2_decap_8 FILLER_25_1563 ();
 sg13g2_decap_8 FILLER_25_1570 ();
 sg13g2_decap_8 FILLER_25_1577 ();
 sg13g2_decap_8 FILLER_25_1584 ();
 sg13g2_decap_8 FILLER_25_1591 ();
 sg13g2_decap_8 FILLER_25_1598 ();
 sg13g2_decap_8 FILLER_25_1605 ();
 sg13g2_decap_8 FILLER_25_1612 ();
 sg13g2_decap_8 FILLER_25_1619 ();
 sg13g2_decap_8 FILLER_25_1626 ();
 sg13g2_decap_8 FILLER_25_1633 ();
 sg13g2_decap_8 FILLER_25_1640 ();
 sg13g2_decap_8 FILLER_25_1647 ();
 sg13g2_decap_8 FILLER_25_1654 ();
 sg13g2_decap_8 FILLER_25_1661 ();
 sg13g2_decap_8 FILLER_25_1668 ();
 sg13g2_decap_8 FILLER_25_1675 ();
 sg13g2_decap_8 FILLER_25_1682 ();
 sg13g2_decap_8 FILLER_25_1689 ();
 sg13g2_decap_8 FILLER_25_1696 ();
 sg13g2_decap_8 FILLER_25_1703 ();
 sg13g2_decap_8 FILLER_25_1710 ();
 sg13g2_decap_8 FILLER_25_1717 ();
 sg13g2_decap_8 FILLER_25_1724 ();
 sg13g2_decap_8 FILLER_25_1731 ();
 sg13g2_decap_8 FILLER_25_1738 ();
 sg13g2_decap_8 FILLER_25_1745 ();
 sg13g2_decap_8 FILLER_25_1752 ();
 sg13g2_decap_8 FILLER_25_1759 ();
 sg13g2_fill_2 FILLER_25_1766 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_178 ();
 sg13g2_fill_1 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_fill_1 FILLER_26_270 ();
 sg13g2_fill_2 FILLER_26_283 ();
 sg13g2_fill_1 FILLER_26_311 ();
 sg13g2_fill_1 FILLER_26_321 ();
 sg13g2_fill_1 FILLER_26_334 ();
 sg13g2_fill_1 FILLER_26_339 ();
 sg13g2_fill_2 FILLER_26_398 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_421 ();
 sg13g2_fill_1 FILLER_26_431 ();
 sg13g2_fill_1 FILLER_26_473 ();
 sg13g2_fill_2 FILLER_26_558 ();
 sg13g2_fill_1 FILLER_26_560 ();
 sg13g2_fill_1 FILLER_26_589 ();
 sg13g2_fill_2 FILLER_26_625 ();
 sg13g2_fill_2 FILLER_26_665 ();
 sg13g2_fill_1 FILLER_26_667 ();
 sg13g2_fill_1 FILLER_26_677 ();
 sg13g2_fill_2 FILLER_26_697 ();
 sg13g2_fill_1 FILLER_26_699 ();
 sg13g2_fill_2 FILLER_26_717 ();
 sg13g2_fill_1 FILLER_26_719 ();
 sg13g2_decap_8 FILLER_26_866 ();
 sg13g2_fill_2 FILLER_26_873 ();
 sg13g2_fill_2 FILLER_26_901 ();
 sg13g2_fill_2 FILLER_26_912 ();
 sg13g2_fill_1 FILLER_26_1036 ();
 sg13g2_fill_2 FILLER_26_1059 ();
 sg13g2_fill_2 FILLER_26_1076 ();
 sg13g2_fill_1 FILLER_26_1172 ();
 sg13g2_fill_2 FILLER_26_1197 ();
 sg13g2_fill_1 FILLER_26_1203 ();
 sg13g2_fill_2 FILLER_26_1229 ();
 sg13g2_fill_1 FILLER_26_1231 ();
 sg13g2_fill_2 FILLER_26_1258 ();
 sg13g2_fill_1 FILLER_26_1260 ();
 sg13g2_fill_1 FILLER_26_1302 ();
 sg13g2_fill_2 FILLER_26_1322 ();
 sg13g2_fill_1 FILLER_26_1334 ();
 sg13g2_fill_2 FILLER_26_1339 ();
 sg13g2_fill_1 FILLER_26_1358 ();
 sg13g2_fill_2 FILLER_26_1364 ();
 sg13g2_fill_2 FILLER_26_1383 ();
 sg13g2_fill_1 FILLER_26_1385 ();
 sg13g2_fill_2 FILLER_26_1444 ();
 sg13g2_fill_2 FILLER_26_1476 ();
 sg13g2_fill_1 FILLER_26_1494 ();
 sg13g2_decap_8 FILLER_26_1542 ();
 sg13g2_decap_8 FILLER_26_1549 ();
 sg13g2_decap_8 FILLER_26_1556 ();
 sg13g2_decap_8 FILLER_26_1563 ();
 sg13g2_decap_8 FILLER_26_1570 ();
 sg13g2_decap_8 FILLER_26_1577 ();
 sg13g2_decap_8 FILLER_26_1584 ();
 sg13g2_decap_8 FILLER_26_1591 ();
 sg13g2_decap_8 FILLER_26_1598 ();
 sg13g2_decap_8 FILLER_26_1605 ();
 sg13g2_decap_8 FILLER_26_1612 ();
 sg13g2_decap_8 FILLER_26_1619 ();
 sg13g2_decap_8 FILLER_26_1626 ();
 sg13g2_decap_8 FILLER_26_1633 ();
 sg13g2_decap_8 FILLER_26_1640 ();
 sg13g2_decap_8 FILLER_26_1647 ();
 sg13g2_decap_8 FILLER_26_1654 ();
 sg13g2_decap_8 FILLER_26_1661 ();
 sg13g2_decap_8 FILLER_26_1668 ();
 sg13g2_decap_8 FILLER_26_1675 ();
 sg13g2_decap_8 FILLER_26_1682 ();
 sg13g2_decap_8 FILLER_26_1689 ();
 sg13g2_decap_8 FILLER_26_1696 ();
 sg13g2_decap_8 FILLER_26_1703 ();
 sg13g2_decap_8 FILLER_26_1710 ();
 sg13g2_decap_8 FILLER_26_1717 ();
 sg13g2_decap_8 FILLER_26_1724 ();
 sg13g2_decap_8 FILLER_26_1731 ();
 sg13g2_decap_8 FILLER_26_1738 ();
 sg13g2_decap_8 FILLER_26_1745 ();
 sg13g2_decap_8 FILLER_26_1752 ();
 sg13g2_decap_8 FILLER_26_1759 ();
 sg13g2_fill_2 FILLER_26_1766 ();
 sg13g2_fill_2 FILLER_27_26 ();
 sg13g2_fill_1 FILLER_27_37 ();
 sg13g2_fill_2 FILLER_27_87 ();
 sg13g2_fill_2 FILLER_27_106 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_1 FILLER_27_126 ();
 sg13g2_fill_2 FILLER_27_210 ();
 sg13g2_fill_1 FILLER_27_212 ();
 sg13g2_fill_2 FILLER_27_236 ();
 sg13g2_fill_1 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_244 ();
 sg13g2_fill_2 FILLER_27_262 ();
 sg13g2_fill_2 FILLER_27_289 ();
 sg13g2_fill_2 FILLER_27_333 ();
 sg13g2_fill_2 FILLER_27_375 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_fill_2 FILLER_27_438 ();
 sg13g2_fill_2 FILLER_27_466 ();
 sg13g2_fill_2 FILLER_27_498 ();
 sg13g2_fill_2 FILLER_27_526 ();
 sg13g2_fill_1 FILLER_27_627 ();
 sg13g2_fill_2 FILLER_27_644 ();
 sg13g2_fill_1 FILLER_27_646 ();
 sg13g2_fill_2 FILLER_27_652 ();
 sg13g2_fill_1 FILLER_27_654 ();
 sg13g2_fill_2 FILLER_27_661 ();
 sg13g2_fill_1 FILLER_27_697 ();
 sg13g2_fill_2 FILLER_27_728 ();
 sg13g2_fill_2 FILLER_27_764 ();
 sg13g2_fill_1 FILLER_27_809 ();
 sg13g2_fill_2 FILLER_27_874 ();
 sg13g2_fill_2 FILLER_27_881 ();
 sg13g2_fill_2 FILLER_27_896 ();
 sg13g2_fill_1 FILLER_27_912 ();
 sg13g2_fill_1 FILLER_27_937 ();
 sg13g2_fill_2 FILLER_27_958 ();
 sg13g2_fill_1 FILLER_27_960 ();
 sg13g2_fill_1 FILLER_27_969 ();
 sg13g2_fill_1 FILLER_27_1020 ();
 sg13g2_fill_2 FILLER_27_1061 ();
 sg13g2_fill_2 FILLER_27_1104 ();
 sg13g2_fill_2 FILLER_27_1177 ();
 sg13g2_fill_1 FILLER_27_1179 ();
 sg13g2_fill_1 FILLER_27_1334 ();
 sg13g2_fill_1 FILLER_27_1364 ();
 sg13g2_decap_8 FILLER_27_1545 ();
 sg13g2_decap_8 FILLER_27_1552 ();
 sg13g2_decap_8 FILLER_27_1559 ();
 sg13g2_decap_8 FILLER_27_1566 ();
 sg13g2_decap_8 FILLER_27_1573 ();
 sg13g2_decap_8 FILLER_27_1580 ();
 sg13g2_decap_8 FILLER_27_1587 ();
 sg13g2_decap_8 FILLER_27_1594 ();
 sg13g2_decap_8 FILLER_27_1601 ();
 sg13g2_decap_8 FILLER_27_1608 ();
 sg13g2_decap_8 FILLER_27_1615 ();
 sg13g2_decap_8 FILLER_27_1622 ();
 sg13g2_decap_8 FILLER_27_1629 ();
 sg13g2_decap_8 FILLER_27_1636 ();
 sg13g2_decap_8 FILLER_27_1643 ();
 sg13g2_decap_8 FILLER_27_1650 ();
 sg13g2_decap_8 FILLER_27_1657 ();
 sg13g2_decap_8 FILLER_27_1664 ();
 sg13g2_decap_8 FILLER_27_1671 ();
 sg13g2_decap_8 FILLER_27_1678 ();
 sg13g2_decap_8 FILLER_27_1685 ();
 sg13g2_decap_8 FILLER_27_1692 ();
 sg13g2_decap_8 FILLER_27_1699 ();
 sg13g2_decap_8 FILLER_27_1706 ();
 sg13g2_decap_8 FILLER_27_1713 ();
 sg13g2_decap_8 FILLER_27_1720 ();
 sg13g2_decap_8 FILLER_27_1727 ();
 sg13g2_decap_8 FILLER_27_1734 ();
 sg13g2_decap_8 FILLER_27_1741 ();
 sg13g2_decap_8 FILLER_27_1748 ();
 sg13g2_decap_8 FILLER_27_1755 ();
 sg13g2_decap_4 FILLER_27_1762 ();
 sg13g2_fill_2 FILLER_27_1766 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_fill_2 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_fill_2 FILLER_28_214 ();
 sg13g2_fill_2 FILLER_28_250 ();
 sg13g2_fill_2 FILLER_28_297 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_407 ();
 sg13g2_fill_2 FILLER_28_434 ();
 sg13g2_fill_1 FILLER_28_436 ();
 sg13g2_fill_2 FILLER_28_538 ();
 sg13g2_fill_1 FILLER_28_550 ();
 sg13g2_fill_2 FILLER_28_567 ();
 sg13g2_fill_1 FILLER_28_592 ();
 sg13g2_fill_2 FILLER_28_622 ();
 sg13g2_fill_1 FILLER_28_647 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_fill_1 FILLER_28_731 ();
 sg13g2_fill_1 FILLER_28_740 ();
 sg13g2_fill_2 FILLER_28_861 ();
 sg13g2_fill_1 FILLER_28_863 ();
 sg13g2_fill_2 FILLER_28_997 ();
 sg13g2_fill_1 FILLER_28_1009 ();
 sg13g2_fill_2 FILLER_28_1066 ();
 sg13g2_fill_1 FILLER_28_1088 ();
 sg13g2_fill_2 FILLER_28_1118 ();
 sg13g2_fill_2 FILLER_28_1158 ();
 sg13g2_fill_1 FILLER_28_1160 ();
 sg13g2_fill_2 FILLER_28_1184 ();
 sg13g2_fill_1 FILLER_28_1199 ();
 sg13g2_fill_2 FILLER_28_1213 ();
 sg13g2_fill_1 FILLER_28_1215 ();
 sg13g2_fill_2 FILLER_28_1236 ();
 sg13g2_fill_1 FILLER_28_1238 ();
 sg13g2_fill_1 FILLER_28_1265 ();
 sg13g2_fill_1 FILLER_28_1315 ();
 sg13g2_fill_2 FILLER_28_1339 ();
 sg13g2_fill_2 FILLER_28_1393 ();
 sg13g2_fill_1 FILLER_28_1395 ();
 sg13g2_fill_2 FILLER_28_1402 ();
 sg13g2_fill_1 FILLER_28_1404 ();
 sg13g2_fill_2 FILLER_28_1451 ();
 sg13g2_fill_2 FILLER_28_1477 ();
 sg13g2_fill_1 FILLER_28_1479 ();
 sg13g2_decap_8 FILLER_28_1541 ();
 sg13g2_decap_8 FILLER_28_1548 ();
 sg13g2_decap_8 FILLER_28_1555 ();
 sg13g2_decap_8 FILLER_28_1562 ();
 sg13g2_decap_8 FILLER_28_1569 ();
 sg13g2_decap_8 FILLER_28_1576 ();
 sg13g2_decap_8 FILLER_28_1583 ();
 sg13g2_decap_8 FILLER_28_1590 ();
 sg13g2_decap_8 FILLER_28_1597 ();
 sg13g2_decap_8 FILLER_28_1604 ();
 sg13g2_decap_8 FILLER_28_1611 ();
 sg13g2_decap_8 FILLER_28_1618 ();
 sg13g2_decap_8 FILLER_28_1625 ();
 sg13g2_decap_8 FILLER_28_1632 ();
 sg13g2_decap_8 FILLER_28_1639 ();
 sg13g2_decap_8 FILLER_28_1646 ();
 sg13g2_decap_8 FILLER_28_1653 ();
 sg13g2_decap_8 FILLER_28_1660 ();
 sg13g2_decap_8 FILLER_28_1667 ();
 sg13g2_decap_8 FILLER_28_1674 ();
 sg13g2_decap_8 FILLER_28_1681 ();
 sg13g2_decap_8 FILLER_28_1688 ();
 sg13g2_decap_8 FILLER_28_1695 ();
 sg13g2_decap_8 FILLER_28_1702 ();
 sg13g2_decap_8 FILLER_28_1709 ();
 sg13g2_decap_8 FILLER_28_1716 ();
 sg13g2_decap_8 FILLER_28_1723 ();
 sg13g2_decap_8 FILLER_28_1730 ();
 sg13g2_decap_8 FILLER_28_1737 ();
 sg13g2_decap_8 FILLER_28_1744 ();
 sg13g2_decap_8 FILLER_28_1751 ();
 sg13g2_decap_8 FILLER_28_1758 ();
 sg13g2_fill_2 FILLER_28_1765 ();
 sg13g2_fill_1 FILLER_28_1767 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_59 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_fill_2 FILLER_29_76 ();
 sg13g2_fill_2 FILLER_29_188 ();
 sg13g2_fill_1 FILLER_29_190 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_251 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_317 ();
 sg13g2_fill_2 FILLER_29_442 ();
 sg13g2_fill_1 FILLER_29_449 ();
 sg13g2_fill_2 FILLER_29_460 ();
 sg13g2_fill_1 FILLER_29_462 ();
 sg13g2_fill_1 FILLER_29_476 ();
 sg13g2_fill_2 FILLER_29_520 ();
 sg13g2_fill_1 FILLER_29_698 ();
 sg13g2_fill_2 FILLER_29_722 ();
 sg13g2_fill_2 FILLER_29_758 ();
 sg13g2_fill_2 FILLER_29_766 ();
 sg13g2_fill_1 FILLER_29_768 ();
 sg13g2_fill_1 FILLER_29_791 ();
 sg13g2_fill_2 FILLER_29_823 ();
 sg13g2_fill_1 FILLER_29_825 ();
 sg13g2_decap_4 FILLER_29_861 ();
 sg13g2_fill_2 FILLER_29_881 ();
 sg13g2_fill_1 FILLER_29_883 ();
 sg13g2_fill_2 FILLER_29_923 ();
 sg13g2_fill_1 FILLER_29_935 ();
 sg13g2_fill_1 FILLER_29_945 ();
 sg13g2_fill_2 FILLER_29_978 ();
 sg13g2_fill_1 FILLER_29_1207 ();
 sg13g2_fill_2 FILLER_29_1247 ();
 sg13g2_fill_1 FILLER_29_1275 ();
 sg13g2_fill_2 FILLER_29_1311 ();
 sg13g2_fill_1 FILLER_29_1366 ();
 sg13g2_fill_2 FILLER_29_1373 ();
 sg13g2_fill_1 FILLER_29_1488 ();
 sg13g2_fill_2 FILLER_29_1509 ();
 sg13g2_fill_1 FILLER_29_1511 ();
 sg13g2_decap_8 FILLER_29_1538 ();
 sg13g2_decap_8 FILLER_29_1545 ();
 sg13g2_decap_8 FILLER_29_1552 ();
 sg13g2_decap_8 FILLER_29_1559 ();
 sg13g2_decap_8 FILLER_29_1566 ();
 sg13g2_decap_8 FILLER_29_1573 ();
 sg13g2_decap_8 FILLER_29_1580 ();
 sg13g2_decap_8 FILLER_29_1587 ();
 sg13g2_decap_8 FILLER_29_1594 ();
 sg13g2_decap_8 FILLER_29_1601 ();
 sg13g2_decap_8 FILLER_29_1608 ();
 sg13g2_decap_8 FILLER_29_1615 ();
 sg13g2_decap_8 FILLER_29_1622 ();
 sg13g2_decap_8 FILLER_29_1629 ();
 sg13g2_decap_8 FILLER_29_1636 ();
 sg13g2_decap_8 FILLER_29_1643 ();
 sg13g2_decap_8 FILLER_29_1650 ();
 sg13g2_decap_8 FILLER_29_1657 ();
 sg13g2_decap_8 FILLER_29_1664 ();
 sg13g2_decap_8 FILLER_29_1671 ();
 sg13g2_decap_8 FILLER_29_1678 ();
 sg13g2_decap_8 FILLER_29_1685 ();
 sg13g2_decap_8 FILLER_29_1692 ();
 sg13g2_decap_8 FILLER_29_1699 ();
 sg13g2_decap_8 FILLER_29_1706 ();
 sg13g2_decap_8 FILLER_29_1713 ();
 sg13g2_decap_8 FILLER_29_1720 ();
 sg13g2_decap_8 FILLER_29_1727 ();
 sg13g2_decap_8 FILLER_29_1734 ();
 sg13g2_decap_8 FILLER_29_1741 ();
 sg13g2_decap_8 FILLER_29_1748 ();
 sg13g2_decap_8 FILLER_29_1755 ();
 sg13g2_decap_4 FILLER_29_1762 ();
 sg13g2_fill_2 FILLER_29_1766 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_71 ();
 sg13g2_fill_2 FILLER_30_82 ();
 sg13g2_fill_2 FILLER_30_89 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_1 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_143 ();
 sg13g2_fill_1 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_fill_2 FILLER_30_339 ();
 sg13g2_fill_2 FILLER_30_391 ();
 sg13g2_fill_2 FILLER_30_456 ();
 sg13g2_fill_1 FILLER_30_458 ();
 sg13g2_fill_1 FILLER_30_467 ();
 sg13g2_fill_2 FILLER_30_481 ();
 sg13g2_fill_1 FILLER_30_523 ();
 sg13g2_fill_2 FILLER_30_533 ();
 sg13g2_fill_1 FILLER_30_544 ();
 sg13g2_fill_2 FILLER_30_565 ();
 sg13g2_decap_8 FILLER_30_601 ();
 sg13g2_fill_1 FILLER_30_608 ();
 sg13g2_fill_1 FILLER_30_631 ();
 sg13g2_fill_1 FILLER_30_638 ();
 sg13g2_fill_1 FILLER_30_661 ();
 sg13g2_fill_2 FILLER_30_681 ();
 sg13g2_fill_1 FILLER_30_683 ();
 sg13g2_decap_4 FILLER_30_693 ();
 sg13g2_fill_1 FILLER_30_697 ();
 sg13g2_fill_2 FILLER_30_728 ();
 sg13g2_decap_4 FILLER_30_804 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_fill_2 FILLER_30_819 ();
 sg13g2_fill_1 FILLER_30_821 ();
 sg13g2_fill_2 FILLER_30_831 ();
 sg13g2_decap_8 FILLER_30_856 ();
 sg13g2_fill_2 FILLER_30_889 ();
 sg13g2_fill_1 FILLER_30_891 ();
 sg13g2_fill_1 FILLER_30_911 ();
 sg13g2_fill_1 FILLER_30_918 ();
 sg13g2_fill_2 FILLER_30_928 ();
 sg13g2_fill_2 FILLER_30_956 ();
 sg13g2_fill_1 FILLER_30_997 ();
 sg13g2_fill_1 FILLER_30_1069 ();
 sg13g2_fill_1 FILLER_30_1123 ();
 sg13g2_fill_2 FILLER_30_1176 ();
 sg13g2_fill_1 FILLER_30_1178 ();
 sg13g2_fill_1 FILLER_30_1234 ();
 sg13g2_fill_2 FILLER_30_1244 ();
 sg13g2_fill_2 FILLER_30_1281 ();
 sg13g2_fill_1 FILLER_30_1283 ();
 sg13g2_fill_2 FILLER_30_1310 ();
 sg13g2_fill_1 FILLER_30_1312 ();
 sg13g2_fill_1 FILLER_30_1426 ();
 sg13g2_fill_1 FILLER_30_1473 ();
 sg13g2_decap_8 FILLER_30_1531 ();
 sg13g2_decap_8 FILLER_30_1538 ();
 sg13g2_decap_8 FILLER_30_1545 ();
 sg13g2_decap_8 FILLER_30_1552 ();
 sg13g2_decap_8 FILLER_30_1559 ();
 sg13g2_decap_8 FILLER_30_1566 ();
 sg13g2_decap_8 FILLER_30_1573 ();
 sg13g2_decap_8 FILLER_30_1580 ();
 sg13g2_decap_8 FILLER_30_1587 ();
 sg13g2_decap_8 FILLER_30_1594 ();
 sg13g2_decap_8 FILLER_30_1601 ();
 sg13g2_decap_8 FILLER_30_1608 ();
 sg13g2_decap_8 FILLER_30_1615 ();
 sg13g2_decap_8 FILLER_30_1622 ();
 sg13g2_decap_8 FILLER_30_1629 ();
 sg13g2_decap_8 FILLER_30_1636 ();
 sg13g2_decap_8 FILLER_30_1643 ();
 sg13g2_decap_8 FILLER_30_1650 ();
 sg13g2_decap_8 FILLER_30_1657 ();
 sg13g2_decap_8 FILLER_30_1664 ();
 sg13g2_decap_8 FILLER_30_1671 ();
 sg13g2_decap_8 FILLER_30_1678 ();
 sg13g2_decap_8 FILLER_30_1685 ();
 sg13g2_decap_8 FILLER_30_1692 ();
 sg13g2_decap_8 FILLER_30_1699 ();
 sg13g2_decap_8 FILLER_30_1706 ();
 sg13g2_decap_8 FILLER_30_1713 ();
 sg13g2_decap_8 FILLER_30_1720 ();
 sg13g2_decap_8 FILLER_30_1727 ();
 sg13g2_decap_8 FILLER_30_1734 ();
 sg13g2_decap_8 FILLER_30_1741 ();
 sg13g2_decap_8 FILLER_30_1748 ();
 sg13g2_decap_8 FILLER_30_1755 ();
 sg13g2_decap_4 FILLER_30_1762 ();
 sg13g2_fill_2 FILLER_30_1766 ();
 sg13g2_fill_1 FILLER_31_67 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_fill_1 FILLER_31_111 ();
 sg13g2_fill_1 FILLER_31_203 ();
 sg13g2_fill_2 FILLER_31_236 ();
 sg13g2_fill_1 FILLER_31_316 ();
 sg13g2_fill_2 FILLER_31_469 ();
 sg13g2_fill_1 FILLER_31_493 ();
 sg13g2_fill_1 FILLER_31_542 ();
 sg13g2_fill_1 FILLER_31_549 ();
 sg13g2_fill_2 FILLER_31_564 ();
 sg13g2_fill_1 FILLER_31_575 ();
 sg13g2_fill_2 FILLER_31_585 ();
 sg13g2_fill_2 FILLER_31_640 ();
 sg13g2_fill_1 FILLER_31_642 ();
 sg13g2_fill_1 FILLER_31_669 ();
 sg13g2_fill_2 FILLER_31_717 ();
 sg13g2_fill_1 FILLER_31_719 ();
 sg13g2_fill_1 FILLER_31_726 ();
 sg13g2_fill_2 FILLER_31_753 ();
 sg13g2_fill_1 FILLER_31_755 ();
 sg13g2_fill_2 FILLER_31_770 ();
 sg13g2_fill_2 FILLER_31_780 ();
 sg13g2_fill_1 FILLER_31_782 ();
 sg13g2_fill_2 FILLER_31_845 ();
 sg13g2_fill_2 FILLER_31_886 ();
 sg13g2_fill_1 FILLER_31_897 ();
 sg13g2_fill_1 FILLER_31_913 ();
 sg13g2_fill_2 FILLER_31_944 ();
 sg13g2_fill_1 FILLER_31_946 ();
 sg13g2_fill_1 FILLER_31_956 ();
 sg13g2_fill_2 FILLER_31_966 ();
 sg13g2_decap_4 FILLER_31_1015 ();
 sg13g2_fill_1 FILLER_31_1019 ();
 sg13g2_fill_2 FILLER_31_1036 ();
 sg13g2_fill_1 FILLER_31_1064 ();
 sg13g2_fill_2 FILLER_31_1137 ();
 sg13g2_fill_1 FILLER_31_1165 ();
 sg13g2_fill_1 FILLER_31_1192 ();
 sg13g2_fill_2 FILLER_31_1208 ();
 sg13g2_fill_1 FILLER_31_1210 ();
 sg13g2_fill_1 FILLER_31_1273 ();
 sg13g2_fill_1 FILLER_31_1305 ();
 sg13g2_fill_2 FILLER_31_1332 ();
 sg13g2_fill_1 FILLER_31_1334 ();
 sg13g2_fill_2 FILLER_31_1367 ();
 sg13g2_fill_1 FILLER_31_1460 ();
 sg13g2_fill_2 FILLER_31_1487 ();
 sg13g2_decap_8 FILLER_31_1550 ();
 sg13g2_decap_8 FILLER_31_1557 ();
 sg13g2_decap_8 FILLER_31_1564 ();
 sg13g2_decap_8 FILLER_31_1571 ();
 sg13g2_decap_8 FILLER_31_1578 ();
 sg13g2_decap_8 FILLER_31_1585 ();
 sg13g2_decap_8 FILLER_31_1592 ();
 sg13g2_decap_8 FILLER_31_1599 ();
 sg13g2_decap_8 FILLER_31_1606 ();
 sg13g2_decap_8 FILLER_31_1613 ();
 sg13g2_decap_8 FILLER_31_1620 ();
 sg13g2_decap_8 FILLER_31_1627 ();
 sg13g2_decap_8 FILLER_31_1634 ();
 sg13g2_decap_8 FILLER_31_1641 ();
 sg13g2_decap_8 FILLER_31_1648 ();
 sg13g2_decap_8 FILLER_31_1655 ();
 sg13g2_decap_8 FILLER_31_1662 ();
 sg13g2_decap_8 FILLER_31_1669 ();
 sg13g2_decap_8 FILLER_31_1676 ();
 sg13g2_decap_8 FILLER_31_1683 ();
 sg13g2_decap_8 FILLER_31_1690 ();
 sg13g2_decap_8 FILLER_31_1697 ();
 sg13g2_decap_8 FILLER_31_1704 ();
 sg13g2_decap_8 FILLER_31_1711 ();
 sg13g2_decap_8 FILLER_31_1718 ();
 sg13g2_decap_8 FILLER_31_1725 ();
 sg13g2_decap_8 FILLER_31_1732 ();
 sg13g2_decap_8 FILLER_31_1739 ();
 sg13g2_decap_8 FILLER_31_1746 ();
 sg13g2_decap_8 FILLER_31_1753 ();
 sg13g2_decap_8 FILLER_31_1760 ();
 sg13g2_fill_1 FILLER_31_1767 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_41 ();
 sg13g2_fill_2 FILLER_32_57 ();
 sg13g2_fill_1 FILLER_32_59 ();
 sg13g2_fill_1 FILLER_32_72 ();
 sg13g2_fill_1 FILLER_32_83 ();
 sg13g2_fill_2 FILLER_32_97 ();
 sg13g2_fill_1 FILLER_32_99 ();
 sg13g2_fill_2 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_130 ();
 sg13g2_fill_2 FILLER_32_152 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_fill_1 FILLER_32_228 ();
 sg13g2_fill_2 FILLER_32_234 ();
 sg13g2_fill_2 FILLER_32_241 ();
 sg13g2_fill_1 FILLER_32_243 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_fill_2 FILLER_32_286 ();
 sg13g2_fill_1 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_fill_2 FILLER_32_368 ();
 sg13g2_fill_2 FILLER_32_438 ();
 sg13g2_fill_2 FILLER_32_495 ();
 sg13g2_fill_1 FILLER_32_518 ();
 sg13g2_fill_2 FILLER_32_585 ();
 sg13g2_fill_1 FILLER_32_587 ();
 sg13g2_fill_2 FILLER_32_668 ();
 sg13g2_decap_4 FILLER_32_681 ();
 sg13g2_fill_1 FILLER_32_787 ();
 sg13g2_fill_2 FILLER_32_797 ();
 sg13g2_fill_2 FILLER_32_816 ();
 sg13g2_decap_8 FILLER_32_822 ();
 sg13g2_fill_1 FILLER_32_829 ();
 sg13g2_decap_8 FILLER_32_834 ();
 sg13g2_fill_2 FILLER_32_841 ();
 sg13g2_fill_2 FILLER_32_878 ();
 sg13g2_fill_1 FILLER_32_880 ();
 sg13g2_fill_2 FILLER_32_916 ();
 sg13g2_fill_1 FILLER_32_918 ();
 sg13g2_fill_1 FILLER_32_927 ();
 sg13g2_fill_2 FILLER_32_968 ();
 sg13g2_fill_2 FILLER_32_975 ();
 sg13g2_fill_1 FILLER_32_977 ();
 sg13g2_fill_1 FILLER_32_991 ();
 sg13g2_fill_1 FILLER_32_1007 ();
 sg13g2_fill_1 FILLER_32_1079 ();
 sg13g2_fill_2 FILLER_32_1090 ();
 sg13g2_fill_1 FILLER_32_1109 ();
 sg13g2_fill_1 FILLER_32_1119 ();
 sg13g2_fill_2 FILLER_32_1224 ();
 sg13g2_fill_1 FILLER_32_1226 ();
 sg13g2_fill_2 FILLER_32_1261 ();
 sg13g2_fill_1 FILLER_32_1263 ();
 sg13g2_fill_2 FILLER_32_1318 ();
 sg13g2_fill_1 FILLER_32_1320 ();
 sg13g2_fill_1 FILLER_32_1363 ();
 sg13g2_fill_2 FILLER_32_1374 ();
 sg13g2_fill_1 FILLER_32_1376 ();
 sg13g2_fill_1 FILLER_32_1411 ();
 sg13g2_fill_2 FILLER_32_1452 ();
 sg13g2_fill_1 FILLER_32_1454 ();
 sg13g2_fill_1 FILLER_32_1477 ();
 sg13g2_decap_4 FILLER_32_1487 ();
 sg13g2_fill_2 FILLER_32_1505 ();
 sg13g2_fill_2 FILLER_32_1524 ();
 sg13g2_fill_1 FILLER_32_1526 ();
 sg13g2_decap_8 FILLER_32_1544 ();
 sg13g2_decap_8 FILLER_32_1551 ();
 sg13g2_decap_8 FILLER_32_1558 ();
 sg13g2_decap_8 FILLER_32_1565 ();
 sg13g2_decap_8 FILLER_32_1572 ();
 sg13g2_decap_8 FILLER_32_1579 ();
 sg13g2_decap_8 FILLER_32_1586 ();
 sg13g2_decap_8 FILLER_32_1593 ();
 sg13g2_decap_8 FILLER_32_1600 ();
 sg13g2_decap_8 FILLER_32_1607 ();
 sg13g2_decap_8 FILLER_32_1614 ();
 sg13g2_decap_8 FILLER_32_1621 ();
 sg13g2_decap_8 FILLER_32_1628 ();
 sg13g2_decap_8 FILLER_32_1635 ();
 sg13g2_decap_8 FILLER_32_1642 ();
 sg13g2_decap_8 FILLER_32_1649 ();
 sg13g2_decap_8 FILLER_32_1656 ();
 sg13g2_decap_8 FILLER_32_1663 ();
 sg13g2_decap_8 FILLER_32_1670 ();
 sg13g2_decap_8 FILLER_32_1677 ();
 sg13g2_decap_8 FILLER_32_1684 ();
 sg13g2_decap_8 FILLER_32_1691 ();
 sg13g2_decap_8 FILLER_32_1698 ();
 sg13g2_decap_8 FILLER_32_1705 ();
 sg13g2_decap_8 FILLER_32_1712 ();
 sg13g2_decap_8 FILLER_32_1719 ();
 sg13g2_decap_8 FILLER_32_1726 ();
 sg13g2_decap_8 FILLER_32_1733 ();
 sg13g2_decap_8 FILLER_32_1740 ();
 sg13g2_decap_8 FILLER_32_1747 ();
 sg13g2_decap_8 FILLER_32_1754 ();
 sg13g2_decap_8 FILLER_32_1761 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_fill_1 FILLER_33_36 ();
 sg13g2_fill_1 FILLER_33_115 ();
 sg13g2_fill_1 FILLER_33_139 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_321 ();
 sg13g2_fill_2 FILLER_33_348 ();
 sg13g2_fill_1 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_410 ();
 sg13g2_fill_2 FILLER_33_417 ();
 sg13g2_fill_2 FILLER_33_467 ();
 sg13g2_fill_1 FILLER_33_561 ();
 sg13g2_fill_2 FILLER_33_579 ();
 sg13g2_fill_2 FILLER_33_595 ();
 sg13g2_fill_2 FILLER_33_629 ();
 sg13g2_fill_2 FILLER_33_637 ();
 sg13g2_fill_2 FILLER_33_772 ();
 sg13g2_fill_1 FILLER_33_774 ();
 sg13g2_fill_2 FILLER_33_831 ();
 sg13g2_fill_2 FILLER_33_846 ();
 sg13g2_fill_2 FILLER_33_878 ();
 sg13g2_fill_2 FILLER_33_894 ();
 sg13g2_fill_2 FILLER_33_968 ();
 sg13g2_fill_2 FILLER_33_982 ();
 sg13g2_fill_1 FILLER_33_984 ();
 sg13g2_decap_8 FILLER_33_1011 ();
 sg13g2_fill_2 FILLER_33_1018 ();
 sg13g2_decap_4 FILLER_33_1028 ();
 sg13g2_fill_2 FILLER_33_1032 ();
 sg13g2_fill_2 FILLER_33_1056 ();
 sg13g2_fill_1 FILLER_33_1058 ();
 sg13g2_fill_2 FILLER_33_1069 ();
 sg13g2_fill_2 FILLER_33_1085 ();
 sg13g2_fill_1 FILLER_33_1117 ();
 sg13g2_fill_2 FILLER_33_1201 ();
 sg13g2_fill_1 FILLER_33_1203 ();
 sg13g2_fill_1 FILLER_33_1218 ();
 sg13g2_fill_2 FILLER_33_1231 ();
 sg13g2_fill_1 FILLER_33_1233 ();
 sg13g2_fill_1 FILLER_33_1276 ();
 sg13g2_fill_1 FILLER_33_1289 ();
 sg13g2_fill_2 FILLER_33_1295 ();
 sg13g2_fill_2 FILLER_33_1313 ();
 sg13g2_fill_2 FILLER_33_1320 ();
 sg13g2_fill_2 FILLER_33_1345 ();
 sg13g2_fill_1 FILLER_33_1347 ();
 sg13g2_fill_1 FILLER_33_1365 ();
 sg13g2_fill_1 FILLER_33_1412 ();
 sg13g2_fill_2 FILLER_33_1421 ();
 sg13g2_decap_4 FILLER_33_1429 ();
 sg13g2_fill_1 FILLER_33_1433 ();
 sg13g2_fill_1 FILLER_33_1473 ();
 sg13g2_fill_1 FILLER_33_1520 ();
 sg13g2_decap_8 FILLER_33_1547 ();
 sg13g2_decap_8 FILLER_33_1554 ();
 sg13g2_decap_8 FILLER_33_1561 ();
 sg13g2_decap_8 FILLER_33_1568 ();
 sg13g2_decap_8 FILLER_33_1575 ();
 sg13g2_decap_8 FILLER_33_1582 ();
 sg13g2_decap_8 FILLER_33_1589 ();
 sg13g2_decap_8 FILLER_33_1596 ();
 sg13g2_decap_8 FILLER_33_1603 ();
 sg13g2_decap_8 FILLER_33_1610 ();
 sg13g2_decap_8 FILLER_33_1617 ();
 sg13g2_decap_8 FILLER_33_1624 ();
 sg13g2_decap_8 FILLER_33_1631 ();
 sg13g2_decap_8 FILLER_33_1638 ();
 sg13g2_decap_8 FILLER_33_1645 ();
 sg13g2_decap_8 FILLER_33_1652 ();
 sg13g2_decap_8 FILLER_33_1659 ();
 sg13g2_decap_8 FILLER_33_1666 ();
 sg13g2_decap_8 FILLER_33_1673 ();
 sg13g2_decap_8 FILLER_33_1680 ();
 sg13g2_decap_8 FILLER_33_1687 ();
 sg13g2_decap_8 FILLER_33_1694 ();
 sg13g2_decap_8 FILLER_33_1701 ();
 sg13g2_decap_8 FILLER_33_1708 ();
 sg13g2_decap_8 FILLER_33_1715 ();
 sg13g2_decap_8 FILLER_33_1722 ();
 sg13g2_decap_8 FILLER_33_1729 ();
 sg13g2_decap_8 FILLER_33_1736 ();
 sg13g2_decap_8 FILLER_33_1743 ();
 sg13g2_decap_8 FILLER_33_1750 ();
 sg13g2_decap_8 FILLER_33_1757 ();
 sg13g2_decap_4 FILLER_33_1764 ();
 sg13g2_fill_2 FILLER_34_25 ();
 sg13g2_fill_1 FILLER_34_27 ();
 sg13g2_fill_1 FILLER_34_43 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_82 ();
 sg13g2_fill_2 FILLER_34_87 ();
 sg13g2_fill_1 FILLER_34_89 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_fill_1 FILLER_34_109 ();
 sg13g2_fill_1 FILLER_34_162 ();
 sg13g2_fill_2 FILLER_34_189 ();
 sg13g2_fill_2 FILLER_34_195 ();
 sg13g2_fill_1 FILLER_34_197 ();
 sg13g2_fill_2 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_215 ();
 sg13g2_fill_2 FILLER_34_224 ();
 sg13g2_fill_1 FILLER_34_226 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_fill_1 FILLER_34_305 ();
 sg13g2_fill_1 FILLER_34_315 ();
 sg13g2_fill_2 FILLER_34_321 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_2 FILLER_34_339 ();
 sg13g2_fill_2 FILLER_34_372 ();
 sg13g2_fill_1 FILLER_34_392 ();
 sg13g2_fill_1 FILLER_34_401 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_fill_2 FILLER_34_417 ();
 sg13g2_fill_1 FILLER_34_419 ();
 sg13g2_fill_2 FILLER_34_449 ();
 sg13g2_fill_1 FILLER_34_451 ();
 sg13g2_fill_2 FILLER_34_470 ();
 sg13g2_fill_1 FILLER_34_472 ();
 sg13g2_fill_2 FILLER_34_486 ();
 sg13g2_fill_1 FILLER_34_488 ();
 sg13g2_fill_2 FILLER_34_506 ();
 sg13g2_fill_1 FILLER_34_508 ();
 sg13g2_fill_2 FILLER_34_573 ();
 sg13g2_fill_1 FILLER_34_575 ();
 sg13g2_fill_1 FILLER_34_602 ();
 sg13g2_fill_1 FILLER_34_638 ();
 sg13g2_fill_2 FILLER_34_661 ();
 sg13g2_fill_1 FILLER_34_663 ();
 sg13g2_fill_1 FILLER_34_704 ();
 sg13g2_fill_1 FILLER_34_734 ();
 sg13g2_fill_1 FILLER_34_761 ();
 sg13g2_fill_1 FILLER_34_775 ();
 sg13g2_fill_2 FILLER_34_803 ();
 sg13g2_fill_1 FILLER_34_805 ();
 sg13g2_fill_2 FILLER_34_815 ();
 sg13g2_fill_2 FILLER_34_821 ();
 sg13g2_fill_2 FILLER_34_874 ();
 sg13g2_fill_1 FILLER_34_876 ();
 sg13g2_fill_1 FILLER_34_903 ();
 sg13g2_fill_1 FILLER_34_912 ();
 sg13g2_fill_2 FILLER_34_955 ();
 sg13g2_fill_1 FILLER_34_957 ();
 sg13g2_fill_2 FILLER_34_1026 ();
 sg13g2_fill_2 FILLER_34_1032 ();
 sg13g2_fill_1 FILLER_34_1159 ();
 sg13g2_fill_1 FILLER_34_1201 ();
 sg13g2_fill_2 FILLER_34_1215 ();
 sg13g2_fill_2 FILLER_34_1222 ();
 sg13g2_fill_1 FILLER_34_1224 ();
 sg13g2_fill_2 FILLER_34_1269 ();
 sg13g2_fill_1 FILLER_34_1271 ();
 sg13g2_fill_2 FILLER_34_1291 ();
 sg13g2_fill_1 FILLER_34_1293 ();
 sg13g2_fill_2 FILLER_34_1370 ();
 sg13g2_fill_1 FILLER_34_1372 ();
 sg13g2_fill_1 FILLER_34_1387 ();
 sg13g2_fill_1 FILLER_34_1406 ();
 sg13g2_fill_1 FILLER_34_1438 ();
 sg13g2_fill_1 FILLER_34_1443 ();
 sg13g2_decap_8 FILLER_34_1544 ();
 sg13g2_decap_8 FILLER_34_1551 ();
 sg13g2_decap_8 FILLER_34_1558 ();
 sg13g2_decap_8 FILLER_34_1565 ();
 sg13g2_decap_8 FILLER_34_1572 ();
 sg13g2_decap_8 FILLER_34_1579 ();
 sg13g2_decap_8 FILLER_34_1586 ();
 sg13g2_decap_8 FILLER_34_1593 ();
 sg13g2_decap_8 FILLER_34_1600 ();
 sg13g2_decap_8 FILLER_34_1607 ();
 sg13g2_decap_8 FILLER_34_1614 ();
 sg13g2_decap_8 FILLER_34_1621 ();
 sg13g2_decap_8 FILLER_34_1628 ();
 sg13g2_decap_8 FILLER_34_1635 ();
 sg13g2_decap_8 FILLER_34_1642 ();
 sg13g2_decap_8 FILLER_34_1649 ();
 sg13g2_decap_8 FILLER_34_1656 ();
 sg13g2_decap_8 FILLER_34_1663 ();
 sg13g2_decap_8 FILLER_34_1670 ();
 sg13g2_decap_8 FILLER_34_1677 ();
 sg13g2_decap_8 FILLER_34_1684 ();
 sg13g2_decap_8 FILLER_34_1691 ();
 sg13g2_decap_8 FILLER_34_1698 ();
 sg13g2_decap_8 FILLER_34_1705 ();
 sg13g2_decap_8 FILLER_34_1712 ();
 sg13g2_decap_8 FILLER_34_1719 ();
 sg13g2_decap_8 FILLER_34_1726 ();
 sg13g2_decap_8 FILLER_34_1733 ();
 sg13g2_decap_8 FILLER_34_1740 ();
 sg13g2_decap_8 FILLER_34_1747 ();
 sg13g2_decap_8 FILLER_34_1754 ();
 sg13g2_decap_8 FILLER_34_1761 ();
 sg13g2_fill_1 FILLER_35_26 ();
 sg13g2_fill_1 FILLER_35_57 ();
 sg13g2_fill_1 FILLER_35_71 ();
 sg13g2_fill_1 FILLER_35_86 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_fill_1 FILLER_35_119 ();
 sg13g2_fill_2 FILLER_35_138 ();
 sg13g2_fill_2 FILLER_35_148 ();
 sg13g2_fill_1 FILLER_35_150 ();
 sg13g2_fill_1 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_190 ();
 sg13g2_fill_2 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_fill_2 FILLER_35_251 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_fill_1 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_333 ();
 sg13g2_fill_1 FILLER_35_335 ();
 sg13g2_fill_1 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_408 ();
 sg13g2_fill_1 FILLER_35_410 ();
 sg13g2_fill_2 FILLER_35_478 ();
 sg13g2_fill_1 FILLER_35_480 ();
 sg13g2_fill_1 FILLER_35_494 ();
 sg13g2_fill_2 FILLER_35_511 ();
 sg13g2_fill_2 FILLER_35_521 ();
 sg13g2_fill_1 FILLER_35_523 ();
 sg13g2_fill_2 FILLER_35_533 ();
 sg13g2_fill_1 FILLER_35_535 ();
 sg13g2_fill_2 FILLER_35_569 ();
 sg13g2_fill_1 FILLER_35_571 ();
 sg13g2_fill_2 FILLER_35_608 ();
 sg13g2_fill_2 FILLER_35_663 ();
 sg13g2_fill_1 FILLER_35_665 ();
 sg13g2_fill_2 FILLER_35_690 ();
 sg13g2_fill_1 FILLER_35_724 ();
 sg13g2_fill_2 FILLER_35_803 ();
 sg13g2_fill_1 FILLER_35_805 ();
 sg13g2_fill_2 FILLER_35_852 ();
 sg13g2_fill_2 FILLER_35_928 ();
 sg13g2_fill_1 FILLER_35_930 ();
 sg13g2_fill_2 FILLER_35_969 ();
 sg13g2_fill_1 FILLER_35_971 ();
 sg13g2_fill_1 FILLER_35_1016 ();
 sg13g2_fill_2 FILLER_35_1052 ();
 sg13g2_fill_2 FILLER_35_1081 ();
 sg13g2_fill_1 FILLER_35_1083 ();
 sg13g2_fill_1 FILLER_35_1089 ();
 sg13g2_fill_1 FILLER_35_1126 ();
 sg13g2_decap_8 FILLER_35_1131 ();
 sg13g2_fill_2 FILLER_35_1143 ();
 sg13g2_fill_1 FILLER_35_1145 ();
 sg13g2_fill_2 FILLER_35_1154 ();
 sg13g2_fill_1 FILLER_35_1156 ();
 sg13g2_decap_4 FILLER_35_1162 ();
 sg13g2_fill_2 FILLER_35_1197 ();
 sg13g2_fill_1 FILLER_35_1234 ();
 sg13g2_fill_2 FILLER_35_1310 ();
 sg13g2_fill_1 FILLER_35_1312 ();
 sg13g2_fill_2 FILLER_35_1322 ();
 sg13g2_fill_2 FILLER_35_1344 ();
 sg13g2_fill_1 FILLER_35_1346 ();
 sg13g2_fill_2 FILLER_35_1383 ();
 sg13g2_fill_2 FILLER_35_1420 ();
 sg13g2_fill_1 FILLER_35_1443 ();
 sg13g2_fill_1 FILLER_35_1478 ();
 sg13g2_fill_2 FILLER_35_1489 ();
 sg13g2_fill_2 FILLER_35_1511 ();
 sg13g2_fill_1 FILLER_35_1513 ();
 sg13g2_decap_8 FILLER_35_1540 ();
 sg13g2_decap_8 FILLER_35_1547 ();
 sg13g2_decap_8 FILLER_35_1554 ();
 sg13g2_decap_8 FILLER_35_1561 ();
 sg13g2_decap_8 FILLER_35_1568 ();
 sg13g2_decap_8 FILLER_35_1575 ();
 sg13g2_decap_8 FILLER_35_1582 ();
 sg13g2_decap_8 FILLER_35_1589 ();
 sg13g2_decap_8 FILLER_35_1596 ();
 sg13g2_decap_8 FILLER_35_1603 ();
 sg13g2_decap_8 FILLER_35_1610 ();
 sg13g2_decap_8 FILLER_35_1617 ();
 sg13g2_decap_8 FILLER_35_1624 ();
 sg13g2_decap_8 FILLER_35_1631 ();
 sg13g2_decap_8 FILLER_35_1638 ();
 sg13g2_decap_8 FILLER_35_1645 ();
 sg13g2_decap_8 FILLER_35_1652 ();
 sg13g2_decap_8 FILLER_35_1659 ();
 sg13g2_decap_8 FILLER_35_1666 ();
 sg13g2_decap_8 FILLER_35_1673 ();
 sg13g2_decap_8 FILLER_35_1680 ();
 sg13g2_decap_8 FILLER_35_1687 ();
 sg13g2_decap_8 FILLER_35_1694 ();
 sg13g2_decap_8 FILLER_35_1701 ();
 sg13g2_decap_8 FILLER_35_1708 ();
 sg13g2_decap_8 FILLER_35_1715 ();
 sg13g2_decap_8 FILLER_35_1722 ();
 sg13g2_decap_8 FILLER_35_1729 ();
 sg13g2_decap_8 FILLER_35_1736 ();
 sg13g2_decap_8 FILLER_35_1743 ();
 sg13g2_decap_8 FILLER_35_1750 ();
 sg13g2_decap_8 FILLER_35_1757 ();
 sg13g2_decap_4 FILLER_35_1764 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_35 ();
 sg13g2_fill_1 FILLER_36_37 ();
 sg13g2_fill_2 FILLER_36_211 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_298 ();
 sg13g2_fill_2 FILLER_36_305 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_329 ();
 sg13g2_fill_2 FILLER_36_336 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_fill_2 FILLER_36_443 ();
 sg13g2_fill_1 FILLER_36_460 ();
 sg13g2_fill_1 FILLER_36_503 ();
 sg13g2_fill_1 FILLER_36_512 ();
 sg13g2_fill_1 FILLER_36_548 ();
 sg13g2_fill_2 FILLER_36_575 ();
 sg13g2_fill_2 FILLER_36_591 ();
 sg13g2_fill_1 FILLER_36_602 ();
 sg13g2_fill_2 FILLER_36_615 ();
 sg13g2_fill_1 FILLER_36_617 ();
 sg13g2_fill_1 FILLER_36_629 ();
 sg13g2_fill_1 FILLER_36_721 ();
 sg13g2_fill_2 FILLER_36_732 ();
 sg13g2_fill_1 FILLER_36_759 ();
 sg13g2_fill_2 FILLER_36_830 ();
 sg13g2_fill_1 FILLER_36_832 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_fill_2 FILLER_36_872 ();
 sg13g2_decap_8 FILLER_36_897 ();
 sg13g2_fill_1 FILLER_36_904 ();
 sg13g2_fill_2 FILLER_36_910 ();
 sg13g2_fill_1 FILLER_36_912 ();
 sg13g2_decap_4 FILLER_36_917 ();
 sg13g2_decap_4 FILLER_36_925 ();
 sg13g2_fill_2 FILLER_36_929 ();
 sg13g2_fill_2 FILLER_36_941 ();
 sg13g2_fill_1 FILLER_36_1026 ();
 sg13g2_fill_1 FILLER_36_1062 ();
 sg13g2_fill_2 FILLER_36_1104 ();
 sg13g2_fill_1 FILLER_36_1132 ();
 sg13g2_fill_2 FILLER_36_1219 ();
 sg13g2_fill_1 FILLER_36_1221 ();
 sg13g2_fill_2 FILLER_36_1266 ();
 sg13g2_fill_2 FILLER_36_1280 ();
 sg13g2_fill_1 FILLER_36_1282 ();
 sg13g2_fill_1 FILLER_36_1359 ();
 sg13g2_fill_1 FILLER_36_1388 ();
 sg13g2_fill_1 FILLER_36_1398 ();
 sg13g2_fill_1 FILLER_36_1402 ();
 sg13g2_fill_2 FILLER_36_1423 ();
 sg13g2_fill_2 FILLER_36_1511 ();
 sg13g2_fill_1 FILLER_36_1513 ();
 sg13g2_decap_8 FILLER_36_1540 ();
 sg13g2_decap_8 FILLER_36_1547 ();
 sg13g2_decap_8 FILLER_36_1554 ();
 sg13g2_decap_8 FILLER_36_1561 ();
 sg13g2_decap_8 FILLER_36_1568 ();
 sg13g2_decap_8 FILLER_36_1575 ();
 sg13g2_decap_8 FILLER_36_1582 ();
 sg13g2_decap_8 FILLER_36_1589 ();
 sg13g2_decap_8 FILLER_36_1596 ();
 sg13g2_decap_8 FILLER_36_1603 ();
 sg13g2_decap_8 FILLER_36_1610 ();
 sg13g2_decap_8 FILLER_36_1617 ();
 sg13g2_decap_8 FILLER_36_1624 ();
 sg13g2_decap_8 FILLER_36_1631 ();
 sg13g2_decap_8 FILLER_36_1638 ();
 sg13g2_decap_8 FILLER_36_1645 ();
 sg13g2_decap_8 FILLER_36_1652 ();
 sg13g2_decap_8 FILLER_36_1659 ();
 sg13g2_decap_8 FILLER_36_1666 ();
 sg13g2_decap_8 FILLER_36_1673 ();
 sg13g2_decap_8 FILLER_36_1680 ();
 sg13g2_decap_8 FILLER_36_1687 ();
 sg13g2_decap_8 FILLER_36_1694 ();
 sg13g2_decap_8 FILLER_36_1701 ();
 sg13g2_decap_8 FILLER_36_1708 ();
 sg13g2_decap_8 FILLER_36_1715 ();
 sg13g2_decap_8 FILLER_36_1722 ();
 sg13g2_decap_8 FILLER_36_1729 ();
 sg13g2_decap_8 FILLER_36_1736 ();
 sg13g2_decap_8 FILLER_36_1743 ();
 sg13g2_decap_8 FILLER_36_1750 ();
 sg13g2_decap_8 FILLER_36_1757 ();
 sg13g2_decap_4 FILLER_36_1764 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_51 ();
 sg13g2_fill_1 FILLER_37_73 ();
 sg13g2_fill_2 FILLER_37_88 ();
 sg13g2_fill_2 FILLER_37_138 ();
 sg13g2_fill_1 FILLER_37_140 ();
 sg13g2_fill_2 FILLER_37_164 ();
 sg13g2_fill_2 FILLER_37_180 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_fill_2 FILLER_37_221 ();
 sg13g2_fill_2 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_1 FILLER_37_297 ();
 sg13g2_fill_2 FILLER_37_354 ();
 sg13g2_fill_1 FILLER_37_356 ();
 sg13g2_fill_1 FILLER_37_383 ();
 sg13g2_decap_4 FILLER_37_414 ();
 sg13g2_fill_1 FILLER_37_418 ();
 sg13g2_fill_1 FILLER_37_459 ();
 sg13g2_fill_2 FILLER_37_469 ();
 sg13g2_fill_1 FILLER_37_471 ();
 sg13g2_fill_2 FILLER_37_504 ();
 sg13g2_fill_2 FILLER_37_514 ();
 sg13g2_fill_1 FILLER_37_516 ();
 sg13g2_fill_1 FILLER_37_534 ();
 sg13g2_fill_2 FILLER_37_550 ();
 sg13g2_fill_1 FILLER_37_566 ();
 sg13g2_fill_1 FILLER_37_694 ();
 sg13g2_fill_2 FILLER_37_712 ();
 sg13g2_fill_2 FILLER_37_720 ();
 sg13g2_decap_4 FILLER_37_748 ();
 sg13g2_fill_2 FILLER_37_795 ();
 sg13g2_fill_1 FILLER_37_807 ();
 sg13g2_fill_1 FILLER_37_848 ();
 sg13g2_fill_1 FILLER_37_863 ();
 sg13g2_fill_1 FILLER_37_895 ();
 sg13g2_fill_2 FILLER_37_904 ();
 sg13g2_fill_2 FILLER_37_914 ();
 sg13g2_fill_1 FILLER_37_916 ();
 sg13g2_fill_2 FILLER_37_923 ();
 sg13g2_fill_2 FILLER_37_951 ();
 sg13g2_fill_1 FILLER_37_953 ();
 sg13g2_fill_2 FILLER_37_968 ();
 sg13g2_fill_1 FILLER_37_970 ();
 sg13g2_fill_2 FILLER_37_976 ();
 sg13g2_fill_2 FILLER_37_991 ();
 sg13g2_fill_2 FILLER_37_1002 ();
 sg13g2_fill_1 FILLER_37_1004 ();
 sg13g2_fill_2 FILLER_37_1055 ();
 sg13g2_decap_4 FILLER_37_1154 ();
 sg13g2_fill_2 FILLER_37_1211 ();
 sg13g2_fill_1 FILLER_37_1213 ();
 sg13g2_fill_1 FILLER_37_1225 ();
 sg13g2_fill_1 FILLER_37_1277 ();
 sg13g2_fill_2 FILLER_37_1292 ();
 sg13g2_fill_2 FILLER_37_1300 ();
 sg13g2_fill_1 FILLER_37_1302 ();
 sg13g2_fill_2 FILLER_37_1322 ();
 sg13g2_fill_1 FILLER_37_1324 ();
 sg13g2_fill_2 FILLER_37_1351 ();
 sg13g2_fill_1 FILLER_37_1353 ();
 sg13g2_fill_2 FILLER_37_1421 ();
 sg13g2_decap_8 FILLER_37_1427 ();
 sg13g2_fill_2 FILLER_37_1447 ();
 sg13g2_fill_1 FILLER_37_1449 ();
 sg13g2_fill_2 FILLER_37_1485 ();
 sg13g2_decap_8 FILLER_37_1545 ();
 sg13g2_decap_8 FILLER_37_1552 ();
 sg13g2_decap_8 FILLER_37_1559 ();
 sg13g2_decap_8 FILLER_37_1566 ();
 sg13g2_decap_8 FILLER_37_1573 ();
 sg13g2_decap_8 FILLER_37_1580 ();
 sg13g2_decap_8 FILLER_37_1587 ();
 sg13g2_decap_8 FILLER_37_1594 ();
 sg13g2_decap_8 FILLER_37_1601 ();
 sg13g2_decap_8 FILLER_37_1608 ();
 sg13g2_decap_8 FILLER_37_1615 ();
 sg13g2_decap_8 FILLER_37_1622 ();
 sg13g2_decap_8 FILLER_37_1629 ();
 sg13g2_decap_8 FILLER_37_1636 ();
 sg13g2_decap_8 FILLER_37_1643 ();
 sg13g2_decap_8 FILLER_37_1650 ();
 sg13g2_decap_8 FILLER_37_1657 ();
 sg13g2_decap_8 FILLER_37_1664 ();
 sg13g2_decap_8 FILLER_37_1671 ();
 sg13g2_decap_8 FILLER_37_1678 ();
 sg13g2_decap_8 FILLER_37_1685 ();
 sg13g2_decap_8 FILLER_37_1692 ();
 sg13g2_decap_8 FILLER_37_1699 ();
 sg13g2_decap_8 FILLER_37_1706 ();
 sg13g2_decap_8 FILLER_37_1713 ();
 sg13g2_decap_8 FILLER_37_1720 ();
 sg13g2_decap_8 FILLER_37_1727 ();
 sg13g2_decap_8 FILLER_37_1734 ();
 sg13g2_decap_8 FILLER_37_1741 ();
 sg13g2_decap_8 FILLER_37_1748 ();
 sg13g2_decap_8 FILLER_37_1755 ();
 sg13g2_decap_4 FILLER_37_1762 ();
 sg13g2_fill_2 FILLER_37_1766 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_69 ();
 sg13g2_fill_1 FILLER_38_71 ();
 sg13g2_fill_2 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_281 ();
 sg13g2_fill_1 FILLER_38_283 ();
 sg13g2_fill_1 FILLER_38_289 ();
 sg13g2_fill_2 FILLER_38_314 ();
 sg13g2_fill_1 FILLER_38_316 ();
 sg13g2_fill_2 FILLER_38_348 ();
 sg13g2_fill_1 FILLER_38_350 ();
 sg13g2_fill_2 FILLER_38_476 ();
 sg13g2_fill_1 FILLER_38_478 ();
 sg13g2_fill_2 FILLER_38_505 ();
 sg13g2_fill_1 FILLER_38_507 ();
 sg13g2_fill_1 FILLER_38_598 ();
 sg13g2_fill_2 FILLER_38_608 ();
 sg13g2_fill_1 FILLER_38_610 ();
 sg13g2_fill_2 FILLER_38_629 ();
 sg13g2_fill_1 FILLER_38_645 ();
 sg13g2_fill_1 FILLER_38_655 ();
 sg13g2_fill_1 FILLER_38_680 ();
 sg13g2_decap_4 FILLER_38_742 ();
 sg13g2_fill_2 FILLER_38_746 ();
 sg13g2_fill_1 FILLER_38_783 ();
 sg13g2_fill_2 FILLER_38_825 ();
 sg13g2_fill_2 FILLER_38_884 ();
 sg13g2_fill_2 FILLER_38_938 ();
 sg13g2_fill_2 FILLER_38_960 ();
 sg13g2_fill_1 FILLER_38_962 ();
 sg13g2_fill_2 FILLER_38_975 ();
 sg13g2_fill_1 FILLER_38_1045 ();
 sg13g2_fill_2 FILLER_38_1060 ();
 sg13g2_fill_1 FILLER_38_1078 ();
 sg13g2_fill_1 FILLER_38_1085 ();
 sg13g2_fill_1 FILLER_38_1100 ();
 sg13g2_fill_1 FILLER_38_1126 ();
 sg13g2_fill_2 FILLER_38_1136 ();
 sg13g2_fill_1 FILLER_38_1138 ();
 sg13g2_fill_1 FILLER_38_1150 ();
 sg13g2_fill_2 FILLER_38_1164 ();
 sg13g2_fill_1 FILLER_38_1171 ();
 sg13g2_fill_2 FILLER_38_1190 ();
 sg13g2_fill_1 FILLER_38_1192 ();
 sg13g2_fill_1 FILLER_38_1228 ();
 sg13g2_fill_2 FILLER_38_1239 ();
 sg13g2_fill_1 FILLER_38_1319 ();
 sg13g2_fill_2 FILLER_38_1332 ();
 sg13g2_fill_1 FILLER_38_1374 ();
 sg13g2_fill_2 FILLER_38_1380 ();
 sg13g2_fill_1 FILLER_38_1413 ();
 sg13g2_decap_8 FILLER_38_1424 ();
 sg13g2_fill_2 FILLER_38_1431 ();
 sg13g2_decap_8 FILLER_38_1437 ();
 sg13g2_fill_2 FILLER_38_1444 ();
 sg13g2_fill_2 FILLER_38_1451 ();
 sg13g2_fill_1 FILLER_38_1457 ();
 sg13g2_fill_2 FILLER_38_1496 ();
 sg13g2_fill_1 FILLER_38_1498 ();
 sg13g2_fill_2 FILLER_38_1517 ();
 sg13g2_fill_1 FILLER_38_1519 ();
 sg13g2_decap_8 FILLER_38_1546 ();
 sg13g2_decap_8 FILLER_38_1553 ();
 sg13g2_decap_8 FILLER_38_1560 ();
 sg13g2_decap_8 FILLER_38_1567 ();
 sg13g2_decap_8 FILLER_38_1574 ();
 sg13g2_decap_8 FILLER_38_1581 ();
 sg13g2_decap_8 FILLER_38_1588 ();
 sg13g2_decap_8 FILLER_38_1595 ();
 sg13g2_decap_8 FILLER_38_1602 ();
 sg13g2_decap_8 FILLER_38_1609 ();
 sg13g2_decap_8 FILLER_38_1616 ();
 sg13g2_decap_8 FILLER_38_1623 ();
 sg13g2_decap_8 FILLER_38_1630 ();
 sg13g2_decap_8 FILLER_38_1637 ();
 sg13g2_decap_8 FILLER_38_1644 ();
 sg13g2_decap_8 FILLER_38_1651 ();
 sg13g2_decap_8 FILLER_38_1658 ();
 sg13g2_decap_8 FILLER_38_1665 ();
 sg13g2_decap_8 FILLER_38_1672 ();
 sg13g2_decap_8 FILLER_38_1679 ();
 sg13g2_decap_8 FILLER_38_1686 ();
 sg13g2_decap_8 FILLER_38_1693 ();
 sg13g2_decap_8 FILLER_38_1700 ();
 sg13g2_decap_8 FILLER_38_1707 ();
 sg13g2_decap_8 FILLER_38_1714 ();
 sg13g2_decap_8 FILLER_38_1721 ();
 sg13g2_decap_8 FILLER_38_1728 ();
 sg13g2_decap_8 FILLER_38_1735 ();
 sg13g2_decap_8 FILLER_38_1742 ();
 sg13g2_decap_8 FILLER_38_1749 ();
 sg13g2_decap_8 FILLER_38_1756 ();
 sg13g2_decap_4 FILLER_38_1763 ();
 sg13g2_fill_1 FILLER_38_1767 ();
 sg13g2_fill_2 FILLER_39_26 ();
 sg13g2_fill_1 FILLER_39_28 ();
 sg13g2_fill_2 FILLER_39_43 ();
 sg13g2_fill_2 FILLER_39_54 ();
 sg13g2_fill_1 FILLER_39_56 ();
 sg13g2_fill_1 FILLER_39_92 ();
 sg13g2_fill_2 FILLER_39_110 ();
 sg13g2_fill_2 FILLER_39_175 ();
 sg13g2_fill_1 FILLER_39_186 ();
 sg13g2_fill_2 FILLER_39_208 ();
 sg13g2_fill_1 FILLER_39_210 ();
 sg13g2_fill_1 FILLER_39_224 ();
 sg13g2_fill_2 FILLER_39_261 ();
 sg13g2_fill_1 FILLER_39_263 ();
 sg13g2_fill_2 FILLER_39_304 ();
 sg13g2_fill_2 FILLER_39_325 ();
 sg13g2_fill_1 FILLER_39_327 ();
 sg13g2_decap_4 FILLER_39_410 ();
 sg13g2_fill_1 FILLER_39_422 ();
 sg13g2_fill_2 FILLER_39_449 ();
 sg13g2_fill_1 FILLER_39_451 ();
 sg13g2_fill_2 FILLER_39_475 ();
 sg13g2_fill_1 FILLER_39_477 ();
 sg13g2_fill_2 FILLER_39_487 ();
 sg13g2_fill_1 FILLER_39_489 ();
 sg13g2_fill_1 FILLER_39_509 ();
 sg13g2_fill_2 FILLER_39_534 ();
 sg13g2_fill_2 FILLER_39_545 ();
 sg13g2_fill_1 FILLER_39_547 ();
 sg13g2_fill_2 FILLER_39_603 ();
 sg13g2_fill_2 FILLER_39_639 ();
 sg13g2_fill_2 FILLER_39_671 ();
 sg13g2_fill_2 FILLER_39_703 ();
 sg13g2_fill_1 FILLER_39_705 ();
 sg13g2_decap_4 FILLER_39_737 ();
 sg13g2_fill_1 FILLER_39_741 ();
 sg13g2_decap_4 FILLER_39_750 ();
 sg13g2_fill_1 FILLER_39_754 ();
 sg13g2_fill_2 FILLER_39_788 ();
 sg13g2_fill_1 FILLER_39_790 ();
 sg13g2_fill_2 FILLER_39_827 ();
 sg13g2_fill_1 FILLER_39_859 ();
 sg13g2_fill_2 FILLER_39_901 ();
 sg13g2_fill_2 FILLER_39_950 ();
 sg13g2_fill_2 FILLER_39_988 ();
 sg13g2_fill_1 FILLER_39_990 ();
 sg13g2_fill_2 FILLER_39_1017 ();
 sg13g2_fill_1 FILLER_39_1024 ();
 sg13g2_fill_2 FILLER_39_1077 ();
 sg13g2_fill_2 FILLER_39_1193 ();
 sg13g2_fill_1 FILLER_39_1195 ();
 sg13g2_fill_2 FILLER_39_1208 ();
 sg13g2_fill_2 FILLER_39_1216 ();
 sg13g2_fill_1 FILLER_39_1218 ();
 sg13g2_fill_2 FILLER_39_1223 ();
 sg13g2_fill_2 FILLER_39_1264 ();
 sg13g2_fill_1 FILLER_39_1266 ();
 sg13g2_fill_2 FILLER_39_1280 ();
 sg13g2_fill_1 FILLER_39_1291 ();
 sg13g2_fill_1 FILLER_39_1302 ();
 sg13g2_fill_2 FILLER_39_1338 ();
 sg13g2_fill_1 FILLER_39_1340 ();
 sg13g2_fill_2 FILLER_39_1474 ();
 sg13g2_fill_2 FILLER_39_1503 ();
 sg13g2_decap_8 FILLER_39_1548 ();
 sg13g2_decap_8 FILLER_39_1555 ();
 sg13g2_decap_8 FILLER_39_1562 ();
 sg13g2_decap_8 FILLER_39_1569 ();
 sg13g2_decap_8 FILLER_39_1576 ();
 sg13g2_decap_8 FILLER_39_1583 ();
 sg13g2_decap_8 FILLER_39_1590 ();
 sg13g2_decap_8 FILLER_39_1597 ();
 sg13g2_decap_8 FILLER_39_1604 ();
 sg13g2_decap_8 FILLER_39_1611 ();
 sg13g2_decap_8 FILLER_39_1618 ();
 sg13g2_decap_8 FILLER_39_1625 ();
 sg13g2_decap_8 FILLER_39_1632 ();
 sg13g2_decap_8 FILLER_39_1639 ();
 sg13g2_decap_8 FILLER_39_1646 ();
 sg13g2_decap_8 FILLER_39_1653 ();
 sg13g2_decap_8 FILLER_39_1660 ();
 sg13g2_decap_8 FILLER_39_1667 ();
 sg13g2_decap_8 FILLER_39_1674 ();
 sg13g2_decap_8 FILLER_39_1681 ();
 sg13g2_decap_8 FILLER_39_1688 ();
 sg13g2_decap_8 FILLER_39_1695 ();
 sg13g2_decap_8 FILLER_39_1702 ();
 sg13g2_decap_8 FILLER_39_1709 ();
 sg13g2_decap_8 FILLER_39_1716 ();
 sg13g2_decap_8 FILLER_39_1723 ();
 sg13g2_decap_8 FILLER_39_1730 ();
 sg13g2_decap_8 FILLER_39_1737 ();
 sg13g2_decap_8 FILLER_39_1744 ();
 sg13g2_decap_8 FILLER_39_1751 ();
 sg13g2_decap_8 FILLER_39_1758 ();
 sg13g2_fill_2 FILLER_39_1765 ();
 sg13g2_fill_1 FILLER_39_1767 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_19 ();
 sg13g2_decap_4 FILLER_40_82 ();
 sg13g2_fill_2 FILLER_40_86 ();
 sg13g2_fill_1 FILLER_40_107 ();
 sg13g2_fill_2 FILLER_40_123 ();
 sg13g2_fill_2 FILLER_40_135 ();
 sg13g2_fill_1 FILLER_40_141 ();
 sg13g2_fill_2 FILLER_40_177 ();
 sg13g2_fill_2 FILLER_40_201 ();
 sg13g2_fill_1 FILLER_40_203 ();
 sg13g2_fill_2 FILLER_40_277 ();
 sg13g2_fill_1 FILLER_40_279 ();
 sg13g2_fill_1 FILLER_40_299 ();
 sg13g2_fill_1 FILLER_40_330 ();
 sg13g2_fill_2 FILLER_40_342 ();
 sg13g2_fill_2 FILLER_40_393 ();
 sg13g2_fill_2 FILLER_40_415 ();
 sg13g2_fill_2 FILLER_40_431 ();
 sg13g2_fill_1 FILLER_40_441 ();
 sg13g2_fill_2 FILLER_40_550 ();
 sg13g2_fill_1 FILLER_40_552 ();
 sg13g2_fill_1 FILLER_40_572 ();
 sg13g2_fill_1 FILLER_40_696 ();
 sg13g2_fill_2 FILLER_40_710 ();
 sg13g2_fill_1 FILLER_40_712 ();
 sg13g2_decap_4 FILLER_40_735 ();
 sg13g2_fill_1 FILLER_40_739 ();
 sg13g2_fill_2 FILLER_40_925 ();
 sg13g2_fill_1 FILLER_40_987 ();
 sg13g2_fill_2 FILLER_40_1035 ();
 sg13g2_fill_1 FILLER_40_1037 ();
 sg13g2_fill_2 FILLER_40_1066 ();
 sg13g2_fill_1 FILLER_40_1068 ();
 sg13g2_fill_2 FILLER_40_1094 ();
 sg13g2_fill_2 FILLER_40_1120 ();
 sg13g2_fill_1 FILLER_40_1122 ();
 sg13g2_fill_2 FILLER_40_1137 ();
 sg13g2_fill_2 FILLER_40_1144 ();
 sg13g2_fill_1 FILLER_40_1146 ();
 sg13g2_fill_2 FILLER_40_1317 ();
 sg13g2_fill_1 FILLER_40_1319 ();
 sg13g2_fill_1 FILLER_40_1366 ();
 sg13g2_decap_4 FILLER_40_1409 ();
 sg13g2_fill_1 FILLER_40_1426 ();
 sg13g2_fill_2 FILLER_40_1433 ();
 sg13g2_decap_4 FILLER_40_1449 ();
 sg13g2_fill_1 FILLER_40_1453 ();
 sg13g2_fill_1 FILLER_40_1463 ();
 sg13g2_fill_2 FILLER_40_1494 ();
 sg13g2_decap_8 FILLER_40_1536 ();
 sg13g2_decap_8 FILLER_40_1543 ();
 sg13g2_decap_8 FILLER_40_1550 ();
 sg13g2_decap_8 FILLER_40_1557 ();
 sg13g2_decap_8 FILLER_40_1564 ();
 sg13g2_decap_8 FILLER_40_1571 ();
 sg13g2_decap_8 FILLER_40_1578 ();
 sg13g2_decap_8 FILLER_40_1585 ();
 sg13g2_decap_8 FILLER_40_1592 ();
 sg13g2_decap_8 FILLER_40_1599 ();
 sg13g2_decap_8 FILLER_40_1606 ();
 sg13g2_decap_8 FILLER_40_1613 ();
 sg13g2_decap_8 FILLER_40_1620 ();
 sg13g2_decap_8 FILLER_40_1627 ();
 sg13g2_decap_8 FILLER_40_1634 ();
 sg13g2_decap_8 FILLER_40_1641 ();
 sg13g2_decap_8 FILLER_40_1648 ();
 sg13g2_decap_8 FILLER_40_1655 ();
 sg13g2_decap_8 FILLER_40_1662 ();
 sg13g2_decap_8 FILLER_40_1669 ();
 sg13g2_decap_8 FILLER_40_1676 ();
 sg13g2_decap_8 FILLER_40_1683 ();
 sg13g2_decap_8 FILLER_40_1690 ();
 sg13g2_decap_8 FILLER_40_1697 ();
 sg13g2_decap_8 FILLER_40_1704 ();
 sg13g2_decap_8 FILLER_40_1711 ();
 sg13g2_decap_8 FILLER_40_1718 ();
 sg13g2_decap_8 FILLER_40_1725 ();
 sg13g2_decap_8 FILLER_40_1732 ();
 sg13g2_decap_8 FILLER_40_1739 ();
 sg13g2_decap_8 FILLER_40_1746 ();
 sg13g2_decap_8 FILLER_40_1753 ();
 sg13g2_decap_8 FILLER_40_1760 ();
 sg13g2_fill_1 FILLER_40_1767 ();
 sg13g2_fill_2 FILLER_41_31 ();
 sg13g2_fill_1 FILLER_41_33 ();
 sg13g2_fill_2 FILLER_41_56 ();
 sg13g2_fill_2 FILLER_41_114 ();
 sg13g2_fill_1 FILLER_41_116 ();
 sg13g2_fill_2 FILLER_41_157 ();
 sg13g2_fill_1 FILLER_41_159 ();
 sg13g2_fill_2 FILLER_41_212 ();
 sg13g2_fill_1 FILLER_41_214 ();
 sg13g2_fill_1 FILLER_41_277 ();
 sg13g2_fill_2 FILLER_41_334 ();
 sg13g2_fill_1 FILLER_41_336 ();
 sg13g2_fill_2 FILLER_41_368 ();
 sg13g2_fill_2 FILLER_41_378 ();
 sg13g2_fill_1 FILLER_41_380 ();
 sg13g2_fill_1 FILLER_41_390 ();
 sg13g2_fill_2 FILLER_41_452 ();
 sg13g2_fill_1 FILLER_41_454 ();
 sg13g2_fill_1 FILLER_41_464 ();
 sg13g2_fill_1 FILLER_41_490 ();
 sg13g2_fill_2 FILLER_41_496 ();
 sg13g2_fill_1 FILLER_41_498 ();
 sg13g2_fill_2 FILLER_41_503 ();
 sg13g2_fill_1 FILLER_41_505 ();
 sg13g2_decap_4 FILLER_41_514 ();
 sg13g2_fill_1 FILLER_41_518 ();
 sg13g2_fill_1 FILLER_41_528 ();
 sg13g2_fill_2 FILLER_41_559 ();
 sg13g2_fill_1 FILLER_41_561 ();
 sg13g2_fill_1 FILLER_41_570 ();
 sg13g2_fill_2 FILLER_41_584 ();
 sg13g2_fill_1 FILLER_41_586 ();
 sg13g2_fill_1 FILLER_41_602 ();
 sg13g2_fill_2 FILLER_41_616 ();
 sg13g2_fill_2 FILLER_41_631 ();
 sg13g2_fill_1 FILLER_41_633 ();
 sg13g2_fill_2 FILLER_41_652 ();
 sg13g2_fill_2 FILLER_41_659 ();
 sg13g2_fill_1 FILLER_41_661 ();
 sg13g2_fill_2 FILLER_41_680 ();
 sg13g2_fill_1 FILLER_41_682 ();
 sg13g2_fill_1 FILLER_41_709 ();
 sg13g2_decap_8 FILLER_41_740 ();
 sg13g2_fill_2 FILLER_41_747 ();
 sg13g2_fill_1 FILLER_41_778 ();
 sg13g2_fill_2 FILLER_41_788 ();
 sg13g2_fill_2 FILLER_41_809 ();
 sg13g2_fill_2 FILLER_41_837 ();
 sg13g2_fill_1 FILLER_41_871 ();
 sg13g2_decap_8 FILLER_41_895 ();
 sg13g2_fill_2 FILLER_41_907 ();
 sg13g2_fill_1 FILLER_41_909 ();
 sg13g2_fill_2 FILLER_41_914 ();
 sg13g2_fill_1 FILLER_41_916 ();
 sg13g2_fill_2 FILLER_41_941 ();
 sg13g2_fill_1 FILLER_41_949 ();
 sg13g2_fill_1 FILLER_41_1076 ();
 sg13g2_fill_2 FILLER_41_1103 ();
 sg13g2_fill_1 FILLER_41_1105 ();
 sg13g2_fill_2 FILLER_41_1138 ();
 sg13g2_fill_1 FILLER_41_1140 ();
 sg13g2_fill_2 FILLER_41_1177 ();
 sg13g2_fill_2 FILLER_41_1204 ();
 sg13g2_fill_2 FILLER_41_1226 ();
 sg13g2_fill_1 FILLER_41_1228 ();
 sg13g2_fill_1 FILLER_41_1246 ();
 sg13g2_fill_2 FILLER_41_1256 ();
 sg13g2_fill_1 FILLER_41_1258 ();
 sg13g2_fill_1 FILLER_41_1274 ();
 sg13g2_fill_2 FILLER_41_1307 ();
 sg13g2_fill_1 FILLER_41_1331 ();
 sg13g2_fill_2 FILLER_41_1370 ();
 sg13g2_fill_1 FILLER_41_1372 ();
 sg13g2_fill_1 FILLER_41_1387 ();
 sg13g2_fill_2 FILLER_41_1419 ();
 sg13g2_fill_1 FILLER_41_1421 ();
 sg13g2_fill_2 FILLER_41_1454 ();
 sg13g2_fill_1 FILLER_41_1469 ();
 sg13g2_decap_8 FILLER_41_1537 ();
 sg13g2_decap_8 FILLER_41_1544 ();
 sg13g2_decap_8 FILLER_41_1551 ();
 sg13g2_decap_8 FILLER_41_1558 ();
 sg13g2_decap_8 FILLER_41_1565 ();
 sg13g2_decap_8 FILLER_41_1572 ();
 sg13g2_decap_8 FILLER_41_1579 ();
 sg13g2_decap_8 FILLER_41_1586 ();
 sg13g2_decap_8 FILLER_41_1593 ();
 sg13g2_decap_8 FILLER_41_1600 ();
 sg13g2_decap_8 FILLER_41_1607 ();
 sg13g2_decap_8 FILLER_41_1614 ();
 sg13g2_decap_8 FILLER_41_1621 ();
 sg13g2_decap_8 FILLER_41_1628 ();
 sg13g2_decap_8 FILLER_41_1635 ();
 sg13g2_decap_8 FILLER_41_1642 ();
 sg13g2_decap_8 FILLER_41_1649 ();
 sg13g2_decap_8 FILLER_41_1656 ();
 sg13g2_decap_8 FILLER_41_1663 ();
 sg13g2_decap_8 FILLER_41_1670 ();
 sg13g2_decap_8 FILLER_41_1677 ();
 sg13g2_decap_8 FILLER_41_1684 ();
 sg13g2_decap_8 FILLER_41_1691 ();
 sg13g2_decap_8 FILLER_41_1698 ();
 sg13g2_decap_8 FILLER_41_1705 ();
 sg13g2_decap_8 FILLER_41_1712 ();
 sg13g2_decap_8 FILLER_41_1719 ();
 sg13g2_decap_8 FILLER_41_1726 ();
 sg13g2_decap_8 FILLER_41_1733 ();
 sg13g2_decap_8 FILLER_41_1740 ();
 sg13g2_decap_8 FILLER_41_1747 ();
 sg13g2_decap_8 FILLER_41_1754 ();
 sg13g2_decap_8 FILLER_41_1761 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_9 ();
 sg13g2_fill_2 FILLER_42_31 ();
 sg13g2_fill_1 FILLER_42_33 ();
 sg13g2_fill_1 FILLER_42_68 ();
 sg13g2_fill_2 FILLER_42_85 ();
 sg13g2_fill_1 FILLER_42_87 ();
 sg13g2_fill_2 FILLER_42_126 ();
 sg13g2_fill_2 FILLER_42_136 ();
 sg13g2_fill_1 FILLER_42_138 ();
 sg13g2_fill_1 FILLER_42_144 ();
 sg13g2_fill_2 FILLER_42_150 ();
 sg13g2_fill_1 FILLER_42_152 ();
 sg13g2_fill_2 FILLER_42_157 ();
 sg13g2_fill_1 FILLER_42_159 ();
 sg13g2_fill_1 FILLER_42_164 ();
 sg13g2_fill_1 FILLER_42_177 ();
 sg13g2_fill_1 FILLER_42_192 ();
 sg13g2_fill_1 FILLER_42_205 ();
 sg13g2_fill_1 FILLER_42_237 ();
 sg13g2_fill_2 FILLER_42_247 ();
 sg13g2_decap_4 FILLER_42_282 ();
 sg13g2_fill_1 FILLER_42_286 ();
 sg13g2_fill_2 FILLER_42_352 ();
 sg13g2_fill_1 FILLER_42_354 ();
 sg13g2_fill_2 FILLER_42_427 ();
 sg13g2_fill_1 FILLER_42_469 ();
 sg13g2_fill_1 FILLER_42_496 ();
 sg13g2_fill_2 FILLER_42_523 ();
 sg13g2_fill_1 FILLER_42_539 ();
 sg13g2_fill_1 FILLER_42_563 ();
 sg13g2_fill_1 FILLER_42_604 ();
 sg13g2_fill_2 FILLER_42_687 ();
 sg13g2_fill_1 FILLER_42_689 ();
 sg13g2_fill_2 FILLER_42_720 ();
 sg13g2_fill_2 FILLER_42_730 ();
 sg13g2_decap_4 FILLER_42_745 ();
 sg13g2_fill_1 FILLER_42_749 ();
 sg13g2_fill_2 FILLER_42_806 ();
 sg13g2_fill_1 FILLER_42_847 ();
 sg13g2_fill_2 FILLER_42_968 ();
 sg13g2_fill_2 FILLER_42_984 ();
 sg13g2_fill_2 FILLER_42_1029 ();
 sg13g2_fill_2 FILLER_42_1044 ();
 sg13g2_decap_8 FILLER_42_1079 ();
 sg13g2_fill_2 FILLER_42_1086 ();
 sg13g2_fill_2 FILLER_42_1108 ();
 sg13g2_fill_1 FILLER_42_1110 ();
 sg13g2_fill_2 FILLER_42_1124 ();
 sg13g2_fill_1 FILLER_42_1126 ();
 sg13g2_fill_1 FILLER_42_1185 ();
 sg13g2_fill_2 FILLER_42_1238 ();
 sg13g2_fill_2 FILLER_42_1266 ();
 sg13g2_fill_1 FILLER_42_1268 ();
 sg13g2_fill_2 FILLER_42_1295 ();
 sg13g2_fill_1 FILLER_42_1495 ();
 sg13g2_decap_8 FILLER_42_1526 ();
 sg13g2_decap_8 FILLER_42_1533 ();
 sg13g2_decap_8 FILLER_42_1540 ();
 sg13g2_decap_8 FILLER_42_1547 ();
 sg13g2_decap_8 FILLER_42_1554 ();
 sg13g2_decap_8 FILLER_42_1561 ();
 sg13g2_decap_8 FILLER_42_1568 ();
 sg13g2_decap_8 FILLER_42_1575 ();
 sg13g2_decap_8 FILLER_42_1582 ();
 sg13g2_decap_8 FILLER_42_1589 ();
 sg13g2_decap_8 FILLER_42_1596 ();
 sg13g2_decap_8 FILLER_42_1603 ();
 sg13g2_decap_8 FILLER_42_1610 ();
 sg13g2_decap_8 FILLER_42_1617 ();
 sg13g2_decap_8 FILLER_42_1624 ();
 sg13g2_decap_8 FILLER_42_1631 ();
 sg13g2_decap_8 FILLER_42_1638 ();
 sg13g2_decap_8 FILLER_42_1645 ();
 sg13g2_decap_8 FILLER_42_1652 ();
 sg13g2_decap_8 FILLER_42_1659 ();
 sg13g2_decap_8 FILLER_42_1666 ();
 sg13g2_decap_8 FILLER_42_1673 ();
 sg13g2_decap_8 FILLER_42_1680 ();
 sg13g2_decap_8 FILLER_42_1687 ();
 sg13g2_decap_8 FILLER_42_1694 ();
 sg13g2_decap_8 FILLER_42_1701 ();
 sg13g2_decap_8 FILLER_42_1708 ();
 sg13g2_decap_8 FILLER_42_1715 ();
 sg13g2_decap_8 FILLER_42_1722 ();
 sg13g2_decap_8 FILLER_42_1729 ();
 sg13g2_decap_8 FILLER_42_1736 ();
 sg13g2_decap_8 FILLER_42_1743 ();
 sg13g2_decap_8 FILLER_42_1750 ();
 sg13g2_decap_8 FILLER_42_1757 ();
 sg13g2_decap_4 FILLER_42_1764 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_48 ();
 sg13g2_fill_2 FILLER_43_105 ();
 sg13g2_fill_1 FILLER_43_107 ();
 sg13g2_fill_2 FILLER_43_234 ();
 sg13g2_fill_1 FILLER_43_236 ();
 sg13g2_fill_2 FILLER_43_263 ();
 sg13g2_decap_4 FILLER_43_274 ();
 sg13g2_fill_1 FILLER_43_308 ();
 sg13g2_fill_2 FILLER_43_339 ();
 sg13g2_fill_1 FILLER_43_341 ();
 sg13g2_fill_1 FILLER_43_368 ();
 sg13g2_fill_2 FILLER_43_388 ();
 sg13g2_fill_1 FILLER_43_390 ();
 sg13g2_fill_2 FILLER_43_417 ();
 sg13g2_fill_2 FILLER_43_477 ();
 sg13g2_fill_1 FILLER_43_479 ();
 sg13g2_decap_8 FILLER_43_499 ();
 sg13g2_fill_2 FILLER_43_506 ();
 sg13g2_decap_8 FILLER_43_512 ();
 sg13g2_fill_2 FILLER_43_519 ();
 sg13g2_fill_1 FILLER_43_521 ();
 sg13g2_decap_4 FILLER_43_537 ();
 sg13g2_fill_2 FILLER_43_541 ();
 sg13g2_decap_4 FILLER_43_547 ();
 sg13g2_fill_2 FILLER_43_561 ();
 sg13g2_fill_1 FILLER_43_572 ();
 sg13g2_decap_8 FILLER_43_588 ();
 sg13g2_fill_2 FILLER_43_595 ();
 sg13g2_fill_1 FILLER_43_597 ();
 sg13g2_fill_2 FILLER_43_624 ();
 sg13g2_fill_1 FILLER_43_626 ();
 sg13g2_fill_2 FILLER_43_653 ();
 sg13g2_fill_2 FILLER_43_673 ();
 sg13g2_fill_2 FILLER_43_783 ();
 sg13g2_fill_1 FILLER_43_785 ();
 sg13g2_fill_2 FILLER_43_824 ();
 sg13g2_fill_1 FILLER_43_834 ();
 sg13g2_fill_1 FILLER_43_844 ();
 sg13g2_fill_2 FILLER_43_876 ();
 sg13g2_fill_2 FILLER_43_896 ();
 sg13g2_decap_8 FILLER_43_916 ();
 sg13g2_fill_2 FILLER_43_923 ();
 sg13g2_fill_1 FILLER_43_925 ();
 sg13g2_fill_2 FILLER_43_931 ();
 sg13g2_decap_4 FILLER_43_941 ();
 sg13g2_fill_1 FILLER_43_945 ();
 sg13g2_fill_2 FILLER_43_1006 ();
 sg13g2_fill_2 FILLER_43_1051 ();
 sg13g2_fill_2 FILLER_43_1074 ();
 sg13g2_fill_1 FILLER_43_1116 ();
 sg13g2_fill_1 FILLER_43_1131 ();
 sg13g2_fill_2 FILLER_43_1171 ();
 sg13g2_fill_2 FILLER_43_1187 ();
 sg13g2_fill_2 FILLER_43_1203 ();
 sg13g2_fill_1 FILLER_43_1226 ();
 sg13g2_fill_2 FILLER_43_1254 ();
 sg13g2_fill_1 FILLER_43_1256 ();
 sg13g2_fill_2 FILLER_43_1262 ();
 sg13g2_fill_2 FILLER_43_1292 ();
 sg13g2_fill_1 FILLER_43_1325 ();
 sg13g2_fill_1 FILLER_43_1387 ();
 sg13g2_decap_8 FILLER_43_1529 ();
 sg13g2_decap_8 FILLER_43_1536 ();
 sg13g2_decap_8 FILLER_43_1543 ();
 sg13g2_decap_8 FILLER_43_1550 ();
 sg13g2_decap_8 FILLER_43_1557 ();
 sg13g2_decap_8 FILLER_43_1564 ();
 sg13g2_decap_8 FILLER_43_1571 ();
 sg13g2_decap_8 FILLER_43_1578 ();
 sg13g2_decap_8 FILLER_43_1585 ();
 sg13g2_decap_8 FILLER_43_1592 ();
 sg13g2_decap_8 FILLER_43_1599 ();
 sg13g2_decap_8 FILLER_43_1606 ();
 sg13g2_decap_8 FILLER_43_1613 ();
 sg13g2_decap_8 FILLER_43_1620 ();
 sg13g2_decap_8 FILLER_43_1627 ();
 sg13g2_decap_8 FILLER_43_1634 ();
 sg13g2_decap_8 FILLER_43_1641 ();
 sg13g2_decap_8 FILLER_43_1648 ();
 sg13g2_decap_8 FILLER_43_1655 ();
 sg13g2_decap_8 FILLER_43_1662 ();
 sg13g2_decap_8 FILLER_43_1669 ();
 sg13g2_decap_8 FILLER_43_1676 ();
 sg13g2_decap_8 FILLER_43_1683 ();
 sg13g2_decap_8 FILLER_43_1690 ();
 sg13g2_decap_8 FILLER_43_1697 ();
 sg13g2_decap_8 FILLER_43_1704 ();
 sg13g2_decap_8 FILLER_43_1711 ();
 sg13g2_decap_8 FILLER_43_1718 ();
 sg13g2_decap_8 FILLER_43_1725 ();
 sg13g2_decap_8 FILLER_43_1732 ();
 sg13g2_decap_8 FILLER_43_1739 ();
 sg13g2_decap_8 FILLER_43_1746 ();
 sg13g2_decap_8 FILLER_43_1753 ();
 sg13g2_decap_8 FILLER_43_1760 ();
 sg13g2_fill_1 FILLER_43_1767 ();
 sg13g2_fill_2 FILLER_44_66 ();
 sg13g2_fill_2 FILLER_44_82 ();
 sg13g2_fill_1 FILLER_44_84 ();
 sg13g2_fill_2 FILLER_44_94 ();
 sg13g2_fill_1 FILLER_44_127 ();
 sg13g2_fill_2 FILLER_44_236 ();
 sg13g2_fill_1 FILLER_44_248 ();
 sg13g2_fill_2 FILLER_44_306 ();
 sg13g2_fill_1 FILLER_44_348 ();
 sg13g2_decap_4 FILLER_44_358 ();
 sg13g2_fill_2 FILLER_44_362 ();
 sg13g2_fill_1 FILLER_44_452 ();
 sg13g2_fill_2 FILLER_44_463 ();
 sg13g2_fill_2 FILLER_44_470 ();
 sg13g2_fill_2 FILLER_44_477 ();
 sg13g2_fill_1 FILLER_44_479 ();
 sg13g2_decap_4 FILLER_44_484 ();
 sg13g2_fill_1 FILLER_44_488 ();
 sg13g2_fill_2 FILLER_44_494 ();
 sg13g2_decap_8 FILLER_44_501 ();
 sg13g2_fill_2 FILLER_44_508 ();
 sg13g2_fill_1 FILLER_44_567 ();
 sg13g2_fill_2 FILLER_44_572 ();
 sg13g2_fill_1 FILLER_44_574 ();
 sg13g2_fill_1 FILLER_44_600 ();
 sg13g2_fill_1 FILLER_44_640 ();
 sg13g2_fill_1 FILLER_44_655 ();
 sg13g2_fill_1 FILLER_44_691 ();
 sg13g2_decap_8 FILLER_44_696 ();
 sg13g2_decap_4 FILLER_44_703 ();
 sg13g2_fill_2 FILLER_44_707 ();
 sg13g2_fill_2 FILLER_44_713 ();
 sg13g2_decap_4 FILLER_44_750 ();
 sg13g2_fill_1 FILLER_44_784 ();
 sg13g2_fill_1 FILLER_44_810 ();
 sg13g2_fill_2 FILLER_44_849 ();
 sg13g2_fill_1 FILLER_44_881 ();
 sg13g2_fill_1 FILLER_44_1016 ();
 sg13g2_decap_8 FILLER_44_1033 ();
 sg13g2_fill_1 FILLER_44_1040 ();
 sg13g2_fill_1 FILLER_44_1158 ();
 sg13g2_fill_1 FILLER_44_1302 ();
 sg13g2_fill_2 FILLER_44_1308 ();
 sg13g2_decap_4 FILLER_44_1369 ();
 sg13g2_fill_2 FILLER_44_1373 ();
 sg13g2_fill_1 FILLER_44_1445 ();
 sg13g2_fill_1 FILLER_44_1485 ();
 sg13g2_fill_1 FILLER_44_1494 ();
 sg13g2_decap_8 FILLER_44_1517 ();
 sg13g2_decap_8 FILLER_44_1524 ();
 sg13g2_decap_4 FILLER_44_1531 ();
 sg13g2_fill_1 FILLER_44_1535 ();
 sg13g2_decap_8 FILLER_44_1540 ();
 sg13g2_decap_8 FILLER_44_1547 ();
 sg13g2_decap_8 FILLER_44_1554 ();
 sg13g2_decap_8 FILLER_44_1561 ();
 sg13g2_decap_8 FILLER_44_1568 ();
 sg13g2_decap_8 FILLER_44_1575 ();
 sg13g2_decap_8 FILLER_44_1582 ();
 sg13g2_decap_8 FILLER_44_1589 ();
 sg13g2_decap_8 FILLER_44_1596 ();
 sg13g2_decap_8 FILLER_44_1603 ();
 sg13g2_decap_8 FILLER_44_1610 ();
 sg13g2_decap_8 FILLER_44_1617 ();
 sg13g2_decap_8 FILLER_44_1624 ();
 sg13g2_decap_8 FILLER_44_1631 ();
 sg13g2_decap_8 FILLER_44_1638 ();
 sg13g2_decap_8 FILLER_44_1645 ();
 sg13g2_decap_8 FILLER_44_1652 ();
 sg13g2_decap_8 FILLER_44_1659 ();
 sg13g2_decap_8 FILLER_44_1666 ();
 sg13g2_decap_8 FILLER_44_1673 ();
 sg13g2_decap_8 FILLER_44_1680 ();
 sg13g2_decap_8 FILLER_44_1687 ();
 sg13g2_decap_8 FILLER_44_1694 ();
 sg13g2_decap_8 FILLER_44_1701 ();
 sg13g2_decap_8 FILLER_44_1708 ();
 sg13g2_decap_8 FILLER_44_1715 ();
 sg13g2_decap_8 FILLER_44_1722 ();
 sg13g2_decap_8 FILLER_44_1729 ();
 sg13g2_decap_8 FILLER_44_1736 ();
 sg13g2_decap_8 FILLER_44_1743 ();
 sg13g2_decap_8 FILLER_44_1750 ();
 sg13g2_decap_8 FILLER_44_1757 ();
 sg13g2_decap_4 FILLER_44_1764 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_fill_2 FILLER_45_33 ();
 sg13g2_fill_2 FILLER_45_61 ();
 sg13g2_fill_2 FILLER_45_81 ();
 sg13g2_fill_1 FILLER_45_83 ();
 sg13g2_fill_2 FILLER_45_117 ();
 sg13g2_fill_2 FILLER_45_127 ();
 sg13g2_fill_1 FILLER_45_249 ();
 sg13g2_fill_1 FILLER_45_254 ();
 sg13g2_fill_1 FILLER_45_269 ();
 sg13g2_fill_1 FILLER_45_288 ();
 sg13g2_fill_1 FILLER_45_302 ();
 sg13g2_fill_2 FILLER_45_312 ();
 sg13g2_fill_1 FILLER_45_314 ();
 sg13g2_fill_1 FILLER_45_332 ();
 sg13g2_decap_8 FILLER_45_359 ();
 sg13g2_fill_2 FILLER_45_378 ();
 sg13g2_fill_1 FILLER_45_380 ();
 sg13g2_fill_2 FILLER_45_389 ();
 sg13g2_fill_2 FILLER_45_425 ();
 sg13g2_fill_2 FILLER_45_475 ();
 sg13g2_fill_1 FILLER_45_477 ();
 sg13g2_fill_1 FILLER_45_528 ();
 sg13g2_fill_2 FILLER_45_569 ();
 sg13g2_fill_1 FILLER_45_571 ();
 sg13g2_fill_1 FILLER_45_588 ();
 sg13g2_decap_8 FILLER_45_600 ();
 sg13g2_decap_4 FILLER_45_607 ();
 sg13g2_fill_2 FILLER_45_611 ();
 sg13g2_fill_2 FILLER_45_635 ();
 sg13g2_fill_1 FILLER_45_637 ();
 sg13g2_fill_2 FILLER_45_672 ();
 sg13g2_decap_4 FILLER_45_678 ();
 sg13g2_fill_1 FILLER_45_682 ();
 sg13g2_fill_1 FILLER_45_725 ();
 sg13g2_decap_4 FILLER_45_732 ();
 sg13g2_fill_1 FILLER_45_758 ();
 sg13g2_fill_2 FILLER_45_777 ();
 sg13g2_fill_1 FILLER_45_805 ();
 sg13g2_fill_2 FILLER_45_837 ();
 sg13g2_fill_1 FILLER_45_870 ();
 sg13g2_decap_8 FILLER_45_906 ();
 sg13g2_fill_2 FILLER_45_913 ();
 sg13g2_fill_2 FILLER_45_923 ();
 sg13g2_decap_4 FILLER_45_955 ();
 sg13g2_fill_2 FILLER_45_994 ();
 sg13g2_fill_1 FILLER_45_996 ();
 sg13g2_decap_8 FILLER_45_1019 ();
 sg13g2_decap_8 FILLER_45_1026 ();
 sg13g2_decap_4 FILLER_45_1033 ();
 sg13g2_decap_8 FILLER_45_1045 ();
 sg13g2_fill_1 FILLER_45_1056 ();
 sg13g2_fill_2 FILLER_45_1065 ();
 sg13g2_fill_1 FILLER_45_1077 ();
 sg13g2_decap_4 FILLER_45_1096 ();
 sg13g2_fill_1 FILLER_45_1100 ();
 sg13g2_fill_2 FILLER_45_1106 ();
 sg13g2_fill_2 FILLER_45_1116 ();
 sg13g2_fill_1 FILLER_45_1118 ();
 sg13g2_fill_2 FILLER_45_1127 ();
 sg13g2_fill_1 FILLER_45_1129 ();
 sg13g2_fill_2 FILLER_45_1135 ();
 sg13g2_fill_2 FILLER_45_1172 ();
 sg13g2_fill_1 FILLER_45_1174 ();
 sg13g2_fill_1 FILLER_45_1189 ();
 sg13g2_fill_2 FILLER_45_1230 ();
 sg13g2_fill_1 FILLER_45_1232 ();
 sg13g2_fill_2 FILLER_45_1270 ();
 sg13g2_decap_8 FILLER_45_1376 ();
 sg13g2_fill_1 FILLER_45_1383 ();
 sg13g2_fill_2 FILLER_45_1443 ();
 sg13g2_fill_2 FILLER_45_1462 ();
 sg13g2_fill_1 FILLER_45_1464 ();
 sg13g2_fill_2 FILLER_45_1491 ();
 sg13g2_fill_2 FILLER_45_1497 ();
 sg13g2_decap_8 FILLER_45_1551 ();
 sg13g2_fill_1 FILLER_45_1558 ();
 sg13g2_fill_2 FILLER_45_1563 ();
 sg13g2_decap_8 FILLER_45_1570 ();
 sg13g2_decap_4 FILLER_45_1577 ();
 sg13g2_fill_2 FILLER_45_1585 ();
 sg13g2_fill_1 FILLER_45_1587 ();
 sg13g2_decap_8 FILLER_45_1597 ();
 sg13g2_decap_8 FILLER_45_1604 ();
 sg13g2_decap_8 FILLER_45_1611 ();
 sg13g2_decap_8 FILLER_45_1618 ();
 sg13g2_decap_8 FILLER_45_1625 ();
 sg13g2_decap_8 FILLER_45_1632 ();
 sg13g2_decap_8 FILLER_45_1639 ();
 sg13g2_decap_8 FILLER_45_1646 ();
 sg13g2_decap_8 FILLER_45_1653 ();
 sg13g2_decap_8 FILLER_45_1660 ();
 sg13g2_decap_8 FILLER_45_1667 ();
 sg13g2_decap_8 FILLER_45_1674 ();
 sg13g2_decap_8 FILLER_45_1681 ();
 sg13g2_decap_8 FILLER_45_1688 ();
 sg13g2_decap_8 FILLER_45_1695 ();
 sg13g2_decap_8 FILLER_45_1702 ();
 sg13g2_decap_8 FILLER_45_1709 ();
 sg13g2_decap_8 FILLER_45_1716 ();
 sg13g2_decap_8 FILLER_45_1723 ();
 sg13g2_decap_8 FILLER_45_1730 ();
 sg13g2_decap_8 FILLER_45_1737 ();
 sg13g2_decap_8 FILLER_45_1744 ();
 sg13g2_decap_8 FILLER_45_1751 ();
 sg13g2_decap_8 FILLER_45_1758 ();
 sg13g2_fill_2 FILLER_45_1765 ();
 sg13g2_fill_1 FILLER_45_1767 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_27 ();
 sg13g2_fill_1 FILLER_46_29 ();
 sg13g2_fill_1 FILLER_46_135 ();
 sg13g2_fill_1 FILLER_46_155 ();
 sg13g2_fill_2 FILLER_46_185 ();
 sg13g2_fill_2 FILLER_46_203 ();
 sg13g2_fill_2 FILLER_46_214 ();
 sg13g2_fill_2 FILLER_46_306 ();
 sg13g2_fill_2 FILLER_46_343 ();
 sg13g2_fill_1 FILLER_46_371 ();
 sg13g2_fill_2 FILLER_46_404 ();
 sg13g2_fill_2 FILLER_46_432 ();
 sg13g2_fill_1 FILLER_46_434 ();
 sg13g2_fill_1 FILLER_46_445 ();
 sg13g2_fill_1 FILLER_46_474 ();
 sg13g2_decap_4 FILLER_46_499 ();
 sg13g2_decap_4 FILLER_46_507 ();
 sg13g2_fill_1 FILLER_46_522 ();
 sg13g2_fill_2 FILLER_46_529 ();
 sg13g2_decap_4 FILLER_46_543 ();
 sg13g2_fill_2 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_fill_2 FILLER_46_567 ();
 sg13g2_fill_1 FILLER_46_569 ();
 sg13g2_fill_1 FILLER_46_606 ();
 sg13g2_decap_8 FILLER_46_637 ();
 sg13g2_fill_1 FILLER_46_644 ();
 sg13g2_fill_2 FILLER_46_660 ();
 sg13g2_fill_1 FILLER_46_662 ();
 sg13g2_fill_1 FILLER_46_689 ();
 sg13g2_fill_1 FILLER_46_711 ();
 sg13g2_decap_8 FILLER_46_762 ();
 sg13g2_fill_2 FILLER_46_769 ();
 sg13g2_fill_1 FILLER_46_771 ();
 sg13g2_fill_2 FILLER_46_797 ();
 sg13g2_fill_1 FILLER_46_799 ();
 sg13g2_fill_1 FILLER_46_848 ();
 sg13g2_fill_2 FILLER_46_857 ();
 sg13g2_fill_1 FILLER_46_894 ();
 sg13g2_fill_2 FILLER_46_978 ();
 sg13g2_fill_1 FILLER_46_984 ();
 sg13g2_fill_2 FILLER_46_1089 ();
 sg13g2_fill_1 FILLER_46_1091 ();
 sg13g2_fill_2 FILLER_46_1148 ();
 sg13g2_fill_2 FILLER_46_1180 ();
 sg13g2_fill_2 FILLER_46_1217 ();
 sg13g2_fill_2 FILLER_46_1276 ();
 sg13g2_fill_2 FILLER_46_1296 ();
 sg13g2_fill_1 FILLER_46_1298 ();
 sg13g2_fill_2 FILLER_46_1341 ();
 sg13g2_fill_2 FILLER_46_1361 ();
 sg13g2_fill_1 FILLER_46_1363 ();
 sg13g2_fill_2 FILLER_46_1416 ();
 sg13g2_fill_2 FILLER_46_1432 ();
 sg13g2_fill_1 FILLER_46_1434 ();
 sg13g2_fill_1 FILLER_46_1502 ();
 sg13g2_fill_1 FILLER_46_1521 ();
 sg13g2_fill_1 FILLER_46_1562 ();
 sg13g2_fill_2 FILLER_46_1589 ();
 sg13g2_decap_8 FILLER_46_1617 ();
 sg13g2_decap_8 FILLER_46_1624 ();
 sg13g2_decap_8 FILLER_46_1631 ();
 sg13g2_decap_8 FILLER_46_1638 ();
 sg13g2_decap_8 FILLER_46_1645 ();
 sg13g2_decap_8 FILLER_46_1652 ();
 sg13g2_decap_8 FILLER_46_1659 ();
 sg13g2_decap_8 FILLER_46_1666 ();
 sg13g2_decap_8 FILLER_46_1673 ();
 sg13g2_decap_8 FILLER_46_1680 ();
 sg13g2_decap_8 FILLER_46_1687 ();
 sg13g2_decap_8 FILLER_46_1694 ();
 sg13g2_decap_8 FILLER_46_1701 ();
 sg13g2_decap_8 FILLER_46_1708 ();
 sg13g2_decap_8 FILLER_46_1715 ();
 sg13g2_decap_8 FILLER_46_1722 ();
 sg13g2_decap_8 FILLER_46_1729 ();
 sg13g2_decap_8 FILLER_46_1736 ();
 sg13g2_decap_8 FILLER_46_1743 ();
 sg13g2_decap_8 FILLER_46_1750 ();
 sg13g2_decap_8 FILLER_46_1757 ();
 sg13g2_decap_4 FILLER_46_1764 ();
 sg13g2_fill_2 FILLER_47_54 ();
 sg13g2_fill_1 FILLER_47_83 ();
 sg13g2_fill_2 FILLER_47_93 ();
 sg13g2_fill_2 FILLER_47_104 ();
 sg13g2_fill_1 FILLER_47_106 ();
 sg13g2_fill_1 FILLER_47_116 ();
 sg13g2_fill_2 FILLER_47_135 ();
 sg13g2_fill_2 FILLER_47_141 ();
 sg13g2_fill_1 FILLER_47_151 ();
 sg13g2_fill_2 FILLER_47_158 ();
 sg13g2_fill_1 FILLER_47_184 ();
 sg13g2_fill_2 FILLER_47_289 ();
 sg13g2_fill_1 FILLER_47_291 ();
 sg13g2_fill_1 FILLER_47_311 ();
 sg13g2_fill_2 FILLER_47_330 ();
 sg13g2_decap_4 FILLER_47_350 ();
 sg13g2_fill_2 FILLER_47_354 ();
 sg13g2_decap_8 FILLER_47_360 ();
 sg13g2_fill_1 FILLER_47_367 ();
 sg13g2_decap_4 FILLER_47_394 ();
 sg13g2_fill_1 FILLER_47_425 ();
 sg13g2_fill_2 FILLER_47_472 ();
 sg13g2_fill_1 FILLER_47_474 ();
 sg13g2_decap_4 FILLER_47_500 ();
 sg13g2_fill_1 FILLER_47_504 ();
 sg13g2_fill_1 FILLER_47_522 ();
 sg13g2_fill_1 FILLER_47_530 ();
 sg13g2_fill_2 FILLER_47_570 ();
 sg13g2_decap_4 FILLER_47_578 ();
 sg13g2_fill_2 FILLER_47_613 ();
 sg13g2_fill_1 FILLER_47_639 ();
 sg13g2_fill_1 FILLER_47_677 ();
 sg13g2_fill_1 FILLER_47_687 ();
 sg13g2_fill_2 FILLER_47_712 ();
 sg13g2_fill_2 FILLER_47_731 ();
 sg13g2_fill_1 FILLER_47_739 ();
 sg13g2_fill_1 FILLER_47_746 ();
 sg13g2_decap_8 FILLER_47_758 ();
 sg13g2_fill_1 FILLER_47_765 ();
 sg13g2_fill_1 FILLER_47_826 ();
 sg13g2_fill_2 FILLER_47_836 ();
 sg13g2_decap_4 FILLER_47_894 ();
 sg13g2_fill_1 FILLER_47_898 ();
 sg13g2_fill_2 FILLER_47_918 ();
 sg13g2_fill_1 FILLER_47_920 ();
 sg13g2_fill_1 FILLER_47_963 ();
 sg13g2_fill_2 FILLER_47_986 ();
 sg13g2_fill_1 FILLER_47_995 ();
 sg13g2_fill_1 FILLER_47_1000 ();
 sg13g2_fill_2 FILLER_47_1018 ();
 sg13g2_fill_1 FILLER_47_1020 ();
 sg13g2_fill_2 FILLER_47_1062 ();
 sg13g2_fill_2 FILLER_47_1076 ();
 sg13g2_fill_2 FILLER_47_1112 ();
 sg13g2_fill_1 FILLER_47_1114 ();
 sg13g2_fill_1 FILLER_47_1184 ();
 sg13g2_fill_1 FILLER_47_1199 ();
 sg13g2_fill_1 FILLER_47_1209 ();
 sg13g2_fill_2 FILLER_47_1245 ();
 sg13g2_fill_2 FILLER_47_1273 ();
 sg13g2_fill_1 FILLER_47_1301 ();
 sg13g2_fill_2 FILLER_47_1332 ();
 sg13g2_fill_2 FILLER_47_1487 ();
 sg13g2_fill_1 FILLER_47_1523 ();
 sg13g2_fill_1 FILLER_47_1528 ();
 sg13g2_fill_2 FILLER_47_1547 ();
 sg13g2_fill_1 FILLER_47_1549 ();
 sg13g2_fill_2 FILLER_47_1567 ();
 sg13g2_fill_2 FILLER_47_1574 ();
 sg13g2_fill_1 FILLER_47_1576 ();
 sg13g2_fill_1 FILLER_47_1590 ();
 sg13g2_fill_1 FILLER_47_1622 ();
 sg13g2_decap_4 FILLER_47_1627 ();
 sg13g2_decap_8 FILLER_47_1635 ();
 sg13g2_decap_8 FILLER_47_1642 ();
 sg13g2_decap_8 FILLER_47_1649 ();
 sg13g2_decap_8 FILLER_47_1656 ();
 sg13g2_decap_8 FILLER_47_1663 ();
 sg13g2_decap_8 FILLER_47_1670 ();
 sg13g2_decap_8 FILLER_47_1677 ();
 sg13g2_decap_8 FILLER_47_1684 ();
 sg13g2_decap_8 FILLER_47_1691 ();
 sg13g2_decap_8 FILLER_47_1698 ();
 sg13g2_decap_8 FILLER_47_1705 ();
 sg13g2_decap_8 FILLER_47_1712 ();
 sg13g2_decap_8 FILLER_47_1719 ();
 sg13g2_decap_8 FILLER_47_1726 ();
 sg13g2_decap_8 FILLER_47_1733 ();
 sg13g2_decap_8 FILLER_47_1740 ();
 sg13g2_decap_8 FILLER_47_1747 ();
 sg13g2_decap_8 FILLER_47_1754 ();
 sg13g2_decap_8 FILLER_47_1761 ();
 sg13g2_fill_2 FILLER_48_121 ();
 sg13g2_fill_1 FILLER_48_156 ();
 sg13g2_fill_2 FILLER_48_176 ();
 sg13g2_fill_1 FILLER_48_183 ();
 sg13g2_fill_2 FILLER_48_205 ();
 sg13g2_fill_2 FILLER_48_246 ();
 sg13g2_fill_1 FILLER_48_252 ();
 sg13g2_fill_1 FILLER_48_302 ();
 sg13g2_fill_1 FILLER_48_329 ();
 sg13g2_fill_1 FILLER_48_335 ();
 sg13g2_decap_4 FILLER_48_367 ();
 sg13g2_fill_2 FILLER_48_380 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_2 FILLER_48_434 ();
 sg13g2_fill_2 FILLER_48_501 ();
 sg13g2_decap_8 FILLER_48_508 ();
 sg13g2_fill_1 FILLER_48_515 ();
 sg13g2_fill_1 FILLER_48_521 ();
 sg13g2_fill_2 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_530 ();
 sg13g2_fill_2 FILLER_48_537 ();
 sg13g2_fill_1 FILLER_48_558 ();
 sg13g2_fill_2 FILLER_48_574 ();
 sg13g2_fill_2 FILLER_48_624 ();
 sg13g2_decap_8 FILLER_48_639 ();
 sg13g2_fill_1 FILLER_48_646 ();
 sg13g2_fill_2 FILLER_48_673 ();
 sg13g2_fill_1 FILLER_48_675 ();
 sg13g2_fill_1 FILLER_48_691 ();
 sg13g2_fill_1 FILLER_48_711 ();
 sg13g2_fill_1 FILLER_48_718 ();
 sg13g2_fill_1 FILLER_48_752 ();
 sg13g2_fill_1 FILLER_48_779 ();
 sg13g2_fill_2 FILLER_48_807 ();
 sg13g2_fill_2 FILLER_48_817 ();
 sg13g2_fill_2 FILLER_48_832 ();
 sg13g2_fill_1 FILLER_48_851 ();
 sg13g2_decap_4 FILLER_48_907 ();
 sg13g2_fill_1 FILLER_48_923 ();
 sg13g2_fill_1 FILLER_48_937 ();
 sg13g2_fill_2 FILLER_48_947 ();
 sg13g2_fill_1 FILLER_48_949 ();
 sg13g2_fill_2 FILLER_48_955 ();
 sg13g2_fill_1 FILLER_48_972 ();
 sg13g2_fill_1 FILLER_48_994 ();
 sg13g2_fill_2 FILLER_48_1013 ();
 sg13g2_fill_1 FILLER_48_1015 ();
 sg13g2_fill_2 FILLER_48_1021 ();
 sg13g2_fill_1 FILLER_48_1034 ();
 sg13g2_fill_2 FILLER_48_1044 ();
 sg13g2_fill_1 FILLER_48_1064 ();
 sg13g2_fill_1 FILLER_48_1095 ();
 sg13g2_fill_1 FILLER_48_1149 ();
 sg13g2_fill_1 FILLER_48_1197 ();
 sg13g2_fill_2 FILLER_48_1213 ();
 sg13g2_fill_2 FILLER_48_1229 ();
 sg13g2_fill_2 FILLER_48_1237 ();
 sg13g2_fill_2 FILLER_48_1276 ();
 sg13g2_fill_1 FILLER_48_1278 ();
 sg13g2_fill_2 FILLER_48_1288 ();
 sg13g2_fill_1 FILLER_48_1342 ();
 sg13g2_fill_2 FILLER_48_1381 ();
 sg13g2_fill_2 FILLER_48_1418 ();
 sg13g2_fill_1 FILLER_48_1420 ();
 sg13g2_fill_1 FILLER_48_1467 ();
 sg13g2_fill_2 FILLER_48_1481 ();
 sg13g2_fill_2 FILLER_48_1488 ();
 sg13g2_fill_2 FILLER_48_1556 ();
 sg13g2_fill_1 FILLER_48_1558 ();
 sg13g2_fill_1 FILLER_48_1569 ();
 sg13g2_fill_1 FILLER_48_1596 ();
 sg13g2_fill_2 FILLER_48_1632 ();
 sg13g2_fill_1 FILLER_48_1634 ();
 sg13g2_decap_8 FILLER_48_1644 ();
 sg13g2_decap_8 FILLER_48_1651 ();
 sg13g2_decap_8 FILLER_48_1658 ();
 sg13g2_decap_8 FILLER_48_1665 ();
 sg13g2_decap_8 FILLER_48_1672 ();
 sg13g2_decap_8 FILLER_48_1679 ();
 sg13g2_decap_8 FILLER_48_1686 ();
 sg13g2_decap_8 FILLER_48_1693 ();
 sg13g2_decap_8 FILLER_48_1700 ();
 sg13g2_decap_8 FILLER_48_1707 ();
 sg13g2_decap_8 FILLER_48_1714 ();
 sg13g2_decap_8 FILLER_48_1721 ();
 sg13g2_decap_8 FILLER_48_1728 ();
 sg13g2_decap_8 FILLER_48_1735 ();
 sg13g2_decap_8 FILLER_48_1742 ();
 sg13g2_decap_8 FILLER_48_1749 ();
 sg13g2_decap_8 FILLER_48_1756 ();
 sg13g2_decap_4 FILLER_48_1763 ();
 sg13g2_fill_1 FILLER_48_1767 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_77 ();
 sg13g2_fill_1 FILLER_49_106 ();
 sg13g2_fill_2 FILLER_49_147 ();
 sg13g2_fill_2 FILLER_49_168 ();
 sg13g2_fill_2 FILLER_49_186 ();
 sg13g2_fill_1 FILLER_49_214 ();
 sg13g2_fill_2 FILLER_49_230 ();
 sg13g2_fill_2 FILLER_49_237 ();
 sg13g2_fill_2 FILLER_49_280 ();
 sg13g2_fill_1 FILLER_49_313 ();
 sg13g2_decap_4 FILLER_49_340 ();
 sg13g2_decap_8 FILLER_49_374 ();
 sg13g2_fill_2 FILLER_49_381 ();
 sg13g2_fill_1 FILLER_49_383 ();
 sg13g2_fill_2 FILLER_49_410 ();
 sg13g2_fill_2 FILLER_49_431 ();
 sg13g2_fill_1 FILLER_49_444 ();
 sg13g2_fill_2 FILLER_49_453 ();
 sg13g2_fill_1 FILLER_49_455 ();
 sg13g2_fill_2 FILLER_49_477 ();
 sg13g2_fill_1 FILLER_49_479 ();
 sg13g2_fill_2 FILLER_49_485 ();
 sg13g2_fill_1 FILLER_49_492 ();
 sg13g2_fill_2 FILLER_49_501 ();
 sg13g2_fill_2 FILLER_49_514 ();
 sg13g2_fill_1 FILLER_49_516 ();
 sg13g2_fill_2 FILLER_49_557 ();
 sg13g2_decap_8 FILLER_49_569 ();
 sg13g2_fill_1 FILLER_49_594 ();
 sg13g2_fill_2 FILLER_49_628 ();
 sg13g2_fill_1 FILLER_49_630 ();
 sg13g2_decap_8 FILLER_49_636 ();
 sg13g2_fill_2 FILLER_49_643 ();
 sg13g2_fill_1 FILLER_49_645 ();
 sg13g2_fill_2 FILLER_49_670 ();
 sg13g2_fill_1 FILLER_49_672 ();
 sg13g2_fill_2 FILLER_49_699 ();
 sg13g2_fill_1 FILLER_49_701 ();
 sg13g2_fill_1 FILLER_49_705 ();
 sg13g2_fill_1 FILLER_49_714 ();
 sg13g2_decap_8 FILLER_49_739 ();
 sg13g2_decap_4 FILLER_49_749 ();
 sg13g2_fill_2 FILLER_49_757 ();
 sg13g2_fill_1 FILLER_49_770 ();
 sg13g2_fill_2 FILLER_49_812 ();
 sg13g2_fill_1 FILLER_49_814 ();
 sg13g2_fill_2 FILLER_49_856 ();
 sg13g2_fill_2 FILLER_49_876 ();
 sg13g2_fill_1 FILLER_49_878 ();
 sg13g2_fill_2 FILLER_49_888 ();
 sg13g2_fill_1 FILLER_49_890 ();
 sg13g2_fill_2 FILLER_49_904 ();
 sg13g2_fill_1 FILLER_49_906 ();
 sg13g2_fill_2 FILLER_49_985 ();
 sg13g2_fill_1 FILLER_49_1013 ();
 sg13g2_fill_1 FILLER_49_1018 ();
 sg13g2_fill_2 FILLER_49_1063 ();
 sg13g2_fill_1 FILLER_49_1065 ();
 sg13g2_fill_2 FILLER_49_1077 ();
 sg13g2_fill_1 FILLER_49_1079 ();
 sg13g2_fill_1 FILLER_49_1089 ();
 sg13g2_fill_2 FILLER_49_1098 ();
 sg13g2_fill_2 FILLER_49_1127 ();
 sg13g2_fill_1 FILLER_49_1129 ();
 sg13g2_fill_1 FILLER_49_1160 ();
 sg13g2_fill_1 FILLER_49_1171 ();
 sg13g2_fill_2 FILLER_49_1220 ();
 sg13g2_fill_2 FILLER_49_1284 ();
 sg13g2_fill_2 FILLER_49_1330 ();
 sg13g2_fill_1 FILLER_49_1337 ();
 sg13g2_fill_2 FILLER_49_1388 ();
 sg13g2_fill_1 FILLER_49_1407 ();
 sg13g2_fill_1 FILLER_49_1429 ();
 sg13g2_fill_2 FILLER_49_1486 ();
 sg13g2_fill_2 FILLER_49_1498 ();
 sg13g2_fill_1 FILLER_49_1519 ();
 sg13g2_fill_2 FILLER_49_1545 ();
 sg13g2_fill_1 FILLER_49_1547 ();
 sg13g2_fill_1 FILLER_49_1557 ();
 sg13g2_fill_2 FILLER_49_1576 ();
 sg13g2_fill_2 FILLER_49_1613 ();
 sg13g2_decap_8 FILLER_49_1646 ();
 sg13g2_decap_8 FILLER_49_1653 ();
 sg13g2_decap_8 FILLER_49_1660 ();
 sg13g2_decap_8 FILLER_49_1667 ();
 sg13g2_decap_8 FILLER_49_1674 ();
 sg13g2_decap_8 FILLER_49_1681 ();
 sg13g2_decap_8 FILLER_49_1688 ();
 sg13g2_decap_8 FILLER_49_1695 ();
 sg13g2_decap_8 FILLER_49_1702 ();
 sg13g2_decap_8 FILLER_49_1709 ();
 sg13g2_decap_8 FILLER_49_1716 ();
 sg13g2_decap_8 FILLER_49_1723 ();
 sg13g2_decap_8 FILLER_49_1730 ();
 sg13g2_decap_8 FILLER_49_1737 ();
 sg13g2_decap_8 FILLER_49_1744 ();
 sg13g2_decap_8 FILLER_49_1751 ();
 sg13g2_decap_8 FILLER_49_1758 ();
 sg13g2_fill_2 FILLER_49_1765 ();
 sg13g2_fill_1 FILLER_49_1767 ();
 sg13g2_fill_1 FILLER_50_149 ();
 sg13g2_fill_2 FILLER_50_163 ();
 sg13g2_fill_1 FILLER_50_180 ();
 sg13g2_fill_2 FILLER_50_207 ();
 sg13g2_fill_2 FILLER_50_276 ();
 sg13g2_fill_2 FILLER_50_287 ();
 sg13g2_fill_1 FILLER_50_298 ();
 sg13g2_decap_8 FILLER_50_329 ();
 sg13g2_decap_8 FILLER_50_336 ();
 sg13g2_fill_2 FILLER_50_365 ();
 sg13g2_fill_2 FILLER_50_376 ();
 sg13g2_fill_1 FILLER_50_412 ();
 sg13g2_fill_1 FILLER_50_418 ();
 sg13g2_decap_8 FILLER_50_432 ();
 sg13g2_fill_1 FILLER_50_439 ();
 sg13g2_decap_4 FILLER_50_453 ();
 sg13g2_fill_1 FILLER_50_457 ();
 sg13g2_decap_8 FILLER_50_466 ();
 sg13g2_fill_2 FILLER_50_473 ();
 sg13g2_fill_2 FILLER_50_504 ();
 sg13g2_fill_1 FILLER_50_506 ();
 sg13g2_fill_1 FILLER_50_533 ();
 sg13g2_decap_8 FILLER_50_553 ();
 sg13g2_decap_8 FILLER_50_560 ();
 sg13g2_decap_8 FILLER_50_567 ();
 sg13g2_fill_1 FILLER_50_593 ();
 sg13g2_fill_2 FILLER_50_648 ();
 sg13g2_fill_1 FILLER_50_650 ();
 sg13g2_fill_1 FILLER_50_695 ();
 sg13g2_decap_8 FILLER_50_712 ();
 sg13g2_fill_2 FILLER_50_719 ();
 sg13g2_fill_1 FILLER_50_721 ();
 sg13g2_fill_2 FILLER_50_731 ();
 sg13g2_fill_1 FILLER_50_773 ();
 sg13g2_fill_2 FILLER_50_782 ();
 sg13g2_fill_1 FILLER_50_847 ();
 sg13g2_fill_1 FILLER_50_911 ();
 sg13g2_fill_1 FILLER_50_923 ();
 sg13g2_fill_2 FILLER_50_929 ();
 sg13g2_fill_1 FILLER_50_931 ();
 sg13g2_fill_2 FILLER_50_951 ();
 sg13g2_fill_1 FILLER_50_953 ();
 sg13g2_fill_2 FILLER_50_960 ();
 sg13g2_decap_4 FILLER_50_970 ();
 sg13g2_fill_1 FILLER_50_974 ();
 sg13g2_decap_4 FILLER_50_983 ();
 sg13g2_fill_2 FILLER_50_1016 ();
 sg13g2_fill_1 FILLER_50_1018 ();
 sg13g2_fill_2 FILLER_50_1027 ();
 sg13g2_fill_1 FILLER_50_1062 ();
 sg13g2_fill_2 FILLER_50_1093 ();
 sg13g2_fill_1 FILLER_50_1095 ();
 sg13g2_fill_1 FILLER_50_1126 ();
 sg13g2_fill_2 FILLER_50_1135 ();
 sg13g2_fill_1 FILLER_50_1137 ();
 sg13g2_fill_2 FILLER_50_1148 ();
 sg13g2_fill_1 FILLER_50_1150 ();
 sg13g2_fill_1 FILLER_50_1165 ();
 sg13g2_fill_1 FILLER_50_1231 ();
 sg13g2_fill_2 FILLER_50_1261 ();
 sg13g2_fill_1 FILLER_50_1263 ();
 sg13g2_fill_1 FILLER_50_1278 ();
 sg13g2_fill_2 FILLER_50_1309 ();
 sg13g2_fill_1 FILLER_50_1311 ();
 sg13g2_fill_2 FILLER_50_1442 ();
 sg13g2_fill_1 FILLER_50_1444 ();
 sg13g2_fill_2 FILLER_50_1477 ();
 sg13g2_fill_1 FILLER_50_1479 ();
 sg13g2_fill_2 FILLER_50_1552 ();
 sg13g2_fill_1 FILLER_50_1554 ();
 sg13g2_fill_2 FILLER_50_1581 ();
 sg13g2_fill_2 FILLER_50_1588 ();
 sg13g2_fill_1 FILLER_50_1590 ();
 sg13g2_fill_2 FILLER_50_1605 ();
 sg13g2_fill_2 FILLER_50_1626 ();
 sg13g2_decap_8 FILLER_50_1658 ();
 sg13g2_decap_8 FILLER_50_1665 ();
 sg13g2_decap_8 FILLER_50_1672 ();
 sg13g2_decap_8 FILLER_50_1679 ();
 sg13g2_decap_8 FILLER_50_1686 ();
 sg13g2_decap_8 FILLER_50_1693 ();
 sg13g2_decap_8 FILLER_50_1700 ();
 sg13g2_decap_8 FILLER_50_1707 ();
 sg13g2_decap_8 FILLER_50_1714 ();
 sg13g2_decap_8 FILLER_50_1721 ();
 sg13g2_decap_8 FILLER_50_1728 ();
 sg13g2_decap_8 FILLER_50_1735 ();
 sg13g2_decap_8 FILLER_50_1742 ();
 sg13g2_decap_8 FILLER_50_1749 ();
 sg13g2_decap_8 FILLER_50_1756 ();
 sg13g2_decap_4 FILLER_50_1763 ();
 sg13g2_fill_1 FILLER_50_1767 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_43 ();
 sg13g2_fill_2 FILLER_51_121 ();
 sg13g2_fill_1 FILLER_51_131 ();
 sg13g2_fill_2 FILLER_51_146 ();
 sg13g2_fill_2 FILLER_51_165 ();
 sg13g2_fill_2 FILLER_51_175 ();
 sg13g2_fill_2 FILLER_51_274 ();
 sg13g2_fill_2 FILLER_51_307 ();
 sg13g2_fill_1 FILLER_51_309 ();
 sg13g2_fill_1 FILLER_51_331 ();
 sg13g2_fill_2 FILLER_51_384 ();
 sg13g2_fill_2 FILLER_51_401 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_fill_1 FILLER_51_446 ();
 sg13g2_decap_4 FILLER_51_461 ();
 sg13g2_fill_2 FILLER_51_465 ();
 sg13g2_decap_4 FILLER_51_490 ();
 sg13g2_fill_1 FILLER_51_494 ();
 sg13g2_decap_8 FILLER_51_505 ();
 sg13g2_fill_1 FILLER_51_512 ();
 sg13g2_fill_2 FILLER_51_530 ();
 sg13g2_fill_1 FILLER_51_532 ();
 sg13g2_decap_8 FILLER_51_536 ();
 sg13g2_fill_2 FILLER_51_543 ();
 sg13g2_fill_1 FILLER_51_545 ();
 sg13g2_fill_2 FILLER_51_581 ();
 sg13g2_fill_2 FILLER_51_593 ();
 sg13g2_fill_1 FILLER_51_595 ();
 sg13g2_decap_4 FILLER_51_602 ();
 sg13g2_decap_4 FILLER_51_622 ();
 sg13g2_decap_8 FILLER_51_632 ();
 sg13g2_fill_2 FILLER_51_644 ();
 sg13g2_fill_2 FILLER_51_665 ();
 sg13g2_fill_1 FILLER_51_679 ();
 sg13g2_fill_1 FILLER_51_748 ();
 sg13g2_fill_2 FILLER_51_767 ();
 sg13g2_fill_2 FILLER_51_818 ();
 sg13g2_fill_2 FILLER_51_836 ();
 sg13g2_fill_1 FILLER_51_875 ();
 sg13g2_decap_4 FILLER_51_880 ();
 sg13g2_fill_2 FILLER_51_884 ();
 sg13g2_fill_2 FILLER_51_907 ();
 sg13g2_decap_8 FILLER_51_939 ();
 sg13g2_fill_2 FILLER_51_946 ();
 sg13g2_fill_1 FILLER_51_948 ();
 sg13g2_fill_2 FILLER_51_990 ();
 sg13g2_fill_1 FILLER_51_992 ();
 sg13g2_fill_2 FILLER_51_999 ();
 sg13g2_fill_1 FILLER_51_1001 ();
 sg13g2_fill_2 FILLER_51_1007 ();
 sg13g2_fill_1 FILLER_51_1022 ();
 sg13g2_fill_2 FILLER_51_1031 ();
 sg13g2_fill_1 FILLER_51_1033 ();
 sg13g2_fill_1 FILLER_51_1047 ();
 sg13g2_fill_1 FILLER_51_1053 ();
 sg13g2_fill_1 FILLER_51_1085 ();
 sg13g2_fill_1 FILLER_51_1137 ();
 sg13g2_fill_1 FILLER_51_1169 ();
 sg13g2_fill_1 FILLER_51_1184 ();
 sg13g2_fill_1 FILLER_51_1234 ();
 sg13g2_fill_2 FILLER_51_1282 ();
 sg13g2_fill_2 FILLER_51_1293 ();
 sg13g2_fill_2 FILLER_51_1309 ();
 sg13g2_fill_1 FILLER_51_1311 ();
 sg13g2_fill_2 FILLER_51_1366 ();
 sg13g2_fill_2 FILLER_51_1382 ();
 sg13g2_fill_2 FILLER_51_1405 ();
 sg13g2_fill_1 FILLER_51_1407 ();
 sg13g2_fill_1 FILLER_51_1439 ();
 sg13g2_fill_2 FILLER_51_1483 ();
 sg13g2_fill_1 FILLER_51_1485 ();
 sg13g2_fill_2 FILLER_51_1503 ();
 sg13g2_fill_1 FILLER_51_1505 ();
 sg13g2_fill_1 FILLER_51_1510 ();
 sg13g2_fill_1 FILLER_51_1525 ();
 sg13g2_fill_2 FILLER_51_1532 ();
 sg13g2_fill_1 FILLER_51_1534 ();
 sg13g2_fill_2 FILLER_51_1578 ();
 sg13g2_fill_1 FILLER_51_1580 ();
 sg13g2_decap_8 FILLER_51_1664 ();
 sg13g2_decap_8 FILLER_51_1671 ();
 sg13g2_decap_8 FILLER_51_1678 ();
 sg13g2_decap_8 FILLER_51_1685 ();
 sg13g2_decap_8 FILLER_51_1692 ();
 sg13g2_decap_8 FILLER_51_1699 ();
 sg13g2_decap_8 FILLER_51_1706 ();
 sg13g2_decap_8 FILLER_51_1713 ();
 sg13g2_decap_8 FILLER_51_1720 ();
 sg13g2_decap_8 FILLER_51_1727 ();
 sg13g2_decap_8 FILLER_51_1734 ();
 sg13g2_decap_8 FILLER_51_1741 ();
 sg13g2_decap_8 FILLER_51_1748 ();
 sg13g2_decap_8 FILLER_51_1755 ();
 sg13g2_decap_4 FILLER_51_1762 ();
 sg13g2_fill_2 FILLER_51_1766 ();
 sg13g2_fill_2 FILLER_52_90 ();
 sg13g2_fill_1 FILLER_52_92 ();
 sg13g2_fill_2 FILLER_52_122 ();
 sg13g2_fill_1 FILLER_52_154 ();
 sg13g2_fill_1 FILLER_52_158 ();
 sg13g2_fill_1 FILLER_52_165 ();
 sg13g2_fill_2 FILLER_52_183 ();
 sg13g2_fill_1 FILLER_52_198 ();
 sg13g2_fill_2 FILLER_52_221 ();
 sg13g2_fill_2 FILLER_52_236 ();
 sg13g2_fill_2 FILLER_52_251 ();
 sg13g2_fill_2 FILLER_52_267 ();
 sg13g2_fill_1 FILLER_52_303 ();
 sg13g2_fill_1 FILLER_52_309 ();
 sg13g2_fill_1 FILLER_52_399 ();
 sg13g2_fill_2 FILLER_52_405 ();
 sg13g2_fill_2 FILLER_52_441 ();
 sg13g2_fill_1 FILLER_52_443 ();
 sg13g2_fill_1 FILLER_52_454 ();
 sg13g2_fill_2 FILLER_52_506 ();
 sg13g2_fill_1 FILLER_52_531 ();
 sg13g2_fill_1 FILLER_52_564 ();
 sg13g2_fill_2 FILLER_52_583 ();
 sg13g2_fill_2 FILLER_52_611 ();
 sg13g2_decap_4 FILLER_52_668 ();
 sg13g2_fill_2 FILLER_52_672 ();
 sg13g2_fill_2 FILLER_52_682 ();
 sg13g2_fill_1 FILLER_52_684 ();
 sg13g2_decap_4 FILLER_52_693 ();
 sg13g2_fill_1 FILLER_52_720 ();
 sg13g2_fill_1 FILLER_52_740 ();
 sg13g2_fill_2 FILLER_52_760 ();
 sg13g2_fill_2 FILLER_52_772 ();
 sg13g2_fill_1 FILLER_52_779 ();
 sg13g2_fill_2 FILLER_52_785 ();
 sg13g2_decap_4 FILLER_52_796 ();
 sg13g2_fill_2 FILLER_52_829 ();
 sg13g2_fill_1 FILLER_52_831 ();
 sg13g2_fill_1 FILLER_52_845 ();
 sg13g2_fill_2 FILLER_52_860 ();
 sg13g2_fill_1 FILLER_52_862 ();
 sg13g2_fill_2 FILLER_52_874 ();
 sg13g2_fill_1 FILLER_52_881 ();
 sg13g2_fill_1 FILLER_52_897 ();
 sg13g2_fill_2 FILLER_52_906 ();
 sg13g2_fill_1 FILLER_52_912 ();
 sg13g2_fill_2 FILLER_52_937 ();
 sg13g2_fill_1 FILLER_52_939 ();
 sg13g2_fill_1 FILLER_52_961 ();
 sg13g2_fill_1 FILLER_52_988 ();
 sg13g2_fill_2 FILLER_52_994 ();
 sg13g2_decap_4 FILLER_52_1001 ();
 sg13g2_fill_1 FILLER_52_1005 ();
 sg13g2_fill_1 FILLER_52_1032 ();
 sg13g2_fill_2 FILLER_52_1038 ();
 sg13g2_fill_2 FILLER_52_1045 ();
 sg13g2_fill_2 FILLER_52_1124 ();
 sg13g2_fill_1 FILLER_52_1126 ();
 sg13g2_fill_1 FILLER_52_1152 ();
 sg13g2_fill_1 FILLER_52_1158 ();
 sg13g2_fill_1 FILLER_52_1185 ();
 sg13g2_fill_1 FILLER_52_1229 ();
 sg13g2_fill_2 FILLER_52_1325 ();
 sg13g2_fill_2 FILLER_52_1362 ();
 sg13g2_fill_1 FILLER_52_1364 ();
 sg13g2_fill_2 FILLER_52_1418 ();
 sg13g2_fill_2 FILLER_52_1450 ();
 sg13g2_fill_2 FILLER_52_1466 ();
 sg13g2_fill_1 FILLER_52_1468 ();
 sg13g2_fill_2 FILLER_52_1507 ();
 sg13g2_fill_1 FILLER_52_1509 ();
 sg13g2_fill_1 FILLER_52_1523 ();
 sg13g2_fill_1 FILLER_52_1554 ();
 sg13g2_fill_1 FILLER_52_1590 ();
 sg13g2_fill_2 FILLER_52_1600 ();
 sg13g2_fill_2 FILLER_52_1623 ();
 sg13g2_fill_1 FILLER_52_1625 ();
 sg13g2_decap_8 FILLER_52_1666 ();
 sg13g2_decap_8 FILLER_52_1673 ();
 sg13g2_decap_8 FILLER_52_1680 ();
 sg13g2_decap_8 FILLER_52_1687 ();
 sg13g2_decap_8 FILLER_52_1694 ();
 sg13g2_decap_8 FILLER_52_1701 ();
 sg13g2_decap_8 FILLER_52_1708 ();
 sg13g2_decap_8 FILLER_52_1715 ();
 sg13g2_decap_8 FILLER_52_1722 ();
 sg13g2_decap_8 FILLER_52_1729 ();
 sg13g2_decap_8 FILLER_52_1736 ();
 sg13g2_decap_8 FILLER_52_1743 ();
 sg13g2_decap_8 FILLER_52_1750 ();
 sg13g2_decap_8 FILLER_52_1757 ();
 sg13g2_decap_4 FILLER_52_1764 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_265 ();
 sg13g2_decap_4 FILLER_53_364 ();
 sg13g2_decap_8 FILLER_53_386 ();
 sg13g2_decap_4 FILLER_53_393 ();
 sg13g2_fill_1 FILLER_53_397 ();
 sg13g2_fill_2 FILLER_53_403 ();
 sg13g2_fill_1 FILLER_53_405 ();
 sg13g2_decap_4 FILLER_53_421 ();
 sg13g2_fill_1 FILLER_53_425 ();
 sg13g2_fill_2 FILLER_53_441 ();
 sg13g2_fill_1 FILLER_53_453 ();
 sg13g2_fill_2 FILLER_53_474 ();
 sg13g2_decap_4 FILLER_53_484 ();
 sg13g2_fill_1 FILLER_53_514 ();
 sg13g2_fill_2 FILLER_53_524 ();
 sg13g2_decap_8 FILLER_53_541 ();
 sg13g2_fill_2 FILLER_53_548 ();
 sg13g2_fill_1 FILLER_53_565 ();
 sg13g2_fill_2 FILLER_53_582 ();
 sg13g2_fill_2 FILLER_53_602 ();
 sg13g2_decap_8 FILLER_53_612 ();
 sg13g2_fill_1 FILLER_53_635 ();
 sg13g2_fill_2 FILLER_53_649 ();
 sg13g2_fill_1 FILLER_53_651 ();
 sg13g2_fill_1 FILLER_53_657 ();
 sg13g2_fill_2 FILLER_53_675 ();
 sg13g2_decap_4 FILLER_53_684 ();
 sg13g2_fill_2 FILLER_53_704 ();
 sg13g2_fill_2 FILLER_53_712 ();
 sg13g2_fill_1 FILLER_53_714 ();
 sg13g2_fill_2 FILLER_53_728 ();
 sg13g2_fill_2 FILLER_53_758 ();
 sg13g2_fill_2 FILLER_53_779 ();
 sg13g2_fill_2 FILLER_53_789 ();
 sg13g2_fill_1 FILLER_53_791 ();
 sg13g2_fill_1 FILLER_53_824 ();
 sg13g2_fill_1 FILLER_53_899 ();
 sg13g2_fill_1 FILLER_53_910 ();
 sg13g2_fill_2 FILLER_53_916 ();
 sg13g2_fill_2 FILLER_53_940 ();
 sg13g2_fill_1 FILLER_53_955 ();
 sg13g2_fill_2 FILLER_53_961 ();
 sg13g2_fill_1 FILLER_53_963 ();
 sg13g2_decap_4 FILLER_53_981 ();
 sg13g2_fill_1 FILLER_53_985 ();
 sg13g2_fill_2 FILLER_53_1003 ();
 sg13g2_fill_2 FILLER_53_1060 ();
 sg13g2_fill_1 FILLER_53_1062 ();
 sg13g2_fill_2 FILLER_53_1085 ();
 sg13g2_fill_2 FILLER_53_1126 ();
 sg13g2_fill_1 FILLER_53_1128 ();
 sg13g2_fill_1 FILLER_53_1169 ();
 sg13g2_fill_2 FILLER_53_1175 ();
 sg13g2_fill_1 FILLER_53_1189 ();
 sg13g2_fill_2 FILLER_53_1219 ();
 sg13g2_fill_1 FILLER_53_1221 ();
 sg13g2_fill_1 FILLER_53_1230 ();
 sg13g2_fill_2 FILLER_53_1269 ();
 sg13g2_fill_2 FILLER_53_1276 ();
 sg13g2_fill_1 FILLER_53_1341 ();
 sg13g2_fill_2 FILLER_53_1372 ();
 sg13g2_fill_1 FILLER_53_1374 ();
 sg13g2_fill_2 FILLER_53_1427 ();
 sg13g2_fill_1 FILLER_53_1495 ();
 sg13g2_fill_1 FILLER_53_1545 ();
 sg13g2_fill_1 FILLER_53_1629 ();
 sg13g2_fill_1 FILLER_53_1635 ();
 sg13g2_decap_8 FILLER_53_1666 ();
 sg13g2_decap_8 FILLER_53_1673 ();
 sg13g2_decap_8 FILLER_53_1680 ();
 sg13g2_decap_8 FILLER_53_1687 ();
 sg13g2_decap_8 FILLER_53_1694 ();
 sg13g2_decap_8 FILLER_53_1701 ();
 sg13g2_decap_8 FILLER_53_1708 ();
 sg13g2_decap_8 FILLER_53_1715 ();
 sg13g2_decap_8 FILLER_53_1722 ();
 sg13g2_decap_8 FILLER_53_1729 ();
 sg13g2_decap_8 FILLER_53_1736 ();
 sg13g2_decap_8 FILLER_53_1743 ();
 sg13g2_decap_8 FILLER_53_1750 ();
 sg13g2_decap_8 FILLER_53_1757 ();
 sg13g2_decap_4 FILLER_53_1764 ();
 sg13g2_fill_1 FILLER_54_110 ();
 sg13g2_fill_1 FILLER_54_144 ();
 sg13g2_fill_1 FILLER_54_160 ();
 sg13g2_decap_8 FILLER_54_166 ();
 sg13g2_fill_2 FILLER_54_173 ();
 sg13g2_fill_1 FILLER_54_275 ();
 sg13g2_fill_2 FILLER_54_306 ();
 sg13g2_decap_4 FILLER_54_343 ();
 sg13g2_fill_2 FILLER_54_373 ();
 sg13g2_fill_1 FILLER_54_390 ();
 sg13g2_fill_1 FILLER_54_417 ();
 sg13g2_decap_8 FILLER_54_423 ();
 sg13g2_fill_2 FILLER_54_430 ();
 sg13g2_fill_1 FILLER_54_432 ();
 sg13g2_decap_4 FILLER_54_444 ();
 sg13g2_fill_1 FILLER_54_456 ();
 sg13g2_decap_8 FILLER_54_478 ();
 sg13g2_decap_8 FILLER_54_485 ();
 sg13g2_fill_1 FILLER_54_504 ();
 sg13g2_decap_8 FILLER_54_513 ();
 sg13g2_decap_4 FILLER_54_520 ();
 sg13g2_decap_4 FILLER_54_536 ();
 sg13g2_fill_2 FILLER_54_540 ();
 sg13g2_fill_1 FILLER_54_592 ();
 sg13g2_decap_8 FILLER_54_597 ();
 sg13g2_fill_2 FILLER_54_604 ();
 sg13g2_fill_2 FILLER_54_622 ();
 sg13g2_fill_1 FILLER_54_624 ();
 sg13g2_fill_2 FILLER_54_633 ();
 sg13g2_fill_1 FILLER_54_643 ();
 sg13g2_fill_2 FILLER_54_683 ();
 sg13g2_fill_1 FILLER_54_685 ();
 sg13g2_fill_2 FILLER_54_701 ();
 sg13g2_fill_1 FILLER_54_703 ();
 sg13g2_fill_2 FILLER_54_712 ();
 sg13g2_fill_1 FILLER_54_714 ();
 sg13g2_decap_8 FILLER_54_720 ();
 sg13g2_decap_4 FILLER_54_727 ();
 sg13g2_fill_1 FILLER_54_731 ();
 sg13g2_fill_2 FILLER_54_777 ();
 sg13g2_fill_2 FILLER_54_788 ();
 sg13g2_fill_1 FILLER_54_790 ();
 sg13g2_fill_2 FILLER_54_795 ();
 sg13g2_fill_1 FILLER_54_797 ();
 sg13g2_fill_1 FILLER_54_832 ();
 sg13g2_fill_2 FILLER_54_840 ();
 sg13g2_fill_1 FILLER_54_881 ();
 sg13g2_fill_1 FILLER_54_895 ();
 sg13g2_fill_1 FILLER_54_901 ();
 sg13g2_fill_1 FILLER_54_933 ();
 sg13g2_fill_2 FILLER_54_938 ();
 sg13g2_fill_1 FILLER_54_984 ();
 sg13g2_fill_2 FILLER_54_1006 ();
 sg13g2_fill_2 FILLER_54_1017 ();
 sg13g2_fill_1 FILLER_54_1019 ();
 sg13g2_fill_2 FILLER_54_1033 ();
 sg13g2_fill_1 FILLER_54_1035 ();
 sg13g2_fill_1 FILLER_54_1047 ();
 sg13g2_fill_1 FILLER_54_1054 ();
 sg13g2_fill_1 FILLER_54_1070 ();
 sg13g2_fill_2 FILLER_54_1088 ();
 sg13g2_fill_2 FILLER_54_1148 ();
 sg13g2_fill_2 FILLER_54_1225 ();
 sg13g2_fill_2 FILLER_54_1266 ();
 sg13g2_fill_1 FILLER_54_1273 ();
 sg13g2_fill_2 FILLER_54_1330 ();
 sg13g2_fill_1 FILLER_54_1342 ();
 sg13g2_fill_1 FILLER_54_1370 ();
 sg13g2_fill_1 FILLER_54_1388 ();
 sg13g2_fill_2 FILLER_54_1398 ();
 sg13g2_fill_2 FILLER_54_1409 ();
 sg13g2_fill_1 FILLER_54_1450 ();
 sg13g2_fill_1 FILLER_54_1467 ();
 sg13g2_fill_2 FILLER_54_1589 ();
 sg13g2_fill_1 FILLER_54_1591 ();
 sg13g2_fill_1 FILLER_54_1637 ();
 sg13g2_decap_8 FILLER_54_1672 ();
 sg13g2_decap_8 FILLER_54_1679 ();
 sg13g2_decap_8 FILLER_54_1686 ();
 sg13g2_decap_8 FILLER_54_1693 ();
 sg13g2_decap_8 FILLER_54_1700 ();
 sg13g2_decap_8 FILLER_54_1707 ();
 sg13g2_decap_8 FILLER_54_1714 ();
 sg13g2_decap_8 FILLER_54_1721 ();
 sg13g2_decap_8 FILLER_54_1728 ();
 sg13g2_decap_8 FILLER_54_1735 ();
 sg13g2_decap_8 FILLER_54_1742 ();
 sg13g2_decap_8 FILLER_54_1749 ();
 sg13g2_decap_8 FILLER_54_1756 ();
 sg13g2_decap_4 FILLER_54_1763 ();
 sg13g2_fill_1 FILLER_54_1767 ();
 sg13g2_fill_1 FILLER_55_65 ();
 sg13g2_fill_1 FILLER_55_98 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_fill_2 FILLER_55_140 ();
 sg13g2_fill_1 FILLER_55_142 ();
 sg13g2_decap_4 FILLER_55_182 ();
 sg13g2_fill_1 FILLER_55_186 ();
 sg13g2_fill_1 FILLER_55_249 ();
 sg13g2_fill_2 FILLER_55_262 ();
 sg13g2_fill_2 FILLER_55_294 ();
 sg13g2_fill_1 FILLER_55_327 ();
 sg13g2_fill_2 FILLER_55_354 ();
 sg13g2_fill_1 FILLER_55_356 ();
 sg13g2_decap_4 FILLER_55_361 ();
 sg13g2_fill_1 FILLER_55_365 ();
 sg13g2_decap_8 FILLER_55_408 ();
 sg13g2_fill_1 FILLER_55_451 ();
 sg13g2_fill_1 FILLER_55_464 ();
 sg13g2_fill_2 FILLER_55_480 ();
 sg13g2_fill_1 FILLER_55_482 ();
 sg13g2_fill_2 FILLER_55_494 ();
 sg13g2_fill_2 FILLER_55_501 ();
 sg13g2_fill_1 FILLER_55_513 ();
 sg13g2_fill_2 FILLER_55_555 ();
 sg13g2_fill_1 FILLER_55_557 ();
 sg13g2_fill_1 FILLER_55_573 ();
 sg13g2_fill_1 FILLER_55_608 ();
 sg13g2_fill_2 FILLER_55_623 ();
 sg13g2_fill_2 FILLER_55_662 ();
 sg13g2_fill_2 FILLER_55_704 ();
 sg13g2_decap_4 FILLER_55_731 ();
 sg13g2_fill_1 FILLER_55_735 ();
 sg13g2_fill_2 FILLER_55_752 ();
 sg13g2_fill_2 FILLER_55_788 ();
 sg13g2_decap_4 FILLER_55_798 ();
 sg13g2_fill_2 FILLER_55_802 ();
 sg13g2_decap_4 FILLER_55_830 ();
 sg13g2_fill_2 FILLER_55_860 ();
 sg13g2_fill_1 FILLER_55_862 ();
 sg13g2_fill_2 FILLER_55_882 ();
 sg13g2_fill_2 FILLER_55_900 ();
 sg13g2_decap_8 FILLER_55_928 ();
 sg13g2_fill_1 FILLER_55_935 ();
 sg13g2_decap_4 FILLER_55_962 ();
 sg13g2_fill_2 FILLER_55_966 ();
 sg13g2_decap_4 FILLER_55_982 ();
 sg13g2_decap_8 FILLER_55_1012 ();
 sg13g2_fill_2 FILLER_55_1019 ();
 sg13g2_fill_2 FILLER_55_1029 ();
 sg13g2_fill_1 FILLER_55_1031 ();
 sg13g2_fill_2 FILLER_55_1036 ();
 sg13g2_fill_1 FILLER_55_1038 ();
 sg13g2_fill_2 FILLER_55_1043 ();
 sg13g2_decap_4 FILLER_55_1059 ();
 sg13g2_fill_2 FILLER_55_1070 ();
 sg13g2_fill_1 FILLER_55_1072 ();
 sg13g2_fill_1 FILLER_55_1078 ();
 sg13g2_fill_2 FILLER_55_1143 ();
 sg13g2_fill_2 FILLER_55_1149 ();
 sg13g2_fill_1 FILLER_55_1151 ();
 sg13g2_fill_1 FILLER_55_1232 ();
 sg13g2_fill_2 FILLER_55_1242 ();
 sg13g2_fill_2 FILLER_55_1250 ();
 sg13g2_fill_1 FILLER_55_1300 ();
 sg13g2_fill_2 FILLER_55_1329 ();
 sg13g2_fill_1 FILLER_55_1458 ();
 sg13g2_fill_2 FILLER_55_1479 ();
 sg13g2_fill_1 FILLER_55_1507 ();
 sg13g2_fill_2 FILLER_55_1533 ();
 sg13g2_fill_1 FILLER_55_1535 ();
 sg13g2_fill_2 FILLER_55_1546 ();
 sg13g2_fill_1 FILLER_55_1585 ();
 sg13g2_fill_1 FILLER_55_1590 ();
 sg13g2_fill_2 FILLER_55_1596 ();
 sg13g2_fill_1 FILLER_55_1598 ();
 sg13g2_fill_2 FILLER_55_1642 ();
 sg13g2_decap_8 FILLER_55_1678 ();
 sg13g2_decap_8 FILLER_55_1685 ();
 sg13g2_decap_8 FILLER_55_1692 ();
 sg13g2_decap_8 FILLER_55_1699 ();
 sg13g2_decap_8 FILLER_55_1706 ();
 sg13g2_decap_8 FILLER_55_1713 ();
 sg13g2_decap_8 FILLER_55_1720 ();
 sg13g2_decap_8 FILLER_55_1727 ();
 sg13g2_decap_8 FILLER_55_1734 ();
 sg13g2_decap_8 FILLER_55_1741 ();
 sg13g2_decap_8 FILLER_55_1748 ();
 sg13g2_decap_8 FILLER_55_1755 ();
 sg13g2_decap_4 FILLER_55_1762 ();
 sg13g2_fill_2 FILLER_55_1766 ();
 sg13g2_fill_2 FILLER_56_83 ();
 sg13g2_fill_2 FILLER_56_134 ();
 sg13g2_fill_1 FILLER_56_136 ();
 sg13g2_fill_1 FILLER_56_176 ();
 sg13g2_fill_1 FILLER_56_213 ();
 sg13g2_fill_1 FILLER_56_246 ();
 sg13g2_fill_2 FILLER_56_337 ();
 sg13g2_decap_4 FILLER_56_346 ();
 sg13g2_fill_2 FILLER_56_350 ();
 sg13g2_fill_1 FILLER_56_388 ();
 sg13g2_fill_1 FILLER_56_425 ();
 sg13g2_decap_8 FILLER_56_508 ();
 sg13g2_decap_4 FILLER_56_515 ();
 sg13g2_fill_1 FILLER_56_519 ();
 sg13g2_fill_1 FILLER_56_534 ();
 sg13g2_decap_4 FILLER_56_543 ();
 sg13g2_fill_2 FILLER_56_558 ();
 sg13g2_fill_1 FILLER_56_560 ();
 sg13g2_fill_1 FILLER_56_602 ();
 sg13g2_decap_4 FILLER_56_624 ();
 sg13g2_fill_2 FILLER_56_628 ();
 sg13g2_fill_1 FILLER_56_685 ();
 sg13g2_fill_2 FILLER_56_703 ();
 sg13g2_fill_2 FILLER_56_730 ();
 sg13g2_fill_1 FILLER_56_779 ();
 sg13g2_fill_2 FILLER_56_811 ();
 sg13g2_fill_1 FILLER_56_813 ();
 sg13g2_decap_4 FILLER_56_821 ();
 sg13g2_fill_2 FILLER_56_834 ();
 sg13g2_fill_1 FILLER_56_836 ();
 sg13g2_decap_8 FILLER_56_882 ();
 sg13g2_decap_4 FILLER_56_889 ();
 sg13g2_fill_1 FILLER_56_893 ();
 sg13g2_fill_1 FILLER_56_899 ();
 sg13g2_decap_4 FILLER_56_909 ();
 sg13g2_fill_2 FILLER_56_917 ();
 sg13g2_fill_1 FILLER_56_919 ();
 sg13g2_decap_4 FILLER_56_938 ();
 sg13g2_fill_2 FILLER_56_942 ();
 sg13g2_fill_1 FILLER_56_959 ();
 sg13g2_fill_1 FILLER_56_974 ();
 sg13g2_fill_2 FILLER_56_994 ();
 sg13g2_fill_1 FILLER_56_996 ();
 sg13g2_fill_2 FILLER_56_1001 ();
 sg13g2_fill_1 FILLER_56_1003 ();
 sg13g2_fill_2 FILLER_56_1130 ();
 sg13g2_fill_2 FILLER_56_1174 ();
 sg13g2_fill_2 FILLER_56_1256 ();
 sg13g2_fill_2 FILLER_56_1301 ();
 sg13g2_fill_1 FILLER_56_1303 ();
 sg13g2_fill_1 FILLER_56_1384 ();
 sg13g2_fill_2 FILLER_56_1399 ();
 sg13g2_fill_1 FILLER_56_1406 ();
 sg13g2_fill_1 FILLER_56_1416 ();
 sg13g2_fill_2 FILLER_56_1441 ();
 sg13g2_fill_1 FILLER_56_1443 ();
 sg13g2_fill_2 FILLER_56_1453 ();
 sg13g2_fill_1 FILLER_56_1455 ();
 sg13g2_fill_1 FILLER_56_1469 ();
 sg13g2_fill_1 FILLER_56_1544 ();
 sg13g2_fill_1 FILLER_56_1567 ();
 sg13g2_fill_2 FILLER_56_1615 ();
 sg13g2_fill_2 FILLER_56_1621 ();
 sg13g2_fill_1 FILLER_56_1623 ();
 sg13g2_fill_1 FILLER_56_1629 ();
 sg13g2_fill_2 FILLER_56_1635 ();
 sg13g2_decap_8 FILLER_56_1672 ();
 sg13g2_decap_8 FILLER_56_1679 ();
 sg13g2_decap_8 FILLER_56_1686 ();
 sg13g2_decap_8 FILLER_56_1693 ();
 sg13g2_decap_8 FILLER_56_1700 ();
 sg13g2_decap_8 FILLER_56_1707 ();
 sg13g2_decap_8 FILLER_56_1714 ();
 sg13g2_decap_8 FILLER_56_1721 ();
 sg13g2_decap_8 FILLER_56_1728 ();
 sg13g2_decap_8 FILLER_56_1735 ();
 sg13g2_decap_8 FILLER_56_1742 ();
 sg13g2_decap_8 FILLER_56_1749 ();
 sg13g2_decap_8 FILLER_56_1756 ();
 sg13g2_decap_4 FILLER_56_1763 ();
 sg13g2_fill_1 FILLER_56_1767 ();
 sg13g2_fill_2 FILLER_57_82 ();
 sg13g2_fill_1 FILLER_57_122 ();
 sg13g2_fill_2 FILLER_57_154 ();
 sg13g2_fill_2 FILLER_57_182 ();
 sg13g2_fill_2 FILLER_57_204 ();
 sg13g2_fill_1 FILLER_57_206 ();
 sg13g2_decap_8 FILLER_57_351 ();
 sg13g2_fill_1 FILLER_57_366 ();
 sg13g2_fill_1 FILLER_57_402 ();
 sg13g2_decap_8 FILLER_57_407 ();
 sg13g2_fill_1 FILLER_57_424 ();
 sg13g2_fill_1 FILLER_57_430 ();
 sg13g2_fill_1 FILLER_57_445 ();
 sg13g2_fill_2 FILLER_57_456 ();
 sg13g2_decap_8 FILLER_57_482 ();
 sg13g2_decap_4 FILLER_57_489 ();
 sg13g2_decap_8 FILLER_57_497 ();
 sg13g2_fill_2 FILLER_57_544 ();
 sg13g2_fill_2 FILLER_57_563 ();
 sg13g2_fill_1 FILLER_57_565 ();
 sg13g2_fill_2 FILLER_57_624 ();
 sg13g2_fill_2 FILLER_57_651 ();
 sg13g2_fill_2 FILLER_57_670 ();
 sg13g2_fill_1 FILLER_57_707 ();
 sg13g2_decap_8 FILLER_57_723 ();
 sg13g2_decap_8 FILLER_57_730 ();
 sg13g2_decap_4 FILLER_57_740 ();
 sg13g2_fill_1 FILLER_57_774 ();
 sg13g2_decap_4 FILLER_57_778 ();
 sg13g2_fill_2 FILLER_57_782 ();
 sg13g2_fill_2 FILLER_57_792 ();
 sg13g2_fill_1 FILLER_57_794 ();
 sg13g2_fill_1 FILLER_57_806 ();
 sg13g2_fill_2 FILLER_57_812 ();
 sg13g2_fill_1 FILLER_57_814 ();
 sg13g2_decap_4 FILLER_57_835 ();
 sg13g2_decap_4 FILLER_57_857 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_fill_2 FILLER_57_866 ();
 sg13g2_fill_1 FILLER_57_868 ();
 sg13g2_decap_4 FILLER_57_885 ();
 sg13g2_fill_2 FILLER_57_889 ();
 sg13g2_fill_2 FILLER_57_910 ();
 sg13g2_fill_1 FILLER_57_912 ();
 sg13g2_decap_4 FILLER_57_933 ();
 sg13g2_fill_2 FILLER_57_937 ();
 sg13g2_fill_2 FILLER_57_944 ();
 sg13g2_fill_1 FILLER_57_946 ();
 sg13g2_decap_8 FILLER_57_968 ();
 sg13g2_decap_4 FILLER_57_980 ();
 sg13g2_decap_8 FILLER_57_995 ();
 sg13g2_fill_2 FILLER_57_1002 ();
 sg13g2_fill_2 FILLER_57_1037 ();
 sg13g2_decap_8 FILLER_57_1110 ();
 sg13g2_decap_4 FILLER_57_1121 ();
 sg13g2_decap_4 FILLER_57_1147 ();
 sg13g2_decap_4 FILLER_57_1177 ();
 sg13g2_fill_1 FILLER_57_1181 ();
 sg13g2_fill_1 FILLER_57_1248 ();
 sg13g2_fill_2 FILLER_57_1312 ();
 sg13g2_fill_1 FILLER_57_1420 ();
 sg13g2_fill_2 FILLER_57_1445 ();
 sg13g2_fill_2 FILLER_57_1465 ();
 sg13g2_fill_1 FILLER_57_1467 ();
 sg13g2_fill_2 FILLER_57_1503 ();
 sg13g2_fill_1 FILLER_57_1505 ();
 sg13g2_fill_1 FILLER_57_1514 ();
 sg13g2_fill_2 FILLER_57_1546 ();
 sg13g2_fill_1 FILLER_57_1548 ();
 sg13g2_decap_8 FILLER_57_1669 ();
 sg13g2_decap_8 FILLER_57_1676 ();
 sg13g2_decap_8 FILLER_57_1683 ();
 sg13g2_decap_8 FILLER_57_1690 ();
 sg13g2_decap_8 FILLER_57_1697 ();
 sg13g2_decap_8 FILLER_57_1704 ();
 sg13g2_decap_8 FILLER_57_1711 ();
 sg13g2_decap_8 FILLER_57_1718 ();
 sg13g2_decap_8 FILLER_57_1725 ();
 sg13g2_decap_8 FILLER_57_1732 ();
 sg13g2_decap_8 FILLER_57_1739 ();
 sg13g2_decap_8 FILLER_57_1746 ();
 sg13g2_decap_8 FILLER_57_1753 ();
 sg13g2_decap_8 FILLER_57_1760 ();
 sg13g2_fill_1 FILLER_57_1767 ();
 sg13g2_fill_1 FILLER_58_26 ();
 sg13g2_fill_2 FILLER_58_75 ();
 sg13g2_fill_1 FILLER_58_77 ();
 sg13g2_fill_2 FILLER_58_140 ();
 sg13g2_fill_2 FILLER_58_176 ();
 sg13g2_fill_2 FILLER_58_214 ();
 sg13g2_fill_1 FILLER_58_216 ();
 sg13g2_fill_2 FILLER_58_284 ();
 sg13g2_fill_1 FILLER_58_335 ();
 sg13g2_decap_4 FILLER_58_373 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_fill_2 FILLER_58_383 ();
 sg13g2_fill_2 FILLER_58_437 ();
 sg13g2_fill_2 FILLER_58_466 ();
 sg13g2_fill_1 FILLER_58_468 ();
 sg13g2_fill_2 FILLER_58_477 ();
 sg13g2_fill_2 FILLER_58_484 ();
 sg13g2_fill_2 FILLER_58_503 ();
 sg13g2_fill_1 FILLER_58_527 ();
 sg13g2_fill_1 FILLER_58_546 ();
 sg13g2_decap_4 FILLER_58_553 ();
 sg13g2_fill_2 FILLER_58_557 ();
 sg13g2_fill_1 FILLER_58_591 ();
 sg13g2_fill_2 FILLER_58_607 ();
 sg13g2_fill_1 FILLER_58_609 ();
 sg13g2_fill_2 FILLER_58_672 ();
 sg13g2_fill_2 FILLER_58_705 ();
 sg13g2_fill_2 FILLER_58_737 ();
 sg13g2_fill_1 FILLER_58_768 ();
 sg13g2_decap_4 FILLER_58_784 ();
 sg13g2_decap_8 FILLER_58_796 ();
 sg13g2_decap_4 FILLER_58_808 ();
 sg13g2_fill_1 FILLER_58_835 ();
 sg13g2_decap_4 FILLER_58_910 ();
 sg13g2_fill_2 FILLER_58_947 ();
 sg13g2_fill_1 FILLER_58_949 ();
 sg13g2_fill_2 FILLER_58_956 ();
 sg13g2_decap_4 FILLER_58_973 ();
 sg13g2_fill_1 FILLER_58_977 ();
 sg13g2_fill_2 FILLER_58_987 ();
 sg13g2_fill_1 FILLER_58_989 ();
 sg13g2_fill_1 FILLER_58_994 ();
 sg13g2_fill_2 FILLER_58_1003 ();
 sg13g2_fill_2 FILLER_58_1011 ();
 sg13g2_fill_1 FILLER_58_1021 ();
 sg13g2_decap_4 FILLER_58_1049 ();
 sg13g2_fill_1 FILLER_58_1053 ();
 sg13g2_fill_1 FILLER_58_1075 ();
 sg13g2_decap_8 FILLER_58_1081 ();
 sg13g2_fill_2 FILLER_58_1088 ();
 sg13g2_fill_1 FILLER_58_1090 ();
 sg13g2_fill_1 FILLER_58_1095 ();
 sg13g2_fill_2 FILLER_58_1150 ();
 sg13g2_fill_1 FILLER_58_1152 ();
 sg13g2_fill_2 FILLER_58_1184 ();
 sg13g2_fill_2 FILLER_58_1217 ();
 sg13g2_fill_1 FILLER_58_1219 ();
 sg13g2_fill_1 FILLER_58_1230 ();
 sg13g2_fill_2 FILLER_58_1239 ();
 sg13g2_fill_1 FILLER_58_1272 ();
 sg13g2_fill_2 FILLER_58_1283 ();
 sg13g2_fill_1 FILLER_58_1285 ();
 sg13g2_fill_1 FILLER_58_1332 ();
 sg13g2_fill_2 FILLER_58_1363 ();
 sg13g2_fill_1 FILLER_58_1365 ();
 sg13g2_fill_2 FILLER_58_1415 ();
 sg13g2_fill_1 FILLER_58_1453 ();
 sg13g2_decap_4 FILLER_58_1468 ();
 sg13g2_fill_1 FILLER_58_1472 ();
 sg13g2_decap_4 FILLER_58_1482 ();
 sg13g2_fill_2 FILLER_58_1526 ();
 sg13g2_fill_2 FILLER_58_1566 ();
 sg13g2_fill_2 FILLER_58_1591 ();
 sg13g2_fill_1 FILLER_58_1593 ();
 sg13g2_fill_1 FILLER_58_1616 ();
 sg13g2_decap_8 FILLER_58_1661 ();
 sg13g2_decap_8 FILLER_58_1668 ();
 sg13g2_decap_8 FILLER_58_1675 ();
 sg13g2_decap_8 FILLER_58_1682 ();
 sg13g2_decap_8 FILLER_58_1689 ();
 sg13g2_decap_8 FILLER_58_1696 ();
 sg13g2_decap_8 FILLER_58_1703 ();
 sg13g2_decap_8 FILLER_58_1710 ();
 sg13g2_decap_8 FILLER_58_1717 ();
 sg13g2_decap_8 FILLER_58_1724 ();
 sg13g2_decap_8 FILLER_58_1731 ();
 sg13g2_decap_8 FILLER_58_1738 ();
 sg13g2_decap_8 FILLER_58_1745 ();
 sg13g2_decap_8 FILLER_58_1752 ();
 sg13g2_decap_8 FILLER_58_1759 ();
 sg13g2_fill_2 FILLER_58_1766 ();
 sg13g2_fill_2 FILLER_59_35 ();
 sg13g2_fill_1 FILLER_59_47 ();
 sg13g2_fill_2 FILLER_59_145 ();
 sg13g2_fill_1 FILLER_59_147 ();
 sg13g2_fill_1 FILLER_59_156 ();
 sg13g2_fill_1 FILLER_59_203 ();
 sg13g2_decap_4 FILLER_59_208 ();
 sg13g2_fill_2 FILLER_59_212 ();
 sg13g2_fill_2 FILLER_59_224 ();
 sg13g2_fill_1 FILLER_59_226 ();
 sg13g2_fill_2 FILLER_59_262 ();
 sg13g2_fill_2 FILLER_59_321 ();
 sg13g2_fill_2 FILLER_59_357 ();
 sg13g2_fill_2 FILLER_59_368 ();
 sg13g2_fill_1 FILLER_59_383 ();
 sg13g2_fill_2 FILLER_59_397 ();
 sg13g2_decap_8 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_417 ();
 sg13g2_decap_4 FILLER_59_426 ();
 sg13g2_decap_4 FILLER_59_484 ();
 sg13g2_fill_2 FILLER_59_488 ();
 sg13g2_fill_1 FILLER_59_493 ();
 sg13g2_fill_2 FILLER_59_507 ();
 sg13g2_fill_2 FILLER_59_557 ();
 sg13g2_fill_1 FILLER_59_631 ();
 sg13g2_fill_1 FILLER_59_640 ();
 sg13g2_fill_1 FILLER_59_645 ();
 sg13g2_fill_2 FILLER_59_651 ();
 sg13g2_fill_2 FILLER_59_708 ();
 sg13g2_fill_1 FILLER_59_760 ();
 sg13g2_fill_1 FILLER_59_786 ();
 sg13g2_decap_4 FILLER_59_791 ();
 sg13g2_fill_1 FILLER_59_795 ();
 sg13g2_fill_1 FILLER_59_800 ();
 sg13g2_fill_2 FILLER_59_820 ();
 sg13g2_fill_1 FILLER_59_851 ();
 sg13g2_fill_2 FILLER_59_867 ();
 sg13g2_fill_1 FILLER_59_869 ();
 sg13g2_fill_2 FILLER_59_883 ();
 sg13g2_fill_1 FILLER_59_885 ();
 sg13g2_fill_2 FILLER_59_897 ();
 sg13g2_fill_2 FILLER_59_911 ();
 sg13g2_fill_1 FILLER_59_913 ();
 sg13g2_fill_1 FILLER_59_918 ();
 sg13g2_fill_2 FILLER_59_924 ();
 sg13g2_fill_1 FILLER_59_943 ();
 sg13g2_decap_8 FILLER_59_979 ();
 sg13g2_fill_1 FILLER_59_1025 ();
 sg13g2_fill_2 FILLER_59_1038 ();
 sg13g2_fill_1 FILLER_59_1044 ();
 sg13g2_fill_2 FILLER_59_1054 ();
 sg13g2_fill_1 FILLER_59_1056 ();
 sg13g2_decap_4 FILLER_59_1062 ();
 sg13g2_fill_1 FILLER_59_1071 ();
 sg13g2_fill_2 FILLER_59_1092 ();
 sg13g2_fill_2 FILLER_59_1133 ();
 sg13g2_fill_2 FILLER_59_1155 ();
 sg13g2_fill_2 FILLER_59_1165 ();
 sg13g2_fill_2 FILLER_59_1234 ();
 sg13g2_fill_1 FILLER_59_1236 ();
 sg13g2_fill_1 FILLER_59_1254 ();
 sg13g2_fill_2 FILLER_59_1261 ();
 sg13g2_fill_1 FILLER_59_1263 ();
 sg13g2_fill_2 FILLER_59_1296 ();
 sg13g2_fill_2 FILLER_59_1302 ();
 sg13g2_fill_1 FILLER_59_1323 ();
 sg13g2_fill_2 FILLER_59_1342 ();
 sg13g2_fill_1 FILLER_59_1357 ();
 sg13g2_fill_2 FILLER_59_1366 ();
 sg13g2_decap_4 FILLER_59_1497 ();
 sg13g2_decap_8 FILLER_59_1509 ();
 sg13g2_fill_1 FILLER_59_1516 ();
 sg13g2_fill_2 FILLER_59_1522 ();
 sg13g2_fill_1 FILLER_59_1524 ();
 sg13g2_fill_2 FILLER_59_1544 ();
 sg13g2_fill_1 FILLER_59_1546 ();
 sg13g2_fill_2 FILLER_59_1622 ();
 sg13g2_fill_2 FILLER_59_1633 ();
 sg13g2_fill_1 FILLER_59_1635 ();
 sg13g2_decap_8 FILLER_59_1658 ();
 sg13g2_decap_8 FILLER_59_1665 ();
 sg13g2_decap_8 FILLER_59_1672 ();
 sg13g2_decap_8 FILLER_59_1679 ();
 sg13g2_decap_8 FILLER_59_1686 ();
 sg13g2_decap_8 FILLER_59_1693 ();
 sg13g2_decap_8 FILLER_59_1700 ();
 sg13g2_decap_8 FILLER_59_1707 ();
 sg13g2_decap_8 FILLER_59_1714 ();
 sg13g2_decap_8 FILLER_59_1721 ();
 sg13g2_decap_8 FILLER_59_1728 ();
 sg13g2_decap_8 FILLER_59_1735 ();
 sg13g2_decap_8 FILLER_59_1742 ();
 sg13g2_decap_8 FILLER_59_1749 ();
 sg13g2_decap_8 FILLER_59_1756 ();
 sg13g2_decap_4 FILLER_59_1763 ();
 sg13g2_fill_1 FILLER_59_1767 ();
 sg13g2_fill_2 FILLER_60_67 ();
 sg13g2_decap_4 FILLER_60_181 ();
 sg13g2_fill_1 FILLER_60_185 ();
 sg13g2_fill_2 FILLER_60_191 ();
 sg13g2_fill_1 FILLER_60_193 ();
 sg13g2_fill_2 FILLER_60_211 ();
 sg13g2_fill_2 FILLER_60_261 ();
 sg13g2_fill_1 FILLER_60_263 ();
 sg13g2_fill_1 FILLER_60_268 ();
 sg13g2_fill_2 FILLER_60_306 ();
 sg13g2_fill_1 FILLER_60_317 ();
 sg13g2_fill_1 FILLER_60_323 ();
 sg13g2_fill_1 FILLER_60_352 ();
 sg13g2_fill_2 FILLER_60_373 ();
 sg13g2_fill_2 FILLER_60_427 ();
 sg13g2_fill_1 FILLER_60_429 ();
 sg13g2_decap_4 FILLER_60_441 ();
 sg13g2_decap_4 FILLER_60_453 ();
 sg13g2_fill_2 FILLER_60_457 ();
 sg13g2_fill_2 FILLER_60_464 ();
 sg13g2_fill_2 FILLER_60_509 ();
 sg13g2_fill_1 FILLER_60_511 ();
 sg13g2_fill_2 FILLER_60_549 ();
 sg13g2_fill_1 FILLER_60_551 ();
 sg13g2_fill_1 FILLER_60_560 ();
 sg13g2_fill_2 FILLER_60_571 ();
 sg13g2_decap_4 FILLER_60_590 ();
 sg13g2_fill_2 FILLER_60_594 ();
 sg13g2_fill_2 FILLER_60_610 ();
 sg13g2_fill_1 FILLER_60_612 ();
 sg13g2_decap_4 FILLER_60_631 ();
 sg13g2_decap_4 FILLER_60_639 ();
 sg13g2_fill_1 FILLER_60_643 ();
 sg13g2_fill_1 FILLER_60_662 ();
 sg13g2_fill_2 FILLER_60_692 ();
 sg13g2_fill_2 FILLER_60_699 ();
 sg13g2_fill_1 FILLER_60_706 ();
 sg13g2_fill_2 FILLER_60_718 ();
 sg13g2_decap_4 FILLER_60_725 ();
 sg13g2_decap_8 FILLER_60_764 ();
 sg13g2_decap_8 FILLER_60_771 ();
 sg13g2_fill_1 FILLER_60_778 ();
 sg13g2_fill_1 FILLER_60_797 ();
 sg13g2_fill_2 FILLER_60_803 ();
 sg13g2_fill_1 FILLER_60_805 ();
 sg13g2_fill_2 FILLER_60_821 ();
 sg13g2_fill_2 FILLER_60_828 ();
 sg13g2_decap_4 FILLER_60_839 ();
 sg13g2_fill_1 FILLER_60_843 ();
 sg13g2_fill_2 FILLER_60_849 ();
 sg13g2_fill_1 FILLER_60_851 ();
 sg13g2_fill_1 FILLER_60_862 ();
 sg13g2_fill_2 FILLER_60_867 ();
 sg13g2_fill_2 FILLER_60_873 ();
 sg13g2_decap_8 FILLER_60_887 ();
 sg13g2_decap_8 FILLER_60_894 ();
 sg13g2_decap_4 FILLER_60_901 ();
 sg13g2_fill_2 FILLER_60_905 ();
 sg13g2_fill_1 FILLER_60_936 ();
 sg13g2_fill_2 FILLER_60_949 ();
 sg13g2_fill_2 FILLER_60_981 ();
 sg13g2_fill_1 FILLER_60_983 ();
 sg13g2_fill_1 FILLER_60_998 ();
 sg13g2_fill_1 FILLER_60_1012 ();
 sg13g2_fill_1 FILLER_60_1021 ();
 sg13g2_fill_2 FILLER_60_1058 ();
 sg13g2_decap_4 FILLER_60_1071 ();
 sg13g2_fill_1 FILLER_60_1075 ();
 sg13g2_decap_4 FILLER_60_1080 ();
 sg13g2_fill_1 FILLER_60_1088 ();
 sg13g2_fill_2 FILLER_60_1098 ();
 sg13g2_fill_1 FILLER_60_1123 ();
 sg13g2_fill_2 FILLER_60_1174 ();
 sg13g2_decap_8 FILLER_60_1181 ();
 sg13g2_fill_2 FILLER_60_1188 ();
 sg13g2_decap_8 FILLER_60_1194 ();
 sg13g2_fill_2 FILLER_60_1201 ();
 sg13g2_fill_1 FILLER_60_1219 ();
 sg13g2_fill_2 FILLER_60_1264 ();
 sg13g2_fill_1 FILLER_60_1284 ();
 sg13g2_fill_1 FILLER_60_1294 ();
 sg13g2_fill_2 FILLER_60_1304 ();
 sg13g2_fill_1 FILLER_60_1324 ();
 sg13g2_fill_2 FILLER_60_1355 ();
 sg13g2_fill_1 FILLER_60_1391 ();
 sg13g2_fill_2 FILLER_60_1422 ();
 sg13g2_fill_2 FILLER_60_1442 ();
 sg13g2_fill_1 FILLER_60_1444 ();
 sg13g2_fill_2 FILLER_60_1453 ();
 sg13g2_fill_1 FILLER_60_1455 ();
 sg13g2_fill_2 FILLER_60_1467 ();
 sg13g2_fill_2 FILLER_60_1477 ();
 sg13g2_fill_1 FILLER_60_1492 ();
 sg13g2_decap_8 FILLER_60_1506 ();
 sg13g2_decap_4 FILLER_60_1513 ();
 sg13g2_fill_1 FILLER_60_1517 ();
 sg13g2_fill_1 FILLER_60_1547 ();
 sg13g2_fill_2 FILLER_60_1569 ();
 sg13g2_fill_2 FILLER_60_1584 ();
 sg13g2_fill_1 FILLER_60_1586 ();
 sg13g2_fill_2 FILLER_60_1596 ();
 sg13g2_decap_8 FILLER_60_1664 ();
 sg13g2_decap_8 FILLER_60_1671 ();
 sg13g2_decap_8 FILLER_60_1678 ();
 sg13g2_decap_8 FILLER_60_1685 ();
 sg13g2_decap_8 FILLER_60_1692 ();
 sg13g2_decap_8 FILLER_60_1699 ();
 sg13g2_decap_8 FILLER_60_1706 ();
 sg13g2_decap_8 FILLER_60_1713 ();
 sg13g2_decap_8 FILLER_60_1720 ();
 sg13g2_decap_8 FILLER_60_1727 ();
 sg13g2_decap_8 FILLER_60_1734 ();
 sg13g2_decap_8 FILLER_60_1741 ();
 sg13g2_decap_8 FILLER_60_1748 ();
 sg13g2_decap_8 FILLER_60_1755 ();
 sg13g2_decap_4 FILLER_60_1762 ();
 sg13g2_fill_2 FILLER_60_1766 ();
 sg13g2_fill_2 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_37 ();
 sg13g2_fill_2 FILLER_61_47 ();
 sg13g2_fill_1 FILLER_61_49 ();
 sg13g2_fill_2 FILLER_61_71 ();
 sg13g2_fill_2 FILLER_61_146 ();
 sg13g2_fill_2 FILLER_61_170 ();
 sg13g2_decap_4 FILLER_61_196 ();
 sg13g2_fill_1 FILLER_61_210 ();
 sg13g2_fill_1 FILLER_61_240 ();
 sg13g2_fill_2 FILLER_61_259 ();
 sg13g2_fill_1 FILLER_61_292 ();
 sg13g2_fill_1 FILLER_61_393 ();
 sg13g2_fill_2 FILLER_61_411 ();
 sg13g2_fill_1 FILLER_61_413 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_fill_1 FILLER_61_430 ();
 sg13g2_fill_1 FILLER_61_441 ();
 sg13g2_fill_1 FILLER_61_463 ();
 sg13g2_fill_2 FILLER_61_477 ();
 sg13g2_fill_1 FILLER_61_479 ();
 sg13g2_fill_2 FILLER_61_502 ();
 sg13g2_fill_2 FILLER_61_530 ();
 sg13g2_fill_1 FILLER_61_536 ();
 sg13g2_fill_1 FILLER_61_567 ();
 sg13g2_fill_1 FILLER_61_586 ();
 sg13g2_fill_1 FILLER_61_613 ();
 sg13g2_fill_1 FILLER_61_619 ();
 sg13g2_fill_1 FILLER_61_668 ();
 sg13g2_decap_4 FILLER_61_736 ();
 sg13g2_decap_8 FILLER_61_756 ();
 sg13g2_decap_4 FILLER_61_837 ();
 sg13g2_fill_2 FILLER_61_841 ();
 sg13g2_fill_2 FILLER_61_879 ();
 sg13g2_decap_8 FILLER_61_898 ();
 sg13g2_decap_4 FILLER_61_905 ();
 sg13g2_fill_1 FILLER_61_953 ();
 sg13g2_decap_4 FILLER_61_971 ();
 sg13g2_fill_2 FILLER_61_975 ();
 sg13g2_fill_2 FILLER_61_996 ();
 sg13g2_fill_2 FILLER_61_1024 ();
 sg13g2_decap_4 FILLER_61_1054 ();
 sg13g2_fill_1 FILLER_61_1058 ();
 sg13g2_fill_2 FILLER_61_1063 ();
 sg13g2_fill_1 FILLER_61_1065 ();
 sg13g2_fill_2 FILLER_61_1143 ();
 sg13g2_decap_8 FILLER_61_1176 ();
 sg13g2_fill_1 FILLER_61_1183 ();
 sg13g2_decap_8 FILLER_61_1195 ();
 sg13g2_decap_4 FILLER_61_1215 ();
 sg13g2_fill_2 FILLER_61_1227 ();
 sg13g2_fill_1 FILLER_61_1281 ();
 sg13g2_fill_2 FILLER_61_1308 ();
 sg13g2_fill_2 FILLER_61_1350 ();
 sg13g2_fill_2 FILLER_61_1372 ();
 sg13g2_fill_2 FILLER_61_1410 ();
 sg13g2_fill_1 FILLER_61_1417 ();
 sg13g2_fill_2 FILLER_61_1460 ();
 sg13g2_fill_2 FILLER_61_1470 ();
 sg13g2_fill_1 FILLER_61_1489 ();
 sg13g2_fill_1 FILLER_61_1568 ();
 sg13g2_fill_1 FILLER_61_1621 ();
 sg13g2_fill_2 FILLER_61_1627 ();
 sg13g2_decap_8 FILLER_61_1667 ();
 sg13g2_decap_8 FILLER_61_1674 ();
 sg13g2_decap_8 FILLER_61_1681 ();
 sg13g2_decap_8 FILLER_61_1688 ();
 sg13g2_decap_8 FILLER_61_1695 ();
 sg13g2_decap_8 FILLER_61_1702 ();
 sg13g2_decap_8 FILLER_61_1709 ();
 sg13g2_decap_8 FILLER_61_1716 ();
 sg13g2_decap_8 FILLER_61_1723 ();
 sg13g2_decap_8 FILLER_61_1730 ();
 sg13g2_decap_8 FILLER_61_1737 ();
 sg13g2_decap_8 FILLER_61_1744 ();
 sg13g2_decap_8 FILLER_61_1751 ();
 sg13g2_decap_8 FILLER_61_1758 ();
 sg13g2_fill_2 FILLER_61_1765 ();
 sg13g2_fill_1 FILLER_61_1767 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_109 ();
 sg13g2_fill_1 FILLER_62_171 ();
 sg13g2_fill_1 FILLER_62_200 ();
 sg13g2_fill_2 FILLER_62_275 ();
 sg13g2_fill_2 FILLER_62_287 ();
 sg13g2_fill_2 FILLER_62_302 ();
 sg13g2_decap_8 FILLER_62_445 ();
 sg13g2_decap_4 FILLER_62_461 ();
 sg13g2_decap_8 FILLER_62_493 ();
 sg13g2_fill_1 FILLER_62_504 ();
 sg13g2_fill_2 FILLER_62_552 ();
 sg13g2_fill_1 FILLER_62_602 ();
 sg13g2_fill_2 FILLER_62_634 ();
 sg13g2_fill_2 FILLER_62_663 ();
 sg13g2_fill_1 FILLER_62_665 ();
 sg13g2_fill_2 FILLER_62_675 ();
 sg13g2_fill_1 FILLER_62_677 ();
 sg13g2_fill_2 FILLER_62_714 ();
 sg13g2_fill_1 FILLER_62_742 ();
 sg13g2_fill_2 FILLER_62_763 ();
 sg13g2_fill_2 FILLER_62_769 ();
 sg13g2_fill_2 FILLER_62_789 ();
 sg13g2_fill_2 FILLER_62_804 ();
 sg13g2_fill_1 FILLER_62_823 ();
 sg13g2_decap_8 FILLER_62_834 ();
 sg13g2_fill_1 FILLER_62_841 ();
 sg13g2_fill_2 FILLER_62_847 ();
 sg13g2_fill_2 FILLER_62_872 ();
 sg13g2_fill_1 FILLER_62_874 ();
 sg13g2_decap_8 FILLER_62_910 ();
 sg13g2_decap_8 FILLER_62_917 ();
 sg13g2_fill_1 FILLER_62_941 ();
 sg13g2_decap_8 FILLER_62_969 ();
 sg13g2_fill_2 FILLER_62_976 ();
 sg13g2_fill_1 FILLER_62_978 ();
 sg13g2_fill_1 FILLER_62_1008 ();
 sg13g2_fill_1 FILLER_62_1022 ();
 sg13g2_fill_2 FILLER_62_1048 ();
 sg13g2_fill_1 FILLER_62_1050 ();
 sg13g2_fill_1 FILLER_62_1062 ();
 sg13g2_decap_8 FILLER_62_1080 ();
 sg13g2_fill_2 FILLER_62_1087 ();
 sg13g2_fill_1 FILLER_62_1089 ();
 sg13g2_fill_2 FILLER_62_1111 ();
 sg13g2_fill_1 FILLER_62_1118 ();
 sg13g2_fill_2 FILLER_62_1222 ();
 sg13g2_fill_1 FILLER_62_1224 ();
 sg13g2_decap_4 FILLER_62_1233 ();
 sg13g2_fill_2 FILLER_62_1278 ();
 sg13g2_fill_1 FILLER_62_1280 ();
 sg13g2_fill_2 FILLER_62_1300 ();
 sg13g2_fill_1 FILLER_62_1302 ();
 sg13g2_fill_2 FILLER_62_1346 ();
 sg13g2_fill_1 FILLER_62_1348 ();
 sg13g2_fill_2 FILLER_62_1354 ();
 sg13g2_fill_2 FILLER_62_1369 ();
 sg13g2_fill_2 FILLER_62_1379 ();
 sg13g2_fill_2 FILLER_62_1407 ();
 sg13g2_fill_2 FILLER_62_1413 ();
 sg13g2_fill_1 FILLER_62_1415 ();
 sg13g2_fill_2 FILLER_62_1421 ();
 sg13g2_fill_1 FILLER_62_1423 ();
 sg13g2_fill_1 FILLER_62_1457 ();
 sg13g2_fill_2 FILLER_62_1463 ();
 sg13g2_fill_1 FILLER_62_1465 ();
 sg13g2_decap_8 FILLER_62_1496 ();
 sg13g2_fill_1 FILLER_62_1509 ();
 sg13g2_fill_2 FILLER_62_1515 ();
 sg13g2_fill_2 FILLER_62_1526 ();
 sg13g2_decap_4 FILLER_62_1538 ();
 sg13g2_fill_1 FILLER_62_1571 ();
 sg13g2_fill_2 FILLER_62_1595 ();
 sg13g2_fill_2 FILLER_62_1632 ();
 sg13g2_decap_8 FILLER_62_1669 ();
 sg13g2_decap_8 FILLER_62_1676 ();
 sg13g2_decap_8 FILLER_62_1683 ();
 sg13g2_decap_8 FILLER_62_1690 ();
 sg13g2_decap_8 FILLER_62_1697 ();
 sg13g2_decap_8 FILLER_62_1704 ();
 sg13g2_decap_8 FILLER_62_1711 ();
 sg13g2_decap_8 FILLER_62_1718 ();
 sg13g2_decap_8 FILLER_62_1725 ();
 sg13g2_decap_8 FILLER_62_1732 ();
 sg13g2_decap_8 FILLER_62_1739 ();
 sg13g2_decap_8 FILLER_62_1746 ();
 sg13g2_decap_8 FILLER_62_1753 ();
 sg13g2_decap_8 FILLER_62_1760 ();
 sg13g2_fill_1 FILLER_62_1767 ();
 sg13g2_fill_1 FILLER_63_26 ();
 sg13g2_fill_2 FILLER_63_56 ();
 sg13g2_fill_1 FILLER_63_58 ();
 sg13g2_fill_2 FILLER_63_105 ();
 sg13g2_fill_1 FILLER_63_141 ();
 sg13g2_fill_1 FILLER_63_173 ();
 sg13g2_fill_1 FILLER_63_178 ();
 sg13g2_fill_1 FILLER_63_196 ();
 sg13g2_fill_1 FILLER_63_202 ();
 sg13g2_fill_1 FILLER_63_228 ();
 sg13g2_fill_2 FILLER_63_350 ();
 sg13g2_decap_4 FILLER_63_417 ();
 sg13g2_fill_2 FILLER_63_421 ();
 sg13g2_fill_1 FILLER_63_431 ();
 sg13g2_fill_2 FILLER_63_486 ();
 sg13g2_fill_1 FILLER_63_488 ();
 sg13g2_fill_2 FILLER_63_515 ();
 sg13g2_fill_1 FILLER_63_553 ();
 sg13g2_fill_2 FILLER_63_605 ();
 sg13g2_fill_2 FILLER_63_619 ();
 sg13g2_fill_1 FILLER_63_621 ();
 sg13g2_fill_2 FILLER_63_631 ();
 sg13g2_fill_1 FILLER_63_633 ();
 sg13g2_fill_1 FILLER_63_646 ();
 sg13g2_fill_1 FILLER_63_673 ();
 sg13g2_fill_2 FILLER_63_705 ();
 sg13g2_fill_2 FILLER_63_735 ();
 sg13g2_fill_2 FILLER_63_740 ();
 sg13g2_fill_1 FILLER_63_742 ();
 sg13g2_fill_1 FILLER_63_748 ();
 sg13g2_fill_2 FILLER_63_754 ();
 sg13g2_fill_1 FILLER_63_756 ();
 sg13g2_decap_4 FILLER_63_776 ();
 sg13g2_fill_1 FILLER_63_780 ();
 sg13g2_decap_8 FILLER_63_801 ();
 sg13g2_fill_1 FILLER_63_808 ();
 sg13g2_decap_4 FILLER_63_846 ();
 sg13g2_fill_2 FILLER_63_855 ();
 sg13g2_fill_1 FILLER_63_857 ();
 sg13g2_decap_8 FILLER_63_877 ();
 sg13g2_decap_4 FILLER_63_884 ();
 sg13g2_fill_2 FILLER_63_888 ();
 sg13g2_fill_1 FILLER_63_905 ();
 sg13g2_decap_8 FILLER_63_911 ();
 sg13g2_fill_2 FILLER_63_938 ();
 sg13g2_decap_8 FILLER_63_959 ();
 sg13g2_decap_8 FILLER_63_966 ();
 sg13g2_fill_1 FILLER_63_973 ();
 sg13g2_fill_2 FILLER_63_989 ();
 sg13g2_fill_1 FILLER_63_991 ();
 sg13g2_decap_8 FILLER_63_1014 ();
 sg13g2_fill_2 FILLER_63_1021 ();
 sg13g2_fill_1 FILLER_63_1023 ();
 sg13g2_decap_4 FILLER_63_1032 ();
 sg13g2_fill_1 FILLER_63_1036 ();
 sg13g2_fill_2 FILLER_63_1041 ();
 sg13g2_fill_1 FILLER_63_1043 ();
 sg13g2_fill_2 FILLER_63_1060 ();
 sg13g2_decap_8 FILLER_63_1087 ();
 sg13g2_fill_2 FILLER_63_1102 ();
 sg13g2_fill_1 FILLER_63_1114 ();
 sg13g2_fill_1 FILLER_63_1190 ();
 sg13g2_fill_1 FILLER_63_1200 ();
 sg13g2_decap_4 FILLER_63_1222 ();
 sg13g2_fill_2 FILLER_63_1226 ();
 sg13g2_fill_1 FILLER_63_1262 ();
 sg13g2_fill_1 FILLER_63_1310 ();
 sg13g2_fill_1 FILLER_63_1363 ();
 sg13g2_fill_1 FILLER_63_1372 ();
 sg13g2_fill_1 FILLER_63_1467 ();
 sg13g2_decap_4 FILLER_63_1525 ();
 sg13g2_fill_2 FILLER_63_1543 ();
 sg13g2_fill_1 FILLER_63_1545 ();
 sg13g2_fill_2 FILLER_63_1597 ();
 sg13g2_fill_1 FILLER_63_1599 ();
 sg13g2_fill_2 FILLER_63_1622 ();
 sg13g2_decap_8 FILLER_63_1659 ();
 sg13g2_decap_8 FILLER_63_1666 ();
 sg13g2_decap_8 FILLER_63_1673 ();
 sg13g2_decap_8 FILLER_63_1680 ();
 sg13g2_decap_8 FILLER_63_1687 ();
 sg13g2_decap_8 FILLER_63_1694 ();
 sg13g2_decap_8 FILLER_63_1701 ();
 sg13g2_decap_8 FILLER_63_1708 ();
 sg13g2_decap_8 FILLER_63_1715 ();
 sg13g2_decap_8 FILLER_63_1722 ();
 sg13g2_decap_8 FILLER_63_1729 ();
 sg13g2_decap_8 FILLER_63_1736 ();
 sg13g2_decap_8 FILLER_63_1743 ();
 sg13g2_decap_8 FILLER_63_1750 ();
 sg13g2_decap_8 FILLER_63_1757 ();
 sg13g2_decap_4 FILLER_63_1764 ();
 sg13g2_fill_1 FILLER_64_42 ();
 sg13g2_fill_2 FILLER_64_92 ();
 sg13g2_fill_2 FILLER_64_155 ();
 sg13g2_fill_1 FILLER_64_157 ();
 sg13g2_fill_2 FILLER_64_166 ();
 sg13g2_fill_1 FILLER_64_168 ();
 sg13g2_fill_1 FILLER_64_173 ();
 sg13g2_fill_2 FILLER_64_179 ();
 sg13g2_fill_1 FILLER_64_201 ();
 sg13g2_fill_1 FILLER_64_254 ();
 sg13g2_fill_2 FILLER_64_356 ();
 sg13g2_fill_1 FILLER_64_441 ();
 sg13g2_fill_1 FILLER_64_453 ();
 sg13g2_fill_1 FILLER_64_469 ();
 sg13g2_decap_4 FILLER_64_482 ();
 sg13g2_fill_1 FILLER_64_486 ();
 sg13g2_fill_2 FILLER_64_497 ();
 sg13g2_decap_4 FILLER_64_506 ();
 sg13g2_fill_1 FILLER_64_510 ();
 sg13g2_fill_2 FILLER_64_613 ();
 sg13g2_fill_2 FILLER_64_641 ();
 sg13g2_fill_1 FILLER_64_658 ();
 sg13g2_fill_2 FILLER_64_664 ();
 sg13g2_fill_2 FILLER_64_708 ();
 sg13g2_fill_2 FILLER_64_729 ();
 sg13g2_fill_2 FILLER_64_762 ();
 sg13g2_fill_1 FILLER_64_764 ();
 sg13g2_fill_2 FILLER_64_769 ();
 sg13g2_decap_8 FILLER_64_801 ();
 sg13g2_fill_1 FILLER_64_808 ();
 sg13g2_decap_4 FILLER_64_842 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_fill_2 FILLER_64_871 ();
 sg13g2_fill_2 FILLER_64_935 ();
 sg13g2_fill_1 FILLER_64_946 ();
 sg13g2_decap_4 FILLER_64_961 ();
 sg13g2_fill_1 FILLER_64_965 ();
 sg13g2_fill_1 FILLER_64_989 ();
 sg13g2_fill_1 FILLER_64_1012 ();
 sg13g2_decap_4 FILLER_64_1016 ();
 sg13g2_fill_2 FILLER_64_1031 ();
 sg13g2_decap_8 FILLER_64_1043 ();
 sg13g2_decap_4 FILLER_64_1050 ();
 sg13g2_fill_1 FILLER_64_1069 ();
 sg13g2_decap_8 FILLER_64_1088 ();
 sg13g2_fill_1 FILLER_64_1095 ();
 sg13g2_fill_2 FILLER_64_1106 ();
 sg13g2_fill_1 FILLER_64_1108 ();
 sg13g2_fill_1 FILLER_64_1141 ();
 sg13g2_fill_2 FILLER_64_1161 ();
 sg13g2_fill_2 FILLER_64_1173 ();
 sg13g2_fill_1 FILLER_64_1175 ();
 sg13g2_fill_2 FILLER_64_1237 ();
 sg13g2_fill_1 FILLER_64_1239 ();
 sg13g2_fill_2 FILLER_64_1257 ();
 sg13g2_fill_1 FILLER_64_1259 ();
 sg13g2_fill_1 FILLER_64_1347 ();
 sg13g2_fill_1 FILLER_64_1369 ();
 sg13g2_fill_1 FILLER_64_1392 ();
 sg13g2_decap_4 FILLER_64_1428 ();
 sg13g2_fill_2 FILLER_64_1437 ();
 sg13g2_fill_2 FILLER_64_1448 ();
 sg13g2_fill_1 FILLER_64_1450 ();
 sg13g2_fill_2 FILLER_64_1455 ();
 sg13g2_fill_2 FILLER_64_1479 ();
 sg13g2_fill_2 FILLER_64_1495 ();
 sg13g2_fill_2 FILLER_64_1506 ();
 sg13g2_fill_1 FILLER_64_1508 ();
 sg13g2_fill_2 FILLER_64_1518 ();
 sg13g2_fill_1 FILLER_64_1520 ();
 sg13g2_fill_2 FILLER_64_1530 ();
 sg13g2_fill_1 FILLER_64_1532 ();
 sg13g2_fill_2 FILLER_64_1561 ();
 sg13g2_fill_2 FILLER_64_1577 ();
 sg13g2_fill_2 FILLER_64_1613 ();
 sg13g2_fill_1 FILLER_64_1615 ();
 sg13g2_fill_2 FILLER_64_1638 ();
 sg13g2_decap_8 FILLER_64_1661 ();
 sg13g2_decap_8 FILLER_64_1668 ();
 sg13g2_decap_8 FILLER_64_1675 ();
 sg13g2_decap_8 FILLER_64_1682 ();
 sg13g2_decap_8 FILLER_64_1689 ();
 sg13g2_decap_8 FILLER_64_1696 ();
 sg13g2_decap_8 FILLER_64_1703 ();
 sg13g2_decap_8 FILLER_64_1710 ();
 sg13g2_decap_8 FILLER_64_1717 ();
 sg13g2_decap_8 FILLER_64_1724 ();
 sg13g2_decap_8 FILLER_64_1731 ();
 sg13g2_decap_8 FILLER_64_1738 ();
 sg13g2_decap_8 FILLER_64_1745 ();
 sg13g2_decap_8 FILLER_64_1752 ();
 sg13g2_decap_8 FILLER_64_1759 ();
 sg13g2_fill_2 FILLER_64_1766 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_106 ();
 sg13g2_fill_1 FILLER_65_134 ();
 sg13g2_fill_2 FILLER_65_170 ();
 sg13g2_fill_1 FILLER_65_172 ();
 sg13g2_fill_2 FILLER_65_191 ();
 sg13g2_fill_1 FILLER_65_193 ();
 sg13g2_fill_2 FILLER_65_199 ();
 sg13g2_fill_1 FILLER_65_254 ();
 sg13g2_fill_2 FILLER_65_269 ();
 sg13g2_fill_1 FILLER_65_311 ();
 sg13g2_fill_1 FILLER_65_335 ();
 sg13g2_fill_1 FILLER_65_417 ();
 sg13g2_fill_2 FILLER_65_449 ();
 sg13g2_fill_1 FILLER_65_478 ();
 sg13g2_fill_2 FILLER_65_503 ();
 sg13g2_fill_1 FILLER_65_505 ();
 sg13g2_fill_2 FILLER_65_549 ();
 sg13g2_fill_1 FILLER_65_560 ();
 sg13g2_fill_2 FILLER_65_642 ();
 sg13g2_fill_2 FILLER_65_653 ();
 sg13g2_fill_1 FILLER_65_663 ();
 sg13g2_fill_2 FILLER_65_690 ();
 sg13g2_fill_2 FILLER_65_700 ();
 sg13g2_fill_2 FILLER_65_742 ();
 sg13g2_fill_2 FILLER_65_752 ();
 sg13g2_fill_2 FILLER_65_767 ();
 sg13g2_fill_1 FILLER_65_769 ();
 sg13g2_fill_2 FILLER_65_778 ();
 sg13g2_fill_1 FILLER_65_780 ();
 sg13g2_decap_4 FILLER_65_809 ();
 sg13g2_fill_2 FILLER_65_813 ();
 sg13g2_decap_4 FILLER_65_841 ();
 sg13g2_fill_1 FILLER_65_883 ();
 sg13g2_fill_2 FILLER_65_888 ();
 sg13g2_fill_2 FILLER_65_931 ();
 sg13g2_fill_1 FILLER_65_933 ();
 sg13g2_fill_2 FILLER_65_953 ();
 sg13g2_fill_1 FILLER_65_955 ();
 sg13g2_fill_1 FILLER_65_965 ();
 sg13g2_decap_8 FILLER_65_975 ();
 sg13g2_decap_8 FILLER_65_982 ();
 sg13g2_decap_8 FILLER_65_989 ();
 sg13g2_decap_4 FILLER_65_1001 ();
 sg13g2_fill_2 FILLER_65_1010 ();
 sg13g2_fill_2 FILLER_65_1038 ();
 sg13g2_decap_4 FILLER_65_1051 ();
 sg13g2_fill_2 FILLER_65_1075 ();
 sg13g2_fill_2 FILLER_65_1097 ();
 sg13g2_fill_2 FILLER_65_1118 ();
 sg13g2_fill_1 FILLER_65_1120 ();
 sg13g2_fill_2 FILLER_65_1147 ();
 sg13g2_decap_8 FILLER_65_1176 ();
 sg13g2_fill_2 FILLER_65_1183 ();
 sg13g2_fill_1 FILLER_65_1185 ();
 sg13g2_fill_2 FILLER_65_1230 ();
 sg13g2_fill_1 FILLER_65_1232 ();
 sg13g2_fill_1 FILLER_65_1250 ();
 sg13g2_fill_2 FILLER_65_1259 ();
 sg13g2_fill_1 FILLER_65_1261 ();
 sg13g2_fill_1 FILLER_65_1266 ();
 sg13g2_fill_1 FILLER_65_1272 ();
 sg13g2_decap_4 FILLER_65_1357 ();
 sg13g2_decap_4 FILLER_65_1366 ();
 sg13g2_fill_1 FILLER_65_1370 ();
 sg13g2_fill_1 FILLER_65_1385 ();
 sg13g2_decap_4 FILLER_65_1394 ();
 sg13g2_fill_1 FILLER_65_1398 ();
 sg13g2_fill_1 FILLER_65_1461 ();
 sg13g2_decap_4 FILLER_65_1477 ();
 sg13g2_fill_1 FILLER_65_1481 ();
 sg13g2_fill_1 FILLER_65_1508 ();
 sg13g2_fill_2 FILLER_65_1529 ();
 sg13g2_fill_1 FILLER_65_1546 ();
 sg13g2_fill_2 FILLER_65_1552 ();
 sg13g2_fill_1 FILLER_65_1594 ();
 sg13g2_decap_8 FILLER_65_1652 ();
 sg13g2_decap_8 FILLER_65_1659 ();
 sg13g2_decap_8 FILLER_65_1666 ();
 sg13g2_decap_8 FILLER_65_1673 ();
 sg13g2_decap_8 FILLER_65_1680 ();
 sg13g2_decap_8 FILLER_65_1687 ();
 sg13g2_decap_8 FILLER_65_1694 ();
 sg13g2_decap_8 FILLER_65_1701 ();
 sg13g2_decap_8 FILLER_65_1708 ();
 sg13g2_decap_8 FILLER_65_1715 ();
 sg13g2_decap_8 FILLER_65_1722 ();
 sg13g2_decap_8 FILLER_65_1729 ();
 sg13g2_decap_8 FILLER_65_1736 ();
 sg13g2_decap_8 FILLER_65_1743 ();
 sg13g2_decap_8 FILLER_65_1750 ();
 sg13g2_decap_8 FILLER_65_1757 ();
 sg13g2_decap_4 FILLER_65_1764 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_32 ();
 sg13g2_fill_2 FILLER_66_52 ();
 sg13g2_fill_1 FILLER_66_54 ();
 sg13g2_fill_2 FILLER_66_153 ();
 sg13g2_fill_1 FILLER_66_180 ();
 sg13g2_fill_2 FILLER_66_190 ();
 sg13g2_fill_2 FILLER_66_218 ();
 sg13g2_fill_1 FILLER_66_238 ();
 sg13g2_fill_2 FILLER_66_244 ();
 sg13g2_fill_2 FILLER_66_261 ();
 sg13g2_fill_1 FILLER_66_289 ();
 sg13g2_fill_1 FILLER_66_304 ();
 sg13g2_fill_1 FILLER_66_346 ();
 sg13g2_fill_2 FILLER_66_482 ();
 sg13g2_fill_1 FILLER_66_484 ();
 sg13g2_fill_2 FILLER_66_489 ();
 sg13g2_fill_2 FILLER_66_501 ();
 sg13g2_fill_1 FILLER_66_528 ();
 sg13g2_fill_1 FILLER_66_542 ();
 sg13g2_fill_2 FILLER_66_554 ();
 sg13g2_fill_1 FILLER_66_565 ();
 sg13g2_fill_1 FILLER_66_592 ();
 sg13g2_fill_2 FILLER_66_605 ();
 sg13g2_fill_2 FILLER_66_613 ();
 sg13g2_fill_2 FILLER_66_655 ();
 sg13g2_fill_1 FILLER_66_657 ();
 sg13g2_fill_2 FILLER_66_668 ();
 sg13g2_fill_1 FILLER_66_670 ();
 sg13g2_decap_8 FILLER_66_684 ();
 sg13g2_fill_1 FILLER_66_691 ();
 sg13g2_decap_8 FILLER_66_714 ();
 sg13g2_fill_1 FILLER_66_721 ();
 sg13g2_fill_1 FILLER_66_726 ();
 sg13g2_fill_1 FILLER_66_731 ();
 sg13g2_fill_2 FILLER_66_771 ();
 sg13g2_fill_1 FILLER_66_773 ();
 sg13g2_fill_2 FILLER_66_800 ();
 sg13g2_fill_2 FILLER_66_818 ();
 sg13g2_fill_1 FILLER_66_820 ();
 sg13g2_fill_1 FILLER_66_833 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_fill_1 FILLER_66_862 ();
 sg13g2_fill_1 FILLER_66_883 ();
 sg13g2_fill_1 FILLER_66_889 ();
 sg13g2_decap_4 FILLER_66_894 ();
 sg13g2_fill_2 FILLER_66_898 ();
 sg13g2_decap_4 FILLER_66_912 ();
 sg13g2_fill_2 FILLER_66_921 ();
 sg13g2_fill_1 FILLER_66_923 ();
 sg13g2_fill_1 FILLER_66_929 ();
 sg13g2_fill_2 FILLER_66_976 ();
 sg13g2_fill_1 FILLER_66_997 ();
 sg13g2_decap_8 FILLER_66_1003 ();
 sg13g2_fill_1 FILLER_66_1010 ();
 sg13g2_fill_1 FILLER_66_1026 ();
 sg13g2_fill_1 FILLER_66_1056 ();
 sg13g2_fill_2 FILLER_66_1065 ();
 sg13g2_fill_1 FILLER_66_1073 ();
 sg13g2_fill_1 FILLER_66_1179 ();
 sg13g2_fill_2 FILLER_66_1192 ();
 sg13g2_fill_1 FILLER_66_1213 ();
 sg13g2_fill_1 FILLER_66_1231 ();
 sg13g2_fill_2 FILLER_66_1269 ();
 sg13g2_fill_1 FILLER_66_1271 ();
 sg13g2_fill_1 FILLER_66_1305 ();
 sg13g2_fill_2 FILLER_66_1310 ();
 sg13g2_fill_1 FILLER_66_1406 ();
 sg13g2_fill_2 FILLER_66_1501 ();
 sg13g2_fill_1 FILLER_66_1503 ();
 sg13g2_fill_2 FILLER_66_1528 ();
 sg13g2_fill_1 FILLER_66_1530 ();
 sg13g2_fill_1 FILLER_66_1539 ();
 sg13g2_fill_2 FILLER_66_1554 ();
 sg13g2_fill_1 FILLER_66_1556 ();
 sg13g2_fill_2 FILLER_66_1597 ();
 sg13g2_fill_1 FILLER_66_1599 ();
 sg13g2_fill_2 FILLER_66_1635 ();
 sg13g2_decap_8 FILLER_66_1650 ();
 sg13g2_decap_8 FILLER_66_1657 ();
 sg13g2_decap_8 FILLER_66_1664 ();
 sg13g2_decap_8 FILLER_66_1671 ();
 sg13g2_decap_8 FILLER_66_1678 ();
 sg13g2_decap_8 FILLER_66_1685 ();
 sg13g2_decap_8 FILLER_66_1692 ();
 sg13g2_decap_8 FILLER_66_1699 ();
 sg13g2_decap_8 FILLER_66_1706 ();
 sg13g2_decap_8 FILLER_66_1713 ();
 sg13g2_decap_8 FILLER_66_1720 ();
 sg13g2_decap_8 FILLER_66_1727 ();
 sg13g2_decap_8 FILLER_66_1734 ();
 sg13g2_decap_8 FILLER_66_1741 ();
 sg13g2_decap_8 FILLER_66_1748 ();
 sg13g2_decap_8 FILLER_66_1755 ();
 sg13g2_decap_4 FILLER_66_1762 ();
 sg13g2_fill_2 FILLER_66_1766 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_31 ();
 sg13g2_fill_2 FILLER_67_58 ();
 sg13g2_fill_1 FILLER_67_60 ();
 sg13g2_fill_1 FILLER_67_74 ();
 sg13g2_fill_2 FILLER_67_89 ();
 sg13g2_fill_2 FILLER_67_104 ();
 sg13g2_fill_2 FILLER_67_125 ();
 sg13g2_fill_2 FILLER_67_136 ();
 sg13g2_fill_1 FILLER_67_138 ();
 sg13g2_fill_1 FILLER_67_184 ();
 sg13g2_fill_1 FILLER_67_221 ();
 sg13g2_fill_2 FILLER_67_242 ();
 sg13g2_fill_1 FILLER_67_244 ();
 sg13g2_fill_1 FILLER_67_257 ();
 sg13g2_fill_2 FILLER_67_268 ();
 sg13g2_fill_1 FILLER_67_270 ();
 sg13g2_fill_1 FILLER_67_394 ();
 sg13g2_fill_1 FILLER_67_417 ();
 sg13g2_fill_2 FILLER_67_428 ();
 sg13g2_fill_2 FILLER_67_472 ();
 sg13g2_fill_2 FILLER_67_554 ();
 sg13g2_fill_2 FILLER_67_603 ();
 sg13g2_fill_2 FILLER_67_631 ();
 sg13g2_fill_1 FILLER_67_638 ();
 sg13g2_fill_2 FILLER_67_665 ();
 sg13g2_fill_2 FILLER_67_675 ();
 sg13g2_fill_1 FILLER_67_677 ();
 sg13g2_fill_2 FILLER_67_684 ();
 sg13g2_decap_4 FILLER_67_693 ();
 sg13g2_fill_1 FILLER_67_710 ();
 sg13g2_fill_2 FILLER_67_739 ();
 sg13g2_fill_2 FILLER_67_746 ();
 sg13g2_fill_1 FILLER_67_748 ();
 sg13g2_fill_2 FILLER_67_754 ();
 sg13g2_fill_1 FILLER_67_761 ();
 sg13g2_fill_2 FILLER_67_770 ();
 sg13g2_fill_1 FILLER_67_772 ();
 sg13g2_decap_8 FILLER_67_790 ();
 sg13g2_fill_2 FILLER_67_797 ();
 sg13g2_fill_1 FILLER_67_804 ();
 sg13g2_fill_1 FILLER_67_818 ();
 sg13g2_decap_8 FILLER_67_833 ();
 sg13g2_decap_4 FILLER_67_840 ();
 sg13g2_fill_1 FILLER_67_844 ();
 sg13g2_fill_1 FILLER_67_849 ();
 sg13g2_fill_2 FILLER_67_872 ();
 sg13g2_fill_1 FILLER_67_874 ();
 sg13g2_fill_1 FILLER_67_907 ();
 sg13g2_decap_8 FILLER_67_916 ();
 sg13g2_decap_8 FILLER_67_923 ();
 sg13g2_fill_2 FILLER_67_930 ();
 sg13g2_fill_1 FILLER_67_932 ();
 sg13g2_fill_2 FILLER_67_954 ();
 sg13g2_fill_1 FILLER_67_956 ();
 sg13g2_decap_8 FILLER_67_983 ();
 sg13g2_fill_1 FILLER_67_990 ();
 sg13g2_decap_4 FILLER_67_1007 ();
 sg13g2_fill_2 FILLER_67_1019 ();
 sg13g2_fill_1 FILLER_67_1021 ();
 sg13g2_fill_2 FILLER_67_1033 ();
 sg13g2_fill_1 FILLER_67_1068 ();
 sg13g2_fill_1 FILLER_67_1094 ();
 sg13g2_fill_2 FILLER_67_1113 ();
 sg13g2_decap_8 FILLER_67_1143 ();
 sg13g2_fill_1 FILLER_67_1150 ();
 sg13g2_fill_2 FILLER_67_1201 ();
 sg13g2_fill_1 FILLER_67_1211 ();
 sg13g2_fill_1 FILLER_67_1226 ();
 sg13g2_fill_1 FILLER_67_1232 ();
 sg13g2_fill_1 FILLER_67_1246 ();
 sg13g2_fill_2 FILLER_67_1265 ();
 sg13g2_fill_2 FILLER_67_1279 ();
 sg13g2_fill_2 FILLER_67_1339 ();
 sg13g2_decap_4 FILLER_67_1373 ();
 sg13g2_fill_2 FILLER_67_1387 ();
 sg13g2_fill_2 FILLER_67_1449 ();
 sg13g2_fill_1 FILLER_67_1451 ();
 sg13g2_fill_2 FILLER_67_1468 ();
 sg13g2_fill_2 FILLER_67_1546 ();
 sg13g2_fill_1 FILLER_67_1548 ();
 sg13g2_fill_1 FILLER_67_1568 ();
 sg13g2_fill_2 FILLER_67_1578 ();
 sg13g2_fill_1 FILLER_67_1592 ();
 sg13g2_decap_8 FILLER_67_1650 ();
 sg13g2_decap_8 FILLER_67_1657 ();
 sg13g2_decap_8 FILLER_67_1664 ();
 sg13g2_decap_8 FILLER_67_1671 ();
 sg13g2_decap_8 FILLER_67_1678 ();
 sg13g2_decap_8 FILLER_67_1685 ();
 sg13g2_decap_8 FILLER_67_1692 ();
 sg13g2_decap_8 FILLER_67_1699 ();
 sg13g2_decap_8 FILLER_67_1706 ();
 sg13g2_decap_8 FILLER_67_1713 ();
 sg13g2_decap_8 FILLER_67_1720 ();
 sg13g2_decap_8 FILLER_67_1727 ();
 sg13g2_decap_8 FILLER_67_1734 ();
 sg13g2_decap_8 FILLER_67_1741 ();
 sg13g2_decap_8 FILLER_67_1748 ();
 sg13g2_decap_8 FILLER_67_1755 ();
 sg13g2_decap_4 FILLER_67_1762 ();
 sg13g2_fill_2 FILLER_67_1766 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_45 ();
 sg13g2_fill_1 FILLER_68_47 ();
 sg13g2_fill_1 FILLER_68_58 ();
 sg13g2_fill_2 FILLER_68_93 ();
 sg13g2_fill_1 FILLER_68_109 ();
 sg13g2_fill_2 FILLER_68_140 ();
 sg13g2_fill_2 FILLER_68_177 ();
 sg13g2_fill_1 FILLER_68_179 ();
 sg13g2_fill_2 FILLER_68_201 ();
 sg13g2_fill_2 FILLER_68_226 ();
 sg13g2_fill_1 FILLER_68_228 ();
 sg13g2_fill_2 FILLER_68_264 ();
 sg13g2_fill_1 FILLER_68_266 ();
 sg13g2_fill_1 FILLER_68_300 ();
 sg13g2_fill_1 FILLER_68_352 ();
 sg13g2_fill_1 FILLER_68_422 ();
 sg13g2_fill_2 FILLER_68_467 ();
 sg13g2_fill_2 FILLER_68_495 ();
 sg13g2_fill_1 FILLER_68_510 ();
 sg13g2_fill_2 FILLER_68_535 ();
 sg13g2_fill_1 FILLER_68_547 ();
 sg13g2_fill_2 FILLER_68_599 ();
 sg13g2_fill_2 FILLER_68_630 ();
 sg13g2_fill_2 FILLER_68_646 ();
 sg13g2_fill_1 FILLER_68_653 ();
 sg13g2_fill_1 FILLER_68_676 ();
 sg13g2_fill_2 FILLER_68_685 ();
 sg13g2_fill_1 FILLER_68_713 ();
 sg13g2_fill_1 FILLER_68_732 ();
 sg13g2_fill_1 FILLER_68_739 ();
 sg13g2_fill_2 FILLER_68_784 ();
 sg13g2_decap_4 FILLER_68_791 ();
 sg13g2_fill_1 FILLER_68_795 ();
 sg13g2_fill_2 FILLER_68_805 ();
 sg13g2_fill_1 FILLER_68_807 ();
 sg13g2_decap_4 FILLER_68_829 ();
 sg13g2_fill_1 FILLER_68_840 ();
 sg13g2_decap_4 FILLER_68_865 ();
 sg13g2_fill_1 FILLER_68_874 ();
 sg13g2_decap_8 FILLER_68_883 ();
 sg13g2_fill_2 FILLER_68_890 ();
 sg13g2_fill_1 FILLER_68_892 ();
 sg13g2_fill_2 FILLER_68_903 ();
 sg13g2_fill_2 FILLER_68_910 ();
 sg13g2_fill_1 FILLER_68_912 ();
 sg13g2_fill_1 FILLER_68_918 ();
 sg13g2_fill_1 FILLER_68_924 ();
 sg13g2_fill_1 FILLER_68_934 ();
 sg13g2_fill_2 FILLER_68_948 ();
 sg13g2_fill_1 FILLER_68_986 ();
 sg13g2_decap_8 FILLER_68_1006 ();
 sg13g2_fill_2 FILLER_68_1013 ();
 sg13g2_decap_4 FILLER_68_1036 ();
 sg13g2_decap_8 FILLER_68_1057 ();
 sg13g2_decap_4 FILLER_68_1064 ();
 sg13g2_fill_2 FILLER_68_1072 ();
 sg13g2_fill_2 FILLER_68_1079 ();
 sg13g2_decap_8 FILLER_68_1086 ();
 sg13g2_fill_1 FILLER_68_1102 ();
 sg13g2_fill_2 FILLER_68_1112 ();
 sg13g2_decap_4 FILLER_68_1137 ();
 sg13g2_fill_2 FILLER_68_1188 ();
 sg13g2_fill_2 FILLER_68_1322 ();
 sg13g2_fill_2 FILLER_68_1381 ();
 sg13g2_fill_2 FILLER_68_1430 ();
 sg13g2_fill_1 FILLER_68_1437 ();
 sg13g2_fill_2 FILLER_68_1447 ();
 sg13g2_fill_1 FILLER_68_1449 ();
 sg13g2_decap_8 FILLER_68_1459 ();
 sg13g2_decap_4 FILLER_68_1466 ();
 sg13g2_fill_1 FILLER_68_1470 ();
 sg13g2_fill_1 FILLER_68_1476 ();
 sg13g2_fill_2 FILLER_68_1496 ();
 sg13g2_fill_1 FILLER_68_1498 ();
 sg13g2_fill_2 FILLER_68_1505 ();
 sg13g2_fill_1 FILLER_68_1507 ();
 sg13g2_fill_2 FILLER_68_1539 ();
 sg13g2_fill_1 FILLER_68_1541 ();
 sg13g2_fill_2 FILLER_68_1594 ();
 sg13g2_decap_8 FILLER_68_1625 ();
 sg13g2_fill_1 FILLER_68_1632 ();
 sg13g2_decap_8 FILLER_68_1642 ();
 sg13g2_decap_8 FILLER_68_1649 ();
 sg13g2_decap_8 FILLER_68_1656 ();
 sg13g2_decap_8 FILLER_68_1663 ();
 sg13g2_decap_8 FILLER_68_1670 ();
 sg13g2_decap_8 FILLER_68_1677 ();
 sg13g2_decap_8 FILLER_68_1684 ();
 sg13g2_decap_8 FILLER_68_1691 ();
 sg13g2_decap_8 FILLER_68_1698 ();
 sg13g2_decap_8 FILLER_68_1705 ();
 sg13g2_decap_8 FILLER_68_1712 ();
 sg13g2_decap_8 FILLER_68_1719 ();
 sg13g2_decap_8 FILLER_68_1726 ();
 sg13g2_decap_8 FILLER_68_1733 ();
 sg13g2_decap_8 FILLER_68_1740 ();
 sg13g2_decap_8 FILLER_68_1747 ();
 sg13g2_decap_8 FILLER_68_1754 ();
 sg13g2_decap_8 FILLER_68_1761 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_68 ();
 sg13g2_fill_1 FILLER_69_70 ();
 sg13g2_fill_2 FILLER_69_80 ();
 sg13g2_fill_1 FILLER_69_82 ();
 sg13g2_fill_1 FILLER_69_122 ();
 sg13g2_fill_1 FILLER_69_132 ();
 sg13g2_fill_2 FILLER_69_185 ();
 sg13g2_fill_1 FILLER_69_187 ();
 sg13g2_fill_2 FILLER_69_211 ();
 sg13g2_fill_1 FILLER_69_213 ();
 sg13g2_fill_1 FILLER_69_227 ();
 sg13g2_fill_2 FILLER_69_237 ();
 sg13g2_fill_2 FILLER_69_268 ();
 sg13g2_fill_1 FILLER_69_270 ();
 sg13g2_fill_2 FILLER_69_364 ();
 sg13g2_fill_2 FILLER_69_516 ();
 sg13g2_fill_2 FILLER_69_562 ();
 sg13g2_fill_2 FILLER_69_656 ();
 sg13g2_decap_8 FILLER_69_664 ();
 sg13g2_fill_2 FILLER_69_671 ();
 sg13g2_fill_1 FILLER_69_673 ();
 sg13g2_fill_2 FILLER_69_683 ();
 sg13g2_fill_1 FILLER_69_685 ();
 sg13g2_fill_2 FILLER_69_690 ();
 sg13g2_fill_1 FILLER_69_692 ();
 sg13g2_decap_4 FILLER_69_706 ();
 sg13g2_fill_1 FILLER_69_710 ();
 sg13g2_decap_4 FILLER_69_716 ();
 sg13g2_fill_1 FILLER_69_720 ();
 sg13g2_decap_4 FILLER_69_738 ();
 sg13g2_fill_2 FILLER_69_742 ();
 sg13g2_fill_2 FILLER_69_749 ();
 sg13g2_fill_1 FILLER_69_751 ();
 sg13g2_decap_4 FILLER_69_757 ();
 sg13g2_fill_2 FILLER_69_785 ();
 sg13g2_decap_8 FILLER_69_792 ();
 sg13g2_fill_2 FILLER_69_799 ();
 sg13g2_fill_1 FILLER_69_801 ();
 sg13g2_fill_1 FILLER_69_824 ();
 sg13g2_decap_4 FILLER_69_830 ();
 sg13g2_fill_2 FILLER_69_834 ();
 sg13g2_decap_4 FILLER_69_841 ();
 sg13g2_fill_2 FILLER_69_875 ();
 sg13g2_fill_1 FILLER_69_924 ();
 sg13g2_decap_4 FILLER_69_950 ();
 sg13g2_fill_1 FILLER_69_954 ();
 sg13g2_fill_2 FILLER_69_976 ();
 sg13g2_decap_4 FILLER_69_997 ();
 sg13g2_fill_2 FILLER_69_1001 ();
 sg13g2_fill_2 FILLER_69_1020 ();
 sg13g2_fill_1 FILLER_69_1022 ();
 sg13g2_fill_2 FILLER_69_1028 ();
 sg13g2_fill_1 FILLER_69_1030 ();
 sg13g2_decap_4 FILLER_69_1036 ();
 sg13g2_fill_2 FILLER_69_1064 ();
 sg13g2_fill_1 FILLER_69_1066 ();
 sg13g2_fill_2 FILLER_69_1107 ();
 sg13g2_decap_4 FILLER_69_1148 ();
 sg13g2_fill_2 FILLER_69_1160 ();
 sg13g2_fill_2 FILLER_69_1327 ();
 sg13g2_fill_1 FILLER_69_1359 ();
 sg13g2_fill_2 FILLER_69_1383 ();
 sg13g2_fill_1 FILLER_69_1412 ();
 sg13g2_fill_2 FILLER_69_1418 ();
 sg13g2_fill_1 FILLER_69_1420 ();
 sg13g2_fill_2 FILLER_69_1431 ();
 sg13g2_fill_1 FILLER_69_1433 ();
 sg13g2_decap_4 FILLER_69_1460 ();
 sg13g2_fill_1 FILLER_69_1464 ();
 sg13g2_fill_2 FILLER_69_1478 ();
 sg13g2_fill_2 FILLER_69_1514 ();
 sg13g2_fill_1 FILLER_69_1516 ();
 sg13g2_fill_2 FILLER_69_1556 ();
 sg13g2_fill_1 FILLER_69_1562 ();
 sg13g2_fill_1 FILLER_69_1581 ();
 sg13g2_decap_8 FILLER_69_1621 ();
 sg13g2_decap_8 FILLER_69_1628 ();
 sg13g2_decap_8 FILLER_69_1635 ();
 sg13g2_decap_8 FILLER_69_1642 ();
 sg13g2_decap_8 FILLER_69_1649 ();
 sg13g2_decap_8 FILLER_69_1656 ();
 sg13g2_decap_8 FILLER_69_1663 ();
 sg13g2_decap_8 FILLER_69_1670 ();
 sg13g2_decap_8 FILLER_69_1677 ();
 sg13g2_decap_8 FILLER_69_1684 ();
 sg13g2_decap_8 FILLER_69_1691 ();
 sg13g2_decap_8 FILLER_69_1698 ();
 sg13g2_decap_8 FILLER_69_1705 ();
 sg13g2_decap_8 FILLER_69_1712 ();
 sg13g2_decap_8 FILLER_69_1719 ();
 sg13g2_decap_8 FILLER_69_1726 ();
 sg13g2_decap_8 FILLER_69_1733 ();
 sg13g2_decap_8 FILLER_69_1740 ();
 sg13g2_decap_8 FILLER_69_1747 ();
 sg13g2_decap_8 FILLER_69_1754 ();
 sg13g2_decap_8 FILLER_69_1761 ();
 sg13g2_fill_2 FILLER_70_35 ();
 sg13g2_fill_1 FILLER_70_37 ();
 sg13g2_fill_2 FILLER_70_83 ();
 sg13g2_fill_1 FILLER_70_85 ();
 sg13g2_fill_1 FILLER_70_100 ();
 sg13g2_fill_1 FILLER_70_148 ();
 sg13g2_fill_1 FILLER_70_158 ();
 sg13g2_fill_2 FILLER_70_194 ();
 sg13g2_fill_1 FILLER_70_211 ();
 sg13g2_fill_2 FILLER_70_319 ();
 sg13g2_fill_1 FILLER_70_352 ();
 sg13g2_fill_2 FILLER_70_362 ();
 sg13g2_fill_1 FILLER_70_441 ();
 sg13g2_fill_1 FILLER_70_459 ();
 sg13g2_fill_1 FILLER_70_584 ();
 sg13g2_fill_1 FILLER_70_588 ();
 sg13g2_decap_4 FILLER_70_599 ();
 sg13g2_fill_2 FILLER_70_612 ();
 sg13g2_fill_2 FILLER_70_623 ();
 sg13g2_fill_2 FILLER_70_646 ();
 sg13g2_decap_4 FILLER_70_671 ();
 sg13g2_fill_1 FILLER_70_675 ();
 sg13g2_fill_2 FILLER_70_694 ();
 sg13g2_fill_1 FILLER_70_706 ();
 sg13g2_fill_2 FILLER_70_743 ();
 sg13g2_fill_1 FILLER_70_745 ();
 sg13g2_fill_1 FILLER_70_751 ();
 sg13g2_fill_2 FILLER_70_760 ();
 sg13g2_fill_1 FILLER_70_762 ();
 sg13g2_fill_2 FILLER_70_774 ();
 sg13g2_fill_2 FILLER_70_788 ();
 sg13g2_decap_8 FILLER_70_802 ();
 sg13g2_decap_8 FILLER_70_809 ();
 sg13g2_fill_2 FILLER_70_833 ();
 sg13g2_fill_2 FILLER_70_873 ();
 sg13g2_decap_8 FILLER_70_885 ();
 sg13g2_decap_8 FILLER_70_892 ();
 sg13g2_decap_4 FILLER_70_904 ();
 sg13g2_fill_2 FILLER_70_908 ();
 sg13g2_decap_4 FILLER_70_915 ();
 sg13g2_decap_8 FILLER_70_949 ();
 sg13g2_fill_2 FILLER_70_956 ();
 sg13g2_fill_1 FILLER_70_958 ();
 sg13g2_fill_1 FILLER_70_972 ();
 sg13g2_fill_2 FILLER_70_1001 ();
 sg13g2_decap_8 FILLER_70_1013 ();
 sg13g2_decap_4 FILLER_70_1020 ();
 sg13g2_decap_4 FILLER_70_1042 ();
 sg13g2_fill_2 FILLER_70_1076 ();
 sg13g2_fill_2 FILLER_70_1090 ();
 sg13g2_fill_1 FILLER_70_1092 ();
 sg13g2_fill_2 FILLER_70_1106 ();
 sg13g2_fill_1 FILLER_70_1108 ();
 sg13g2_fill_2 FILLER_70_1116 ();
 sg13g2_decap_4 FILLER_70_1123 ();
 sg13g2_fill_1 FILLER_70_1127 ();
 sg13g2_decap_8 FILLER_70_1152 ();
 sg13g2_fill_2 FILLER_70_1176 ();
 sg13g2_fill_2 FILLER_70_1182 ();
 sg13g2_fill_1 FILLER_70_1184 ();
 sg13g2_fill_2 FILLER_70_1202 ();
 sg13g2_fill_2 FILLER_70_1260 ();
 sg13g2_fill_2 FILLER_70_1288 ();
 sg13g2_fill_1 FILLER_70_1290 ();
 sg13g2_fill_1 FILLER_70_1340 ();
 sg13g2_fill_2 FILLER_70_1394 ();
 sg13g2_fill_1 FILLER_70_1396 ();
 sg13g2_fill_2 FILLER_70_1416 ();
 sg13g2_fill_1 FILLER_70_1434 ();
 sg13g2_decap_8 FILLER_70_1452 ();
 sg13g2_decap_8 FILLER_70_1485 ();
 sg13g2_fill_2 FILLER_70_1560 ();
 sg13g2_fill_2 FILLER_70_1566 ();
 sg13g2_fill_1 FILLER_70_1568 ();
 sg13g2_decap_8 FILLER_70_1604 ();
 sg13g2_decap_8 FILLER_70_1611 ();
 sg13g2_decap_8 FILLER_70_1618 ();
 sg13g2_decap_8 FILLER_70_1625 ();
 sg13g2_decap_8 FILLER_70_1632 ();
 sg13g2_decap_8 FILLER_70_1639 ();
 sg13g2_decap_8 FILLER_70_1646 ();
 sg13g2_decap_8 FILLER_70_1653 ();
 sg13g2_decap_8 FILLER_70_1660 ();
 sg13g2_decap_8 FILLER_70_1667 ();
 sg13g2_decap_8 FILLER_70_1674 ();
 sg13g2_decap_8 FILLER_70_1681 ();
 sg13g2_decap_8 FILLER_70_1688 ();
 sg13g2_decap_8 FILLER_70_1695 ();
 sg13g2_decap_8 FILLER_70_1702 ();
 sg13g2_decap_8 FILLER_70_1709 ();
 sg13g2_decap_8 FILLER_70_1716 ();
 sg13g2_decap_8 FILLER_70_1723 ();
 sg13g2_decap_8 FILLER_70_1730 ();
 sg13g2_decap_8 FILLER_70_1737 ();
 sg13g2_decap_8 FILLER_70_1744 ();
 sg13g2_decap_8 FILLER_70_1751 ();
 sg13g2_decap_8 FILLER_70_1758 ();
 sg13g2_fill_2 FILLER_70_1765 ();
 sg13g2_fill_1 FILLER_70_1767 ();
 sg13g2_fill_2 FILLER_71_26 ();
 sg13g2_fill_1 FILLER_71_54 ();
 sg13g2_fill_2 FILLER_71_69 ();
 sg13g2_fill_1 FILLER_71_71 ();
 sg13g2_fill_1 FILLER_71_81 ();
 sg13g2_fill_1 FILLER_71_99 ();
 sg13g2_fill_2 FILLER_71_118 ();
 sg13g2_fill_1 FILLER_71_138 ();
 sg13g2_fill_2 FILLER_71_143 ();
 sg13g2_fill_1 FILLER_71_177 ();
 sg13g2_fill_2 FILLER_71_198 ();
 sg13g2_fill_1 FILLER_71_200 ();
 sg13g2_fill_2 FILLER_71_217 ();
 sg13g2_fill_2 FILLER_71_245 ();
 sg13g2_fill_1 FILLER_71_247 ();
 sg13g2_fill_1 FILLER_71_289 ();
 sg13g2_fill_2 FILLER_71_327 ();
 sg13g2_fill_1 FILLER_71_373 ();
 sg13g2_fill_2 FILLER_71_427 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_fill_2 FILLER_71_465 ();
 sg13g2_fill_1 FILLER_71_480 ();
 sg13g2_fill_1 FILLER_71_504 ();
 sg13g2_fill_1 FILLER_71_547 ();
 sg13g2_fill_1 FILLER_71_562 ();
 sg13g2_fill_1 FILLER_71_581 ();
 sg13g2_fill_1 FILLER_71_631 ();
 sg13g2_decap_8 FILLER_71_665 ();
 sg13g2_decap_8 FILLER_71_672 ();
 sg13g2_fill_1 FILLER_71_679 ();
 sg13g2_decap_4 FILLER_71_706 ();
 sg13g2_fill_1 FILLER_71_710 ();
 sg13g2_decap_8 FILLER_71_736 ();
 sg13g2_fill_2 FILLER_71_743 ();
 sg13g2_fill_2 FILLER_71_755 ();
 sg13g2_fill_2 FILLER_71_771 ();
 sg13g2_fill_1 FILLER_71_783 ();
 sg13g2_fill_1 FILLER_71_789 ();
 sg13g2_decap_8 FILLER_71_794 ();
 sg13g2_fill_1 FILLER_71_801 ();
 sg13g2_fill_2 FILLER_71_807 ();
 sg13g2_fill_1 FILLER_71_829 ();
 sg13g2_decap_8 FILLER_71_843 ();
 sg13g2_fill_2 FILLER_71_850 ();
 sg13g2_fill_1 FILLER_71_852 ();
 sg13g2_decap_4 FILLER_71_857 ();
 sg13g2_fill_2 FILLER_71_866 ();
 sg13g2_decap_4 FILLER_71_882 ();
 sg13g2_fill_1 FILLER_71_886 ();
 sg13g2_fill_2 FILLER_71_891 ();
 sg13g2_fill_2 FILLER_71_903 ();
 sg13g2_decap_8 FILLER_71_919 ();
 sg13g2_decap_4 FILLER_71_926 ();
 sg13g2_decap_4 FILLER_71_950 ();
 sg13g2_fill_2 FILLER_71_982 ();
 sg13g2_decap_4 FILLER_71_993 ();
 sg13g2_fill_1 FILLER_71_1019 ();
 sg13g2_fill_1 FILLER_71_1028 ();
 sg13g2_decap_8 FILLER_71_1045 ();
 sg13g2_fill_1 FILLER_71_1052 ();
 sg13g2_fill_2 FILLER_71_1063 ();
 sg13g2_fill_1 FILLER_71_1065 ();
 sg13g2_decap_4 FILLER_71_1071 ();
 sg13g2_fill_2 FILLER_71_1075 ();
 sg13g2_fill_2 FILLER_71_1091 ();
 sg13g2_fill_1 FILLER_71_1093 ();
 sg13g2_fill_2 FILLER_71_1103 ();
 sg13g2_fill_1 FILLER_71_1113 ();
 sg13g2_decap_4 FILLER_71_1120 ();
 sg13g2_fill_1 FILLER_71_1156 ();
 sg13g2_fill_2 FILLER_71_1165 ();
 sg13g2_fill_1 FILLER_71_1263 ();
 sg13g2_fill_2 FILLER_71_1278 ();
 sg13g2_fill_2 FILLER_71_1289 ();
 sg13g2_fill_1 FILLER_71_1291 ();
 sg13g2_fill_2 FILLER_71_1386 ();
 sg13g2_fill_1 FILLER_71_1415 ();
 sg13g2_decap_4 FILLER_71_1446 ();
 sg13g2_decap_4 FILLER_71_1520 ();
 sg13g2_fill_2 FILLER_71_1576 ();
 sg13g2_decap_8 FILLER_71_1591 ();
 sg13g2_decap_8 FILLER_71_1598 ();
 sg13g2_decap_8 FILLER_71_1605 ();
 sg13g2_decap_8 FILLER_71_1612 ();
 sg13g2_decap_8 FILLER_71_1619 ();
 sg13g2_decap_8 FILLER_71_1626 ();
 sg13g2_decap_8 FILLER_71_1633 ();
 sg13g2_decap_8 FILLER_71_1640 ();
 sg13g2_decap_8 FILLER_71_1647 ();
 sg13g2_decap_8 FILLER_71_1654 ();
 sg13g2_decap_8 FILLER_71_1661 ();
 sg13g2_decap_8 FILLER_71_1668 ();
 sg13g2_decap_8 FILLER_71_1675 ();
 sg13g2_decap_8 FILLER_71_1682 ();
 sg13g2_decap_8 FILLER_71_1689 ();
 sg13g2_decap_8 FILLER_71_1696 ();
 sg13g2_decap_8 FILLER_71_1703 ();
 sg13g2_decap_8 FILLER_71_1710 ();
 sg13g2_decap_8 FILLER_71_1717 ();
 sg13g2_decap_8 FILLER_71_1724 ();
 sg13g2_decap_8 FILLER_71_1731 ();
 sg13g2_decap_8 FILLER_71_1738 ();
 sg13g2_decap_8 FILLER_71_1745 ();
 sg13g2_decap_8 FILLER_71_1752 ();
 sg13g2_decap_8 FILLER_71_1759 ();
 sg13g2_fill_2 FILLER_71_1766 ();
 sg13g2_fill_1 FILLER_72_65 ();
 sg13g2_fill_2 FILLER_72_82 ();
 sg13g2_fill_2 FILLER_72_97 ();
 sg13g2_fill_1 FILLER_72_119 ();
 sg13g2_fill_2 FILLER_72_160 ();
 sg13g2_fill_1 FILLER_72_162 ();
 sg13g2_fill_1 FILLER_72_168 ();
 sg13g2_fill_2 FILLER_72_194 ();
 sg13g2_fill_1 FILLER_72_196 ();
 sg13g2_fill_1 FILLER_72_245 ();
 sg13g2_fill_2 FILLER_72_259 ();
 sg13g2_fill_1 FILLER_72_305 ();
 sg13g2_fill_2 FILLER_72_333 ();
 sg13g2_fill_2 FILLER_72_505 ();
 sg13g2_fill_1 FILLER_72_542 ();
 sg13g2_fill_2 FILLER_72_587 ();
 sg13g2_fill_1 FILLER_72_594 ();
 sg13g2_fill_1 FILLER_72_609 ();
 sg13g2_decap_4 FILLER_72_664 ();
 sg13g2_fill_1 FILLER_72_668 ();
 sg13g2_fill_1 FILLER_72_682 ();
 sg13g2_fill_2 FILLER_72_688 ();
 sg13g2_fill_1 FILLER_72_690 ();
 sg13g2_decap_4 FILLER_72_696 ();
 sg13g2_fill_1 FILLER_72_700 ();
 sg13g2_fill_1 FILLER_72_743 ();
 sg13g2_decap_8 FILLER_72_759 ();
 sg13g2_fill_1 FILLER_72_766 ();
 sg13g2_fill_2 FILLER_72_786 ();
 sg13g2_fill_1 FILLER_72_788 ();
 sg13g2_fill_2 FILLER_72_794 ();
 sg13g2_fill_1 FILLER_72_796 ();
 sg13g2_fill_1 FILLER_72_816 ();
 sg13g2_fill_2 FILLER_72_834 ();
 sg13g2_decap_4 FILLER_72_841 ();
 sg13g2_fill_1 FILLER_72_862 ();
 sg13g2_decap_4 FILLER_72_879 ();
 sg13g2_decap_8 FILLER_72_925 ();
 sg13g2_decap_4 FILLER_72_953 ();
 sg13g2_fill_1 FILLER_72_957 ();
 sg13g2_fill_1 FILLER_72_982 ();
 sg13g2_decap_8 FILLER_72_996 ();
 sg13g2_decap_8 FILLER_72_1020 ();
 sg13g2_decap_8 FILLER_72_1035 ();
 sg13g2_decap_4 FILLER_72_1055 ();
 sg13g2_fill_1 FILLER_72_1107 ();
 sg13g2_fill_2 FILLER_72_1127 ();
 sg13g2_fill_1 FILLER_72_1129 ();
 sg13g2_fill_2 FILLER_72_1151 ();
 sg13g2_fill_2 FILLER_72_1244 ();
 sg13g2_fill_1 FILLER_72_1246 ();
 sg13g2_fill_2 FILLER_72_1261 ();
 sg13g2_fill_1 FILLER_72_1263 ();
 sg13g2_fill_2 FILLER_72_1312 ();
 sg13g2_fill_1 FILLER_72_1314 ();
 sg13g2_fill_1 FILLER_72_1393 ();
 sg13g2_fill_2 FILLER_72_1421 ();
 sg13g2_fill_1 FILLER_72_1423 ();
 sg13g2_fill_1 FILLER_72_1429 ();
 sg13g2_fill_1 FILLER_72_1443 ();
 sg13g2_fill_2 FILLER_72_1467 ();
 sg13g2_fill_1 FILLER_72_1469 ();
 sg13g2_fill_2 FILLER_72_1485 ();
 sg13g2_fill_1 FILLER_72_1487 ();
 sg13g2_fill_2 FILLER_72_1518 ();
 sg13g2_decap_4 FILLER_72_1523 ();
 sg13g2_fill_1 FILLER_72_1527 ();
 sg13g2_fill_2 FILLER_72_1553 ();
 sg13g2_fill_1 FILLER_72_1555 ();
 sg13g2_fill_2 FILLER_72_1560 ();
 sg13g2_fill_1 FILLER_72_1562 ();
 sg13g2_fill_1 FILLER_72_1576 ();
 sg13g2_decap_8 FILLER_72_1581 ();
 sg13g2_decap_8 FILLER_72_1588 ();
 sg13g2_decap_8 FILLER_72_1595 ();
 sg13g2_decap_8 FILLER_72_1602 ();
 sg13g2_decap_8 FILLER_72_1609 ();
 sg13g2_decap_8 FILLER_72_1616 ();
 sg13g2_decap_8 FILLER_72_1623 ();
 sg13g2_decap_8 FILLER_72_1630 ();
 sg13g2_decap_8 FILLER_72_1637 ();
 sg13g2_decap_8 FILLER_72_1644 ();
 sg13g2_decap_8 FILLER_72_1651 ();
 sg13g2_decap_8 FILLER_72_1658 ();
 sg13g2_decap_8 FILLER_72_1665 ();
 sg13g2_decap_8 FILLER_72_1672 ();
 sg13g2_decap_8 FILLER_72_1679 ();
 sg13g2_decap_8 FILLER_72_1686 ();
 sg13g2_decap_8 FILLER_72_1693 ();
 sg13g2_decap_8 FILLER_72_1700 ();
 sg13g2_decap_8 FILLER_72_1707 ();
 sg13g2_decap_8 FILLER_72_1714 ();
 sg13g2_decap_8 FILLER_72_1721 ();
 sg13g2_decap_8 FILLER_72_1728 ();
 sg13g2_decap_8 FILLER_72_1735 ();
 sg13g2_decap_8 FILLER_72_1742 ();
 sg13g2_decap_8 FILLER_72_1749 ();
 sg13g2_decap_8 FILLER_72_1756 ();
 sg13g2_decap_4 FILLER_72_1763 ();
 sg13g2_fill_1 FILLER_72_1767 ();
 sg13g2_fill_2 FILLER_73_70 ();
 sg13g2_fill_2 FILLER_73_118 ();
 sg13g2_fill_2 FILLER_73_165 ();
 sg13g2_fill_1 FILLER_73_175 ();
 sg13g2_fill_2 FILLER_73_205 ();
 sg13g2_fill_1 FILLER_73_221 ();
 sg13g2_fill_2 FILLER_73_278 ();
 sg13g2_fill_1 FILLER_73_387 ();
 sg13g2_fill_2 FILLER_73_442 ();
 sg13g2_fill_2 FILLER_73_480 ();
 sg13g2_fill_1 FILLER_73_486 ();
 sg13g2_fill_1 FILLER_73_542 ();
 sg13g2_fill_1 FILLER_73_548 ();
 sg13g2_fill_1 FILLER_73_553 ();
 sg13g2_fill_1 FILLER_73_558 ();
 sg13g2_fill_1 FILLER_73_567 ();
 sg13g2_fill_1 FILLER_73_583 ();
 sg13g2_decap_4 FILLER_73_592 ();
 sg13g2_fill_2 FILLER_73_601 ();
 sg13g2_fill_2 FILLER_73_616 ();
 sg13g2_fill_2 FILLER_73_630 ();
 sg13g2_fill_1 FILLER_73_632 ();
 sg13g2_fill_2 FILLER_73_667 ();
 sg13g2_fill_1 FILLER_73_669 ();
 sg13g2_fill_2 FILLER_73_703 ();
 sg13g2_fill_2 FILLER_73_710 ();
 sg13g2_fill_1 FILLER_73_712 ();
 sg13g2_fill_2 FILLER_73_744 ();
 sg13g2_fill_1 FILLER_73_746 ();
 sg13g2_decap_4 FILLER_73_752 ();
 sg13g2_fill_2 FILLER_73_776 ();
 sg13g2_fill_1 FILLER_73_778 ();
 sg13g2_fill_2 FILLER_73_789 ();
 sg13g2_fill_1 FILLER_73_791 ();
 sg13g2_fill_2 FILLER_73_797 ();
 sg13g2_fill_1 FILLER_73_826 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_4 FILLER_73_843 ();
 sg13g2_fill_1 FILLER_73_855 ();
 sg13g2_fill_2 FILLER_73_864 ();
 sg13g2_fill_1 FILLER_73_866 ();
 sg13g2_fill_1 FILLER_73_872 ();
 sg13g2_decap_4 FILLER_73_878 ();
 sg13g2_fill_1 FILLER_73_882 ();
 sg13g2_decap_4 FILLER_73_888 ();
 sg13g2_decap_8 FILLER_73_902 ();
 sg13g2_decap_4 FILLER_73_909 ();
 sg13g2_fill_1 FILLER_73_913 ();
 sg13g2_decap_8 FILLER_73_919 ();
 sg13g2_fill_2 FILLER_73_926 ();
 sg13g2_fill_2 FILLER_73_934 ();
 sg13g2_fill_1 FILLER_73_941 ();
 sg13g2_decap_4 FILLER_73_956 ();
 sg13g2_fill_2 FILLER_73_973 ();
 sg13g2_fill_2 FILLER_73_983 ();
 sg13g2_fill_1 FILLER_73_985 ();
 sg13g2_decap_8 FILLER_73_1002 ();
 sg13g2_fill_1 FILLER_73_1009 ();
 sg13g2_fill_2 FILLER_73_1018 ();
 sg13g2_fill_1 FILLER_73_1025 ();
 sg13g2_decap_4 FILLER_73_1044 ();
 sg13g2_fill_2 FILLER_73_1048 ();
 sg13g2_fill_2 FILLER_73_1058 ();
 sg13g2_fill_1 FILLER_73_1060 ();
 sg13g2_fill_1 FILLER_73_1066 ();
 sg13g2_decap_8 FILLER_73_1096 ();
 sg13g2_fill_1 FILLER_73_1103 ();
 sg13g2_decap_4 FILLER_73_1109 ();
 sg13g2_fill_2 FILLER_73_1113 ();
 sg13g2_fill_2 FILLER_73_1123 ();
 sg13g2_fill_1 FILLER_73_1156 ();
 sg13g2_fill_1 FILLER_73_1171 ();
 sg13g2_fill_1 FILLER_73_1186 ();
 sg13g2_fill_2 FILLER_73_1222 ();
 sg13g2_fill_1 FILLER_73_1224 ();
 sg13g2_fill_2 FILLER_73_1272 ();
 sg13g2_fill_1 FILLER_73_1299 ();
 sg13g2_fill_1 FILLER_73_1344 ();
 sg13g2_fill_2 FILLER_73_1389 ();
 sg13g2_fill_2 FILLER_73_1447 ();
 sg13g2_fill_1 FILLER_73_1449 ();
 sg13g2_fill_2 FILLER_73_1499 ();
 sg13g2_decap_8 FILLER_73_1536 ();
 sg13g2_decap_8 FILLER_73_1543 ();
 sg13g2_decap_8 FILLER_73_1550 ();
 sg13g2_decap_8 FILLER_73_1557 ();
 sg13g2_decap_8 FILLER_73_1564 ();
 sg13g2_decap_8 FILLER_73_1571 ();
 sg13g2_decap_8 FILLER_73_1578 ();
 sg13g2_decap_8 FILLER_73_1585 ();
 sg13g2_decap_8 FILLER_73_1592 ();
 sg13g2_decap_8 FILLER_73_1599 ();
 sg13g2_decap_8 FILLER_73_1606 ();
 sg13g2_decap_8 FILLER_73_1613 ();
 sg13g2_decap_8 FILLER_73_1620 ();
 sg13g2_decap_8 FILLER_73_1627 ();
 sg13g2_decap_8 FILLER_73_1634 ();
 sg13g2_decap_8 FILLER_73_1641 ();
 sg13g2_decap_8 FILLER_73_1648 ();
 sg13g2_decap_8 FILLER_73_1655 ();
 sg13g2_decap_8 FILLER_73_1662 ();
 sg13g2_decap_8 FILLER_73_1669 ();
 sg13g2_decap_8 FILLER_73_1676 ();
 sg13g2_decap_8 FILLER_73_1683 ();
 sg13g2_decap_8 FILLER_73_1690 ();
 sg13g2_decap_8 FILLER_73_1697 ();
 sg13g2_decap_8 FILLER_73_1704 ();
 sg13g2_decap_8 FILLER_73_1711 ();
 sg13g2_decap_8 FILLER_73_1718 ();
 sg13g2_decap_8 FILLER_73_1725 ();
 sg13g2_decap_8 FILLER_73_1732 ();
 sg13g2_decap_8 FILLER_73_1739 ();
 sg13g2_decap_8 FILLER_73_1746 ();
 sg13g2_decap_8 FILLER_73_1753 ();
 sg13g2_decap_8 FILLER_73_1760 ();
 sg13g2_fill_1 FILLER_73_1767 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_2 ();
 sg13g2_fill_1 FILLER_74_28 ();
 sg13g2_fill_1 FILLER_74_34 ();
 sg13g2_fill_2 FILLER_74_40 ();
 sg13g2_fill_1 FILLER_74_42 ();
 sg13g2_fill_2 FILLER_74_57 ();
 sg13g2_fill_1 FILLER_74_59 ();
 sg13g2_fill_2 FILLER_74_69 ();
 sg13g2_fill_1 FILLER_74_71 ();
 sg13g2_fill_1 FILLER_74_80 ();
 sg13g2_fill_1 FILLER_74_95 ();
 sg13g2_decap_4 FILLER_74_167 ();
 sg13g2_fill_1 FILLER_74_193 ();
 sg13g2_fill_2 FILLER_74_203 ();
 sg13g2_fill_1 FILLER_74_211 ();
 sg13g2_fill_1 FILLER_74_235 ();
 sg13g2_fill_1 FILLER_74_266 ();
 sg13g2_fill_1 FILLER_74_301 ();
 sg13g2_fill_1 FILLER_74_308 ();
 sg13g2_fill_2 FILLER_74_329 ();
 sg13g2_fill_2 FILLER_74_349 ();
 sg13g2_fill_2 FILLER_74_477 ();
 sg13g2_fill_1 FILLER_74_503 ();
 sg13g2_fill_1 FILLER_74_532 ();
 sg13g2_fill_1 FILLER_74_553 ();
 sg13g2_decap_4 FILLER_74_591 ();
 sg13g2_decap_4 FILLER_74_639 ();
 sg13g2_fill_1 FILLER_74_643 ();
 sg13g2_fill_2 FILLER_74_663 ();
 sg13g2_fill_2 FILLER_74_690 ();
 sg13g2_fill_1 FILLER_74_692 ();
 sg13g2_fill_1 FILLER_74_745 ();
 sg13g2_decap_4 FILLER_74_751 ();
 sg13g2_fill_1 FILLER_74_759 ();
 sg13g2_decap_4 FILLER_74_781 ();
 sg13g2_fill_2 FILLER_74_785 ();
 sg13g2_fill_2 FILLER_74_810 ();
 sg13g2_fill_2 FILLER_74_820 ();
 sg13g2_fill_1 FILLER_74_822 ();
 sg13g2_decap_4 FILLER_74_832 ();
 sg13g2_fill_1 FILLER_74_836 ();
 sg13g2_fill_2 FILLER_74_859 ();
 sg13g2_fill_1 FILLER_74_866 ();
 sg13g2_decap_8 FILLER_74_911 ();
 sg13g2_decap_4 FILLER_74_933 ();
 sg13g2_fill_1 FILLER_74_956 ();
 sg13g2_fill_2 FILLER_74_988 ();
 sg13g2_fill_2 FILLER_74_1006 ();
 sg13g2_fill_2 FILLER_74_1037 ();
 sg13g2_fill_1 FILLER_74_1039 ();
 sg13g2_decap_8 FILLER_74_1055 ();
 sg13g2_decap_4 FILLER_74_1062 ();
 sg13g2_decap_8 FILLER_74_1084 ();
 sg13g2_fill_1 FILLER_74_1112 ();
 sg13g2_fill_2 FILLER_74_1148 ();
 sg13g2_fill_2 FILLER_74_1186 ();
 sg13g2_fill_1 FILLER_74_1188 ();
 sg13g2_fill_2 FILLER_74_1291 ();
 sg13g2_fill_2 FILLER_74_1328 ();
 sg13g2_fill_2 FILLER_74_1361 ();
 sg13g2_fill_1 FILLER_74_1389 ();
 sg13g2_fill_2 FILLER_74_1466 ();
 sg13g2_fill_1 FILLER_74_1468 ();
 sg13g2_fill_2 FILLER_74_1479 ();
 sg13g2_fill_1 FILLER_74_1511 ();
 sg13g2_decap_8 FILLER_74_1516 ();
 sg13g2_decap_8 FILLER_74_1523 ();
 sg13g2_decap_8 FILLER_74_1530 ();
 sg13g2_decap_8 FILLER_74_1537 ();
 sg13g2_decap_8 FILLER_74_1544 ();
 sg13g2_decap_8 FILLER_74_1551 ();
 sg13g2_decap_8 FILLER_74_1558 ();
 sg13g2_decap_8 FILLER_74_1565 ();
 sg13g2_decap_8 FILLER_74_1572 ();
 sg13g2_decap_8 FILLER_74_1579 ();
 sg13g2_decap_8 FILLER_74_1586 ();
 sg13g2_decap_8 FILLER_74_1593 ();
 sg13g2_decap_8 FILLER_74_1600 ();
 sg13g2_decap_8 FILLER_74_1607 ();
 sg13g2_decap_8 FILLER_74_1614 ();
 sg13g2_decap_8 FILLER_74_1621 ();
 sg13g2_decap_8 FILLER_74_1628 ();
 sg13g2_decap_8 FILLER_74_1635 ();
 sg13g2_decap_8 FILLER_74_1642 ();
 sg13g2_decap_8 FILLER_74_1649 ();
 sg13g2_decap_8 FILLER_74_1656 ();
 sg13g2_decap_8 FILLER_74_1663 ();
 sg13g2_decap_8 FILLER_74_1670 ();
 sg13g2_decap_8 FILLER_74_1677 ();
 sg13g2_decap_8 FILLER_74_1684 ();
 sg13g2_decap_8 FILLER_74_1691 ();
 sg13g2_decap_8 FILLER_74_1698 ();
 sg13g2_decap_8 FILLER_74_1705 ();
 sg13g2_decap_8 FILLER_74_1712 ();
 sg13g2_decap_8 FILLER_74_1719 ();
 sg13g2_decap_8 FILLER_74_1726 ();
 sg13g2_decap_8 FILLER_74_1733 ();
 sg13g2_decap_8 FILLER_74_1740 ();
 sg13g2_decap_8 FILLER_74_1747 ();
 sg13g2_decap_8 FILLER_74_1754 ();
 sg13g2_decap_8 FILLER_74_1761 ();
 sg13g2_fill_1 FILLER_75_32 ();
 sg13g2_fill_1 FILLER_75_65 ();
 sg13g2_fill_2 FILLER_75_74 ();
 sg13g2_fill_1 FILLER_75_88 ();
 sg13g2_fill_2 FILLER_75_138 ();
 sg13g2_fill_1 FILLER_75_146 ();
 sg13g2_fill_1 FILLER_75_154 ();
 sg13g2_fill_1 FILLER_75_164 ();
 sg13g2_decap_4 FILLER_75_171 ();
 sg13g2_fill_1 FILLER_75_175 ();
 sg13g2_fill_1 FILLER_75_194 ();
 sg13g2_fill_1 FILLER_75_200 ();
 sg13g2_fill_1 FILLER_75_217 ();
 sg13g2_fill_2 FILLER_75_279 ();
 sg13g2_fill_1 FILLER_75_362 ();
 sg13g2_fill_1 FILLER_75_403 ();
 sg13g2_fill_2 FILLER_75_417 ();
 sg13g2_fill_1 FILLER_75_419 ();
 sg13g2_fill_2 FILLER_75_455 ();
 sg13g2_fill_1 FILLER_75_487 ();
 sg13g2_fill_2 FILLER_75_528 ();
 sg13g2_fill_2 FILLER_75_538 ();
 sg13g2_fill_1 FILLER_75_597 ();
 sg13g2_fill_1 FILLER_75_624 ();
 sg13g2_decap_8 FILLER_75_664 ();
 sg13g2_fill_2 FILLER_75_671 ();
 sg13g2_fill_1 FILLER_75_673 ();
 sg13g2_fill_2 FILLER_75_679 ();
 sg13g2_decap_4 FILLER_75_691 ();
 sg13g2_fill_1 FILLER_75_710 ();
 sg13g2_decap_8 FILLER_75_727 ();
 sg13g2_fill_1 FILLER_75_734 ();
 sg13g2_decap_4 FILLER_75_739 ();
 sg13g2_fill_1 FILLER_75_748 ();
 sg13g2_decap_4 FILLER_75_770 ();
 sg13g2_fill_2 FILLER_75_787 ();
 sg13g2_fill_1 FILLER_75_789 ();
 sg13g2_fill_2 FILLER_75_805 ();
 sg13g2_fill_1 FILLER_75_812 ();
 sg13g2_fill_2 FILLER_75_827 ();
 sg13g2_fill_2 FILLER_75_842 ();
 sg13g2_fill_2 FILLER_75_849 ();
 sg13g2_fill_2 FILLER_75_860 ();
 sg13g2_fill_1 FILLER_75_862 ();
 sg13g2_fill_2 FILLER_75_878 ();
 sg13g2_fill_1 FILLER_75_880 ();
 sg13g2_decap_8 FILLER_75_896 ();
 sg13g2_decap_8 FILLER_75_908 ();
 sg13g2_decap_8 FILLER_75_930 ();
 sg13g2_fill_2 FILLER_75_937 ();
 sg13g2_fill_1 FILLER_75_939 ();
 sg13g2_fill_2 FILLER_75_959 ();
 sg13g2_fill_1 FILLER_75_961 ();
 sg13g2_fill_2 FILLER_75_966 ();
 sg13g2_fill_1 FILLER_75_968 ();
 sg13g2_fill_1 FILLER_75_1003 ();
 sg13g2_fill_2 FILLER_75_1008 ();
 sg13g2_decap_4 FILLER_75_1029 ();
 sg13g2_fill_2 FILLER_75_1033 ();
 sg13g2_fill_1 FILLER_75_1040 ();
 sg13g2_decap_8 FILLER_75_1051 ();
 sg13g2_decap_8 FILLER_75_1058 ();
 sg13g2_decap_4 FILLER_75_1065 ();
 sg13g2_fill_2 FILLER_75_1247 ();
 sg13g2_fill_1 FILLER_75_1257 ();
 sg13g2_fill_2 FILLER_75_1325 ();
 sg13g2_fill_2 FILLER_75_1353 ();
 sg13g2_fill_1 FILLER_75_1355 ();
 sg13g2_fill_2 FILLER_75_1382 ();
 sg13g2_fill_1 FILLER_75_1384 ();
 sg13g2_fill_2 FILLER_75_1398 ();
 sg13g2_decap_8 FILLER_75_1501 ();
 sg13g2_decap_8 FILLER_75_1508 ();
 sg13g2_decap_8 FILLER_75_1515 ();
 sg13g2_decap_8 FILLER_75_1522 ();
 sg13g2_decap_8 FILLER_75_1529 ();
 sg13g2_decap_8 FILLER_75_1536 ();
 sg13g2_decap_8 FILLER_75_1543 ();
 sg13g2_decap_8 FILLER_75_1550 ();
 sg13g2_decap_8 FILLER_75_1557 ();
 sg13g2_decap_8 FILLER_75_1564 ();
 sg13g2_decap_8 FILLER_75_1571 ();
 sg13g2_decap_8 FILLER_75_1578 ();
 sg13g2_decap_8 FILLER_75_1585 ();
 sg13g2_decap_8 FILLER_75_1592 ();
 sg13g2_decap_8 FILLER_75_1599 ();
 sg13g2_decap_8 FILLER_75_1606 ();
 sg13g2_decap_8 FILLER_75_1613 ();
 sg13g2_decap_8 FILLER_75_1620 ();
 sg13g2_decap_8 FILLER_75_1627 ();
 sg13g2_decap_8 FILLER_75_1634 ();
 sg13g2_decap_8 FILLER_75_1641 ();
 sg13g2_decap_8 FILLER_75_1648 ();
 sg13g2_decap_8 FILLER_75_1655 ();
 sg13g2_decap_8 FILLER_75_1662 ();
 sg13g2_decap_8 FILLER_75_1669 ();
 sg13g2_decap_8 FILLER_75_1676 ();
 sg13g2_decap_8 FILLER_75_1683 ();
 sg13g2_decap_8 FILLER_75_1690 ();
 sg13g2_decap_8 FILLER_75_1697 ();
 sg13g2_decap_8 FILLER_75_1704 ();
 sg13g2_decap_8 FILLER_75_1711 ();
 sg13g2_decap_8 FILLER_75_1718 ();
 sg13g2_decap_8 FILLER_75_1725 ();
 sg13g2_decap_8 FILLER_75_1732 ();
 sg13g2_decap_8 FILLER_75_1739 ();
 sg13g2_decap_8 FILLER_75_1746 ();
 sg13g2_decap_8 FILLER_75_1753 ();
 sg13g2_decap_8 FILLER_75_1760 ();
 sg13g2_fill_1 FILLER_75_1767 ();
 sg13g2_fill_2 FILLER_76_30 ();
 sg13g2_fill_2 FILLER_76_63 ();
 sg13g2_fill_2 FILLER_76_96 ();
 sg13g2_fill_1 FILLER_76_98 ();
 sg13g2_fill_2 FILLER_76_122 ();
 sg13g2_fill_2 FILLER_76_140 ();
 sg13g2_fill_1 FILLER_76_142 ();
 sg13g2_fill_2 FILLER_76_148 ();
 sg13g2_fill_1 FILLER_76_150 ();
 sg13g2_fill_1 FILLER_76_173 ();
 sg13g2_fill_1 FILLER_76_196 ();
 sg13g2_fill_1 FILLER_76_211 ();
 sg13g2_fill_2 FILLER_76_230 ();
 sg13g2_fill_1 FILLER_76_273 ();
 sg13g2_fill_1 FILLER_76_283 ();
 sg13g2_fill_1 FILLER_76_293 ();
 sg13g2_decap_4 FILLER_76_308 ();
 sg13g2_fill_2 FILLER_76_348 ();
 sg13g2_fill_2 FILLER_76_380 ();
 sg13g2_fill_2 FILLER_76_482 ();
 sg13g2_fill_1 FILLER_76_532 ();
 sg13g2_fill_1 FILLER_76_538 ();
 sg13g2_fill_1 FILLER_76_554 ();
 sg13g2_fill_2 FILLER_76_560 ();
 sg13g2_fill_2 FILLER_76_567 ();
 sg13g2_fill_1 FILLER_76_584 ();
 sg13g2_decap_4 FILLER_76_638 ();
 sg13g2_fill_2 FILLER_76_653 ();
 sg13g2_fill_1 FILLER_76_655 ();
 sg13g2_fill_2 FILLER_76_667 ();
 sg13g2_fill_1 FILLER_76_669 ();
 sg13g2_fill_2 FILLER_76_701 ();
 sg13g2_fill_2 FILLER_76_728 ();
 sg13g2_fill_2 FILLER_76_749 ();
 sg13g2_fill_2 FILLER_76_756 ();
 sg13g2_fill_1 FILLER_76_764 ();
 sg13g2_fill_2 FILLER_76_780 ();
 sg13g2_fill_1 FILLER_76_782 ();
 sg13g2_fill_1 FILLER_76_792 ();
 sg13g2_fill_2 FILLER_76_798 ();
 sg13g2_fill_1 FILLER_76_800 ();
 sg13g2_fill_1 FILLER_76_832 ();
 sg13g2_decap_4 FILLER_76_877 ();
 sg13g2_fill_1 FILLER_76_881 ();
 sg13g2_fill_1 FILLER_76_892 ();
 sg13g2_decap_4 FILLER_76_898 ();
 sg13g2_fill_1 FILLER_76_902 ();
 sg13g2_fill_1 FILLER_76_907 ();
 sg13g2_fill_2 FILLER_76_921 ();
 sg13g2_decap_4 FILLER_76_928 ();
 sg13g2_fill_1 FILLER_76_932 ();
 sg13g2_fill_2 FILLER_76_953 ();
 sg13g2_fill_1 FILLER_76_981 ();
 sg13g2_fill_2 FILLER_76_1021 ();
 sg13g2_fill_1 FILLER_76_1023 ();
 sg13g2_fill_1 FILLER_76_1031 ();
 sg13g2_fill_2 FILLER_76_1056 ();
 sg13g2_fill_2 FILLER_76_1070 ();
 sg13g2_fill_1 FILLER_76_1072 ();
 sg13g2_fill_2 FILLER_76_1113 ();
 sg13g2_fill_1 FILLER_76_1133 ();
 sg13g2_fill_2 FILLER_76_1197 ();
 sg13g2_fill_1 FILLER_76_1199 ();
 sg13g2_fill_2 FILLER_76_1223 ();
 sg13g2_fill_1 FILLER_76_1225 ();
 sg13g2_fill_1 FILLER_76_1259 ();
 sg13g2_fill_1 FILLER_76_1278 ();
 sg13g2_fill_1 FILLER_76_1334 ();
 sg13g2_fill_1 FILLER_76_1361 ();
 sg13g2_fill_1 FILLER_76_1422 ();
 sg13g2_fill_2 FILLER_76_1432 ();
 sg13g2_fill_1 FILLER_76_1461 ();
 sg13g2_decap_8 FILLER_76_1485 ();
 sg13g2_decap_8 FILLER_76_1492 ();
 sg13g2_decap_8 FILLER_76_1499 ();
 sg13g2_decap_8 FILLER_76_1506 ();
 sg13g2_decap_8 FILLER_76_1513 ();
 sg13g2_decap_8 FILLER_76_1520 ();
 sg13g2_decap_8 FILLER_76_1527 ();
 sg13g2_decap_8 FILLER_76_1534 ();
 sg13g2_decap_8 FILLER_76_1541 ();
 sg13g2_decap_8 FILLER_76_1548 ();
 sg13g2_decap_8 FILLER_76_1555 ();
 sg13g2_decap_8 FILLER_76_1562 ();
 sg13g2_decap_8 FILLER_76_1569 ();
 sg13g2_decap_8 FILLER_76_1576 ();
 sg13g2_decap_8 FILLER_76_1583 ();
 sg13g2_decap_8 FILLER_76_1590 ();
 sg13g2_decap_8 FILLER_76_1597 ();
 sg13g2_decap_8 FILLER_76_1604 ();
 sg13g2_decap_8 FILLER_76_1611 ();
 sg13g2_decap_8 FILLER_76_1618 ();
 sg13g2_decap_8 FILLER_76_1625 ();
 sg13g2_decap_8 FILLER_76_1632 ();
 sg13g2_decap_8 FILLER_76_1639 ();
 sg13g2_decap_8 FILLER_76_1646 ();
 sg13g2_decap_8 FILLER_76_1653 ();
 sg13g2_decap_8 FILLER_76_1660 ();
 sg13g2_decap_8 FILLER_76_1667 ();
 sg13g2_decap_8 FILLER_76_1674 ();
 sg13g2_decap_8 FILLER_76_1681 ();
 sg13g2_decap_8 FILLER_76_1688 ();
 sg13g2_decap_8 FILLER_76_1695 ();
 sg13g2_decap_8 FILLER_76_1702 ();
 sg13g2_decap_8 FILLER_76_1709 ();
 sg13g2_decap_8 FILLER_76_1716 ();
 sg13g2_decap_8 FILLER_76_1723 ();
 sg13g2_decap_8 FILLER_76_1730 ();
 sg13g2_decap_8 FILLER_76_1737 ();
 sg13g2_decap_8 FILLER_76_1744 ();
 sg13g2_decap_8 FILLER_76_1751 ();
 sg13g2_decap_8 FILLER_76_1758 ();
 sg13g2_fill_2 FILLER_76_1765 ();
 sg13g2_fill_1 FILLER_76_1767 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_27 ();
 sg13g2_fill_2 FILLER_77_43 ();
 sg13g2_fill_1 FILLER_77_45 ();
 sg13g2_fill_2 FILLER_77_54 ();
 sg13g2_fill_1 FILLER_77_64 ();
 sg13g2_fill_2 FILLER_77_97 ();
 sg13g2_fill_2 FILLER_77_106 ();
 sg13g2_fill_1 FILLER_77_108 ();
 sg13g2_fill_2 FILLER_77_125 ();
 sg13g2_fill_1 FILLER_77_127 ();
 sg13g2_fill_2 FILLER_77_156 ();
 sg13g2_fill_1 FILLER_77_158 ();
 sg13g2_fill_1 FILLER_77_165 ();
 sg13g2_fill_1 FILLER_77_169 ();
 sg13g2_fill_1 FILLER_77_175 ();
 sg13g2_fill_1 FILLER_77_189 ();
 sg13g2_fill_1 FILLER_77_213 ();
 sg13g2_fill_2 FILLER_77_240 ();
 sg13g2_fill_2 FILLER_77_332 ();
 sg13g2_fill_2 FILLER_77_399 ();
 sg13g2_fill_2 FILLER_77_468 ();
 sg13g2_fill_1 FILLER_77_489 ();
 sg13g2_fill_2 FILLER_77_516 ();
 sg13g2_fill_2 FILLER_77_553 ();
 sg13g2_fill_2 FILLER_77_564 ();
 sg13g2_decap_8 FILLER_77_663 ();
 sg13g2_decap_4 FILLER_77_675 ();
 sg13g2_decap_4 FILLER_77_702 ();
 sg13g2_fill_2 FILLER_77_706 ();
 sg13g2_fill_1 FILLER_77_712 ();
 sg13g2_fill_1 FILLER_77_728 ();
 sg13g2_decap_4 FILLER_77_734 ();
 sg13g2_fill_2 FILLER_77_738 ();
 sg13g2_fill_2 FILLER_77_757 ();
 sg13g2_fill_1 FILLER_77_759 ();
 sg13g2_fill_1 FILLER_77_770 ();
 sg13g2_fill_1 FILLER_77_781 ();
 sg13g2_fill_2 FILLER_77_805 ();
 sg13g2_decap_4 FILLER_77_840 ();
 sg13g2_fill_1 FILLER_77_844 ();
 sg13g2_fill_1 FILLER_77_859 ();
 sg13g2_decap_4 FILLER_77_864 ();
 sg13g2_fill_1 FILLER_77_868 ();
 sg13g2_fill_2 FILLER_77_874 ();
 sg13g2_fill_2 FILLER_77_886 ();
 sg13g2_decap_4 FILLER_77_961 ();
 sg13g2_fill_1 FILLER_77_965 ();
 sg13g2_decap_8 FILLER_77_975 ();
 sg13g2_decap_8 FILLER_77_982 ();
 sg13g2_fill_1 FILLER_77_994 ();
 sg13g2_fill_2 FILLER_77_1008 ();
 sg13g2_decap_8 FILLER_77_1015 ();
 sg13g2_fill_1 FILLER_77_1022 ();
 sg13g2_decap_8 FILLER_77_1050 ();
 sg13g2_fill_2 FILLER_77_1085 ();
 sg13g2_fill_1 FILLER_77_1087 ();
 sg13g2_fill_2 FILLER_77_1131 ();
 sg13g2_fill_1 FILLER_77_1142 ();
 sg13g2_fill_1 FILLER_77_1175 ();
 sg13g2_fill_1 FILLER_77_1197 ();
 sg13g2_fill_1 FILLER_77_1250 ();
 sg13g2_fill_1 FILLER_77_1278 ();
 sg13g2_decap_8 FILLER_77_1358 ();
 sg13g2_decap_4 FILLER_77_1365 ();
 sg13g2_fill_2 FILLER_77_1388 ();
 sg13g2_fill_1 FILLER_77_1399 ();
 sg13g2_fill_1 FILLER_77_1409 ();
 sg13g2_decap_8 FILLER_77_1493 ();
 sg13g2_decap_8 FILLER_77_1500 ();
 sg13g2_decap_8 FILLER_77_1507 ();
 sg13g2_decap_8 FILLER_77_1514 ();
 sg13g2_decap_8 FILLER_77_1521 ();
 sg13g2_decap_8 FILLER_77_1528 ();
 sg13g2_decap_8 FILLER_77_1535 ();
 sg13g2_decap_8 FILLER_77_1542 ();
 sg13g2_decap_8 FILLER_77_1549 ();
 sg13g2_decap_8 FILLER_77_1556 ();
 sg13g2_decap_8 FILLER_77_1563 ();
 sg13g2_decap_8 FILLER_77_1570 ();
 sg13g2_decap_8 FILLER_77_1577 ();
 sg13g2_decap_8 FILLER_77_1584 ();
 sg13g2_decap_8 FILLER_77_1591 ();
 sg13g2_decap_8 FILLER_77_1598 ();
 sg13g2_decap_8 FILLER_77_1605 ();
 sg13g2_decap_8 FILLER_77_1612 ();
 sg13g2_decap_8 FILLER_77_1619 ();
 sg13g2_decap_8 FILLER_77_1626 ();
 sg13g2_decap_8 FILLER_77_1633 ();
 sg13g2_decap_8 FILLER_77_1640 ();
 sg13g2_decap_8 FILLER_77_1647 ();
 sg13g2_decap_8 FILLER_77_1654 ();
 sg13g2_decap_8 FILLER_77_1661 ();
 sg13g2_decap_8 FILLER_77_1668 ();
 sg13g2_decap_8 FILLER_77_1675 ();
 sg13g2_decap_8 FILLER_77_1682 ();
 sg13g2_decap_8 FILLER_77_1689 ();
 sg13g2_decap_8 FILLER_77_1696 ();
 sg13g2_decap_8 FILLER_77_1703 ();
 sg13g2_decap_8 FILLER_77_1710 ();
 sg13g2_decap_8 FILLER_77_1717 ();
 sg13g2_decap_8 FILLER_77_1724 ();
 sg13g2_decap_8 FILLER_77_1731 ();
 sg13g2_decap_8 FILLER_77_1738 ();
 sg13g2_decap_8 FILLER_77_1745 ();
 sg13g2_decap_8 FILLER_77_1752 ();
 sg13g2_decap_8 FILLER_77_1759 ();
 sg13g2_fill_2 FILLER_77_1766 ();
 sg13g2_decap_4 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_4 ();
 sg13g2_fill_2 FILLER_78_28 ();
 sg13g2_fill_1 FILLER_78_75 ();
 sg13g2_fill_1 FILLER_78_103 ();
 sg13g2_fill_2 FILLER_78_131 ();
 sg13g2_fill_2 FILLER_78_162 ();
 sg13g2_decap_8 FILLER_78_178 ();
 sg13g2_fill_1 FILLER_78_185 ();
 sg13g2_decap_4 FILLER_78_229 ();
 sg13g2_fill_1 FILLER_78_233 ();
 sg13g2_fill_1 FILLER_78_275 ();
 sg13g2_fill_2 FILLER_78_378 ();
 sg13g2_fill_2 FILLER_78_425 ();
 sg13g2_fill_1 FILLER_78_427 ();
 sg13g2_fill_1 FILLER_78_471 ();
 sg13g2_fill_2 FILLER_78_512 ();
 sg13g2_fill_1 FILLER_78_541 ();
 sg13g2_fill_1 FILLER_78_625 ();
 sg13g2_fill_2 FILLER_78_667 ();
 sg13g2_fill_2 FILLER_78_702 ();
 sg13g2_fill_1 FILLER_78_704 ();
 sg13g2_fill_1 FILLER_78_721 ();
 sg13g2_decap_4 FILLER_78_733 ();
 sg13g2_fill_2 FILLER_78_741 ();
 sg13g2_decap_4 FILLER_78_760 ();
 sg13g2_fill_2 FILLER_78_764 ();
 sg13g2_decap_4 FILLER_78_770 ();
 sg13g2_fill_1 FILLER_78_774 ();
 sg13g2_fill_2 FILLER_78_785 ();
 sg13g2_fill_2 FILLER_78_792 ();
 sg13g2_decap_4 FILLER_78_808 ();
 sg13g2_fill_1 FILLER_78_812 ();
 sg13g2_fill_1 FILLER_78_823 ();
 sg13g2_fill_1 FILLER_78_828 ();
 sg13g2_decap_8 FILLER_78_837 ();
 sg13g2_fill_1 FILLER_78_844 ();
 sg13g2_fill_2 FILLER_78_855 ();
 sg13g2_fill_2 FILLER_78_862 ();
 sg13g2_fill_2 FILLER_78_869 ();
 sg13g2_fill_1 FILLER_78_871 ();
 sg13g2_decap_4 FILLER_78_876 ();
 sg13g2_fill_1 FILLER_78_880 ();
 sg13g2_fill_2 FILLER_78_886 ();
 sg13g2_decap_4 FILLER_78_893 ();
 sg13g2_fill_1 FILLER_78_897 ();
 sg13g2_fill_2 FILLER_78_912 ();
 sg13g2_decap_8 FILLER_78_922 ();
 sg13g2_fill_2 FILLER_78_929 ();
 sg13g2_fill_1 FILLER_78_940 ();
 sg13g2_fill_2 FILLER_78_951 ();
 sg13g2_fill_1 FILLER_78_953 ();
 sg13g2_decap_4 FILLER_78_958 ();
 sg13g2_fill_1 FILLER_78_988 ();
 sg13g2_decap_4 FILLER_78_993 ();
 sg13g2_fill_2 FILLER_78_1005 ();
 sg13g2_fill_1 FILLER_78_1007 ();
 sg13g2_fill_1 FILLER_78_1013 ();
 sg13g2_fill_2 FILLER_78_1019 ();
 sg13g2_fill_1 FILLER_78_1021 ();
 sg13g2_fill_2 FILLER_78_1027 ();
 sg13g2_decap_8 FILLER_78_1080 ();
 sg13g2_fill_1 FILLER_78_1087 ();
 sg13g2_fill_2 FILLER_78_1193 ();
 sg13g2_fill_1 FILLER_78_1195 ();
 sg13g2_fill_2 FILLER_78_1288 ();
 sg13g2_fill_1 FILLER_78_1290 ();
 sg13g2_fill_2 FILLER_78_1321 ();
 sg13g2_fill_1 FILLER_78_1323 ();
 sg13g2_fill_1 FILLER_78_1333 ();
 sg13g2_decap_8 FILLER_78_1347 ();
 sg13g2_decap_8 FILLER_78_1354 ();
 sg13g2_decap_8 FILLER_78_1361 ();
 sg13g2_decap_4 FILLER_78_1368 ();
 sg13g2_decap_8 FILLER_78_1442 ();
 sg13g2_fill_2 FILLER_78_1449 ();
 sg13g2_decap_4 FILLER_78_1455 ();
 sg13g2_fill_2 FILLER_78_1459 ();
 sg13g2_decap_4 FILLER_78_1471 ();
 sg13g2_decap_8 FILLER_78_1488 ();
 sg13g2_decap_8 FILLER_78_1495 ();
 sg13g2_decap_8 FILLER_78_1502 ();
 sg13g2_decap_8 FILLER_78_1509 ();
 sg13g2_decap_8 FILLER_78_1516 ();
 sg13g2_decap_8 FILLER_78_1523 ();
 sg13g2_decap_8 FILLER_78_1530 ();
 sg13g2_decap_8 FILLER_78_1537 ();
 sg13g2_decap_8 FILLER_78_1544 ();
 sg13g2_decap_8 FILLER_78_1551 ();
 sg13g2_decap_8 FILLER_78_1558 ();
 sg13g2_decap_8 FILLER_78_1565 ();
 sg13g2_decap_8 FILLER_78_1572 ();
 sg13g2_decap_8 FILLER_78_1579 ();
 sg13g2_decap_8 FILLER_78_1586 ();
 sg13g2_decap_8 FILLER_78_1593 ();
 sg13g2_decap_8 FILLER_78_1600 ();
 sg13g2_decap_8 FILLER_78_1607 ();
 sg13g2_decap_8 FILLER_78_1614 ();
 sg13g2_decap_8 FILLER_78_1621 ();
 sg13g2_decap_8 FILLER_78_1628 ();
 sg13g2_decap_8 FILLER_78_1635 ();
 sg13g2_decap_8 FILLER_78_1642 ();
 sg13g2_decap_8 FILLER_78_1649 ();
 sg13g2_decap_8 FILLER_78_1656 ();
 sg13g2_decap_8 FILLER_78_1663 ();
 sg13g2_decap_8 FILLER_78_1670 ();
 sg13g2_decap_8 FILLER_78_1677 ();
 sg13g2_decap_8 FILLER_78_1684 ();
 sg13g2_decap_8 FILLER_78_1691 ();
 sg13g2_decap_8 FILLER_78_1698 ();
 sg13g2_decap_8 FILLER_78_1705 ();
 sg13g2_decap_8 FILLER_78_1712 ();
 sg13g2_decap_8 FILLER_78_1719 ();
 sg13g2_decap_8 FILLER_78_1726 ();
 sg13g2_decap_8 FILLER_78_1733 ();
 sg13g2_decap_8 FILLER_78_1740 ();
 sg13g2_decap_8 FILLER_78_1747 ();
 sg13g2_decap_8 FILLER_78_1754 ();
 sg13g2_decap_8 FILLER_78_1761 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_fill_1 FILLER_79_21 ();
 sg13g2_fill_1 FILLER_79_35 ();
 sg13g2_fill_2 FILLER_79_64 ();
 sg13g2_fill_2 FILLER_79_110 ();
 sg13g2_fill_1 FILLER_79_112 ();
 sg13g2_fill_1 FILLER_79_122 ();
 sg13g2_fill_2 FILLER_79_153 ();
 sg13g2_fill_1 FILLER_79_195 ();
 sg13g2_decap_8 FILLER_79_212 ();
 sg13g2_decap_8 FILLER_79_219 ();
 sg13g2_fill_1 FILLER_79_230 ();
 sg13g2_fill_1 FILLER_79_235 ();
 sg13g2_fill_2 FILLER_79_291 ();
 sg13g2_fill_1 FILLER_79_338 ();
 sg13g2_fill_1 FILLER_79_370 ();
 sg13g2_fill_1 FILLER_79_406 ();
 sg13g2_fill_2 FILLER_79_421 ();
 sg13g2_fill_2 FILLER_79_437 ();
 sg13g2_fill_2 FILLER_79_478 ();
 sg13g2_fill_1 FILLER_79_563 ();
 sg13g2_fill_1 FILLER_79_630 ();
 sg13g2_fill_2 FILLER_79_657 ();
 sg13g2_fill_1 FILLER_79_659 ();
 sg13g2_fill_2 FILLER_79_673 ();
 sg13g2_fill_1 FILLER_79_675 ();
 sg13g2_fill_1 FILLER_79_691 ();
 sg13g2_fill_1 FILLER_79_697 ();
 sg13g2_fill_2 FILLER_79_708 ();
 sg13g2_fill_2 FILLER_79_807 ();
 sg13g2_fill_1 FILLER_79_809 ();
 sg13g2_fill_1 FILLER_79_819 ();
 sg13g2_fill_2 FILLER_79_878 ();
 sg13g2_fill_1 FILLER_79_880 ();
 sg13g2_fill_1 FILLER_79_891 ();
 sg13g2_fill_2 FILLER_79_938 ();
 sg13g2_fill_1 FILLER_79_981 ();
 sg13g2_fill_2 FILLER_79_992 ();
 sg13g2_fill_1 FILLER_79_1020 ();
 sg13g2_fill_1 FILLER_79_1050 ();
 sg13g2_fill_2 FILLER_79_1068 ();
 sg13g2_fill_2 FILLER_79_1089 ();
 sg13g2_fill_1 FILLER_79_1103 ();
 sg13g2_fill_1 FILLER_79_1255 ();
 sg13g2_fill_1 FILLER_79_1261 ();
 sg13g2_fill_2 FILLER_79_1280 ();
 sg13g2_fill_1 FILLER_79_1322 ();
 sg13g2_decap_8 FILLER_79_1327 ();
 sg13g2_decap_8 FILLER_79_1334 ();
 sg13g2_decap_8 FILLER_79_1341 ();
 sg13g2_decap_8 FILLER_79_1348 ();
 sg13g2_decap_8 FILLER_79_1355 ();
 sg13g2_decap_8 FILLER_79_1362 ();
 sg13g2_decap_8 FILLER_79_1369 ();
 sg13g2_decap_8 FILLER_79_1376 ();
 sg13g2_decap_8 FILLER_79_1395 ();
 sg13g2_decap_8 FILLER_79_1402 ();
 sg13g2_decap_8 FILLER_79_1409 ();
 sg13g2_decap_4 FILLER_79_1416 ();
 sg13g2_decap_4 FILLER_79_1424 ();
 sg13g2_fill_2 FILLER_79_1428 ();
 sg13g2_decap_8 FILLER_79_1438 ();
 sg13g2_decap_8 FILLER_79_1445 ();
 sg13g2_decap_8 FILLER_79_1452 ();
 sg13g2_decap_8 FILLER_79_1459 ();
 sg13g2_decap_8 FILLER_79_1466 ();
 sg13g2_decap_8 FILLER_79_1473 ();
 sg13g2_decap_8 FILLER_79_1480 ();
 sg13g2_decap_8 FILLER_79_1487 ();
 sg13g2_decap_8 FILLER_79_1494 ();
 sg13g2_decap_8 FILLER_79_1501 ();
 sg13g2_decap_8 FILLER_79_1508 ();
 sg13g2_decap_8 FILLER_79_1515 ();
 sg13g2_decap_8 FILLER_79_1522 ();
 sg13g2_decap_8 FILLER_79_1529 ();
 sg13g2_decap_8 FILLER_79_1536 ();
 sg13g2_decap_8 FILLER_79_1543 ();
 sg13g2_decap_8 FILLER_79_1550 ();
 sg13g2_decap_8 FILLER_79_1557 ();
 sg13g2_decap_8 FILLER_79_1564 ();
 sg13g2_decap_8 FILLER_79_1571 ();
 sg13g2_decap_8 FILLER_79_1578 ();
 sg13g2_decap_8 FILLER_79_1585 ();
 sg13g2_decap_8 FILLER_79_1592 ();
 sg13g2_decap_8 FILLER_79_1599 ();
 sg13g2_decap_8 FILLER_79_1606 ();
 sg13g2_decap_8 FILLER_79_1613 ();
 sg13g2_decap_8 FILLER_79_1620 ();
 sg13g2_decap_8 FILLER_79_1627 ();
 sg13g2_decap_8 FILLER_79_1634 ();
 sg13g2_decap_8 FILLER_79_1641 ();
 sg13g2_decap_8 FILLER_79_1648 ();
 sg13g2_decap_8 FILLER_79_1655 ();
 sg13g2_decap_8 FILLER_79_1662 ();
 sg13g2_decap_8 FILLER_79_1669 ();
 sg13g2_decap_8 FILLER_79_1676 ();
 sg13g2_decap_8 FILLER_79_1683 ();
 sg13g2_decap_8 FILLER_79_1690 ();
 sg13g2_decap_8 FILLER_79_1697 ();
 sg13g2_decap_8 FILLER_79_1704 ();
 sg13g2_decap_8 FILLER_79_1711 ();
 sg13g2_decap_8 FILLER_79_1718 ();
 sg13g2_decap_8 FILLER_79_1725 ();
 sg13g2_decap_8 FILLER_79_1732 ();
 sg13g2_decap_8 FILLER_79_1739 ();
 sg13g2_decap_8 FILLER_79_1746 ();
 sg13g2_decap_8 FILLER_79_1753 ();
 sg13g2_decap_8 FILLER_79_1760 ();
 sg13g2_fill_1 FILLER_79_1767 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_4 FILLER_80_35 ();
 sg13g2_fill_2 FILLER_80_39 ();
 sg13g2_decap_8 FILLER_80_45 ();
 sg13g2_fill_2 FILLER_80_52 ();
 sg13g2_fill_2 FILLER_80_83 ();
 sg13g2_fill_1 FILLER_80_85 ();
 sg13g2_decap_8 FILLER_80_164 ();
 sg13g2_decap_8 FILLER_80_175 ();
 sg13g2_decap_8 FILLER_80_182 ();
 sg13g2_decap_8 FILLER_80_189 ();
 sg13g2_decap_8 FILLER_80_196 ();
 sg13g2_decap_8 FILLER_80_203 ();
 sg13g2_decap_8 FILLER_80_210 ();
 sg13g2_fill_1 FILLER_80_217 ();
 sg13g2_fill_2 FILLER_80_308 ();
 sg13g2_fill_1 FILLER_80_310 ();
 sg13g2_fill_2 FILLER_80_390 ();
 sg13g2_fill_1 FILLER_80_444 ();
 sg13g2_fill_2 FILLER_80_507 ();
 sg13g2_fill_1 FILLER_80_533 ();
 sg13g2_decap_4 FILLER_80_538 ();
 sg13g2_fill_2 FILLER_80_542 ();
 sg13g2_decap_8 FILLER_80_552 ();
 sg13g2_fill_2 FILLER_80_559 ();
 sg13g2_fill_1 FILLER_80_561 ();
 sg13g2_fill_2 FILLER_80_579 ();
 sg13g2_decap_4 FILLER_80_590 ();
 sg13g2_fill_2 FILLER_80_594 ();
 sg13g2_fill_2 FILLER_80_605 ();
 sg13g2_decap_4 FILLER_80_620 ();
 sg13g2_fill_1 FILLER_80_624 ();
 sg13g2_fill_2 FILLER_80_639 ();
 sg13g2_decap_8 FILLER_80_660 ();
 sg13g2_decap_8 FILLER_80_684 ();
 sg13g2_decap_8 FILLER_80_700 ();
 sg13g2_decap_4 FILLER_80_707 ();
 sg13g2_fill_2 FILLER_80_711 ();
 sg13g2_fill_2 FILLER_80_722 ();
 sg13g2_fill_1 FILLER_80_724 ();
 sg13g2_decap_8 FILLER_80_734 ();
 sg13g2_decap_4 FILLER_80_741 ();
 sg13g2_fill_2 FILLER_80_745 ();
 sg13g2_decap_4 FILLER_80_760 ();
 sg13g2_decap_4 FILLER_80_769 ();
 sg13g2_fill_1 FILLER_80_773 ();
 sg13g2_fill_1 FILLER_80_782 ();
 sg13g2_decap_4 FILLER_80_788 ();
 sg13g2_fill_2 FILLER_80_792 ();
 sg13g2_decap_8 FILLER_80_804 ();
 sg13g2_fill_2 FILLER_80_821 ();
 sg13g2_fill_1 FILLER_80_831 ();
 sg13g2_decap_8 FILLER_80_840 ();
 sg13g2_decap_8 FILLER_80_855 ();
 sg13g2_fill_1 FILLER_80_862 ();
 sg13g2_fill_1 FILLER_80_875 ();
 sg13g2_fill_1 FILLER_80_883 ();
 sg13g2_decap_8 FILLER_80_888 ();
 sg13g2_fill_1 FILLER_80_895 ();
 sg13g2_fill_1 FILLER_80_900 ();
 sg13g2_decap_4 FILLER_80_906 ();
 sg13g2_decap_4 FILLER_80_926 ();
 sg13g2_fill_2 FILLER_80_930 ();
 sg13g2_decap_8 FILLER_80_948 ();
 sg13g2_fill_1 FILLER_80_955 ();
 sg13g2_decap_4 FILLER_80_960 ();
 sg13g2_decap_4 FILLER_80_977 ();
 sg13g2_fill_2 FILLER_80_981 ();
 sg13g2_decap_8 FILLER_80_995 ();
 sg13g2_fill_2 FILLER_80_1002 ();
 sg13g2_fill_1 FILLER_80_1004 ();
 sg13g2_decap_8 FILLER_80_1014 ();
 sg13g2_fill_2 FILLER_80_1029 ();
 sg13g2_decap_8 FILLER_80_1040 ();
 sg13g2_decap_4 FILLER_80_1047 ();
 sg13g2_fill_1 FILLER_80_1051 ();
 sg13g2_fill_2 FILLER_80_1057 ();
 sg13g2_fill_1 FILLER_80_1059 ();
 sg13g2_decap_8 FILLER_80_1080 ();
 sg13g2_decap_4 FILLER_80_1087 ();
 sg13g2_fill_2 FILLER_80_1091 ();
 sg13g2_fill_2 FILLER_80_1154 ();
 sg13g2_fill_1 FILLER_80_1156 ();
 sg13g2_fill_2 FILLER_80_1224 ();
 sg13g2_fill_1 FILLER_80_1226 ();
 sg13g2_fill_2 FILLER_80_1254 ();
 sg13g2_fill_1 FILLER_80_1256 ();
 sg13g2_decap_8 FILLER_80_1312 ();
 sg13g2_decap_8 FILLER_80_1319 ();
 sg13g2_decap_8 FILLER_80_1326 ();
 sg13g2_decap_8 FILLER_80_1333 ();
 sg13g2_decap_8 FILLER_80_1340 ();
 sg13g2_decap_8 FILLER_80_1347 ();
 sg13g2_decap_8 FILLER_80_1354 ();
 sg13g2_decap_8 FILLER_80_1361 ();
 sg13g2_decap_8 FILLER_80_1368 ();
 sg13g2_decap_8 FILLER_80_1375 ();
 sg13g2_decap_8 FILLER_80_1382 ();
 sg13g2_decap_8 FILLER_80_1389 ();
 sg13g2_decap_8 FILLER_80_1396 ();
 sg13g2_decap_8 FILLER_80_1403 ();
 sg13g2_decap_8 FILLER_80_1410 ();
 sg13g2_decap_8 FILLER_80_1417 ();
 sg13g2_decap_8 FILLER_80_1424 ();
 sg13g2_decap_8 FILLER_80_1431 ();
 sg13g2_decap_8 FILLER_80_1438 ();
 sg13g2_decap_8 FILLER_80_1445 ();
 sg13g2_decap_8 FILLER_80_1452 ();
 sg13g2_decap_8 FILLER_80_1459 ();
 sg13g2_decap_8 FILLER_80_1466 ();
 sg13g2_decap_8 FILLER_80_1473 ();
 sg13g2_decap_8 FILLER_80_1480 ();
 sg13g2_decap_8 FILLER_80_1487 ();
 sg13g2_decap_8 FILLER_80_1494 ();
 sg13g2_decap_8 FILLER_80_1501 ();
 sg13g2_decap_8 FILLER_80_1508 ();
 sg13g2_decap_8 FILLER_80_1515 ();
 sg13g2_decap_8 FILLER_80_1522 ();
 sg13g2_decap_8 FILLER_80_1529 ();
 sg13g2_decap_8 FILLER_80_1536 ();
 sg13g2_decap_8 FILLER_80_1543 ();
 sg13g2_decap_8 FILLER_80_1550 ();
 sg13g2_decap_8 FILLER_80_1557 ();
 sg13g2_decap_8 FILLER_80_1564 ();
 sg13g2_decap_8 FILLER_80_1571 ();
 sg13g2_decap_8 FILLER_80_1578 ();
 sg13g2_decap_8 FILLER_80_1585 ();
 sg13g2_decap_8 FILLER_80_1592 ();
 sg13g2_decap_8 FILLER_80_1599 ();
 sg13g2_decap_8 FILLER_80_1606 ();
 sg13g2_decap_8 FILLER_80_1613 ();
 sg13g2_decap_8 FILLER_80_1620 ();
 sg13g2_decap_8 FILLER_80_1627 ();
 sg13g2_decap_8 FILLER_80_1634 ();
 sg13g2_decap_8 FILLER_80_1641 ();
 sg13g2_decap_8 FILLER_80_1648 ();
 sg13g2_decap_8 FILLER_80_1655 ();
 sg13g2_decap_8 FILLER_80_1662 ();
 sg13g2_decap_8 FILLER_80_1669 ();
 sg13g2_decap_8 FILLER_80_1676 ();
 sg13g2_decap_8 FILLER_80_1683 ();
 sg13g2_decap_8 FILLER_80_1690 ();
 sg13g2_decap_8 FILLER_80_1697 ();
 sg13g2_decap_8 FILLER_80_1704 ();
 sg13g2_decap_8 FILLER_80_1711 ();
 sg13g2_decap_8 FILLER_80_1718 ();
 sg13g2_decap_8 FILLER_80_1725 ();
 sg13g2_decap_8 FILLER_80_1732 ();
 sg13g2_decap_8 FILLER_80_1739 ();
 sg13g2_decap_8 FILLER_80_1746 ();
 sg13g2_decap_8 FILLER_80_1753 ();
 sg13g2_decap_8 FILLER_80_1760 ();
 sg13g2_fill_1 FILLER_80_1767 ();
endmodule
