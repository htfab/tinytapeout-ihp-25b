module tt_um_wokwi_434925031692840961 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net109;
 wire net110;
 wire params_ready;
 wire spike_out;
 wire \system_inst.leak_cycles[0] ;
 wire \system_inst.leak_cycles[1] ;
 wire \system_inst.leak_cycles[2] ;
 wire \system_inst.leak_cycles[3] ;
 wire \system_inst.leak_rate[0] ;
 wire \system_inst.leak_rate[1] ;
 wire \system_inst.leak_rate[2] ;
 wire \system_inst.leak_rate[3] ;
 wire \system_inst.leak_rate[4] ;
 wire \system_inst.leak_rate[5] ;
 wire \system_inst.leak_rate[6] ;
 wire \system_inst.leak_rate[7] ;
 wire \system_inst.loader.bit_count[0] ;
 wire \system_inst.loader.bit_count[1] ;
 wire \system_inst.loader.bit_count[2] ;
 wire \system_inst.loader.current_state[0] ;
 wire \system_inst.loader.current_state[1] ;
 wire \system_inst.loader.current_state[2] ;
 wire \system_inst.loader.current_state[3] ;
 wire \system_inst.loader.current_state[5] ;
 wire \system_inst.loader.shift_reg[0] ;
 wire \system_inst.loader.shift_reg[1] ;
 wire \system_inst.loader.shift_reg[2] ;
 wire \system_inst.loader.shift_reg[3] ;
 wire \system_inst.loader.shift_reg[4] ;
 wire \system_inst.loader.shift_reg[5] ;
 wire \system_inst.loader.shift_reg[6] ;
 wire \system_inst.loader.threshold[0] ;
 wire \system_inst.loader.threshold[1] ;
 wire \system_inst.loader.threshold[2] ;
 wire \system_inst.loader.threshold[3] ;
 wire \system_inst.loader.threshold[4] ;
 wire \system_inst.loader.threshold[5] ;
 wire \system_inst.loader.threshold[6] ;
 wire \system_inst.loader.threshold[7] ;
 wire \system_inst.loader.weight_a[0] ;
 wire \system_inst.loader.weight_a[1] ;
 wire \system_inst.loader.weight_a[2] ;
 wire \system_inst.neuron.leak_counter[0] ;
 wire \system_inst.neuron.leak_counter[1] ;
 wire \system_inst.neuron.leak_counter[2] ;
 wire \system_inst.neuron.leak_counter[3] ;
 wire \system_inst.neuron.refr_cnt[0] ;
 wire \system_inst.neuron.refr_cnt[1] ;
 wire \system_inst.neuron.refr_cnt[2] ;
 wire \system_inst.neuron.refr_cnt[3] ;
 wire \system_inst.neuron.v_mem[0] ;
 wire \system_inst.neuron.v_mem[1] ;
 wire \system_inst.neuron.v_mem[2] ;
 wire \system_inst.neuron.v_mem[3] ;
 wire \system_inst.neuron.v_mem[4] ;
 wire \system_inst.neuron.v_mem[5] ;
 wire \system_inst.neuron.v_mem[6] ;
 wire \system_inst.neuron.v_mem[7] ;
 wire \system_inst.neuron.v_mem[8] ;
 wire clknet_0_clk;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;

 sg13g2_inv_1 _0515_ (.Y(_0060_),
    .A(net199));
 sg13g2_inv_2 _0516_ (.Y(_0061_),
    .A(net162));
 sg13g2_inv_1 _0517_ (.Y(_0062_),
    .A(net148));
 sg13g2_inv_1 _0518_ (.Y(_0063_),
    .A(net145));
 sg13g2_inv_1 _0519_ (.Y(_0064_),
    .A(net117));
 sg13g2_inv_1 _0520_ (.Y(_0065_),
    .A(net150));
 sg13g2_inv_1 _0521_ (.Y(_0066_),
    .A(net138));
 sg13g2_inv_1 _0522_ (.Y(_0067_),
    .A(net129));
 sg13g2_inv_1 _0523_ (.Y(_0068_),
    .A(net156));
 sg13g2_inv_1 _0524_ (.Y(_0069_),
    .A(net179));
 sg13g2_inv_1 _0525_ (.Y(_0070_),
    .A(net142));
 sg13g2_inv_1 _0526_ (.Y(_0071_),
    .A(\system_inst.loader.threshold[1] ));
 sg13g2_inv_1 _0527_ (.Y(_0072_),
    .A(net136));
 sg13g2_inv_1 _0528_ (.Y(_0073_),
    .A(net154));
 sg13g2_inv_1 _0529_ (.Y(_0074_),
    .A(net133));
 sg13g2_inv_1 _0530_ (.Y(_0075_),
    .A(net167));
 sg13g2_inv_1 _0531_ (.Y(_0076_),
    .A(net165));
 sg13g2_inv_1 _0532_ (.Y(_0077_),
    .A(net160));
 sg13g2_inv_1 _0533_ (.Y(_0078_),
    .A(net183));
 sg13g2_inv_1 _0534_ (.Y(_0079_),
    .A(net121));
 sg13g2_inv_1 _0535_ (.Y(_0080_),
    .A(net115));
 sg13g2_inv_1 _0536_ (.Y(_0081_),
    .A(net128));
 sg13g2_inv_1 _0537_ (.Y(_0082_),
    .A(net107));
 sg13g2_inv_1 _0538_ (.Y(_0083_),
    .A(net152));
 sg13g2_inv_1 _0539_ (.Y(_0084_),
    .A(\system_inst.loader.current_state[0] ));
 sg13g2_nand2b_1 _0540_ (.Y(_0085_),
    .B(net106),
    .A_N(net1));
 sg13g2_nand2_1 _0541_ (.Y(_0086_),
    .A(net131),
    .B(\system_inst.loader.bit_count[0] ));
 sg13g2_nor2_1 _0542_ (.A(_0005_),
    .B(_0086_),
    .Y(_0087_));
 sg13g2_and2_2 _0543_ (.A(net4),
    .B(net1),
    .X(_0088_));
 sg13g2_nand2_1 _0544_ (.Y(_0089_),
    .A(net106),
    .B(_0088_));
 sg13g2_o21ai_1 _0545_ (.B1(_0085_),
    .Y(_0090_),
    .A1(_0087_),
    .A2(_0089_));
 sg13g2_and3_2 _0546_ (.X(_0091_),
    .A(net172),
    .B(net94),
    .C(_0088_));
 sg13g2_nand3_1 _0547_ (.B(net94),
    .C(_0088_),
    .A(\system_inst.loader.current_state[5] ),
    .Y(_0092_));
 sg13g2_a22oi_1 _0548_ (.Y(_0093_),
    .B1(_0091_),
    .B2(net106),
    .A2(_0090_),
    .A1(net152));
 sg13g2_inv_1 _0549_ (.Y(_0001_),
    .A(net153));
 sg13g2_and3_1 _0550_ (.X(_0094_),
    .A(\system_inst.loader.current_state[2] ),
    .B(_0087_),
    .C(_0088_));
 sg13g2_nand3_1 _0551_ (.B(net94),
    .C(_0088_),
    .A(\system_inst.loader.current_state[2] ),
    .Y(_0095_));
 sg13g2_a22oi_1 _0552_ (.Y(_0096_),
    .B1(_0094_),
    .B2(net106),
    .A2(_0090_),
    .A1(net172));
 sg13g2_inv_1 _0553_ (.Y(_0004_),
    .A(net173));
 sg13g2_nor2_1 _0554_ (.A(net127),
    .B(_0085_),
    .Y(_0097_));
 sg13g2_a21oi_1 _0555_ (.A1(net106),
    .A2(_0088_),
    .Y(_0000_),
    .B1(_0097_));
 sg13g2_nand3_1 _0556_ (.B(net94),
    .C(_0088_),
    .A(net122),
    .Y(_0098_));
 sg13g2_inv_1 _0557_ (.Y(_0099_),
    .A(_0098_));
 sg13g2_a22oi_1 _0558_ (.Y(_0100_),
    .B1(_0099_),
    .B2(net106),
    .A2(_0090_),
    .A1(net174));
 sg13g2_inv_1 _0559_ (.Y(_0002_),
    .A(_0100_));
 sg13g2_nand2_1 _0560_ (.Y(_0101_),
    .A(net122),
    .B(_0090_));
 sg13g2_o21ai_1 _0561_ (.B1(_0101_),
    .Y(_0003_),
    .A1(_0084_),
    .A2(_0089_));
 sg13g2_nor2b_1 _0562_ (.A(net95),
    .B_N(\system_inst.neuron.v_mem[0] ),
    .Y(uo_out[1]));
 sg13g2_nor2b_1 _0563_ (.A(net95),
    .B_N(\system_inst.neuron.v_mem[1] ),
    .Y(uo_out[2]));
 sg13g2_nor2b_1 _0564_ (.A(net95),
    .B_N(\system_inst.neuron.v_mem[2] ),
    .Y(uo_out[3]));
 sg13g2_nor2b_1 _0565_ (.A(\system_inst.neuron.v_mem[8] ),
    .B_N(\system_inst.neuron.v_mem[3] ),
    .Y(uo_out[4]));
 sg13g2_nor2b_1 _0566_ (.A(net95),
    .B_N(\system_inst.neuron.v_mem[4] ),
    .Y(uo_out[5]));
 sg13g2_nor2b_1 _0567_ (.A(net95),
    .B_N(\system_inst.neuron.v_mem[5] ),
    .Y(uo_out[6]));
 sg13g2_nor2b_1 _0568_ (.A(net95),
    .B_N(\system_inst.neuron.v_mem[6] ),
    .Y(uo_out[7]));
 sg13g2_nor3_2 _0569_ (.A(\system_inst.loader.current_state[2] ),
    .B(\system_inst.loader.current_state[5] ),
    .C(\system_inst.loader.current_state[3] ),
    .Y(_0102_));
 sg13g2_nand2_1 _0570_ (.Y(_0103_),
    .A(_0007_),
    .B(_0102_));
 sg13g2_nor2_1 _0571_ (.A(net127),
    .B(_0103_),
    .Y(_0104_));
 sg13g2_o21ai_1 _0572_ (.B1(net1),
    .Y(_0105_),
    .A1(net4),
    .A2(_0084_));
 sg13g2_nor2_1 _0573_ (.A(_0104_),
    .B(_0105_),
    .Y(_0106_));
 sg13g2_o21ai_1 _0574_ (.B1(_0102_),
    .Y(_0107_),
    .A1(_0007_),
    .A2(net94));
 sg13g2_nand2_1 _0575_ (.Y(_0108_),
    .A(net4),
    .B(_0107_));
 sg13g2_nand2_1 _0576_ (.Y(_0109_),
    .A(_0106_),
    .B(_0108_));
 sg13g2_and2_2 _0577_ (.A(_0083_),
    .B(_0102_),
    .X(_0110_));
 sg13g2_a21oi_1 _0578_ (.A1(net187),
    .A2(_0109_),
    .Y(_0111_),
    .B1(net102));
 sg13g2_o21ai_1 _0579_ (.B1(_0111_),
    .Y(_0008_),
    .A1(_0109_),
    .A2(_0110_));
 sg13g2_o21ai_1 _0580_ (.B1(net108),
    .Y(_0112_),
    .A1(net5),
    .A2(_0098_));
 sg13g2_a21oi_1 _0581_ (.A1(_0081_),
    .A2(_0098_),
    .Y(_0009_),
    .B1(_0112_));
 sg13g2_a21oi_1 _0582_ (.A1(net98),
    .A2(_0098_),
    .Y(_0113_),
    .B1(net103));
 sg13g2_o21ai_1 _0583_ (.B1(_0113_),
    .Y(_0010_),
    .A1(_0061_),
    .A2(_0098_));
 sg13g2_o21ai_1 _0584_ (.B1(net106),
    .Y(_0114_),
    .A1(\system_inst.loader.shift_reg[1] ),
    .A2(_0098_));
 sg13g2_a21oi_1 _0585_ (.A1(_0080_),
    .A2(_0098_),
    .Y(_0011_),
    .B1(_0114_));
 sg13g2_o21ai_1 _0586_ (.B1(net107),
    .Y(_0115_),
    .A1(net5),
    .A2(net92));
 sg13g2_a21oi_1 _0587_ (.A1(_0079_),
    .A2(net92),
    .Y(_0012_),
    .B1(_0115_));
 sg13g2_a21oi_1 _0588_ (.A1(net191),
    .A2(net92),
    .Y(_0116_),
    .B1(net102));
 sg13g2_o21ai_1 _0589_ (.B1(_0116_),
    .Y(_0013_),
    .A1(_0061_),
    .A2(net92));
 sg13g2_o21ai_1 _0590_ (.B1(net107),
    .Y(_0117_),
    .A1(\system_inst.loader.shift_reg[1] ),
    .A2(net92));
 sg13g2_a21oi_1 _0591_ (.A1(_0078_),
    .A2(net92),
    .Y(_0014_),
    .B1(_0117_));
 sg13g2_o21ai_1 _0592_ (.B1(net105),
    .Y(_0118_),
    .A1(\system_inst.loader.shift_reg[2] ),
    .A2(net92));
 sg13g2_a21oi_1 _0593_ (.A1(_0077_),
    .A2(net92),
    .Y(_0015_),
    .B1(_0118_));
 sg13g2_o21ai_1 _0594_ (.B1(net105),
    .Y(_0119_),
    .A1(\system_inst.loader.shift_reg[3] ),
    .A2(net91));
 sg13g2_a21oi_1 _0595_ (.A1(_0076_),
    .A2(net91),
    .Y(_0016_),
    .B1(_0119_));
 sg13g2_o21ai_1 _0596_ (.B1(net104),
    .Y(_0120_),
    .A1(\system_inst.loader.shift_reg[4] ),
    .A2(net91));
 sg13g2_a21oi_1 _0597_ (.A1(_0075_),
    .A2(net91),
    .Y(_0017_),
    .B1(_0120_));
 sg13g2_o21ai_1 _0598_ (.B1(net105),
    .Y(_0121_),
    .A1(\system_inst.loader.shift_reg[5] ),
    .A2(net91));
 sg13g2_a21oi_1 _0599_ (.A1(_0074_),
    .A2(net91),
    .Y(_0018_),
    .B1(_0121_));
 sg13g2_o21ai_1 _0600_ (.B1(net104),
    .Y(_0122_),
    .A1(\system_inst.loader.shift_reg[6] ),
    .A2(net91));
 sg13g2_a21oi_1 _0601_ (.A1(_0073_),
    .A2(net91),
    .Y(_0019_),
    .B1(_0122_));
 sg13g2_o21ai_1 _0602_ (.B1(net107),
    .Y(_0123_),
    .A1(net5),
    .A2(_0092_));
 sg13g2_a21oi_1 _0603_ (.A1(_0072_),
    .A2(_0092_),
    .Y(_0020_),
    .B1(_0123_));
 sg13g2_a21oi_1 _0604_ (.A1(net140),
    .A2(net93),
    .Y(_0124_),
    .B1(net102));
 sg13g2_o21ai_1 _0605_ (.B1(_0124_),
    .Y(_0021_),
    .A1(_0061_),
    .A2(net93));
 sg13g2_a21oi_1 _0606_ (.A1(\system_inst.loader.shift_reg[1] ),
    .A2(_0091_),
    .Y(_0125_),
    .B1(net101));
 sg13g2_o21ai_1 _0607_ (.B1(_0125_),
    .Y(_0022_),
    .A1(_0070_),
    .A2(_0091_));
 sg13g2_a21oi_1 _0608_ (.A1(\system_inst.loader.shift_reg[2] ),
    .A2(_0091_),
    .Y(_0126_),
    .B1(net101));
 sg13g2_o21ai_1 _0609_ (.B1(_0126_),
    .Y(_0023_),
    .A1(_0069_),
    .A2(_0091_));
 sg13g2_a21oi_1 _0610_ (.A1(\system_inst.loader.shift_reg[3] ),
    .A2(_0091_),
    .Y(_0127_),
    .B1(net101));
 sg13g2_o21ai_1 _0611_ (.B1(_0127_),
    .Y(_0024_),
    .A1(_0068_),
    .A2(_0091_));
 sg13g2_o21ai_1 _0612_ (.B1(net104),
    .Y(_0128_),
    .A1(\system_inst.loader.shift_reg[4] ),
    .A2(net93));
 sg13g2_a21oi_1 _0613_ (.A1(_0067_),
    .A2(net93),
    .Y(_0025_),
    .B1(_0128_));
 sg13g2_o21ai_1 _0614_ (.B1(net104),
    .Y(_0129_),
    .A1(\system_inst.loader.shift_reg[5] ),
    .A2(net93));
 sg13g2_a21oi_1 _0615_ (.A1(_0066_),
    .A2(net93),
    .Y(_0026_),
    .B1(_0129_));
 sg13g2_o21ai_1 _0616_ (.B1(net104),
    .Y(_0130_),
    .A1(\system_inst.loader.shift_reg[6] ),
    .A2(net93));
 sg13g2_a21oi_1 _0617_ (.A1(_0065_),
    .A2(net93),
    .Y(_0027_),
    .B1(_0130_));
 sg13g2_nand3_1 _0618_ (.B(net94),
    .C(_0088_),
    .A(net152),
    .Y(_0131_));
 sg13g2_o21ai_1 _0619_ (.B1(net108),
    .Y(_0132_),
    .A1(net5),
    .A2(_0131_));
 sg13g2_a21oi_1 _0620_ (.A1(_0064_),
    .A2(_0131_),
    .Y(_0028_),
    .B1(_0132_));
 sg13g2_a21oi_1 _0621_ (.A1(net171),
    .A2(_0131_),
    .Y(_0133_),
    .B1(net102));
 sg13g2_o21ai_1 _0622_ (.B1(_0133_),
    .Y(_0029_),
    .A1(_0061_),
    .A2(_0131_));
 sg13g2_o21ai_1 _0623_ (.B1(net108),
    .Y(_0134_),
    .A1(\system_inst.loader.shift_reg[1] ),
    .A2(_0131_));
 sg13g2_a21oi_1 _0624_ (.A1(_0063_),
    .A2(_0131_),
    .Y(_0030_),
    .B1(_0134_));
 sg13g2_o21ai_1 _0625_ (.B1(net106),
    .Y(_0135_),
    .A1(\system_inst.loader.shift_reg[2] ),
    .A2(_0131_));
 sg13g2_a21oi_1 _0626_ (.A1(_0062_),
    .A2(_0131_),
    .Y(_0031_),
    .B1(_0135_));
 sg13g2_nor2_1 _0627_ (.A(net4),
    .B(_0110_),
    .Y(_0136_));
 sg13g2_nor2b_2 _0628_ (.A(_0136_),
    .B_N(_0106_),
    .Y(_0137_));
 sg13g2_nand2b_1 _0629_ (.Y(_0138_),
    .B(_0106_),
    .A_N(_0136_));
 sg13g2_a21oi_2 _0630_ (.B1(_0110_),
    .Y(_0139_),
    .A2(net94),
    .A1(_0083_));
 sg13g2_a21oi_1 _0631_ (.A1(net5),
    .A2(_0139_),
    .Y(_0140_),
    .B1(_0138_));
 sg13g2_o21ai_1 _0632_ (.B1(net107),
    .Y(_0141_),
    .A1(net162),
    .A2(_0137_));
 sg13g2_nor2_1 _0633_ (.A(_0140_),
    .B(_0141_),
    .Y(_0032_));
 sg13g2_a21oi_1 _0634_ (.A1(net162),
    .A2(_0139_),
    .Y(_0142_),
    .B1(_0138_));
 sg13g2_o21ai_1 _0635_ (.B1(net107),
    .Y(_0143_),
    .A1(\system_inst.loader.shift_reg[1] ),
    .A2(_0137_));
 sg13g2_nor2_1 _0636_ (.A(_0142_),
    .B(_0143_),
    .Y(_0033_));
 sg13g2_a21oi_1 _0637_ (.A1(net198),
    .A2(_0139_),
    .Y(_0144_),
    .B1(net86));
 sg13g2_o21ai_1 _0638_ (.B1(net105),
    .Y(_0145_),
    .A1(net192),
    .A2(_0137_));
 sg13g2_nor2_1 _0639_ (.A(_0144_),
    .B(_0145_),
    .Y(_0034_));
 sg13g2_a21oi_1 _0640_ (.A1(net192),
    .A2(_0139_),
    .Y(_0146_),
    .B1(net86));
 sg13g2_o21ai_1 _0641_ (.B1(net105),
    .Y(_0147_),
    .A1(net189),
    .A2(_0137_));
 sg13g2_nor2_1 _0642_ (.A(_0146_),
    .B(_0147_),
    .Y(_0035_));
 sg13g2_a21oi_1 _0643_ (.A1(net189),
    .A2(_0139_),
    .Y(_0148_),
    .B1(net86));
 sg13g2_o21ai_1 _0644_ (.B1(net104),
    .Y(_0149_),
    .A1(net178),
    .A2(_0137_));
 sg13g2_nor2_1 _0645_ (.A(_0148_),
    .B(_0149_),
    .Y(_0036_));
 sg13g2_a21oi_1 _0646_ (.A1(net178),
    .A2(_0139_),
    .Y(_0150_),
    .B1(net86));
 sg13g2_o21ai_1 _0647_ (.B1(net104),
    .Y(_0151_),
    .A1(net169),
    .A2(_0137_));
 sg13g2_nor2_1 _0648_ (.A(_0150_),
    .B(_0151_),
    .Y(_0037_));
 sg13g2_a21oi_1 _0649_ (.A1(net169),
    .A2(_0139_),
    .Y(_0152_),
    .B1(net86));
 sg13g2_o21ai_1 _0650_ (.B1(net104),
    .Y(_0153_),
    .A1(\system_inst.loader.shift_reg[6] ),
    .A2(_0137_));
 sg13g2_nor2_1 _0651_ (.A(_0152_),
    .B(_0153_),
    .Y(_0038_));
 sg13g2_nor2_2 _0652_ (.A(_0110_),
    .B(net86),
    .Y(_0154_));
 sg13g2_o21ai_1 _0653_ (.B1(net107),
    .Y(_0155_),
    .A1(net119),
    .A2(_0154_));
 sg13g2_a21oi_1 _0654_ (.A1(net119),
    .A2(_0137_),
    .Y(_0039_),
    .B1(_0155_));
 sg13g2_o21ai_1 _0655_ (.B1(_0103_),
    .Y(_0156_),
    .A1(net131),
    .A2(net119));
 sg13g2_nor2b_1 _0656_ (.A(_0156_),
    .B_N(_0086_),
    .Y(_0157_));
 sg13g2_a22oi_1 _0657_ (.Y(_0158_),
    .B1(_0154_),
    .B2(_0157_),
    .A2(net86),
    .A1(net131));
 sg13g2_nor2_1 _0658_ (.A(net102),
    .B(net132),
    .Y(_0040_));
 sg13g2_a22oi_1 _0659_ (.Y(_0159_),
    .B1(_0102_),
    .B2(_0007_),
    .A2(_0086_),
    .A1(_0005_));
 sg13g2_nor2b_1 _0660_ (.A(net94),
    .B_N(_0159_),
    .Y(_0160_));
 sg13g2_a22oi_1 _0661_ (.Y(_0161_),
    .B1(_0154_),
    .B2(_0160_),
    .A2(net86),
    .A1(net113));
 sg13g2_nor2_1 _0662_ (.A(net102),
    .B(net114),
    .Y(_0041_));
 sg13g2_nand3_1 _0663_ (.B(net97),
    .C(net7),
    .A(\system_inst.neuron.v_mem[3] ),
    .Y(_0162_));
 sg13g2_and2_1 _0664_ (.A(\system_inst.loader.weight_a[1] ),
    .B(net8),
    .X(_0163_));
 sg13g2_a21o_1 _0665_ (.A2(net7),
    .A1(net97),
    .B1(\system_inst.neuron.v_mem[3] ),
    .X(_0164_));
 sg13g2_nand3_1 _0666_ (.B(_0163_),
    .C(_0164_),
    .A(_0162_),
    .Y(_0165_));
 sg13g2_nand2_1 _0667_ (.Y(_0166_),
    .A(_0162_),
    .B(_0165_));
 sg13g2_nand2_1 _0668_ (.Y(_0167_),
    .A(net98),
    .B(net9));
 sg13g2_and3_1 _0669_ (.X(_0168_),
    .A(\system_inst.neuron.v_mem[4] ),
    .B(net96),
    .C(net8));
 sg13g2_nand3_1 _0670_ (.B(net97),
    .C(net8),
    .A(\system_inst.neuron.v_mem[4] ),
    .Y(_0169_));
 sg13g2_a21oi_1 _0671_ (.A1(net97),
    .A2(net8),
    .Y(_0170_),
    .B1(\system_inst.neuron.v_mem[4] ));
 sg13g2_nor2_1 _0672_ (.A(_0168_),
    .B(_0170_),
    .Y(_0171_));
 sg13g2_xnor2_1 _0673_ (.Y(_0172_),
    .A(_0167_),
    .B(_0171_));
 sg13g2_nand2_1 _0674_ (.Y(_0173_),
    .A(_0166_),
    .B(_0172_));
 sg13g2_nand2_1 _0675_ (.Y(_0174_),
    .A(net99),
    .B(net10));
 sg13g2_xnor2_1 _0676_ (.Y(_0175_),
    .A(_0166_),
    .B(_0172_));
 sg13g2_o21ai_1 _0677_ (.B1(_0173_),
    .Y(_0176_),
    .A1(_0174_),
    .A2(_0175_));
 sg13g2_nand2_1 _0678_ (.Y(_0177_),
    .A(net99),
    .B(net11));
 sg13g2_o21ai_1 _0679_ (.B1(_0169_),
    .Y(_0178_),
    .A1(_0167_),
    .A2(_0170_));
 sg13g2_nand2_1 _0680_ (.Y(_0179_),
    .A(net98),
    .B(net10));
 sg13g2_nand3_1 _0681_ (.B(net96),
    .C(net9),
    .A(\system_inst.neuron.v_mem[5] ),
    .Y(_0180_));
 sg13g2_a21o_1 _0682_ (.A2(net9),
    .A1(net96),
    .B1(\system_inst.neuron.v_mem[5] ),
    .X(_0181_));
 sg13g2_nand2_1 _0683_ (.Y(_0182_),
    .A(_0180_),
    .B(_0181_));
 sg13g2_xor2_1 _0684_ (.B(_0182_),
    .A(_0179_),
    .X(_0183_));
 sg13g2_nand2_1 _0685_ (.Y(_0184_),
    .A(_0178_),
    .B(_0183_));
 sg13g2_xnor2_1 _0686_ (.Y(_0185_),
    .A(_0178_),
    .B(_0183_));
 sg13g2_xor2_1 _0687_ (.B(_0185_),
    .A(_0177_),
    .X(_0186_));
 sg13g2_and2_1 _0688_ (.A(_0176_),
    .B(_0186_),
    .X(_0187_));
 sg13g2_nand3_1 _0689_ (.B(net97),
    .C(net6),
    .A(\system_inst.neuron.v_mem[2] ),
    .Y(_0188_));
 sg13g2_nand2_1 _0690_ (.Y(_0189_),
    .A(net98),
    .B(net7));
 sg13g2_a21oi_1 _0691_ (.A1(net97),
    .A2(net6),
    .Y(_0190_),
    .B1(\system_inst.neuron.v_mem[2] ));
 sg13g2_a21o_1 _0692_ (.A2(net6),
    .A1(net97),
    .B1(\system_inst.neuron.v_mem[2] ),
    .X(_0191_));
 sg13g2_and4_1 _0693_ (.A(net98),
    .B(net7),
    .C(_0188_),
    .D(_0191_),
    .X(_0192_));
 sg13g2_o21ai_1 _0694_ (.B1(_0188_),
    .Y(_0193_),
    .A1(_0189_),
    .A2(_0190_));
 sg13g2_a21o_1 _0695_ (.A2(_0164_),
    .A1(_0162_),
    .B1(_0163_),
    .X(_0194_));
 sg13g2_nand3_1 _0696_ (.B(_0193_),
    .C(_0194_),
    .A(_0165_),
    .Y(_0195_));
 sg13g2_a21o_1 _0697_ (.A2(_0194_),
    .A1(_0165_),
    .B1(_0193_),
    .X(_0196_));
 sg13g2_and4_1 _0698_ (.A(net99),
    .B(net9),
    .C(_0195_),
    .D(_0196_),
    .X(_0197_));
 sg13g2_nand4_1 _0699_ (.B(net9),
    .C(_0195_),
    .A(net99),
    .Y(_0198_),
    .D(_0196_));
 sg13g2_nand2_1 _0700_ (.Y(_0199_),
    .A(_0195_),
    .B(_0198_));
 sg13g2_xor2_1 _0701_ (.B(_0175_),
    .A(_0174_),
    .X(_0200_));
 sg13g2_nand2_1 _0702_ (.Y(_0201_),
    .A(_0199_),
    .B(_0200_));
 sg13g2_nand3_1 _0703_ (.B(\system_inst.loader.weight_a[1] ),
    .C(net6),
    .A(\system_inst.neuron.v_mem[1] ),
    .Y(_0202_));
 sg13g2_a22oi_1 _0704_ (.Y(_0203_),
    .B1(_0188_),
    .B2(_0191_),
    .A2(net7),
    .A1(net98));
 sg13g2_nor3_1 _0705_ (.A(_0192_),
    .B(_0202_),
    .C(_0203_),
    .Y(_0204_));
 sg13g2_or3_1 _0706_ (.A(_0192_),
    .B(_0202_),
    .C(_0203_),
    .X(_0205_));
 sg13g2_and2_1 _0707_ (.A(net99),
    .B(net8),
    .X(_0206_));
 sg13g2_nand2_1 _0708_ (.Y(_0207_),
    .A(net99),
    .B(net8));
 sg13g2_o21ai_1 _0709_ (.B1(_0202_),
    .Y(_0208_),
    .A1(_0192_),
    .A2(_0203_));
 sg13g2_a21oi_1 _0710_ (.A1(_0206_),
    .A2(_0208_),
    .Y(_0209_),
    .B1(_0204_));
 sg13g2_a22oi_1 _0711_ (.Y(_0210_),
    .B1(_0195_),
    .B2(_0196_),
    .A2(net9),
    .A1(net99));
 sg13g2_nor3_1 _0712_ (.A(_0197_),
    .B(_0209_),
    .C(_0210_),
    .Y(_0211_));
 sg13g2_nand2_1 _0713_ (.Y(_0212_),
    .A(net99),
    .B(net7));
 sg13g2_a21o_1 _0714_ (.A2(net6),
    .A1(net98),
    .B1(\system_inst.neuron.v_mem[1] ),
    .X(_0213_));
 sg13g2_nand2_1 _0715_ (.Y(_0214_),
    .A(_0202_),
    .B(_0213_));
 sg13g2_or2_1 _0716_ (.X(_0215_),
    .B(_0214_),
    .A(_0212_));
 sg13g2_nand3_1 _0717_ (.B(_0207_),
    .C(_0208_),
    .A(_0205_),
    .Y(_0216_));
 sg13g2_a21o_1 _0718_ (.A2(_0208_),
    .A1(_0205_),
    .B1(_0207_),
    .X(_0217_));
 sg13g2_a21o_1 _0719_ (.A2(_0217_),
    .A1(_0216_),
    .B1(_0215_),
    .X(_0218_));
 sg13g2_xor2_1 _0720_ (.B(_0214_),
    .A(_0212_),
    .X(_0219_));
 sg13g2_nand2_1 _0721_ (.Y(_0220_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net6));
 sg13g2_nor2_1 _0722_ (.A(_0006_),
    .B(_0220_),
    .Y(_0221_));
 sg13g2_nand2_1 _0723_ (.Y(_0222_),
    .A(_0219_),
    .B(_0221_));
 sg13g2_a21oi_1 _0724_ (.A1(_0216_),
    .A2(_0217_),
    .Y(_0223_),
    .B1(_0222_));
 sg13g2_a22oi_1 _0725_ (.Y(_0224_),
    .B1(_0222_),
    .B2(_0215_),
    .A2(_0217_),
    .A1(_0216_));
 sg13g2_o21ai_1 _0726_ (.B1(_0209_),
    .Y(_0225_),
    .A1(_0197_),
    .A2(_0210_));
 sg13g2_nor2b_1 _0727_ (.A(_0211_),
    .B_N(_0225_),
    .Y(_0226_));
 sg13g2_a21oi_1 _0728_ (.A1(_0224_),
    .A2(_0225_),
    .Y(_0227_),
    .B1(_0211_));
 sg13g2_xnor2_1 _0729_ (.Y(_0228_),
    .A(_0199_),
    .B(_0200_));
 sg13g2_o21ai_1 _0730_ (.B1(_0201_),
    .Y(_0229_),
    .A1(_0227_),
    .A2(_0228_));
 sg13g2_xnor2_1 _0731_ (.Y(_0230_),
    .A(_0176_),
    .B(_0186_));
 sg13g2_inv_1 _0732_ (.Y(_0231_),
    .A(_0230_));
 sg13g2_a21oi_1 _0733_ (.A1(_0229_),
    .A2(_0231_),
    .Y(_0232_),
    .B1(_0187_));
 sg13g2_o21ai_1 _0734_ (.B1(_0184_),
    .Y(_0233_),
    .A1(_0177_),
    .A2(_0185_));
 sg13g2_o21ai_1 _0735_ (.B1(_0180_),
    .Y(_0234_),
    .A1(_0179_),
    .A2(_0182_));
 sg13g2_nand2_1 _0736_ (.Y(_0235_),
    .A(net98),
    .B(net11));
 sg13g2_and3_1 _0737_ (.X(_0236_),
    .A(\system_inst.neuron.v_mem[6] ),
    .B(net96),
    .C(net10));
 sg13g2_nand3_1 _0738_ (.B(net96),
    .C(net10),
    .A(\system_inst.neuron.v_mem[6] ),
    .Y(_0237_));
 sg13g2_a21oi_1 _0739_ (.A1(net96),
    .A2(net10),
    .Y(_0238_),
    .B1(\system_inst.neuron.v_mem[6] ));
 sg13g2_nor2_1 _0740_ (.A(_0236_),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_xnor2_1 _0741_ (.Y(_0240_),
    .A(_0235_),
    .B(_0239_));
 sg13g2_nand2_1 _0742_ (.Y(_0241_),
    .A(_0234_),
    .B(_0240_));
 sg13g2_xnor2_1 _0743_ (.Y(_0242_),
    .A(_0234_),
    .B(_0240_));
 sg13g2_nand2b_1 _0744_ (.Y(_0243_),
    .B(_0233_),
    .A_N(_0242_));
 sg13g2_xor2_1 _0745_ (.B(_0242_),
    .A(_0233_),
    .X(_0244_));
 sg13g2_xnor2_1 _0746_ (.Y(_0245_),
    .A(_0232_),
    .B(_0244_));
 sg13g2_nand2b_1 _0747_ (.Y(_0246_),
    .B(_0074_),
    .A_N(_0245_));
 sg13g2_xnor2_1 _0748_ (.Y(_0247_),
    .A(\system_inst.leak_rate[6] ),
    .B(_0245_));
 sg13g2_xnor2_1 _0749_ (.Y(_0248_),
    .A(_0229_),
    .B(_0231_));
 sg13g2_nand2b_1 _0750_ (.Y(_0249_),
    .B(_0075_),
    .A_N(_0248_));
 sg13g2_inv_1 _0751_ (.Y(_0250_),
    .A(_0249_));
 sg13g2_xor2_1 _0752_ (.B(_0228_),
    .A(_0227_),
    .X(_0251_));
 sg13g2_nand2_1 _0753_ (.Y(_0252_),
    .A(_0076_),
    .B(_0251_));
 sg13g2_xnor2_1 _0754_ (.Y(_0253_),
    .A(_0076_),
    .B(_0251_));
 sg13g2_xor2_1 _0755_ (.B(_0226_),
    .A(_0224_),
    .X(_0254_));
 sg13g2_and2_1 _0756_ (.A(_0077_),
    .B(_0254_),
    .X(_0255_));
 sg13g2_and3_1 _0757_ (.X(_0256_),
    .A(_0216_),
    .B(_0217_),
    .C(_0222_));
 sg13g2_o21ai_1 _0758_ (.B1(_0215_),
    .Y(_0257_),
    .A1(_0223_),
    .A2(_0256_));
 sg13g2_and2_1 _0759_ (.A(_0218_),
    .B(_0257_),
    .X(_0258_));
 sg13g2_nand3_1 _0760_ (.B(_0218_),
    .C(_0257_),
    .A(_0078_),
    .Y(_0259_));
 sg13g2_a21oi_1 _0761_ (.A1(_0218_),
    .A2(_0257_),
    .Y(_0260_),
    .B1(_0078_));
 sg13g2_xnor2_1 _0762_ (.Y(_0261_),
    .A(_0078_),
    .B(_0258_));
 sg13g2_xnor2_1 _0763_ (.Y(_0262_),
    .A(_0219_),
    .B(_0221_));
 sg13g2_nor2_1 _0764_ (.A(\system_inst.leak_rate[1] ),
    .B(_0262_),
    .Y(_0263_));
 sg13g2_xor2_1 _0765_ (.B(_0220_),
    .A(_0006_),
    .X(_0264_));
 sg13g2_nand2b_1 _0766_ (.Y(_0265_),
    .B(\system_inst.leak_rate[0] ),
    .A_N(_0264_));
 sg13g2_xor2_1 _0767_ (.B(_0262_),
    .A(\system_inst.leak_rate[1] ),
    .X(_0266_));
 sg13g2_a21oi_1 _0768_ (.A1(_0265_),
    .A2(_0266_),
    .Y(_0267_),
    .B1(_0263_));
 sg13g2_o21ai_1 _0769_ (.B1(_0259_),
    .Y(_0268_),
    .A1(_0260_),
    .A2(_0267_));
 sg13g2_xnor2_1 _0770_ (.Y(_0269_),
    .A(\system_inst.leak_rate[3] ),
    .B(_0254_));
 sg13g2_a21oi_1 _0771_ (.A1(_0268_),
    .A2(_0269_),
    .Y(_0270_),
    .B1(_0255_));
 sg13g2_o21ai_1 _0772_ (.B1(_0252_),
    .Y(_0271_),
    .A1(_0253_),
    .A2(_0270_));
 sg13g2_xnor2_1 _0773_ (.Y(_0272_),
    .A(_0075_),
    .B(_0248_));
 sg13g2_a21oi_1 _0774_ (.A1(_0271_),
    .A2(_0272_),
    .Y(_0273_),
    .B1(_0250_));
 sg13g2_o21ai_1 _0775_ (.B1(_0246_),
    .Y(_0274_),
    .A1(_0247_),
    .A2(_0273_));
 sg13g2_o21ai_1 _0776_ (.B1(_0243_),
    .Y(_0275_),
    .A1(_0232_),
    .A2(_0244_));
 sg13g2_o21ai_1 _0777_ (.B1(_0237_),
    .Y(_0276_),
    .A1(_0235_),
    .A2(_0238_));
 sg13g2_nand3_1 _0778_ (.B(net96),
    .C(net11),
    .A(\system_inst.neuron.v_mem[7] ),
    .Y(_0277_));
 sg13g2_a21o_1 _0779_ (.A2(net11),
    .A1(net96),
    .B1(\system_inst.neuron.v_mem[7] ),
    .X(_0278_));
 sg13g2_and2_1 _0780_ (.A(_0277_),
    .B(_0278_),
    .X(_0279_));
 sg13g2_nand2_1 _0781_ (.Y(_0280_),
    .A(_0276_),
    .B(_0279_));
 sg13g2_xnor2_1 _0782_ (.Y(_0281_),
    .A(_0276_),
    .B(_0279_));
 sg13g2_nor2_1 _0783_ (.A(_0241_),
    .B(_0281_),
    .Y(_0282_));
 sg13g2_xor2_1 _0784_ (.B(_0281_),
    .A(_0241_),
    .X(_0283_));
 sg13g2_xnor2_1 _0785_ (.Y(_0284_),
    .A(_0275_),
    .B(_0283_));
 sg13g2_xnor2_1 _0786_ (.Y(_0285_),
    .A(_0073_),
    .B(_0284_));
 sg13g2_nor2b_1 _0787_ (.A(\system_inst.leak_cycles[1] ),
    .B_N(\system_inst.neuron.leak_counter[1] ),
    .Y(_0286_));
 sg13g2_nor3_1 _0788_ (.A(\system_inst.neuron.leak_counter[0] ),
    .B(_0064_),
    .C(_0286_),
    .Y(_0287_));
 sg13g2_nand2b_1 _0789_ (.Y(_0288_),
    .B(\system_inst.leak_cycles[1] ),
    .A_N(\system_inst.neuron.leak_counter[1] ));
 sg13g2_o21ai_1 _0790_ (.B1(_0288_),
    .Y(_0289_),
    .A1(\system_inst.neuron.leak_counter[2] ),
    .A2(_0063_));
 sg13g2_a22oi_1 _0791_ (.Y(_0290_),
    .B1(_0063_),
    .B2(\system_inst.neuron.leak_counter[2] ),
    .A2(_0062_),
    .A1(\system_inst.neuron.leak_counter[3] ));
 sg13g2_o21ai_1 _0792_ (.B1(_0290_),
    .Y(_0291_),
    .A1(_0287_),
    .A2(_0289_));
 sg13g2_o21ai_1 _0793_ (.B1(_0291_),
    .Y(_0292_),
    .A1(\system_inst.neuron.leak_counter[3] ),
    .A2(_0062_));
 sg13g2_inv_2 _0794_ (.Y(_0293_),
    .A(net87));
 sg13g2_o21ai_1 _0795_ (.B1(_0293_),
    .Y(_0294_),
    .A1(\system_inst.leak_rate[7] ),
    .A2(_0284_));
 sg13g2_a21oi_2 _0796_ (.B1(_0294_),
    .Y(_0295_),
    .A2(_0285_),
    .A1(_0274_));
 sg13g2_a21oi_1 _0797_ (.A1(_0275_),
    .A2(_0283_),
    .Y(_0296_),
    .B1(_0282_));
 sg13g2_xnor2_1 _0798_ (.Y(_0297_),
    .A(net95),
    .B(_0277_));
 sg13g2_xnor2_1 _0799_ (.Y(_0298_),
    .A(_0280_),
    .B(_0297_));
 sg13g2_xor2_1 _0800_ (.B(_0298_),
    .A(_0296_),
    .X(_0299_));
 sg13g2_xor2_1 _0801_ (.B(_0299_),
    .A(_0295_),
    .X(_0300_));
 sg13g2_xnor2_1 _0802_ (.Y(_0301_),
    .A(_0295_),
    .B(_0299_));
 sg13g2_xnor2_1 _0803_ (.Y(_0302_),
    .A(_0247_),
    .B(_0273_));
 sg13g2_nand2_1 _0804_ (.Y(_0303_),
    .A(_0293_),
    .B(_0302_));
 sg13g2_nand2_1 _0805_ (.Y(_0304_),
    .A(_0245_),
    .B(net87));
 sg13g2_nand3_1 _0806_ (.B(_0303_),
    .C(_0304_),
    .A(net85),
    .Y(_0305_));
 sg13g2_nand2_1 _0807_ (.Y(_0306_),
    .A(\system_inst.loader.threshold[6] ),
    .B(_0305_));
 sg13g2_xor2_1 _0808_ (.B(_0285_),
    .A(_0274_),
    .X(_0307_));
 sg13g2_nand2_1 _0809_ (.Y(_0308_),
    .A(_0284_),
    .B(net87));
 sg13g2_o21ai_1 _0810_ (.B1(_0308_),
    .Y(_0309_),
    .A1(net87),
    .A2(_0307_));
 sg13g2_o21ai_1 _0811_ (.B1(\system_inst.loader.threshold[7] ),
    .Y(_0310_),
    .A1(net83),
    .A2(_0309_));
 sg13g2_xor2_1 _0812_ (.B(_0272_),
    .A(_0271_),
    .X(_0311_));
 sg13g2_nand2_1 _0813_ (.Y(_0312_),
    .A(_0248_),
    .B(net87));
 sg13g2_o21ai_1 _0814_ (.B1(_0312_),
    .Y(_0313_),
    .A1(net87),
    .A2(_0311_));
 sg13g2_or2_1 _0815_ (.X(_0314_),
    .B(_0313_),
    .A(net83));
 sg13g2_nor3_2 _0816_ (.A(\system_inst.loader.threshold[7] ),
    .B(net83),
    .C(_0309_),
    .Y(_0315_));
 sg13g2_xnor2_1 _0817_ (.Y(_0316_),
    .A(\system_inst.loader.threshold[6] ),
    .B(_0305_));
 sg13g2_o21ai_1 _0818_ (.B1(_0310_),
    .Y(_0317_),
    .A1(\system_inst.loader.threshold[5] ),
    .A2(_0314_));
 sg13g2_nor3_1 _0819_ (.A(_0315_),
    .B(_0316_),
    .C(_0317_),
    .Y(_0318_));
 sg13g2_o21ai_1 _0820_ (.B1(\system_inst.loader.threshold[5] ),
    .Y(_0319_),
    .A1(net83),
    .A2(_0313_));
 sg13g2_xnor2_1 _0821_ (.Y(_0320_),
    .A(_0253_),
    .B(_0270_));
 sg13g2_nor2_1 _0822_ (.A(_0251_),
    .B(_0293_),
    .Y(_0321_));
 sg13g2_a21oi_1 _0823_ (.A1(_0293_),
    .A2(_0320_),
    .Y(_0322_),
    .B1(_0321_));
 sg13g2_inv_1 _0824_ (.Y(_0323_),
    .A(_0322_));
 sg13g2_o21ai_1 _0825_ (.B1(\system_inst.loader.threshold[4] ),
    .Y(_0324_),
    .A1(net83),
    .A2(_0323_));
 sg13g2_nand2_1 _0826_ (.Y(_0325_),
    .A(_0319_),
    .B(_0324_));
 sg13g2_nand3_1 _0827_ (.B(net85),
    .C(_0322_),
    .A(_0068_),
    .Y(_0326_));
 sg13g2_nand3_1 _0828_ (.B(_0324_),
    .C(_0326_),
    .A(_0319_),
    .Y(_0327_));
 sg13g2_nor4_2 _0829_ (.A(_0315_),
    .B(_0316_),
    .C(_0317_),
    .Y(_0328_),
    .D(_0327_));
 sg13g2_xnor2_1 _0830_ (.Y(_0329_),
    .A(_0268_),
    .B(_0269_));
 sg13g2_nor2_1 _0831_ (.A(_0254_),
    .B(_0293_),
    .Y(_0330_));
 sg13g2_a21oi_1 _0832_ (.A1(_0293_),
    .A2(_0329_),
    .Y(_0331_),
    .B1(_0330_));
 sg13g2_inv_1 _0833_ (.Y(_0332_),
    .A(_0331_));
 sg13g2_a21oi_1 _0834_ (.A1(_0300_),
    .A2(_0331_),
    .Y(_0333_),
    .B1(_0069_));
 sg13g2_xnor2_1 _0835_ (.Y(_0334_),
    .A(_0261_),
    .B(_0267_));
 sg13g2_nand2_1 _0836_ (.Y(_0335_),
    .A(_0258_),
    .B(net87));
 sg13g2_o21ai_1 _0837_ (.B1(_0335_),
    .Y(_0336_),
    .A1(net88),
    .A2(_0334_));
 sg13g2_inv_1 _0838_ (.Y(_0337_),
    .A(_0336_));
 sg13g2_a21oi_1 _0839_ (.A1(net85),
    .A2(_0336_),
    .Y(_0338_),
    .B1(_0070_));
 sg13g2_nor3_1 _0840_ (.A(\system_inst.loader.threshold[2] ),
    .B(net84),
    .C(_0337_),
    .Y(_0339_));
 sg13g2_nor3_1 _0841_ (.A(\system_inst.loader.threshold[3] ),
    .B(net84),
    .C(_0332_),
    .Y(_0340_));
 sg13g2_nand3_1 _0842_ (.B(net85),
    .C(_0331_),
    .A(_0069_),
    .Y(_0341_));
 sg13g2_or4_1 _0843_ (.A(_0333_),
    .B(_0338_),
    .C(_0339_),
    .D(_0340_),
    .X(_0342_));
 sg13g2_nand2b_1 _0844_ (.Y(_0343_),
    .B(net88),
    .A_N(_0262_));
 sg13g2_xnor2_1 _0845_ (.Y(_0344_),
    .A(_0265_),
    .B(_0266_));
 sg13g2_o21ai_1 _0846_ (.B1(_0343_),
    .Y(_0345_),
    .A1(net87),
    .A2(_0344_));
 sg13g2_nand2_1 _0847_ (.Y(_0346_),
    .A(net85),
    .B(_0345_));
 sg13g2_a21oi_1 _0848_ (.A1(net85),
    .A2(_0345_),
    .Y(_0347_),
    .B1(_0071_));
 sg13g2_nand3_1 _0849_ (.B(net85),
    .C(_0345_),
    .A(_0071_),
    .Y(_0348_));
 sg13g2_nor2_1 _0850_ (.A(_0079_),
    .B(net88),
    .Y(_0349_));
 sg13g2_xnor2_1 _0851_ (.Y(_0350_),
    .A(_0264_),
    .B(_0349_));
 sg13g2_or2_1 _0852_ (.X(_0351_),
    .B(_0350_),
    .A(net84));
 sg13g2_nand3b_1 _0853_ (.B(_0072_),
    .C(net85),
    .Y(_0352_),
    .A_N(_0350_));
 sg13g2_nand2_1 _0854_ (.Y(_0353_),
    .A(_0348_),
    .B(_0352_));
 sg13g2_a21oi_1 _0855_ (.A1(_0348_),
    .A2(_0352_),
    .Y(_0354_),
    .B1(_0347_));
 sg13g2_o21ai_1 _0856_ (.B1(_0341_),
    .Y(_0355_),
    .A1(_0333_),
    .A2(_0338_));
 sg13g2_o21ai_1 _0857_ (.B1(_0355_),
    .Y(_0356_),
    .A1(_0342_),
    .A2(_0354_));
 sg13g2_o21ai_1 _0858_ (.B1(_0310_),
    .Y(_0357_),
    .A1(_0306_),
    .A2(_0315_));
 sg13g2_a221oi_1 _0859_ (.B2(_0356_),
    .C1(_0357_),
    .B1(_0328_),
    .A1(_0318_),
    .Y(_0358_),
    .A2(_0325_));
 sg13g2_nand2_1 _0860_ (.Y(_0359_),
    .A(\system_inst.loader.threshold[0] ),
    .B(_0351_));
 sg13g2_nor3_1 _0861_ (.A(_0342_),
    .B(_0347_),
    .C(_0353_),
    .Y(_0360_));
 sg13g2_and3_1 _0862_ (.X(_0361_),
    .A(_0328_),
    .B(_0359_),
    .C(_0360_));
 sg13g2_nor2_1 _0863_ (.A(_0358_),
    .B(_0361_),
    .Y(_0362_));
 sg13g2_or2_1 _0864_ (.X(_0363_),
    .B(_0361_),
    .A(_0358_));
 sg13g2_or3_1 _0865_ (.A(net193),
    .B(\system_inst.neuron.refr_cnt[1] ),
    .C(\system_inst.neuron.refr_cnt[0] ),
    .X(_0364_));
 sg13g2_or2_2 _0866_ (.X(_0365_),
    .B(_0364_),
    .A(net111));
 sg13g2_and2_2 _0867_ (.A(params_ready),
    .B(net1),
    .X(_0366_));
 sg13g2_nand2_2 _0868_ (.Y(_0367_),
    .A(params_ready),
    .B(net1));
 sg13g2_and2_1 _0869_ (.A(net3),
    .B(_0366_),
    .X(_0368_));
 sg13g2_nand2b_2 _0870_ (.Y(_0369_),
    .B(_0368_),
    .A_N(_0365_));
 sg13g2_nor3_1 _0871_ (.A(net100),
    .B(net82),
    .C(net90),
    .Y(_0042_));
 sg13g2_nor2_1 _0872_ (.A(_0351_),
    .B(_0369_),
    .Y(_0370_));
 sg13g2_a22oi_1 _0873_ (.Y(_0371_),
    .B1(_0370_),
    .B2(_0362_),
    .A2(_0369_),
    .A1(net120));
 sg13g2_nor2_1 _0874_ (.A(net101),
    .B(_0371_),
    .Y(_0043_));
 sg13g2_nor2_1 _0875_ (.A(_0346_),
    .B(net90),
    .Y(_0372_));
 sg13g2_a22oi_1 _0876_ (.Y(_0373_),
    .B1(_0372_),
    .B2(net82),
    .A2(net90),
    .A1(net147));
 sg13g2_nor2_1 _0877_ (.A(net100),
    .B(_0373_),
    .Y(_0044_));
 sg13g2_nor3_1 _0878_ (.A(net84),
    .B(_0337_),
    .C(net90),
    .Y(_0374_));
 sg13g2_a22oi_1 _0879_ (.Y(_0375_),
    .B1(_0374_),
    .B2(net82),
    .A2(_0369_),
    .A1(net177));
 sg13g2_nor2_1 _0880_ (.A(net100),
    .B(_0375_),
    .Y(_0045_));
 sg13g2_nor3_1 _0881_ (.A(net83),
    .B(_0332_),
    .C(net90),
    .Y(_0376_));
 sg13g2_a22oi_1 _0882_ (.Y(_0377_),
    .B1(_0376_),
    .B2(net82),
    .A2(net89),
    .A1(net158));
 sg13g2_nor2_1 _0883_ (.A(net100),
    .B(_0377_),
    .Y(_0046_));
 sg13g2_nor3_1 _0884_ (.A(net83),
    .B(_0323_),
    .C(net89),
    .Y(_0378_));
 sg13g2_a22oi_1 _0885_ (.Y(_0379_),
    .B1(_0378_),
    .B2(net82),
    .A2(net90),
    .A1(net159));
 sg13g2_nor2_1 _0886_ (.A(net100),
    .B(_0379_),
    .Y(_0047_));
 sg13g2_nor2_1 _0887_ (.A(_0314_),
    .B(net89),
    .Y(_0380_));
 sg13g2_a22oi_1 _0888_ (.Y(_0381_),
    .B1(_0380_),
    .B2(net82),
    .A2(net89),
    .A1(net144));
 sg13g2_nor2_1 _0889_ (.A(net100),
    .B(_0381_),
    .Y(_0048_));
 sg13g2_nor2_1 _0890_ (.A(_0305_),
    .B(net89),
    .Y(_0382_));
 sg13g2_a22oi_1 _0891_ (.Y(_0383_),
    .B1(_0382_),
    .B2(net82),
    .A2(net89),
    .A1(net164));
 sg13g2_nor2_1 _0892_ (.A(net100),
    .B(_0383_),
    .Y(_0049_));
 sg13g2_nor3_1 _0893_ (.A(net83),
    .B(_0309_),
    .C(net89),
    .Y(_0384_));
 sg13g2_a22oi_1 _0894_ (.Y(_0385_),
    .B1(_0384_),
    .B2(net82),
    .A2(net89),
    .A1(net135));
 sg13g2_nor2_1 _0895_ (.A(net100),
    .B(_0385_),
    .Y(_0050_));
 sg13g2_and3_1 _0896_ (.X(_0051_),
    .A(net95),
    .B(net2),
    .C(net90));
 sg13g2_nand2_1 _0897_ (.Y(_0386_),
    .A(_0365_),
    .B(_0366_));
 sg13g2_o21ai_1 _0898_ (.B1(_0368_),
    .Y(_0387_),
    .A1(_0358_),
    .A2(_0361_));
 sg13g2_and3_1 _0899_ (.X(_0388_),
    .A(_0060_),
    .B(_0386_),
    .C(_0387_));
 sg13g2_a22oi_1 _0900_ (.Y(_0389_),
    .B1(_0386_),
    .B2(_0387_),
    .A2(_0365_),
    .A1(_0060_));
 sg13g2_nor3_1 _0901_ (.A(net103),
    .B(_0388_),
    .C(_0389_),
    .Y(_0052_));
 sg13g2_xnor2_1 _0902_ (.Y(_0390_),
    .A(net196),
    .B(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_a22oi_1 _0903_ (.Y(_0391_),
    .B1(_0390_),
    .B2(_0365_),
    .A2(_0387_),
    .A1(_0386_));
 sg13g2_a221oi_1 _0904_ (.B2(_0363_),
    .C1(net196),
    .B1(_0368_),
    .A1(_0365_),
    .Y(_0392_),
    .A2(_0366_));
 sg13g2_nor3_1 _0905_ (.A(net103),
    .B(_0391_),
    .C(_0392_),
    .Y(_0053_));
 sg13g2_a221oi_1 _0906_ (.B2(_0363_),
    .C1(net193),
    .B1(_0368_),
    .A1(_0365_),
    .Y(_0393_),
    .A2(_0366_));
 sg13g2_o21ai_1 _0907_ (.B1(net193),
    .Y(_0394_),
    .A1(\system_inst.neuron.refr_cnt[1] ),
    .A2(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_and3_1 _0908_ (.X(_0395_),
    .A(_0364_),
    .B(_0366_),
    .C(_0394_));
 sg13g2_nor3_1 _0909_ (.A(net102),
    .B(_0393_),
    .C(_0395_),
    .Y(_0054_));
 sg13g2_o21ai_1 _0910_ (.B1(net111),
    .Y(_0396_),
    .A1(_0364_),
    .A2(_0367_));
 sg13g2_nor2_1 _0911_ (.A(net102),
    .B(net112),
    .Y(_0055_));
 sg13g2_o21ai_1 _0912_ (.B1(net108),
    .Y(_0397_),
    .A1(net88),
    .A2(_0367_));
 sg13g2_xnor2_1 _0913_ (.Y(_0398_),
    .A(net185),
    .B(_0366_));
 sg13g2_nor2_1 _0914_ (.A(_0397_),
    .B(net186),
    .Y(_0056_));
 sg13g2_and3_1 _0915_ (.X(_0399_),
    .A(net124),
    .B(\system_inst.neuron.leak_counter[0] ),
    .C(_0366_));
 sg13g2_a21oi_1 _0916_ (.A1(\system_inst.neuron.leak_counter[0] ),
    .A2(_0366_),
    .Y(_0400_),
    .B1(net124));
 sg13g2_nor3_1 _0917_ (.A(_0397_),
    .B(_0399_),
    .C(net125),
    .Y(_0057_));
 sg13g2_nand2_1 _0918_ (.Y(_0401_),
    .A(\system_inst.neuron.leak_counter[2] ),
    .B(_0399_));
 sg13g2_xnor2_1 _0919_ (.Y(_0402_),
    .A(net181),
    .B(_0399_));
 sg13g2_nor2_1 _0920_ (.A(_0397_),
    .B(net182),
    .Y(_0058_));
 sg13g2_xor2_1 _0921_ (.B(_0401_),
    .A(net175),
    .X(_0403_));
 sg13g2_nor2_1 _0922_ (.A(_0397_),
    .B(net176),
    .Y(_0059_));
 sg13g2_dfrbp_1 _0923_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net60),
    .D(net188),
    .Q_N(_0454_),
    .Q(params_ready));
 sg13g2_dfrbp_1 _0924_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net67),
    .D(_0009_),
    .Q_N(_0453_),
    .Q(\system_inst.loader.weight_a[0] ));
 sg13g2_dfrbp_1 _0925_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net65),
    .D(_0010_),
    .Q_N(_0452_),
    .Q(\system_inst.loader.weight_a[1] ));
 sg13g2_dfrbp_1 _0926_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net58),
    .D(net116),
    .Q_N(_0451_),
    .Q(\system_inst.loader.weight_a[2] ));
 sg13g2_dfrbp_1 _0927_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net56),
    .D(_0012_),
    .Q_N(_0450_),
    .Q(\system_inst.leak_rate[0] ));
 sg13g2_dfrbp_1 _0928_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net54),
    .D(_0013_),
    .Q_N(_0449_),
    .Q(\system_inst.leak_rate[1] ));
 sg13g2_dfrbp_1 _0929_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net52),
    .D(net184),
    .Q_N(_0448_),
    .Q(\system_inst.leak_rate[2] ));
 sg13g2_dfrbp_1 _0930_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net50),
    .D(net161),
    .Q_N(_0447_),
    .Q(\system_inst.leak_rate[3] ));
 sg13g2_dfrbp_1 _0931_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net48),
    .D(net166),
    .Q_N(_0446_),
    .Q(\system_inst.leak_rate[4] ));
 sg13g2_dfrbp_1 _0932_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net46),
    .D(net168),
    .Q_N(_0445_),
    .Q(\system_inst.leak_rate[5] ));
 sg13g2_dfrbp_1 _0933_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net44),
    .D(net134),
    .Q_N(_0444_),
    .Q(\system_inst.leak_rate[6] ));
 sg13g2_dfrbp_1 _0934_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net42),
    .D(net155),
    .Q_N(_0443_),
    .Q(\system_inst.leak_rate[7] ));
 sg13g2_dfrbp_1 _0935_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net40),
    .D(net137),
    .Q_N(_0442_),
    .Q(\system_inst.loader.threshold[0] ));
 sg13g2_dfrbp_1 _0936_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net38),
    .D(net141),
    .Q_N(_0441_),
    .Q(\system_inst.loader.threshold[1] ));
 sg13g2_dfrbp_1 _0937_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net36),
    .D(net143),
    .Q_N(_0440_),
    .Q(\system_inst.loader.threshold[2] ));
 sg13g2_dfrbp_1 _0938_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net34),
    .D(net180),
    .Q_N(_0439_),
    .Q(\system_inst.loader.threshold[3] ));
 sg13g2_dfrbp_1 _0939_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net32),
    .D(net157),
    .Q_N(_0438_),
    .Q(\system_inst.loader.threshold[4] ));
 sg13g2_dfrbp_1 _0940_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net30),
    .D(net130),
    .Q_N(_0437_),
    .Q(\system_inst.loader.threshold[5] ));
 sg13g2_dfrbp_1 _0941_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net28),
    .D(net139),
    .Q_N(_0436_),
    .Q(\system_inst.loader.threshold[6] ));
 sg13g2_dfrbp_1 _0942_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net26),
    .D(net151),
    .Q_N(_0435_),
    .Q(\system_inst.loader.threshold[7] ));
 sg13g2_dfrbp_1 _0943_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net81),
    .D(net118),
    .Q_N(_0434_),
    .Q(\system_inst.leak_cycles[0] ));
 sg13g2_dfrbp_1 _0944_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net79),
    .D(_0029_),
    .Q_N(_0433_),
    .Q(\system_inst.leak_cycles[1] ));
 sg13g2_dfrbp_1 _0945_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net77),
    .D(net146),
    .Q_N(_0432_),
    .Q(\system_inst.leak_cycles[2] ));
 sg13g2_dfrbp_1 _0946_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net75),
    .D(net149),
    .Q_N(_0431_),
    .Q(\system_inst.leak_cycles[3] ));
 sg13g2_dfrbp_1 _0947_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net73),
    .D(_0032_),
    .Q_N(_0430_),
    .Q(\system_inst.loader.shift_reg[0] ));
 sg13g2_dfrbp_1 _0948_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net71),
    .D(net163),
    .Q_N(_0429_),
    .Q(\system_inst.loader.shift_reg[1] ));
 sg13g2_dfrbp_1 _0949_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net69),
    .D(_0034_),
    .Q_N(_0428_),
    .Q(\system_inst.loader.shift_reg[2] ));
 sg13g2_dfrbp_1 _0950_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net66),
    .D(_0035_),
    .Q_N(_0427_),
    .Q(\system_inst.loader.shift_reg[3] ));
 sg13g2_dfrbp_1 _0951_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net57),
    .D(_0036_),
    .Q_N(_0426_),
    .Q(\system_inst.loader.shift_reg[4] ));
 sg13g2_dfrbp_1 _0952_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net53),
    .D(_0037_),
    .Q_N(_0425_),
    .Q(\system_inst.loader.shift_reg[5] ));
 sg13g2_dfrbp_1 _0953_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net49),
    .D(net170),
    .Q_N(_0424_),
    .Q(\system_inst.loader.shift_reg[6] ));
 sg13g2_dfrbp_1 _0954_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net45),
    .D(_0039_),
    .Q_N(_0423_),
    .Q(\system_inst.loader.bit_count[0] ));
 sg13g2_dfrbp_1 _0955_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net41),
    .D(_0040_),
    .Q_N(_0422_),
    .Q(\system_inst.loader.bit_count[1] ));
 sg13g2_dfrbp_1 _0956_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net61),
    .D(_0041_),
    .Q_N(_0005_),
    .Q(\system_inst.loader.bit_count[2] ));
 sg13g2_dfrbp_1 _0957_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net62),
    .D(_0000_),
    .Q_N(_0455_),
    .Q(\system_inst.loader.current_state[0] ));
 sg13g2_dfrbp_1 _0958_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net63),
    .D(_0001_),
    .Q_N(_0007_),
    .Q(\system_inst.loader.current_state[1] ));
 sg13g2_dfrbp_1 _0959_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net64),
    .D(_0002_),
    .Q_N(_0456_),
    .Q(\system_inst.loader.current_state[2] ));
 sg13g2_dfrbp_1 _0960_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net109),
    .D(net123),
    .Q_N(_0457_),
    .Q(\system_inst.loader.current_state[3] ));
 sg13g2_dfrbp_1 _0961_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net37),
    .D(_0004_),
    .Q_N(_0421_),
    .Q(\system_inst.loader.current_state[5] ));
 sg13g2_dfrbp_1 _0962_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net33),
    .D(_0042_),
    .Q_N(_0420_),
    .Q(spike_out));
 sg13g2_dfrbp_1 _0963_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net31),
    .D(_0043_),
    .Q_N(_0006_),
    .Q(\system_inst.neuron.v_mem[0] ));
 sg13g2_dfrbp_1 _0964_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net27),
    .D(_0044_),
    .Q_N(_0419_),
    .Q(\system_inst.neuron.v_mem[1] ));
 sg13g2_dfrbp_1 _0965_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net80),
    .D(_0045_),
    .Q_N(_0418_),
    .Q(\system_inst.neuron.v_mem[2] ));
 sg13g2_dfrbp_1 _0966_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net76),
    .D(_0046_),
    .Q_N(_0417_),
    .Q(\system_inst.neuron.v_mem[3] ));
 sg13g2_dfrbp_1 _0967_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net72),
    .D(_0047_),
    .Q_N(_0416_),
    .Q(\system_inst.neuron.v_mem[4] ));
 sg13g2_dfrbp_1 _0968_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net68),
    .D(_0048_),
    .Q_N(_0415_),
    .Q(\system_inst.neuron.v_mem[5] ));
 sg13g2_dfrbp_1 _0969_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net55),
    .D(_0049_),
    .Q_N(_0414_),
    .Q(\system_inst.neuron.v_mem[6] ));
 sg13g2_dfrbp_1 _0970_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net47),
    .D(_0050_),
    .Q_N(_0413_),
    .Q(\system_inst.neuron.v_mem[7] ));
 sg13g2_dfrbp_1 _0971_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net39),
    .D(_0051_),
    .Q_N(_0412_),
    .Q(\system_inst.neuron.v_mem[8] ));
 sg13g2_dfrbp_1 _0972_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net29),
    .D(_0052_),
    .Q_N(_0411_),
    .Q(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_dfrbp_1 _0973_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net78),
    .D(net197),
    .Q_N(_0410_),
    .Q(\system_inst.neuron.refr_cnt[1] ));
 sg13g2_dfrbp_1 _0974_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net70),
    .D(net194),
    .Q_N(_0409_),
    .Q(\system_inst.neuron.refr_cnt[2] ));
 sg13g2_dfrbp_1 _0975_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net51),
    .D(_0055_),
    .Q_N(_0408_),
    .Q(\system_inst.neuron.refr_cnt[3] ));
 sg13g2_dfrbp_1 _0976_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net35),
    .D(_0056_),
    .Q_N(_0407_),
    .Q(\system_inst.neuron.leak_counter[0] ));
 sg13g2_dfrbp_1 _0977_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net74),
    .D(net126),
    .Q_N(_0406_),
    .Q(\system_inst.neuron.leak_counter[1] ));
 sg13g2_dfrbp_1 _0978_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net43),
    .D(_0058_),
    .Q_N(_0405_),
    .Q(\system_inst.neuron.leak_counter[2] ));
 sg13g2_dfrbp_1 _0979_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net59),
    .D(_0059_),
    .Q_N(_0404_),
    .Q(\system_inst.neuron.leak_counter[3] ));
 sg13g2_tiehi _0964__27 (.L_HI(net27));
 sg13g2_tiehi _0941__28 (.L_HI(net28));
 sg13g2_tiehi _0972__29 (.L_HI(net29));
 sg13g2_tiehi _0940__30 (.L_HI(net30));
 sg13g2_tiehi _0963__31 (.L_HI(net31));
 sg13g2_tiehi _0939__32 (.L_HI(net32));
 sg13g2_tiehi _0962__33 (.L_HI(net33));
 sg13g2_tiehi _0938__34 (.L_HI(net34));
 sg13g2_tiehi _0976__35 (.L_HI(net35));
 sg13g2_tiehi _0937__36 (.L_HI(net36));
 sg13g2_tiehi _0961__37 (.L_HI(net37));
 sg13g2_tiehi _0936__38 (.L_HI(net38));
 sg13g2_tiehi _0971__39 (.L_HI(net39));
 sg13g2_tiehi _0935__40 (.L_HI(net40));
 sg13g2_tiehi _0955__41 (.L_HI(net41));
 sg13g2_tiehi _0934__42 (.L_HI(net42));
 sg13g2_tiehi _0978__43 (.L_HI(net43));
 sg13g2_tiehi _0933__44 (.L_HI(net44));
 sg13g2_tiehi _0954__45 (.L_HI(net45));
 sg13g2_tiehi _0932__46 (.L_HI(net46));
 sg13g2_tiehi _0970__47 (.L_HI(net47));
 sg13g2_tiehi _0931__48 (.L_HI(net48));
 sg13g2_tiehi _0953__49 (.L_HI(net49));
 sg13g2_tiehi _0930__50 (.L_HI(net50));
 sg13g2_tiehi _0975__51 (.L_HI(net51));
 sg13g2_tiehi _0929__52 (.L_HI(net52));
 sg13g2_tiehi _0952__53 (.L_HI(net53));
 sg13g2_tiehi _0928__54 (.L_HI(net54));
 sg13g2_tiehi _0969__55 (.L_HI(net55));
 sg13g2_tiehi _0927__56 (.L_HI(net56));
 sg13g2_tiehi _0951__57 (.L_HI(net57));
 sg13g2_tiehi _0926__58 (.L_HI(net58));
 sg13g2_tiehi _0979__59 (.L_HI(net59));
 sg13g2_tiehi _0923__60 (.L_HI(net60));
 sg13g2_tiehi _0956__61 (.L_HI(net61));
 sg13g2_tiehi _0957__62 (.L_HI(net62));
 sg13g2_tiehi _0958__63 (.L_HI(net63));
 sg13g2_tiehi _0959__64 (.L_HI(net64));
 sg13g2_tiehi _0925__65 (.L_HI(net65));
 sg13g2_tiehi _0950__66 (.L_HI(net66));
 sg13g2_tiehi _0924__67 (.L_HI(net67));
 sg13g2_tiehi _0968__68 (.L_HI(net68));
 sg13g2_tiehi _0949__69 (.L_HI(net69));
 sg13g2_tiehi _0974__70 (.L_HI(net70));
 sg13g2_tiehi _0948__71 (.L_HI(net71));
 sg13g2_tiehi _0967__72 (.L_HI(net72));
 sg13g2_tiehi _0947__73 (.L_HI(net73));
 sg13g2_tiehi _0977__74 (.L_HI(net74));
 sg13g2_tiehi _0946__75 (.L_HI(net75));
 sg13g2_tiehi _0966__76 (.L_HI(net76));
 sg13g2_tiehi _0945__77 (.L_HI(net77));
 sg13g2_tiehi _0973__78 (.L_HI(net78));
 sg13g2_tiehi _0944__79 (.L_HI(net79));
 sg13g2_tiehi _0965__80 (.L_HI(net80));
 sg13g2_tiehi _0943__81 (.L_HI(net81));
 sg13g2_tiehi _0960__82 (.L_HI(net109));
 sg13g2_tiehi tt_um_wokwi_434925031692840961_83 (.L_HI(net110));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_wokwi_434925031692840961_13 (.L_LO(net13));
 sg13g2_tielo tt_um_wokwi_434925031692840961_14 (.L_LO(net14));
 sg13g2_tielo tt_um_wokwi_434925031692840961_15 (.L_LO(net15));
 sg13g2_tielo tt_um_wokwi_434925031692840961_16 (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_434925031692840961_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_434925031692840961_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_434925031692840961_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_434925031692840961_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_434925031692840961_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_434925031692840961_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_434925031692840961_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_434925031692840961_24 (.L_LO(net24));
 sg13g2_tielo tt_um_wokwi_434925031692840961_25 (.L_LO(net25));
 sg13g2_tiehi _0942__26 (.L_HI(net26));
 sg13g2_buf_2 _1052_ (.A(params_ready),
    .X(uio_out[0]));
 sg13g2_buf_1 _1053_ (.A(spike_out),
    .X(uo_out[0]));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_0362_));
 sg13g2_buf_2 fanout83 (.A(_0301_),
    .X(net83));
 sg13g2_buf_1 fanout84 (.A(_0301_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0300_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0138_),
    .X(net86));
 sg13g2_buf_4 fanout87 (.X(net87),
    .A(_0292_));
 sg13g2_buf_1 fanout88 (.A(_0292_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(net90),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0369_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0095_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0095_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0092_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0087_),
    .X(net94));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(net195));
 sg13g2_buf_2 fanout96 (.A(net97),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(\system_inst.loader.weight_a[2] ),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(net190),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(\system_inst.loader.weight_a[0] ),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(net103),
    .X(net101));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(net103));
 sg13g2_buf_2 fanout103 (.A(_0082_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(net2),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(net107),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(net108),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(net2),
    .X(net108));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_2 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[0]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[1]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[2]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[3]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[4]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[5]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(ui_in[6]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(ui_in[7]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[0]),
    .X(net11));
 sg13g2_tielo tt_um_wokwi_434925031692840961_12 (.L_LO(net12));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\system_inst.neuron.refr_cnt[3] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0396_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold3 (.A(\system_inst.loader.bit_count[2] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0161_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold5 (.A(\system_inst.loader.weight_a[2] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0011_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold7 (.A(\system_inst.leak_cycles[0] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0028_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold9 (.A(\system_inst.loader.bit_count[0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold10 (.A(\system_inst.neuron.v_mem[0] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold11 (.A(\system_inst.leak_rate[0] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold12 (.A(\system_inst.loader.current_state[3] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0003_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold14 (.A(\system_inst.neuron.leak_counter[1] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0400_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0057_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold17 (.A(\system_inst.loader.current_state[0] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold18 (.A(\system_inst.loader.weight_a[0] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold19 (.A(\system_inst.loader.threshold[5] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0025_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold21 (.A(\system_inst.loader.bit_count[1] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0158_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold23 (.A(\system_inst.leak_rate[6] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0018_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold25 (.A(\system_inst.neuron.v_mem[7] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold26 (.A(\system_inst.loader.threshold[0] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0020_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold28 (.A(\system_inst.loader.threshold[6] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0026_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold30 (.A(\system_inst.loader.threshold[1] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0021_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold32 (.A(\system_inst.loader.threshold[2] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0022_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold34 (.A(\system_inst.neuron.v_mem[5] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold35 (.A(\system_inst.leak_cycles[2] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0030_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold37 (.A(\system_inst.neuron.v_mem[1] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold38 (.A(\system_inst.leak_cycles[3] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0031_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold40 (.A(\system_inst.loader.threshold[7] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0027_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold42 (.A(\system_inst.loader.current_state[1] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0093_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold44 (.A(\system_inst.leak_rate[7] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0019_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold46 (.A(\system_inst.loader.threshold[4] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0024_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold48 (.A(\system_inst.neuron.v_mem[3] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold49 (.A(\system_inst.neuron.v_mem[4] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold50 (.A(\system_inst.leak_rate[3] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0015_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold52 (.A(\system_inst.loader.shift_reg[0] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0033_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold54 (.A(\system_inst.neuron.v_mem[6] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold55 (.A(\system_inst.leak_rate[4] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0016_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold57 (.A(\system_inst.leak_rate[5] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0017_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold59 (.A(\system_inst.loader.shift_reg[5] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0038_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold61 (.A(\system_inst.leak_cycles[1] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold62 (.A(\system_inst.loader.current_state[5] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0096_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold64 (.A(\system_inst.loader.current_state[2] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold65 (.A(\system_inst.neuron.leak_counter[3] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0403_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold67 (.A(\system_inst.neuron.v_mem[2] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold68 (.A(\system_inst.loader.shift_reg[4] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold69 (.A(\system_inst.loader.threshold[3] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0023_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold71 (.A(\system_inst.neuron.leak_counter[2] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0402_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold73 (.A(\system_inst.leak_rate[2] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0014_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold75 (.A(\system_inst.neuron.leak_counter[0] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0398_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold77 (.A(params_ready),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0008_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold79 (.A(\system_inst.loader.shift_reg[3] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold80 (.A(\system_inst.loader.weight_a[1] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold81 (.A(\system_inst.leak_rate[1] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold82 (.A(\system_inst.loader.shift_reg[2] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold83 (.A(\system_inst.neuron.refr_cnt[2] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0054_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold85 (.A(\system_inst.neuron.v_mem[8] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold86 (.A(\system_inst.neuron.refr_cnt[1] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0053_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold88 (.A(\system_inst.loader.shift_reg[1] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold89 (.A(\system_inst.neuron.refr_cnt[0] ),
    .X(net199));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_4 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_246 ();
 sg13g2_decap_8 FILLER_17_253 ();
 sg13g2_decap_8 FILLER_17_260 ();
 sg13g2_decap_4 FILLER_17_267 ();
 sg13g2_fill_2 FILLER_17_271 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_fill_1 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_217 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_fill_2 FILLER_18_250 ();
 sg13g2_fill_1 FILLER_18_252 ();
 sg13g2_fill_2 FILLER_18_279 ();
 sg13g2_fill_1 FILLER_18_285 ();
 sg13g2_fill_1 FILLER_18_312 ();
 sg13g2_decap_4 FILLER_18_337 ();
 sg13g2_fill_2 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_fill_1 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_146 ();
 sg13g2_decap_8 FILLER_19_153 ();
 sg13g2_decap_8 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_decap_4 FILLER_19_301 ();
 sg13g2_fill_2 FILLER_19_305 ();
 sg13g2_decap_4 FILLER_19_314 ();
 sg13g2_fill_2 FILLER_19_318 ();
 sg13g2_fill_2 FILLER_19_334 ();
 sg13g2_fill_1 FILLER_19_336 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_fill_1 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_110 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_fill_2 FILLER_20_137 ();
 sg13g2_fill_1 FILLER_20_139 ();
 sg13g2_decap_4 FILLER_20_144 ();
 sg13g2_fill_2 FILLER_20_148 ();
 sg13g2_decap_4 FILLER_20_179 ();
 sg13g2_fill_2 FILLER_20_209 ();
 sg13g2_fill_1 FILLER_20_211 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_decap_4 FILLER_20_283 ();
 sg13g2_fill_1 FILLER_20_287 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_fill_2 FILLER_20_332 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_fill_2 FILLER_20_369 ();
 sg13g2_fill_1 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_4 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_121 ();
 sg13g2_fill_1 FILLER_21_137 ();
 sg13g2_decap_4 FILLER_21_148 ();
 sg13g2_fill_2 FILLER_21_166 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_decap_4 FILLER_21_174 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_212 ();
 sg13g2_decap_4 FILLER_21_221 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_4 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_242 ();
 sg13g2_fill_2 FILLER_21_248 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_fill_2 FILLER_21_277 ();
 sg13g2_fill_2 FILLER_21_289 ();
 sg13g2_decap_8 FILLER_21_314 ();
 sg13g2_decap_8 FILLER_21_321 ();
 sg13g2_fill_2 FILLER_21_328 ();
 sg13g2_fill_2 FILLER_21_342 ();
 sg13g2_fill_1 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_4 FILLER_22_77 ();
 sg13g2_fill_2 FILLER_22_81 ();
 sg13g2_decap_4 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_2 FILLER_22_152 ();
 sg13g2_fill_1 FILLER_22_154 ();
 sg13g2_fill_2 FILLER_22_159 ();
 sg13g2_decap_4 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_1 FILLER_22_194 ();
 sg13g2_fill_1 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_fill_2 FILLER_22_260 ();
 sg13g2_fill_2 FILLER_22_266 ();
 sg13g2_fill_1 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_fill_2 FILLER_22_332 ();
 sg13g2_fill_1 FILLER_22_334 ();
 sg13g2_decap_4 FILLER_22_339 ();
 sg13g2_fill_2 FILLER_22_353 ();
 sg13g2_fill_1 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_4 FILLER_23_84 ();
 sg13g2_fill_2 FILLER_23_88 ();
 sg13g2_decap_4 FILLER_23_107 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_1 FILLER_23_128 ();
 sg13g2_fill_2 FILLER_23_170 ();
 sg13g2_fill_1 FILLER_23_198 ();
 sg13g2_decap_8 FILLER_23_230 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_decap_4 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_254 ();
 sg13g2_decap_8 FILLER_23_261 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_fill_2 FILLER_23_279 ();
 sg13g2_fill_2 FILLER_23_299 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_fill_2 FILLER_23_341 ();
 sg13g2_fill_2 FILLER_23_369 ();
 sg13g2_fill_2 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_fill_1 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_fill_2 FILLER_24_77 ();
 sg13g2_fill_2 FILLER_24_105 ();
 sg13g2_fill_2 FILLER_24_124 ();
 sg13g2_fill_1 FILLER_24_126 ();
 sg13g2_decap_4 FILLER_24_132 ();
 sg13g2_fill_2 FILLER_24_160 ();
 sg13g2_fill_1 FILLER_24_162 ();
 sg13g2_fill_2 FILLER_24_172 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_decap_4 FILLER_24_186 ();
 sg13g2_fill_2 FILLER_24_190 ();
 sg13g2_decap_8 FILLER_24_197 ();
 sg13g2_fill_1 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_223 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_fill_1 FILLER_24_279 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_fill_2 FILLER_24_347 ();
 sg13g2_fill_1 FILLER_24_349 ();
 sg13g2_fill_1 FILLER_24_376 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_fill_2 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_fill_1 FILLER_25_165 ();
 sg13g2_fill_2 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_decap_4 FILLER_25_218 ();
 sg13g2_decap_4 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_232 ();
 sg13g2_decap_4 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_248 ();
 sg13g2_decap_4 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_274 ();
 sg13g2_fill_1 FILLER_25_285 ();
 sg13g2_fill_2 FILLER_25_299 ();
 sg13g2_fill_1 FILLER_25_301 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_321 ();
 sg13g2_decap_4 FILLER_25_328 ();
 sg13g2_fill_2 FILLER_25_332 ();
 sg13g2_fill_2 FILLER_25_339 ();
 sg13g2_fill_1 FILLER_25_360 ();
 sg13g2_fill_2 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_367 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_fill_2 FILLER_25_390 ();
 sg13g2_fill_1 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_117 ();
 sg13g2_fill_2 FILLER_26_154 ();
 sg13g2_decap_4 FILLER_26_170 ();
 sg13g2_fill_2 FILLER_26_195 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_264 ();
 sg13g2_fill_1 FILLER_26_268 ();
 sg13g2_decap_4 FILLER_26_300 ();
 sg13g2_fill_2 FILLER_26_330 ();
 sg13g2_fill_1 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_338 ();
 sg13g2_fill_2 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_decap_4 FILLER_26_364 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_4 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_94 ();
 sg13g2_decap_4 FILLER_27_101 ();
 sg13g2_decap_8 FILLER_27_118 ();
 sg13g2_fill_2 FILLER_27_125 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_decap_4 FILLER_27_149 ();
 sg13g2_fill_2 FILLER_27_174 ();
 sg13g2_fill_1 FILLER_27_176 ();
 sg13g2_decap_4 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_201 ();
 sg13g2_decap_4 FILLER_27_211 ();
 sg13g2_fill_1 FILLER_27_228 ();
 sg13g2_fill_1 FILLER_27_251 ();
 sg13g2_fill_2 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_283 ();
 sg13g2_decap_8 FILLER_27_289 ();
 sg13g2_decap_8 FILLER_27_296 ();
 sg13g2_fill_2 FILLER_27_303 ();
 sg13g2_decap_4 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_314 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_324 ();
 sg13g2_fill_2 FILLER_27_334 ();
 sg13g2_fill_1 FILLER_27_376 ();
 sg13g2_fill_2 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_102 ();
 sg13g2_fill_2 FILLER_28_128 ();
 sg13g2_decap_4 FILLER_28_135 ();
 sg13g2_decap_8 FILLER_28_146 ();
 sg13g2_decap_4 FILLER_28_153 ();
 sg13g2_fill_2 FILLER_28_157 ();
 sg13g2_decap_8 FILLER_28_171 ();
 sg13g2_decap_4 FILLER_28_178 ();
 sg13g2_fill_1 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_fill_1 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_229 ();
 sg13g2_fill_2 FILLER_28_236 ();
 sg13g2_fill_2 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_decap_8 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_278 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_decap_8 FILLER_28_291 ();
 sg13g2_fill_2 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_319 ();
 sg13g2_decap_4 FILLER_28_325 ();
 sg13g2_fill_2 FILLER_28_329 ();
 sg13g2_fill_1 FILLER_28_341 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_decap_4 FILLER_28_366 ();
 sg13g2_fill_2 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_decap_4 FILLER_29_121 ();
 sg13g2_fill_2 FILLER_29_125 ();
 sg13g2_decap_4 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_136 ();
 sg13g2_decap_4 FILLER_29_151 ();
 sg13g2_decap_4 FILLER_29_160 ();
 sg13g2_decap_8 FILLER_29_174 ();
 sg13g2_decap_4 FILLER_29_181 ();
 sg13g2_fill_1 FILLER_29_185 ();
 sg13g2_decap_4 FILLER_29_199 ();
 sg13g2_fill_2 FILLER_29_203 ();
 sg13g2_fill_2 FILLER_29_215 ();
 sg13g2_decap_4 FILLER_29_225 ();
 sg13g2_fill_1 FILLER_29_229 ();
 sg13g2_decap_8 FILLER_29_271 ();
 sg13g2_decap_4 FILLER_29_278 ();
 sg13g2_fill_1 FILLER_29_282 ();
 sg13g2_fill_2 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_340 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_374 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_4 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_135 ();
 sg13g2_fill_2 FILLER_30_142 ();
 sg13g2_fill_2 FILLER_30_148 ();
 sg13g2_fill_2 FILLER_30_167 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_187 ();
 sg13g2_fill_2 FILLER_30_193 ();
 sg13g2_decap_4 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_207 ();
 sg13g2_decap_4 FILLER_30_217 ();
 sg13g2_fill_1 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_227 ();
 sg13g2_decap_8 FILLER_30_234 ();
 sg13g2_decap_4 FILLER_30_241 ();
 sg13g2_fill_1 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_decap_8 FILLER_30_274 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_4 FILLER_30_294 ();
 sg13g2_decap_4 FILLER_30_302 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_decap_4 FILLER_30_319 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_fill_2 FILLER_30_354 ();
 sg13g2_fill_1 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_4 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_95 ();
 sg13g2_decap_8 FILLER_31_117 ();
 sg13g2_fill_2 FILLER_31_124 ();
 sg13g2_decap_8 FILLER_31_143 ();
 sg13g2_decap_8 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_157 ();
 sg13g2_decap_8 FILLER_31_170 ();
 sg13g2_decap_8 FILLER_31_177 ();
 sg13g2_fill_2 FILLER_31_184 ();
 sg13g2_decap_8 FILLER_31_198 ();
 sg13g2_decap_4 FILLER_31_205 ();
 sg13g2_fill_1 FILLER_31_209 ();
 sg13g2_decap_8 FILLER_31_228 ();
 sg13g2_decap_4 FILLER_31_235 ();
 sg13g2_fill_2 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_260 ();
 sg13g2_decap_8 FILLER_31_267 ();
 sg13g2_decap_4 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_fill_2 FILLER_31_324 ();
 sg13g2_decap_4 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_100 ();
 sg13g2_decap_8 FILLER_32_113 ();
 sg13g2_decap_8 FILLER_32_141 ();
 sg13g2_fill_1 FILLER_32_148 ();
 sg13g2_decap_8 FILLER_32_170 ();
 sg13g2_decap_4 FILLER_32_177 ();
 sg13g2_fill_2 FILLER_32_181 ();
 sg13g2_decap_4 FILLER_32_200 ();
 sg13g2_fill_2 FILLER_32_204 ();
 sg13g2_fill_1 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_226 ();
 sg13g2_fill_1 FILLER_32_233 ();
 sg13g2_fill_2 FILLER_32_260 ();
 sg13g2_fill_2 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_290 ();
 sg13g2_fill_2 FILLER_32_297 ();
 sg13g2_fill_1 FILLER_32_299 ();
 sg13g2_decap_8 FILLER_32_313 ();
 sg13g2_decap_4 FILLER_32_320 ();
 sg13g2_fill_1 FILLER_32_324 ();
 sg13g2_fill_1 FILLER_32_342 ();
 sg13g2_fill_2 FILLER_32_360 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_4 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_115 ();
 sg13g2_decap_4 FILLER_33_122 ();
 sg13g2_decap_4 FILLER_33_142 ();
 sg13g2_decap_8 FILLER_33_163 ();
 sg13g2_decap_4 FILLER_33_195 ();
 sg13g2_fill_1 FILLER_33_199 ();
 sg13g2_fill_2 FILLER_33_223 ();
 sg13g2_fill_1 FILLER_33_229 ();
 sg13g2_fill_2 FILLER_33_235 ();
 sg13g2_fill_1 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_244 ();
 sg13g2_decap_4 FILLER_33_249 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_292 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_307 ();
 sg13g2_decap_4 FILLER_33_321 ();
 sg13g2_fill_1 FILLER_33_335 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_91 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_decap_4 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_123 ();
 sg13g2_decap_8 FILLER_34_143 ();
 sg13g2_fill_1 FILLER_34_150 ();
 sg13g2_decap_8 FILLER_34_163 ();
 sg13g2_decap_8 FILLER_34_170 ();
 sg13g2_fill_2 FILLER_34_193 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_decap_8 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_226 ();
 sg13g2_fill_1 FILLER_34_251 ();
 sg13g2_fill_2 FILLER_34_267 ();
 sg13g2_fill_2 FILLER_34_298 ();
 sg13g2_decap_4 FILLER_34_315 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_fill_1 FILLER_34_392 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_111 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_fill_2 FILLER_35_125 ();
 sg13g2_fill_1 FILLER_35_127 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_176 ();
 sg13g2_decap_4 FILLER_35_183 ();
 sg13g2_fill_1 FILLER_35_187 ();
 sg13g2_decap_8 FILLER_35_209 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_decap_8 FILLER_35_228 ();
 sg13g2_decap_8 FILLER_35_235 ();
 sg13g2_decap_8 FILLER_35_242 ();
 sg13g2_fill_2 FILLER_35_249 ();
 sg13g2_fill_1 FILLER_35_251 ();
 sg13g2_decap_4 FILLER_35_260 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_fill_1 FILLER_35_280 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_fill_2 FILLER_35_340 ();
 sg13g2_fill_2 FILLER_35_353 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_fill_1 FILLER_35_374 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_4 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_95 ();
 sg13g2_decap_4 FILLER_36_100 ();
 sg13g2_fill_2 FILLER_36_113 ();
 sg13g2_fill_1 FILLER_36_115 ();
 sg13g2_decap_8 FILLER_36_120 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_fill_2 FILLER_36_151 ();
 sg13g2_fill_1 FILLER_36_157 ();
 sg13g2_decap_4 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_decap_8 FILLER_36_194 ();
 sg13g2_decap_4 FILLER_36_201 ();
 sg13g2_fill_1 FILLER_36_224 ();
 sg13g2_decap_4 FILLER_36_232 ();
 sg13g2_fill_2 FILLER_36_236 ();
 sg13g2_decap_8 FILLER_36_242 ();
 sg13g2_decap_4 FILLER_36_249 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_fill_2 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_114 ();
 sg13g2_fill_1 FILLER_37_145 ();
 sg13g2_fill_2 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_261 ();
 sg13g2_decap_4 FILLER_37_286 ();
 sg13g2_fill_2 FILLER_37_333 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_1 FILLER_37_354 ();
 sg13g2_fill_2 FILLER_37_364 ();
 sg13g2_fill_1 FILLER_37_366 ();
 sg13g2_fill_2 FILLER_37_381 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_124 ();
 sg13g2_fill_2 FILLER_38_133 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_165 ();
 sg13g2_fill_1 FILLER_38_167 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_fill_2 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_decap_8 FILLER_38_193 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_fill_1 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_decap_4 FILLER_38_249 ();
 sg13g2_fill_2 FILLER_38_262 ();
 sg13g2_decap_8 FILLER_38_290 ();
 sg13g2_fill_2 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_fill_2 FILLER_38_309 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_1 FILLER_38_381 ();
 assign uio_oe[0] = net110;
 assign uio_oe[1] = net12;
 assign uio_oe[2] = net13;
 assign uio_oe[3] = net14;
 assign uio_oe[4] = net15;
 assign uio_oe[5] = net16;
 assign uio_oe[6] = net17;
 assign uio_oe[7] = net18;
 assign uio_out[1] = net19;
 assign uio_out[2] = net20;
 assign uio_out[3] = net21;
 assign uio_out[4] = net22;
 assign uio_out[5] = net23;
 assign uio_out[6] = net24;
 assign uio_out[7] = net25;
endmodule
