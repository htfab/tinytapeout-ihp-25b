module tt_um_2048_vga_game (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire clknet_leaf_0_clk;
 wire \btn_down_debounce.button_sync_0 ;
 wire \btn_down_debounce.button_sync_1 ;
 wire \btn_down_debounce.debounce_counter[0] ;
 wire \btn_down_debounce.debounce_counter[10] ;
 wire \btn_down_debounce.debounce_counter[11] ;
 wire \btn_down_debounce.debounce_counter[12] ;
 wire \btn_down_debounce.debounce_counter[13] ;
 wire \btn_down_debounce.debounce_counter[14] ;
 wire \btn_down_debounce.debounce_counter[15] ;
 wire \btn_down_debounce.debounce_counter[16] ;
 wire \btn_down_debounce.debounce_counter[17] ;
 wire \btn_down_debounce.debounce_counter[1] ;
 wire \btn_down_debounce.debounce_counter[2] ;
 wire \btn_down_debounce.debounce_counter[3] ;
 wire \btn_down_debounce.debounce_counter[4] ;
 wire \btn_down_debounce.debounce_counter[5] ;
 wire \btn_down_debounce.debounce_counter[6] ;
 wire \btn_down_debounce.debounce_counter[7] ;
 wire \btn_down_debounce.debounce_counter[8] ;
 wire \btn_down_debounce.debounce_counter[9] ;
 wire \btn_down_debounce.debounced ;
 wire \btn_left_debounce.button_sync_0 ;
 wire \btn_left_debounce.button_sync_1 ;
 wire \btn_left_debounce.debounce_counter[0] ;
 wire \btn_left_debounce.debounce_counter[10] ;
 wire \btn_left_debounce.debounce_counter[11] ;
 wire \btn_left_debounce.debounce_counter[12] ;
 wire \btn_left_debounce.debounce_counter[13] ;
 wire \btn_left_debounce.debounce_counter[14] ;
 wire \btn_left_debounce.debounce_counter[15] ;
 wire \btn_left_debounce.debounce_counter[16] ;
 wire \btn_left_debounce.debounce_counter[17] ;
 wire \btn_left_debounce.debounce_counter[1] ;
 wire \btn_left_debounce.debounce_counter[2] ;
 wire \btn_left_debounce.debounce_counter[3] ;
 wire \btn_left_debounce.debounce_counter[4] ;
 wire \btn_left_debounce.debounce_counter[5] ;
 wire \btn_left_debounce.debounce_counter[6] ;
 wire \btn_left_debounce.debounce_counter[7] ;
 wire \btn_left_debounce.debounce_counter[8] ;
 wire \btn_left_debounce.debounce_counter[9] ;
 wire \btn_left_debounce.debounced ;
 wire \btn_right_debounce.button_sync_0 ;
 wire \btn_right_debounce.button_sync_1 ;
 wire \btn_right_debounce.debounce_counter[0] ;
 wire \btn_right_debounce.debounce_counter[10] ;
 wire \btn_right_debounce.debounce_counter[11] ;
 wire \btn_right_debounce.debounce_counter[12] ;
 wire \btn_right_debounce.debounce_counter[13] ;
 wire \btn_right_debounce.debounce_counter[14] ;
 wire \btn_right_debounce.debounce_counter[15] ;
 wire \btn_right_debounce.debounce_counter[16] ;
 wire \btn_right_debounce.debounce_counter[17] ;
 wire \btn_right_debounce.debounce_counter[1] ;
 wire \btn_right_debounce.debounce_counter[2] ;
 wire \btn_right_debounce.debounce_counter[3] ;
 wire \btn_right_debounce.debounce_counter[4] ;
 wire \btn_right_debounce.debounce_counter[5] ;
 wire \btn_right_debounce.debounce_counter[6] ;
 wire \btn_right_debounce.debounce_counter[7] ;
 wire \btn_right_debounce.debounce_counter[8] ;
 wire \btn_right_debounce.debounce_counter[9] ;
 wire \btn_right_debounce.debounced ;
 wire btn_select_prev;
 wire \btn_up_debounce.button_sync_0 ;
 wire \btn_up_debounce.button_sync_1 ;
 wire \btn_up_debounce.debounce_counter[0] ;
 wire \btn_up_debounce.debounce_counter[10] ;
 wire \btn_up_debounce.debounce_counter[11] ;
 wire \btn_up_debounce.debounce_counter[12] ;
 wire \btn_up_debounce.debounce_counter[13] ;
 wire \btn_up_debounce.debounce_counter[14] ;
 wire \btn_up_debounce.debounce_counter[15] ;
 wire \btn_up_debounce.debounce_counter[16] ;
 wire \btn_up_debounce.debounce_counter[17] ;
 wire \btn_up_debounce.debounce_counter[1] ;
 wire \btn_up_debounce.debounce_counter[2] ;
 wire \btn_up_debounce.debounce_counter[3] ;
 wire \btn_up_debounce.debounce_counter[4] ;
 wire \btn_up_debounce.debounce_counter[5] ;
 wire \btn_up_debounce.debounce_counter[6] ;
 wire \btn_up_debounce.debounce_counter[7] ;
 wire \btn_up_debounce.debounce_counter[8] ;
 wire \btn_up_debounce.debounce_counter[9] ;
 wire \btn_up_debounce.debounced ;
 wire debug_btn_down;
 wire debug_btn_left;
 wire debug_btn_right;
 wire debug_btn_up;
 wire \debug_controller_inst.data_out_en ;
 wire \debug_controller_inst.grid_addr[0] ;
 wire \debug_controller_inst.grid_addr[1] ;
 wire \debug_controller_inst.grid_addr[2] ;
 wire \debug_controller_inst.grid_addr[3] ;
 wire \debug_controller_inst.grid_in[0] ;
 wire \debug_controller_inst.grid_in[10] ;
 wire \debug_controller_inst.grid_in[11] ;
 wire \debug_controller_inst.grid_in[12] ;
 wire \debug_controller_inst.grid_in[13] ;
 wire \debug_controller_inst.grid_in[14] ;
 wire \debug_controller_inst.grid_in[15] ;
 wire \debug_controller_inst.grid_in[16] ;
 wire \debug_controller_inst.grid_in[17] ;
 wire \debug_controller_inst.grid_in[18] ;
 wire \debug_controller_inst.grid_in[19] ;
 wire \debug_controller_inst.grid_in[1] ;
 wire \debug_controller_inst.grid_in[20] ;
 wire \debug_controller_inst.grid_in[21] ;
 wire \debug_controller_inst.grid_in[22] ;
 wire \debug_controller_inst.grid_in[23] ;
 wire \debug_controller_inst.grid_in[24] ;
 wire \debug_controller_inst.grid_in[25] ;
 wire \debug_controller_inst.grid_in[26] ;
 wire \debug_controller_inst.grid_in[27] ;
 wire \debug_controller_inst.grid_in[28] ;
 wire \debug_controller_inst.grid_in[29] ;
 wire \debug_controller_inst.grid_in[2] ;
 wire \debug_controller_inst.grid_in[30] ;
 wire \debug_controller_inst.grid_in[31] ;
 wire \debug_controller_inst.grid_in[32] ;
 wire \debug_controller_inst.grid_in[33] ;
 wire \debug_controller_inst.grid_in[34] ;
 wire \debug_controller_inst.grid_in[35] ;
 wire \debug_controller_inst.grid_in[36] ;
 wire \debug_controller_inst.grid_in[37] ;
 wire \debug_controller_inst.grid_in[38] ;
 wire \debug_controller_inst.grid_in[39] ;
 wire \debug_controller_inst.grid_in[3] ;
 wire \debug_controller_inst.grid_in[40] ;
 wire \debug_controller_inst.grid_in[41] ;
 wire \debug_controller_inst.grid_in[42] ;
 wire \debug_controller_inst.grid_in[43] ;
 wire \debug_controller_inst.grid_in[44] ;
 wire \debug_controller_inst.grid_in[45] ;
 wire \debug_controller_inst.grid_in[46] ;
 wire \debug_controller_inst.grid_in[47] ;
 wire \debug_controller_inst.grid_in[48] ;
 wire \debug_controller_inst.grid_in[49] ;
 wire \debug_controller_inst.grid_in[4] ;
 wire \debug_controller_inst.grid_in[50] ;
 wire \debug_controller_inst.grid_in[51] ;
 wire \debug_controller_inst.grid_in[52] ;
 wire \debug_controller_inst.grid_in[53] ;
 wire \debug_controller_inst.grid_in[54] ;
 wire \debug_controller_inst.grid_in[55] ;
 wire \debug_controller_inst.grid_in[56] ;
 wire \debug_controller_inst.grid_in[57] ;
 wire \debug_controller_inst.grid_in[58] ;
 wire \debug_controller_inst.grid_in[59] ;
 wire \debug_controller_inst.grid_in[5] ;
 wire \debug_controller_inst.grid_in[60] ;
 wire \debug_controller_inst.grid_in[61] ;
 wire \debug_controller_inst.grid_in[62] ;
 wire \debug_controller_inst.grid_in[63] ;
 wire \debug_controller_inst.grid_in[6] ;
 wire \debug_controller_inst.grid_in[7] ;
 wire \debug_controller_inst.grid_in[8] ;
 wire \debug_controller_inst.grid_in[9] ;
 wire \debug_controller_inst.grid_out_addr[0] ;
 wire \debug_controller_inst.grid_out_addr[1] ;
 wire \debug_controller_inst.grid_out_addr[2] ;
 wire \debug_controller_inst.grid_out_addr[3] ;
 wire \debug_controller_inst.grid_out_data[0] ;
 wire \debug_controller_inst.grid_out_data[1] ;
 wire \debug_controller_inst.grid_out_data[2] ;
 wire \debug_controller_inst.grid_out_data[3] ;
 wire \debug_controller_inst.grid_out_valid ;
 wire \draw_game_inst.board_x[0] ;
 wire \draw_game_inst.board_x[1] ;
 wire \draw_game_inst.board_x[2] ;
 wire \draw_game_inst.board_x[3] ;
 wire \draw_game_inst.board_x[4] ;
 wire \draw_game_inst.board_x[5] ;
 wire \draw_game_inst.board_y[0] ;
 wire \draw_game_inst.board_y[1] ;
 wire \draw_game_inst.board_y[2] ;
 wire \draw_game_inst.board_y[3] ;
 wire \draw_game_inst.board_y[4] ;
 wire \draw_game_inst.board_y[5] ;
 wire \draw_game_inst.board_y[6] ;
 wire \draw_game_inst.grid[0] ;
 wire \draw_game_inst.grid[10] ;
 wire \draw_game_inst.grid[11] ;
 wire \draw_game_inst.grid[12] ;
 wire \draw_game_inst.grid[13] ;
 wire \draw_game_inst.grid[14] ;
 wire \draw_game_inst.grid[15] ;
 wire \draw_game_inst.grid[16] ;
 wire \draw_game_inst.grid[17] ;
 wire \draw_game_inst.grid[18] ;
 wire \draw_game_inst.grid[19] ;
 wire \draw_game_inst.grid[1] ;
 wire \draw_game_inst.grid[20] ;
 wire \draw_game_inst.grid[21] ;
 wire \draw_game_inst.grid[22] ;
 wire \draw_game_inst.grid[23] ;
 wire \draw_game_inst.grid[24] ;
 wire \draw_game_inst.grid[25] ;
 wire \draw_game_inst.grid[26] ;
 wire \draw_game_inst.grid[27] ;
 wire \draw_game_inst.grid[28] ;
 wire \draw_game_inst.grid[29] ;
 wire \draw_game_inst.grid[2] ;
 wire \draw_game_inst.grid[30] ;
 wire \draw_game_inst.grid[31] ;
 wire \draw_game_inst.grid[32] ;
 wire \draw_game_inst.grid[33] ;
 wire \draw_game_inst.grid[34] ;
 wire \draw_game_inst.grid[35] ;
 wire \draw_game_inst.grid[36] ;
 wire \draw_game_inst.grid[37] ;
 wire \draw_game_inst.grid[38] ;
 wire \draw_game_inst.grid[39] ;
 wire \draw_game_inst.grid[3] ;
 wire \draw_game_inst.grid[40] ;
 wire \draw_game_inst.grid[41] ;
 wire \draw_game_inst.grid[42] ;
 wire \draw_game_inst.grid[43] ;
 wire \draw_game_inst.grid[44] ;
 wire \draw_game_inst.grid[45] ;
 wire \draw_game_inst.grid[46] ;
 wire \draw_game_inst.grid[47] ;
 wire \draw_game_inst.grid[48] ;
 wire \draw_game_inst.grid[49] ;
 wire \draw_game_inst.grid[4] ;
 wire \draw_game_inst.grid[50] ;
 wire \draw_game_inst.grid[51] ;
 wire \draw_game_inst.grid[52] ;
 wire \draw_game_inst.grid[53] ;
 wire \draw_game_inst.grid[54] ;
 wire \draw_game_inst.grid[55] ;
 wire \draw_game_inst.grid[56] ;
 wire \draw_game_inst.grid[57] ;
 wire \draw_game_inst.grid[58] ;
 wire \draw_game_inst.grid[59] ;
 wire \draw_game_inst.grid[5] ;
 wire \draw_game_inst.grid[60] ;
 wire \draw_game_inst.grid[61] ;
 wire \draw_game_inst.grid[62] ;
 wire \draw_game_inst.grid[63] ;
 wire \draw_game_inst.grid[6] ;
 wire \draw_game_inst.grid[7] ;
 wire \draw_game_inst.grid[8] ;
 wire \draw_game_inst.grid[9] ;
 wire \draw_game_inst.new_tiles[0] ;
 wire \draw_game_inst.new_tiles[10] ;
 wire \draw_game_inst.new_tiles[11] ;
 wire \draw_game_inst.new_tiles[12] ;
 wire \draw_game_inst.new_tiles[13] ;
 wire \draw_game_inst.new_tiles[14] ;
 wire \draw_game_inst.new_tiles[15] ;
 wire \draw_game_inst.new_tiles[1] ;
 wire \draw_game_inst.new_tiles[2] ;
 wire \draw_game_inst.new_tiles[3] ;
 wire \draw_game_inst.new_tiles[4] ;
 wire \draw_game_inst.new_tiles[5] ;
 wire \draw_game_inst.new_tiles[6] ;
 wire \draw_game_inst.new_tiles[7] ;
 wire \draw_game_inst.new_tiles[8] ;
 wire \draw_game_inst.new_tiles[9] ;
 wire \draw_game_inst.new_tiles_counter[0] ;
 wire \draw_game_inst.new_tiles_counter[1] ;
 wire \draw_game_inst.new_tiles_counter[2] ;
 wire \draw_game_inst.x[6] ;
 wire \draw_game_inst.x[7] ;
 wire \draw_game_inst.x[8] ;
 wire \draw_game_inst.x[9] ;
 wire \draw_game_inst.y[7] ;
 wire \draw_game_inst.y[8] ;
 wire \draw_game_inst.y[9] ;
 wire \game_logic_inst.add_new_tiles[0] ;
 wire \game_logic_inst.add_new_tiles[1] ;
 wire \game_logic_inst.added_tile_index[0] ;
 wire \game_logic_inst.added_tile_index[1] ;
 wire \game_logic_inst.added_tile_index[2] ;
 wire \game_logic_inst.added_tile_index[3] ;
 wire \game_logic_inst.calculate_move ;
 wire \game_logic_inst.current_direction[1] ;
 wire \game_logic_inst.current_direction[2] ;
 wire \game_logic_inst.current_direction[3] ;
 wire \game_logic_inst.current_row_index[0] ;
 wire \game_logic_inst.current_row_index[1] ;
 wire \game_logic_inst.debug_move_reg ;
 wire \game_logic_inst.game_started ;
 wire \game_logic_inst.lfsr_shift[0] ;
 wire \game_logic_inst.lfsr_shift[1] ;
 wire \game_logic_inst.lfsr_value[0] ;
 wire \game_logic_inst.lfsr_value[10] ;
 wire \game_logic_inst.lfsr_value[11] ;
 wire \game_logic_inst.lfsr_value[12] ;
 wire \game_logic_inst.lfsr_value[13] ;
 wire \game_logic_inst.lfsr_value[14] ;
 wire \game_logic_inst.lfsr_value[15] ;
 wire \game_logic_inst.lfsr_value[1] ;
 wire \game_logic_inst.lfsr_value[2] ;
 wire \game_logic_inst.lfsr_value[3] ;
 wire \game_logic_inst.lfsr_value[4] ;
 wire \game_logic_inst.lfsr_value[5] ;
 wire \game_logic_inst.lfsr_value[6] ;
 wire \game_logic_inst.lfsr_value[7] ;
 wire \game_logic_inst.lfsr_value[8] ;
 wire \game_logic_inst.lfsr_value[9] ;
 wire \game_logic_inst.prev_any_button_pressed ;
 wire \game_logic_inst.should_transpose ;
 wire \game_logic_inst.valid_move ;
 wire \gamepad_pmod.decoder.data_reg[0] ;
 wire \gamepad_pmod.decoder.data_reg[10] ;
 wire \gamepad_pmod.decoder.data_reg[11] ;
 wire \gamepad_pmod.decoder.data_reg[1] ;
 wire \gamepad_pmod.decoder.data_reg[2] ;
 wire \gamepad_pmod.decoder.data_reg[3] ;
 wire \gamepad_pmod.decoder.data_reg[4] ;
 wire \gamepad_pmod.decoder.data_reg[5] ;
 wire \gamepad_pmod.decoder.data_reg[6] ;
 wire \gamepad_pmod.decoder.data_reg[7] ;
 wire \gamepad_pmod.decoder.data_reg[8] ;
 wire \gamepad_pmod.decoder.data_reg[9] ;
 wire \gamepad_pmod.driver.pmod_clk_prev ;
 wire \gamepad_pmod.driver.pmod_clk_sync[0] ;
 wire \gamepad_pmod.driver.pmod_clk_sync[1] ;
 wire \gamepad_pmod.driver.pmod_data_sync[0] ;
 wire \gamepad_pmod.driver.pmod_data_sync[1] ;
 wire \gamepad_pmod.driver.pmod_latch_prev ;
 wire \gamepad_pmod.driver.pmod_latch_sync[0] ;
 wire \gamepad_pmod.driver.pmod_latch_sync[1] ;
 wire \gamepad_pmod.driver.shift_reg[0] ;
 wire \gamepad_pmod.driver.shift_reg[10] ;
 wire \gamepad_pmod.driver.shift_reg[11] ;
 wire \gamepad_pmod.driver.shift_reg[1] ;
 wire \gamepad_pmod.driver.shift_reg[2] ;
 wire \gamepad_pmod.driver.shift_reg[3] ;
 wire \gamepad_pmod.driver.shift_reg[4] ;
 wire \gamepad_pmod.driver.shift_reg[5] ;
 wire \gamepad_pmod.driver.shift_reg[6] ;
 wire \gamepad_pmod.driver.shift_reg[7] ;
 wire \gamepad_pmod.driver.shift_reg[8] ;
 wire \gamepad_pmod.driver.shift_reg[9] ;
 wire hsync;
 wire \lfsr_inst.lfsr[16] ;
 wire \lfsr_inst.lfsr[17] ;
 wire \lfsr_inst.lfsr[18] ;
 wire \lfsr_inst.lfsr[19] ;
 wire \lfsr_inst.lfsr[20] ;
 wire \lfsr_inst.lfsr[21] ;
 wire \lfsr_inst.lfsr[22] ;
 wire \lfsr_inst.lfsr[23] ;
 wire \lfsr_inst.lfsr[24] ;
 wire \lfsr_inst.lfsr[25] ;
 wire \lfsr_inst.lfsr[26] ;
 wire \lfsr_inst.lfsr[27] ;
 wire \lfsr_inst.lfsr[28] ;
 wire \lfsr_inst.lfsr[29] ;
 wire \lfsr_inst.lfsr[30] ;
 wire \lfsr_inst.lfsr[31] ;
 wire \new_tiles_counter[0] ;
 wire \new_tiles_counter[4] ;
 wire retro_colors;
 wire show_welcome_screen;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire \vga_sync_gen.vsync ;
 wire vsync_prev;
 wire \welcome_screen_grid[0] ;
 wire \welcome_screen_grid[11] ;
 wire \welcome_screen_grid[12] ;
 wire \welcome_screen_grid[16] ;
 wire \welcome_screen_grid[20] ;
 wire \welcome_screen_grid[24] ;
 wire \welcome_screen_grid[28] ;
 wire \welcome_screen_grid[32] ;
 wire \welcome_screen_grid[36] ;
 wire \welcome_screen_grid[40] ;
 wire \welcome_screen_grid[44] ;
 wire \welcome_screen_grid[48] ;
 wire \welcome_screen_grid[4] ;
 wire \welcome_screen_grid[52] ;
 wire \welcome_screen_grid[56] ;
 wire \welcome_screen_grid[60] ;
 wire \welcome_screen_inst.welcome_counter[0] ;
 wire \welcome_screen_inst.welcome_counter[1] ;
 wire \welcome_screen_inst.welcome_counter[2] ;
 wire \welcome_screen_inst.welcome_counter[3] ;
 wire \welcome_screen_inst.welcome_counter[4] ;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;

 sg13g2_inv_2 _4755_ (.Y(_3975_),
    .A(net955));
 sg13g2_inv_1 _4756_ (.Y(_3976_),
    .A(net2127));
 sg13g2_inv_1 _4757_ (.Y(_3977_),
    .A(net2130));
 sg13g2_inv_1 _4758_ (.Y(_3978_),
    .A(net2136));
 sg13g2_inv_1 _4759_ (.Y(_3979_),
    .A(net2142));
 sg13g2_inv_1 _4760_ (.Y(_3980_),
    .A(net16));
 sg13g2_inv_1 _4761_ (.Y(_3981_),
    .A(net15));
 sg13g2_inv_1 _4762_ (.Y(_3982_),
    .A(net2146));
 sg13g2_inv_1 _4763_ (.Y(_3983_),
    .A(net14));
 sg13g2_inv_1 _4764_ (.Y(_3984_),
    .A(net2149));
 sg13g2_inv_1 _4765_ (.Y(_3985_),
    .A(net13));
 sg13g2_inv_2 _4766_ (.Y(_3986_),
    .A(net2178));
 sg13g2_inv_1 _4767_ (.Y(_3987_),
    .A(net954));
 sg13g2_inv_1 _4768_ (.Y(_3988_),
    .A(net676));
 sg13g2_inv_1 _4769_ (.Y(_3989_),
    .A(net742));
 sg13g2_inv_2 _4770_ (.Y(_3990_),
    .A(net837));
 sg13g2_inv_1 _4771_ (.Y(_3991_),
    .A(net540));
 sg13g2_inv_1 _4772_ (.Y(_3992_),
    .A(\gamepad_pmod.driver.shift_reg[10] ));
 sg13g2_inv_1 _4773_ (.Y(_3993_),
    .A(net467));
 sg13g2_inv_1 _4774_ (.Y(_3994_),
    .A(net591));
 sg13g2_inv_1 _4775_ (.Y(_3995_),
    .A(net595));
 sg13g2_inv_1 _4776_ (.Y(_3996_),
    .A(net607));
 sg13g2_inv_1 _4777_ (.Y(_3997_),
    .A(net614));
 sg13g2_inv_1 _4778_ (.Y(_3998_),
    .A(net655));
 sg13g2_inv_1 _4779_ (.Y(_3999_),
    .A(net605));
 sg13g2_inv_1 _4780_ (.Y(_4000_),
    .A(\gamepad_pmod.driver.shift_reg[2] ));
 sg13g2_inv_1 _4781_ (.Y(_4001_),
    .A(net469));
 sg13g2_inv_1 _4782_ (.Y(_4002_),
    .A(net586));
 sg13g2_inv_1 _4783_ (.Y(_4003_),
    .A(net512));
 sg13g2_inv_1 _4784_ (.Y(_4004_),
    .A(net645));
 sg13g2_inv_1 _4785_ (.Y(_4005_),
    .A(\btn_left_debounce.debounced ));
 sg13g2_inv_1 _4786_ (.Y(_4006_),
    .A(\btn_down_debounce.debounced ));
 sg13g2_inv_1 _4787_ (.Y(_4007_),
    .A(net616));
 sg13g2_inv_1 _4788_ (.Y(_4008_),
    .A(net465));
 sg13g2_inv_1 _4789_ (.Y(_4009_),
    .A(net2275));
 sg13g2_inv_1 _4790_ (.Y(_4010_),
    .A(net490));
 sg13g2_inv_1 _4791_ (.Y(_4011_),
    .A(net510));
 sg13g2_inv_1 _4792_ (.Y(_4012_),
    .A(net518));
 sg13g2_inv_1 _4793_ (.Y(_4013_),
    .A(net506));
 sg13g2_inv_1 _4794_ (.Y(_4014_),
    .A(net602));
 sg13g2_inv_1 _4795_ (.Y(_4015_),
    .A(net560));
 sg13g2_inv_1 _4796_ (.Y(_4016_),
    .A(net550));
 sg13g2_inv_1 _4797_ (.Y(_4017_),
    .A(net557));
 sg13g2_inv_1 _4798_ (.Y(_4018_),
    .A(net559));
 sg13g2_inv_1 _4799_ (.Y(_4019_),
    .A(net682));
 sg13g2_inv_1 _4800_ (.Y(_4020_),
    .A(net508));
 sg13g2_inv_1 _4801_ (.Y(_4021_),
    .A(net534));
 sg13g2_inv_1 _4802_ (.Y(_4022_),
    .A(net2268));
 sg13g2_inv_1 _4803_ (.Y(_4023_),
    .A(net2161));
 sg13g2_inv_1 _4804_ (.Y(_4024_),
    .A(net2319));
 sg13g2_inv_1 _4805_ (.Y(_4025_),
    .A(net916));
 sg13g2_inv_1 _4806_ (.Y(_4026_),
    .A(\lfsr_inst.lfsr[31] ));
 sg13g2_inv_1 _4807_ (.Y(_4027_),
    .A(\debug_controller_inst.grid_in[20] ));
 sg13g2_inv_1 _4808_ (.Y(_4028_),
    .A(\debug_controller_inst.grid_in[52] ));
 sg13g2_inv_1 _4809_ (.Y(_4029_),
    .A(\debug_controller_inst.grid_in[21] ));
 sg13g2_inv_1 _4810_ (.Y(_4030_),
    .A(\debug_controller_inst.grid_in[53] ));
 sg13g2_inv_1 _4811_ (.Y(_4031_),
    .A(\debug_controller_inst.grid_in[22] ));
 sg13g2_inv_1 _4812_ (.Y(_4032_),
    .A(\debug_controller_inst.grid_in[54] ));
 sg13g2_inv_1 _4813_ (.Y(_4033_),
    .A(\debug_controller_inst.grid_in[23] ));
 sg13g2_inv_1 _4814_ (.Y(_4034_),
    .A(\debug_controller_inst.grid_in[55] ));
 sg13g2_inv_1 _4815_ (.Y(_4035_),
    .A(\btn_up_debounce.debounce_counter[13] ));
 sg13g2_inv_1 _4816_ (.Y(_4036_),
    .A(\btn_right_debounce.debounce_counter[13] ));
 sg13g2_inv_1 _4817_ (.Y(_4037_),
    .A(\btn_left_debounce.debounce_counter[14] ));
 sg13g2_inv_1 _4818_ (.Y(_4038_),
    .A(\btn_down_debounce.debounce_counter[7] ));
 sg13g2_inv_1 _4819_ (.Y(_4039_),
    .A(\draw_game_inst.x[8] ));
 sg13g2_inv_1 _4820_ (.Y(_4040_),
    .A(\draw_game_inst.y[9] ));
 sg13g2_inv_1 _4821_ (.Y(_4041_),
    .A(net2179));
 sg13g2_inv_2 _4822_ (.Y(_4042_),
    .A(net2184));
 sg13g2_inv_1 _4823_ (.Y(_4043_),
    .A(net2195));
 sg13g2_inv_2 _4824_ (.Y(_4044_),
    .A(net2211));
 sg13g2_inv_1 _4825_ (.Y(_4045_),
    .A(net2246));
 sg13g2_inv_2 _4826_ (.Y(_4046_),
    .A(net2300));
 sg13g2_inv_1 _4827_ (.Y(_4047_),
    .A(net2287));
 sg13g2_inv_2 _4828_ (.Y(_4048_),
    .A(net2290));
 sg13g2_inv_1 _4829_ (.Y(_4049_),
    .A(net2282));
 sg13g2_inv_2 _4830_ (.Y(_4050_),
    .A(net2158));
 sg13g2_inv_1 _4831_ (.Y(_4051_),
    .A(\game_logic_inst.added_tile_index[1] ));
 sg13g2_inv_1 _4832_ (.Y(_4052_),
    .A(\game_logic_inst.added_tile_index[0] ));
 sg13g2_inv_1 _4833_ (.Y(_4053_),
    .A(net456));
 sg13g2_inv_1 _4834_ (.Y(_4054_),
    .A(net982));
 sg13g2_inv_4 _4835_ (.A(net2284),
    .Y(_4055_));
 sg13g2_inv_1 _4836_ (.Y(_4056_),
    .A(_0099_));
 sg13g2_inv_1 _4837_ (.Y(_4057_),
    .A(\debug_controller_inst.grid_out_valid ));
 sg13g2_inv_1 _4838_ (.Y(_4058_),
    .A(net1004));
 sg13g2_inv_1 _4839_ (.Y(_4059_),
    .A(net991));
 sg13g2_inv_1 _4840_ (.Y(_4060_),
    .A(net993));
 sg13g2_inv_1 _4841_ (.Y(_4061_),
    .A(_0110_));
 sg13g2_inv_1 _4842_ (.Y(_4062_),
    .A(net952));
 sg13g2_inv_1 _4843_ (.Y(_4063_),
    .A(net1016));
 sg13g2_inv_1 _4844_ (.Y(_4064_),
    .A(net1014));
 sg13g2_inv_1 _4845_ (.Y(_4065_),
    .A(_0118_));
 sg13g2_inv_1 _4846_ (.Y(_4066_),
    .A(net1002));
 sg13g2_inv_1 _4847_ (.Y(_4067_),
    .A(net1012));
 sg13g2_inv_1 _4848_ (.Y(_4068_),
    .A(net1024));
 sg13g2_inv_1 _4849_ (.Y(_4069_),
    .A(net1001));
 sg13g2_inv_1 _4850_ (.Y(_4070_),
    .A(net913));
 sg13g2_inv_1 _4851_ (.Y(_4071_),
    .A(net1022));
 sg13g2_inv_1 _4852_ (.Y(_4072_),
    .A(net1018));
 sg13g2_inv_1 _4853_ (.Y(_4073_),
    .A(net999));
 sg13g2_inv_1 _4854_ (.Y(_4074_),
    .A(net889));
 sg13g2_inv_1 _4855_ (.Y(_4075_),
    .A(net443));
 sg13g2_inv_1 _4856_ (.Y(_4076_),
    .A(net441));
 sg13g2_nand4_1 _4857_ (.B(\gamepad_pmod.decoder.data_reg[8] ),
    .C(\gamepad_pmod.decoder.data_reg[11] ),
    .A(\gamepad_pmod.decoder.data_reg[9] ),
    .Y(_4077_),
    .D(\gamepad_pmod.decoder.data_reg[10] ));
 sg13g2_nand4_1 _4858_ (.B(\gamepad_pmod.decoder.data_reg[4] ),
    .C(\gamepad_pmod.decoder.data_reg[7] ),
    .A(\gamepad_pmod.decoder.data_reg[5] ),
    .Y(_4078_),
    .D(\gamepad_pmod.decoder.data_reg[6] ));
 sg13g2_nand4_1 _4859_ (.B(\gamepad_pmod.decoder.data_reg[0] ),
    .C(\gamepad_pmod.decoder.data_reg[3] ),
    .A(\gamepad_pmod.decoder.data_reg[1] ),
    .Y(_0495_),
    .D(\gamepad_pmod.decoder.data_reg[2] ));
 sg13g2_or3_2 _4860_ (.A(_4077_),
    .B(_4078_),
    .C(_0495_),
    .X(_0496_));
 sg13g2_a21o_1 _4861_ (.A2(_0496_),
    .A1(\gamepad_pmod.decoder.data_reg[6] ),
    .B1(\btn_down_debounce.debounced ),
    .X(_0497_));
 sg13g2_a21oi_2 _4862_ (.B1(debug_btn_down),
    .Y(_0498_),
    .A2(_0497_),
    .A1(_0165_));
 sg13g2_a21o_2 _4863_ (.A2(_0496_),
    .A1(\gamepad_pmod.decoder.data_reg[7] ),
    .B1(\btn_up_debounce.debounced ),
    .X(_0499_));
 sg13g2_a21oi_2 _4864_ (.B1(net844),
    .Y(_0500_),
    .A2(_0499_),
    .A1(_0165_));
 sg13g2_a21o_1 _4865_ (.A2(_0496_),
    .A1(\gamepad_pmod.decoder.data_reg[5] ),
    .B1(\btn_left_debounce.debounced ),
    .X(_0501_));
 sg13g2_a21oi_1 _4866_ (.A1(_0165_),
    .A2(_0501_),
    .Y(_0502_),
    .B1(net1025));
 sg13g2_a21o_2 _4867_ (.A2(_0496_),
    .A1(\gamepad_pmod.decoder.data_reg[4] ),
    .B1(\btn_right_debounce.debounced ),
    .X(_0503_));
 sg13g2_a21oi_1 _4868_ (.A1(_0165_),
    .A2(_0503_),
    .Y(_0504_),
    .B1(debug_btn_right));
 sg13g2_a21o_1 _4869_ (.A2(_0503_),
    .A1(_0165_),
    .B1(debug_btn_right),
    .X(_0505_));
 sg13g2_nand4_1 _4870_ (.B(_0500_),
    .C(_0502_),
    .A(_0498_),
    .Y(_0506_),
    .D(_0504_));
 sg13g2_nor2b_1 _4871_ (.A(\game_logic_inst.prev_any_button_pressed ),
    .B_N(_0506_),
    .Y(_0507_));
 sg13g2_nand2b_2 _4872_ (.Y(_0508_),
    .B(_0506_),
    .A_N(\game_logic_inst.prev_any_button_pressed ));
 sg13g2_o21ai_1 _4873_ (.B1(net2170),
    .Y(_0509_),
    .A1(net851),
    .A2(_0507_));
 sg13g2_and2_1 _4874_ (.A(net2314),
    .B(_0509_),
    .X(_0510_));
 sg13g2_nor2_2 _4875_ (.A(net2302),
    .B(net851),
    .Y(_0511_));
 sg13g2_nand3_1 _4876_ (.B(_0507_),
    .C(_0511_),
    .A(_0502_),
    .Y(_0512_));
 sg13g2_nor3_1 _4877_ (.A(_0498_),
    .B(_0505_),
    .C(_0512_),
    .Y(_0513_));
 sg13g2_a22oi_1 _4878_ (.Y(_0514_),
    .B1(_0513_),
    .B2(net845),
    .A2(_0510_),
    .A1(\game_logic_inst.current_direction[3] ));
 sg13g2_inv_1 _4879_ (.Y(_0002_),
    .A(net846));
 sg13g2_nand2_1 _4880_ (.Y(_0515_),
    .A(net863),
    .B(_0510_));
 sg13g2_o21ai_1 _4881_ (.B1(_0515_),
    .Y(_0001_),
    .A1(_0504_),
    .A2(_0512_));
 sg13g2_nor3_1 _4882_ (.A(_0500_),
    .B(_0505_),
    .C(_0512_),
    .Y(_0516_));
 sg13g2_a21o_1 _4883_ (.A2(_0510_),
    .A1(net555),
    .B1(_0516_),
    .X(_0000_));
 sg13g2_nor2_1 _4884_ (.A(net2139),
    .B(net2140),
    .Y(_0517_));
 sg13g2_nor3_2 _4885_ (.A(net2137),
    .B(net2139),
    .C(net2140),
    .Y(_0518_));
 sg13g2_nand2b_2 _4886_ (.Y(_0519_),
    .B(_0518_),
    .A_N(\debug_controller_inst.grid_out_addr[3] ));
 sg13g2_nor2_2 _4887_ (.A(_4057_),
    .B(_0519_),
    .Y(_0520_));
 sg13g2_nor2_1 _4888_ (.A(net2153),
    .B(net2157),
    .Y(_0521_));
 sg13g2_nor2_1 _4889_ (.A(\game_logic_inst.current_direction[3] ),
    .B(\game_logic_inst.current_direction[2] ),
    .Y(_0522_));
 sg13g2_or2_1 _4890_ (.X(_0523_),
    .B(\game_logic_inst.current_direction[2] ),
    .A(\game_logic_inst.current_direction[3] ));
 sg13g2_nor2b_1 _4891_ (.A(net2153),
    .B_N(net2157),
    .Y(_0524_));
 sg13g2_nor2b_1 _4892_ (.A(net2157),
    .B_N(net2153),
    .Y(_0525_));
 sg13g2_nand2b_2 _4893_ (.Y(_0526_),
    .B(net2153),
    .A_N(net2157));
 sg13g2_and2_1 _4894_ (.A(net2153),
    .B(net2157),
    .X(_0527_));
 sg13g2_nand2_1 _4895_ (.Y(_0528_),
    .A(net2153),
    .B(net2157));
 sg13g2_mux4_1 _4896_ (.S0(net2154),
    .A0(\debug_controller_inst.grid_in[0] ),
    .A1(\debug_controller_inst.grid_in[16] ),
    .A2(\debug_controller_inst.grid_in[32] ),
    .A3(\debug_controller_inst.grid_in[48] ),
    .S1(net2150),
    .X(_0529_));
 sg13g2_and2_1 _4897_ (.A(net2053),
    .B(_0529_),
    .X(_0530_));
 sg13g2_mux4_1 _4898_ (.S0(net2156),
    .A0(\debug_controller_inst.grid_in[12] ),
    .A1(\debug_controller_inst.grid_in[28] ),
    .A2(\debug_controller_inst.grid_in[44] ),
    .A3(\debug_controller_inst.grid_in[60] ),
    .S1(net2152),
    .X(_0531_));
 sg13g2_a21oi_2 _4899_ (.B1(_0530_),
    .Y(_0532_),
    .A2(_0531_),
    .A1(net2056));
 sg13g2_a21o_2 _4900_ (.A2(_0531_),
    .A1(net2056),
    .B1(_0530_),
    .X(_0533_));
 sg13g2_mux4_1 _4901_ (.S0(net2154),
    .A0(\debug_controller_inst.grid_in[5] ),
    .A1(\debug_controller_inst.grid_in[21] ),
    .A2(\debug_controller_inst.grid_in[37] ),
    .A3(\debug_controller_inst.grid_in[53] ),
    .S1(net2150),
    .X(_0534_));
 sg13g2_mux4_1 _4902_ (.S0(net2155),
    .A0(\debug_controller_inst.grid_in[9] ),
    .A1(\debug_controller_inst.grid_in[25] ),
    .A2(\debug_controller_inst.grid_in[41] ),
    .A3(\debug_controller_inst.grid_in[57] ),
    .S1(net2151),
    .X(_0535_));
 sg13g2_mux2_1 _4903_ (.A0(_0534_),
    .A1(_0535_),
    .S(net2055),
    .X(_0536_));
 sg13g2_mux4_1 _4904_ (.S0(net2156),
    .A0(\debug_controller_inst.grid_in[4] ),
    .A1(\debug_controller_inst.grid_in[20] ),
    .A2(\debug_controller_inst.grid_in[36] ),
    .A3(\debug_controller_inst.grid_in[52] ),
    .S1(net2152),
    .X(_0537_));
 sg13g2_inv_2 _4905_ (.Y(_0538_),
    .A(_0537_));
 sg13g2_nand2_1 _4906_ (.Y(_0539_),
    .A(net2051),
    .B(_0537_));
 sg13g2_mux4_1 _4907_ (.S0(net2156),
    .A0(\debug_controller_inst.grid_in[8] ),
    .A1(\debug_controller_inst.grid_in[24] ),
    .A2(\debug_controller_inst.grid_in[40] ),
    .A3(\debug_controller_inst.grid_in[56] ),
    .S1(net2152),
    .X(_0540_));
 sg13g2_nand2_1 _4908_ (.Y(_0541_),
    .A(net2055),
    .B(_0540_));
 sg13g2_nand2_2 _4909_ (.Y(_0542_),
    .A(_0539_),
    .B(_0541_));
 sg13g2_inv_2 _4910_ (.Y(_0543_),
    .A(_0542_));
 sg13g2_mux4_1 _4911_ (.S0(net2155),
    .A0(\debug_controller_inst.grid_in[6] ),
    .A1(\debug_controller_inst.grid_in[22] ),
    .A2(\debug_controller_inst.grid_in[38] ),
    .A3(\debug_controller_inst.grid_in[54] ),
    .S1(net2150),
    .X(_0544_));
 sg13g2_nand2_1 _4912_ (.Y(_0545_),
    .A(net2052),
    .B(_0544_));
 sg13g2_mux4_1 _4913_ (.S0(net2155),
    .A0(\debug_controller_inst.grid_in[10] ),
    .A1(\debug_controller_inst.grid_in[26] ),
    .A2(\debug_controller_inst.grid_in[42] ),
    .A3(\debug_controller_inst.grid_in[58] ),
    .S1(net2151),
    .X(_0546_));
 sg13g2_nand2_1 _4914_ (.Y(_0547_),
    .A(net2055),
    .B(_0546_));
 sg13g2_nand2_2 _4915_ (.Y(_0548_),
    .A(_0545_),
    .B(_0547_));
 sg13g2_mux4_1 _4916_ (.S0(net2154),
    .A0(\debug_controller_inst.grid_in[7] ),
    .A1(\debug_controller_inst.grid_in[23] ),
    .A2(\debug_controller_inst.grid_in[39] ),
    .A3(\debug_controller_inst.grid_in[55] ),
    .S1(net2150),
    .X(_0549_));
 sg13g2_mux4_1 _4917_ (.S0(net2155),
    .A0(\debug_controller_inst.grid_in[11] ),
    .A1(\debug_controller_inst.grid_in[27] ),
    .A2(\debug_controller_inst.grid_in[43] ),
    .A3(\debug_controller_inst.grid_in[59] ),
    .S1(net2151),
    .X(_0550_));
 sg13g2_mux2_1 _4918_ (.A0(_0549_),
    .A1(_0550_),
    .S(net2056),
    .X(_0551_));
 sg13g2_nor4_2 _4919_ (.A(_0536_),
    .B(_0542_),
    .C(_0548_),
    .Y(_0552_),
    .D(_0551_));
 sg13g2_mux4_1 _4920_ (.S0(net2154),
    .A0(\debug_controller_inst.grid_in[14] ),
    .A1(\debug_controller_inst.grid_in[30] ),
    .A2(\debug_controller_inst.grid_in[46] ),
    .A3(\debug_controller_inst.grid_in[62] ),
    .S1(net2151),
    .X(_0553_));
 sg13g2_mux4_1 _4921_ (.S0(net2154),
    .A0(\debug_controller_inst.grid_in[2] ),
    .A1(\debug_controller_inst.grid_in[18] ),
    .A2(\debug_controller_inst.grid_in[34] ),
    .A3(\debug_controller_inst.grid_in[50] ),
    .S1(net2150),
    .X(_0554_));
 sg13g2_mux2_2 _4922_ (.A0(_0553_),
    .A1(_0554_),
    .S(net2056),
    .X(_0555_));
 sg13g2_mux4_1 _4923_ (.S0(net2154),
    .A0(\debug_controller_inst.grid_in[15] ),
    .A1(\debug_controller_inst.grid_in[31] ),
    .A2(\debug_controller_inst.grid_in[47] ),
    .A3(\debug_controller_inst.grid_in[63] ),
    .S1(net2150),
    .X(_0556_));
 sg13g2_mux4_1 _4924_ (.S0(net2154),
    .A0(\debug_controller_inst.grid_in[3] ),
    .A1(\debug_controller_inst.grid_in[19] ),
    .A2(\debug_controller_inst.grid_in[35] ),
    .A3(\debug_controller_inst.grid_in[51] ),
    .S1(net2150),
    .X(_0557_));
 sg13g2_mux2_2 _4925_ (.A0(_0556_),
    .A1(_0557_),
    .S(net2055),
    .X(_0558_));
 sg13g2_mux2_2 _4926_ (.A0(_0529_),
    .A1(_0531_),
    .S(net2052),
    .X(_0559_));
 sg13g2_inv_1 _4927_ (.Y(_0560_),
    .A(_0559_));
 sg13g2_mux4_1 _4928_ (.S0(net2155),
    .A0(\debug_controller_inst.grid_in[1] ),
    .A1(\debug_controller_inst.grid_in[17] ),
    .A2(\debug_controller_inst.grid_in[33] ),
    .A3(\debug_controller_inst.grid_in[49] ),
    .S1(net2151),
    .X(_0561_));
 sg13g2_mux4_1 _4929_ (.S0(net2154),
    .A0(\debug_controller_inst.grid_in[13] ),
    .A1(\debug_controller_inst.grid_in[29] ),
    .A2(\debug_controller_inst.grid_in[45] ),
    .A3(\debug_controller_inst.grid_in[61] ),
    .S1(net2150),
    .X(_0562_));
 sg13g2_mux2_2 _4930_ (.A0(_0561_),
    .A1(_0562_),
    .S(net2051),
    .X(_0563_));
 sg13g2_inv_1 _4931_ (.Y(_0564_),
    .A(_0563_));
 sg13g2_nor4_2 _4932_ (.A(_0555_),
    .B(_0558_),
    .C(_0559_),
    .Y(_0565_),
    .D(_0563_));
 sg13g2_or4_2 _4933_ (.A(_0555_),
    .B(_0558_),
    .C(_0559_),
    .D(_0563_),
    .X(_0566_));
 sg13g2_mux2_2 _4934_ (.A0(_0544_),
    .A1(_0546_),
    .S(net2052),
    .X(_0567_));
 sg13g2_mux2_2 _4935_ (.A0(_0534_),
    .A1(_0535_),
    .S(net2051),
    .X(_0568_));
 sg13g2_mux2_2 _4936_ (.A0(_0537_),
    .A1(_0540_),
    .S(net2051),
    .X(_0569_));
 sg13g2_mux2_2 _4937_ (.A0(_0549_),
    .A1(_0550_),
    .S(net2052),
    .X(_0570_));
 sg13g2_inv_1 _4938_ (.Y(_0571_),
    .A(_0570_));
 sg13g2_nor4_2 _4939_ (.A(_0567_),
    .B(_0568_),
    .C(_0569_),
    .Y(_0572_),
    .D(_0570_));
 sg13g2_and2_2 _4940_ (.A(_0565_),
    .B(_0572_),
    .X(_0573_));
 sg13g2_xnor2_1 _4941_ (.Y(_0574_),
    .A(_0555_),
    .B(_0567_));
 sg13g2_xnor2_1 _4942_ (.Y(_0575_),
    .A(_0559_),
    .B(_0569_));
 sg13g2_xnor2_1 _4943_ (.Y(_0576_),
    .A(_0563_),
    .B(_0568_));
 sg13g2_xnor2_1 _4944_ (.Y(_0577_),
    .A(_0558_),
    .B(_0570_));
 sg13g2_and4_2 _4945_ (.A(_0574_),
    .B(_0575_),
    .C(_0576_),
    .D(_0577_),
    .X(_0578_));
 sg13g2_nand4_1 _4946_ (.B(_0575_),
    .C(_0576_),
    .A(_0574_),
    .Y(_0579_),
    .D(_0577_));
 sg13g2_nor3_2 _4947_ (.A(_0565_),
    .B(_0572_),
    .C(_0578_),
    .Y(_0580_));
 sg13g2_inv_1 _4948_ (.Y(_0581_),
    .A(_0580_));
 sg13g2_or2_2 _4949_ (.X(_0582_),
    .B(_0580_),
    .A(_0573_));
 sg13g2_and2_1 _4950_ (.A(_0559_),
    .B(_0563_),
    .X(_0583_));
 sg13g2_and2_1 _4951_ (.A(_0578_),
    .B(_0583_),
    .X(_0584_));
 sg13g2_a21oi_1 _4952_ (.A1(_0578_),
    .A2(_0583_),
    .Y(_0585_),
    .B1(_0555_));
 sg13g2_nand2_1 _4953_ (.Y(_0586_),
    .A(_0555_),
    .B(_0583_));
 sg13g2_o21ai_1 _4954_ (.B1(_0566_),
    .Y(_0587_),
    .A1(net1816),
    .A2(_0586_));
 sg13g2_nand2_1 _4955_ (.Y(_0588_),
    .A(_0565_),
    .B(_0567_));
 sg13g2_o21ai_1 _4956_ (.B1(_0588_),
    .Y(_0589_),
    .A1(_0585_),
    .A2(_0587_));
 sg13g2_xnor2_1 _4957_ (.Y(_0590_),
    .A(_0548_),
    .B(_0589_));
 sg13g2_nand2_1 _4958_ (.Y(_0591_),
    .A(_0560_),
    .B(net1816));
 sg13g2_a21oi_1 _4959_ (.A1(_0559_),
    .A2(_0578_),
    .Y(_0592_),
    .B1(_0565_));
 sg13g2_a22oi_1 _4960_ (.Y(_0593_),
    .B1(_0591_),
    .B2(_0592_),
    .A2(_0569_),
    .A1(_0565_));
 sg13g2_xnor2_1 _4961_ (.Y(_0594_),
    .A(_0543_),
    .B(_0593_));
 sg13g2_or3_1 _4962_ (.A(_0558_),
    .B(net1816),
    .C(_0586_),
    .X(_0595_));
 sg13g2_nand2_1 _4963_ (.Y(_0596_),
    .A(_0565_),
    .B(_0570_));
 sg13g2_o21ai_1 _4964_ (.B1(_0558_),
    .Y(_0597_),
    .A1(net1816),
    .A2(_0586_));
 sg13g2_nand3_1 _4965_ (.B(_0596_),
    .C(_0597_),
    .A(_0595_),
    .Y(_0598_));
 sg13g2_xnor2_1 _4966_ (.Y(_0599_),
    .A(net1955),
    .B(_0598_));
 sg13g2_nand2_1 _4967_ (.Y(_0600_),
    .A(_0565_),
    .B(_0568_));
 sg13g2_a21oi_1 _4968_ (.A1(_0559_),
    .A2(_0578_),
    .Y(_0601_),
    .B1(_0563_));
 sg13g2_o21ai_1 _4969_ (.B1(_0600_),
    .Y(_0602_),
    .A1(_0584_),
    .A2(_0601_));
 sg13g2_xnor2_1 _4970_ (.Y(_0603_),
    .A(net1956),
    .B(_0602_));
 sg13g2_and4_1 _4971_ (.A(_0590_),
    .B(_0594_),
    .C(_0599_),
    .D(_0603_),
    .X(_0604_));
 sg13g2_nand4_1 _4972_ (.B(_0594_),
    .C(_0599_),
    .A(_0590_),
    .Y(_0605_),
    .D(_0603_));
 sg13g2_nor2_2 _4973_ (.A(_0572_),
    .B(_0579_),
    .Y(_0606_));
 sg13g2_nand2b_1 _4974_ (.Y(_0607_),
    .B(_0578_),
    .A_N(_0572_));
 sg13g2_a21oi_2 _4975_ (.B1(_0582_),
    .Y(_0608_),
    .A2(_0607_),
    .A1(_0604_));
 sg13g2_nand3_1 _4976_ (.B(_0570_),
    .C(net1816),
    .A(_0566_),
    .Y(_0609_));
 sg13g2_xor2_1 _4977_ (.B(_0609_),
    .A(net1955),
    .X(_0610_));
 sg13g2_nand3_1 _4978_ (.B(_0569_),
    .C(_0579_),
    .A(_0566_),
    .Y(_0611_));
 sg13g2_xnor2_1 _4979_ (.Y(_0612_),
    .A(_0543_),
    .B(_0611_));
 sg13g2_nand3_1 _4980_ (.B(_0568_),
    .C(net1816),
    .A(_0566_),
    .Y(_0613_));
 sg13g2_xor2_1 _4981_ (.B(_0613_),
    .A(net1956),
    .X(_0614_));
 sg13g2_nand3_1 _4982_ (.B(_0567_),
    .C(net1816),
    .A(_0566_),
    .Y(_0615_));
 sg13g2_xor2_1 _4983_ (.B(_0615_),
    .A(_0548_),
    .X(_0616_));
 sg13g2_and4_1 _4984_ (.A(_0610_),
    .B(_0612_),
    .C(_0614_),
    .D(_0616_),
    .X(_0617_));
 sg13g2_nand4_1 _4985_ (.B(_0612_),
    .C(_0614_),
    .A(_0610_),
    .Y(_0618_),
    .D(_0616_));
 sg13g2_nor2_1 _4986_ (.A(_0573_),
    .B(_0618_),
    .Y(_0619_));
 sg13g2_nor2_1 _4987_ (.A(_0608_),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_nor3_1 _4988_ (.A(_0552_),
    .B(_0608_),
    .C(_0619_),
    .Y(_0621_));
 sg13g2_xor2_1 _4989_ (.B(_0620_),
    .A(_0552_),
    .X(_0622_));
 sg13g2_nand2_2 _4990_ (.Y(_0623_),
    .A(net1810),
    .B(net1796));
 sg13g2_nor2b_1 _4991_ (.A(net1810),
    .B_N(_0552_),
    .Y(_0624_));
 sg13g2_nor2_2 _4992_ (.A(_0621_),
    .B(_0624_),
    .Y(_0625_));
 sg13g2_or2_1 _4993_ (.X(_0626_),
    .B(_0624_),
    .A(_0621_));
 sg13g2_nand2_1 _4994_ (.Y(_0627_),
    .A(_0623_),
    .B(_0626_));
 sg13g2_nand2_1 _4995_ (.Y(_0628_),
    .A(_0622_),
    .B(_0627_));
 sg13g2_inv_1 _4996_ (.Y(_0629_),
    .A(_0628_));
 sg13g2_mux2_1 _4997_ (.A0(_0556_),
    .A1(_0557_),
    .S(net2051),
    .X(_0630_));
 sg13g2_nor2b_1 _4998_ (.A(_0623_),
    .B_N(net1955),
    .Y(_0631_));
 sg13g2_nand3_1 _4999_ (.B(net1810),
    .C(net1796),
    .A(net1955),
    .Y(_0632_));
 sg13g2_xnor2_1 _5000_ (.Y(_0633_),
    .A(net1954),
    .B(_0632_));
 sg13g2_nor3_2 _5001_ (.A(_0543_),
    .B(_0581_),
    .C(_0617_),
    .Y(_0634_));
 sg13g2_xnor2_1 _5002_ (.Y(_0635_),
    .A(_0532_),
    .B(_0634_));
 sg13g2_and2_1 _5003_ (.A(net2052),
    .B(_0554_),
    .X(_0636_));
 sg13g2_and2_1 _5004_ (.A(net2055),
    .B(_0553_),
    .X(_0637_));
 sg13g2_nor2_2 _5005_ (.A(_0636_),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_or2_2 _5006_ (.X(_0639_),
    .B(_0637_),
    .A(_0636_));
 sg13g2_nor2b_1 _5007_ (.A(_0623_),
    .B_N(_0548_),
    .Y(_0640_));
 sg13g2_nand3_1 _5008_ (.B(net1810),
    .C(net1796),
    .A(_0548_),
    .Y(_0641_));
 sg13g2_xnor2_1 _5009_ (.Y(_0642_),
    .A(_0639_),
    .B(_0641_));
 sg13g2_nor2b_1 _5010_ (.A(_0623_),
    .B_N(net1956),
    .Y(_0643_));
 sg13g2_nand3_1 _5011_ (.B(net1810),
    .C(net1796),
    .A(net1956),
    .Y(_0644_));
 sg13g2_mux2_2 _5012_ (.A0(_0561_),
    .A1(_0562_),
    .S(net2054),
    .X(_0645_));
 sg13g2_inv_1 _5013_ (.Y(_0646_),
    .A(_0645_));
 sg13g2_xnor2_1 _5014_ (.Y(_0647_),
    .A(_0644_),
    .B(_0645_));
 sg13g2_nor4_2 _5015_ (.A(_0633_),
    .B(_0635_),
    .C(_0642_),
    .Y(_0648_),
    .D(_0647_));
 sg13g2_or2_2 _5016_ (.X(_0649_),
    .B(_0648_),
    .A(_0628_));
 sg13g2_nor2_1 _5017_ (.A(_0532_),
    .B(_0649_),
    .Y(_0650_));
 sg13g2_and2_1 _5018_ (.A(_0542_),
    .B(_0573_),
    .X(_0651_));
 sg13g2_nor4_2 _5019_ (.A(_0543_),
    .B(net1810),
    .C(_0605_),
    .Y(_0652_),
    .D(_0606_));
 sg13g2_or4_1 _5020_ (.A(_0552_),
    .B(_0580_),
    .C(_0605_),
    .D(_0606_),
    .X(_0653_));
 sg13g2_a21oi_2 _5021_ (.B1(_0652_),
    .Y(_0654_),
    .A2(_0653_),
    .A1(_0593_));
 sg13g2_nor2_2 _5022_ (.A(_0651_),
    .B(_0654_),
    .Y(_0655_));
 sg13g2_or2_1 _5023_ (.X(_0656_),
    .B(_0654_),
    .A(_0651_));
 sg13g2_nand2_1 _5024_ (.Y(_0657_),
    .A(_0548_),
    .B(_0573_));
 sg13g2_nand2b_1 _5025_ (.Y(_0658_),
    .B(_0602_),
    .A_N(_0593_));
 sg13g2_nand2_1 _5026_ (.Y(_0659_),
    .A(_0581_),
    .B(_0589_));
 sg13g2_nor4_2 _5027_ (.A(_0605_),
    .B(_0606_),
    .C(_0658_),
    .Y(_0660_),
    .D(_0659_));
 sg13g2_a21oi_1 _5028_ (.A1(_0602_),
    .A2(_0652_),
    .Y(_0661_),
    .B1(_0589_));
 sg13g2_o21ai_1 _5029_ (.B1(_0657_),
    .Y(_0662_),
    .A1(_0660_),
    .A2(_0661_));
 sg13g2_nand2_1 _5030_ (.Y(_0663_),
    .A(net1956),
    .B(_0573_));
 sg13g2_xnor2_1 _5031_ (.Y(_0664_),
    .A(_0602_),
    .B(_0652_));
 sg13g2_and2_1 _5032_ (.A(_0663_),
    .B(_0664_),
    .X(_0665_));
 sg13g2_and3_1 _5033_ (.X(_0666_),
    .A(_0645_),
    .B(_0663_),
    .C(_0664_));
 sg13g2_a21oi_1 _5034_ (.A1(net1816),
    .A2(_0605_),
    .Y(_0667_),
    .B1(_0582_));
 sg13g2_nand2_1 _5035_ (.Y(_0668_),
    .A(net1955),
    .B(_0573_));
 sg13g2_inv_1 _5036_ (.Y(_0669_),
    .A(_0668_));
 sg13g2_xor2_1 _5037_ (.B(_0660_),
    .A(_0598_),
    .X(_0670_));
 sg13g2_xnor2_1 _5038_ (.Y(_0671_),
    .A(_0598_),
    .B(_0660_));
 sg13g2_nand2_1 _5039_ (.Y(_0672_),
    .A(_0668_),
    .B(_0671_));
 sg13g2_nand3b_1 _5040_ (.B(_0668_),
    .C(_0671_),
    .Y(_0673_),
    .A_N(_0630_));
 sg13g2_o21ai_1 _5041_ (.B1(net1954),
    .Y(_0674_),
    .A1(_0669_),
    .A2(_0670_));
 sg13g2_nor3_1 _5042_ (.A(_0532_),
    .B(_0651_),
    .C(_0654_),
    .Y(_0675_));
 sg13g2_a21oi_1 _5043_ (.A1(_0663_),
    .A2(_0664_),
    .Y(_0676_),
    .B1(_0645_));
 sg13g2_a221oi_1 _5044_ (.B2(_0674_),
    .C1(_0667_),
    .B1(_0673_),
    .A1(_0532_),
    .Y(_0677_),
    .A2(_0656_));
 sg13g2_xnor2_1 _5045_ (.Y(_0678_),
    .A(_0639_),
    .B(_0662_));
 sg13g2_nor3_1 _5046_ (.A(_0666_),
    .B(_0675_),
    .C(_0676_),
    .Y(_0679_));
 sg13g2_nand3_1 _5047_ (.B(_0678_),
    .C(_0679_),
    .A(_0677_),
    .Y(_0680_));
 sg13g2_and2_1 _5048_ (.A(_0622_),
    .B(_0623_),
    .X(_0681_));
 sg13g2_nand2_2 _5049_ (.Y(_0682_),
    .A(_0622_),
    .B(_0623_));
 sg13g2_xnor2_1 _5050_ (.Y(_0683_),
    .A(_0655_),
    .B(_0680_));
 sg13g2_nor4_1 _5051_ (.A(_0533_),
    .B(net1954),
    .C(_0639_),
    .D(_0645_),
    .Y(_0684_));
 sg13g2_inv_1 _5052_ (.Y(_0685_),
    .A(_0684_));
 sg13g2_nand3_1 _5053_ (.B(_0626_),
    .C(_0685_),
    .A(_0623_),
    .Y(_0686_));
 sg13g2_and2_1 _5054_ (.A(_0620_),
    .B(_0624_),
    .X(_0687_));
 sg13g2_a21oi_1 _5055_ (.A1(_0533_),
    .A2(_0687_),
    .Y(_0688_),
    .B1(_0686_));
 sg13g2_o21ai_1 _5056_ (.B1(_0688_),
    .Y(_0689_),
    .A1(_0682_),
    .A2(_0683_));
 sg13g2_nand2_2 _5057_ (.Y(_0690_),
    .A(_0655_),
    .B(_0686_));
 sg13g2_and2_1 _5058_ (.A(_0689_),
    .B(_0690_),
    .X(_0691_));
 sg13g2_nor2_2 _5059_ (.A(net2054),
    .B(_0650_),
    .Y(_0692_));
 sg13g2_a21oi_2 _5060_ (.B1(net2050),
    .Y(_0693_),
    .A2(_0690_),
    .A1(_0689_));
 sg13g2_nor2_2 _5061_ (.A(_0692_),
    .B(_0693_),
    .Y(_0694_));
 sg13g2_o21ai_1 _5062_ (.B1(net2176),
    .Y(_0695_),
    .A1(_0099_),
    .A2(net2059));
 sg13g2_a21oi_1 _5063_ (.A1(net2059),
    .A2(_0694_),
    .Y(_0696_),
    .B1(_0695_));
 sg13g2_nor2_1 _5064_ (.A(\game_logic_inst.should_transpose ),
    .B(net1809),
    .Y(_0697_));
 sg13g2_nand2b_1 _5065_ (.Y(_0698_),
    .B(net1808),
    .A_N(\game_logic_inst.should_transpose ));
 sg13g2_mux4_1 _5066_ (.S0(\game_logic_inst.lfsr_shift[0] ),
    .A0(\game_logic_inst.lfsr_value[3] ),
    .A1(\game_logic_inst.lfsr_value[7] ),
    .A2(\game_logic_inst.lfsr_value[11] ),
    .A3(\game_logic_inst.lfsr_value[15] ),
    .S1(\game_logic_inst.lfsr_shift[1] ),
    .X(_0699_));
 sg13g2_inv_1 _5067_ (.Y(_0700_),
    .A(_0699_));
 sg13g2_mux4_1 _5068_ (.S0(\game_logic_inst.lfsr_shift[0] ),
    .A0(\game_logic_inst.lfsr_value[2] ),
    .A1(\game_logic_inst.lfsr_value[6] ),
    .A2(\game_logic_inst.lfsr_value[10] ),
    .A3(\game_logic_inst.lfsr_value[14] ),
    .S1(\game_logic_inst.lfsr_shift[1] ),
    .X(_0701_));
 sg13g2_inv_4 _5069_ (.A(net2035),
    .Y(_0702_));
 sg13g2_mux4_1 _5070_ (.S0(\game_logic_inst.lfsr_shift[0] ),
    .A0(\game_logic_inst.lfsr_value[1] ),
    .A1(\game_logic_inst.lfsr_value[5] ),
    .A2(\game_logic_inst.lfsr_value[9] ),
    .A3(\game_logic_inst.lfsr_value[13] ),
    .S1(\game_logic_inst.lfsr_shift[1] ),
    .X(_0703_));
 sg13g2_mux4_1 _5071_ (.S0(\game_logic_inst.lfsr_shift[0] ),
    .A0(\game_logic_inst.lfsr_value[0] ),
    .A1(\game_logic_inst.lfsr_value[4] ),
    .A2(\game_logic_inst.lfsr_value[8] ),
    .A3(\game_logic_inst.lfsr_value[12] ),
    .S1(\game_logic_inst.lfsr_shift[1] ),
    .X(_0704_));
 sg13g2_nand2_2 _5072_ (.Y(_0705_),
    .A(_0703_),
    .B(_0704_));
 sg13g2_nor4_2 _5073_ (.A(\debug_controller_inst.grid_in[28] ),
    .B(\debug_controller_inst.grid_in[29] ),
    .C(\debug_controller_inst.grid_in[30] ),
    .Y(_0706_),
    .D(\debug_controller_inst.grid_in[31] ));
 sg13g2_or2_2 _5074_ (.X(_0707_),
    .B(_0704_),
    .A(_0703_));
 sg13g2_nor4_2 _5075_ (.A(\debug_controller_inst.grid_in[16] ),
    .B(\debug_controller_inst.grid_in[17] ),
    .C(\debug_controller_inst.grid_in[18] ),
    .Y(_0708_),
    .D(\debug_controller_inst.grid_in[19] ));
 sg13g2_nor2_1 _5076_ (.A(_0707_),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_nand2b_2 _5077_ (.Y(_0710_),
    .B(_0704_),
    .A_N(_0703_));
 sg13g2_nor4_1 _5078_ (.A(\debug_controller_inst.grid_in[20] ),
    .B(\debug_controller_inst.grid_in[21] ),
    .C(\debug_controller_inst.grid_in[22] ),
    .D(\debug_controller_inst.grid_in[23] ),
    .Y(_0711_));
 sg13g2_nand2b_2 _5079_ (.Y(_0712_),
    .B(_0703_),
    .A_N(_0704_));
 sg13g2_nor4_1 _5080_ (.A(\debug_controller_inst.grid_in[24] ),
    .B(\debug_controller_inst.grid_in[25] ),
    .C(\debug_controller_inst.grid_in[26] ),
    .D(\debug_controller_inst.grid_in[27] ),
    .Y(_0713_));
 sg13g2_nor2_1 _5081_ (.A(_0712_),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_o21ai_1 _5082_ (.B1(net2035),
    .Y(_0715_),
    .A1(_0710_),
    .A2(_0711_));
 sg13g2_nor3_1 _5083_ (.A(_0709_),
    .B(_0714_),
    .C(_0715_),
    .Y(_0716_));
 sg13g2_o21ai_1 _5084_ (.B1(_0716_),
    .Y(_0717_),
    .A1(_0705_),
    .A2(_0706_));
 sg13g2_nor4_2 _5085_ (.A(\debug_controller_inst.grid_in[12] ),
    .B(\debug_controller_inst.grid_in[13] ),
    .C(\debug_controller_inst.grid_in[14] ),
    .Y(_0718_),
    .D(\debug_controller_inst.grid_in[15] ));
 sg13g2_o21ai_1 _5086_ (.B1(_0702_),
    .Y(_0719_),
    .A1(_0705_),
    .A2(_0718_));
 sg13g2_nor4_1 _5087_ (.A(\debug_controller_inst.grid_in[0] ),
    .B(\debug_controller_inst.grid_in[1] ),
    .C(\debug_controller_inst.grid_in[2] ),
    .D(\debug_controller_inst.grid_in[3] ),
    .Y(_0720_));
 sg13g2_nor2_1 _5088_ (.A(_0707_),
    .B(_0720_),
    .Y(_0721_));
 sg13g2_nor4_1 _5089_ (.A(\debug_controller_inst.grid_in[8] ),
    .B(\debug_controller_inst.grid_in[9] ),
    .C(\debug_controller_inst.grid_in[10] ),
    .D(\debug_controller_inst.grid_in[11] ),
    .Y(_0722_));
 sg13g2_nor2_1 _5090_ (.A(_0712_),
    .B(_0722_),
    .Y(_0723_));
 sg13g2_nor4_2 _5091_ (.A(\debug_controller_inst.grid_in[4] ),
    .B(\debug_controller_inst.grid_in[5] ),
    .C(\debug_controller_inst.grid_in[6] ),
    .Y(_0724_),
    .D(\debug_controller_inst.grid_in[7] ));
 sg13g2_nor2_1 _5092_ (.A(_0710_),
    .B(_0724_),
    .Y(_0725_));
 sg13g2_nor4_1 _5093_ (.A(_0719_),
    .B(_0721_),
    .C(_0723_),
    .D(_0725_),
    .Y(_0726_));
 sg13g2_nor2_1 _5094_ (.A(_0699_),
    .B(_0726_),
    .Y(_0727_));
 sg13g2_nor4_1 _5095_ (.A(\debug_controller_inst.grid_in[32] ),
    .B(\debug_controller_inst.grid_in[33] ),
    .C(\debug_controller_inst.grid_in[34] ),
    .D(\debug_controller_inst.grid_in[35] ),
    .Y(_0728_));
 sg13g2_o21ai_1 _5096_ (.B1(_0702_),
    .Y(_0729_),
    .A1(_0707_),
    .A2(_0728_));
 sg13g2_nor4_1 _5097_ (.A(\debug_controller_inst.grid_in[40] ),
    .B(\debug_controller_inst.grid_in[41] ),
    .C(\debug_controller_inst.grid_in[42] ),
    .D(\debug_controller_inst.grid_in[43] ),
    .Y(_0730_));
 sg13g2_nor2_1 _5098_ (.A(_0712_),
    .B(_0730_),
    .Y(_0731_));
 sg13g2_nor4_1 _5099_ (.A(\debug_controller_inst.grid_in[36] ),
    .B(\debug_controller_inst.grid_in[37] ),
    .C(\debug_controller_inst.grid_in[38] ),
    .D(\debug_controller_inst.grid_in[39] ),
    .Y(_0732_));
 sg13g2_nor2_1 _5100_ (.A(_0710_),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_nor4_1 _5101_ (.A(\debug_controller_inst.grid_in[44] ),
    .B(\debug_controller_inst.grid_in[45] ),
    .C(\debug_controller_inst.grid_in[46] ),
    .D(\debug_controller_inst.grid_in[47] ),
    .Y(_0734_));
 sg13g2_nor2_1 _5102_ (.A(_0705_),
    .B(_0734_),
    .Y(_0735_));
 sg13g2_nor4_1 _5103_ (.A(_0729_),
    .B(_0731_),
    .C(_0733_),
    .D(_0735_),
    .Y(_0736_));
 sg13g2_nor3_1 _5104_ (.A(\debug_controller_inst.grid_in[52] ),
    .B(\debug_controller_inst.grid_in[53] ),
    .C(\debug_controller_inst.grid_in[54] ),
    .Y(_0737_));
 sg13g2_a21oi_1 _5105_ (.A1(_4034_),
    .A2(_0737_),
    .Y(_0738_),
    .B1(_0710_));
 sg13g2_nor4_1 _5106_ (.A(\debug_controller_inst.grid_in[60] ),
    .B(\debug_controller_inst.grid_in[61] ),
    .C(\debug_controller_inst.grid_in[62] ),
    .D(\debug_controller_inst.grid_in[63] ),
    .Y(_0739_));
 sg13g2_nor2_1 _5107_ (.A(_0705_),
    .B(_0739_),
    .Y(_0740_));
 sg13g2_nor4_2 _5108_ (.A(\debug_controller_inst.grid_in[48] ),
    .B(\debug_controller_inst.grid_in[49] ),
    .C(\debug_controller_inst.grid_in[50] ),
    .Y(_0741_),
    .D(\debug_controller_inst.grid_in[51] ));
 sg13g2_nor4_1 _5109_ (.A(\debug_controller_inst.grid_in[56] ),
    .B(\debug_controller_inst.grid_in[57] ),
    .C(\debug_controller_inst.grid_in[58] ),
    .D(\debug_controller_inst.grid_in[59] ),
    .Y(_0742_));
 sg13g2_nor2_1 _5110_ (.A(_0712_),
    .B(_0742_),
    .Y(_0743_));
 sg13g2_o21ai_1 _5111_ (.B1(net2035),
    .Y(_0744_),
    .A1(_0707_),
    .A2(_0741_));
 sg13g2_nor4_1 _5112_ (.A(_0738_),
    .B(_0740_),
    .C(_0743_),
    .D(_0744_),
    .Y(_0745_));
 sg13g2_nor3_1 _5113_ (.A(_0700_),
    .B(_0736_),
    .C(_0745_),
    .Y(_0746_));
 sg13g2_nor2_2 _5114_ (.A(\game_logic_inst.add_new_tiles[1] ),
    .B(\game_logic_inst.add_new_tiles[0] ),
    .Y(_0747_));
 sg13g2_a21oi_2 _5115_ (.B1(_0746_),
    .Y(_0748_),
    .A2(_0727_),
    .A1(_0717_));
 sg13g2_nand2b_1 _5116_ (.Y(_0749_),
    .B(_0748_),
    .A_N(_0747_));
 sg13g2_inv_1 _5117_ (.Y(_0750_),
    .A(_0749_));
 sg13g2_nor2_1 _5118_ (.A(_0699_),
    .B(_0749_),
    .Y(_0751_));
 sg13g2_nor2_2 _5119_ (.A(net2035),
    .B(_0707_),
    .Y(_0752_));
 sg13g2_and2_1 _5120_ (.A(_0751_),
    .B(_0752_),
    .X(_0753_));
 sg13g2_nor3_1 _5121_ (.A(net2176),
    .B(_4056_),
    .C(_0753_),
    .Y(_0754_));
 sg13g2_nor3_1 _5122_ (.A(_0696_),
    .B(net1791),
    .C(_0754_),
    .Y(_0755_));
 sg13g2_o21ai_1 _5123_ (.B1(net2170),
    .Y(_0756_),
    .A1(_0099_),
    .A2(net1794));
 sg13g2_nor2_2 _5124_ (.A(net2301),
    .B(_0520_),
    .Y(_0757_));
 sg13g2_o21ai_1 _5125_ (.B1(_0757_),
    .Y(_0758_),
    .A1(_0755_),
    .A2(_0756_));
 sg13g2_a21oi_1 _5126_ (.A1(net2102),
    .A2(net942),
    .Y(_0759_),
    .B1(_0758_));
 sg13g2_a21o_1 _5127_ (.A2(_0520_),
    .A1(net2149),
    .B1(_0759_),
    .X(_0003_));
 sg13g2_nor2_1 _5128_ (.A(_3986_),
    .B(net1791),
    .Y(_0760_));
 sg13g2_nand2_1 _5129_ (.Y(_0761_),
    .A(net2178),
    .B(net1795));
 sg13g2_or3_1 _5130_ (.A(_0100_),
    .B(net1791),
    .C(_0753_),
    .X(_0762_));
 sg13g2_nor2_1 _5131_ (.A(_0646_),
    .B(_0649_),
    .Y(_0763_));
 sg13g2_nand2_1 _5132_ (.Y(_0764_),
    .A(_0665_),
    .B(_0686_));
 sg13g2_o21ai_1 _5133_ (.B1(_0665_),
    .Y(_0765_),
    .A1(_0655_),
    .A2(_0680_));
 sg13g2_nor2_1 _5134_ (.A(_0655_),
    .B(_0665_),
    .Y(_0766_));
 sg13g2_and4_1 _5135_ (.A(_0677_),
    .B(_0678_),
    .C(_0679_),
    .D(_0766_),
    .X(_0767_));
 sg13g2_nor2_1 _5136_ (.A(_0682_),
    .B(_0767_),
    .Y(_0768_));
 sg13g2_a21o_1 _5137_ (.A2(_0687_),
    .A1(_0645_),
    .B1(_0686_),
    .X(_0769_));
 sg13g2_a21o_1 _5138_ (.A2(_0768_),
    .A1(_0765_),
    .B1(_0769_),
    .X(_0770_));
 sg13g2_and2_1 _5139_ (.A(_0764_),
    .B(_0770_),
    .X(_0771_));
 sg13g2_nor2_1 _5140_ (.A(net2054),
    .B(_0763_),
    .Y(_0772_));
 sg13g2_a21oi_1 _5141_ (.A1(_0764_),
    .A2(_0770_),
    .Y(_0773_),
    .B1(net2050));
 sg13g2_nor2_2 _5142_ (.A(_0772_),
    .B(_0773_),
    .Y(_0774_));
 sg13g2_nor2_1 _5143_ (.A(_0100_),
    .B(net2059),
    .Y(_0775_));
 sg13g2_a21oi_1 _5144_ (.A1(net2059),
    .A2(_0774_),
    .Y(_0776_),
    .B1(_0775_));
 sg13g2_a22oi_1 _5145_ (.Y(_0777_),
    .B1(_0776_),
    .B2(net2176),
    .A2(_0762_),
    .A1(net1759));
 sg13g2_o21ai_1 _5146_ (.B1(net2170),
    .Y(_0778_),
    .A1(net873),
    .A2(net1794));
 sg13g2_o21ai_1 _5147_ (.B1(_0757_),
    .Y(_0779_),
    .A1(_0777_),
    .A2(_0778_));
 sg13g2_a21oi_1 _5148_ (.A1(net2102),
    .A2(net873),
    .Y(_0780_),
    .B1(_0779_));
 sg13g2_a21o_1 _5149_ (.A2(_0520_),
    .A1(net2145),
    .B1(_0780_),
    .X(_0014_));
 sg13g2_or3_1 _5150_ (.A(_0101_),
    .B(net1792),
    .C(_0753_),
    .X(_0781_));
 sg13g2_nor2_1 _5151_ (.A(_0638_),
    .B(_0649_),
    .Y(_0782_));
 sg13g2_a21oi_1 _5152_ (.A1(_0662_),
    .A2(_0767_),
    .Y(_0783_),
    .B1(_0682_));
 sg13g2_o21ai_1 _5153_ (.B1(_0662_),
    .Y(_0784_),
    .A1(_0686_),
    .A2(_0783_));
 sg13g2_a22oi_1 _5154_ (.Y(_0785_),
    .B1(_0767_),
    .B2(_0783_),
    .A2(_0687_),
    .A1(_0639_));
 sg13g2_nand2_1 _5155_ (.Y(_0786_),
    .A(_0784_),
    .B(_0785_));
 sg13g2_mux2_2 _5156_ (.A0(_0782_),
    .A1(_0786_),
    .S(net2055),
    .X(_0787_));
 sg13g2_nor2_1 _5157_ (.A(_0101_),
    .B(net2059),
    .Y(_0788_));
 sg13g2_a21oi_1 _5158_ (.A1(net2059),
    .A2(_0787_),
    .Y(_0789_),
    .B1(_0788_));
 sg13g2_a22oi_1 _5159_ (.Y(_0790_),
    .B1(_0789_),
    .B2(net2178),
    .A2(_0781_),
    .A1(net1760));
 sg13g2_o21ai_1 _5160_ (.B1(net2172),
    .Y(_0791_),
    .A1(net870),
    .A2(net1795));
 sg13g2_o21ai_1 _5161_ (.B1(_0757_),
    .Y(_0792_),
    .A1(_0790_),
    .A2(_0791_));
 sg13g2_a21oi_1 _5162_ (.A1(net2099),
    .A2(net870),
    .Y(_0793_),
    .B1(_0792_));
 sg13g2_a21o_1 _5163_ (.A2(_0520_),
    .A1(net2143),
    .B1(_0793_),
    .X(_0025_));
 sg13g2_or3_1 _5164_ (.A(_0102_),
    .B(net1791),
    .C(_0753_),
    .X(_0794_));
 sg13g2_o21ai_1 _5165_ (.B1(_0672_),
    .Y(_0795_),
    .A1(_0686_),
    .A2(_0783_));
 sg13g2_nor2_1 _5166_ (.A(_0672_),
    .B(_0682_),
    .Y(_0796_));
 sg13g2_nand3_1 _5167_ (.B(_0767_),
    .C(_0796_),
    .A(_0662_),
    .Y(_0797_));
 sg13g2_nand2_1 _5168_ (.Y(_0798_),
    .A(net1954),
    .B(_0687_));
 sg13g2_and2_1 _5169_ (.A(_0797_),
    .B(_0798_),
    .X(_0799_));
 sg13g2_a21o_1 _5170_ (.A2(_0799_),
    .A1(_0795_),
    .B1(net2051),
    .X(_0800_));
 sg13g2_nor2b_1 _5171_ (.A(_0649_),
    .B_N(net1954),
    .Y(_0801_));
 sg13g2_nand2_1 _5172_ (.Y(_0802_),
    .A(net2051),
    .B(_0801_));
 sg13g2_and2_2 _5173_ (.A(_0800_),
    .B(_0802_),
    .X(_0803_));
 sg13g2_mux2_1 _5174_ (.A0(_0102_),
    .A1(_0803_),
    .S(net2059),
    .X(_0804_));
 sg13g2_a22oi_1 _5175_ (.Y(_0805_),
    .B1(_0804_),
    .B2(net2176),
    .A2(_0794_),
    .A1(net1759));
 sg13g2_o21ai_1 _5176_ (.B1(net2170),
    .Y(_0806_),
    .A1(_0102_),
    .A2(net1794));
 sg13g2_o21ai_1 _5177_ (.B1(_0757_),
    .Y(_0807_),
    .A1(_0805_),
    .A2(_0806_));
 sg13g2_a21oi_1 _5178_ (.A1(net2102),
    .A2(net905),
    .Y(_0808_),
    .B1(_0807_));
 sg13g2_a21o_1 _5179_ (.A2(_0520_),
    .A1(net2142),
    .B1(net906),
    .X(_0036_));
 sg13g2_xnor2_1 _5180_ (.Y(_0809_),
    .A(\debug_controller_inst.grid_out_addr[3] ),
    .B(_0518_));
 sg13g2_nand2_2 _5181_ (.Y(_0810_),
    .A(\debug_controller_inst.grid_out_valid ),
    .B(_0809_));
 sg13g2_nor2b_1 _5182_ (.A(net2139),
    .B_N(net2140),
    .Y(_0811_));
 sg13g2_nand2b_1 _5183_ (.Y(_0812_),
    .B(net2140),
    .A_N(net2139));
 sg13g2_nor3_2 _5184_ (.A(net2137),
    .B(_0810_),
    .C(_0812_),
    .Y(_0813_));
 sg13g2_nand2b_1 _5185_ (.Y(_0814_),
    .B(_0617_),
    .A_N(_0552_));
 sg13g2_nor3_2 _5186_ (.A(_0538_),
    .B(_0552_),
    .C(net1796),
    .Y(_0815_));
 sg13g2_nor4_2 _5187_ (.A(_0538_),
    .B(_0552_),
    .C(_0613_),
    .Y(_0816_),
    .D(net1796));
 sg13g2_and2_1 _5188_ (.A(_0567_),
    .B(_0816_),
    .X(_0817_));
 sg13g2_xnor2_1 _5189_ (.Y(_0818_),
    .A(_0615_),
    .B(_0816_));
 sg13g2_a221oi_1 _5190_ (.B2(_0607_),
    .C1(_0582_),
    .B1(_0604_),
    .A1(_0545_),
    .Y(_0819_),
    .A2(_0547_));
 sg13g2_or2_1 _5191_ (.X(_0820_),
    .B(_0819_),
    .A(_0818_));
 sg13g2_o21ai_1 _5192_ (.B1(_0638_),
    .Y(_0821_),
    .A1(_0818_),
    .A2(_0819_));
 sg13g2_or3_1 _5193_ (.A(_0638_),
    .B(_0818_),
    .C(_0819_),
    .X(_0822_));
 sg13g2_and3_1 _5194_ (.X(_0823_),
    .A(_0814_),
    .B(_0821_),
    .C(_0822_));
 sg13g2_nand2_1 _5195_ (.Y(_0824_),
    .A(_0571_),
    .B(_0817_));
 sg13g2_a21oi_1 _5196_ (.A1(_0567_),
    .A2(_0816_),
    .Y(_0825_),
    .B1(_0609_));
 sg13g2_a21oi_1 _5197_ (.A1(net1955),
    .A2(_0608_),
    .Y(_0826_),
    .B1(_0825_));
 sg13g2_a221oi_1 _5198_ (.B2(_0571_),
    .C1(_0825_),
    .B1(_0817_),
    .A1(net1955),
    .Y(_0827_),
    .A2(_0608_));
 sg13g2_nand2_1 _5199_ (.Y(_0828_),
    .A(_0824_),
    .B(_0826_));
 sg13g2_xor2_1 _5200_ (.B(_0827_),
    .A(net1954),
    .X(_0829_));
 sg13g2_a221oi_1 _5201_ (.B2(_0607_),
    .C1(_0582_),
    .B1(_0604_),
    .A1(_0539_),
    .Y(_0830_),
    .A2(_0541_));
 sg13g2_a21oi_1 _5202_ (.A1(_0611_),
    .A2(_0814_),
    .Y(_0831_),
    .B1(_0815_));
 sg13g2_a21o_1 _5203_ (.A2(_0814_),
    .A1(_0611_),
    .B1(_0815_),
    .X(_0832_));
 sg13g2_nand2b_1 _5204_ (.Y(_0833_),
    .B(_0832_),
    .A_N(_0830_));
 sg13g2_nand3b_1 _5205_ (.B(_0832_),
    .C(_0532_),
    .Y(_0834_),
    .A_N(_0830_));
 sg13g2_o21ai_1 _5206_ (.B1(_0533_),
    .Y(_0835_),
    .A1(_0830_),
    .A2(_0831_));
 sg13g2_nor2b_1 _5207_ (.A(_0582_),
    .B_N(net1956),
    .Y(_0836_));
 sg13g2_o21ai_1 _5208_ (.B1(_0836_),
    .Y(_0837_),
    .A1(_0605_),
    .A2(_0606_));
 sg13g2_xor2_1 _5209_ (.B(_0815_),
    .A(_0613_),
    .X(_0838_));
 sg13g2_nand2_2 _5210_ (.Y(_0839_),
    .A(_0837_),
    .B(_0838_));
 sg13g2_inv_1 _5211_ (.Y(_0840_),
    .A(_0839_));
 sg13g2_nand3_1 _5212_ (.B(_0837_),
    .C(_0838_),
    .A(_0646_),
    .Y(_0841_));
 sg13g2_a21o_1 _5213_ (.A2(_0838_),
    .A1(_0837_),
    .B1(_0646_),
    .X(_0842_));
 sg13g2_a22oi_1 _5214_ (.Y(_0843_),
    .B1(_0841_),
    .B2(_0842_),
    .A2(_0835_),
    .A1(_0834_));
 sg13g2_nand3_1 _5215_ (.B(_0829_),
    .C(_0843_),
    .A(_0823_),
    .Y(_0844_));
 sg13g2_and2_1 _5216_ (.A(_0625_),
    .B(_0844_),
    .X(_0845_));
 sg13g2_nand2_1 _5217_ (.Y(_0846_),
    .A(_0634_),
    .B(_0648_));
 sg13g2_xor2_1 _5218_ (.B(_0648_),
    .A(_0634_),
    .X(_0847_));
 sg13g2_a22oi_1 _5219_ (.Y(_0848_),
    .B1(_0847_),
    .B2(_0629_),
    .A2(_0845_),
    .A1(_0533_));
 sg13g2_and2_1 _5220_ (.A(_0680_),
    .B(_0681_),
    .X(_0849_));
 sg13g2_a21oi_1 _5221_ (.A1(_0626_),
    .A2(_0682_),
    .Y(_0850_),
    .B1(_0684_));
 sg13g2_nand4_1 _5222_ (.B(_0678_),
    .C(_0679_),
    .A(_0677_),
    .Y(_0851_),
    .D(_0681_));
 sg13g2_nand3b_1 _5223_ (.B(_0850_),
    .C(_0851_),
    .Y(_0852_),
    .A_N(_0845_));
 sg13g2_nand4_1 _5224_ (.B(_0823_),
    .C(_0829_),
    .A(_0625_),
    .Y(_0853_),
    .D(_0843_));
 sg13g2_nor2_1 _5225_ (.A(_0833_),
    .B(_0853_),
    .Y(_0854_));
 sg13g2_a221oi_1 _5226_ (.B2(_0833_),
    .C1(_0854_),
    .B1(_0852_),
    .A1(_0533_),
    .Y(_0855_),
    .A2(_0849_));
 sg13g2_mux2_2 _5227_ (.A0(_0848_),
    .A1(_0855_),
    .S(net2054),
    .X(_0856_));
 sg13g2_nor2b_1 _5228_ (.A(_0856_),
    .B_N(net2058),
    .Y(_0857_));
 sg13g2_o21ai_1 _5229_ (.B1(net1765),
    .Y(_0858_),
    .A1(_0103_),
    .A2(net2058));
 sg13g2_and2_1 _5230_ (.A(\game_logic_inst.should_transpose ),
    .B(net1808),
    .X(_0859_));
 sg13g2_nor2_1 _5231_ (.A(net2035),
    .B(_0710_),
    .Y(_0860_));
 sg13g2_nor3_2 _5232_ (.A(net1809),
    .B(_0699_),
    .C(_0749_),
    .Y(_0861_));
 sg13g2_nand2_2 _5233_ (.Y(_0862_),
    .A(_0860_),
    .B(net1758));
 sg13g2_nor2_2 _5234_ (.A(\game_logic_inst.should_transpose ),
    .B(net2176),
    .Y(_0863_));
 sg13g2_or2_1 _5235_ (.X(_0864_),
    .B(net2176),
    .A(\game_logic_inst.should_transpose ));
 sg13g2_nand2_1 _5236_ (.Y(_0865_),
    .A(net1808),
    .B(net2033));
 sg13g2_and2_1 _5237_ (.A(_0103_),
    .B(net1778),
    .X(_0866_));
 sg13g2_a22oi_1 _5238_ (.Y(_0867_),
    .B1(_0862_),
    .B2(_0866_),
    .A2(net1785),
    .A1(_0104_));
 sg13g2_o21ai_1 _5239_ (.B1(_0867_),
    .Y(_0868_),
    .A1(_0857_),
    .A2(_0858_));
 sg13g2_nand2_1 _5240_ (.Y(_0869_),
    .A(net2165),
    .B(_0868_));
 sg13g2_nand2b_2 _5241_ (.Y(_0870_),
    .B(net2311),
    .A_N(_0813_));
 sg13g2_a21oi_1 _5242_ (.A1(net2098),
    .A2(net878),
    .Y(_0871_),
    .B1(_0870_));
 sg13g2_a22oi_1 _5243_ (.Y(_0872_),
    .B1(_0869_),
    .B2(_0871_),
    .A2(_0813_),
    .A1(net2148));
 sg13g2_inv_1 _5244_ (.Y(_0047_),
    .A(net879));
 sg13g2_nand3_1 _5245_ (.B(_0634_),
    .C(_0648_),
    .A(net1956),
    .Y(_0873_));
 sg13g2_nand4_1 _5246_ (.B(net1796),
    .C(_0622_),
    .A(net1810),
    .Y(_0874_),
    .D(_0873_));
 sg13g2_nand4_1 _5247_ (.B(_0685_),
    .C(_0853_),
    .A(_0627_),
    .Y(_0875_),
    .D(_0874_));
 sg13g2_nor2_1 _5248_ (.A(_0846_),
    .B(_0874_),
    .Y(_0876_));
 sg13g2_a221oi_1 _5249_ (.B2(_0643_),
    .C1(_0876_),
    .B1(_0875_),
    .A1(_0645_),
    .Y(_0877_),
    .A2(_0845_));
 sg13g2_or2_1 _5250_ (.X(_0878_),
    .B(_0877_),
    .A(net2054));
 sg13g2_nand4_1 _5251_ (.B(_0829_),
    .C(_0833_),
    .A(_0823_),
    .Y(_0879_),
    .D(_0843_));
 sg13g2_o21ai_1 _5252_ (.B1(_0625_),
    .Y(_0880_),
    .A1(_0840_),
    .A2(_0879_));
 sg13g2_nand3_1 _5253_ (.B(_0851_),
    .C(_0880_),
    .A(_0850_),
    .Y(_0881_));
 sg13g2_nor2_1 _5254_ (.A(_0879_),
    .B(_0880_),
    .Y(_0882_));
 sg13g2_a221oi_1 _5255_ (.B2(_0839_),
    .C1(_0882_),
    .B1(_0881_),
    .A1(_0645_),
    .Y(_0883_),
    .A2(_0849_));
 sg13g2_o21ai_1 _5256_ (.B1(_0878_),
    .Y(_0884_),
    .A1(net2050),
    .A2(_0883_));
 sg13g2_o21ai_1 _5257_ (.B1(net1765),
    .Y(_0885_),
    .A1(_0105_),
    .A2(net2058));
 sg13g2_a21oi_1 _5258_ (.A1(net2058),
    .A2(_0884_),
    .Y(_0886_),
    .B1(_0885_));
 sg13g2_a22oi_1 _5259_ (.Y(_0887_),
    .B1(net1778),
    .B2(net900),
    .A2(net1785),
    .A1(_0106_));
 sg13g2_nor2_1 _5260_ (.A(net1809),
    .B(net2033),
    .Y(_0888_));
 sg13g2_o21ai_1 _5261_ (.B1(_0887_),
    .Y(_0889_),
    .A1(_0862_),
    .A2(net2032));
 sg13g2_o21ai_1 _5262_ (.B1(net2165),
    .Y(_0890_),
    .A1(_0886_),
    .A2(_0889_));
 sg13g2_a21oi_1 _5263_ (.A1(net2098),
    .A2(net900),
    .Y(_0891_),
    .B1(_0870_));
 sg13g2_a22oi_1 _5264_ (.Y(_0892_),
    .B1(_0890_),
    .B2(_0891_),
    .A2(_0813_),
    .A1(net2145));
 sg13g2_inv_1 _5265_ (.Y(_0058_),
    .A(net901));
 sg13g2_nand4_1 _5266_ (.B(_0634_),
    .C(_0640_),
    .A(net1956),
    .Y(_0893_),
    .D(_0648_));
 sg13g2_nand4_1 _5267_ (.B(net1796),
    .C(_0622_),
    .A(net1810),
    .Y(_0894_),
    .D(_0893_));
 sg13g2_nor2_1 _5268_ (.A(_0873_),
    .B(_0894_),
    .Y(_0895_));
 sg13g2_a221oi_1 _5269_ (.B2(_0640_),
    .C1(_0895_),
    .B1(_0875_),
    .A1(_0639_),
    .Y(_0896_),
    .A2(_0845_));
 sg13g2_nand2_1 _5270_ (.Y(_0897_),
    .A(_0820_),
    .B(_0839_));
 sg13g2_o21ai_1 _5271_ (.B1(_0625_),
    .Y(_0898_),
    .A1(_0879_),
    .A2(_0897_));
 sg13g2_nand3_1 _5272_ (.B(_0851_),
    .C(_0898_),
    .A(_0850_),
    .Y(_0899_));
 sg13g2_nor3_1 _5273_ (.A(_0840_),
    .B(_0879_),
    .C(_0898_),
    .Y(_0900_));
 sg13g2_a221oi_1 _5274_ (.B2(_0820_),
    .C1(_0900_),
    .B1(_0881_),
    .A1(_0639_),
    .Y(_0901_),
    .A2(_0849_));
 sg13g2_mux2_2 _5275_ (.A0(_0896_),
    .A1(_0901_),
    .S(net2054),
    .X(_0902_));
 sg13g2_inv_1 _5276_ (.Y(_0903_),
    .A(_0902_));
 sg13g2_o21ai_1 _5277_ (.B1(net1765),
    .Y(_0904_),
    .A1(_0107_),
    .A2(net2058));
 sg13g2_a21oi_1 _5278_ (.A1(net2058),
    .A2(_0903_),
    .Y(_0905_),
    .B1(_0904_));
 sg13g2_a22oi_1 _5279_ (.Y(_0906_),
    .B1(net1778),
    .B2(_0107_),
    .A2(net1785),
    .A1(_0108_));
 sg13g2_o21ai_1 _5280_ (.B1(_0906_),
    .Y(_0907_),
    .A1(_0862_),
    .A2(net2032));
 sg13g2_o21ai_1 _5281_ (.B1(net2164),
    .Y(_0908_),
    .A1(_0905_),
    .A2(_0907_));
 sg13g2_a21oi_1 _5282_ (.A1(net2097),
    .A2(net947),
    .Y(_0909_),
    .B1(_0870_));
 sg13g2_a22oi_1 _5283_ (.Y(_0910_),
    .B1(_0908_),
    .B2(_0909_),
    .A2(_0813_),
    .A1(net2143));
 sg13g2_inv_1 _5284_ (.Y(_0063_),
    .A(net948));
 sg13g2_nand4_1 _5285_ (.B(_0685_),
    .C(_0853_),
    .A(_0627_),
    .Y(_0911_),
    .D(_0894_));
 sg13g2_nor2_1 _5286_ (.A(net1955),
    .B(_0893_),
    .Y(_0912_));
 sg13g2_a221oi_1 _5287_ (.B2(_0631_),
    .C1(_0912_),
    .B1(_0911_),
    .A1(net1954),
    .Y(_0913_),
    .A2(_0845_));
 sg13g2_or2_1 _5288_ (.X(_0914_),
    .B(_0913_),
    .A(net2054));
 sg13g2_nor4_1 _5289_ (.A(_0626_),
    .B(_0828_),
    .C(_0879_),
    .D(_0897_),
    .Y(_0915_));
 sg13g2_a221oi_1 _5290_ (.B2(_0828_),
    .C1(_0915_),
    .B1(_0899_),
    .A1(net1954),
    .Y(_0916_),
    .A2(_0849_));
 sg13g2_o21ai_1 _5291_ (.B1(_0914_),
    .Y(_0917_),
    .A1(net2050),
    .A2(_0916_));
 sg13g2_o21ai_1 _5292_ (.B1(net1765),
    .Y(_0918_),
    .A1(net865),
    .A2(net2058));
 sg13g2_a21oi_1 _5293_ (.A1(net2058),
    .A2(_0917_),
    .Y(_0919_),
    .B1(_0918_));
 sg13g2_a22oi_1 _5294_ (.Y(_0920_),
    .B1(net1777),
    .B2(net865),
    .A2(net1785),
    .A1(_0110_));
 sg13g2_o21ai_1 _5295_ (.B1(_0920_),
    .Y(_0921_),
    .A1(_0862_),
    .A2(net2032));
 sg13g2_o21ai_1 _5296_ (.B1(net2164),
    .Y(_0922_),
    .A1(_0919_),
    .A2(_0921_));
 sg13g2_a21oi_1 _5297_ (.A1(net2097),
    .A2(net865),
    .Y(_0923_),
    .B1(_0870_));
 sg13g2_a22oi_1 _5298_ (.Y(_0924_),
    .B1(_0922_),
    .B2(_0923_),
    .A2(_0813_),
    .A1(net2141));
 sg13g2_inv_1 _5299_ (.Y(_0064_),
    .A(net866));
 sg13g2_mux2_2 _5300_ (.A0(_0848_),
    .A1(_0855_),
    .S(net2050),
    .X(_0925_));
 sg13g2_nor2b_1 _5301_ (.A(_0925_),
    .B_N(net2057),
    .Y(_0926_));
 sg13g2_o21ai_1 _5302_ (.B1(net1761),
    .Y(_0927_),
    .A1(_0111_),
    .A2(net2057));
 sg13g2_nor2_1 _5303_ (.A(net2035),
    .B(_0712_),
    .Y(_0928_));
 sg13g2_nand2_1 _5304_ (.Y(_0929_),
    .A(_0111_),
    .B(net1775));
 sg13g2_a21oi_1 _5305_ (.A1(net1758),
    .A2(_0928_),
    .Y(_0930_),
    .B1(_0929_));
 sg13g2_a21oi_1 _5306_ (.A1(_0112_),
    .A2(net1782),
    .Y(_0931_),
    .B1(_0930_));
 sg13g2_o21ai_1 _5307_ (.B1(_0931_),
    .Y(_0932_),
    .A1(_0926_),
    .A2(_0927_));
 sg13g2_nand2_1 _5308_ (.Y(_0933_),
    .A(net2162),
    .B(_0932_));
 sg13g2_nand2_1 _5309_ (.Y(_0934_),
    .A(net2095),
    .B(net929));
 sg13g2_nor2b_1 _5310_ (.A(net2140),
    .B_N(net2139),
    .Y(_0935_));
 sg13g2_nor2b_2 _5311_ (.A(net2137),
    .B_N(_0935_),
    .Y(_0936_));
 sg13g2_nand3_1 _5312_ (.B(_0809_),
    .C(_0936_),
    .A(\debug_controller_inst.grid_out_valid ),
    .Y(_0937_));
 sg13g2_and2_1 _5313_ (.A(net2309),
    .B(_0937_),
    .X(_0938_));
 sg13g2_nand3_1 _5314_ (.B(_0934_),
    .C(_0938_),
    .A(_0933_),
    .Y(_0939_));
 sg13g2_nand2_2 _5315_ (.Y(_0940_),
    .A(net2148),
    .B(_0519_));
 sg13g2_o21ai_1 _5316_ (.B1(net930),
    .Y(_0065_),
    .A1(_0937_),
    .A2(_0940_));
 sg13g2_nand2_2 _5317_ (.Y(_0941_),
    .A(net2145),
    .B(_0519_));
 sg13g2_mux2_2 _5318_ (.A0(_0877_),
    .A1(_0883_),
    .S(net2050),
    .X(_0942_));
 sg13g2_inv_1 _5319_ (.Y(_0943_),
    .A(_0942_));
 sg13g2_o21ai_1 _5320_ (.B1(net1761),
    .Y(_0944_),
    .A1(_0113_),
    .A2(net2057));
 sg13g2_a21oi_1 _5321_ (.A1(net2057),
    .A2(_0943_),
    .Y(_0945_),
    .B1(_0944_));
 sg13g2_a22oi_1 _5322_ (.Y(_0946_),
    .B1(net1775),
    .B2(net957),
    .A2(net1782),
    .A1(_0114_));
 sg13g2_nand3_1 _5323_ (.B(net2034),
    .C(_0928_),
    .A(net1758),
    .Y(_0947_));
 sg13g2_nand2_1 _5324_ (.Y(_0948_),
    .A(_0946_),
    .B(_0947_));
 sg13g2_o21ai_1 _5325_ (.B1(net2161),
    .Y(_0949_),
    .A1(_0945_),
    .A2(_0948_));
 sg13g2_nand2_1 _5326_ (.Y(_0950_),
    .A(net2095),
    .B(net957));
 sg13g2_nand3_1 _5327_ (.B(_0949_),
    .C(_0950_),
    .A(_0938_),
    .Y(_0951_));
 sg13g2_o21ai_1 _5328_ (.B1(net958),
    .Y(_0066_),
    .A1(_0937_),
    .A2(_0941_));
 sg13g2_nand2_2 _5329_ (.Y(_0952_),
    .A(net2143),
    .B(_0519_));
 sg13g2_mux2_2 _5330_ (.A0(_0896_),
    .A1(_0901_),
    .S(net2050),
    .X(_0953_));
 sg13g2_inv_1 _5331_ (.Y(_0954_),
    .A(_0953_));
 sg13g2_o21ai_1 _5332_ (.B1(net1761),
    .Y(_0955_),
    .A1(_0115_),
    .A2(net2057));
 sg13g2_a21oi_1 _5333_ (.A1(net2057),
    .A2(_0954_),
    .Y(_0956_),
    .B1(_0955_));
 sg13g2_a22oi_1 _5334_ (.Y(_0957_),
    .B1(net1775),
    .B2(net935),
    .A2(net1782),
    .A1(_0116_));
 sg13g2_nand2_1 _5335_ (.Y(_0958_),
    .A(_0947_),
    .B(_0957_));
 sg13g2_o21ai_1 _5336_ (.B1(net2161),
    .Y(_0959_),
    .A1(_0956_),
    .A2(_0958_));
 sg13g2_nand2_1 _5337_ (.Y(_0960_),
    .A(net2095),
    .B(net935));
 sg13g2_nand3_1 _5338_ (.B(_0959_),
    .C(_0960_),
    .A(_0938_),
    .Y(_0961_));
 sg13g2_o21ai_1 _5339_ (.B1(net936),
    .Y(_0004_),
    .A1(_0937_),
    .A2(_0952_));
 sg13g2_nand2_2 _5340_ (.Y(_0962_),
    .A(net2141),
    .B(_0519_));
 sg13g2_mux2_2 _5341_ (.A0(_0913_),
    .A1(_0916_),
    .S(net2050),
    .X(_0963_));
 sg13g2_inv_1 _5342_ (.Y(_0964_),
    .A(_0963_));
 sg13g2_o21ai_1 _5343_ (.B1(net1761),
    .Y(_0965_),
    .A1(_0117_),
    .A2(net2057));
 sg13g2_a21oi_1 _5344_ (.A1(net2057),
    .A2(_0964_),
    .Y(_0966_),
    .B1(_0965_));
 sg13g2_a22oi_1 _5345_ (.Y(_0967_),
    .B1(net1775),
    .B2(_0117_),
    .A2(net1782),
    .A1(_0118_));
 sg13g2_nand2_1 _5346_ (.Y(_0968_),
    .A(_0947_),
    .B(_0967_));
 sg13g2_o21ai_1 _5347_ (.B1(net2162),
    .Y(_0969_),
    .A1(_0966_),
    .A2(_0968_));
 sg13g2_nand2_1 _5348_ (.Y(_0970_),
    .A(net2095),
    .B(net897));
 sg13g2_nand3_1 _5349_ (.B(_0969_),
    .C(_0970_),
    .A(_0938_),
    .Y(_0971_));
 sg13g2_o21ai_1 _5350_ (.B1(net898),
    .Y(_0005_),
    .A1(_0937_),
    .A2(_0962_));
 sg13g2_nand2_1 _5351_ (.Y(_0972_),
    .A(net2139),
    .B(net2140));
 sg13g2_nor3_2 _5352_ (.A(net2137),
    .B(_0810_),
    .C(_0972_),
    .Y(_0973_));
 sg13g2_nor2_2 _5353_ (.A(net2053),
    .B(_0650_),
    .Y(_0974_));
 sg13g2_a21oi_2 _5354_ (.B1(net2054),
    .Y(_0975_),
    .A2(_0690_),
    .A1(_0689_));
 sg13g2_nor2_1 _5355_ (.A(_0974_),
    .B(_0975_),
    .Y(_0976_));
 sg13g2_o21ai_1 _5356_ (.B1(net1767),
    .Y(_0977_),
    .A1(_0119_),
    .A2(net2060));
 sg13g2_a21oi_1 _5357_ (.A1(net2060),
    .A2(_0976_),
    .Y(_0978_),
    .B1(_0977_));
 sg13g2_nor2_2 _5358_ (.A(_0701_),
    .B(_0705_),
    .Y(_0979_));
 sg13g2_nand2_1 _5359_ (.Y(_0980_),
    .A(_0119_),
    .B(net1780));
 sg13g2_a21oi_1 _5360_ (.A1(net1758),
    .A2(_0979_),
    .Y(_0981_),
    .B1(_0980_));
 sg13g2_a21o_1 _5361_ (.A2(net1788),
    .A1(_0120_),
    .B1(_0981_),
    .X(_0982_));
 sg13g2_o21ai_1 _5362_ (.B1(net2175),
    .Y(_0983_),
    .A1(_0978_),
    .A2(_0982_));
 sg13g2_nand2b_1 _5363_ (.Y(_0984_),
    .B(net2311),
    .A_N(_0973_));
 sg13g2_a21oi_1 _5364_ (.A1(net2101),
    .A2(net880),
    .Y(_0985_),
    .B1(_0984_));
 sg13g2_a22oi_1 _5365_ (.Y(_0986_),
    .B1(_0983_),
    .B2(_0985_),
    .A2(_0973_),
    .A1(net2148));
 sg13g2_inv_1 _5366_ (.Y(_0006_),
    .A(net881));
 sg13g2_nor2_1 _5367_ (.A(net2053),
    .B(_0763_),
    .Y(_0987_));
 sg13g2_a21oi_1 _5368_ (.A1(_0764_),
    .A2(_0770_),
    .Y(_0988_),
    .B1(net2056));
 sg13g2_nor2_2 _5369_ (.A(_0987_),
    .B(_0988_),
    .Y(_0989_));
 sg13g2_o21ai_1 _5370_ (.B1(net1767),
    .Y(_0990_),
    .A1(_0121_),
    .A2(net2060));
 sg13g2_a21oi_1 _5371_ (.A1(net2060),
    .A2(_0989_),
    .Y(_0991_),
    .B1(_0990_));
 sg13g2_nand3_1 _5372_ (.B(_0863_),
    .C(_0979_),
    .A(net1758),
    .Y(_0992_));
 sg13g2_a22oi_1 _5373_ (.Y(_0993_),
    .B1(net1780),
    .B2(net924),
    .A2(net1788),
    .A1(_0122_));
 sg13g2_nand2_1 _5374_ (.Y(_0994_),
    .A(_0992_),
    .B(_0993_));
 sg13g2_o21ai_1 _5375_ (.B1(net2175),
    .Y(_0995_),
    .A1(_0991_),
    .A2(_0994_));
 sg13g2_a21oi_1 _5376_ (.A1(net2101),
    .A2(net924),
    .Y(_0996_),
    .B1(_0984_));
 sg13g2_a22oi_1 _5377_ (.Y(_0997_),
    .B1(_0995_),
    .B2(_0996_),
    .A2(_0973_),
    .A1(net2146));
 sg13g2_inv_1 _5378_ (.Y(_0007_),
    .A(net925));
 sg13g2_mux2_2 _5379_ (.A0(_0782_),
    .A1(_0786_),
    .S(net2051),
    .X(_0998_));
 sg13g2_o21ai_1 _5380_ (.B1(net1767),
    .Y(_0999_),
    .A1(_0123_),
    .A2(net2060));
 sg13g2_a21oi_1 _5381_ (.A1(net2061),
    .A2(_0998_),
    .Y(_1000_),
    .B1(_0999_));
 sg13g2_a22oi_1 _5382_ (.Y(_1001_),
    .B1(net1780),
    .B2(net933),
    .A2(net1788),
    .A1(_0124_));
 sg13g2_nand2_1 _5383_ (.Y(_1002_),
    .A(_0992_),
    .B(_1001_));
 sg13g2_o21ai_1 _5384_ (.B1(net2175),
    .Y(_1003_),
    .A1(_1000_),
    .A2(_1002_));
 sg13g2_a21oi_1 _5385_ (.A1(net2101),
    .A2(net933),
    .Y(_1004_),
    .B1(_0984_));
 sg13g2_a22oi_1 _5386_ (.Y(_1005_),
    .B1(_1003_),
    .B2(_1004_),
    .A2(_0973_),
    .A1(net2144));
 sg13g2_inv_1 _5387_ (.Y(_0008_),
    .A(net934));
 sg13g2_a21oi_1 _5388_ (.A1(_0795_),
    .A2(_0799_),
    .Y(_1006_),
    .B1(net2055));
 sg13g2_a21oi_2 _5389_ (.B1(_1006_),
    .Y(_1007_),
    .A2(_0801_),
    .A1(net2055));
 sg13g2_nor2b_1 _5390_ (.A(_1007_),
    .B_N(net2061),
    .Y(_1008_));
 sg13g2_o21ai_1 _5391_ (.B1(net1766),
    .Y(_1009_),
    .A1(_0125_),
    .A2(net2061));
 sg13g2_a22oi_1 _5392_ (.Y(_1010_),
    .B1(net1778),
    .B2(_0125_),
    .A2(net1787),
    .A1(_0126_));
 sg13g2_and2_1 _5393_ (.A(_0992_),
    .B(_1010_),
    .X(_1011_));
 sg13g2_o21ai_1 _5394_ (.B1(_1011_),
    .Y(_1012_),
    .A1(_1008_),
    .A2(_1009_));
 sg13g2_nand2_1 _5395_ (.Y(_1013_),
    .A(net2168),
    .B(_1012_));
 sg13g2_a21oi_1 _5396_ (.A1(net2098),
    .A2(net885),
    .Y(_1014_),
    .B1(_0984_));
 sg13g2_a22oi_1 _5397_ (.Y(_1015_),
    .B1(_1013_),
    .B2(_1014_),
    .A2(_0973_),
    .A1(net2141));
 sg13g2_inv_1 _5398_ (.Y(_0009_),
    .A(net886));
 sg13g2_nand2_1 _5399_ (.Y(_1016_),
    .A(net2137),
    .B(_0517_));
 sg13g2_nor2_2 _5400_ (.A(_0810_),
    .B(_1016_),
    .Y(_1017_));
 sg13g2_nor2_2 _5401_ (.A(_0098_),
    .B(net2059),
    .Y(_1018_));
 sg13g2_or2_1 _5402_ (.X(_1019_),
    .B(net2060),
    .A(_0098_));
 sg13g2_nor4_1 _5403_ (.A(net2039),
    .B(_0692_),
    .C(_0693_),
    .D(net1951),
    .Y(_1020_));
 sg13g2_o21ai_1 _5404_ (.B1(net1764),
    .Y(_1021_),
    .A1(_0104_),
    .A2(net2048));
 sg13g2_nor2_2 _5405_ (.A(_0702_),
    .B(_0707_),
    .Y(_1022_));
 sg13g2_nand2_1 _5406_ (.Y(_1023_),
    .A(net1758),
    .B(_1022_));
 sg13g2_a21oi_1 _5407_ (.A1(net1808),
    .A2(net2032),
    .Y(_1024_),
    .B1(_4058_));
 sg13g2_a22oi_1 _5408_ (.Y(_1025_),
    .B1(_1023_),
    .B2(_1024_),
    .A2(net1785),
    .A1(_0103_));
 sg13g2_o21ai_1 _5409_ (.B1(_1025_),
    .Y(_1026_),
    .A1(_1020_),
    .A2(_1021_));
 sg13g2_nor2_2 _5410_ (.A(net2307),
    .B(_1017_),
    .Y(_1027_));
 sg13g2_o21ai_1 _5411_ (.B1(_1027_),
    .Y(_1028_),
    .A1(net2165),
    .A2(_4058_));
 sg13g2_a21oi_1 _5412_ (.A1(net2165),
    .A2(_1026_),
    .Y(_1029_),
    .B1(_1028_));
 sg13g2_a21o_1 _5413_ (.A2(_1017_),
    .A1(net2148),
    .B1(net1005),
    .X(_0010_));
 sg13g2_nand3_1 _5414_ (.B(_0774_),
    .C(net1953),
    .A(net2036),
    .Y(_1030_));
 sg13g2_o21ai_1 _5415_ (.B1(net1765),
    .Y(_1031_),
    .A1(_0106_),
    .A2(net2048));
 sg13g2_nand2b_1 _5416_ (.Y(_1032_),
    .B(_1030_),
    .A_N(_1031_));
 sg13g2_nand3_1 _5417_ (.B(net2034),
    .C(_1022_),
    .A(net1758),
    .Y(_1033_));
 sg13g2_a22oi_1 _5418_ (.Y(_1034_),
    .B1(net1777),
    .B2(_0106_),
    .A2(net1785),
    .A1(_0105_));
 sg13g2_nand3_1 _5419_ (.B(_1033_),
    .C(_1034_),
    .A(_1032_),
    .Y(_1035_));
 sg13g2_o21ai_1 _5420_ (.B1(_1027_),
    .Y(_1036_),
    .A1(net2164),
    .A2(_4059_));
 sg13g2_a21oi_1 _5421_ (.A1(net2164),
    .A2(_1035_),
    .Y(_1037_),
    .B1(_1036_));
 sg13g2_a21o_1 _5422_ (.A2(_1017_),
    .A1(net2147),
    .B1(net992),
    .X(_0011_));
 sg13g2_nand3_1 _5423_ (.B(_0787_),
    .C(net1953),
    .A(net2036),
    .Y(_1038_));
 sg13g2_o21ai_1 _5424_ (.B1(net1764),
    .Y(_1039_),
    .A1(_0108_),
    .A2(net2048));
 sg13g2_nand2b_1 _5425_ (.Y(_1040_),
    .B(_1038_),
    .A_N(_1039_));
 sg13g2_a22oi_1 _5426_ (.Y(_1041_),
    .B1(net1777),
    .B2(_0108_),
    .A2(net1785),
    .A1(_0107_));
 sg13g2_nand3_1 _5427_ (.B(_1040_),
    .C(_1041_),
    .A(_1033_),
    .Y(_1042_));
 sg13g2_o21ai_1 _5428_ (.B1(_1027_),
    .Y(_1043_),
    .A1(net2164),
    .A2(_4060_));
 sg13g2_a21oi_1 _5429_ (.A1(net2164),
    .A2(_1042_),
    .Y(_1044_),
    .B1(_1043_));
 sg13g2_a21o_1 _5430_ (.A2(_1017_),
    .A1(net2144),
    .B1(_1044_),
    .X(_0012_));
 sg13g2_nor2_1 _5431_ (.A(_0803_),
    .B(net1951),
    .Y(_1045_));
 sg13g2_o21ai_1 _5432_ (.B1(net1764),
    .Y(_1046_),
    .A1(_0110_),
    .A2(net2048));
 sg13g2_a21o_1 _5433_ (.A2(_1045_),
    .A1(net2036),
    .B1(_1046_),
    .X(_1047_));
 sg13g2_a22oi_1 _5434_ (.Y(_1048_),
    .B1(net1777),
    .B2(_0110_),
    .A2(net1785),
    .A1(net1006));
 sg13g2_nand3_1 _5435_ (.B(_1047_),
    .C(net1007),
    .A(_1033_),
    .Y(_1049_));
 sg13g2_o21ai_1 _5436_ (.B1(_1027_),
    .Y(_1050_),
    .A1(net2164),
    .A2(_4061_));
 sg13g2_a21oi_1 _5437_ (.A1(net2164),
    .A2(_1049_),
    .Y(_1051_),
    .B1(_1050_));
 sg13g2_a21o_1 _5438_ (.A2(_1017_),
    .A1(net2141),
    .B1(net1008),
    .X(_0013_));
 sg13g2_nand2_1 _5439_ (.Y(_1052_),
    .A(net2138),
    .B(_0811_));
 sg13g2_nor2_1 _5440_ (.A(_0810_),
    .B(_1052_),
    .Y(_1053_));
 sg13g2_nor2_1 _5441_ (.A(_0856_),
    .B(net1952),
    .Y(_1054_));
 sg13g2_o21ai_1 _5442_ (.B1(net2177),
    .Y(_1055_),
    .A1(_0127_),
    .A2(net2049));
 sg13g2_a21oi_1 _5443_ (.A1(net2037),
    .A2(_1054_),
    .Y(_1056_),
    .B1(_1055_));
 sg13g2_nor2_1 _5444_ (.A(_0702_),
    .B(_0710_),
    .Y(_1057_));
 sg13g2_and2_1 _5445_ (.A(_0751_),
    .B(_1057_),
    .X(_1058_));
 sg13g2_nor3_1 _5446_ (.A(net2177),
    .B(_4070_),
    .C(_1058_),
    .Y(_1059_));
 sg13g2_or3_1 _5447_ (.A(net1792),
    .B(_1056_),
    .C(_1059_),
    .X(_1060_));
 sg13g2_a21oi_1 _5448_ (.A1(_4070_),
    .A2(net1791),
    .Y(_1061_),
    .B1(net2100));
 sg13g2_o21ai_1 _5449_ (.B1(net2316),
    .Y(_1062_),
    .A1(_0810_),
    .A2(_1052_));
 sg13g2_a221oi_1 _5450_ (.B2(_1061_),
    .C1(_1062_),
    .B1(_1060_),
    .A1(net2100),
    .Y(_1063_),
    .A2(net913));
 sg13g2_a21o_1 _5451_ (.A2(_1053_),
    .A1(net2149),
    .B1(_1063_),
    .X(_0015_));
 sg13g2_nand2b_1 _5452_ (.Y(_1064_),
    .B(net1793),
    .A_N(_0128_));
 sg13g2_o21ai_1 _5453_ (.B1(_0761_),
    .Y(_1065_),
    .A1(_1058_),
    .A2(_1064_));
 sg13g2_nand3_1 _5454_ (.B(_0884_),
    .C(net1953),
    .A(net2037),
    .Y(_1066_));
 sg13g2_o21ai_1 _5455_ (.B1(_1066_),
    .Y(_1067_),
    .A1(_0128_),
    .A2(net2049));
 sg13g2_o21ai_1 _5456_ (.B1(_1065_),
    .Y(_1068_),
    .A1(_3986_),
    .A2(_1067_));
 sg13g2_o21ai_1 _5457_ (.B1(net2171),
    .Y(_1069_),
    .A1(net976),
    .A2(net1793));
 sg13g2_inv_1 _5458_ (.Y(_1070_),
    .A(_1069_));
 sg13g2_a221oi_1 _5459_ (.B2(_1070_),
    .C1(_1062_),
    .B1(_1068_),
    .A1(net2100),
    .Y(_1071_),
    .A2(net976));
 sg13g2_a21o_1 _5460_ (.A2(_1053_),
    .A1(net2146),
    .B1(_1071_),
    .X(_0016_));
 sg13g2_or3_1 _5461_ (.A(_0129_),
    .B(net1792),
    .C(_1058_),
    .X(_1072_));
 sg13g2_nor2_1 _5462_ (.A(_0902_),
    .B(net1952),
    .Y(_1073_));
 sg13g2_nor2_1 _5463_ (.A(_0129_),
    .B(net2049),
    .Y(_1074_));
 sg13g2_a21oi_1 _5464_ (.A1(net2037),
    .A2(_1073_),
    .Y(_1075_),
    .B1(_1074_));
 sg13g2_a22oi_1 _5465_ (.Y(_1076_),
    .B1(_1075_),
    .B2(net2177),
    .A2(_1072_),
    .A1(net1759));
 sg13g2_o21ai_1 _5466_ (.B1(net2173),
    .Y(_1077_),
    .A1(net903),
    .A2(net1793));
 sg13g2_a21oi_1 _5467_ (.A1(net2100),
    .A2(net903),
    .Y(_1078_),
    .B1(_1062_));
 sg13g2_o21ai_1 _5468_ (.B1(_1078_),
    .Y(_1079_),
    .A1(_1076_),
    .A2(_1077_));
 sg13g2_nand3_1 _5469_ (.B(net2144),
    .C(_0811_),
    .A(net2138),
    .Y(_1080_));
 sg13g2_o21ai_1 _5470_ (.B1(_1079_),
    .Y(_0017_),
    .A1(_0810_),
    .A2(_1080_));
 sg13g2_nor3_1 _5471_ (.A(_0130_),
    .B(net1792),
    .C(_1058_),
    .Y(_1081_));
 sg13g2_nand2_2 _5472_ (.Y(_1082_),
    .A(_0917_),
    .B(net1953));
 sg13g2_o21ai_1 _5473_ (.B1(net2177),
    .Y(_1083_),
    .A1(_0130_),
    .A2(net2049));
 sg13g2_inv_1 _5474_ (.Y(_1084_),
    .A(_1083_));
 sg13g2_o21ai_1 _5475_ (.B1(_1084_),
    .Y(_1085_),
    .A1(net2042),
    .A2(_1082_));
 sg13g2_o21ai_1 _5476_ (.B1(_1085_),
    .Y(_1086_),
    .A1(net1768),
    .A2(_1081_));
 sg13g2_o21ai_1 _5477_ (.B1(net2173),
    .Y(_1087_),
    .A1(_0130_),
    .A2(net1793));
 sg13g2_inv_1 _5478_ (.Y(_1088_),
    .A(_1087_));
 sg13g2_a221oi_1 _5479_ (.B2(_1088_),
    .C1(_1062_),
    .B1(_1086_),
    .A1(net2100),
    .Y(_1089_),
    .A2(net973));
 sg13g2_a21o_1 _5480_ (.A2(_1053_),
    .A1(net2142),
    .B1(net974),
    .X(_0018_));
 sg13g2_nand4_1 _5481_ (.B(\debug_controller_inst.grid_out_valid ),
    .C(_0809_),
    .A(net2137),
    .Y(_1090_),
    .D(_0935_));
 sg13g2_nor2_1 _5482_ (.A(_0925_),
    .B(net1951),
    .Y(_1091_));
 sg13g2_o21ai_1 _5483_ (.B1(net1764),
    .Y(_1092_),
    .A1(_0131_),
    .A2(net2048));
 sg13g2_a21oi_1 _5484_ (.A1(net2036),
    .A2(_1091_),
    .Y(_1093_),
    .B1(_1092_));
 sg13g2_nor2_2 _5485_ (.A(_0702_),
    .B(_0712_),
    .Y(_1094_));
 sg13g2_nand2_1 _5486_ (.Y(_1095_),
    .A(_0131_),
    .B(net1777));
 sg13g2_a21oi_1 _5487_ (.A1(_0861_),
    .A2(_1094_),
    .Y(_1096_),
    .B1(_1095_));
 sg13g2_a21o_1 _5488_ (.A2(net1784),
    .A1(net810),
    .B1(_1096_),
    .X(_1097_));
 sg13g2_o21ai_1 _5489_ (.B1(net2166),
    .Y(_1098_),
    .A1(_1093_),
    .A2(_1097_));
 sg13g2_nand2_1 _5490_ (.Y(_1099_),
    .A(net2097),
    .B(net887));
 sg13g2_and2_1 _5491_ (.A(net2311),
    .B(_1090_),
    .X(_1100_));
 sg13g2_nand3_1 _5492_ (.B(_1099_),
    .C(_1100_),
    .A(_1098_),
    .Y(_1101_));
 sg13g2_o21ai_1 _5493_ (.B1(net888),
    .Y(_0019_),
    .A1(_0940_),
    .A2(_1090_));
 sg13g2_nor2_1 _5494_ (.A(_0942_),
    .B(net1951),
    .Y(_1102_));
 sg13g2_o21ai_1 _5495_ (.B1(net1762),
    .Y(_1103_),
    .A1(_0133_),
    .A2(net2048));
 sg13g2_a21oi_1 _5496_ (.A1(net2036),
    .A2(_1102_),
    .Y(_1104_),
    .B1(_1103_));
 sg13g2_nand3_1 _5497_ (.B(net2034),
    .C(_1094_),
    .A(_0861_),
    .Y(_1105_));
 sg13g2_a22oi_1 _5498_ (.Y(_1106_),
    .B1(net1776),
    .B2(_0133_),
    .A2(net1784),
    .A1(_0134_));
 sg13g2_nand2_1 _5499_ (.Y(_1107_),
    .A(_1105_),
    .B(_1106_));
 sg13g2_o21ai_1 _5500_ (.B1(net2162),
    .Y(_1108_),
    .A1(_1104_),
    .A2(_1107_));
 sg13g2_nand2_1 _5501_ (.Y(_1109_),
    .A(net2096),
    .B(net945));
 sg13g2_nand3_1 _5502_ (.B(_1108_),
    .C(_1109_),
    .A(_1100_),
    .Y(_1110_));
 sg13g2_o21ai_1 _5503_ (.B1(net946),
    .Y(_0020_),
    .A1(_0941_),
    .A2(_1090_));
 sg13g2_nor2_1 _5504_ (.A(_0953_),
    .B(net1951),
    .Y(_1111_));
 sg13g2_o21ai_1 _5505_ (.B1(net1762),
    .Y(_1112_),
    .A1(_0135_),
    .A2(net2048));
 sg13g2_a21oi_1 _5506_ (.A1(net2036),
    .A2(_1111_),
    .Y(_1113_),
    .B1(_1112_));
 sg13g2_a22oi_1 _5507_ (.Y(_1114_),
    .B1(net1776),
    .B2(net931),
    .A2(net1784),
    .A1(net927));
 sg13g2_nand2_1 _5508_ (.Y(_1115_),
    .A(_1105_),
    .B(_1114_));
 sg13g2_o21ai_1 _5509_ (.B1(net2163),
    .Y(_1116_),
    .A1(_1113_),
    .A2(_1115_));
 sg13g2_nand2_1 _5510_ (.Y(_1117_),
    .A(net2095),
    .B(net931));
 sg13g2_nand3_1 _5511_ (.B(_1116_),
    .C(_1117_),
    .A(_1100_),
    .Y(_1118_));
 sg13g2_o21ai_1 _5512_ (.B1(net932),
    .Y(_0021_),
    .A1(_0952_),
    .A2(_1090_));
 sg13g2_nor2_1 _5513_ (.A(_0963_),
    .B(net1951),
    .Y(_1119_));
 sg13g2_o21ai_1 _5514_ (.B1(net1762),
    .Y(_1120_),
    .A1(_0137_),
    .A2(net2048));
 sg13g2_a21oi_1 _5515_ (.A1(net2036),
    .A2(_1119_),
    .Y(_1121_),
    .B1(_1120_));
 sg13g2_a22oi_1 _5516_ (.Y(_1122_),
    .B1(net1776),
    .B2(_0137_),
    .A2(net1784),
    .A1(net883));
 sg13g2_nand2_1 _5517_ (.Y(_1123_),
    .A(_1105_),
    .B(_1122_));
 sg13g2_o21ai_1 _5518_ (.B1(net2162),
    .Y(_1124_),
    .A1(_1121_),
    .A2(_1123_));
 sg13g2_nand2_1 _5519_ (.Y(_1125_),
    .A(net2095),
    .B(net963));
 sg13g2_nand3_1 _5520_ (.B(_1124_),
    .C(_1125_),
    .A(_1100_),
    .Y(_1126_));
 sg13g2_o21ai_1 _5521_ (.B1(_1126_),
    .Y(_0022_),
    .A1(_0962_),
    .A2(_1090_));
 sg13g2_nand3_1 _5522_ (.B(net2139),
    .C(net2140),
    .A(net2138),
    .Y(_1127_));
 sg13g2_nor2_2 _5523_ (.A(_0810_),
    .B(_1127_),
    .Y(_1128_));
 sg13g2_nor4_1 _5524_ (.A(net2043),
    .B(_0974_),
    .C(_0975_),
    .D(net1952),
    .Y(_1129_));
 sg13g2_o21ai_1 _5525_ (.B1(net1767),
    .Y(_1130_),
    .A1(_0139_),
    .A2(net2049));
 sg13g2_nand4_1 _5526_ (.B(_0703_),
    .C(_0704_),
    .A(net2035),
    .Y(_1131_),
    .D(net1758));
 sg13g2_a21oi_1 _5527_ (.A1(_0508_),
    .A2(net2033),
    .Y(_1132_),
    .B1(_4071_));
 sg13g2_a22oi_1 _5528_ (.Y(_1133_),
    .B1(_1131_),
    .B2(_1132_),
    .A2(net1788),
    .A1(_0140_));
 sg13g2_o21ai_1 _5529_ (.B1(_1133_),
    .Y(_1134_),
    .A1(_1129_),
    .A2(_1130_));
 sg13g2_nor2_2 _5530_ (.A(net2302),
    .B(_1128_),
    .Y(_1135_));
 sg13g2_o21ai_1 _5531_ (.B1(_1135_),
    .Y(_1136_),
    .A1(net2174),
    .A2(_4071_));
 sg13g2_a21oi_1 _5532_ (.A1(net2174),
    .A2(_1134_),
    .Y(_1137_),
    .B1(_1136_));
 sg13g2_a21o_1 _5533_ (.A2(_1128_),
    .A1(net2149),
    .B1(net1023),
    .X(_0023_));
 sg13g2_nand3_1 _5534_ (.B(_0989_),
    .C(_1018_),
    .A(net2037),
    .Y(_1138_));
 sg13g2_o21ai_1 _5535_ (.B1(net1768),
    .Y(_1139_),
    .A1(_0141_),
    .A2(net2049));
 sg13g2_nand2b_1 _5536_ (.Y(_1140_),
    .B(_1138_),
    .A_N(_1139_));
 sg13g2_or2_1 _5537_ (.X(_1141_),
    .B(_1131_),
    .A(net2033));
 sg13g2_a22oi_1 _5538_ (.Y(_1142_),
    .B1(net1780),
    .B2(_0141_),
    .A2(net1789),
    .A1(_0142_));
 sg13g2_nand3_1 _5539_ (.B(_1141_),
    .C(_1142_),
    .A(_1140_),
    .Y(_1143_));
 sg13g2_o21ai_1 _5540_ (.B1(_1135_),
    .Y(_1144_),
    .A1(net2174),
    .A2(_4072_));
 sg13g2_a21oi_1 _5541_ (.A1(net2173),
    .A2(_1143_),
    .Y(_1145_),
    .B1(_1144_));
 sg13g2_a21o_1 _5542_ (.A2(_1128_),
    .A1(net2146),
    .B1(net1019),
    .X(_0024_));
 sg13g2_and2_1 _5543_ (.A(_0998_),
    .B(net1953),
    .X(_1146_));
 sg13g2_o21ai_1 _5544_ (.B1(net1767),
    .Y(_1147_),
    .A1(_0143_),
    .A2(net2049));
 sg13g2_a21oi_1 _5545_ (.A1(net2037),
    .A2(_1146_),
    .Y(_1148_),
    .B1(_1147_));
 sg13g2_a22oi_1 _5546_ (.Y(_1149_),
    .B1(net1781),
    .B2(_0143_),
    .A2(net1789),
    .A1(_0144_));
 sg13g2_nand2_1 _5547_ (.Y(_1150_),
    .A(_1141_),
    .B(_1149_));
 sg13g2_o21ai_1 _5548_ (.B1(net2174),
    .Y(_1151_),
    .A1(_1148_),
    .A2(_1150_));
 sg13g2_nand2_1 _5549_ (.Y(_1152_),
    .A(net2101),
    .B(net959));
 sg13g2_nand3_1 _5550_ (.B(_1151_),
    .C(_1152_),
    .A(_1135_),
    .Y(_1153_));
 sg13g2_nand4_1 _5551_ (.B(net2139),
    .C(net2140),
    .A(net2138),
    .Y(_1154_),
    .D(net2143));
 sg13g2_o21ai_1 _5552_ (.B1(net960),
    .Y(_0026_),
    .A1(_0810_),
    .A2(_1154_));
 sg13g2_nor2_1 _5553_ (.A(_1007_),
    .B(net1952),
    .Y(_1155_));
 sg13g2_o21ai_1 _5554_ (.B1(net1768),
    .Y(_1156_),
    .A1(_0145_),
    .A2(net2049));
 sg13g2_a21o_1 _5555_ (.A2(_1155_),
    .A1(net2038),
    .B1(_1156_),
    .X(_1157_));
 sg13g2_a22oi_1 _5556_ (.Y(_1158_),
    .B1(net1780),
    .B2(_0145_),
    .A2(net1789),
    .A1(_0146_));
 sg13g2_nand3_1 _5557_ (.B(_1157_),
    .C(_1158_),
    .A(_1141_),
    .Y(_1159_));
 sg13g2_o21ai_1 _5558_ (.B1(_1135_),
    .Y(_1160_),
    .A1(net2173),
    .A2(_4073_));
 sg13g2_a21oi_1 _5559_ (.A1(net2173),
    .A2(_1159_),
    .Y(_1161_),
    .B1(_1160_));
 sg13g2_a21o_1 _5560_ (.A2(_1128_),
    .A1(net2142),
    .B1(net1000),
    .X(_0027_));
 sg13g2_o21ai_1 _5561_ (.B1(net1763),
    .Y(_1162_),
    .A1(net952),
    .A2(net2044));
 sg13g2_a21oi_1 _5562_ (.A1(net2044),
    .A2(_0694_),
    .Y(_1163_),
    .B1(_1162_));
 sg13g2_or3_2 _5563_ (.A(_0700_),
    .B(_0746_),
    .C(_0747_),
    .X(_1164_));
 sg13g2_nor2_1 _5564_ (.A(net1809),
    .B(_1164_),
    .Y(_1165_));
 sg13g2_nand2_1 _5565_ (.Y(_1166_),
    .A(_0752_),
    .B(net1773));
 sg13g2_a21oi_1 _5566_ (.A1(net1808),
    .A2(net2032),
    .Y(_1167_),
    .B1(_4062_));
 sg13g2_a221oi_1 _5567_ (.B2(_1167_),
    .C1(_1163_),
    .B1(_1166_),
    .A1(net929),
    .Y(_1168_),
    .A2(net1783));
 sg13g2_nor2_1 _5568_ (.A(net2095),
    .B(_1168_),
    .Y(_1169_));
 sg13g2_and3_2 _5569_ (.X(_1170_),
    .A(\debug_controller_inst.grid_out_addr[3] ),
    .B(\debug_controller_inst.grid_out_valid ),
    .C(_0518_));
 sg13g2_nor2_2 _5570_ (.A(net2301),
    .B(_1170_),
    .Y(_1171_));
 sg13g2_o21ai_1 _5571_ (.B1(_1171_),
    .Y(_1172_),
    .A1(net2162),
    .A2(_4062_));
 sg13g2_nand2_1 _5572_ (.Y(_1173_),
    .A(net2148),
    .B(_1170_));
 sg13g2_o21ai_1 _5573_ (.B1(_1173_),
    .Y(_0028_),
    .A1(_1169_),
    .A2(_1172_));
 sg13g2_o21ai_1 _5574_ (.B1(net1761),
    .Y(_1174_),
    .A1(_0114_),
    .A2(net2045));
 sg13g2_a21o_1 _5575_ (.A2(_0774_),
    .A1(net2045),
    .B1(_1174_),
    .X(_1175_));
 sg13g2_nand3_1 _5576_ (.B(net2034),
    .C(net1773),
    .A(_0752_),
    .Y(_1176_));
 sg13g2_a22oi_1 _5577_ (.Y(_1177_),
    .B1(net1775),
    .B2(net1016),
    .A2(net1782),
    .A1(_0113_));
 sg13g2_nand3_1 _5578_ (.B(_1176_),
    .C(_1177_),
    .A(_1175_),
    .Y(_1178_));
 sg13g2_o21ai_1 _5579_ (.B1(_1171_),
    .Y(_1179_),
    .A1(net2161),
    .A2(_4063_));
 sg13g2_a21oi_1 _5580_ (.A1(net2161),
    .A2(_1178_),
    .Y(_1180_),
    .B1(_1179_));
 sg13g2_a21o_1 _5581_ (.A2(_1170_),
    .A1(net2145),
    .B1(net1017),
    .X(_0029_));
 sg13g2_o21ai_1 _5582_ (.B1(net1761),
    .Y(_1181_),
    .A1(_0116_),
    .A2(net2045));
 sg13g2_a21o_1 _5583_ (.A2(_0787_),
    .A1(net2045),
    .B1(_1181_),
    .X(_1182_));
 sg13g2_a22oi_1 _5584_ (.Y(_1183_),
    .B1(net1775),
    .B2(_0116_),
    .A2(net1782),
    .A1(_0115_));
 sg13g2_nand3_1 _5585_ (.B(_1182_),
    .C(_1183_),
    .A(_1176_),
    .Y(_1184_));
 sg13g2_o21ai_1 _5586_ (.B1(_1171_),
    .Y(_1185_),
    .A1(net2161),
    .A2(_4064_));
 sg13g2_a21oi_1 _5587_ (.A1(net2161),
    .A2(_1184_),
    .Y(_1186_),
    .B1(_1185_));
 sg13g2_a21o_1 _5588_ (.A2(_1170_),
    .A1(net2143),
    .B1(net1015),
    .X(_0030_));
 sg13g2_o21ai_1 _5589_ (.B1(net1761),
    .Y(_1187_),
    .A1(_0118_),
    .A2(net2045));
 sg13g2_inv_1 _5590_ (.Y(_1188_),
    .A(_1187_));
 sg13g2_o21ai_1 _5591_ (.B1(_1188_),
    .Y(_1189_),
    .A1(_0526_),
    .A2(_0803_));
 sg13g2_a22oi_1 _5592_ (.Y(_1190_),
    .B1(net1775),
    .B2(_0118_),
    .A2(net1782),
    .A1(_0117_));
 sg13g2_nand3_1 _5593_ (.B(_1189_),
    .C(_1190_),
    .A(_1176_),
    .Y(_1191_));
 sg13g2_o21ai_1 _5594_ (.B1(_1171_),
    .Y(_1192_),
    .A1(net2161),
    .A2(_4065_));
 sg13g2_a21oi_1 _5595_ (.A1(net2163),
    .A2(_1191_),
    .Y(_1193_),
    .B1(_1192_));
 sg13g2_a21o_1 _5596_ (.A2(_1170_),
    .A1(net2141),
    .B1(_1193_),
    .X(_0031_));
 sg13g2_nor2_1 _5597_ (.A(_0526_),
    .B(_0856_),
    .Y(_1194_));
 sg13g2_o21ai_1 _5598_ (.B1(net1764),
    .Y(_1195_),
    .A1(_0132_),
    .A2(net2046));
 sg13g2_nand2_1 _5599_ (.Y(_1196_),
    .A(_0132_),
    .B(net1777));
 sg13g2_a21oi_1 _5600_ (.A1(_0860_),
    .A2(net1774),
    .Y(_1197_),
    .B1(_1196_));
 sg13g2_a21oi_1 _5601_ (.A1(_0131_),
    .A2(net1784),
    .Y(_1198_),
    .B1(_1197_));
 sg13g2_o21ai_1 _5602_ (.B1(_1198_),
    .Y(_1199_),
    .A1(_1194_),
    .A2(_1195_));
 sg13g2_nand2_1 _5603_ (.Y(_1200_),
    .A(net2097),
    .B(net810));
 sg13g2_nor2_2 _5604_ (.A(_4057_),
    .B(_0809_),
    .Y(_1201_));
 sg13g2_nand2b_2 _5605_ (.Y(_1202_),
    .B(\debug_controller_inst.grid_out_valid ),
    .A_N(_0809_));
 sg13g2_nor3_2 _5606_ (.A(net2138),
    .B(_0812_),
    .C(_1202_),
    .Y(_1203_));
 sg13g2_nand2b_1 _5607_ (.Y(_1204_),
    .B(net2311),
    .A_N(_1203_));
 sg13g2_a21oi_1 _5608_ (.A1(net2166),
    .A2(_1199_),
    .Y(_1205_),
    .B1(_1204_));
 sg13g2_a22oi_1 _5609_ (.Y(_1206_),
    .B1(_1205_),
    .B2(_1200_),
    .A2(_1203_),
    .A1(net2148));
 sg13g2_inv_1 _5610_ (.Y(_0032_),
    .A(_1206_));
 sg13g2_o21ai_1 _5611_ (.B1(net1764),
    .Y(_1207_),
    .A1(_0134_),
    .A2(net2046));
 sg13g2_a21oi_1 _5612_ (.A1(net2046),
    .A2(_0884_),
    .Y(_1208_),
    .B1(_1207_));
 sg13g2_nand3_1 _5613_ (.B(net2034),
    .C(net1773),
    .A(_0860_),
    .Y(_1209_));
 sg13g2_a22oi_1 _5614_ (.Y(_1210_),
    .B1(net1775),
    .B2(net922),
    .A2(net1784),
    .A1(_0133_));
 sg13g2_nand2_1 _5615_ (.Y(_1211_),
    .A(_1209_),
    .B(_1210_));
 sg13g2_o21ai_1 _5616_ (.B1(net2166),
    .Y(_1212_),
    .A1(_1208_),
    .A2(_1211_));
 sg13g2_a21oi_1 _5617_ (.A1(net2097),
    .A2(net922),
    .Y(_1213_),
    .B1(_1204_));
 sg13g2_a22oi_1 _5618_ (.Y(_1214_),
    .B1(_1212_),
    .B2(_1213_),
    .A2(_1203_),
    .A1(net2145));
 sg13g2_inv_1 _5619_ (.Y(_0033_),
    .A(net923));
 sg13g2_o21ai_1 _5620_ (.B1(net1764),
    .Y(_1215_),
    .A1(_0136_),
    .A2(net2046));
 sg13g2_a21oi_1 _5621_ (.A1(net2046),
    .A2(_0903_),
    .Y(_1216_),
    .B1(_1215_));
 sg13g2_a22oi_1 _5622_ (.Y(_1217_),
    .B1(net1777),
    .B2(_0136_),
    .A2(net1784),
    .A1(_0135_));
 sg13g2_nand2_1 _5623_ (.Y(_1218_),
    .A(_1209_),
    .B(_1217_));
 sg13g2_o21ai_1 _5624_ (.B1(net2166),
    .Y(_1219_),
    .A1(_1216_),
    .A2(_1218_));
 sg13g2_a21oi_1 _5625_ (.A1(net2097),
    .A2(net927),
    .Y(_1220_),
    .B1(_1204_));
 sg13g2_a22oi_1 _5626_ (.Y(_1221_),
    .B1(_1219_),
    .B2(_1220_),
    .A2(_1203_),
    .A1(net2143));
 sg13g2_inv_1 _5627_ (.Y(_0034_),
    .A(net928));
 sg13g2_o21ai_1 _5628_ (.B1(net1764),
    .Y(_1222_),
    .A1(_0138_),
    .A2(net2046));
 sg13g2_a21oi_1 _5629_ (.A1(net2046),
    .A2(_0917_),
    .Y(_1223_),
    .B1(_1222_));
 sg13g2_a22oi_1 _5630_ (.Y(_1224_),
    .B1(net1777),
    .B2(net883),
    .A2(net1784),
    .A1(_0137_));
 sg13g2_nand2_1 _5631_ (.Y(_1225_),
    .A(_1209_),
    .B(_1224_));
 sg13g2_o21ai_1 _5632_ (.B1(net2166),
    .Y(_1226_),
    .A1(_1223_),
    .A2(_1225_));
 sg13g2_a21oi_1 _5633_ (.A1(net2097),
    .A2(net883),
    .Y(_1227_),
    .B1(_1204_));
 sg13g2_a22oi_1 _5634_ (.Y(_1228_),
    .B1(_1226_),
    .B2(_1227_),
    .A2(_1203_),
    .A1(net2141));
 sg13g2_inv_1 _5635_ (.Y(_0035_),
    .A(net884));
 sg13g2_nand2_2 _5636_ (.Y(_1229_),
    .A(_0936_),
    .B(_1201_));
 sg13g2_mux2_1 _5637_ (.A0(_0147_),
    .A1(_0925_),
    .S(net2044),
    .X(_1230_));
 sg13g2_nor3_2 _5638_ (.A(net2035),
    .B(_0712_),
    .C(_1164_),
    .Y(_1231_));
 sg13g2_nand2_1 _5639_ (.Y(_1232_),
    .A(_3986_),
    .B(_0147_));
 sg13g2_o21ai_1 _5640_ (.B1(net1795),
    .Y(_1233_),
    .A1(_1231_),
    .A2(_1232_));
 sg13g2_a21oi_1 _5641_ (.A1(net2178),
    .A2(_1230_),
    .Y(_1234_),
    .B1(_1233_));
 sg13g2_o21ai_1 _5642_ (.B1(net2163),
    .Y(_1235_),
    .A1(net895),
    .A2(net1795));
 sg13g2_a21oi_2 _5643_ (.B1(net2301),
    .Y(_1236_),
    .A2(_1201_),
    .A1(_0936_));
 sg13g2_o21ai_1 _5644_ (.B1(_1236_),
    .Y(_1237_),
    .A1(_1234_),
    .A2(_1235_));
 sg13g2_a21o_1 _5645_ (.A2(net895),
    .A1(net2096),
    .B1(_1237_),
    .X(_1238_));
 sg13g2_o21ai_1 _5646_ (.B1(_1238_),
    .Y(_0037_),
    .A1(_0940_),
    .A2(_1229_));
 sg13g2_or3_1 _5647_ (.A(_0148_),
    .B(net1792),
    .C(_1231_),
    .X(_1239_));
 sg13g2_nor2_1 _5648_ (.A(_0148_),
    .B(net2045),
    .Y(_1240_));
 sg13g2_a21oi_1 _5649_ (.A1(net2044),
    .A2(_0943_),
    .Y(_1241_),
    .B1(_1240_));
 sg13g2_a22oi_1 _5650_ (.Y(_1242_),
    .B1(_1241_),
    .B2(net2178),
    .A2(_1239_),
    .A1(net1760));
 sg13g2_o21ai_1 _5651_ (.B1(net2163),
    .Y(_1243_),
    .A1(net875),
    .A2(net1795));
 sg13g2_o21ai_1 _5652_ (.B1(_1236_),
    .Y(_1244_),
    .A1(_1242_),
    .A2(_1243_));
 sg13g2_a21o_1 _5653_ (.A2(net875),
    .A1(net2103),
    .B1(_1244_),
    .X(_1245_));
 sg13g2_o21ai_1 _5654_ (.B1(_1245_),
    .Y(_0038_),
    .A1(_0941_),
    .A2(_1229_));
 sg13g2_or3_1 _5655_ (.A(_0149_),
    .B(net1792),
    .C(_1231_),
    .X(_1246_));
 sg13g2_nor2_1 _5656_ (.A(_0149_),
    .B(net2044),
    .Y(_1247_));
 sg13g2_a21oi_1 _5657_ (.A1(net2044),
    .A2(_0954_),
    .Y(_1248_),
    .B1(_1247_));
 sg13g2_a22oi_1 _5658_ (.Y(_1249_),
    .B1(_1248_),
    .B2(net2178),
    .A2(_1246_),
    .A1(net1760));
 sg13g2_o21ai_1 _5659_ (.B1(net2163),
    .Y(_1250_),
    .A1(net872),
    .A2(net1795));
 sg13g2_o21ai_1 _5660_ (.B1(_1236_),
    .Y(_1251_),
    .A1(_1249_),
    .A2(_1250_));
 sg13g2_a21o_1 _5661_ (.A2(net872),
    .A1(net2096),
    .B1(_1251_),
    .X(_1252_));
 sg13g2_o21ai_1 _5662_ (.B1(_1252_),
    .Y(_0039_),
    .A1(_0952_),
    .A2(_1229_));
 sg13g2_or3_1 _5663_ (.A(_0150_),
    .B(net1792),
    .C(_1231_),
    .X(_1253_));
 sg13g2_nor2_1 _5664_ (.A(_0150_),
    .B(net2044),
    .Y(_1254_));
 sg13g2_a21oi_1 _5665_ (.A1(net2044),
    .A2(_0964_),
    .Y(_1255_),
    .B1(_1254_));
 sg13g2_a22oi_1 _5666_ (.Y(_1256_),
    .B1(_1255_),
    .B2(net2178),
    .A2(_1253_),
    .A1(net1760));
 sg13g2_o21ai_1 _5667_ (.B1(net2163),
    .Y(_1257_),
    .A1(net908),
    .A2(net1795));
 sg13g2_o21ai_1 _5668_ (.B1(_1236_),
    .Y(_1258_),
    .A1(_1256_),
    .A2(_1257_));
 sg13g2_a21o_1 _5669_ (.A2(net908),
    .A1(net2096),
    .B1(_1258_),
    .X(_1259_));
 sg13g2_o21ai_1 _5670_ (.B1(_1259_),
    .Y(_0040_),
    .A1(_0962_),
    .A2(_1229_));
 sg13g2_nor3_2 _5671_ (.A(net2137),
    .B(_0972_),
    .C(_1202_),
    .Y(_1260_));
 sg13g2_o21ai_1 _5672_ (.B1(net1766),
    .Y(_1261_),
    .A1(net861),
    .A2(net2047));
 sg13g2_a21oi_1 _5673_ (.A1(net2047),
    .A2(_0976_),
    .Y(_1262_),
    .B1(_1261_));
 sg13g2_nand2_1 _5674_ (.Y(_1263_),
    .A(_0152_),
    .B(net1786));
 sg13g2_nand2_2 _5675_ (.Y(_1264_),
    .A(_0979_),
    .B(net1773));
 sg13g2_nand3_1 _5676_ (.B(net1779),
    .C(_1264_),
    .A(net861),
    .Y(_1265_));
 sg13g2_nand2_1 _5677_ (.Y(_1266_),
    .A(_1263_),
    .B(_1265_));
 sg13g2_o21ai_1 _5678_ (.B1(net2167),
    .Y(_1267_),
    .A1(_1262_),
    .A2(_1266_));
 sg13g2_nand2b_2 _5679_ (.Y(_1268_),
    .B(net2311),
    .A_N(_1260_));
 sg13g2_a21oi_1 _5680_ (.A1(net2098),
    .A2(net861),
    .Y(_1269_),
    .B1(_1268_));
 sg13g2_a22oi_1 _5681_ (.Y(_1270_),
    .B1(_1267_),
    .B2(_1269_),
    .A2(_1260_),
    .A1(net2148));
 sg13g2_inv_1 _5682_ (.Y(_0041_),
    .A(net862));
 sg13g2_o21ai_1 _5683_ (.B1(net1763),
    .Y(_1271_),
    .A1(_0153_),
    .A2(net2047));
 sg13g2_a21oi_1 _5684_ (.A1(net2047),
    .A2(_0989_),
    .Y(_1272_),
    .B1(_1271_));
 sg13g2_nor2_1 _5685_ (.A(net2032),
    .B(_1264_),
    .Y(_1273_));
 sg13g2_a22oi_1 _5686_ (.Y(_1274_),
    .B1(net1779),
    .B2(net914),
    .A2(net1783),
    .A1(_0154_));
 sg13g2_o21ai_1 _5687_ (.B1(_1274_),
    .Y(_1275_),
    .A1(net2032),
    .A2(_1264_));
 sg13g2_o21ai_1 _5688_ (.B1(net2169),
    .Y(_1276_),
    .A1(_1272_),
    .A2(_1275_));
 sg13g2_a21oi_1 _5689_ (.A1(net2096),
    .A2(net914),
    .Y(_1277_),
    .B1(_1268_));
 sg13g2_a22oi_1 _5690_ (.Y(_1278_),
    .B1(_1276_),
    .B2(_1277_),
    .A2(_1260_),
    .A1(net2145));
 sg13g2_inv_1 _5691_ (.Y(_0042_),
    .A(net915));
 sg13g2_o21ai_1 _5692_ (.B1(net1769),
    .Y(_1279_),
    .A1(net867),
    .A2(net2046));
 sg13g2_a21oi_1 _5693_ (.A1(net2047),
    .A2(_0998_),
    .Y(_1280_),
    .B1(_1279_));
 sg13g2_a22oi_1 _5694_ (.Y(_1281_),
    .B1(net1776),
    .B2(net867),
    .A2(net1786),
    .A1(net1026));
 sg13g2_o21ai_1 _5695_ (.B1(_1281_),
    .Y(_1282_),
    .A1(net2032),
    .A2(_1264_));
 sg13g2_o21ai_1 _5696_ (.B1(net2167),
    .Y(_1283_),
    .A1(_1280_),
    .A2(_1282_));
 sg13g2_a21oi_1 _5697_ (.A1(net2098),
    .A2(net867),
    .Y(_1284_),
    .B1(_1268_));
 sg13g2_a22oi_1 _5698_ (.Y(_1285_),
    .B1(_1283_),
    .B2(_1284_),
    .A2(_1260_),
    .A1(net2143));
 sg13g2_inv_1 _5699_ (.Y(_0043_),
    .A(_1285_));
 sg13g2_nor2_1 _5700_ (.A(_0526_),
    .B(_1007_),
    .Y(_1286_));
 sg13g2_o21ai_1 _5701_ (.B1(net1763),
    .Y(_1287_),
    .A1(_0157_),
    .A2(net2045));
 sg13g2_a221oi_1 _5702_ (.B2(net868),
    .C1(_1273_),
    .B1(net1776),
    .A1(_0158_),
    .Y(_1288_),
    .A2(net1783));
 sg13g2_o21ai_1 _5703_ (.B1(_1288_),
    .Y(_1289_),
    .A1(_1286_),
    .A2(_1287_));
 sg13g2_nand2_1 _5704_ (.Y(_1290_),
    .A(net2096),
    .B(net868));
 sg13g2_a21oi_1 _5705_ (.A1(net2163),
    .A2(_1289_),
    .Y(_1291_),
    .B1(_1268_));
 sg13g2_a22oi_1 _5706_ (.Y(_1292_),
    .B1(_1290_),
    .B2(_1291_),
    .A2(_1260_),
    .A1(net2141));
 sg13g2_inv_1 _5707_ (.Y(_0044_),
    .A(net869));
 sg13g2_nor2_2 _5708_ (.A(_1016_),
    .B(_1202_),
    .Y(_1293_));
 sg13g2_nand3_1 _5709_ (.B(_0694_),
    .C(_1018_),
    .A(net2040),
    .Y(_1294_));
 sg13g2_o21ai_1 _5710_ (.B1(_1294_),
    .Y(_1295_),
    .A1(_0120_),
    .A2(net2040));
 sg13g2_nand2_1 _5711_ (.Y(_1296_),
    .A(_1022_),
    .B(net1773));
 sg13g2_a21oi_1 _5712_ (.A1(net1808),
    .A2(net2033),
    .Y(_1297_),
    .B1(_4066_));
 sg13g2_a22oi_1 _5713_ (.Y(_1298_),
    .B1(_1296_),
    .B2(_1297_),
    .A2(net1788),
    .A1(_0119_));
 sg13g2_o21ai_1 _5714_ (.B1(_1298_),
    .Y(_1299_),
    .A1(net1760),
    .A2(_1295_));
 sg13g2_nor2_2 _5715_ (.A(net2301),
    .B(_1293_),
    .Y(_1300_));
 sg13g2_o21ai_1 _5716_ (.B1(_1300_),
    .Y(_1301_),
    .A1(net2167),
    .A2(_4066_));
 sg13g2_a21oi_1 _5717_ (.A1(net2167),
    .A2(_1299_),
    .Y(_1302_),
    .B1(_1301_));
 sg13g2_a21o_1 _5718_ (.A2(_1293_),
    .A1(net2148),
    .B1(_1302_),
    .X(_0045_));
 sg13g2_nand3_1 _5719_ (.B(_0774_),
    .C(net1953),
    .A(net2039),
    .Y(_1303_));
 sg13g2_nand2_1 _5720_ (.Y(_1304_),
    .A(_4067_),
    .B(net2036));
 sg13g2_nand3_1 _5721_ (.B(_1303_),
    .C(_1304_),
    .A(net1766),
    .Y(_1305_));
 sg13g2_nand3_1 _5722_ (.B(_1022_),
    .C(net1773),
    .A(net2034),
    .Y(_1306_));
 sg13g2_a22oi_1 _5723_ (.Y(_1307_),
    .B1(net1778),
    .B2(net1012),
    .A2(net1786),
    .A1(_0121_));
 sg13g2_nand3_1 _5724_ (.B(_1306_),
    .C(_1307_),
    .A(_1305_),
    .Y(_1308_));
 sg13g2_o21ai_1 _5725_ (.B1(_1300_),
    .Y(_1309_),
    .A1(net2168),
    .A2(_4067_));
 sg13g2_a21oi_1 _5726_ (.A1(net2167),
    .A2(_1308_),
    .Y(_1310_),
    .B1(_1309_));
 sg13g2_a21o_1 _5727_ (.A2(_1293_),
    .A1(net2145),
    .B1(net1013),
    .X(_0046_));
 sg13g2_nand3_1 _5728_ (.B(_0787_),
    .C(net1953),
    .A(net2039),
    .Y(_1311_));
 sg13g2_nand2_1 _5729_ (.Y(_1312_),
    .A(_4068_),
    .B(net2038));
 sg13g2_nand3_1 _5730_ (.B(_1311_),
    .C(_1312_),
    .A(net1766),
    .Y(_1313_));
 sg13g2_a22oi_1 _5731_ (.Y(_1314_),
    .B1(net1778),
    .B2(net1024),
    .A2(net1786),
    .A1(_0123_));
 sg13g2_nand3_1 _5732_ (.B(_1313_),
    .C(_1314_),
    .A(_1306_),
    .Y(_1315_));
 sg13g2_o21ai_1 _5733_ (.B1(_1300_),
    .Y(_1316_),
    .A1(net2168),
    .A2(_4068_));
 sg13g2_a21oi_1 _5734_ (.A1(net2168),
    .A2(_1315_),
    .Y(_1317_),
    .B1(_1316_));
 sg13g2_a21o_1 _5735_ (.A2(_1293_),
    .A1(net2143),
    .B1(_1317_),
    .X(_0048_));
 sg13g2_nor3_1 _5736_ (.A(net2038),
    .B(_0803_),
    .C(net1951),
    .Y(_1318_));
 sg13g2_o21ai_1 _5737_ (.B1(net1766),
    .Y(_1319_),
    .A1(_0126_),
    .A2(net2039));
 sg13g2_a22oi_1 _5738_ (.Y(_1320_),
    .B1(net1778),
    .B2(_0126_),
    .A2(net1787),
    .A1(_0125_));
 sg13g2_and2_1 _5739_ (.A(_1306_),
    .B(_1320_),
    .X(_1321_));
 sg13g2_o21ai_1 _5740_ (.B1(_1321_),
    .Y(_1322_),
    .A1(_1318_),
    .A2(_1319_));
 sg13g2_o21ai_1 _5741_ (.B1(_1300_),
    .Y(_1323_),
    .A1(net2167),
    .A2(_4069_));
 sg13g2_a21oi_1 _5742_ (.A1(net2167),
    .A2(_1322_),
    .Y(_1324_),
    .B1(_1323_));
 sg13g2_a21o_1 _5743_ (.A2(_1293_),
    .A1(net2141),
    .B1(_1324_),
    .X(_0049_));
 sg13g2_nand2b_2 _5744_ (.Y(_1325_),
    .B(_1201_),
    .A_N(_1052_));
 sg13g2_o21ai_1 _5745_ (.B1(net1767),
    .Y(_1326_),
    .A1(_0140_),
    .A2(net2042));
 sg13g2_a21oi_1 _5746_ (.A1(net2042),
    .A2(_1054_),
    .Y(_1327_),
    .B1(_1326_));
 sg13g2_nand2_1 _5747_ (.Y(_1328_),
    .A(_0140_),
    .B(net1781));
 sg13g2_a21oi_1 _5748_ (.A1(_1057_),
    .A2(net1774),
    .Y(_1329_),
    .B1(_1328_));
 sg13g2_a21o_1 _5749_ (.A2(net1789),
    .A1(_0139_),
    .B1(_1329_),
    .X(_1330_));
 sg13g2_o21ai_1 _5750_ (.B1(net2173),
    .Y(_1331_),
    .A1(_1327_),
    .A2(_1330_));
 sg13g2_nand2_1 _5751_ (.Y(_1332_),
    .A(net2100),
    .B(net926));
 sg13g2_and2_1 _5752_ (.A(net2316),
    .B(_1325_),
    .X(_1333_));
 sg13g2_nand3_1 _5753_ (.B(_1332_),
    .C(_1333_),
    .A(_1331_),
    .Y(_1334_));
 sg13g2_o21ai_1 _5754_ (.B1(_1334_),
    .Y(_0050_),
    .A1(_3984_),
    .A2(_1325_));
 sg13g2_nand3_1 _5755_ (.B(_0884_),
    .C(net1953),
    .A(net2043),
    .Y(_1335_));
 sg13g2_o21ai_1 _5756_ (.B1(_1335_),
    .Y(_1336_),
    .A1(_0142_),
    .A2(net2042));
 sg13g2_nor2_1 _5757_ (.A(net1759),
    .B(_1336_),
    .Y(_1337_));
 sg13g2_nand3_1 _5758_ (.B(_1057_),
    .C(net1774),
    .A(net2034),
    .Y(_1338_));
 sg13g2_a22oi_1 _5759_ (.Y(_1339_),
    .B1(net1780),
    .B2(_0142_),
    .A2(net1788),
    .A1(_0141_));
 sg13g2_nand2_1 _5760_ (.Y(_1340_),
    .A(_1338_),
    .B(_1339_));
 sg13g2_o21ai_1 _5761_ (.B1(net2174),
    .Y(_1341_),
    .A1(_1337_),
    .A2(_1340_));
 sg13g2_nand2_1 _5762_ (.Y(_1342_),
    .A(net2101),
    .B(net940));
 sg13g2_nand3_1 _5763_ (.B(_1341_),
    .C(_1342_),
    .A(_1333_),
    .Y(_1343_));
 sg13g2_o21ai_1 _5764_ (.B1(net941),
    .Y(_0051_),
    .A1(_3982_),
    .A2(_1325_));
 sg13g2_o21ai_1 _5765_ (.B1(net1767),
    .Y(_1344_),
    .A1(_0144_),
    .A2(net2042));
 sg13g2_a21oi_1 _5766_ (.A1(net2042),
    .A2(_1073_),
    .Y(_1345_),
    .B1(_1344_));
 sg13g2_a22oi_1 _5767_ (.Y(_1346_),
    .B1(net1780),
    .B2(_0144_),
    .A2(net1788),
    .A1(_0143_));
 sg13g2_nand2_1 _5768_ (.Y(_1347_),
    .A(_1338_),
    .B(_1346_));
 sg13g2_o21ai_1 _5769_ (.B1(net2173),
    .Y(_1348_),
    .A1(_1345_),
    .A2(_1347_));
 sg13g2_nand2_1 _5770_ (.Y(_1349_),
    .A(net2100),
    .B(net980));
 sg13g2_nand3_1 _5771_ (.B(_1348_),
    .C(_1349_),
    .A(_1333_),
    .Y(_1350_));
 sg13g2_o21ai_1 _5772_ (.B1(_1350_),
    .Y(_0052_),
    .A1(_1080_),
    .A2(_1202_));
 sg13g2_nor2_1 _5773_ (.A(net2037),
    .B(_1082_),
    .Y(_1351_));
 sg13g2_o21ai_1 _5774_ (.B1(net1767),
    .Y(_1352_),
    .A1(_0146_),
    .A2(net2042));
 sg13g2_nor2_1 _5775_ (.A(_1351_),
    .B(_1352_),
    .Y(_1353_));
 sg13g2_a22oi_1 _5776_ (.Y(_1354_),
    .B1(net1780),
    .B2(_0146_),
    .A2(net1788),
    .A1(_0145_));
 sg13g2_nand2_1 _5777_ (.Y(_1355_),
    .A(_1338_),
    .B(_1354_));
 sg13g2_o21ai_1 _5778_ (.B1(net2173),
    .Y(_1356_),
    .A1(_1353_),
    .A2(_1355_));
 sg13g2_nand2_1 _5779_ (.Y(_1357_),
    .A(net2100),
    .B(net949));
 sg13g2_nand3_1 _5780_ (.B(_1356_),
    .C(_1357_),
    .A(_1333_),
    .Y(_1358_));
 sg13g2_o21ai_1 _5781_ (.B1(net950),
    .Y(_0053_),
    .A1(_3979_),
    .A2(_1325_));
 sg13g2_nand3_1 _5782_ (.B(_0935_),
    .C(_1201_),
    .A(net2137),
    .Y(_1359_));
 sg13g2_o21ai_1 _5783_ (.B1(net1766),
    .Y(_1360_),
    .A1(_0152_),
    .A2(net2039));
 sg13g2_a21oi_1 _5784_ (.A1(net2039),
    .A2(_1091_),
    .Y(_1361_),
    .B1(_1360_));
 sg13g2_nand2_1 _5785_ (.Y(_1362_),
    .A(_0152_),
    .B(net1779));
 sg13g2_a21oi_1 _5786_ (.A1(_1094_),
    .A2(net1773),
    .Y(_1363_),
    .B1(_1362_));
 sg13g2_a21o_1 _5787_ (.A2(net1786),
    .A1(net861),
    .B1(_1363_),
    .X(_1364_));
 sg13g2_o21ai_1 _5788_ (.B1(net2167),
    .Y(_1365_),
    .A1(_1361_),
    .A2(_1364_));
 sg13g2_nand2_1 _5789_ (.Y(_1366_),
    .A(net2098),
    .B(net876));
 sg13g2_and2_1 _5790_ (.A(net2311),
    .B(_1359_),
    .X(_1367_));
 sg13g2_nand3_1 _5791_ (.B(_1366_),
    .C(_1367_),
    .A(_1365_),
    .Y(_1368_));
 sg13g2_o21ai_1 _5792_ (.B1(net877),
    .Y(_0054_),
    .A1(_0940_),
    .A2(_1359_));
 sg13g2_o21ai_1 _5793_ (.B1(net1761),
    .Y(_1369_),
    .A1(_0154_),
    .A2(net2040));
 sg13g2_a21oi_1 _5794_ (.A1(net2040),
    .A2(_1102_),
    .Y(_1370_),
    .B1(_1369_));
 sg13g2_nand3_1 _5795_ (.B(_1094_),
    .C(net1773),
    .A(net2034),
    .Y(_1371_));
 sg13g2_a22oi_1 _5796_ (.Y(_1372_),
    .B1(net1779),
    .B2(net911),
    .A2(net1783),
    .A1(_0153_));
 sg13g2_nand2_1 _5797_ (.Y(_1373_),
    .A(_1371_),
    .B(_1372_));
 sg13g2_o21ai_1 _5798_ (.B1(net2162),
    .Y(_1374_),
    .A1(_1370_),
    .A2(_1373_));
 sg13g2_nand2_1 _5799_ (.Y(_1375_),
    .A(net2095),
    .B(net911));
 sg13g2_nand3_1 _5800_ (.B(_1374_),
    .C(_1375_),
    .A(_1367_),
    .Y(_1376_));
 sg13g2_o21ai_1 _5801_ (.B1(net912),
    .Y(_0055_),
    .A1(_0941_),
    .A2(_1359_));
 sg13g2_o21ai_1 _5802_ (.B1(net1762),
    .Y(_1377_),
    .A1(_0156_),
    .A2(net2039));
 sg13g2_a21oi_1 _5803_ (.A1(net2039),
    .A2(_1111_),
    .Y(_1378_),
    .B1(_1377_));
 sg13g2_a22oi_1 _5804_ (.Y(_1379_),
    .B1(net1776),
    .B2(net891),
    .A2(net1786),
    .A1(net867));
 sg13g2_nand2_1 _5805_ (.Y(_1380_),
    .A(_1371_),
    .B(_1379_));
 sg13g2_o21ai_1 _5806_ (.B1(net2162),
    .Y(_1381_),
    .A1(_1378_),
    .A2(_1380_));
 sg13g2_nand2_1 _5807_ (.Y(_1382_),
    .A(net2097),
    .B(net891));
 sg13g2_nand3_1 _5808_ (.B(_1381_),
    .C(_1382_),
    .A(_1367_),
    .Y(_1383_));
 sg13g2_o21ai_1 _5809_ (.B1(net892),
    .Y(_0056_),
    .A1(_0952_),
    .A2(_1359_));
 sg13g2_o21ai_1 _5810_ (.B1(net1762),
    .Y(_1384_),
    .A1(_0158_),
    .A2(net2040));
 sg13g2_a21oi_1 _5811_ (.A1(net2040),
    .A2(_1119_),
    .Y(_1385_),
    .B1(_1384_));
 sg13g2_a22oi_1 _5812_ (.Y(_1386_),
    .B1(net1776),
    .B2(net917),
    .A2(net1782),
    .A1(_0157_));
 sg13g2_nand2_1 _5813_ (.Y(_1387_),
    .A(_1371_),
    .B(_1386_));
 sg13g2_o21ai_1 _5814_ (.B1(net2169),
    .Y(_1388_),
    .A1(_1385_),
    .A2(_1387_));
 sg13g2_nand2_1 _5815_ (.Y(_1389_),
    .A(net2096),
    .B(net917));
 sg13g2_nand3_1 _5816_ (.B(_1388_),
    .C(_1389_),
    .A(_1367_),
    .Y(_1390_));
 sg13g2_o21ai_1 _5817_ (.B1(net918),
    .Y(_0057_),
    .A1(_0962_),
    .A2(_1359_));
 sg13g2_nor2_1 _5818_ (.A(_1127_),
    .B(_1202_),
    .Y(_1391_));
 sg13g2_nor4_2 _5819_ (.A(net2037),
    .B(_0974_),
    .C(_0975_),
    .Y(_1392_),
    .D(net1951));
 sg13g2_o21ai_1 _5820_ (.B1(net2177),
    .Y(_1393_),
    .A1(_0159_),
    .A2(net2041));
 sg13g2_nor3_2 _5821_ (.A(_0702_),
    .B(_0705_),
    .C(_1164_),
    .Y(_1394_));
 sg13g2_nor3_1 _5822_ (.A(net2177),
    .B(_4074_),
    .C(_1394_),
    .Y(_1395_));
 sg13g2_nor2_1 _5823_ (.A(net1791),
    .B(_1395_),
    .Y(_1396_));
 sg13g2_o21ai_1 _5824_ (.B1(_1396_),
    .Y(_1397_),
    .A1(_1392_),
    .A2(_1393_));
 sg13g2_a21oi_1 _5825_ (.A1(_4074_),
    .A2(net1791),
    .Y(_1398_),
    .B1(net2099));
 sg13g2_o21ai_1 _5826_ (.B1(net2316),
    .Y(_1399_),
    .A1(_1127_),
    .A2(_1202_));
 sg13g2_a221oi_1 _5827_ (.B2(_1398_),
    .C1(_1399_),
    .B1(_1397_),
    .A1(net2099),
    .Y(_1400_),
    .A2(net889));
 sg13g2_a21o_1 _5828_ (.A2(_1391_),
    .A1(net2149),
    .B1(_1400_),
    .X(_0059_));
 sg13g2_nand2b_1 _5829_ (.Y(_1401_),
    .B(net1794),
    .A_N(_0160_));
 sg13g2_o21ai_1 _5830_ (.B1(net1759),
    .Y(_1402_),
    .A1(_1394_),
    .A2(_1401_));
 sg13g2_nand3_1 _5831_ (.B(_0989_),
    .C(_1018_),
    .A(net2041),
    .Y(_1403_));
 sg13g2_o21ai_1 _5832_ (.B1(_1403_),
    .Y(_1404_),
    .A1(_0160_),
    .A2(net2041));
 sg13g2_o21ai_1 _5833_ (.B1(_1402_),
    .Y(_1405_),
    .A1(_3986_),
    .A2(_1404_));
 sg13g2_o21ai_1 _5834_ (.B1(net2171),
    .Y(_1406_),
    .A1(net938),
    .A2(net1793));
 sg13g2_inv_1 _5835_ (.Y(_1407_),
    .A(_1406_));
 sg13g2_a221oi_1 _5836_ (.B2(_1407_),
    .C1(_1399_),
    .B1(_1405_),
    .A1(net2099),
    .Y(_1408_),
    .A2(net938));
 sg13g2_a21o_1 _5837_ (.A2(_1391_),
    .A1(net2145),
    .B1(_1408_),
    .X(_0060_));
 sg13g2_or3_1 _5838_ (.A(_0161_),
    .B(net1791),
    .C(_1394_),
    .X(_1409_));
 sg13g2_nand2_1 _5839_ (.Y(_1410_),
    .A(net2042),
    .B(_1146_));
 sg13g2_o21ai_1 _5840_ (.B1(net2177),
    .Y(_1411_),
    .A1(_0161_),
    .A2(net2041));
 sg13g2_inv_1 _5841_ (.Y(_1412_),
    .A(_1411_));
 sg13g2_a22oi_1 _5842_ (.Y(_1413_),
    .B1(_1410_),
    .B2(_1412_),
    .A2(_1409_),
    .A1(net1759));
 sg13g2_o21ai_1 _5843_ (.B1(net2171),
    .Y(_1414_),
    .A1(net871),
    .A2(net1793));
 sg13g2_a21oi_1 _5844_ (.A1(net2099),
    .A2(net871),
    .Y(_1415_),
    .B1(_1399_));
 sg13g2_o21ai_1 _5845_ (.B1(_1415_),
    .Y(_1416_),
    .A1(_1413_),
    .A2(_1414_));
 sg13g2_o21ai_1 _5846_ (.B1(_1416_),
    .Y(_0061_),
    .A1(_1154_),
    .A2(_1202_));
 sg13g2_nand2b_1 _5847_ (.Y(_1417_),
    .B(net1793),
    .A_N(_0162_));
 sg13g2_o21ai_1 _5848_ (.B1(net1759),
    .Y(_1418_),
    .A1(_1394_),
    .A2(_1417_));
 sg13g2_nor3_1 _5849_ (.A(net2037),
    .B(_1007_),
    .C(net1952),
    .Y(_1419_));
 sg13g2_o21ai_1 _5850_ (.B1(net2176),
    .Y(_1420_),
    .A1(_0162_),
    .A2(net2041));
 sg13g2_o21ai_1 _5851_ (.B1(_1418_),
    .Y(_1421_),
    .A1(_1419_),
    .A2(_1420_));
 sg13g2_o21ai_1 _5852_ (.B1(net2171),
    .Y(_1422_),
    .A1(_0162_),
    .A2(net1793));
 sg13g2_inv_1 _5853_ (.Y(_1423_),
    .A(_1422_));
 sg13g2_a221oi_1 _5854_ (.B2(_1423_),
    .C1(_1399_),
    .B1(_1421_),
    .A1(net2099),
    .Y(_1424_),
    .A2(net969));
 sg13g2_a21o_1 _5855_ (.A2(_1391_),
    .A1(net2142),
    .B1(net970),
    .X(_0062_));
 sg13g2_and2_1 _5856_ (.A(\draw_game_inst.y[7] ),
    .B(\draw_game_inst.board_y[6] ),
    .X(_1425_));
 sg13g2_nand2_1 _5857_ (.Y(_1426_),
    .A(net858),
    .B(net2031));
 sg13g2_nand2_1 _5858_ (.Y(_1427_),
    .A(net2189),
    .B(net2222));
 sg13g2_nor2_2 _5859_ (.A(net2085),
    .B(net2205),
    .Y(_1428_));
 sg13g2_nand2_1 _5860_ (.Y(_1429_),
    .A(net2196),
    .B(net2082));
 sg13g2_nand2_2 _5861_ (.Y(_1430_),
    .A(net2228),
    .B(net1947));
 sg13g2_inv_1 _5862_ (.Y(_1431_),
    .A(_1430_));
 sg13g2_nor2_1 _5863_ (.A(net2091),
    .B(net2184),
    .Y(_1432_));
 sg13g2_nand2_2 _5864_ (.Y(_1433_),
    .A(net2179),
    .B(_4042_));
 sg13g2_or4_1 _5865_ (.A(net994),
    .B(_1426_),
    .C(_1430_),
    .D(net1934),
    .X(_0068_));
 sg13g2_nor2_2 _5866_ (.A(net2286),
    .B(net2291),
    .Y(_1434_));
 sg13g2_or2_2 _5867_ (.X(_1435_),
    .B(net2292),
    .A(net2287));
 sg13g2_nor2_2 _5868_ (.A(net2063),
    .B(net2062),
    .Y(_1436_));
 sg13g2_nand2_2 _5869_ (.Y(_1437_),
    .A(net2286),
    .B(net2291));
 sg13g2_and2_1 _5870_ (.A(net2276),
    .B(net2280),
    .X(_1438_));
 sg13g2_a22oi_1 _5871_ (.Y(_1439_),
    .B1(_1436_),
    .B2(net2027),
    .A2(net2029),
    .A1(_4049_));
 sg13g2_nand4_1 _5872_ (.B(net2278),
    .C(net920),
    .A(_4039_),
    .Y(_0067_),
    .D(_1439_));
 sg13g2_and2_1 _5873_ (.A(net2322),
    .B(net543),
    .X(_0175_));
 sg13g2_and2_2 _5874_ (.A(\draw_game_inst.board_x[0] ),
    .B(\draw_game_inst.board_x[1] ),
    .X(_1440_));
 sg13g2_nand3_1 _5875_ (.B(\draw_game_inst.board_x[2] ),
    .C(_1440_),
    .A(net2296),
    .Y(_1441_));
 sg13g2_nor2b_1 _5876_ (.A(net2286),
    .B_N(net2291),
    .Y(_1442_));
 sg13g2_nand2b_2 _5877_ (.Y(_1443_),
    .B(net2293),
    .A_N(net2288));
 sg13g2_nor2_1 _5878_ (.A(net2276),
    .B(net2280),
    .Y(_1444_));
 sg13g2_nand4_1 _5879_ (.B(\draw_game_inst.x[9] ),
    .C(net2022),
    .A(\draw_game_inst.x[8] ),
    .Y(_1445_),
    .D(net2020));
 sg13g2_nor2_1 _5880_ (.A(_1441_),
    .B(_1445_),
    .Y(_1446_));
 sg13g2_nor2_1 _5881_ (.A(net2306),
    .B(_1446_),
    .Y(_1447_));
 sg13g2_o21ai_1 _5882_ (.B1(net2335),
    .Y(_1448_),
    .A1(_1441_),
    .A2(_1445_));
 sg13g2_and2_1 _5883_ (.A(net439),
    .B(net1815),
    .X(_0176_));
 sg13g2_nor2_1 _5884_ (.A(\draw_game_inst.board_x[0] ),
    .B(net987),
    .Y(_1449_));
 sg13g2_nor2b_1 _5885_ (.A(\draw_game_inst.board_x[0] ),
    .B_N(\draw_game_inst.board_x[1] ),
    .Y(_1450_));
 sg13g2_nor3_1 _5886_ (.A(net2306),
    .B(_1440_),
    .C(_1449_),
    .Y(_0177_));
 sg13g2_o21ai_1 _5887_ (.B1(net2335),
    .Y(_1451_),
    .A1(net939),
    .A2(_1440_));
 sg13g2_a21oi_1 _5888_ (.A1(net939),
    .A2(_1440_),
    .Y(_0178_),
    .B1(_1451_));
 sg13g2_a21oi_1 _5889_ (.A1(net939),
    .A2(_1440_),
    .Y(_1452_),
    .B1(net2296));
 sg13g2_nand2_1 _5890_ (.Y(_1453_),
    .A(net2336),
    .B(_1441_));
 sg13g2_nor2_2 _5891_ (.A(_1452_),
    .B(_1453_),
    .Y(_0179_));
 sg13g2_xnor2_1 _5892_ (.Y(_1454_),
    .A(net2062),
    .B(_1441_));
 sg13g2_nor2_1 _5893_ (.A(_1448_),
    .B(_1454_),
    .Y(_0180_));
 sg13g2_nor2_1 _5894_ (.A(_0096_),
    .B(_1441_),
    .Y(_1455_));
 sg13g2_xnor2_1 _5895_ (.Y(_1456_),
    .A(net2286),
    .B(_1455_));
 sg13g2_nor2_1 _5896_ (.A(_1448_),
    .B(_1456_),
    .Y(_0181_));
 sg13g2_nor2_2 _5897_ (.A(net2066),
    .B(net2064),
    .Y(_1457_));
 sg13g2_nand2_2 _5898_ (.Y(_1458_),
    .A(net2299),
    .B(net2289));
 sg13g2_and2_1 _5899_ (.A(net2296),
    .B(net2291),
    .X(_1459_));
 sg13g2_nand2_2 _5900_ (.Y(_1460_),
    .A(net2298),
    .B(net2292));
 sg13g2_nand2_2 _5901_ (.Y(_1461_),
    .A(net2287),
    .B(net2018));
 sg13g2_nor2_2 _5902_ (.A(_1437_),
    .B(_1441_),
    .Y(_1462_));
 sg13g2_xnor2_1 _5903_ (.Y(_1463_),
    .A(net2282),
    .B(_1462_));
 sg13g2_nor2_1 _5904_ (.A(_1448_),
    .B(_1463_),
    .Y(_0182_));
 sg13g2_a21oi_1 _5905_ (.A1(net2282),
    .A2(_1462_),
    .Y(_1464_),
    .B1(net2278));
 sg13g2_and2_1 _5906_ (.A(net2027),
    .B(_1462_),
    .X(_1465_));
 sg13g2_nor3_1 _5907_ (.A(_1448_),
    .B(_1464_),
    .C(_1465_),
    .Y(_0183_));
 sg13g2_nand2_1 _5908_ (.Y(_1466_),
    .A(net972),
    .B(_1465_));
 sg13g2_o21ai_1 _5909_ (.B1(net1815),
    .Y(_1467_),
    .A1(net972),
    .A2(_1465_));
 sg13g2_nor2b_1 _5910_ (.A(_1467_),
    .B_N(_1466_),
    .Y(_0184_));
 sg13g2_xor2_1 _5911_ (.B(_1466_),
    .A(net920),
    .X(_1468_));
 sg13g2_nor2_1 _5912_ (.A(_1448_),
    .B(_1468_),
    .Y(_0185_));
 sg13g2_nand3_1 _5913_ (.B(net2181),
    .C(net2031),
    .A(net874),
    .Y(_1469_));
 sg13g2_or2_1 _5914_ (.X(_1470_),
    .B(net2278),
    .A(\draw_game_inst.x[8] ));
 sg13g2_nand2_1 _5915_ (.Y(_1471_),
    .A(net984),
    .B(_1470_));
 sg13g2_nor2_1 _5916_ (.A(net2306),
    .B(net994),
    .Y(_1472_));
 sg13g2_nand3_1 _5917_ (.B(_1471_),
    .C(_1472_),
    .A(_1469_),
    .Y(_1473_));
 sg13g2_nor2_1 _5918_ (.A(net2195),
    .B(net2210),
    .Y(_1474_));
 sg13g2_nand2_2 _5919_ (.Y(_1475_),
    .A(net2089),
    .B(net2082));
 sg13g2_nor2_1 _5920_ (.A(net2268),
    .B(net2246),
    .Y(_1476_));
 sg13g2_nand2_1 _5921_ (.Y(_1477_),
    .A(net2105),
    .B(net2069));
 sg13g2_nor3_1 _5922_ (.A(net2179),
    .B(net2184),
    .C(net1925),
    .Y(_1478_));
 sg13g2_nand2_1 _5923_ (.Y(_1479_),
    .A(net2014),
    .B(_1478_));
 sg13g2_nand2b_2 _5924_ (.Y(_1480_),
    .B(\draw_game_inst.y[7] ),
    .A_N(\draw_game_inst.board_y[6] ));
 sg13g2_o21ai_1 _5925_ (.B1(_0088_),
    .Y(_1481_),
    .A1(_1479_),
    .A2(_1480_));
 sg13g2_nor2_1 _5926_ (.A(\draw_game_inst.y[9] ),
    .B(\draw_game_inst.y[8] ),
    .Y(_1482_));
 sg13g2_xnor2_1 _5927_ (.Y(_1483_),
    .A(\draw_game_inst.x[8] ),
    .B(net2027));
 sg13g2_mux2_1 _5928_ (.A0(_1482_),
    .A1(\draw_game_inst.y[8] ),
    .S(_1481_),
    .X(_1484_));
 sg13g2_or4_2 _5929_ (.A(\draw_game_inst.x[9] ),
    .B(\draw_game_inst.y[9] ),
    .C(_1483_),
    .D(_1484_),
    .X(_1485_));
 sg13g2_nor2_2 _5930_ (.A(\draw_game_inst.y[7] ),
    .B(\draw_game_inst.board_y[6] ),
    .Y(_1486_));
 sg13g2_a22oi_1 _5931_ (.Y(_1487_),
    .B1(net2281),
    .B2(\draw_game_inst.grid[43] ),
    .A2(net2277),
    .A1(\draw_game_inst.grid[47] ));
 sg13g2_a22oi_1 _5932_ (.Y(_1488_),
    .B1(net2019),
    .B2(\draw_game_inst.grid[39] ),
    .A2(net2025),
    .A1(\draw_game_inst.grid[35] ));
 sg13g2_o21ai_1 _5933_ (.B1(_1488_),
    .Y(_1489_),
    .A1(net2025),
    .A2(_1487_));
 sg13g2_nor2b_2 _5934_ (.A(\draw_game_inst.y[7] ),
    .B_N(\draw_game_inst.board_y[6] ),
    .Y(_1490_));
 sg13g2_a22oi_1 _5935_ (.Y(_1491_),
    .B1(net2281),
    .B2(\draw_game_inst.grid[59] ),
    .A2(net2277),
    .A1(\draw_game_inst.grid[63] ));
 sg13g2_a22oi_1 _5936_ (.Y(_1492_),
    .B1(net2019),
    .B2(\draw_game_inst.grid[55] ),
    .A2(net2025),
    .A1(\draw_game_inst.grid[51] ));
 sg13g2_o21ai_1 _5937_ (.B1(_1492_),
    .Y(_1493_),
    .A1(net2025),
    .A2(_1491_));
 sg13g2_a22oi_1 _5938_ (.Y(_1494_),
    .B1(net2282),
    .B2(\draw_game_inst.grid[11] ),
    .A2(net2277),
    .A1(\draw_game_inst.grid[15] ));
 sg13g2_or2_1 _5939_ (.X(_1495_),
    .B(_1494_),
    .A(net2026));
 sg13g2_a22oi_1 _5940_ (.Y(_1496_),
    .B1(net2019),
    .B2(\draw_game_inst.grid[7] ),
    .A2(net2026),
    .A1(\draw_game_inst.grid[3] ));
 sg13g2_a21oi_1 _5941_ (.A1(_1495_),
    .A2(_1496_),
    .Y(_1497_),
    .B1(_1480_));
 sg13g2_a22oi_1 _5942_ (.Y(_1498_),
    .B1(net2282),
    .B2(\draw_game_inst.grid[27] ),
    .A2(net2279),
    .A1(\draw_game_inst.grid[31] ));
 sg13g2_a22oi_1 _5943_ (.Y(_1499_),
    .B1(net2019),
    .B2(\draw_game_inst.grid[23] ),
    .A2(net2026),
    .A1(\draw_game_inst.grid[19] ));
 sg13g2_o21ai_1 _5944_ (.B1(_1499_),
    .Y(_1500_),
    .A1(net2026),
    .A2(_1498_));
 sg13g2_a21o_1 _5945_ (.A2(_1500_),
    .A1(_1425_),
    .B1(_1497_),
    .X(_1501_));
 sg13g2_a221oi_1 _5946_ (.B2(_1493_),
    .C1(_1501_),
    .B1(_1490_),
    .A1(_1486_),
    .Y(_1502_),
    .A2(_1489_));
 sg13g2_a22oi_1 _5947_ (.Y(_1503_),
    .B1(net2280),
    .B2(\draw_game_inst.grid[58] ),
    .A2(net2279),
    .A1(\draw_game_inst.grid[62] ));
 sg13g2_a22oi_1 _5948_ (.Y(_1504_),
    .B1(net2021),
    .B2(\draw_game_inst.grid[54] ),
    .A2(net2024),
    .A1(\draw_game_inst.grid[50] ));
 sg13g2_o21ai_1 _5949_ (.B1(_1504_),
    .Y(_1505_),
    .A1(net2024),
    .A2(_1503_));
 sg13g2_a22oi_1 _5950_ (.Y(_1506_),
    .B1(net2283),
    .B2(\draw_game_inst.grid[10] ),
    .A2(net2276),
    .A1(\draw_game_inst.grid[14] ));
 sg13g2_or2_1 _5951_ (.X(_1507_),
    .B(_1506_),
    .A(net2024));
 sg13g2_a22oi_1 _5952_ (.Y(_1508_),
    .B1(net2021),
    .B2(\draw_game_inst.grid[6] ),
    .A2(net2024),
    .A1(\draw_game_inst.grid[2] ));
 sg13g2_a21oi_1 _5953_ (.A1(_1507_),
    .A2(_1508_),
    .Y(_1509_),
    .B1(_1480_));
 sg13g2_a22oi_1 _5954_ (.Y(_1510_),
    .B1(net2280),
    .B2(\draw_game_inst.grid[42] ),
    .A2(net2276),
    .A1(\draw_game_inst.grid[46] ));
 sg13g2_a22oi_1 _5955_ (.Y(_1511_),
    .B1(net2021),
    .B2(\draw_game_inst.grid[38] ),
    .A2(net2024),
    .A1(\draw_game_inst.grid[34] ));
 sg13g2_o21ai_1 _5956_ (.B1(_1511_),
    .Y(_1512_),
    .A1(net2024),
    .A2(_1510_));
 sg13g2_a22oi_1 _5957_ (.Y(_1513_),
    .B1(net2283),
    .B2(\draw_game_inst.grid[26] ),
    .A2(net2279),
    .A1(\draw_game_inst.grid[30] ));
 sg13g2_a22oi_1 _5958_ (.Y(_1514_),
    .B1(net2020),
    .B2(\draw_game_inst.grid[22] ),
    .A2(net2027),
    .A1(\draw_game_inst.grid[18] ));
 sg13g2_o21ai_1 _5959_ (.B1(_1514_),
    .Y(_1515_),
    .A1(net2027),
    .A2(_1513_));
 sg13g2_a21o_1 _5960_ (.A2(_1515_),
    .A1(net2031),
    .B1(_1509_),
    .X(_1516_));
 sg13g2_a221oi_1 _5961_ (.B2(_1486_),
    .C1(_1516_),
    .B1(_1512_),
    .A1(_1490_),
    .Y(_1517_),
    .A2(_1505_));
 sg13g2_mux4_1 _5962_ (.S0(net2281),
    .A0(\draw_game_inst.grid[53] ),
    .A1(\draw_game_inst.grid[57] ),
    .A2(\draw_game_inst.grid[61] ),
    .A3(\draw_game_inst.grid[49] ),
    .S1(net2277),
    .X(_1518_));
 sg13g2_nand2_1 _5963_ (.Y(_1519_),
    .A(_1490_),
    .B(_1518_));
 sg13g2_a22oi_1 _5964_ (.Y(_1520_),
    .B1(net2282),
    .B2(\draw_game_inst.grid[25] ),
    .A2(net2278),
    .A1(\draw_game_inst.grid[29] ));
 sg13g2_a22oi_1 _5965_ (.Y(_1521_),
    .B1(net2020),
    .B2(\draw_game_inst.grid[21] ),
    .A2(net2027),
    .A1(\draw_game_inst.grid[17] ));
 sg13g2_o21ai_1 _5966_ (.B1(_1521_),
    .Y(_1522_),
    .A1(net2028),
    .A2(_1520_));
 sg13g2_a22oi_1 _5967_ (.Y(_1523_),
    .B1(net2281),
    .B2(\draw_game_inst.grid[9] ),
    .A2(net2278),
    .A1(\draw_game_inst.grid[13] ));
 sg13g2_or2_1 _5968_ (.X(_1524_),
    .B(_1523_),
    .A(net2026));
 sg13g2_a22oi_1 _5969_ (.Y(_1525_),
    .B1(net2019),
    .B2(\draw_game_inst.grid[5] ),
    .A2(net2026),
    .A1(\draw_game_inst.grid[1] ));
 sg13g2_a21oi_1 _5970_ (.A1(_1524_),
    .A2(_1525_),
    .Y(_1526_),
    .B1(_1480_));
 sg13g2_a21oi_1 _5971_ (.A1(net2031),
    .A2(_1522_),
    .Y(_1527_),
    .B1(_1526_));
 sg13g2_mux4_1 _5972_ (.S0(net2281),
    .A0(\draw_game_inst.grid[37] ),
    .A1(\draw_game_inst.grid[41] ),
    .A2(\draw_game_inst.grid[45] ),
    .A3(\draw_game_inst.grid[33] ),
    .S1(net2277),
    .X(_1528_));
 sg13g2_nand2_1 _5973_ (.Y(_1529_),
    .A(_1486_),
    .B(_1528_));
 sg13g2_and3_1 _5974_ (.X(_1530_),
    .A(_1519_),
    .B(_1527_),
    .C(_1529_));
 sg13g2_nand3_1 _5975_ (.B(_1527_),
    .C(_1529_),
    .A(_1519_),
    .Y(_1531_));
 sg13g2_and2_1 _5976_ (.A(_1502_),
    .B(_1517_),
    .X(_1532_));
 sg13g2_nor2b_1 _5977_ (.A(_1517_),
    .B_N(_1502_),
    .Y(_1533_));
 sg13g2_nand2b_1 _5978_ (.Y(_1534_),
    .B(_1502_),
    .A_N(_1517_));
 sg13g2_nand2b_2 _5979_ (.Y(_1535_),
    .B(_1517_),
    .A_N(_1502_));
 sg13g2_nand2_1 _5980_ (.Y(_1536_),
    .A(_1534_),
    .B(_1535_));
 sg13g2_a21o_1 _5981_ (.A2(_1531_),
    .A1(_1502_),
    .B1(_1536_),
    .X(_1537_));
 sg13g2_a21oi_2 _5982_ (.B1(_1536_),
    .Y(_1538_),
    .A2(_1531_),
    .A1(_1502_));
 sg13g2_nor2b_2 _5983_ (.A(net2290),
    .B_N(\draw_game_inst.board_x[5] ),
    .Y(_1539_));
 sg13g2_nand2b_1 _5984_ (.Y(_1540_),
    .B(net2286),
    .A_N(net2290));
 sg13g2_nor2_1 _5985_ (.A(net2297),
    .B(net2063),
    .Y(_1541_));
 sg13g2_nand2_1 _5986_ (.Y(_1542_),
    .A(net2065),
    .B(net2286));
 sg13g2_nor2_1 _5987_ (.A(net2296),
    .B(net2004),
    .Y(_1543_));
 sg13g2_nand2_1 _5988_ (.Y(_1544_),
    .A(net2065),
    .B(net2006));
 sg13g2_nor2_2 _5989_ (.A(net2296),
    .B(net2290),
    .Y(_1545_));
 sg13g2_nand2_2 _5990_ (.Y(_1546_),
    .A(net2065),
    .B(net2062));
 sg13g2_nor2_1 _5991_ (.A(net2223),
    .B(net1911),
    .Y(_1547_));
 sg13g2_nand2_2 _5992_ (.Y(_1548_),
    .A(net2067),
    .B(net1916));
 sg13g2_nor2_1 _5993_ (.A(net2082),
    .B(net2071),
    .Y(_1549_));
 sg13g2_nand2_2 _5994_ (.Y(_1550_),
    .A(net2210),
    .B(net2236));
 sg13g2_nor2_1 _5995_ (.A(net2195),
    .B(net2082),
    .Y(_1551_));
 sg13g2_nand2_2 _5996_ (.Y(_1552_),
    .A(net2089),
    .B(net2211));
 sg13g2_nor2b_1 _5997_ (.A(net2221),
    .B_N(net2250),
    .Y(_1553_));
 sg13g2_nand2_2 _5998_ (.Y(_1554_),
    .A(net2252),
    .B(net2072));
 sg13g2_nor2_2 _5999_ (.A(net2200),
    .B(net2246),
    .Y(_1555_));
 sg13g2_nand2_2 _6000_ (.Y(_1556_),
    .A(net2087),
    .B(net2069));
 sg13g2_nor2_2 _6001_ (.A(net2236),
    .B(_1475_),
    .Y(_1557_));
 sg13g2_nand2_2 _6002_ (.Y(_1558_),
    .A(net2067),
    .B(net2013));
 sg13g2_a21oi_2 _6003_ (.B1(net2182),
    .Y(_1559_),
    .A2(net2000),
    .A1(net2013));
 sg13g2_nor2_2 _6004_ (.A(_4046_),
    .B(net2289),
    .Y(_1560_));
 sg13g2_nand2_1 _6005_ (.Y(_1561_),
    .A(net2297),
    .B(net2063));
 sg13g2_nor2_2 _6006_ (.A(_4048_),
    .B(net1901),
    .Y(_1562_));
 sg13g2_nand2_1 _6007_ (.Y(_1563_),
    .A(net2063),
    .B(net2018));
 sg13g2_nand2_2 _6008_ (.Y(_1564_),
    .A(net1912),
    .B(net1898));
 sg13g2_nand2_2 _6009_ (.Y(_1565_),
    .A(net2086),
    .B(net1913));
 sg13g2_nand2_1 _6010_ (.Y(_1566_),
    .A(_1559_),
    .B(_1565_));
 sg13g2_nor2_1 _6011_ (.A(net2205),
    .B(net1839),
    .Y(_1567_));
 sg13g2_o21ai_1 _6012_ (.B1(_1559_),
    .Y(_1568_),
    .A1(net1929),
    .A2(_1564_));
 sg13g2_a21oi_1 _6013_ (.A1(_1548_),
    .A2(net1905),
    .Y(_1569_),
    .B1(_1568_));
 sg13g2_nand2b_1 _6014_ (.Y(_1570_),
    .B(net1916),
    .A_N(net2250));
 sg13g2_nor2_1 _6015_ (.A(_0093_),
    .B(net2204),
    .Y(_1571_));
 sg13g2_or2_1 _6016_ (.X(_1572_),
    .B(net2204),
    .A(_0093_));
 sg13g2_o21ai_1 _6017_ (.B1(net2189),
    .Y(_1573_),
    .A1(_1570_),
    .A2(_1572_));
 sg13g2_a21oi_1 _6018_ (.A1(_1569_),
    .A2(_1573_),
    .Y(_1574_),
    .B1(net2180));
 sg13g2_nor2_2 _6019_ (.A(net2091),
    .B(_4042_),
    .Y(_1575_));
 sg13g2_nand2_2 _6020_ (.Y(_1576_),
    .A(net2180),
    .B(net2185));
 sg13g2_nand2_2 _6021_ (.Y(_1577_),
    .A(_1443_),
    .B(net2004));
 sg13g2_nor2_1 _6022_ (.A(net2029),
    .B(_1457_),
    .Y(_1578_));
 sg13g2_nand2_1 _6023_ (.Y(_1579_),
    .A(_1458_),
    .B(_1577_));
 sg13g2_inv_1 _6024_ (.Y(_1580_),
    .A(_1579_));
 sg13g2_nor2_1 _6025_ (.A(net2210),
    .B(net2237),
    .Y(_1581_));
 sg13g2_nand2_2 _6026_ (.Y(_1582_),
    .A(net2079),
    .B(net2068));
 sg13g2_a21oi_1 _6027_ (.A1(net1840),
    .A2(_1580_),
    .Y(_1583_),
    .B1(_1576_));
 sg13g2_and3_2 _6028_ (.X(_1584_),
    .A(net2250),
    .B(_0093_),
    .C(net1916));
 sg13g2_nor2_1 _6029_ (.A(net2107),
    .B(net2076),
    .Y(_1585_));
 sg13g2_nand2_2 _6030_ (.Y(_1586_),
    .A(net2266),
    .B(net2246));
 sg13g2_nor2_1 _6031_ (.A(net1902),
    .B(net1995),
    .Y(_1587_));
 sg13g2_nor2_2 _6032_ (.A(net1897),
    .B(net1993),
    .Y(_1588_));
 sg13g2_nor2_1 _6033_ (.A(_1584_),
    .B(_1588_),
    .Y(_1589_));
 sg13g2_nor2_2 _6034_ (.A(net1946),
    .B(net1838),
    .Y(_1590_));
 sg13g2_a21oi_1 _6035_ (.A1(net2013),
    .A2(net1912),
    .Y(_1591_),
    .B1(_1590_));
 sg13g2_nor2_2 _6036_ (.A(net2085),
    .B(net2079),
    .Y(_1592_));
 sg13g2_nand2_2 _6037_ (.Y(_1593_),
    .A(net2200),
    .B(net2217));
 sg13g2_nor2_1 _6038_ (.A(net2250),
    .B(_0093_),
    .Y(_1594_));
 sg13g2_nand2_1 _6039_ (.Y(_1595_),
    .A(_1580_),
    .B(_1594_));
 sg13g2_a22oi_1 _6040_ (.Y(_1596_),
    .B1(net1885),
    .B2(_1595_),
    .A2(_1589_),
    .A1(net1905));
 sg13g2_a21oi_1 _6041_ (.A1(_1591_),
    .A2(_1596_),
    .Y(_1597_),
    .B1(net1932));
 sg13g2_nor3_1 _6042_ (.A(_1574_),
    .B(_1583_),
    .C(_1597_),
    .Y(_1598_));
 sg13g2_a22oi_1 _6043_ (.Y(_1599_),
    .B1(net2282),
    .B2(\draw_game_inst.grid[24] ),
    .A2(net2278),
    .A1(\draw_game_inst.grid[28] ));
 sg13g2_a22oi_1 _6044_ (.Y(_1600_),
    .B1(net2020),
    .B2(\draw_game_inst.grid[20] ),
    .A2(net2027),
    .A1(\draw_game_inst.grid[16] ));
 sg13g2_o21ai_1 _6045_ (.B1(_1600_),
    .Y(_1601_),
    .A1(net2027),
    .A2(_1599_));
 sg13g2_a22oi_1 _6046_ (.Y(_1602_),
    .B1(net2281),
    .B2(\draw_game_inst.grid[56] ),
    .A2(net2277),
    .A1(\draw_game_inst.grid[60] ));
 sg13g2_a22oi_1 _6047_ (.Y(_1603_),
    .B1(net2019),
    .B2(\draw_game_inst.grid[52] ),
    .A2(net2025),
    .A1(\draw_game_inst.grid[48] ));
 sg13g2_o21ai_1 _6048_ (.B1(_1603_),
    .Y(_1604_),
    .A1(net2025),
    .A2(_1602_));
 sg13g2_a22oi_1 _6049_ (.Y(_1605_),
    .B1(net2281),
    .B2(\draw_game_inst.grid[8] ),
    .A2(net2277),
    .A1(\draw_game_inst.grid[12] ));
 sg13g2_or2_1 _6050_ (.X(_1606_),
    .B(_1605_),
    .A(net2026));
 sg13g2_a22oi_1 _6051_ (.Y(_1607_),
    .B1(net2019),
    .B2(\draw_game_inst.grid[4] ),
    .A2(net2026),
    .A1(\draw_game_inst.grid[0] ));
 sg13g2_a21oi_1 _6052_ (.A1(_1606_),
    .A2(_1607_),
    .Y(_1608_),
    .B1(_1480_));
 sg13g2_a22oi_1 _6053_ (.Y(_1609_),
    .B1(net2281),
    .B2(\draw_game_inst.grid[40] ),
    .A2(net2277),
    .A1(\draw_game_inst.grid[44] ));
 sg13g2_a22oi_1 _6054_ (.Y(_1610_),
    .B1(net2019),
    .B2(\draw_game_inst.grid[36] ),
    .A2(net2025),
    .A1(\draw_game_inst.grid[32] ));
 sg13g2_o21ai_1 _6055_ (.B1(_1610_),
    .Y(_1611_),
    .A1(net2025),
    .A2(_1609_));
 sg13g2_a21o_1 _6056_ (.A2(_1601_),
    .A1(net2031),
    .B1(_1608_),
    .X(_1612_));
 sg13g2_a221oi_1 _6057_ (.B2(_1486_),
    .C1(_1612_),
    .B1(_1611_),
    .A1(_1490_),
    .Y(_1613_),
    .A2(_1604_));
 sg13g2_nor2_2 _6058_ (.A(_1531_),
    .B(_1613_),
    .Y(_1614_));
 sg13g2_and2_2 _6059_ (.A(_1533_),
    .B(_1614_),
    .X(_1615_));
 sg13g2_nor2_1 _6060_ (.A(net2298),
    .B(net2062),
    .Y(_1616_));
 sg13g2_nand2_1 _6061_ (.Y(_1617_),
    .A(net2065),
    .B(net2290));
 sg13g2_nor2_1 _6062_ (.A(_0094_),
    .B(net1879),
    .Y(_1618_));
 sg13g2_nand2_2 _6063_ (.Y(_1619_),
    .A(_4055_),
    .B(net1882));
 sg13g2_nor2_2 _6064_ (.A(net2266),
    .B(net1881),
    .Y(_1620_));
 sg13g2_nor2_1 _6065_ (.A(net2297),
    .B(_1443_),
    .Y(_1621_));
 sg13g2_nand2_1 _6066_ (.Y(_1622_),
    .A(net2065),
    .B(net2022));
 sg13g2_nand2_1 _6067_ (.Y(_1623_),
    .A(net2262),
    .B(net1875));
 sg13g2_a21oi_2 _6068_ (.B1(net1879),
    .Y(_1624_),
    .A2(net2288),
    .A1(net2263));
 sg13g2_nor2_2 _6069_ (.A(net2235),
    .B(_1624_),
    .Y(_1625_));
 sg13g2_nor2_1 _6070_ (.A(net2225),
    .B(net1836),
    .Y(_1626_));
 sg13g2_nand2_2 _6071_ (.Y(_1627_),
    .A(_1619_),
    .B(_1625_));
 sg13g2_nor2_2 _6072_ (.A(net2212),
    .B(_1627_),
    .Y(_1628_));
 sg13g2_nor2_1 _6073_ (.A(net2065),
    .B(net2290),
    .Y(_1629_));
 sg13g2_nand2_1 _6074_ (.Y(_1630_),
    .A(net2296),
    .B(net2062));
 sg13g2_nand2_1 _6075_ (.Y(_1631_),
    .A(net2299),
    .B(_4055_));
 sg13g2_nor2_2 _6076_ (.A(net2284),
    .B(net1869),
    .Y(_1632_));
 sg13g2_nand2_1 _6077_ (.Y(_1633_),
    .A(_4055_),
    .B(net1871));
 sg13g2_nand2_2 _6078_ (.Y(_1634_),
    .A(_1554_),
    .B(net1834));
 sg13g2_a21oi_2 _6079_ (.B1(net2188),
    .Y(_1635_),
    .A2(_1634_),
    .A1(net2207));
 sg13g2_nor2_1 _6080_ (.A(net2210),
    .B(net2071),
    .Y(_1636_));
 sg13g2_nand2_2 _6081_ (.Y(_1637_),
    .A(net2233),
    .B(net1873));
 sg13g2_a21oi_1 _6082_ (.A1(net1874),
    .A2(net1866),
    .Y(_1638_),
    .B1(_1628_));
 sg13g2_nor2_2 _6083_ (.A(net1922),
    .B(net1903),
    .Y(_1639_));
 sg13g2_nand2_2 _6084_ (.Y(_1640_),
    .A(net1921),
    .B(net1901));
 sg13g2_nor2_1 _6085_ (.A(net2293),
    .B(net1901),
    .Y(_1641_));
 sg13g2_nand2_2 _6086_ (.Y(_1642_),
    .A(_4048_),
    .B(net1903));
 sg13g2_nand2_1 _6087_ (.Y(_1643_),
    .A(net1914),
    .B(_1642_));
 sg13g2_nor2_2 _6088_ (.A(net1919),
    .B(net1830),
    .Y(_1644_));
 sg13g2_nor2_1 _6089_ (.A(net1881),
    .B(net1872),
    .Y(_1645_));
 sg13g2_nand2_1 _6090_ (.Y(_1646_),
    .A(net1879),
    .B(net1870));
 sg13g2_nand2_2 _6091_ (.Y(_1647_),
    .A(net2263),
    .B(net2005));
 sg13g2_nor2_2 _6092_ (.A(net2107),
    .B(net1922),
    .Y(_1648_));
 sg13g2_nand2_2 _6093_ (.Y(_1649_),
    .A(net2253),
    .B(net1920));
 sg13g2_nor2_1 _6094_ (.A(net1826),
    .B(_1649_),
    .Y(_1650_));
 sg13g2_a21oi_1 _6095_ (.A1(net2110),
    .A2(_1644_),
    .Y(_1651_),
    .B1(_1650_));
 sg13g2_nand2_1 _6096_ (.Y(_1652_),
    .A(net2234),
    .B(_1651_));
 sg13g2_o21ai_1 _6097_ (.B1(_1652_),
    .Y(_1653_),
    .A1(net2252),
    .A2(_1548_));
 sg13g2_nor2_2 _6098_ (.A(net2210),
    .B(net1892),
    .Y(_1654_));
 sg13g2_nand2_2 _6099_ (.Y(_1655_),
    .A(net2083),
    .B(net1994));
 sg13g2_nor2_1 _6100_ (.A(net2090),
    .B(net1890),
    .Y(_1656_));
 sg13g2_nor2_2 _6101_ (.A(net1946),
    .B(net1892),
    .Y(_1657_));
 sg13g2_nand2_2 _6102_ (.Y(_1658_),
    .A(net1947),
    .B(net1991));
 sg13g2_a221oi_1 _6103_ (.B2(net1886),
    .C1(net2185),
    .B1(_1653_),
    .A1(_1635_),
    .Y(_1659_),
    .A2(_1638_));
 sg13g2_o21ai_1 _6104_ (.B1(_1659_),
    .Y(_1660_),
    .A1(net1833),
    .A2(_1658_));
 sg13g2_nand2_1 _6105_ (.Y(_1661_),
    .A(net1772),
    .B(_1660_));
 sg13g2_and2_2 _6106_ (.A(_1531_),
    .B(_1613_),
    .X(_1662_));
 sg13g2_nor2b_2 _6107_ (.A(_1535_),
    .B_N(_1662_),
    .Y(_1663_));
 sg13g2_o21ai_1 _6108_ (.B1(_1657_),
    .Y(_1664_),
    .A1(net2007),
    .A2(_1637_));
 sg13g2_nor2_2 _6109_ (.A(net2253),
    .B(net2066),
    .Y(_1665_));
 sg13g2_nand2_2 _6110_ (.Y(_1666_),
    .A(net2110),
    .B(net2297));
 sg13g2_nor2_2 _6111_ (.A(net2254),
    .B(net2006),
    .Y(_1667_));
 sg13g2_nand2_2 _6112_ (.Y(_1668_),
    .A(net2110),
    .B(net1915));
 sg13g2_nor2_1 _6113_ (.A(net1918),
    .B(net1877),
    .Y(_1669_));
 sg13g2_nand2_2 _6114_ (.Y(_1670_),
    .A(net1915),
    .B(net1873));
 sg13g2_nor2_1 _6115_ (.A(net2260),
    .B(_1670_),
    .Y(_1671_));
 sg13g2_nor2_1 _6116_ (.A(net1876),
    .B(_1647_),
    .Y(_1672_));
 sg13g2_a21oi_1 _6117_ (.A1(_1647_),
    .A2(_1668_),
    .Y(_1673_),
    .B1(net1876));
 sg13g2_a21oi_1 _6118_ (.A1(net2073),
    .A2(_1673_),
    .Y(_1674_),
    .B1(_1664_));
 sg13g2_nor2_2 _6119_ (.A(_1567_),
    .B(net1996),
    .Y(_1675_));
 sg13g2_nor2_2 _6120_ (.A(net2298),
    .B(_1437_),
    .Y(_1676_));
 sg13g2_nand2_1 _6121_ (.Y(_1677_),
    .A(net2293),
    .B(net1922));
 sg13g2_nand2_2 _6122_ (.Y(_1678_),
    .A(net2293),
    .B(_1640_));
 sg13g2_inv_1 _6123_ (.Y(_1679_),
    .A(net1814));
 sg13g2_nand2_1 _6124_ (.Y(_1680_),
    .A(net2262),
    .B(net1814));
 sg13g2_nor2_2 _6125_ (.A(net2007),
    .B(net1922),
    .Y(_1681_));
 sg13g2_nor2_2 _6126_ (.A(net2063),
    .B(net2018),
    .Y(_1682_));
 sg13g2_nor2_2 _6127_ (.A(_1545_),
    .B(_1681_),
    .Y(_1683_));
 sg13g2_nand2_2 _6128_ (.Y(_1684_),
    .A(net2289),
    .B(net1825));
 sg13g2_nor2_2 _6129_ (.A(net2261),
    .B(net1838),
    .Y(_1685_));
 sg13g2_nand2_2 _6130_ (.Y(_1686_),
    .A(net2106),
    .B(net1898));
 sg13g2_o21ai_1 _6131_ (.B1(_1680_),
    .Y(_1687_),
    .A1(_1683_),
    .A2(_1686_));
 sg13g2_nor2_1 _6132_ (.A(net2235),
    .B(_1687_),
    .Y(_1688_));
 sg13g2_nand2_1 _6133_ (.Y(_1689_),
    .A(net2289),
    .B(_0096_));
 sg13g2_nor2_2 _6134_ (.A(net2297),
    .B(net2287),
    .Y(_1690_));
 sg13g2_nand2_2 _6135_ (.Y(_1691_),
    .A(net2064),
    .B(_1460_));
 sg13g2_and2_2 _6136_ (.A(_1689_),
    .B(_1691_),
    .X(_1692_));
 sg13g2_nand2_2 _6137_ (.Y(_1693_),
    .A(net2223),
    .B(net2290));
 sg13g2_nor2_2 _6138_ (.A(net2072),
    .B(net1923),
    .Y(_1694_));
 sg13g2_nor2_2 _6139_ (.A(net2067),
    .B(net1916),
    .Y(_1695_));
 sg13g2_nand2_1 _6140_ (.Y(_1696_),
    .A(net1900),
    .B(_1695_));
 sg13g2_o21ai_1 _6141_ (.B1(_1696_),
    .Y(_1697_),
    .A1(net2235),
    .A2(_1692_));
 sg13g2_a21oi_1 _6142_ (.A1(net2214),
    .A2(_1697_),
    .Y(_1698_),
    .B1(net2194));
 sg13g2_o21ai_1 _6143_ (.B1(_1698_),
    .Y(_1699_),
    .A1(_1675_),
    .A2(_1688_));
 sg13g2_nand2b_1 _6144_ (.Y(_1700_),
    .B(_1699_),
    .A_N(_1674_));
 sg13g2_nor2_2 _6145_ (.A(_1530_),
    .B(_1613_),
    .Y(_1701_));
 sg13g2_nor2b_2 _6146_ (.A(_1535_),
    .B_N(_1701_),
    .Y(_1702_));
 sg13g2_nand2b_2 _6147_ (.Y(_1703_),
    .B(_1701_),
    .A_N(_1535_));
 sg13g2_nand2_1 _6148_ (.Y(_1704_),
    .A(net2265),
    .B(net2030));
 sg13g2_nor2_1 _6149_ (.A(net2231),
    .B(net1903),
    .Y(_1705_));
 sg13g2_nand2_1 _6150_ (.Y(_1706_),
    .A(net1921),
    .B(_1705_));
 sg13g2_a21oi_1 _6151_ (.A1(_1640_),
    .A2(_1704_),
    .Y(_1707_),
    .B1(net2240));
 sg13g2_nand2_2 _6152_ (.Y(_1708_),
    .A(net2109),
    .B(net2287));
 sg13g2_nor2_1 _6153_ (.A(net2215),
    .B(_1460_),
    .Y(_1709_));
 sg13g2_a21oi_2 _6154_ (.B1(net1997),
    .Y(_1710_),
    .A2(_1709_),
    .A1(_1708_));
 sg13g2_nor3_1 _6155_ (.A(net2202),
    .B(_1707_),
    .C(_1710_),
    .Y(_1711_));
 sg13g2_nor2_2 _6156_ (.A(net1925),
    .B(net1985),
    .Y(_1712_));
 sg13g2_nand2_2 _6157_ (.Y(_1713_),
    .A(_1460_),
    .B(net2005));
 sg13g2_o21ai_1 _6158_ (.B1(net2242),
    .Y(_1714_),
    .A1(net2265),
    .A2(_1713_));
 sg13g2_nand2_2 _6159_ (.Y(_1715_),
    .A(net2265),
    .B(net1880));
 sg13g2_nor2_2 _6160_ (.A(net2224),
    .B(net2029),
    .Y(_1716_));
 sg13g2_a221oi_1 _6161_ (.B2(net1927),
    .C1(net1824),
    .B1(_1713_),
    .A1(_1461_),
    .Y(_1717_),
    .A2(_1712_));
 sg13g2_nor2b_1 _6162_ (.A(net2292),
    .B_N(net2285),
    .Y(_1718_));
 sg13g2_a21oi_2 _6163_ (.B1(_1718_),
    .Y(_1719_),
    .A2(net2295),
    .A1(net2292));
 sg13g2_o21ai_1 _6164_ (.B1(net1907),
    .Y(_1720_),
    .A1(net2241),
    .A2(_1719_));
 sg13g2_nand2_2 _6165_ (.Y(_1721_),
    .A(net2062),
    .B(net1985));
 sg13g2_nand2_1 _6166_ (.Y(_1722_),
    .A(net2230),
    .B(_1460_));
 sg13g2_nor2b_1 _6167_ (.A(_1722_),
    .B_N(_1721_),
    .Y(_1723_));
 sg13g2_nor2_1 _6168_ (.A(_1711_),
    .B(_1717_),
    .Y(_1724_));
 sg13g2_o21ai_1 _6169_ (.B1(_1724_),
    .Y(_1725_),
    .A1(_1720_),
    .A2(_1723_));
 sg13g2_a22oi_1 _6170_ (.Y(_1726_),
    .B1(_1702_),
    .B2(_1725_),
    .A2(_1700_),
    .A1(net1771));
 sg13g2_o21ai_1 _6171_ (.B1(_1661_),
    .Y(_1727_),
    .A1(net2185),
    .A2(_1726_));
 sg13g2_nor2_2 _6172_ (.A(net2228),
    .B(net2017),
    .Y(_1728_));
 sg13g2_nand2_1 _6173_ (.Y(_1729_),
    .A(net2070),
    .B(_1460_));
 sg13g2_nand3_1 _6174_ (.B(_1721_),
    .C(_1728_),
    .A(net2016),
    .Y(_1730_));
 sg13g2_and2_1 _6175_ (.A(net2185),
    .B(_1730_),
    .X(_1731_));
 sg13g2_nand3b_1 _6176_ (.B(net2180),
    .C(_1727_),
    .Y(_1732_),
    .A_N(_1731_));
 sg13g2_and2_2 _6177_ (.A(_1533_),
    .B(_1701_),
    .X(_1733_));
 sg13g2_nand2_1 _6178_ (.Y(_1734_),
    .A(net2246),
    .B(net1870));
 sg13g2_nor2_2 _6179_ (.A(net2246),
    .B(net1830),
    .Y(_1735_));
 sg13g2_nand2_2 _6180_ (.Y(_1736_),
    .A(net2076),
    .B(_1642_));
 sg13g2_nor2_2 _6181_ (.A(net2266),
    .B(_1677_),
    .Y(_1737_));
 sg13g2_nand2b_1 _6182_ (.Y(_1738_),
    .B(_1735_),
    .A_N(_1737_));
 sg13g2_a21oi_1 _6183_ (.A1(_1734_),
    .A2(_1738_),
    .Y(_1739_),
    .B1(net1931));
 sg13g2_nor2b_2 _6184_ (.A(net2288),
    .B_N(_0095_),
    .Y(_1740_));
 sg13g2_nand2_2 _6185_ (.Y(_1741_),
    .A(net2063),
    .B(net2295));
 sg13g2_nand2_1 _6186_ (.Y(_1742_),
    .A(net1921),
    .B(_1741_));
 sg13g2_nor2_2 _6187_ (.A(_1436_),
    .B(_1742_),
    .Y(_1743_));
 sg13g2_nand3_1 _6188_ (.B(net1921),
    .C(_1741_),
    .A(_1437_),
    .Y(_1744_));
 sg13g2_nand2_2 _6189_ (.Y(_1745_),
    .A(net2107),
    .B(_1744_));
 sg13g2_nor2_2 _6190_ (.A(net2107),
    .B(net1872),
    .Y(_1746_));
 sg13g2_nor2_1 _6191_ (.A(net2245),
    .B(_1746_),
    .Y(_1747_));
 sg13g2_nand2_2 _6192_ (.Y(_1748_),
    .A(net2261),
    .B(net1902));
 sg13g2_nand2_2 _6193_ (.Y(_1749_),
    .A(net1901),
    .B(_1648_));
 sg13g2_nor2_2 _6194_ (.A(net2266),
    .B(net1872),
    .Y(_1750_));
 sg13g2_nor2_1 _6195_ (.A(net2075),
    .B(_1750_),
    .Y(_1751_));
 sg13g2_a221oi_1 _6196_ (.B2(_1751_),
    .C1(net1944),
    .B1(_1749_),
    .A1(_1745_),
    .Y(_1752_),
    .A2(_1747_));
 sg13g2_a21oi_1 _6197_ (.A1(net2011),
    .A2(_1640_),
    .Y(_1753_),
    .B1(net1990));
 sg13g2_nor2_1 _6198_ (.A(net1936),
    .B(_1753_),
    .Y(_1754_));
 sg13g2_nor2_1 _6199_ (.A(net2011),
    .B(_1744_),
    .Y(_1755_));
 sg13g2_o21ai_1 _6200_ (.B1(net1908),
    .Y(_1756_),
    .A1(net1926),
    .A2(net1870));
 sg13g2_o21ai_1 _6201_ (.B1(_1754_),
    .Y(_1757_),
    .A1(_1755_),
    .A2(_1756_));
 sg13g2_nor3_1 _6202_ (.A(_1739_),
    .B(_1752_),
    .C(_1757_),
    .Y(_1758_));
 sg13g2_nor2_1 _6203_ (.A(net2179),
    .B(net2182),
    .Y(_1759_));
 sg13g2_or2_1 _6204_ (.X(_1760_),
    .B(net2182),
    .A(net2179));
 sg13g2_nor2_2 _6205_ (.A(net2086),
    .B(net1980),
    .Y(_1761_));
 sg13g2_nand2_1 _6206_ (.Y(_1762_),
    .A(net2201),
    .B(net1984));
 sg13g2_nor2_1 _6207_ (.A(net2267),
    .B(_1560_),
    .Y(_1763_));
 sg13g2_nand2_2 _6208_ (.Y(_1764_),
    .A(net2108),
    .B(net1901));
 sg13g2_nand2_1 _6209_ (.Y(_1765_),
    .A(net2264),
    .B(_1644_));
 sg13g2_o21ai_1 _6210_ (.B1(_1765_),
    .Y(_1766_),
    .A1(net1919),
    .A2(_1764_));
 sg13g2_nand2_2 _6211_ (.Y(_1767_),
    .A(net2240),
    .B(_1766_));
 sg13g2_nor2_2 _6212_ (.A(_1457_),
    .B(net2007),
    .Y(_1768_));
 sg13g2_nor3_2 _6213_ (.A(_1457_),
    .B(net2006),
    .C(_1740_),
    .Y(_1769_));
 sg13g2_nand2_2 _6214_ (.Y(_1770_),
    .A(_1741_),
    .B(_1768_));
 sg13g2_nand2_2 _6215_ (.Y(_1771_),
    .A(net2107),
    .B(_1770_));
 sg13g2_a21o_1 _6216_ (.A2(_1771_),
    .A1(_1749_),
    .B1(net2245),
    .X(_1772_));
 sg13g2_nor2_1 _6217_ (.A(net2203),
    .B(net1981),
    .Y(_1773_));
 sg13g2_nand3_1 _6218_ (.B(_1772_),
    .C(net1862),
    .A(_1767_),
    .Y(_1774_));
 sg13g2_and2_2 _6219_ (.A(net2265),
    .B(net1985),
    .X(_1775_));
 sg13g2_a21oi_1 _6220_ (.A1(net1893),
    .A2(_1690_),
    .Y(_1776_),
    .B1(net2292));
 sg13g2_nand2_1 _6221_ (.Y(_1777_),
    .A(net1923),
    .B(net1892));
 sg13g2_nand3_1 _6222_ (.B(_1644_),
    .C(_1777_),
    .A(net1886),
    .Y(_1778_));
 sg13g2_o21ai_1 _6223_ (.B1(_1778_),
    .Y(_1779_),
    .A1(net1945),
    .A2(_1776_));
 sg13g2_a21oi_1 _6224_ (.A1(net1864),
    .A2(_1774_),
    .Y(_1780_),
    .B1(_1779_));
 sg13g2_o21ai_1 _6225_ (.B1(_1733_),
    .Y(_1781_),
    .A1(_1758_),
    .A2(_1780_));
 sg13g2_nand2b_2 _6226_ (.Y(_1782_),
    .B(_1614_),
    .A_N(_1535_));
 sg13g2_nor2_1 _6227_ (.A(_4055_),
    .B(net1911),
    .Y(_1783_));
 sg13g2_nand2_1 _6228_ (.Y(_1784_),
    .A(net2284),
    .B(_1545_));
 sg13g2_nor2_1 _6229_ (.A(net2297),
    .B(net2029),
    .Y(_1785_));
 sg13g2_nand2_2 _6230_ (.Y(_1786_),
    .A(_4046_),
    .B(_1435_));
 sg13g2_nor2_2 _6231_ (.A(_1442_),
    .B(net1985),
    .Y(_1787_));
 sg13g2_nor2_2 _6232_ (.A(net2287),
    .B(net1872),
    .Y(_1788_));
 sg13g2_nor2_2 _6233_ (.A(net2066),
    .B(_1577_),
    .Y(_1789_));
 sg13g2_nand2_2 _6234_ (.Y(_1790_),
    .A(_1681_),
    .B(_1787_));
 sg13g2_o21ai_1 _6235_ (.B1(net2008),
    .Y(_1791_),
    .A1(net1858),
    .A2(_1789_));
 sg13g2_nand2_2 _6236_ (.Y(_1792_),
    .A(net1924),
    .B(net1832));
 sg13g2_a21oi_2 _6237_ (.B1(net1942),
    .Y(_1793_),
    .A2(_1792_),
    .A1(_1791_));
 sg13g2_o21ai_1 _6238_ (.B1(net1947),
    .Y(_1794_),
    .A1(net2008),
    .A2(net1860));
 sg13g2_o21ai_1 _6239_ (.B1(_1793_),
    .Y(_1795_),
    .A1(net2008),
    .A2(net1860));
 sg13g2_nand2_1 _6240_ (.Y(_1796_),
    .A(net2064),
    .B(net1829));
 sg13g2_a22oi_1 _6241_ (.Y(_1797_),
    .B1(_1796_),
    .B2(net2231),
    .A2(_1716_),
    .A1(net1821));
 sg13g2_a21oi_1 _6242_ (.A1(net1862),
    .A2(_1797_),
    .Y(_1798_),
    .B1(_1761_));
 sg13g2_nor2_1 _6243_ (.A(net2069),
    .B(net2029),
    .Y(_1799_));
 sg13g2_nor2_1 _6244_ (.A(net2266),
    .B(net2076),
    .Y(_1800_));
 sg13g2_nand2_2 _6245_ (.Y(_1801_),
    .A(net2104),
    .B(net2227));
 sg13g2_nor2_2 _6246_ (.A(net2030),
    .B(_1801_),
    .Y(_1802_));
 sg13g2_nand2_1 _6247_ (.Y(_1803_),
    .A(_1435_),
    .B(net1857));
 sg13g2_nor2_2 _6248_ (.A(net2070),
    .B(net1820),
    .Y(_1804_));
 sg13g2_nand2_2 _6249_ (.Y(_1805_),
    .A(net2231),
    .B(net1860));
 sg13g2_o21ai_1 _6250_ (.B1(_1803_),
    .Y(_1806_),
    .A1(net1992),
    .A2(_1783_));
 sg13g2_o21ai_1 _6251_ (.B1(net1884),
    .Y(_1807_),
    .A1(_1716_),
    .A2(_1806_));
 sg13g2_nand2_1 _6252_ (.Y(_1808_),
    .A(_1795_),
    .B(_1807_));
 sg13g2_nor2_2 _6253_ (.A(net2261),
    .B(net1923),
    .Y(_1809_));
 sg13g2_nand2_2 _6254_ (.Y(_1810_),
    .A(net2105),
    .B(net1920));
 sg13g2_nand2_1 _6255_ (.Y(_1811_),
    .A(net2225),
    .B(_1810_));
 sg13g2_nand2_2 _6256_ (.Y(_1812_),
    .A(net2289),
    .B(net1829));
 sg13g2_nor2_2 _6257_ (.A(net2107),
    .B(net2022),
    .Y(_1813_));
 sg13g2_a22oi_1 _6258_ (.Y(_1814_),
    .B1(_1812_),
    .B2(_1813_),
    .A2(_1811_),
    .A1(_1693_));
 sg13g2_nand2_1 _6259_ (.Y(_1815_),
    .A(net1947),
    .B(_1814_));
 sg13g2_nor2_2 _6260_ (.A(net2250),
    .B(net2067),
    .Y(_1816_));
 sg13g2_nand2b_1 _6261_ (.Y(_1817_),
    .B(net2237),
    .A_N(net2252));
 sg13g2_nor2_1 _6262_ (.A(net2221),
    .B(net1835),
    .Y(_1818_));
 sg13g2_a21oi_1 _6263_ (.A1(net1820),
    .A2(_1816_),
    .Y(_1819_),
    .B1(_1818_));
 sg13g2_nor2_1 _6264_ (.A(net2074),
    .B(net2292),
    .Y(_1820_));
 sg13g2_o21ai_1 _6265_ (.B1(net2242),
    .Y(_1821_),
    .A1(net2297),
    .A2(_0094_));
 sg13g2_nor2_2 _6266_ (.A(net2068),
    .B(net1836),
    .Y(_1822_));
 sg13g2_nand2_1 _6267_ (.Y(_1823_),
    .A(net1825),
    .B(_1712_));
 sg13g2_a22oi_1 _6268_ (.Y(_1824_),
    .B1(_1822_),
    .B2(net2014),
    .A2(net1859),
    .A1(net1997));
 sg13g2_a22oi_1 _6269_ (.Y(_1825_),
    .B1(_1823_),
    .B2(net1884),
    .A2(_1819_),
    .A1(net1905));
 sg13g2_nand4_1 _6270_ (.B(_1815_),
    .C(_1824_),
    .A(net1937),
    .Y(_1826_),
    .D(_1825_));
 sg13g2_o21ai_1 _6271_ (.B1(_1826_),
    .Y(_1827_),
    .A1(_1798_),
    .A2(_1808_));
 sg13g2_nand2b_1 _6272_ (.Y(_1828_),
    .B(_1827_),
    .A_N(_1782_));
 sg13g2_and2_2 _6273_ (.A(_1532_),
    .B(_1662_),
    .X(_1829_));
 sg13g2_o21ai_1 _6274_ (.B1(_1575_),
    .Y(_1830_),
    .A1(net1913),
    .A2(_1558_));
 sg13g2_and2_1 _6275_ (.A(_1829_),
    .B(_1830_),
    .X(_1831_));
 sg13g2_nand2_2 _6276_ (.Y(_1832_),
    .A(net2189),
    .B(net1912));
 sg13g2_a21o_1 _6277_ (.A2(net1996),
    .A1(_1580_),
    .B1(_1832_),
    .X(_1833_));
 sg13g2_nor2_2 _6278_ (.A(net2195),
    .B(net2002),
    .Y(_1834_));
 sg13g2_a21oi_1 _6279_ (.A1(net1918),
    .A2(net2003),
    .Y(_1835_),
    .B1(net2190));
 sg13g2_nand2_1 _6280_ (.Y(_1836_),
    .A(_1580_),
    .B(_1666_));
 sg13g2_o21ai_1 _6281_ (.B1(_1835_),
    .Y(_1837_),
    .A1(net2003),
    .A2(_1836_));
 sg13g2_a21oi_1 _6282_ (.A1(_1833_),
    .A2(_1837_),
    .Y(_1838_),
    .B1(net1935));
 sg13g2_nand2_2 _6283_ (.Y(_1839_),
    .A(_1560_),
    .B(_1693_));
 sg13g2_o21ai_1 _6284_ (.B1(_1564_),
    .Y(_1840_),
    .A1(net1943),
    .A2(_1839_));
 sg13g2_o21ai_1 _6285_ (.B1(net2093),
    .Y(_1841_),
    .A1(_1566_),
    .A2(_1840_));
 sg13g2_nand2_1 _6286_ (.Y(_1842_),
    .A(_1831_),
    .B(_1841_));
 sg13g2_nor2_1 _6287_ (.A(_1838_),
    .B(_1842_),
    .Y(_1843_));
 sg13g2_nand2_2 _6288_ (.Y(_1844_),
    .A(net2261),
    .B(net1876));
 sg13g2_inv_1 _6289_ (.Y(_1845_),
    .A(_1844_));
 sg13g2_a22oi_1 _6290_ (.Y(_1846_),
    .B1(net1902),
    .B2(_1437_),
    .A2(net2022),
    .A1(net2260));
 sg13g2_o21ai_1 _6291_ (.B1(net1866),
    .Y(_1847_),
    .A1(_1845_),
    .A2(_1846_));
 sg13g2_nor2_1 _6292_ (.A(net2217),
    .B(net1877),
    .Y(_1848_));
 sg13g2_nand2_1 _6293_ (.Y(_1849_),
    .A(net2257),
    .B(_1545_));
 sg13g2_nand2_2 _6294_ (.Y(_1850_),
    .A(net2261),
    .B(net1918));
 sg13g2_nand3_1 _6295_ (.B(net1873),
    .C(_1850_),
    .A(net1998),
    .Y(_1851_));
 sg13g2_nand3_1 _6296_ (.B(_1680_),
    .C(_1686_),
    .A(net2235),
    .Y(_1852_));
 sg13g2_a21oi_2 _6297_ (.B1(net2066),
    .Y(_1853_),
    .A2(net2004),
    .A1(_1443_));
 sg13g2_nand2_2 _6298_ (.Y(_1854_),
    .A(net2300),
    .B(_1577_));
 sg13g2_nand3_1 _6299_ (.B(_1852_),
    .C(_1854_),
    .A(net2214),
    .Y(_1855_));
 sg13g2_nor2_2 _6300_ (.A(_0091_),
    .B(net1981),
    .Y(_1856_));
 sg13g2_nand2b_2 _6301_ (.Y(_1857_),
    .B(net1983),
    .A_N(_0091_));
 sg13g2_nand2_1 _6302_ (.Y(_1858_),
    .A(net1771),
    .B(_1856_));
 sg13g2_nand2_2 _6303_ (.Y(_1859_),
    .A(_1530_),
    .B(_1613_));
 sg13g2_nor2_2 _6304_ (.A(_1534_),
    .B(_1859_),
    .Y(_1860_));
 sg13g2_or2_2 _6305_ (.X(_1861_),
    .B(_1859_),
    .A(_1534_));
 sg13g2_nor2_2 _6306_ (.A(net2247),
    .B(net1877),
    .Y(_1862_));
 sg13g2_nor2_2 _6307_ (.A(net2001),
    .B(_1862_),
    .Y(_1863_));
 sg13g2_nor2_2 _6308_ (.A(net2294),
    .B(_1458_),
    .Y(_1864_));
 sg13g2_nand2_2 _6309_ (.Y(_1865_),
    .A(_4048_),
    .B(_1457_));
 sg13g2_nor2_2 _6310_ (.A(net1878),
    .B(_1864_),
    .Y(_1866_));
 sg13g2_nand2_2 _6311_ (.Y(_1867_),
    .A(net1875),
    .B(net1818));
 sg13g2_o21ai_1 _6312_ (.B1(net2071),
    .Y(_1868_),
    .A1(net2252),
    .A2(_1866_));
 sg13g2_or2_1 _6313_ (.X(_1869_),
    .B(_1868_),
    .A(net2210));
 sg13g2_nor2_1 _6314_ (.A(_1715_),
    .B(_1864_),
    .Y(_1870_));
 sg13g2_nor2_2 _6315_ (.A(net2260),
    .B(_1867_),
    .Y(_1871_));
 sg13g2_o21ai_1 _6316_ (.B1(net1865),
    .Y(_1872_),
    .A1(_1870_),
    .A2(_1871_));
 sg13g2_a21o_1 _6317_ (.A2(_1872_),
    .A1(_1869_),
    .B1(net2194),
    .X(_1873_));
 sg13g2_nor2_1 _6318_ (.A(net2236),
    .B(net1858),
    .Y(_1874_));
 sg13g2_nand2_2 _6319_ (.Y(_1875_),
    .A(net2107),
    .B(net1831));
 sg13g2_a22oi_1 _6320_ (.Y(_1876_),
    .B1(_1874_),
    .B2(_1875_),
    .A2(net1822),
    .A1(net2236));
 sg13g2_nor2_1 _6321_ (.A(net1946),
    .B(_1876_),
    .Y(_1877_));
 sg13g2_nor2_1 _6322_ (.A(net2082),
    .B(net2236),
    .Y(_1878_));
 sg13g2_nand2_2 _6323_ (.Y(_1879_),
    .A(net2211),
    .B(net2071));
 sg13g2_nand2_2 _6324_ (.Y(_1880_),
    .A(net2071),
    .B(net1886));
 sg13g2_nor3_1 _6325_ (.A(net2007),
    .B(net1876),
    .C(_1880_),
    .Y(_1881_));
 sg13g2_or2_2 _6326_ (.X(_1882_),
    .B(_1718_),
    .A(net2018));
 sg13g2_nor2_2 _6327_ (.A(net2068),
    .B(net1987),
    .Y(_1883_));
 sg13g2_nand2_2 _6328_ (.Y(_1884_),
    .A(net2233),
    .B(net1886));
 sg13g2_a22oi_1 _6329_ (.Y(_1885_),
    .B1(net1855),
    .B2(_1882_),
    .A2(_1786_),
    .A1(net1892));
 sg13g2_nor2_1 _6330_ (.A(net1989),
    .B(_1885_),
    .Y(_1886_));
 sg13g2_nor3_1 _6331_ (.A(_1877_),
    .B(_1881_),
    .C(_1886_),
    .Y(_1887_));
 sg13g2_nor2_2 _6332_ (.A(net2007),
    .B(net1827),
    .Y(_1888_));
 sg13g2_nand2_2 _6333_ (.Y(_1889_),
    .A(net2011),
    .B(_1888_));
 sg13g2_nor2_2 _6334_ (.A(net2196),
    .B(_1879_),
    .Y(_1890_));
 sg13g2_nand3_1 _6335_ (.B(net1879),
    .C(_1644_),
    .A(net1907),
    .Y(_1891_));
 sg13g2_o21ai_1 _6336_ (.B1(net1927),
    .Y(_1892_),
    .A1(net1881),
    .A2(_1643_));
 sg13g2_nand3_1 _6337_ (.B(_1889_),
    .C(_1892_),
    .A(net1907),
    .Y(_1893_));
 sg13g2_nand4_1 _6338_ (.B(_1873_),
    .C(_1887_),
    .A(_1860_),
    .Y(_1894_),
    .D(_1893_));
 sg13g2_nor2_2 _6339_ (.A(net2081),
    .B(_1626_),
    .Y(_1895_));
 sg13g2_nor2_2 _6340_ (.A(net1837),
    .B(net1877),
    .Y(_1896_));
 sg13g2_nand2_2 _6341_ (.Y(_1897_),
    .A(net2237),
    .B(_1896_));
 sg13g2_nand2_1 _6342_ (.Y(_1898_),
    .A(_1895_),
    .B(_1897_));
 sg13g2_nor2_2 _6343_ (.A(net2108),
    .B(net1837),
    .Y(_1899_));
 sg13g2_a21oi_1 _6344_ (.A1(net1921),
    .A2(net1994),
    .Y(_1900_),
    .B1(net2212));
 sg13g2_o21ai_1 _6345_ (.B1(_1900_),
    .Y(_1901_),
    .A1(net1994),
    .A2(net1837));
 sg13g2_nand3_1 _6346_ (.B(_1898_),
    .C(_1901_),
    .A(net2196),
    .Y(_1902_));
 sg13g2_a21oi_2 _6347_ (.B1(_1899_),
    .Y(_1903_),
    .A2(_1642_),
    .A1(_1620_));
 sg13g2_nor2_1 _6348_ (.A(net2238),
    .B(_1903_),
    .Y(_1904_));
 sg13g2_o21ai_1 _6349_ (.B1(net2213),
    .Y(_1905_),
    .A1(net2238),
    .A2(_1903_));
 sg13g2_a21oi_1 _6350_ (.A1(_1554_),
    .A2(net1871),
    .Y(_1906_),
    .B1(_1863_));
 sg13g2_nand2_1 _6351_ (.Y(_1907_),
    .A(net2236),
    .B(net1827));
 sg13g2_a21oi_1 _6352_ (.A1(net2237),
    .A2(net1827),
    .Y(_1908_),
    .B1(net2210));
 sg13g2_nor2b_1 _6353_ (.A(_1906_),
    .B_N(_1908_),
    .Y(_1909_));
 sg13g2_nor2_1 _6354_ (.A(net2196),
    .B(_1909_),
    .Y(_1910_));
 sg13g2_o21ai_1 _6355_ (.B1(_1910_),
    .Y(_1911_),
    .A1(_1694_),
    .A2(_1905_));
 sg13g2_nand3_1 _6356_ (.B(_1902_),
    .C(_1911_),
    .A(net1772),
    .Y(_1912_));
 sg13g2_a21oi_1 _6357_ (.A1(_1894_),
    .A2(_1912_),
    .Y(_1913_),
    .B1(net1982));
 sg13g2_nand2_2 _6358_ (.Y(_1914_),
    .A(_1532_),
    .B(_1701_));
 sg13g2_a21oi_1 _6359_ (.A1(net1912),
    .A2(net1899),
    .Y(_1915_),
    .B1(net2193));
 sg13g2_a21oi_1 _6360_ (.A1(net1840),
    .A2(_1564_),
    .Y(_1916_),
    .B1(_1576_));
 sg13g2_or2_1 _6361_ (.X(_1917_),
    .B(_1916_),
    .A(_1914_));
 sg13g2_inv_1 _6362_ (.Y(_1918_),
    .A(_1917_));
 sg13g2_nand2_2 _6363_ (.Y(_1919_),
    .A(net2255),
    .B(net1898));
 sg13g2_o21ai_1 _6364_ (.B1(_1918_),
    .Y(_1920_),
    .A1(_1576_),
    .A2(_1919_));
 sg13g2_nor2_2 _6365_ (.A(net1913),
    .B(net2000),
    .Y(_1921_));
 sg13g2_nor2_1 _6366_ (.A(_1588_),
    .B(_1921_),
    .Y(_1922_));
 sg13g2_o21ai_1 _6367_ (.B1(net2189),
    .Y(_1923_),
    .A1(net2204),
    .A2(_1922_));
 sg13g2_nand2_1 _6368_ (.Y(_1924_),
    .A(_1569_),
    .B(_1923_));
 sg13g2_nand3_1 _6369_ (.B(_1850_),
    .C(net1852),
    .A(net1873),
    .Y(_1925_));
 sg13g2_o21ai_1 _6370_ (.B1(net2193),
    .Y(_1926_),
    .A1(net2214),
    .A2(net1876));
 sg13g2_nor2_2 _6371_ (.A(net2106),
    .B(net1897),
    .Y(_1927_));
 sg13g2_nor3_1 _6372_ (.A(net1918),
    .B(net2002),
    .C(_1927_),
    .Y(_1928_));
 sg13g2_nor2_1 _6373_ (.A(_1926_),
    .B(_1928_),
    .Y(_1929_));
 sg13g2_nand2_1 _6374_ (.Y(_1930_),
    .A(net2067),
    .B(net1839));
 sg13g2_nor2_1 _6375_ (.A(net2205),
    .B(net1916),
    .Y(_1931_));
 sg13g2_a21oi_1 _6376_ (.A1(_1930_),
    .A2(_1931_),
    .Y(_1932_),
    .B1(net2187));
 sg13g2_o21ai_1 _6377_ (.B1(_1932_),
    .Y(_1933_),
    .A1(net2080),
    .A2(net1878));
 sg13g2_a21oi_1 _6378_ (.A1(_1925_),
    .A2(_1929_),
    .Y(_1934_),
    .B1(net1935));
 sg13g2_a221oi_1 _6379_ (.B2(_1934_),
    .C1(_1920_),
    .B1(_1933_),
    .A1(net2093),
    .Y(_1935_),
    .A2(_1924_));
 sg13g2_nand2_2 _6380_ (.Y(_1936_),
    .A(_1533_),
    .B(_1662_));
 sg13g2_nand2_2 _6381_ (.Y(_1937_),
    .A(net2089),
    .B(net1984));
 sg13g2_nor2_2 _6382_ (.A(net1830),
    .B(_1676_),
    .Y(_1938_));
 sg13g2_nand2_2 _6383_ (.Y(_1939_),
    .A(_1642_),
    .B(net1821));
 sg13g2_nor2_1 _6384_ (.A(net2285),
    .B(net1828),
    .Y(_1940_));
 sg13g2_o21ai_1 _6385_ (.B1(net2238),
    .Y(_1941_),
    .A1(net2285),
    .A2(net1827));
 sg13g2_nand2_1 _6386_ (.Y(_1942_),
    .A(net2212),
    .B(_1941_));
 sg13g2_a221oi_1 _6387_ (.B2(net2072),
    .C1(_1942_),
    .B1(_1938_),
    .A1(net1879),
    .Y(_1943_),
    .A2(net1855));
 sg13g2_nor2_2 _6388_ (.A(net2076),
    .B(_1560_),
    .Y(_1944_));
 sg13g2_nand3_1 _6389_ (.B(net1879),
    .C(_1642_),
    .A(net2239),
    .Y(_1945_));
 sg13g2_nor2_2 _6390_ (.A(net2252),
    .B(_1896_),
    .Y(_1946_));
 sg13g2_nor2_1 _6391_ (.A(net2239),
    .B(_1946_),
    .Y(_1947_));
 sg13g2_o21ai_1 _6392_ (.B1(_1945_),
    .Y(_1948_),
    .A1(net2239),
    .A2(_1946_));
 sg13g2_nor2_2 _6393_ (.A(net2212),
    .B(_1947_),
    .Y(_1949_));
 sg13g2_a21oi_1 _6394_ (.A1(_1945_),
    .A2(_1949_),
    .Y(_1950_),
    .B1(_1943_));
 sg13g2_o21ai_1 _6395_ (.B1(_1777_),
    .Y(_1951_),
    .A1(net1892),
    .A2(_1619_));
 sg13g2_nand3_1 _6396_ (.B(net2007),
    .C(_1666_),
    .A(net2237),
    .Y(_1952_));
 sg13g2_nor2_1 _6397_ (.A(net1923),
    .B(_1552_),
    .Y(_1953_));
 sg13g2_a21oi_1 _6398_ (.A1(_1952_),
    .A2(_1953_),
    .Y(_1954_),
    .B1(net1935));
 sg13g2_o21ai_1 _6399_ (.B1(_1954_),
    .Y(_1955_),
    .A1(net1931),
    .A2(_1951_));
 sg13g2_o21ai_1 _6400_ (.B1(_1955_),
    .Y(_1956_),
    .A1(_1937_),
    .A2(_1950_));
 sg13g2_nand2_1 _6401_ (.Y(_1957_),
    .A(_1895_),
    .B(_1945_));
 sg13g2_nor2_2 _6402_ (.A(net2208),
    .B(_1822_),
    .Y(_1958_));
 sg13g2_o21ai_1 _6403_ (.B1(_1958_),
    .Y(_1959_),
    .A1(net2238),
    .A2(_1682_));
 sg13g2_nand3_1 _6404_ (.B(_1957_),
    .C(_1959_),
    .A(net2197),
    .Y(_1960_));
 sg13g2_nor2_2 _6405_ (.A(net2091),
    .B(_1558_),
    .Y(_1961_));
 sg13g2_nor2_2 _6406_ (.A(_4042_),
    .B(_1558_),
    .Y(_1962_));
 sg13g2_nand2_1 _6407_ (.Y(_1963_),
    .A(net2186),
    .B(net1840));
 sg13g2_nor2_2 _6408_ (.A(_1558_),
    .B(_1576_),
    .Y(_1964_));
 sg13g2_nand2_2 _6409_ (.Y(_1965_),
    .A(net1880),
    .B(_1746_));
 sg13g2_nand2_2 _6410_ (.Y(_1966_),
    .A(_1620_),
    .B(_1865_));
 sg13g2_a21oi_1 _6411_ (.A1(_1965_),
    .A2(_1966_),
    .Y(_1967_),
    .B1(_1879_));
 sg13g2_nor2_2 _6412_ (.A(net2206),
    .B(net1834),
    .Y(_1968_));
 sg13g2_nor2_1 _6413_ (.A(net2212),
    .B(_1940_),
    .Y(_1969_));
 sg13g2_nor2_1 _6414_ (.A(_1550_),
    .B(net1830),
    .Y(_1970_));
 sg13g2_nor2_1 _6415_ (.A(net2082),
    .B(_1945_),
    .Y(_1971_));
 sg13g2_nor4_1 _6416_ (.A(net1864),
    .B(_1967_),
    .C(_1969_),
    .D(_1971_),
    .Y(_1972_));
 sg13g2_a221oi_1 _6417_ (.B2(_1888_),
    .C1(_1972_),
    .B1(_1964_),
    .A1(_1956_),
    .Y(_1973_),
    .A2(_1960_));
 sg13g2_nor2_1 _6418_ (.A(_1936_),
    .B(_1973_),
    .Y(_1974_));
 sg13g2_a21oi_1 _6419_ (.A1(_1867_),
    .A2(_1961_),
    .Y(_1975_),
    .B1(net1939));
 sg13g2_nor2_1 _6420_ (.A(net1988),
    .B(_1874_),
    .Y(_1976_));
 sg13g2_nor2_2 _6421_ (.A(net1882),
    .B(_1810_),
    .Y(_1977_));
 sg13g2_o21ai_1 _6422_ (.B1(net2234),
    .Y(_1978_),
    .A1(_1870_),
    .A2(_1977_));
 sg13g2_a221oi_1 _6423_ (.B2(_1978_),
    .C1(net2186),
    .B1(_1976_),
    .A1(net1988),
    .Y(_1979_),
    .A2(net1858));
 sg13g2_nor3_1 _6424_ (.A(_1861_),
    .B(_1975_),
    .C(_1979_),
    .Y(_1980_));
 sg13g2_nor2_2 _6425_ (.A(_1535_),
    .B(_1859_),
    .Y(_1981_));
 sg13g2_nand2_2 _6426_ (.Y(_1982_),
    .A(_1577_),
    .B(net1880));
 sg13g2_nand2_2 _6427_ (.Y(_1983_),
    .A(net1900),
    .B(_1809_));
 sg13g2_a221oi_1 _6428_ (.B2(net2005),
    .C1(_1550_),
    .B1(_1746_),
    .A1(_1681_),
    .Y(_1984_),
    .A2(_1685_));
 sg13g2_a21oi_1 _6429_ (.A1(net2009),
    .A2(net1834),
    .Y(_1985_),
    .B1(net2206));
 sg13g2_inv_1 _6430_ (.Y(_1986_),
    .A(_1985_));
 sg13g2_o21ai_1 _6431_ (.B1(_1985_),
    .Y(_1987_),
    .A1(net1834),
    .A2(net1820));
 sg13g2_nand3_1 _6432_ (.B(_1812_),
    .C(net1853),
    .A(_1691_),
    .Y(_1988_));
 sg13g2_nand2_1 _6433_ (.Y(_1989_),
    .A(_1987_),
    .B(_1988_));
 sg13g2_o21ai_1 _6434_ (.B1(_1761_),
    .Y(_1990_),
    .A1(_1984_),
    .A2(_1989_));
 sg13g2_nand3_1 _6435_ (.B(_1705_),
    .C(_1849_),
    .A(net1920),
    .Y(_1991_));
 sg13g2_nand2_2 _6436_ (.Y(_1992_),
    .A(net2087),
    .B(net1862));
 sg13g2_inv_2 _6437_ (.Y(_1993_),
    .A(_1992_));
 sg13g2_nand2_1 _6438_ (.Y(_1994_),
    .A(_1991_),
    .B(_1993_));
 sg13g2_nor2_1 _6439_ (.A(_1806_),
    .B(_1994_),
    .Y(_1995_));
 sg13g2_nor3_1 _6440_ (.A(_1457_),
    .B(net2006),
    .C(net1878),
    .Y(_1996_));
 sg13g2_nand2_2 _6441_ (.Y(_1997_),
    .A(net1875),
    .B(_1768_));
 sg13g2_nand2_2 _6442_ (.Y(_1998_),
    .A(net2256),
    .B(_1997_));
 sg13g2_nand2_2 _6443_ (.Y(_1999_),
    .A(net2105),
    .B(net1911));
 sg13g2_a21oi_2 _6444_ (.B1(net2069),
    .Y(_2000_),
    .A2(net1911),
    .A1(net2106));
 sg13g2_a21oi_2 _6445_ (.B1(net2227),
    .Y(_2001_),
    .A2(net1911),
    .A1(net2259));
 sg13g2_nand2_1 _6446_ (.Y(_2002_),
    .A(_1667_),
    .B(net1859));
 sg13g2_a221oi_1 _6447_ (.B2(_2002_),
    .C1(net1942),
    .B1(_2001_),
    .A1(_1998_),
    .Y(_2003_),
    .A2(_2000_));
 sg13g2_a21oi_2 _6448_ (.B1(net1986),
    .Y(_2004_),
    .A2(_1996_),
    .A1(net2012));
 sg13g2_nor2_1 _6449_ (.A(net1934),
    .B(_2004_),
    .Y(_2005_));
 sg13g2_nand2b_1 _6450_ (.Y(_2006_),
    .B(net1937),
    .A_N(_2004_));
 sg13g2_nor2_1 _6451_ (.A(net2209),
    .B(net1869),
    .Y(_2007_));
 sg13g2_nand2_1 _6452_ (.Y(_2008_),
    .A(net2090),
    .B(net2004));
 sg13g2_o21ai_1 _6453_ (.B1(_2005_),
    .Y(_2009_),
    .A1(_2007_),
    .A2(_2008_));
 sg13g2_o21ai_1 _6454_ (.B1(_1990_),
    .Y(_2010_),
    .A1(_2003_),
    .A2(_2009_));
 sg13g2_o21ai_1 _6455_ (.B1(_1981_),
    .Y(_2011_),
    .A1(_1995_),
    .A2(_2010_));
 sg13g2_a21oi_1 _6456_ (.A1(net2292),
    .A2(net2295),
    .Y(_2012_),
    .B1(_1647_));
 sg13g2_nor2_1 _6457_ (.A(net2243),
    .B(net1881),
    .Y(_2013_));
 sg13g2_nand2b_1 _6458_ (.Y(_2014_),
    .B(_2013_),
    .A_N(_1775_));
 sg13g2_o21ai_1 _6459_ (.B1(_2014_),
    .Y(_2015_),
    .A1(_1714_),
    .A2(_2012_));
 sg13g2_nor2_1 _6460_ (.A(net2216),
    .B(_2015_),
    .Y(_2016_));
 sg13g2_nor2_2 _6461_ (.A(_1682_),
    .B(_1740_),
    .Y(_2017_));
 sg13g2_nand2_2 _6462_ (.Y(_2018_),
    .A(_1681_),
    .B(_1741_));
 sg13g2_a21oi_1 _6463_ (.A1(net2109),
    .A2(_2018_),
    .Y(_2019_),
    .B1(_1550_));
 sg13g2_nand2_1 _6464_ (.Y(_2020_),
    .A(_1749_),
    .B(_2019_));
 sg13g2_o21ai_1 _6465_ (.B1(_2020_),
    .Y(_2021_),
    .A1(net1851),
    .A2(_2018_));
 sg13g2_o21ai_1 _6466_ (.B1(_1702_),
    .Y(_2022_),
    .A1(_2016_),
    .A2(_2021_));
 sg13g2_nand4_1 _6467_ (.B(_1781_),
    .C(_1828_),
    .A(net1757),
    .Y(_2023_),
    .D(_2011_));
 sg13g2_nor3_1 _6468_ (.A(_1843_),
    .B(_1980_),
    .C(_2023_),
    .Y(_2024_));
 sg13g2_nand4_1 _6469_ (.B(_1847_),
    .C(_1851_),
    .A(_1663_),
    .Y(_2025_),
    .D(_1855_));
 sg13g2_a21oi_1 _6470_ (.A1(_2022_),
    .A2(_2025_),
    .Y(_2026_),
    .B1(_1857_));
 sg13g2_nor4_1 _6471_ (.A(_1913_),
    .B(_1935_),
    .C(_1974_),
    .D(_2026_),
    .Y(_2027_));
 sg13g2_nand3_1 _6472_ (.B(_2024_),
    .C(_2027_),
    .A(_1732_),
    .Y(_2028_));
 sg13g2_o21ai_1 _6473_ (.B1(_2028_),
    .Y(_2029_),
    .A1(net1757),
    .A2(_1598_));
 sg13g2_nand3b_1 _6474_ (.B(_2029_),
    .C(\draw_game_inst.board_x[0] ),
    .Y(_2030_),
    .A_N(\draw_game_inst.board_x[1] ));
 sg13g2_nor2_2 _6475_ (.A(net2264),
    .B(_1457_),
    .Y(_2031_));
 sg13g2_nor2_2 _6476_ (.A(net2285),
    .B(_1460_),
    .Y(_2032_));
 sg13g2_nand2_1 _6477_ (.Y(_2033_),
    .A(_4055_),
    .B(net2017));
 sg13g2_nand2_2 _6478_ (.Y(_2034_),
    .A(net2256),
    .B(net1850));
 sg13g2_nor2_1 _6479_ (.A(net2070),
    .B(_2031_),
    .Y(_2035_));
 sg13g2_nand2_2 _6480_ (.Y(_2036_),
    .A(net2287),
    .B(net2295));
 sg13g2_nand2_2 _6481_ (.Y(_2037_),
    .A(_1787_),
    .B(_2036_));
 sg13g2_nand2_1 _6482_ (.Y(_2038_),
    .A(net2105),
    .B(_2037_));
 sg13g2_a21oi_1 _6483_ (.A1(net2257),
    .A2(_1458_),
    .Y(_2039_),
    .B1(net2230));
 sg13g2_a221oi_1 _6484_ (.B2(_2039_),
    .C1(net2080),
    .B1(_2038_),
    .A1(_2034_),
    .Y(_2040_),
    .A2(_2035_));
 sg13g2_nand2_2 _6485_ (.Y(_2041_),
    .A(net2065),
    .B(net2004));
 sg13g2_nand2_1 _6486_ (.Y(_2042_),
    .A(_4055_),
    .B(_1620_));
 sg13g2_a22oi_1 _6487_ (.Y(_2043_),
    .B1(_1813_),
    .B2(_2041_),
    .A2(_1620_),
    .A1(_4055_));
 sg13g2_a221oi_1 _6488_ (.B2(net1997),
    .C1(_2040_),
    .B1(_2043_),
    .A1(net1868),
    .Y(_2044_),
    .A2(_2037_));
 sg13g2_nor2_1 _6489_ (.A(net2284),
    .B(net1871),
    .Y(_2045_));
 sg13g2_nor2_2 _6490_ (.A(net2285),
    .B(net1825),
    .Y(_2046_));
 sg13g2_inv_1 _6491_ (.Y(_2047_),
    .A(_2046_));
 sg13g2_o21ai_1 _6492_ (.B1(_2001_),
    .Y(_2048_),
    .A1(net2259),
    .A2(_2046_));
 sg13g2_a22oi_1 _6493_ (.Y(_2049_),
    .B1(net1825),
    .B2(net2104),
    .A2(_1639_),
    .A1(net1911));
 sg13g2_nand2_1 _6494_ (.Y(_2050_),
    .A(net2227),
    .B(_2049_));
 sg13g2_nand3_1 _6495_ (.B(_2048_),
    .C(_2050_),
    .A(net1948),
    .Y(_2051_));
 sg13g2_o21ai_1 _6496_ (.B1(_2051_),
    .Y(_2052_),
    .A1(net2191),
    .A2(_2044_));
 sg13g2_nor2_1 _6497_ (.A(_2006_),
    .B(_2052_),
    .Y(_2053_));
 sg13g2_nand3_1 _6498_ (.B(net1861),
    .C(_1805_),
    .A(_1706_),
    .Y(_2054_));
 sg13g2_nor2_1 _6499_ (.A(net2222),
    .B(net1850),
    .Y(_2055_));
 sg13g2_nand2_2 _6500_ (.Y(_2056_),
    .A(net1949),
    .B(net1859));
 sg13g2_a21oi_1 _6501_ (.A1(net1993),
    .A2(_2032_),
    .Y(_2057_),
    .B1(_2056_));
 sg13g2_a21oi_1 _6502_ (.A1(_1883_),
    .A2(_1982_),
    .Y(_2058_),
    .B1(_2057_));
 sg13g2_nor2_1 _6503_ (.A(net2255),
    .B(net1813),
    .Y(_2059_));
 sg13g2_nand2_1 _6504_ (.Y(_2060_),
    .A(_1648_),
    .B(_1982_));
 sg13g2_nor2b_1 _6505_ (.A(_2059_),
    .B_N(_2060_),
    .Y(_2061_));
 sg13g2_o21ai_1 _6506_ (.B1(_2058_),
    .Y(_2062_),
    .A1(_1880_),
    .A2(_2061_));
 sg13g2_a21oi_1 _6507_ (.A1(net1863),
    .A2(_2054_),
    .Y(_2063_),
    .B1(_2062_));
 sg13g2_o21ai_1 _6508_ (.B1(_1981_),
    .Y(_2064_),
    .A1(_2053_),
    .A2(_2063_));
 sg13g2_nand2_1 _6509_ (.Y(_2065_),
    .A(net2180),
    .B(_1731_));
 sg13g2_nand2_1 _6510_ (.Y(_2066_),
    .A(_1615_),
    .B(_2065_));
 sg13g2_nand3_1 _6511_ (.B(_1654_),
    .C(_1897_),
    .A(_1627_),
    .Y(_2067_));
 sg13g2_nor2_1 _6512_ (.A(net2104),
    .B(net2227),
    .Y(_2068_));
 sg13g2_nand2_2 _6513_ (.Y(_2069_),
    .A(net2264),
    .B(net2074));
 sg13g2_nor2_1 _6514_ (.A(net1899),
    .B(_2069_),
    .Y(_2070_));
 sg13g2_a221oi_1 _6515_ (.B2(net2214),
    .C1(net2193),
    .B1(_2070_),
    .A1(net1910),
    .Y(_2071_),
    .A2(_1853_));
 sg13g2_o21ai_1 _6516_ (.B1(net1950),
    .Y(_2072_),
    .A1(net1892),
    .A2(net1819));
 sg13g2_o21ai_1 _6517_ (.B1(net2208),
    .Y(_2073_),
    .A1(net1924),
    .A2(net1897));
 sg13g2_o21ai_1 _6518_ (.B1(net1887),
    .Y(_2074_),
    .A1(net1926),
    .A2(net1899));
 sg13g2_nand2b_1 _6519_ (.Y(_2075_),
    .B(_1652_),
    .A_N(_2074_));
 sg13g2_o21ai_1 _6520_ (.B1(_2075_),
    .Y(_2076_),
    .A1(_1588_),
    .A2(_2072_));
 sg13g2_a21oi_1 _6521_ (.A1(_2067_),
    .A2(_2071_),
    .Y(_2077_),
    .B1(_2076_));
 sg13g2_a21oi_1 _6522_ (.A1(_1868_),
    .A2(_1907_),
    .Y(_2078_),
    .B1(net1931));
 sg13g2_a21oi_1 _6523_ (.A1(_1619_),
    .A2(_1844_),
    .Y(_2079_),
    .B1(net2001));
 sg13g2_nor2_1 _6524_ (.A(net2000),
    .B(_1626_),
    .Y(_2080_));
 sg13g2_nor3_2 _6525_ (.A(net2208),
    .B(net1912),
    .C(_1816_),
    .Y(_2081_));
 sg13g2_nand2b_1 _6526_ (.Y(_2082_),
    .B(net2195),
    .A_N(_2081_));
 sg13g2_a21oi_1 _6527_ (.A1(_1895_),
    .A2(_2079_),
    .Y(_2083_),
    .B1(_2082_));
 sg13g2_a21oi_1 _6528_ (.A1(_1817_),
    .A2(_1939_),
    .Y(_2084_),
    .B1(net1904));
 sg13g2_or4_1 _6529_ (.A(net2183),
    .B(_2078_),
    .C(_2083_),
    .D(_2084_),
    .X(_2085_));
 sg13g2_a21oi_1 _6530_ (.A1(net2093),
    .A2(_2085_),
    .Y(_2086_),
    .B1(_2066_));
 sg13g2_o21ai_1 _6531_ (.B1(_2086_),
    .Y(_2087_),
    .A1(net1935),
    .A2(_2077_));
 sg13g2_nand2_1 _6532_ (.Y(_2088_),
    .A(_1577_),
    .B(_2000_));
 sg13g2_nand3_1 _6533_ (.B(_1548_),
    .C(_2088_),
    .A(net2205),
    .Y(_2089_));
 sg13g2_nand2_1 _6534_ (.Y(_2090_),
    .A(_1932_),
    .B(_2089_));
 sg13g2_nand3_1 _6535_ (.B(_1443_),
    .C(net2004),
    .A(net2079),
    .Y(_2091_));
 sg13g2_a221oi_1 _6536_ (.B2(net2206),
    .C1(net2085),
    .B1(net1913),
    .A1(net2222),
    .Y(_2092_),
    .A2(net1920));
 sg13g2_nand2_1 _6537_ (.Y(_2093_),
    .A(_2091_),
    .B(_2092_));
 sg13g2_nand3_1 _6538_ (.B(_2090_),
    .C(_2093_),
    .A(net1938),
    .Y(_2094_));
 sg13g2_a21oi_1 _6539_ (.A1(net2208),
    .A2(net1839),
    .Y(_2095_),
    .B1(_1832_));
 sg13g2_o21ai_1 _6540_ (.B1(net2092),
    .Y(_2096_),
    .A1(_1566_),
    .A2(_2095_));
 sg13g2_nand3_1 _6541_ (.B(_2094_),
    .C(_2096_),
    .A(_1831_),
    .Y(_2097_));
 sg13g2_nand2_1 _6542_ (.Y(_2098_),
    .A(net2261),
    .B(_1866_));
 sg13g2_nand3_1 _6543_ (.B(_1966_),
    .C(_2098_),
    .A(net1840),
    .Y(_2099_));
 sg13g2_a21oi_1 _6544_ (.A1(_1575_),
    .A2(_2099_),
    .Y(_2100_),
    .B1(_1861_));
 sg13g2_nand2_1 _6545_ (.Y(_2101_),
    .A(net1994),
    .B(_1897_));
 sg13g2_o21ai_1 _6546_ (.B1(_2101_),
    .Y(_2102_),
    .A1(net1827),
    .A2(_1748_));
 sg13g2_nand2b_1 _6547_ (.Y(_2103_),
    .B(_2102_),
    .A_N(_1874_));
 sg13g2_nor2_2 _6548_ (.A(net2227),
    .B(_1437_),
    .Y(_2104_));
 sg13g2_nand2b_2 _6549_ (.Y(_2105_),
    .B(net1858),
    .A_N(_2104_));
 sg13g2_nand2_1 _6550_ (.Y(_2106_),
    .A(net2212),
    .B(_1436_));
 sg13g2_a21oi_1 _6551_ (.A1(_1785_),
    .A2(_2106_),
    .Y(_2107_),
    .B1(net2197));
 sg13g2_a221oi_1 _6552_ (.B2(net1950),
    .C1(_2107_),
    .B1(_2105_),
    .A1(net1887),
    .Y(_2108_),
    .A2(_2103_));
 sg13g2_nor2_2 _6553_ (.A(net2030),
    .B(net1828),
    .Y(_2109_));
 sg13g2_nand2_2 _6554_ (.Y(_2110_),
    .A(_1435_),
    .B(net1826));
 sg13g2_nand2_1 _6555_ (.Y(_2111_),
    .A(net1865),
    .B(_2110_));
 sg13g2_nand2_1 _6556_ (.Y(_2112_),
    .A(_1666_),
    .B(_1888_));
 sg13g2_nor2_2 _6557_ (.A(net2288),
    .B(net1828),
    .Y(_2113_));
 sg13g2_nand2_2 _6558_ (.Y(_2114_),
    .A(net2064),
    .B(net1826));
 sg13g2_a22oi_1 _6559_ (.Y(_2115_),
    .B1(_1648_),
    .B2(_2114_),
    .A2(_1642_),
    .A1(_1620_));
 sg13g2_o21ai_1 _6560_ (.B1(_1869_),
    .Y(_2116_),
    .A1(net2002),
    .A2(_2115_));
 sg13g2_a221oi_1 _6561_ (.B2(net1852),
    .C1(_2116_),
    .B1(_2112_),
    .A1(net1866),
    .Y(_2117_),
    .A2(_2110_));
 sg13g2_nand2_2 _6562_ (.Y(_2118_),
    .A(net1950),
    .B(net1823));
 sg13g2_nor2_2 _6563_ (.A(net2106),
    .B(net1916),
    .Y(_2119_));
 sg13g2_a221oi_1 _6564_ (.B2(net1873),
    .C1(net2234),
    .B1(_2119_),
    .A1(net2110),
    .Y(_2120_),
    .A2(_1644_));
 sg13g2_nand2_1 _6565_ (.Y(_2121_),
    .A(net1874),
    .B(_1667_));
 sg13g2_a22oi_1 _6566_ (.Y(_2122_),
    .B1(_1882_),
    .B2(net2263),
    .A2(_1667_),
    .A1(net1873));
 sg13g2_nor2_1 _6567_ (.A(_1880_),
    .B(_2122_),
    .Y(_2123_));
 sg13g2_nor3_1 _6568_ (.A(net2183),
    .B(_1886_),
    .C(_2123_),
    .Y(_2124_));
 sg13g2_o21ai_1 _6569_ (.B1(_2124_),
    .Y(_2125_),
    .A1(_2118_),
    .A2(_2120_));
 sg13g2_inv_1 _6570_ (.Y(_2126_),
    .A(_2125_));
 sg13g2_o21ai_1 _6571_ (.B1(_2126_),
    .Y(_2127_),
    .A1(net2195),
    .A2(_2117_));
 sg13g2_a221oi_1 _6572_ (.B2(net2092),
    .C1(_1861_),
    .B1(_2127_),
    .A1(_1575_),
    .Y(_2128_),
    .A2(_2099_));
 sg13g2_o21ai_1 _6573_ (.B1(_2128_),
    .Y(_2129_),
    .A1(net1935),
    .A2(_2108_));
 sg13g2_nor2_1 _6574_ (.A(net2257),
    .B(net1831),
    .Y(_2130_));
 sg13g2_nor2_2 _6575_ (.A(net2262),
    .B(_1939_),
    .Y(_2131_));
 sg13g2_o21ai_1 _6576_ (.B1(net1998),
    .Y(_2132_),
    .A1(_1899_),
    .A2(_2131_));
 sg13g2_a21oi_2 _6577_ (.B1(net2003),
    .Y(_2133_),
    .A2(_2060_),
    .A1(_1983_));
 sg13g2_nor2_2 _6578_ (.A(_1562_),
    .B(net1851),
    .Y(_2134_));
 sg13g2_nor2_2 _6579_ (.A(net2234),
    .B(net1838),
    .Y(_2135_));
 sg13g2_nand2_2 _6580_ (.Y(_2136_),
    .A(net2068),
    .B(net1897));
 sg13g2_a221oi_1 _6581_ (.B2(net1921),
    .C1(_2133_),
    .B1(_2134_),
    .A1(net1866),
    .Y(_2137_),
    .A2(net1814));
 sg13g2_a21oi_1 _6582_ (.A1(_2132_),
    .A2(_2137_),
    .Y(_2138_),
    .B1(net2197));
 sg13g2_o21ai_1 _6583_ (.B1(_1590_),
    .Y(_2139_),
    .A1(_1681_),
    .A2(_1820_));
 sg13g2_nor2_2 _6584_ (.A(net1994),
    .B(_1888_),
    .Y(_2140_));
 sg13g2_a21oi_1 _6585_ (.A1(net1855),
    .A2(_1938_),
    .Y(_2141_),
    .B1(_2140_));
 sg13g2_o21ai_1 _6586_ (.B1(_2139_),
    .Y(_2142_),
    .A1(net1989),
    .A2(_2141_));
 sg13g2_nor2_2 _6587_ (.A(net2110),
    .B(net1830),
    .Y(_2143_));
 sg13g2_a22oi_1 _6588_ (.Y(_2144_),
    .B1(net1821),
    .B2(_2143_),
    .A2(net1835),
    .A1(net2110));
 sg13g2_o21ai_1 _6589_ (.B1(net1940),
    .Y(_2145_),
    .A1(_1880_),
    .A2(_2144_));
 sg13g2_nor3_1 _6590_ (.A(_2138_),
    .B(_2142_),
    .C(_2145_),
    .Y(_2146_));
 sg13g2_nand2_1 _6591_ (.Y(_2147_),
    .A(net2254),
    .B(net1819));
 sg13g2_nor2_2 _6592_ (.A(_1683_),
    .B(_1919_),
    .Y(_2148_));
 sg13g2_nor2_1 _6593_ (.A(net2262),
    .B(_1679_),
    .Y(_2149_));
 sg13g2_o21ai_1 _6594_ (.B1(net2071),
    .Y(_2150_),
    .A1(_2148_),
    .A2(_2149_));
 sg13g2_nand2_1 _6595_ (.Y(_2151_),
    .A(_1941_),
    .B(_2150_));
 sg13g2_nor2_2 _6596_ (.A(net1994),
    .B(_1939_),
    .Y(_2152_));
 sg13g2_a221oi_1 _6597_ (.B2(_2013_),
    .C1(_2152_),
    .B1(_1865_),
    .A1(net1828),
    .Y(_2153_),
    .A2(net1855));
 sg13g2_nand2_1 _6598_ (.Y(_2154_),
    .A(net1896),
    .B(net1814));
 sg13g2_o21ai_1 _6599_ (.B1(_2154_),
    .Y(_2155_),
    .A1(net1896),
    .A2(_1939_));
 sg13g2_a21oi_1 _6600_ (.A1(net1907),
    .A2(_2155_),
    .Y(_2156_),
    .B1(net1982));
 sg13g2_o21ai_1 _6601_ (.B1(_2156_),
    .Y(_2157_),
    .A1(net1989),
    .A2(_2153_));
 sg13g2_a221oi_1 _6602_ (.B2(net1950),
    .C1(_2157_),
    .B1(_2151_),
    .A1(net2015),
    .Y(_2158_),
    .A2(_1948_));
 sg13g2_o21ai_1 _6603_ (.B1(_1557_),
    .Y(_2159_),
    .A1(net1876),
    .A2(_1903_));
 sg13g2_o21ai_1 _6604_ (.B1(_1964_),
    .Y(_2160_),
    .A1(net1877),
    .A2(_1903_));
 sg13g2_nand2b_1 _6605_ (.Y(_2161_),
    .B(_2160_),
    .A_N(_2146_));
 sg13g2_nor2_1 _6606_ (.A(_2158_),
    .B(_2161_),
    .Y(_2162_));
 sg13g2_o21ai_1 _6607_ (.B1(_2129_),
    .Y(_2163_),
    .A1(_1936_),
    .A2(_2162_));
 sg13g2_nor2_2 _6608_ (.A(net2210),
    .B(net2001),
    .Y(_2164_));
 sg13g2_nor2_2 _6609_ (.A(net2260),
    .B(net1851),
    .Y(_2165_));
 sg13g2_o21ai_1 _6610_ (.B1(_1915_),
    .Y(_2166_),
    .A1(_2164_),
    .A2(_2165_));
 sg13g2_inv_1 _6611_ (.Y(_2167_),
    .A(_2166_));
 sg13g2_nand3_1 _6612_ (.B(_1564_),
    .C(_1571_),
    .A(net2193),
    .Y(_2168_));
 sg13g2_a21oi_1 _6613_ (.A1(_2166_),
    .A2(_2168_),
    .Y(_2169_),
    .B1(net2183));
 sg13g2_a21oi_1 _6614_ (.A1(net1912),
    .A2(net1898),
    .Y(_2170_),
    .B1(_0093_));
 sg13g2_a21oi_1 _6615_ (.A1(_1668_),
    .A2(_2170_),
    .Y(_2171_),
    .B1(net1988));
 sg13g2_nand2b_2 _6616_ (.Y(_2172_),
    .B(net2214),
    .A_N(_0093_));
 sg13g2_o21ai_1 _6617_ (.B1(_1926_),
    .Y(_2173_),
    .A1(net1873),
    .A2(_2172_));
 sg13g2_a21oi_1 _6618_ (.A1(_1654_),
    .A2(_1915_),
    .Y(_2174_),
    .B1(_2173_));
 sg13g2_o21ai_1 _6619_ (.B1(net1939),
    .Y(_2175_),
    .A1(_2171_),
    .A2(_2174_));
 sg13g2_o21ai_1 _6620_ (.B1(_2175_),
    .Y(_2176_),
    .A1(net2180),
    .A2(_2169_));
 sg13g2_nor2_1 _6621_ (.A(_1917_),
    .B(_2176_),
    .Y(_2177_));
 sg13g2_nor2b_1 _6622_ (.A(net2288),
    .B_N(_0096_),
    .Y(_2178_));
 sg13g2_nand2_2 _6623_ (.Y(_2179_),
    .A(net2063),
    .B(_0096_));
 sg13g2_nor2_1 _6624_ (.A(net2266),
    .B(_2178_),
    .Y(_2180_));
 sg13g2_a221oi_1 _6625_ (.B2(_1677_),
    .C1(net2075),
    .B1(_2180_),
    .A1(net2266),
    .Y(_2181_),
    .A2(_1938_));
 sg13g2_nand3_1 _6626_ (.B(net1901),
    .C(_2036_),
    .A(_1435_),
    .Y(_2182_));
 sg13g2_a221oi_1 _6627_ (.B2(_2182_),
    .C1(_2181_),
    .B1(net1849),
    .A1(net2010),
    .Y(_2183_),
    .A2(net1850));
 sg13g2_nand2_1 _6628_ (.Y(_2184_),
    .A(_1691_),
    .B(_2036_));
 sg13g2_nand2_1 _6629_ (.Y(_2185_),
    .A(net2241),
    .B(_2184_));
 sg13g2_inv_1 _6630_ (.Y(_2186_),
    .A(_2185_));
 sg13g2_o21ai_1 _6631_ (.B1(_2185_),
    .Y(_2187_),
    .A1(_1719_),
    .A2(_2069_));
 sg13g2_nand2b_1 _6632_ (.Y(_2188_),
    .B(_1889_),
    .A_N(_2187_));
 sg13g2_a21oi_1 _6633_ (.A1(net2215),
    .A2(_2188_),
    .Y(_2189_),
    .B1(_1857_));
 sg13g2_o21ai_1 _6634_ (.B1(_2189_),
    .Y(_2190_),
    .A1(net2215),
    .A2(_2183_));
 sg13g2_nor2_2 _6635_ (.A(net2104),
    .B(net2017),
    .Y(_2191_));
 sg13g2_nor2_2 _6636_ (.A(net2258),
    .B(_1692_),
    .Y(_2192_));
 sg13g2_o21ai_1 _6637_ (.B1(net2229),
    .Y(_2193_),
    .A1(_2191_),
    .A2(_2192_));
 sg13g2_nor2_2 _6638_ (.A(net2068),
    .B(net1929),
    .Y(_2194_));
 sg13g2_nand2_2 _6639_ (.Y(_2195_),
    .A(net2228),
    .B(net2014));
 sg13g2_nand3_1 _6640_ (.B(net1911),
    .C(_1691_),
    .A(net2014),
    .Y(_2196_));
 sg13g2_nand2_1 _6641_ (.Y(_2197_),
    .A(_2195_),
    .B(_2196_));
 sg13g2_nand2_1 _6642_ (.Y(_2198_),
    .A(_1684_),
    .B(_2179_));
 sg13g2_nand2_1 _6643_ (.Y(_2199_),
    .A(_1996_),
    .B(net1848));
 sg13g2_a221oi_1 _6644_ (.B2(net2008),
    .C1(net1943),
    .B1(_2198_),
    .A1(net2230),
    .Y(_2200_),
    .A2(_2042_));
 sg13g2_o21ai_1 _6645_ (.B1(net1906),
    .Y(_2201_),
    .A1(net2229),
    .A2(_1692_));
 sg13g2_a221oi_1 _6646_ (.B2(net1890),
    .C1(_2201_),
    .B1(_2198_),
    .A1(_1460_),
    .Y(_2202_),
    .A2(net1857));
 sg13g2_a221oi_1 _6647_ (.B2(_2200_),
    .C1(_2202_),
    .B1(_2199_),
    .A1(_2193_),
    .Y(_2203_),
    .A2(_2197_));
 sg13g2_o21ai_1 _6648_ (.B1(_2190_),
    .Y(_2204_),
    .A1(net1936),
    .A2(_2203_));
 sg13g2_a21o_1 _6649_ (.A2(_2204_),
    .A1(net1771),
    .B1(_2177_),
    .X(_2205_));
 sg13g2_a21oi_1 _6650_ (.A1(net2070),
    .A2(net1859),
    .Y(_2206_),
    .B1(net2209));
 sg13g2_nor2_2 _6651_ (.A(net2253),
    .B(net1859),
    .Y(_2207_));
 sg13g2_nand2_1 _6652_ (.Y(_2208_),
    .A(net1992),
    .B(_1805_));
 sg13g2_or2_1 _6653_ (.X(_2209_),
    .B(_0095_),
    .A(net2293));
 sg13g2_o21ai_1 _6654_ (.B1(_2209_),
    .Y(_2210_),
    .A1(net2062),
    .A2(net2285));
 sg13g2_a22oi_1 _6655_ (.Y(_2211_),
    .B1(_2210_),
    .B2(net2257),
    .A2(_1805_),
    .A1(net1992));
 sg13g2_inv_1 _6656_ (.Y(_2212_),
    .A(_2211_));
 sg13g2_a22oi_1 _6657_ (.Y(_2213_),
    .B1(_2212_),
    .B2(_2206_),
    .A2(_2210_),
    .A1(_2165_));
 sg13g2_o21ai_1 _6658_ (.B1(net2231),
    .Y(_2214_),
    .A1(net2251),
    .A2(net1835));
 sg13g2_o21ai_1 _6659_ (.B1(_1804_),
    .Y(_2215_),
    .A1(net2257),
    .A2(net1835));
 sg13g2_a221oi_1 _6660_ (.B2(_1895_),
    .C1(net2191),
    .B1(_2215_),
    .A1(_2206_),
    .Y(_2216_),
    .A2(_2214_));
 sg13g2_a21oi_1 _6661_ (.A1(net2191),
    .A2(_2213_),
    .Y(_2217_),
    .B1(net1934));
 sg13g2_nand2b_1 _6662_ (.Y(_2218_),
    .B(_2217_),
    .A_N(_2216_));
 sg13g2_nor3_1 _6663_ (.A(net2258),
    .B(_1790_),
    .C(_1802_),
    .Y(_2219_));
 sg13g2_o21ai_1 _6664_ (.B1(_2208_),
    .Y(_2220_),
    .A1(_1715_),
    .A2(_1787_));
 sg13g2_a21oi_1 _6665_ (.A1(net1821),
    .A2(_1716_),
    .Y(_2221_),
    .B1(net2204));
 sg13g2_a21oi_1 _6666_ (.A1(_2220_),
    .A2(_2221_),
    .Y(_2222_),
    .B1(net2191));
 sg13g2_and3_1 _6667_ (.X(_2223_),
    .A(net1948),
    .B(_1721_),
    .C(_1728_));
 sg13g2_nand2_2 _6668_ (.Y(_2224_),
    .A(net1947),
    .B(net1850));
 sg13g2_nor2_1 _6669_ (.A(_1805_),
    .B(_2224_),
    .Y(_2225_));
 sg13g2_nor4_1 _6670_ (.A(net1980),
    .B(_2222_),
    .C(_2223_),
    .D(_2225_),
    .Y(_2226_));
 sg13g2_o21ai_1 _6671_ (.B1(_2226_),
    .Y(_2227_),
    .A1(_1807_),
    .A2(_2219_));
 sg13g2_a21oi_2 _6672_ (.B1(_1782_),
    .Y(_2228_),
    .A2(_2227_),
    .A1(_2218_));
 sg13g2_nand3b_1 _6673_ (.B(_1706_),
    .C(_1767_),
    .Y(_2229_),
    .A_N(_0092_));
 sg13g2_nand2_1 _6674_ (.Y(_2230_),
    .A(_1684_),
    .B(_1787_));
 sg13g2_a21oi_1 _6675_ (.A1(_1684_),
    .A2(_1787_),
    .Y(_2231_),
    .B1(net2264));
 sg13g2_a21oi_1 _6676_ (.A1(net2264),
    .A2(_1644_),
    .Y(_2232_),
    .B1(_2231_));
 sg13g2_a21oi_1 _6677_ (.A1(_1640_),
    .A2(_1802_),
    .Y(_2233_),
    .B1(_2230_));
 sg13g2_o21ai_1 _6678_ (.B1(_1644_),
    .Y(_2234_),
    .A1(_1694_),
    .A2(net1856));
 sg13g2_o21ai_1 _6679_ (.B1(_2234_),
    .Y(_2235_),
    .A1(net2240),
    .A2(_2232_));
 sg13g2_o21ai_1 _6680_ (.B1(net1984),
    .Y(_2236_),
    .A1(net1944),
    .A2(_2233_));
 sg13g2_a221oi_1 _6681_ (.B2(net1888),
    .C1(_2236_),
    .B1(_2235_),
    .A1(net2088),
    .Y(_2237_),
    .A2(_2229_));
 sg13g2_nand2_2 _6682_ (.Y(_2238_),
    .A(_1642_),
    .B(_1809_));
 sg13g2_a21oi_1 _6683_ (.A1(_1765_),
    .A2(_2238_),
    .Y(_2239_),
    .B1(_1582_));
 sg13g2_and2_1 _6684_ (.A(net2240),
    .B(net2295),
    .X(_2240_));
 sg13g2_a221oi_1 _6685_ (.B2(net2216),
    .C1(_2239_),
    .B1(_2240_),
    .A1(net1853),
    .Y(_2241_),
    .A2(_2037_));
 sg13g2_nor2_1 _6686_ (.A(net2199),
    .B(_2241_),
    .Y(_2242_));
 sg13g2_o21ai_1 _6687_ (.B1(_1875_),
    .Y(_2243_),
    .A1(net2108),
    .A2(_2037_));
 sg13g2_o21ai_1 _6688_ (.B1(_1754_),
    .Y(_2244_),
    .A1(_2195_),
    .A2(_2243_));
 sg13g2_a22oi_1 _6689_ (.Y(_2245_),
    .B1(_2018_),
    .B2(net1849),
    .A2(net2010),
    .A1(net2295));
 sg13g2_a21oi_1 _6690_ (.A1(net1921),
    .A2(_1944_),
    .Y(_2246_),
    .B1(_1802_));
 sg13g2_a21oi_1 _6691_ (.A1(_2245_),
    .A2(_2246_),
    .Y(_2247_),
    .B1(net1944));
 sg13g2_nor3_1 _6692_ (.A(_2242_),
    .B(_2244_),
    .C(_2247_),
    .Y(_2248_));
 sg13g2_o21ai_1 _6693_ (.B1(net1770),
    .Y(_2249_),
    .A1(_2237_),
    .A2(_2248_));
 sg13g2_nand2_1 _6694_ (.Y(_2250_),
    .A(_1461_),
    .B(_1741_));
 sg13g2_a22oi_1 _6695_ (.Y(_2251_),
    .B1(_2250_),
    .B2(net2077),
    .A2(_2186_),
    .A1(_1708_));
 sg13g2_nor2_1 _6696_ (.A(_1775_),
    .B(_2185_),
    .Y(_2252_));
 sg13g2_nand3_1 _6697_ (.B(_1693_),
    .C(_1811_),
    .A(net1947),
    .Y(_2253_));
 sg13g2_a21oi_2 _6698_ (.B1(net2242),
    .Y(_2254_),
    .A2(net1903),
    .A1(net2260));
 sg13g2_a221oi_1 _6699_ (.B2(_1643_),
    .C1(_2253_),
    .B1(_2254_),
    .A1(net1838),
    .Y(_2255_),
    .A2(net1849));
 sg13g2_a21oi_1 _6700_ (.A1(net2016),
    .A2(_2251_),
    .Y(_2256_),
    .B1(_2255_));
 sg13g2_o21ai_1 _6701_ (.B1(_2256_),
    .Y(_2257_),
    .A1(_1720_),
    .A2(_2252_));
 sg13g2_nor3_1 _6702_ (.A(net1919),
    .B(net2002),
    .C(_1740_),
    .Y(_2258_));
 sg13g2_nor2_1 _6703_ (.A(net2233),
    .B(_1670_),
    .Y(_2259_));
 sg13g2_o21ai_1 _6704_ (.B1(net2214),
    .Y(_2260_),
    .A1(net2233),
    .A2(_1670_));
 sg13g2_nor2_1 _6705_ (.A(net2216),
    .B(net1826),
    .Y(_2261_));
 sg13g2_nor2_2 _6706_ (.A(net2255),
    .B(_1632_),
    .Y(_2262_));
 sg13g2_a22oi_1 _6707_ (.Y(_2263_),
    .B1(_2262_),
    .B2(net1999),
    .A2(_2261_),
    .A1(_1821_));
 sg13g2_a21o_1 _6708_ (.A2(_2263_),
    .A1(_2260_),
    .B1(_2258_),
    .X(_2264_));
 sg13g2_a22oi_1 _6709_ (.Y(_2265_),
    .B1(_2264_),
    .B2(_1856_),
    .A2(_2257_),
    .A1(net1940));
 sg13g2_o21ai_1 _6710_ (.B1(_2249_),
    .Y(_2266_),
    .A1(_1703_),
    .A2(_2265_));
 sg13g2_nor4_1 _6711_ (.A(_2163_),
    .B(_2205_),
    .C(_2228_),
    .D(_2266_),
    .Y(_2267_));
 sg13g2_nand4_1 _6712_ (.B(_2087_),
    .C(_2097_),
    .A(_2064_),
    .Y(_2268_),
    .D(_2267_));
 sg13g2_a21oi_1 _6713_ (.A1(_1564_),
    .A2(_1816_),
    .Y(_2269_),
    .B1(_2074_));
 sg13g2_nor4_1 _6714_ (.A(net1935),
    .B(_1590_),
    .C(_1835_),
    .D(_2269_),
    .Y(_2270_));
 sg13g2_a221oi_1 _6715_ (.B2(net1983),
    .C1(_2270_),
    .B1(_2167_),
    .A1(_1564_),
    .Y(_2271_),
    .A2(net1817));
 sg13g2_o21ai_1 _6716_ (.B1(_1449_),
    .Y(_2272_),
    .A1(net1756),
    .A2(_2271_));
 sg13g2_nor2_1 _6717_ (.A(_2268_),
    .B(_2272_),
    .Y(_2273_));
 sg13g2_nand3_1 _6718_ (.B(_1564_),
    .C(_2136_),
    .A(net1924),
    .Y(_2274_));
 sg13g2_a21oi_2 _6719_ (.B1(net2182),
    .Y(_2275_),
    .A2(_2274_),
    .A1(net2013));
 sg13g2_a21oi_2 _6720_ (.B1(net2082),
    .Y(_2276_),
    .A2(_1817_),
    .A1(net1918));
 sg13g2_a21oi_1 _6721_ (.A1(net2205),
    .A2(net1913),
    .Y(_2277_),
    .B1(net2187));
 sg13g2_nor2_1 _6722_ (.A(net2187),
    .B(_2276_),
    .Y(_2278_));
 sg13g2_a221oi_1 _6723_ (.B2(net1885),
    .C1(_2278_),
    .B1(_1921_),
    .A1(net1878),
    .Y(_2279_),
    .A2(_1657_));
 sg13g2_nand2b_1 _6724_ (.Y(_2280_),
    .B(_2275_),
    .A_N(_2279_));
 sg13g2_o21ai_1 _6725_ (.B1(net2193),
    .Y(_2281_),
    .A1(net1899),
    .A2(_1655_));
 sg13g2_inv_1 _6726_ (.Y(_2282_),
    .A(_2281_));
 sg13g2_nand2_2 _6727_ (.Y(_2283_),
    .A(net2022),
    .B(_1666_));
 sg13g2_a21oi_1 _6728_ (.A1(_1850_),
    .A2(_2283_),
    .Y(_2284_),
    .B1(_2172_));
 sg13g2_a21oi_1 _6729_ (.A1(net1910),
    .A2(net1838),
    .Y(_2285_),
    .B1(_2081_));
 sg13g2_nand2_1 _6730_ (.Y(_2286_),
    .A(net2089),
    .B(_2285_));
 sg13g2_o21ai_1 _6731_ (.B1(_2286_),
    .Y(_2287_),
    .A1(_2281_),
    .A2(_2284_));
 sg13g2_a221oi_1 _6732_ (.B2(net1938),
    .C1(_1583_),
    .B1(_2287_),
    .A1(net2092),
    .Y(_2288_),
    .A2(_2280_));
 sg13g2_nor2_1 _6733_ (.A(net1756),
    .B(_2288_),
    .Y(_2289_));
 sg13g2_nor2_1 _6734_ (.A(net2253),
    .B(net2029),
    .Y(_2290_));
 sg13g2_nand2_1 _6735_ (.Y(_2291_),
    .A(net1821),
    .B(_2290_));
 sg13g2_a21oi_1 _6736_ (.A1(_1998_),
    .A2(_2291_),
    .Y(_2292_),
    .B1(net2223));
 sg13g2_a21oi_1 _6737_ (.A1(_1786_),
    .A2(_1790_),
    .Y(_2293_),
    .B1(net2069));
 sg13g2_nor3_1 _6738_ (.A(net2203),
    .B(_2292_),
    .C(_2293_),
    .Y(_2294_));
 sg13g2_nor2_1 _6739_ (.A(net2192),
    .B(_2294_),
    .Y(_2295_));
 sg13g2_nor3_1 _6740_ (.A(net2000),
    .B(_1735_),
    .C(_1799_),
    .Y(_2296_));
 sg13g2_nor3_1 _6741_ (.A(net1980),
    .B(_1793_),
    .C(_2295_),
    .Y(_2297_));
 sg13g2_o21ai_1 _6742_ (.B1(_2297_),
    .Y(_2298_),
    .A1(net1986),
    .A2(_2296_));
 sg13g2_a21oi_2 _6743_ (.B1(net2243),
    .Y(_2299_),
    .A2(net1837),
    .A1(net2267));
 sg13g2_nand2_1 _6744_ (.Y(_2300_),
    .A(net1837),
    .B(_2165_));
 sg13g2_nand2b_1 _6745_ (.Y(_2301_),
    .B(_2299_),
    .A_N(_2207_));
 sg13g2_a22oi_1 _6746_ (.Y(_2302_),
    .B1(_2301_),
    .B2(_1958_),
    .A2(_2165_),
    .A1(net1836));
 sg13g2_a21o_1 _6747_ (.A2(_1716_),
    .A1(net1869),
    .B1(net2000),
    .X(_2303_));
 sg13g2_nor3_1 _6748_ (.A(net1942),
    .B(_1814_),
    .C(_2303_),
    .Y(_2304_));
 sg13g2_nor2_2 _6749_ (.A(net1925),
    .B(net1986),
    .Y(_2305_));
 sg13g2_o21ai_1 _6750_ (.B1(_2305_),
    .Y(_2306_),
    .A1(net2029),
    .A2(_1683_));
 sg13g2_o21ai_1 _6751_ (.B1(_2306_),
    .Y(_2307_),
    .A1(net2192),
    .A2(_2302_));
 sg13g2_o21ai_1 _6752_ (.B1(net1937),
    .Y(_2308_),
    .A1(_2304_),
    .A2(_2307_));
 sg13g2_a21o_2 _6753_ (.A2(_2308_),
    .A1(_2298_),
    .B1(_1782_),
    .X(_2309_));
 sg13g2_nand2_1 _6754_ (.Y(_2310_),
    .A(net1855),
    .B(_1896_));
 sg13g2_nor2b_2 _6755_ (.A(_2140_),
    .B_N(_2310_),
    .Y(_2311_));
 sg13g2_or3_1 _6756_ (.A(net2235),
    .B(_1682_),
    .C(_2207_),
    .X(_2312_));
 sg13g2_a22oi_1 _6757_ (.Y(_2313_),
    .B1(_2312_),
    .B2(_1958_),
    .A2(_2311_),
    .A1(_1895_));
 sg13g2_a22oi_1 _6758_ (.Y(_2314_),
    .B1(net1820),
    .B2(net1926),
    .A2(_1667_),
    .A1(net2066));
 sg13g2_a22oi_1 _6759_ (.Y(_2315_),
    .B1(_2299_),
    .B2(_2314_),
    .A2(_1804_),
    .A1(net1920));
 sg13g2_nand3_1 _6760_ (.B(net1859),
    .C(_1952_),
    .A(net1920),
    .Y(_2316_));
 sg13g2_a22oi_1 _6761_ (.Y(_2317_),
    .B1(_2316_),
    .B2(net1905),
    .A2(_2315_),
    .A1(net2015));
 sg13g2_o21ai_1 _6762_ (.B1(_2317_),
    .Y(_2318_),
    .A1(net2089),
    .A2(_2313_));
 sg13g2_a21oi_1 _6763_ (.A1(_1888_),
    .A2(_2164_),
    .Y(_2319_),
    .B1(net2197));
 sg13g2_o21ai_1 _6764_ (.B1(_2319_),
    .Y(_2320_),
    .A1(_1904_),
    .A2(_1942_));
 sg13g2_nand2_1 _6765_ (.Y(_2321_),
    .A(net2009),
    .B(net1880));
 sg13g2_a21oi_1 _6766_ (.A1(net2030),
    .A2(net1926),
    .Y(_2322_),
    .B1(net1881));
 sg13g2_a221oi_1 _6767_ (.B2(net1887),
    .C1(net1982),
    .B1(_2322_),
    .A1(net2197),
    .Y(_2323_),
    .A2(_1969_));
 sg13g2_and2_1 _6768_ (.A(_2320_),
    .B(_2323_),
    .X(_2324_));
 sg13g2_a221oi_1 _6769_ (.B2(net1939),
    .C1(_2324_),
    .B1(_2318_),
    .A1(_1888_),
    .Y(_2325_),
    .A2(net1817));
 sg13g2_o21ai_1 _6770_ (.B1(_2309_),
    .Y(_2326_),
    .A1(_1936_),
    .A2(_2325_));
 sg13g2_o21ai_1 _6771_ (.B1(net2233),
    .Y(_2327_),
    .A1(_1650_),
    .A2(_1671_));
 sg13g2_o21ai_1 _6772_ (.B1(_2327_),
    .Y(_2328_),
    .A1(net2233),
    .A2(net1918));
 sg13g2_nor2_1 _6773_ (.A(net2222),
    .B(net1833),
    .Y(_2329_));
 sg13g2_a22oi_1 _6774_ (.Y(_2330_),
    .B1(net1865),
    .B2(net1874),
    .A2(net1833),
    .A1(net2208));
 sg13g2_o21ai_1 _6775_ (.B1(_2330_),
    .Y(_2331_),
    .A1(_1582_),
    .A2(_1624_));
 sg13g2_nand2_1 _6776_ (.Y(_2332_),
    .A(net2089),
    .B(_2331_));
 sg13g2_o21ai_1 _6777_ (.B1(_2332_),
    .Y(_2333_),
    .A1(_2056_),
    .A2(_2329_));
 sg13g2_a21o_1 _6778_ (.A2(_2328_),
    .A1(net1886),
    .B1(_2333_),
    .X(_2334_));
 sg13g2_nand2_1 _6779_ (.Y(_2335_),
    .A(net1873),
    .B(_1750_));
 sg13g2_a21oi_1 _6780_ (.A1(_1965_),
    .A2(_2335_),
    .Y(_2336_),
    .B1(_2195_));
 sg13g2_nor2_1 _6781_ (.A(net2183),
    .B(_2336_),
    .Y(_2337_));
 sg13g2_nand3_1 _6782_ (.B(net1879),
    .C(_1644_),
    .A(net2011),
    .Y(_2338_));
 sg13g2_o21ai_1 _6783_ (.B1(_2338_),
    .Y(_2339_),
    .A1(net2011),
    .A2(net1923));
 sg13g2_a22oi_1 _6784_ (.Y(_2340_),
    .B1(_2339_),
    .B2(net1907),
    .A2(_1906_),
    .A1(net2015));
 sg13g2_nand3_1 _6785_ (.B(_2337_),
    .C(_2340_),
    .A(_1902_),
    .Y(_2341_));
 sg13g2_a221oi_1 _6786_ (.B2(net2093),
    .C1(_2066_),
    .B1(_2341_),
    .A1(net1939),
    .Y(_2342_),
    .A2(_2334_));
 sg13g2_o21ai_1 _6787_ (.B1(net1858),
    .Y(_2343_),
    .A1(net2071),
    .A2(_1437_));
 sg13g2_a21oi_1 _6788_ (.A1(net1950),
    .A2(_2343_),
    .Y(_2344_),
    .B1(net1982));
 sg13g2_o21ai_1 _6789_ (.B1(_2121_),
    .Y(_2345_),
    .A1(net1881),
    .A2(_1649_));
 sg13g2_a21oi_1 _6790_ (.A1(_1883_),
    .A2(_2345_),
    .Y(_2346_),
    .B1(_1881_));
 sg13g2_nand4_1 _6791_ (.B(_1891_),
    .C(_2344_),
    .A(_1873_),
    .Y(_2347_),
    .D(_2346_));
 sg13g2_o21ai_1 _6792_ (.B1(net2234),
    .Y(_2348_),
    .A1(_1672_),
    .A2(_1977_));
 sg13g2_a221oi_1 _6793_ (.B2(_2348_),
    .C1(net2186),
    .B1(_1976_),
    .A1(net1988),
    .Y(_2349_),
    .A2(net1858));
 sg13g2_or2_1 _6794_ (.X(_2350_),
    .B(_2349_),
    .A(_1975_));
 sg13g2_a21oi_1 _6795_ (.A1(_2347_),
    .A2(_2350_),
    .Y(_2351_),
    .B1(_1861_));
 sg13g2_nor3_1 _6796_ (.A(net2001),
    .B(net1824),
    .C(_1713_),
    .Y(_2352_));
 sg13g2_a21oi_2 _6797_ (.B1(_1805_),
    .Y(_2353_),
    .A2(_2032_),
    .A1(net2105));
 sg13g2_a221oi_1 _6798_ (.B2(_1888_),
    .C1(_2353_),
    .B1(net1848),
    .A1(net2009),
    .Y(_2354_),
    .A2(_1982_));
 sg13g2_nor2_1 _6799_ (.A(net2081),
    .B(_2354_),
    .Y(_2355_));
 sg13g2_a21oi_2 _6800_ (.B1(net2238),
    .Y(_2356_),
    .A2(net1814),
    .A1(net2262));
 sg13g2_a21oi_1 _6801_ (.A1(_1983_),
    .A2(_2356_),
    .Y(_2357_),
    .B1(_1675_));
 sg13g2_nor3_1 _6802_ (.A(net2191),
    .B(_2355_),
    .C(_2357_),
    .Y(_2358_));
 sg13g2_o21ai_1 _6803_ (.B1(net1941),
    .Y(_2359_),
    .A1(_2352_),
    .A2(_2358_));
 sg13g2_a21oi_1 _6804_ (.A1(_1764_),
    .A2(_1919_),
    .Y(_2360_),
    .B1(net1917));
 sg13g2_nand2_1 _6805_ (.Y(_2361_),
    .A(net1909),
    .B(_2360_));
 sg13g2_a21o_1 _6806_ (.A2(_2041_),
    .A1(net2080),
    .B1(net1868),
    .X(_2362_));
 sg13g2_o21ai_1 _6807_ (.B1(net2231),
    .Y(_2363_),
    .A1(net2255),
    .A2(net1820));
 sg13g2_o21ai_1 _6808_ (.B1(_2362_),
    .Y(_2364_),
    .A1(_2143_),
    .A2(_2363_));
 sg13g2_nor2_1 _6809_ (.A(net1917),
    .B(net1903),
    .Y(_2365_));
 sg13g2_o21ai_1 _6810_ (.B1(net1853),
    .Y(_2366_),
    .A1(_2130_),
    .A2(_2365_));
 sg13g2_nand4_1 _6811_ (.B(_2361_),
    .C(_2364_),
    .A(_1856_),
    .Y(_2367_),
    .D(_2366_));
 sg13g2_a21oi_1 _6812_ (.A1(_2359_),
    .A2(_2367_),
    .Y(_2368_),
    .B1(_1703_));
 sg13g2_nor2_2 _6813_ (.A(net1822),
    .B(_2119_),
    .Y(_2369_));
 sg13g2_nor3_1 _6814_ (.A(_1427_),
    .B(_1927_),
    .C(_2369_),
    .Y(_2370_));
 sg13g2_nor2_1 _6815_ (.A(net2193),
    .B(_1637_),
    .Y(_2371_));
 sg13g2_or3_1 _6816_ (.A(_2260_),
    .B(_2370_),
    .C(_2371_),
    .X(_2372_));
 sg13g2_a221oi_1 _6817_ (.B2(_2135_),
    .C1(_1475_),
    .B1(_1850_),
    .A1(_1695_),
    .Y(_2373_),
    .A2(_1844_));
 sg13g2_a21oi_1 _6818_ (.A1(net1918),
    .A2(net1892),
    .Y(_2374_),
    .B1(net1876));
 sg13g2_o21ai_1 _6819_ (.B1(net1939),
    .Y(_2375_),
    .A1(net1946),
    .A2(_2374_));
 sg13g2_nor2_1 _6820_ (.A(_2373_),
    .B(_2375_),
    .Y(_2376_));
 sg13g2_a22oi_1 _6821_ (.Y(_2377_),
    .B1(net1822),
    .B2(_1834_),
    .A2(net1886),
    .A1(net2073));
 sg13g2_nand2_1 _6822_ (.Y(_2378_),
    .A(net2193),
    .B(_1928_));
 sg13g2_nand3_1 _6823_ (.B(_1844_),
    .C(_1890_),
    .A(net1912),
    .Y(_2379_));
 sg13g2_and4_1 _6824_ (.A(_2118_),
    .B(_2275_),
    .C(_2378_),
    .D(_2379_),
    .X(_2380_));
 sg13g2_o21ai_1 _6825_ (.B1(_2380_),
    .Y(_2381_),
    .A1(_2369_),
    .A2(_2377_));
 sg13g2_a221oi_1 _6826_ (.B2(net2092),
    .C1(_1920_),
    .B1(_2381_),
    .A1(_2372_),
    .Y(_2382_),
    .A2(_2376_));
 sg13g2_nor2_1 _6827_ (.A(_2368_),
    .B(_2382_),
    .Y(_2383_));
 sg13g2_a221oi_1 _6828_ (.B2(net1875),
    .C1(net1824),
    .B1(net2004),
    .A1(net2252),
    .Y(_2384_),
    .A2(net2074));
 sg13g2_or2_2 _6829_ (.X(_2385_),
    .B(_1737_),
    .A(net1838));
 sg13g2_nor2_2 _6830_ (.A(net2218),
    .B(_1944_),
    .Y(_2386_));
 sg13g2_nand2_2 _6831_ (.Y(_2387_),
    .A(_2385_),
    .B(_2386_));
 sg13g2_mux2_2 _6832_ (.A0(net2284),
    .A1(_0096_),
    .S(net2296),
    .X(_2388_));
 sg13g2_a21oi_2 _6833_ (.B1(_2192_),
    .Y(_2389_),
    .A2(_2388_),
    .A1(net2256));
 sg13g2_a22oi_1 _6834_ (.Y(_2390_),
    .B1(net1853),
    .B2(_2389_),
    .A2(net1909),
    .A1(net1917));
 sg13g2_a21oi_1 _6835_ (.A1(_2387_),
    .A2(_2390_),
    .Y(_2391_),
    .B1(net2199));
 sg13g2_o21ai_1 _6836_ (.B1(net1940),
    .Y(_2392_),
    .A1(_2384_),
    .A2(_2391_));
 sg13g2_o21ai_1 _6837_ (.B1(net1853),
    .Y(_2393_),
    .A1(_2148_),
    .A2(_2262_));
 sg13g2_nand2_2 _6838_ (.Y(_2394_),
    .A(net2255),
    .B(net1833));
 sg13g2_o21ai_1 _6839_ (.B1(_1999_),
    .Y(_2395_),
    .A1(net1820),
    .A2(_2394_));
 sg13g2_a21oi_1 _6840_ (.A1(net1865),
    .A2(_2395_),
    .Y(_2396_),
    .B1(_1857_));
 sg13g2_nor2_2 _6841_ (.A(_1775_),
    .B(_2369_),
    .Y(_2397_));
 sg13g2_a22oi_1 _6842_ (.Y(_2398_),
    .B1(_2397_),
    .B2(net1996),
    .A2(_1687_),
    .A1(net1910));
 sg13g2_nand3_1 _6843_ (.B(_2396_),
    .C(_2398_),
    .A(_2393_),
    .Y(_2399_));
 sg13g2_nand2_1 _6844_ (.Y(_2400_),
    .A(_2392_),
    .B(_2399_));
 sg13g2_nand3_1 _6845_ (.B(_1642_),
    .C(_1809_),
    .A(net2244),
    .Y(_2401_));
 sg13g2_nor2_1 _6846_ (.A(net2292),
    .B(_1690_),
    .Y(_2402_));
 sg13g2_o21ai_1 _6847_ (.B1(_2401_),
    .Y(_2403_),
    .A1(net2243),
    .A2(_2402_));
 sg13g2_nor2_1 _6848_ (.A(_2152_),
    .B(_2403_),
    .Y(_2404_));
 sg13g2_nor2_1 _6849_ (.A(net1990),
    .B(_2404_),
    .Y(_2405_));
 sg13g2_nor2_2 _6850_ (.A(net2243),
    .B(_1769_),
    .Y(_2406_));
 sg13g2_nand2_1 _6851_ (.Y(_2407_),
    .A(net1985),
    .B(net1855));
 sg13g2_nand3_1 _6852_ (.B(net1862),
    .C(_2407_),
    .A(_1693_),
    .Y(_2408_));
 sg13g2_o21ai_1 _6853_ (.B1(net1864),
    .Y(_2409_),
    .A1(_2406_),
    .A2(_2408_));
 sg13g2_o21ai_1 _6854_ (.B1(_2409_),
    .Y(_2410_),
    .A1(net1945),
    .A2(_1776_));
 sg13g2_o21ai_1 _6855_ (.B1(net1998),
    .Y(_2411_),
    .A1(_1746_),
    .A2(_2131_));
 sg13g2_o21ai_1 _6856_ (.B1(_2411_),
    .Y(_2412_),
    .A1(net2217),
    .A2(_1734_));
 sg13g2_a21oi_1 _6857_ (.A1(net2217),
    .A2(_1744_),
    .Y(_2413_),
    .B1(_2412_));
 sg13g2_nor2_2 _6858_ (.A(net1942),
    .B(net1991),
    .Y(_2414_));
 sg13g2_a22oi_1 _6859_ (.Y(_2415_),
    .B1(_2250_),
    .B2(_2414_),
    .A2(_1657_),
    .A1(net1870));
 sg13g2_and2_1 _6860_ (.A(_1754_),
    .B(_2415_),
    .X(_2416_));
 sg13g2_o21ai_1 _6861_ (.B1(_2416_),
    .Y(_2417_),
    .A1(net2200),
    .A2(_2413_));
 sg13g2_o21ai_1 _6862_ (.B1(_2417_),
    .Y(_2418_),
    .A1(_2405_),
    .A2(_2410_));
 sg13g2_a221oi_1 _6863_ (.B2(net1770),
    .C1(_1538_),
    .B1(_2418_),
    .A1(net1771),
    .Y(_2419_),
    .A2(_2400_));
 sg13g2_nand3_1 _6864_ (.B(net1833),
    .C(net1859),
    .A(net1891),
    .Y(_2420_));
 sg13g2_nand4_1 _6865_ (.B(_1803_),
    .C(_1991_),
    .A(net1861),
    .Y(_2421_),
    .D(_2420_));
 sg13g2_nand2_1 _6866_ (.Y(_2422_),
    .A(_1770_),
    .B(net1818));
 sg13g2_nor2_1 _6867_ (.A(net2267),
    .B(_2422_),
    .Y(_2423_));
 sg13g2_a21oi_1 _6868_ (.A1(net2005),
    .A2(_1746_),
    .Y(_2424_),
    .B1(_2423_));
 sg13g2_nand2_1 _6869_ (.Y(_2425_),
    .A(net2074),
    .B(_2207_));
 sg13g2_a22oi_1 _6870_ (.Y(_2426_),
    .B1(_2425_),
    .B2(_1968_),
    .A2(_2134_),
    .A1(_1684_));
 sg13g2_o21ai_1 _6871_ (.B1(_2426_),
    .Y(_2427_),
    .A1(net2003),
    .A2(_2424_));
 sg13g2_a22oi_1 _6872_ (.Y(_2428_),
    .B1(_2427_),
    .B2(net2191),
    .A2(_2421_),
    .A1(net1863));
 sg13g2_o21ai_1 _6873_ (.B1(net1906),
    .Y(_2429_),
    .A1(net1993),
    .A2(net1860));
 sg13g2_nand3_1 _6874_ (.B(net1948),
    .C(net1859),
    .A(net2070),
    .Y(_2430_));
 sg13g2_o21ai_1 _6875_ (.B1(net2014),
    .Y(_2431_),
    .A1(net1890),
    .A2(net1869));
 sg13g2_nand3_1 _6876_ (.B(_2430_),
    .C(_2431_),
    .A(_2429_),
    .Y(_2432_));
 sg13g2_a22oi_1 _6877_ (.Y(_2433_),
    .B1(_2262_),
    .B2(_1804_),
    .A2(_1997_),
    .A1(net1890));
 sg13g2_o21ai_1 _6878_ (.B1(_2005_),
    .Y(_2434_),
    .A1(net1943),
    .A2(_2433_));
 sg13g2_a21oi_1 _6879_ (.A1(net2005),
    .A2(_2432_),
    .Y(_2435_),
    .B1(_2434_));
 sg13g2_o21ai_1 _6880_ (.B1(_1981_),
    .Y(_2436_),
    .A1(_2428_),
    .A2(_2435_));
 sg13g2_a21oi_1 _6881_ (.A1(net2233),
    .A2(_1836_),
    .Y(_2437_),
    .B1(_2259_));
 sg13g2_nor2_1 _6882_ (.A(net1904),
    .B(_2437_),
    .Y(_2438_));
 sg13g2_o21ai_1 _6883_ (.B1(_1833_),
    .Y(_2439_),
    .A1(net1929),
    .A2(net1917));
 sg13g2_o21ai_1 _6884_ (.B1(net1938),
    .Y(_2440_),
    .A1(_2438_),
    .A2(_2439_));
 sg13g2_o21ai_1 _6885_ (.B1(net2080),
    .Y(_2441_),
    .A1(net2009),
    .A2(net1897));
 sg13g2_o21ai_1 _6886_ (.B1(net2208),
    .Y(_2442_),
    .A1(net1897),
    .A2(net1891));
 sg13g2_a21oi_1 _6887_ (.A1(_2441_),
    .A2(_2442_),
    .Y(_2443_),
    .B1(_1832_));
 sg13g2_o21ai_1 _6888_ (.B1(net2091),
    .Y(_2444_),
    .A1(_1566_),
    .A2(_2443_));
 sg13g2_nand3_1 _6889_ (.B(_2440_),
    .C(_2444_),
    .A(_1831_),
    .Y(_2445_));
 sg13g2_nand4_1 _6890_ (.B(_2419_),
    .C(_2436_),
    .A(_2383_),
    .Y(_2446_),
    .D(_2445_));
 sg13g2_nor4_2 _6891_ (.A(_2326_),
    .B(_2342_),
    .C(_2351_),
    .Y(_2447_),
    .D(_2446_));
 sg13g2_o21ai_1 _6892_ (.B1(_1450_),
    .Y(_2448_),
    .A1(_2289_),
    .A2(_2447_));
 sg13g2_o21ai_1 _6893_ (.B1(_2007_),
    .Y(_2449_),
    .A1(_4055_),
    .A2(net1854));
 sg13g2_o21ai_1 _6894_ (.B1(_2406_),
    .Y(_2450_),
    .A1(net2267),
    .A2(net1818));
 sg13g2_a22oi_1 _6895_ (.Y(_2451_),
    .B1(net1855),
    .B2(_1938_),
    .A2(net1869),
    .A1(net1893));
 sg13g2_nand3_1 _6896_ (.B(_2450_),
    .C(_2451_),
    .A(net2217),
    .Y(_2452_));
 sg13g2_a21oi_1 _6897_ (.A1(_2449_),
    .A2(_2452_),
    .Y(_2453_),
    .B1(net1863));
 sg13g2_nor2_2 _6898_ (.A(net1871),
    .B(_1998_),
    .Y(_2454_));
 sg13g2_o21ai_1 _6899_ (.B1(_1431_),
    .Y(_2455_),
    .A1(_2059_),
    .A2(_2454_));
 sg13g2_a21oi_2 _6900_ (.B1(_1667_),
    .Y(_2456_),
    .A2(net1832),
    .A1(net2255));
 sg13g2_nor2_1 _6901_ (.A(_2430_),
    .B(_2456_),
    .Y(_2457_));
 sg13g2_nand3_1 _6902_ (.B(_1764_),
    .C(_1965_),
    .A(net2245),
    .Y(_2458_));
 sg13g2_a21oi_2 _6903_ (.B1(net1931),
    .Y(_2459_),
    .A2(_2458_),
    .A1(_2402_));
 sg13g2_a221oi_1 _6904_ (.B2(_1437_),
    .C1(net1904),
    .B1(_1944_),
    .A1(net2074),
    .Y(_2460_),
    .A2(net1919));
 sg13g2_nor4_1 _6905_ (.A(_2006_),
    .B(_2457_),
    .C(_2459_),
    .D(_2460_),
    .Y(_2461_));
 sg13g2_nand3_1 _6906_ (.B(_1684_),
    .C(net1857),
    .A(_1435_),
    .Y(_2462_));
 sg13g2_a221oi_1 _6907_ (.B2(net2069),
    .C1(_1992_),
    .B1(_1997_),
    .A1(net1891),
    .Y(_2463_),
    .A2(net1869));
 sg13g2_a221oi_1 _6908_ (.B2(_2463_),
    .C1(_2453_),
    .B1(_2462_),
    .A1(_2455_),
    .Y(_2464_),
    .A2(_2461_));
 sg13g2_nor2_1 _6909_ (.A(_1859_),
    .B(_2464_),
    .Y(_2465_));
 sg13g2_nor2_2 _6910_ (.A(net2081),
    .B(net1890),
    .Y(_2466_));
 sg13g2_a22oi_1 _6911_ (.Y(_2467_),
    .B1(_2466_),
    .B2(net1836),
    .A2(_2207_),
    .A1(net1868));
 sg13g2_o21ai_1 _6912_ (.B1(_2467_),
    .Y(_2468_),
    .A1(_1582_),
    .A2(_2397_));
 sg13g2_nor2_1 _6913_ (.A(_2276_),
    .B(_2362_),
    .Y(_2469_));
 sg13g2_a22oi_1 _6914_ (.Y(_2470_),
    .B1(_2469_),
    .B2(_1701_),
    .A2(_2468_),
    .A1(_1662_));
 sg13g2_nor2_1 _6915_ (.A(_1857_),
    .B(_2470_),
    .Y(_2471_));
 sg13g2_nor3_1 _6916_ (.A(net2001),
    .B(net1824),
    .C(net1823),
    .Y(_2472_));
 sg13g2_nor4_1 _6917_ (.A(net2188),
    .B(net2204),
    .C(net1920),
    .D(_1816_),
    .Y(_2473_));
 sg13g2_a21o_1 _6918_ (.A2(_2473_),
    .A1(_1693_),
    .B1(_2472_),
    .X(_2474_));
 sg13g2_o21ai_1 _6919_ (.B1(net2209),
    .Y(_2475_),
    .A1(_1547_),
    .A2(_2207_));
 sg13g2_nor2_1 _6920_ (.A(net2000),
    .B(_2041_),
    .Y(_2476_));
 sg13g2_a22oi_1 _6921_ (.Y(_2477_),
    .B1(_1656_),
    .B2(_2476_),
    .A2(net1836),
    .A1(net1840));
 sg13g2_a21oi_1 _6922_ (.A1(_2475_),
    .A2(_2477_),
    .Y(_2478_),
    .B1(net1883));
 sg13g2_a22oi_1 _6923_ (.Y(_2479_),
    .B1(_2478_),
    .B2(_1701_),
    .A2(_2474_),
    .A1(_1662_));
 sg13g2_nor2_1 _6924_ (.A(net1933),
    .B(_2479_),
    .Y(_2480_));
 sg13g2_nor3_1 _6925_ (.A(_2465_),
    .B(_2471_),
    .C(_2480_),
    .Y(_2481_));
 sg13g2_or2_1 _6926_ (.X(_2482_),
    .B(_2481_),
    .A(_1535_));
 sg13g2_a21oi_1 _6927_ (.A1(net2294),
    .A2(_1639_),
    .Y(_2483_),
    .B1(net1992));
 sg13g2_a22oi_1 _6928_ (.Y(_2484_),
    .B1(_2483_),
    .B2(net1914),
    .A2(_2230_),
    .A1(net1995));
 sg13g2_nor2_1 _6929_ (.A(net1929),
    .B(_2484_),
    .Y(_2485_));
 sg13g2_o21ai_1 _6930_ (.B1(_1833_),
    .Y(_2486_),
    .A1(net2189),
    .A2(_2437_));
 sg13g2_o21ai_1 _6931_ (.B1(net1938),
    .Y(_2487_),
    .A1(_2485_),
    .A2(_2486_));
 sg13g2_nor2_1 _6932_ (.A(net1909),
    .B(net1897),
    .Y(_2488_));
 sg13g2_a21oi_1 _6933_ (.A1(net2208),
    .A2(_1588_),
    .Y(_2489_),
    .B1(_1565_));
 sg13g2_o21ai_1 _6934_ (.B1(_1559_),
    .Y(_2490_),
    .A1(_1832_),
    .A2(_2488_));
 sg13g2_o21ai_1 _6935_ (.B1(net2092),
    .Y(_2491_),
    .A1(_2489_),
    .A2(_2490_));
 sg13g2_nand3_1 _6936_ (.B(_2487_),
    .C(_2491_),
    .A(_1831_),
    .Y(_2492_));
 sg13g2_o21ai_1 _6937_ (.B1(net1947),
    .Y(_2493_),
    .A1(net2224),
    .A2(net1871));
 sg13g2_a221oi_1 _6938_ (.B2(_1735_),
    .C1(net1930),
    .B1(net1821),
    .A1(net2225),
    .Y(_2494_),
    .A2(net1835));
 sg13g2_nand2_2 _6939_ (.Y(_2495_),
    .A(_1684_),
    .B(_1721_));
 sg13g2_a21oi_1 _6940_ (.A1(_2305_),
    .A2(_2495_),
    .Y(_2496_),
    .B1(_2494_));
 sg13g2_o21ai_1 _6941_ (.B1(_2496_),
    .Y(_2497_),
    .A1(_1814_),
    .A2(_2493_));
 sg13g2_a21oi_2 _6942_ (.B1(net2029),
    .Y(_2498_),
    .A2(_1676_),
    .A1(net2256));
 sg13g2_o21ai_1 _6943_ (.B1(net1883),
    .Y(_2499_),
    .A1(_2303_),
    .A2(_2498_));
 sg13g2_a21oi_1 _6944_ (.A1(net1821),
    .A2(_2290_),
    .Y(_2500_),
    .B1(_2454_));
 sg13g2_o21ai_1 _6945_ (.B1(_2147_),
    .Y(_2501_),
    .A1(_1683_),
    .A2(_1686_));
 sg13g2_a21oi_1 _6946_ (.A1(net2225),
    .A2(_2501_),
    .Y(_2502_),
    .B1(_1992_));
 sg13g2_o21ai_1 _6947_ (.B1(_2502_),
    .Y(_2503_),
    .A1(net2223),
    .A2(_2500_));
 sg13g2_o21ai_1 _6948_ (.B1(_2503_),
    .Y(_2504_),
    .A1(net1863),
    .A2(_1968_));
 sg13g2_a22oi_1 _6949_ (.Y(_2505_),
    .B1(_2499_),
    .B2(_2504_),
    .A2(_2497_),
    .A1(net1937));
 sg13g2_or2_1 _6950_ (.X(_2506_),
    .B(_2505_),
    .A(_1782_));
 sg13g2_a21oi_1 _6951_ (.A1(net1878),
    .A2(_1654_),
    .Y(_2507_),
    .B1(_1832_));
 sg13g2_a221oi_1 _6952_ (.B2(net1912),
    .C1(_2507_),
    .B1(_1890_),
    .A1(net1905),
    .Y(_2508_),
    .A2(net1823));
 sg13g2_a21oi_1 _6953_ (.A1(_2275_),
    .A2(_2508_),
    .Y(_2509_),
    .B1(net2180));
 sg13g2_nand3_1 _6954_ (.B(_1850_),
    .C(_2283_),
    .A(net2237),
    .Y(_2510_));
 sg13g2_nand3_1 _6955_ (.B(_1863_),
    .C(_2510_),
    .A(net2211),
    .Y(_2511_));
 sg13g2_a21oi_1 _6956_ (.A1(net1926),
    .A2(net1838),
    .Y(_2512_),
    .B1(_1552_));
 sg13g2_a221oi_1 _6957_ (.B2(_2511_),
    .C1(_2512_),
    .B1(_2282_),
    .A1(net2015),
    .Y(_2513_),
    .A2(_1548_));
 sg13g2_nor3_1 _6958_ (.A(net1757),
    .B(_1583_),
    .C(_2509_),
    .Y(_2514_));
 sg13g2_o21ai_1 _6959_ (.B1(_2514_),
    .Y(_2515_),
    .A1(net1932),
    .A2(_2513_));
 sg13g2_nor2_1 _6960_ (.A(net2254),
    .B(_1853_),
    .Y(_2516_));
 sg13g2_nor2_1 _6961_ (.A(net1851),
    .B(_2516_),
    .Y(_2517_));
 sg13g2_nand2_1 _6962_ (.Y(_2518_),
    .A(net1868),
    .B(_2147_));
 sg13g2_nand3_1 _6963_ (.B(_1686_),
    .C(_2394_),
    .A(net1909),
    .Y(_2519_));
 sg13g2_o21ai_1 _6964_ (.B1(_2519_),
    .Y(_2520_),
    .A1(_2262_),
    .A2(_2518_));
 sg13g2_a221oi_1 _6965_ (.B2(_1919_),
    .C1(_2520_),
    .B1(_2517_),
    .A1(net1996),
    .Y(_2521_),
    .A2(net1813));
 sg13g2_nor2_1 _6966_ (.A(net2190),
    .B(_2521_),
    .Y(_2522_));
 sg13g2_nand2_1 _6967_ (.Y(_2523_),
    .A(_1461_),
    .B(_2414_));
 sg13g2_nand3_1 _6968_ (.B(_2179_),
    .C(_2414_),
    .A(_1461_),
    .Y(_2524_));
 sg13g2_a221oi_1 _6969_ (.B2(_1578_),
    .C1(_2522_),
    .B1(_2305_),
    .A1(net1834),
    .Y(_2525_),
    .A2(_1657_));
 sg13g2_a21oi_1 _6970_ (.A1(_2524_),
    .A2(_2525_),
    .Y(_2526_),
    .B1(net1932));
 sg13g2_nand2_1 _6971_ (.Y(_2527_),
    .A(_1822_),
    .B(_2262_));
 sg13g2_nand4_1 _6972_ (.B(_2150_),
    .C(_2420_),
    .A(net1861),
    .Y(_2528_),
    .D(_2527_));
 sg13g2_nand2_1 _6973_ (.Y(_2529_),
    .A(_1430_),
    .B(_2056_));
 sg13g2_nor2_2 _6974_ (.A(net2253),
    .B(net1832),
    .Y(_2530_));
 sg13g2_nor2_1 _6975_ (.A(net1837),
    .B(_2530_),
    .Y(_2531_));
 sg13g2_a22oi_1 _6976_ (.Y(_2532_),
    .B1(_2531_),
    .B2(_1883_),
    .A2(_2529_),
    .A1(net2005));
 sg13g2_o21ai_1 _6977_ (.B1(_2532_),
    .Y(_2533_),
    .A1(_1880_),
    .A2(_2456_));
 sg13g2_a21oi_1 _6978_ (.A1(net1863),
    .A2(_2528_),
    .Y(_2534_),
    .B1(_2533_));
 sg13g2_o21ai_1 _6979_ (.B1(net1770),
    .Y(_2535_),
    .A1(_2526_),
    .A2(_2534_));
 sg13g2_a221oi_1 _6980_ (.B2(_1834_),
    .C1(net1980),
    .B1(net1833),
    .A1(net2251),
    .Y(_2536_),
    .A2(_1557_));
 sg13g2_o21ai_1 _6981_ (.B1(_2536_),
    .Y(_2537_),
    .A1(net1929),
    .A2(_2113_));
 sg13g2_nand2_1 _6982_ (.Y(_2538_),
    .A(_1708_),
    .B(_1867_));
 sg13g2_and2_1 _6983_ (.A(_1890_),
    .B(_2538_),
    .X(_2539_));
 sg13g2_a21oi_1 _6984_ (.A1(net1993),
    .A2(net1834),
    .Y(_2540_),
    .B1(_1794_));
 sg13g2_nor3_1 _6985_ (.A(net1895),
    .B(_1691_),
    .C(_1716_),
    .Y(_2541_));
 sg13g2_nor3_1 _6986_ (.A(net1988),
    .B(_1775_),
    .C(_2541_),
    .Y(_2542_));
 sg13g2_nor4_1 _6987_ (.A(_2537_),
    .B(_2539_),
    .C(_2540_),
    .D(_2542_),
    .Y(_2543_));
 sg13g2_nor2_1 _6988_ (.A(net2224),
    .B(_1545_),
    .Y(_2544_));
 sg13g2_nand2_1 _6989_ (.Y(_2545_),
    .A(net2073),
    .B(net1911));
 sg13g2_o21ai_1 _6990_ (.B1(_1804_),
    .Y(_2546_),
    .A1(net2106),
    .A2(_1681_));
 sg13g2_a21oi_1 _6991_ (.A1(_2545_),
    .A2(_2546_),
    .Y(_2547_),
    .B1(net1904));
 sg13g2_a21oi_1 _6992_ (.A1(_1666_),
    .A2(_2113_),
    .Y(_2548_),
    .B1(_1884_));
 sg13g2_a21oi_1 _6993_ (.A1(net2289),
    .A2(_1728_),
    .Y(_2549_),
    .B1(_2056_));
 sg13g2_nand2_1 _6994_ (.Y(_2550_),
    .A(net2075),
    .B(net1985));
 sg13g2_nand3_1 _6995_ (.B(_1546_),
    .C(_2550_),
    .A(net2015),
    .Y(_2551_));
 sg13g2_o21ai_1 _6996_ (.B1(_2551_),
    .Y(_2552_),
    .A1(net1877),
    .A2(_1880_));
 sg13g2_nor4_1 _6997_ (.A(_2547_),
    .B(_2548_),
    .C(_2549_),
    .D(_2552_),
    .Y(_2553_));
 sg13g2_nor2_1 _6998_ (.A(net2257),
    .B(_2113_),
    .Y(_2554_));
 sg13g2_nor2_1 _6999_ (.A(_2114_),
    .B(_2143_),
    .Y(_2555_));
 sg13g2_a221oi_1 _7000_ (.B2(net1817),
    .C1(_2543_),
    .B1(_2555_),
    .A1(net1939),
    .Y(_2556_),
    .A2(_2553_));
 sg13g2_or2_1 _7001_ (.X(_2557_),
    .B(_2556_),
    .A(_1936_));
 sg13g2_o21ai_1 _7002_ (.B1(_1884_),
    .Y(_2558_),
    .A1(net1840),
    .A2(_1670_));
 sg13g2_o21ai_1 _7003_ (.B1(_2558_),
    .Y(_2559_),
    .A1(_1836_),
    .A2(_1884_));
 sg13g2_nand2_2 _7004_ (.Y(_2560_),
    .A(net1899),
    .B(_1850_));
 sg13g2_inv_1 _7005_ (.Y(_2561_),
    .A(_2560_));
 sg13g2_a22oi_1 _7006_ (.Y(_2562_),
    .B1(_2561_),
    .B2(net1840),
    .A2(_1839_),
    .A1(net2185));
 sg13g2_nand3_1 _7007_ (.B(_2559_),
    .C(_2562_),
    .A(net2180),
    .Y(_2563_));
 sg13g2_nor2_1 _7008_ (.A(net1931),
    .B(_2070_),
    .Y(_2564_));
 sg13g2_o21ai_1 _7009_ (.B1(_2564_),
    .Y(_2565_),
    .A1(net2073),
    .A2(_2561_));
 sg13g2_nand3_1 _7010_ (.B(net2002),
    .C(net1822),
    .A(net2193),
    .Y(_2566_));
 sg13g2_a21oi_1 _7011_ (.A1(net1907),
    .A2(net1822),
    .Y(_2567_),
    .B1(net1981));
 sg13g2_nand4_1 _7012_ (.B(_2565_),
    .C(_2566_),
    .A(_2378_),
    .Y(_2568_),
    .D(_2567_));
 sg13g2_a21o_1 _7013_ (.A2(_2568_),
    .A1(_2563_),
    .B1(_1914_),
    .X(_2569_));
 sg13g2_nand3_1 _7014_ (.B(_2098_),
    .C(_2121_),
    .A(_1962_),
    .Y(_2570_));
 sg13g2_nand2_1 _7015_ (.Y(_2571_),
    .A(net2234),
    .B(_1673_));
 sg13g2_o21ai_1 _7016_ (.B1(_1896_),
    .Y(_2572_),
    .A1(net2198),
    .A2(_1901_));
 sg13g2_a22oi_1 _7017_ (.Y(_2573_),
    .B1(_2572_),
    .B2(net1988),
    .A2(_2571_),
    .A1(_1976_));
 sg13g2_o21ai_1 _7018_ (.B1(_2570_),
    .Y(_2574_),
    .A1(net2185),
    .A2(_2573_));
 sg13g2_o21ai_1 _7019_ (.B1(_1746_),
    .Y(_2575_),
    .A1(net2297),
    .A2(net2285));
 sg13g2_a21oi_1 _7020_ (.A1(net1828),
    .A2(_1809_),
    .Y(_2576_),
    .B1(_1963_));
 sg13g2_o21ai_1 _7021_ (.B1(_2327_),
    .Y(_2577_),
    .A1(_1775_),
    .A2(_2545_));
 sg13g2_nand2_1 _7022_ (.Y(_2578_),
    .A(net1888),
    .B(_2577_));
 sg13g2_a21oi_1 _7023_ (.A1(net2209),
    .A2(_1792_),
    .Y(_2579_),
    .B1(net2192));
 sg13g2_a21oi_1 _7024_ (.A1(_1555_),
    .A2(_1871_),
    .Y(_2580_),
    .B1(_2579_));
 sg13g2_nor2b_2 _7025_ (.A(_1862_),
    .B_N(_2164_),
    .Y(_2581_));
 sg13g2_nand2_1 _7026_ (.Y(_2582_),
    .A(net2242),
    .B(_2538_));
 sg13g2_a21oi_1 _7027_ (.A1(_2581_),
    .A2(_2582_),
    .Y(_2583_),
    .B1(_2580_));
 sg13g2_nor2_1 _7028_ (.A(_2430_),
    .B(_2530_),
    .Y(_2584_));
 sg13g2_and3_1 _7029_ (.X(_2585_),
    .A(net1948),
    .B(_1849_),
    .C(_2208_));
 sg13g2_nor4_1 _7030_ (.A(net2186),
    .B(_2583_),
    .C(_2584_),
    .D(_2585_),
    .Y(_2586_));
 sg13g2_a22oi_1 _7031_ (.Y(_2587_),
    .B1(_2578_),
    .B2(_2586_),
    .A2(_2576_),
    .A1(_2575_));
 sg13g2_inv_1 _7032_ (.Y(_2588_),
    .A(_2587_));
 sg13g2_a22oi_1 _7033_ (.Y(_2589_),
    .B1(_2588_),
    .B2(_1615_),
    .A2(_2574_),
    .A1(_1860_));
 sg13g2_nor2_1 _7034_ (.A(net2091),
    .B(_2589_),
    .Y(_2590_));
 sg13g2_o21ai_1 _7035_ (.B1(net2214),
    .Y(_2591_),
    .A1(net2233),
    .A2(_1866_));
 sg13g2_o21ai_1 _7036_ (.B1(net2235),
    .Y(_2592_),
    .A1(net2260),
    .A2(_1867_));
 sg13g2_a21oi_1 _7037_ (.A1(net2260),
    .A2(net1822),
    .Y(_2593_),
    .B1(_2592_));
 sg13g2_nand2_1 _7038_ (.Y(_2594_),
    .A(_1715_),
    .B(net1858));
 sg13g2_a22oi_1 _7039_ (.Y(_2595_),
    .B1(_2594_),
    .B2(net1996),
    .A2(net1865),
    .A1(net1874));
 sg13g2_o21ai_1 _7040_ (.B1(_2595_),
    .Y(_2596_),
    .A1(_2591_),
    .A2(_2593_));
 sg13g2_and2_1 _7041_ (.A(net2194),
    .B(_2596_),
    .X(_2597_));
 sg13g2_nor2_1 _7042_ (.A(_1647_),
    .B(_2113_),
    .Y(_2598_));
 sg13g2_o21ai_1 _7043_ (.B1(net1865),
    .Y(_2599_),
    .A1(_1871_),
    .A2(_2598_));
 sg13g2_a21oi_1 _7044_ (.A1(net2110),
    .A2(net1830),
    .Y(_2600_),
    .B1(net2002));
 sg13g2_a21oi_1 _7045_ (.A1(_1649_),
    .A2(_1668_),
    .Y(_2601_),
    .B1(net1851));
 sg13g2_a22oi_1 _7046_ (.Y(_2602_),
    .B1(_2601_),
    .B2(_2114_),
    .A2(_2600_),
    .A1(_1786_));
 sg13g2_nand3_1 _7047_ (.B(_2599_),
    .C(_2602_),
    .A(_1869_),
    .Y(_2603_));
 sg13g2_a21oi_1 _7048_ (.A1(net2089),
    .A2(_2603_),
    .Y(_2604_),
    .B1(_2597_));
 sg13g2_o21ai_1 _7049_ (.B1(_2335_),
    .Y(_2605_),
    .A1(_1647_),
    .A2(_2113_));
 sg13g2_nor2_1 _7050_ (.A(_1763_),
    .B(_1813_),
    .Y(_2606_));
 sg13g2_o21ai_1 _7051_ (.B1(_1897_),
    .Y(_2607_),
    .A1(net2238),
    .A2(net1881));
 sg13g2_nor2_1 _7052_ (.A(net2213),
    .B(_1906_),
    .Y(_2608_));
 sg13g2_a21oi_1 _7053_ (.A1(net2212),
    .A2(net1858),
    .Y(_2609_),
    .B1(_2608_));
 sg13g2_a221oi_1 _7054_ (.B2(net1910),
    .C1(_2609_),
    .B1(_2606_),
    .A1(net1865),
    .Y(_2610_),
    .A2(_2605_));
 sg13g2_nand2_1 _7055_ (.Y(_2611_),
    .A(net1891),
    .B(net1836));
 sg13g2_o21ai_1 _7056_ (.B1(net1993),
    .Y(_2612_),
    .A1(net1922),
    .A2(net1820));
 sg13g2_nand3_1 _7057_ (.B(_2611_),
    .C(_2612_),
    .A(net1949),
    .Y(_2613_));
 sg13g2_o21ai_1 _7058_ (.B1(_2613_),
    .Y(_2614_),
    .A1(net2197),
    .A2(_2610_));
 sg13g2_a21oi_1 _7059_ (.A1(net1886),
    .A2(_2607_),
    .Y(_2615_),
    .B1(_2614_));
 sg13g2_a22oi_1 _7060_ (.Y(_2616_),
    .B1(_2615_),
    .B2(net1772),
    .A2(_2604_),
    .A1(_1860_));
 sg13g2_o21ai_1 _7061_ (.B1(_2506_),
    .Y(_2617_),
    .A1(net1980),
    .A2(_2616_));
 sg13g2_nand4_1 _7062_ (.B(_2535_),
    .C(_2557_),
    .A(_2492_),
    .Y(_2618_),
    .D(_2569_));
 sg13g2_nand3_1 _7063_ (.B(_2482_),
    .C(_2515_),
    .A(_1440_),
    .Y(_2619_));
 sg13g2_nor4_1 _7064_ (.A(_2590_),
    .B(_2617_),
    .C(_2618_),
    .D(_2619_),
    .Y(_2620_));
 sg13g2_nor2_1 _7065_ (.A(_2273_),
    .B(_2620_),
    .Y(_2621_));
 sg13g2_nand4_1 _7066_ (.B(_2030_),
    .C(_2448_),
    .A(\draw_game_inst.board_x[2] ),
    .Y(_2622_),
    .D(_2621_));
 sg13g2_a21oi_2 _7067_ (.B1(_1917_),
    .Y(_2623_),
    .A2(_2119_),
    .A1(_1575_));
 sg13g2_nor4_2 _7068_ (.A(net2222),
    .B(net1929),
    .C(net1916),
    .Y(_2624_),
    .D(_1927_));
 sg13g2_a21oi_1 _7069_ (.A1(net2254),
    .A2(net2006),
    .Y(_2625_),
    .B1(net1839));
 sg13g2_nor2_1 _7070_ (.A(net2067),
    .B(_2625_),
    .Y(_2626_));
 sg13g2_a221oi_1 _7071_ (.B2(_2626_),
    .C1(_1853_),
    .B1(net1885),
    .A1(net2067),
    .Y(_2627_),
    .A2(net2013));
 sg13g2_o21ai_1 _7072_ (.B1(net1938),
    .Y(_2628_),
    .A1(_2624_),
    .A2(_2627_));
 sg13g2_nand2_1 _7073_ (.Y(_2629_),
    .A(_2623_),
    .B(_2628_));
 sg13g2_o21ai_1 _7074_ (.B1(_1962_),
    .Y(_2630_),
    .A1(net1836),
    .A2(_2530_));
 sg13g2_nand2_1 _7075_ (.Y(_2631_),
    .A(net2206),
    .B(net1850));
 sg13g2_a221oi_1 _7076_ (.B2(_1986_),
    .C1(net2188),
    .B1(_2631_),
    .A1(net2221),
    .Y(_2632_),
    .A2(_2032_));
 sg13g2_nand3_1 _7077_ (.B(_1634_),
    .C(_2611_),
    .A(net1885),
    .Y(_2633_));
 sg13g2_nand3_1 _7078_ (.B(_2224_),
    .C(_2633_),
    .A(_4042_),
    .Y(_2634_));
 sg13g2_o21ai_1 _7079_ (.B1(_2630_),
    .Y(_2635_),
    .A1(_2632_),
    .A2(_2634_));
 sg13g2_nand2_1 _7080_ (.Y(_2636_),
    .A(_1860_),
    .B(_2635_));
 sg13g2_nand2_1 _7081_ (.Y(_2637_),
    .A(_1768_),
    .B(_2179_));
 sg13g2_a22oi_1 _7082_ (.Y(_2638_),
    .B1(net1856),
    .B2(_2637_),
    .A2(_1678_),
    .A1(net1894));
 sg13g2_nand2_1 _7083_ (.Y(_2639_),
    .A(net1995),
    .B(_1678_));
 sg13g2_or2_1 _7084_ (.X(_2640_),
    .B(_2638_),
    .A(net2218));
 sg13g2_o21ai_1 _7085_ (.B1(_2639_),
    .Y(_2641_),
    .A1(net1995),
    .A2(_1618_));
 sg13g2_a22oi_1 _7086_ (.Y(_2642_),
    .B1(_2641_),
    .B2(net2218),
    .A2(_2283_),
    .A1(net1998));
 sg13g2_a21oi_1 _7087_ (.A1(_2640_),
    .A2(_2642_),
    .Y(_2643_),
    .B1(net2200));
 sg13g2_nor2_1 _7088_ (.A(net1894),
    .B(_1744_),
    .Y(_2644_));
 sg13g2_nor3_1 _7089_ (.A(net1919),
    .B(net1995),
    .C(_2178_),
    .Y(_2645_));
 sg13g2_nor3_1 _7090_ (.A(net1990),
    .B(_2644_),
    .C(_2645_),
    .Y(_2646_));
 sg13g2_a21oi_1 _7091_ (.A1(_1734_),
    .A2(_1736_),
    .Y(_2647_),
    .B1(net1944));
 sg13g2_nor4_2 _7092_ (.A(net2186),
    .B(_2643_),
    .C(_2646_),
    .Y(_2648_),
    .D(_2647_));
 sg13g2_o21ai_1 _7093_ (.B1(_1631_),
    .Y(_2649_),
    .A1(net2299),
    .A2(_0096_));
 sg13g2_a21oi_1 _7094_ (.A1(net1915),
    .A2(_2179_),
    .Y(_2650_),
    .B1(net2265));
 sg13g2_nor2_1 _7095_ (.A(net2109),
    .B(_2649_),
    .Y(_2651_));
 sg13g2_nor3_1 _7096_ (.A(_1963_),
    .B(_2650_),
    .C(_2651_),
    .Y(_2652_));
 sg13g2_o21ai_1 _7097_ (.B1(net1772),
    .Y(_2653_),
    .A1(_2648_),
    .A2(_2652_));
 sg13g2_nand3_1 _7098_ (.B(_2636_),
    .C(_2653_),
    .A(_2629_),
    .Y(_2654_));
 sg13g2_nand2_1 _7099_ (.Y(_2655_),
    .A(net2179),
    .B(_2654_));
 sg13g2_nor2_1 _7100_ (.A(net1909),
    .B(_1853_),
    .Y(_2656_));
 sg13g2_nor2_1 _7101_ (.A(net2085),
    .B(_2656_),
    .Y(_2657_));
 sg13g2_o21ai_1 _7102_ (.B1(net1909),
    .Y(_2658_),
    .A1(_2119_),
    .A2(_2516_));
 sg13g2_o21ai_1 _7103_ (.B1(net1868),
    .Y(_2659_),
    .A1(_1665_),
    .A2(_1982_));
 sg13g2_a221oi_1 _7104_ (.B2(net2207),
    .C1(net2187),
    .B1(net1819),
    .A1(_1570_),
    .Y(_2660_),
    .A2(net1996));
 sg13g2_a22oi_1 _7105_ (.Y(_2661_),
    .B1(_2659_),
    .B2(_2660_),
    .A2(_2658_),
    .A1(_2657_));
 sg13g2_nor3_1 _7106_ (.A(net2182),
    .B(_2629_),
    .C(_2661_),
    .Y(_2662_));
 sg13g2_o21ai_1 _7107_ (.B1(_2195_),
    .Y(_2663_),
    .A1(net1904),
    .A2(_2626_));
 sg13g2_nand2_1 _7108_ (.Y(_2664_),
    .A(net1819),
    .B(_2663_));
 sg13g2_o21ai_1 _7109_ (.B1(net2188),
    .Y(_2665_),
    .A1(_1582_),
    .A2(_1982_));
 sg13g2_o21ai_1 _7110_ (.B1(_2664_),
    .Y(_2666_),
    .A1(_1582_),
    .A2(_2665_));
 sg13g2_a21oi_1 _7111_ (.A1(_1558_),
    .A2(_2665_),
    .Y(_2667_),
    .B1(net1834));
 sg13g2_o21ai_1 _7112_ (.B1(net1938),
    .Y(_2668_),
    .A1(_2666_),
    .A2(_2667_));
 sg13g2_o21ai_1 _7113_ (.B1(_1575_),
    .Y(_2669_),
    .A1(_1558_),
    .A2(net1832));
 sg13g2_a21oi_1 _7114_ (.A1(net2222),
    .A2(net2006),
    .Y(_2670_),
    .B1(net1904));
 sg13g2_o21ai_1 _7115_ (.B1(_2670_),
    .Y(_2671_),
    .A1(net2221),
    .A2(net1832));
 sg13g2_a21oi_1 _7116_ (.A1(net1885),
    .A2(net1832),
    .Y(_2672_),
    .B1(net2182));
 sg13g2_a22oi_1 _7117_ (.Y(_2673_),
    .B1(_1634_),
    .B2(net2013),
    .A2(net2004),
    .A1(net1949));
 sg13g2_nand3_1 _7118_ (.B(_2672_),
    .C(_2673_),
    .A(_2671_),
    .Y(_2674_));
 sg13g2_nand2_1 _7119_ (.Y(_2675_),
    .A(net2091),
    .B(_2674_));
 sg13g2_nand4_1 _7120_ (.B(_2668_),
    .C(_2669_),
    .A(_1829_),
    .Y(_2676_),
    .D(_2675_));
 sg13g2_o21ai_1 _7121_ (.B1(net2257),
    .Y(_2677_),
    .A1(_1788_),
    .A2(_1864_));
 sg13g2_nand3_1 _7122_ (.B(_1668_),
    .C(_2677_),
    .A(net2226),
    .Y(_2678_));
 sg13g2_nand4_1 _7123_ (.B(net2014),
    .C(_1639_),
    .A(net2290),
    .Y(_2679_),
    .D(_2678_));
 sg13g2_and2_2 _7124_ (.A(_1689_),
    .B(_1787_),
    .X(_2680_));
 sg13g2_nand2_1 _7125_ (.Y(_2681_),
    .A(_1689_),
    .B(_1787_));
 sg13g2_o21ai_1 _7126_ (.B1(_2680_),
    .Y(_2682_),
    .A1(_2305_),
    .A2(_2414_));
 sg13g2_o21ai_1 _7127_ (.B1(net1875),
    .Y(_2683_),
    .A1(net1991),
    .A2(net1835));
 sg13g2_a22oi_1 _7128_ (.Y(_2684_),
    .B1(_2683_),
    .B2(net1906),
    .A2(_1657_),
    .A1(net1882));
 sg13g2_nand3_1 _7129_ (.B(_2682_),
    .C(_2684_),
    .A(_2679_),
    .Y(_2685_));
 sg13g2_o21ai_1 _7130_ (.B1(net1948),
    .Y(_2686_),
    .A1(net1925),
    .A2(net1835));
 sg13g2_nand2_1 _7131_ (.Y(_2687_),
    .A(_1461_),
    .B(_2114_));
 sg13g2_o21ai_1 _7132_ (.B1(_1736_),
    .Y(_2688_),
    .A1(net1854),
    .A2(_2687_));
 sg13g2_o21ai_1 _7133_ (.B1(net1888),
    .Y(_2689_),
    .A1(_2483_),
    .A2(_2688_));
 sg13g2_nor2_2 _7134_ (.A(net1878),
    .B(_2677_),
    .Y(_2690_));
 sg13g2_a21oi_1 _7135_ (.A1(_1812_),
    .A2(_2554_),
    .Y(_2691_),
    .B1(_2690_));
 sg13g2_nor2_1 _7136_ (.A(net2256),
    .B(_2045_),
    .Y(_2692_));
 sg13g2_o21ai_1 _7137_ (.B1(net2225),
    .Y(_2693_),
    .A1(_1648_),
    .A2(_2692_));
 sg13g2_a21oi_1 _7138_ (.A1(net1861),
    .A2(_2693_),
    .Y(_2694_),
    .B1(_1761_));
 sg13g2_o21ai_1 _7139_ (.B1(_2686_),
    .Y(_2695_),
    .A1(_1556_),
    .A2(_2691_));
 sg13g2_nor2_1 _7140_ (.A(_2694_),
    .B(_2695_),
    .Y(_2696_));
 sg13g2_a22oi_1 _7141_ (.Y(_2697_),
    .B1(_2689_),
    .B2(_2696_),
    .A2(_2685_),
    .A1(net1937));
 sg13g2_o21ai_1 _7142_ (.B1(net1756),
    .Y(_2698_),
    .A1(_1782_),
    .A2(_2697_));
 sg13g2_nand2b_1 _7143_ (.Y(_2699_),
    .B(_2676_),
    .A_N(_2698_));
 sg13g2_nor2_1 _7144_ (.A(net1878),
    .B(_2680_),
    .Y(_2700_));
 sg13g2_a221oi_1 _7145_ (.B2(_2700_),
    .C1(net2203),
    .B1(net1857),
    .A1(net1895),
    .Y(_2701_),
    .A2(net1880));
 sg13g2_o21ai_1 _7146_ (.B1(net2074),
    .Y(_2702_),
    .A1(_2231_),
    .A2(_2690_));
 sg13g2_a21oi_1 _7147_ (.A1(_2701_),
    .A2(_2702_),
    .Y(_2703_),
    .B1(net2199));
 sg13g2_a21oi_1 _7148_ (.A1(net2240),
    .A2(_2283_),
    .Y(_2704_),
    .B1(_1625_));
 sg13g2_nor2_2 _7149_ (.A(net2266),
    .B(net2022),
    .Y(_2705_));
 sg13g2_nand3_1 _7150_ (.B(net1915),
    .C(_2705_),
    .A(net2074),
    .Y(_2706_));
 sg13g2_a22oi_1 _7151_ (.Y(_2707_),
    .B1(net1848),
    .B2(_2198_),
    .A2(_0096_),
    .A1(net2230));
 sg13g2_a21oi_1 _7152_ (.A1(_2706_),
    .A2(_2707_),
    .Y(_2708_),
    .B1(net1990));
 sg13g2_o21ai_1 _7153_ (.B1(net1983),
    .Y(_2709_),
    .A1(net1944),
    .A2(_2704_));
 sg13g2_nor3_1 _7154_ (.A(_2703_),
    .B(_2708_),
    .C(_2709_),
    .Y(_2710_));
 sg13g2_o21ai_1 _7155_ (.B1(net2191),
    .Y(_2711_),
    .A1(net2081),
    .A2(_1791_));
 sg13g2_o21ai_1 _7156_ (.B1(net2227),
    .Y(_2712_),
    .A1(net2256),
    .A2(_1436_));
 sg13g2_nor3_1 _7157_ (.A(net2220),
    .B(_2690_),
    .C(_2712_),
    .Y(_2713_));
 sg13g2_o21ai_1 _7158_ (.B1(_1764_),
    .Y(_2714_),
    .A1(net2105),
    .A2(_1692_));
 sg13g2_nor2_1 _7159_ (.A(_1582_),
    .B(_2714_),
    .Y(_2715_));
 sg13g2_nor3_1 _7160_ (.A(_2711_),
    .B(_2713_),
    .C(_2715_),
    .Y(_2716_));
 sg13g2_nor3_1 _7161_ (.A(net2001),
    .B(_1735_),
    .C(_1944_),
    .Y(_2717_));
 sg13g2_nor2_1 _7162_ (.A(_2387_),
    .B(_2717_),
    .Y(_2718_));
 sg13g2_nor2_2 _7163_ (.A(net2084),
    .B(_1944_),
    .Y(_2719_));
 sg13g2_o21ai_1 _7164_ (.B1(net2217),
    .Y(_2720_),
    .A1(net2075),
    .A2(net1903));
 sg13g2_nor3_1 _7165_ (.A(net2001),
    .B(_1735_),
    .C(_2720_),
    .Y(_2721_));
 sg13g2_nor3_2 _7166_ (.A(net2200),
    .B(_2718_),
    .C(_2721_),
    .Y(_2722_));
 sg13g2_nor3_1 _7167_ (.A(net1936),
    .B(_2716_),
    .C(_2722_),
    .Y(_2723_));
 sg13g2_o21ai_1 _7168_ (.B1(_1981_),
    .Y(_2724_),
    .A1(_2710_),
    .A2(_2723_));
 sg13g2_a21oi_2 _7169_ (.B1(net1995),
    .Y(_2725_),
    .A2(_2179_),
    .A1(_1768_));
 sg13g2_a21oi_1 _7170_ (.A1(net2247),
    .A2(_2705_),
    .Y(_2726_),
    .B1(_2725_));
 sg13g2_a21oi_1 _7171_ (.A1(net1893),
    .A2(_1770_),
    .Y(_2727_),
    .B1(net2084));
 sg13g2_a221oi_1 _7172_ (.B2(_2639_),
    .C1(net2200),
    .B1(_2727_),
    .A1(_2581_),
    .Y(_2728_),
    .A2(_2726_));
 sg13g2_o21ai_1 _7173_ (.B1(net2244),
    .Y(_2729_),
    .A1(net2107),
    .A2(_1743_));
 sg13g2_a21oi_1 _7174_ (.A1(_1443_),
    .A2(_1763_),
    .Y(_2730_),
    .B1(_2729_));
 sg13g2_o21ai_1 _7175_ (.B1(net2075),
    .Y(_2731_),
    .A1(net2267),
    .A2(_2113_));
 sg13g2_a21oi_1 _7176_ (.A1(net1901),
    .A2(_1813_),
    .Y(_2732_),
    .B1(_2731_));
 sg13g2_nor3_1 _7177_ (.A(net1990),
    .B(_2730_),
    .C(_2732_),
    .Y(_2733_));
 sg13g2_a221oi_1 _7178_ (.B2(net2076),
    .C1(net1945),
    .B1(_1737_),
    .A1(net2064),
    .Y(_2734_),
    .A2(net1871));
 sg13g2_nor4_1 _7179_ (.A(net1981),
    .B(_2728_),
    .C(_2733_),
    .D(_2734_),
    .Y(_2735_));
 sg13g2_a21oi_1 _7180_ (.A1(net2267),
    .A2(net2298),
    .Y(_2736_),
    .B1(_1443_));
 sg13g2_o21ai_1 _7181_ (.B1(net2218),
    .Y(_2737_),
    .A1(net2243),
    .A2(net1903));
 sg13g2_o21ai_1 _7182_ (.B1(net2244),
    .Y(_2738_),
    .A1(_1685_),
    .A2(_1813_));
 sg13g2_nand2b_1 _7183_ (.Y(_2739_),
    .B(_2738_),
    .A_N(_2737_));
 sg13g2_o21ai_1 _7184_ (.B1(_2386_),
    .Y(_2740_),
    .A1(net2243),
    .A2(_2210_));
 sg13g2_nand3_1 _7185_ (.B(_2739_),
    .C(_2740_),
    .A(net2200),
    .Y(_2741_));
 sg13g2_a221oi_1 _7186_ (.B2(net2267),
    .C1(net2002),
    .B1(_2210_),
    .A1(net2030),
    .Y(_2742_),
    .A2(_1665_));
 sg13g2_o21ai_1 _7187_ (.B1(net1852),
    .Y(_2743_),
    .A1(_1750_),
    .A2(_2143_));
 sg13g2_o21ai_1 _7188_ (.B1(_2743_),
    .Y(_2744_),
    .A1(net2217),
    .A2(_1743_));
 sg13g2_o21ai_1 _7189_ (.B1(net2088),
    .Y(_2745_),
    .A1(_2742_),
    .A2(_2744_));
 sg13g2_nand2_1 _7190_ (.Y(_2746_),
    .A(_2741_),
    .B(_2745_));
 sg13g2_inv_1 _7191_ (.Y(_2747_),
    .A(_2746_));
 sg13g2_a221oi_1 _7192_ (.B2(net1940),
    .C1(_2735_),
    .B1(_2747_),
    .A1(net1817),
    .Y(_2748_),
    .A2(_2736_));
 sg13g2_o21ai_1 _7193_ (.B1(_2724_),
    .Y(_2749_),
    .A1(_1936_),
    .A2(_2748_));
 sg13g2_nor3_1 _7194_ (.A(net2074),
    .B(net1838),
    .C(_2034_),
    .Y(_2750_));
 sg13g2_a21oi_1 _7195_ (.A1(net1856),
    .A2(_2018_),
    .Y(_2751_),
    .B1(_2750_));
 sg13g2_nand3_1 _7196_ (.B(_2245_),
    .C(_2751_),
    .A(_1428_),
    .Y(_2752_));
 sg13g2_a22oi_1 _7197_ (.Y(_2753_),
    .B1(net1848),
    .B2(_2184_),
    .A2(_1854_),
    .A1(net2010));
 sg13g2_nand3b_1 _7198_ (.B(_2753_),
    .C(net1908),
    .Y(_2754_),
    .A_N(_2240_));
 sg13g2_a21oi_1 _7199_ (.A1(net2246),
    .A2(net2287),
    .Y(_2755_),
    .B1(_1460_));
 sg13g2_nand3_1 _7200_ (.B(net1818),
    .C(_2637_),
    .A(net2247),
    .Y(_2756_));
 sg13g2_o21ai_1 _7201_ (.B1(_2164_),
    .Y(_2757_),
    .A1(net2247),
    .A2(net1881));
 sg13g2_nor2_1 _7202_ (.A(net2200),
    .B(_2757_),
    .Y(_2758_));
 sg13g2_a22oi_1 _7203_ (.Y(_2759_),
    .B1(_2756_),
    .B2(_2758_),
    .A2(_2755_),
    .A1(net1888));
 sg13g2_nand3_1 _7204_ (.B(_2754_),
    .C(_2759_),
    .A(_2752_),
    .Y(_2760_));
 sg13g2_o21ai_1 _7205_ (.B1(net1998),
    .Y(_2761_),
    .A1(net2252),
    .A2(net1835));
 sg13g2_and2_1 _7206_ (.A(_2111_),
    .B(_2761_),
    .X(_2762_));
 sg13g2_a21oi_1 _7207_ (.A1(_2591_),
    .A2(_2762_),
    .Y(_2763_),
    .B1(net2194));
 sg13g2_nand3b_1 _7208_ (.B(_2762_),
    .C(_2034_),
    .Y(_2764_),
    .A_N(_2592_));
 sg13g2_nor2_1 _7209_ (.A(net1943),
    .B(_2055_),
    .Y(_2765_));
 sg13g2_o21ai_1 _7210_ (.B1(net1813),
    .Y(_2766_),
    .A1(_1822_),
    .A2(_2262_));
 sg13g2_nor2_1 _7211_ (.A(net1987),
    .B(_1818_),
    .Y(_2767_));
 sg13g2_a221oi_1 _7212_ (.B2(_2767_),
    .C1(_2765_),
    .B1(_2766_),
    .A1(_2763_),
    .Y(_2768_),
    .A2(_2764_));
 sg13g2_a22oi_1 _7213_ (.Y(_2769_),
    .B1(_2768_),
    .B2(_1860_),
    .A2(_2760_),
    .A1(net1772));
 sg13g2_nand2b_1 _7214_ (.Y(_2770_),
    .B(net1983),
    .A_N(_2769_));
 sg13g2_nand3_1 _7215_ (.B(_1657_),
    .C(_1853_),
    .A(net1924),
    .Y(_2771_));
 sg13g2_and2_1 _7216_ (.A(net2013),
    .B(_1594_),
    .X(_2772_));
 sg13g2_a22oi_1 _7217_ (.Y(_2773_),
    .B1(_2772_),
    .B2(_1632_),
    .A2(_1890_),
    .A1(_1457_));
 sg13g2_a21oi_1 _7218_ (.A1(_2771_),
    .A2(_2773_),
    .Y(_2774_),
    .B1(net1933));
 sg13g2_o21ai_1 _7219_ (.B1(_2034_),
    .Y(_2775_),
    .A1(net2253),
    .A2(net1831));
 sg13g2_nand3_1 _7220_ (.B(_1856_),
    .C(_2631_),
    .A(net2003),
    .Y(_2776_));
 sg13g2_a221oi_1 _7221_ (.B2(net2221),
    .C1(_2776_),
    .B1(_2775_),
    .A1(net1997),
    .Y(_2777_),
    .A2(_1744_));
 sg13g2_o21ai_1 _7222_ (.B1(net1771),
    .Y(_2778_),
    .A1(_2774_),
    .A2(_2777_));
 sg13g2_nand2b_1 _7223_ (.Y(_2779_),
    .B(net2225),
    .A_N(_2389_));
 sg13g2_a21oi_1 _7224_ (.A1(_2080_),
    .A2(_2779_),
    .Y(_2780_),
    .B1(net1942));
 sg13g2_nor2_1 _7225_ (.A(_1809_),
    .B(_2119_),
    .Y(_2781_));
 sg13g2_o21ai_1 _7226_ (.B1(net2014),
    .Y(_2782_),
    .A1(_1811_),
    .A2(_2119_));
 sg13g2_o21ai_1 _7227_ (.B1(net2000),
    .Y(_2783_),
    .A1(net2017),
    .A2(net1922));
 sg13g2_a221oi_1 _7228_ (.B2(_2783_),
    .C1(net1934),
    .B1(net1884),
    .A1(_1548_),
    .Y(_2784_),
    .A2(net1906));
 sg13g2_o21ai_1 _7229_ (.B1(_2784_),
    .Y(_2785_),
    .A1(_2104_),
    .A2(_2782_));
 sg13g2_nand3_1 _7230_ (.B(_1771_),
    .C(_1919_),
    .A(net2073),
    .Y(_2786_));
 sg13g2_nand3_1 _7231_ (.B(_1852_),
    .C(_2786_),
    .A(net2083),
    .Y(_2787_));
 sg13g2_a221oi_1 _7232_ (.B2(net2106),
    .C1(net2079),
    .B1(_1818_),
    .A1(_1436_),
    .Y(_2788_),
    .A2(net1924));
 sg13g2_nor2_1 _7233_ (.A(net1863),
    .B(_2788_),
    .Y(_2789_));
 sg13g2_and2_1 _7234_ (.A(_2787_),
    .B(_2789_),
    .X(_2790_));
 sg13g2_o21ai_1 _7235_ (.B1(_1993_),
    .Y(_2791_),
    .A1(net2225),
    .A2(_2045_));
 sg13g2_nor2_1 _7236_ (.A(_2152_),
    .B(_2791_),
    .Y(_2792_));
 sg13g2_o21ai_1 _7237_ (.B1(_2792_),
    .Y(_2793_),
    .A1(net1854),
    .A2(_2680_));
 sg13g2_o21ai_1 _7238_ (.B1(_2793_),
    .Y(_2794_),
    .A1(_2780_),
    .A2(_2785_));
 sg13g2_o21ai_1 _7239_ (.B1(net1770),
    .Y(_2795_),
    .A1(_2790_),
    .A2(_2794_));
 sg13g2_nand3_1 _7240_ (.B(_1657_),
    .C(_2017_),
    .A(_1554_),
    .Y(_2796_));
 sg13g2_o21ai_1 _7241_ (.B1(net1930),
    .Y(_2797_),
    .A1(_1556_),
    .A2(net1869));
 sg13g2_a21o_1 _7242_ (.A2(_1816_),
    .A1(net1831),
    .B1(_2055_),
    .X(_2798_));
 sg13g2_o21ai_1 _7243_ (.B1(_2797_),
    .Y(_2799_),
    .A1(net2206),
    .A2(_2798_));
 sg13g2_a21oi_1 _7244_ (.A1(_2796_),
    .A2(_2799_),
    .Y(_2800_),
    .B1(net1932));
 sg13g2_a221oi_1 _7245_ (.B2(net2068),
    .C1(net2206),
    .B1(_2017_),
    .A1(_1632_),
    .Y(_2801_),
    .A2(_1816_));
 sg13g2_nor2_1 _7246_ (.A(net2080),
    .B(_2329_),
    .Y(_2802_));
 sg13g2_nor3_1 _7247_ (.A(_1857_),
    .B(_2801_),
    .C(_2802_),
    .Y(_2803_));
 sg13g2_o21ai_1 _7248_ (.B1(_1702_),
    .Y(_2804_),
    .A1(_2800_),
    .A2(_2803_));
 sg13g2_nand4_1 _7249_ (.B(_2778_),
    .C(_2795_),
    .A(_2770_),
    .Y(_2805_),
    .D(_2804_));
 sg13g2_nor4_1 _7250_ (.A(_2662_),
    .B(_2699_),
    .C(_2749_),
    .D(_2805_),
    .Y(_2806_));
 sg13g2_nand3_1 _7251_ (.B(net1880),
    .C(_1961_),
    .A(_1577_),
    .Y(_2807_));
 sg13g2_and2_1 _7252_ (.A(net1932),
    .B(_2807_),
    .X(_2808_));
 sg13g2_nand2_2 _7253_ (.Y(_2809_),
    .A(net2205),
    .B(_1930_));
 sg13g2_nor2_1 _7254_ (.A(_2626_),
    .B(_2809_),
    .Y(_2810_));
 sg13g2_nor2_1 _7255_ (.A(net2085),
    .B(_2810_),
    .Y(_2811_));
 sg13g2_nand2_1 _7256_ (.Y(_2812_),
    .A(net2079),
    .B(_1548_));
 sg13g2_a22oi_1 _7257_ (.Y(_2813_),
    .B1(_2811_),
    .B2(_2812_),
    .A2(_2277_),
    .A1(_1986_));
 sg13g2_a21oi_1 _7258_ (.A1(_4042_),
    .A2(_2813_),
    .Y(_2814_),
    .B1(_2808_));
 sg13g2_nand3b_1 _7259_ (.B(net2232),
    .C(_2394_),
    .Y(_2815_),
    .A_N(_2516_));
 sg13g2_a21oi_1 _7260_ (.A1(net2067),
    .A2(_1853_),
    .Y(_2816_),
    .B1(net1943));
 sg13g2_nand2_1 _7261_ (.Y(_2817_),
    .A(net2091),
    .B(_2672_));
 sg13g2_a221oi_1 _7262_ (.B2(_2816_),
    .C1(_2817_),
    .B1(_2815_),
    .A1(net1905),
    .Y(_2818_),
    .A2(net1819));
 sg13g2_and2_1 _7263_ (.A(net2013),
    .B(_1952_),
    .X(_2819_));
 sg13g2_o21ai_1 _7264_ (.B1(_2819_),
    .Y(_2820_),
    .A1(net2250),
    .A2(_1548_));
 sg13g2_a21oi_1 _7265_ (.A1(_2818_),
    .A2(_2820_),
    .Y(_2821_),
    .B1(_2814_));
 sg13g2_a221oi_1 _7266_ (.B2(_1538_),
    .C1(\draw_game_inst.board_x[0] ),
    .B1(_2821_),
    .A1(_2655_),
    .Y(_2822_),
    .A2(_2806_));
 sg13g2_nand3_1 _7267_ (.B(net1997),
    .C(_1639_),
    .A(net2294),
    .Y(_2823_));
 sg13g2_and4_1 _7268_ (.A(net1865),
    .B(net1825),
    .C(_1708_),
    .D(net1818),
    .X(_2824_));
 sg13g2_o21ai_1 _7269_ (.B1(_2823_),
    .Y(_2825_),
    .A1(net2080),
    .A2(_1822_));
 sg13g2_a22oi_1 _7270_ (.Y(_2826_),
    .B1(_1882_),
    .B2(net2260),
    .A2(_1809_),
    .A1(net1827));
 sg13g2_nand2b_1 _7271_ (.Y(_2827_),
    .B(net1852),
    .A_N(_2826_));
 sg13g2_o21ai_1 _7272_ (.B1(_2827_),
    .Y(_2828_),
    .A1(_2824_),
    .A2(_2825_));
 sg13g2_o21ai_1 _7273_ (.B1(_2796_),
    .Y(_2829_),
    .A1(net2187),
    .A2(_2828_));
 sg13g2_a21oi_1 _7274_ (.A1(net2010),
    .A2(net1830),
    .Y(_2830_),
    .B1(_1755_));
 sg13g2_a22oi_1 _7275_ (.Y(_2831_),
    .B1(_2700_),
    .B2(net2264),
    .A2(_2031_),
    .A1(net1829));
 sg13g2_nor3_1 _7276_ (.A(net2216),
    .B(net2063),
    .C(_1820_),
    .Y(_2832_));
 sg13g2_nor4_1 _7277_ (.A(net2199),
    .B(_1970_),
    .C(_2261_),
    .D(_2832_),
    .Y(_2833_));
 sg13g2_o21ai_1 _7278_ (.B1(_2833_),
    .Y(_2834_),
    .A1(net1851),
    .A2(_2831_));
 sg13g2_o21ai_1 _7279_ (.B1(_2834_),
    .Y(_2835_),
    .A1(net1824),
    .A2(_2830_));
 sg13g2_a22oi_1 _7280_ (.Y(_2836_),
    .B1(_2835_),
    .B2(net1771),
    .A2(_2829_),
    .A1(_1702_));
 sg13g2_a22oi_1 _7281_ (.Y(_2837_),
    .B1(_2179_),
    .B2(net1818),
    .A2(_2069_),
    .A1(net1854));
 sg13g2_o21ai_1 _7282_ (.B1(_2706_),
    .Y(_2838_),
    .A1(net1995),
    .A2(_1692_));
 sg13g2_o21ai_1 _7283_ (.B1(net1888),
    .Y(_2839_),
    .A1(_2837_),
    .A2(_2838_));
 sg13g2_nand2_1 _7284_ (.Y(_2840_),
    .A(_1741_),
    .B(net1818));
 sg13g2_o21ai_1 _7285_ (.B1(_1555_),
    .Y(_2841_),
    .A1(_1737_),
    .A2(_2840_));
 sg13g2_nand3_1 _7286_ (.B(_1681_),
    .C(_2179_),
    .A(net2010),
    .Y(_2842_));
 sg13g2_a21oi_1 _7287_ (.A1(net2022),
    .A2(net1927),
    .Y(_2843_),
    .B1(net1944));
 sg13g2_a21o_1 _7288_ (.A2(_0096_),
    .A1(net2241),
    .B1(net2204),
    .X(_2844_));
 sg13g2_a22oi_1 _7289_ (.Y(_2845_),
    .B1(_2844_),
    .B2(net2088),
    .A2(_2843_),
    .A1(_2842_));
 sg13g2_nand4_1 _7290_ (.B(_2839_),
    .C(_2841_),
    .A(_1981_),
    .Y(_2846_),
    .D(_2845_));
 sg13g2_nand2_2 _7291_ (.Y(_2847_),
    .A(net2264),
    .B(net2295));
 sg13g2_o21ai_1 _7292_ (.B1(_2847_),
    .Y(_2848_),
    .A1(net2254),
    .A2(_2017_));
 sg13g2_o21ai_1 _7293_ (.B1(net2206),
    .Y(_2849_),
    .A1(net2009),
    .A2(net1874));
 sg13g2_a21oi_1 _7294_ (.A1(net2009),
    .A2(net1834),
    .Y(_2850_),
    .B1(_2849_));
 sg13g2_a21oi_1 _7295_ (.A1(net1832),
    .A2(net1868),
    .Y(_2851_),
    .B1(_0091_));
 sg13g2_a21oi_1 _7296_ (.A1(net1997),
    .A2(_2848_),
    .Y(_2852_),
    .B1(_2850_));
 sg13g2_nand3_1 _7297_ (.B(_2851_),
    .C(_2852_),
    .A(_1702_),
    .Y(_2853_));
 sg13g2_a21oi_1 _7298_ (.A1(_2846_),
    .A2(_2853_),
    .Y(_2854_),
    .B1(net1981));
 sg13g2_nor3_1 _7299_ (.A(net2187),
    .B(_1675_),
    .C(_1921_),
    .Y(_2855_));
 sg13g2_nor2_1 _7300_ (.A(net2003),
    .B(_2560_),
    .Y(_2856_));
 sg13g2_o21ai_1 _7301_ (.B1(net2187),
    .Y(_2857_),
    .A1(_2656_),
    .A2(_2856_));
 sg13g2_a21oi_1 _7302_ (.A1(net1905),
    .A2(net1819),
    .Y(_2858_),
    .B1(net2182));
 sg13g2_nand3b_1 _7303_ (.B(_2857_),
    .C(_2858_),
    .Y(_2859_),
    .A_N(_2855_));
 sg13g2_nor3_1 _7304_ (.A(net1916),
    .B(_1884_),
    .C(_1919_),
    .Y(_2860_));
 sg13g2_nand2_1 _7305_ (.Y(_2861_),
    .A(net1949),
    .B(net1832));
 sg13g2_nand2_2 _7306_ (.Y(_2862_),
    .A(net1994),
    .B(net1887));
 sg13g2_o21ai_1 _7307_ (.B1(_2861_),
    .Y(_2863_),
    .A1(_1853_),
    .A2(_2862_));
 sg13g2_nor3_1 _7308_ (.A(_2624_),
    .B(_2860_),
    .C(_2863_),
    .Y(_2864_));
 sg13g2_nand2_1 _7309_ (.Y(_2865_),
    .A(_1686_),
    .B(_2147_));
 sg13g2_nand2_1 _7310_ (.Y(_2866_),
    .A(net2222),
    .B(_2865_));
 sg13g2_o21ai_1 _7311_ (.B1(_1792_),
    .Y(_2867_),
    .A1(net1924),
    .A2(_1853_));
 sg13g2_a22oi_1 _7312_ (.Y(_2868_),
    .B1(_2867_),
    .B2(net1905),
    .A2(_2865_),
    .A1(_2194_));
 sg13g2_a21oi_1 _7313_ (.A1(_2864_),
    .A2(_2868_),
    .Y(_2869_),
    .B1(net1932));
 sg13g2_a21oi_1 _7314_ (.A1(net2091),
    .A2(_2859_),
    .Y(_2870_),
    .B1(_2869_));
 sg13g2_nand2_1 _7315_ (.Y(_2871_),
    .A(net2253),
    .B(_2047_));
 sg13g2_o21ai_1 _7316_ (.B1(_2045_),
    .Y(_2872_),
    .A1(net2104),
    .A2(net1880));
 sg13g2_a21oi_1 _7317_ (.A1(net2224),
    .A2(_2872_),
    .Y(_2873_),
    .B1(net2203));
 sg13g2_or2_1 _7318_ (.X(_2874_),
    .B(_2873_),
    .A(net2192));
 sg13g2_nand3_1 _7319_ (.B(_1786_),
    .C(_1790_),
    .A(_1555_),
    .Y(_2875_));
 sg13g2_o21ai_1 _7320_ (.B1(net1948),
    .Y(_2876_),
    .A1(net1914),
    .A2(net1854));
 sg13g2_a21oi_1 _7321_ (.A1(net1854),
    .A2(_2046_),
    .Y(_2877_),
    .B1(_2876_));
 sg13g2_o21ai_1 _7322_ (.B1(_2875_),
    .Y(_2878_),
    .A1(net1986),
    .A2(_2484_));
 sg13g2_nor3_1 _7323_ (.A(net1980),
    .B(_2877_),
    .C(_2878_),
    .Y(_2879_));
 sg13g2_nor3_1 _7324_ (.A(net1925),
    .B(_1788_),
    .C(_1864_),
    .Y(_2880_));
 sg13g2_o21ai_1 _7325_ (.B1(net1937),
    .Y(_2881_),
    .A1(net1986),
    .A2(_2880_));
 sg13g2_a21oi_1 _7326_ (.A1(net1906),
    .A2(_2105_),
    .Y(_2882_),
    .B1(_2881_));
 sg13g2_nand2_1 _7327_ (.Y(_2883_),
    .A(net1947),
    .B(_2678_));
 sg13g2_a21oi_1 _7328_ (.A1(net2065),
    .A2(_1716_),
    .Y(_2884_),
    .B1(_2883_));
 sg13g2_a22oi_1 _7329_ (.Y(_2885_),
    .B1(_1812_),
    .B2(_1862_),
    .A2(net1823),
    .A1(net2223));
 sg13g2_nor2_1 _7330_ (.A(net1930),
    .B(_2885_),
    .Y(_2886_));
 sg13g2_nor2_1 _7331_ (.A(_2884_),
    .B(_2886_),
    .Y(_2887_));
 sg13g2_a22oi_1 _7332_ (.Y(_2888_),
    .B1(_2882_),
    .B2(_2887_),
    .A2(_2879_),
    .A1(_2874_));
 sg13g2_o21ai_1 _7333_ (.B1(net2229),
    .Y(_2889_),
    .A1(_2192_),
    .A2(_2690_));
 sg13g2_nor2_1 _7334_ (.A(net2209),
    .B(_1728_),
    .Y(_2890_));
 sg13g2_a21oi_1 _7335_ (.A1(_2889_),
    .A2(_2890_),
    .Y(_2891_),
    .B1(_2711_));
 sg13g2_nand3_1 _7336_ (.B(_1729_),
    .C(_2889_),
    .A(net1883),
    .Y(_2892_));
 sg13g2_a22oi_1 _7337_ (.Y(_2893_),
    .B1(_1736_),
    .B2(_2719_),
    .A2(net1998),
    .A1(net2017));
 sg13g2_a21oi_1 _7338_ (.A1(net2087),
    .A2(_2893_),
    .Y(_2894_),
    .B1(_2891_));
 sg13g2_nand4_1 _7339_ (.B(_1981_),
    .C(_2892_),
    .A(net1937),
    .Y(_2895_),
    .D(_2894_));
 sg13g2_o21ai_1 _7340_ (.B1(_2895_),
    .Y(_2896_),
    .A1(_1782_),
    .A2(_2888_));
 sg13g2_nand2_1 _7341_ (.Y(_2897_),
    .A(_1745_),
    .B(_2847_));
 sg13g2_o21ai_1 _7342_ (.B1(net2084),
    .Y(_2898_),
    .A1(net2073),
    .A2(_1789_));
 sg13g2_nor2_2 _7343_ (.A(net2084),
    .B(net2011),
    .Y(_2899_));
 sg13g2_a22oi_1 _7344_ (.Y(_2900_),
    .B1(_2899_),
    .B2(_2113_),
    .A2(_2165_),
    .A1(_1789_));
 sg13g2_a221oi_1 _7345_ (.B2(_2900_),
    .C1(_1858_),
    .B1(_2898_),
    .A1(net1999),
    .Y(_2901_),
    .A2(_2897_));
 sg13g2_a221oi_1 _7346_ (.B2(net1818),
    .C1(_2757_),
    .B1(_2725_),
    .A1(net1856),
    .Y(_2902_),
    .A2(_2110_));
 sg13g2_a22oi_1 _7347_ (.Y(_2903_),
    .B1(_2720_),
    .B2(net2088),
    .A2(_1744_),
    .A1(_1555_));
 sg13g2_nor2_1 _7348_ (.A(_2902_),
    .B(_2903_),
    .Y(_2904_));
 sg13g2_o21ai_1 _7349_ (.B1(net1889),
    .Y(_2905_),
    .A1(net1900),
    .A2(net1894));
 sg13g2_a21oi_2 _7350_ (.B1(net1901),
    .Y(_2906_),
    .A2(net1894),
    .A1(net2062));
 sg13g2_o21ai_1 _7351_ (.B1(_2905_),
    .Y(_2907_),
    .A1(net1944),
    .A2(_2906_));
 sg13g2_nor3_2 _7352_ (.A(net2183),
    .B(_2904_),
    .C(_2907_),
    .Y(_2908_));
 sg13g2_nor2_1 _7353_ (.A(net2002),
    .B(_2385_),
    .Y(_2909_));
 sg13g2_a221oi_1 _7354_ (.B2(_1848_),
    .C1(_2909_),
    .B1(_2299_),
    .A1(net1814),
    .Y(_2910_),
    .A2(net1852));
 sg13g2_a21oi_1 _7355_ (.A1(_2640_),
    .A2(_2910_),
    .Y(_2911_),
    .B1(net2201));
 sg13g2_a21oi_1 _7356_ (.A1(_1546_),
    .A2(net1894),
    .Y(_2912_),
    .B1(_2644_));
 sg13g2_a21oi_1 _7357_ (.A1(net2011),
    .A2(net1903),
    .Y(_2913_),
    .B1(_1755_));
 sg13g2_a221oi_1 _7358_ (.B2(net1950),
    .C1(net2186),
    .B1(_2913_),
    .A1(net1888),
    .Y(_2914_),
    .A2(_2912_));
 sg13g2_nand2b_1 _7359_ (.Y(_2915_),
    .B(_2914_),
    .A_N(_2911_));
 sg13g2_a21oi_2 _7360_ (.B1(net2092),
    .Y(_2916_),
    .A2(_2649_),
    .A1(_1962_));
 sg13g2_o21ai_1 _7361_ (.B1(net1772),
    .Y(_2917_),
    .A1(net2181),
    .A2(_2908_));
 sg13g2_a21oi_2 _7362_ (.B1(_2917_),
    .Y(_2918_),
    .A2(_2916_),
    .A1(_2915_));
 sg13g2_o21ai_1 _7363_ (.B1(net2267),
    .Y(_2919_),
    .A1(net1918),
    .A2(_1740_));
 sg13g2_nand3_1 _7364_ (.B(_1764_),
    .C(_2919_),
    .A(net2088),
    .Y(_2920_));
 sg13g2_a21oi_1 _7365_ (.A1(net2244),
    .A2(_2920_),
    .Y(_2921_),
    .B1(_2737_));
 sg13g2_o21ai_1 _7366_ (.B1(net2075),
    .Y(_2922_),
    .A1(net1919),
    .A2(_1740_));
 sg13g2_nor3_1 _7367_ (.A(_1763_),
    .B(_1813_),
    .C(_2737_),
    .Y(_2923_));
 sg13g2_a21oi_1 _7368_ (.A1(_2386_),
    .A2(_2922_),
    .Y(_2924_),
    .B1(_2923_));
 sg13g2_o21ai_1 _7369_ (.B1(net2016),
    .Y(_2925_),
    .A1(_1587_),
    .A2(_2644_));
 sg13g2_o21ai_1 _7370_ (.B1(_2925_),
    .Y(_2926_),
    .A1(net2088),
    .A2(_2924_));
 sg13g2_o21ai_1 _7371_ (.B1(net1940),
    .Y(_2927_),
    .A1(_2921_),
    .A2(_2926_));
 sg13g2_a21oi_1 _7372_ (.A1(_2209_),
    .A2(_2705_),
    .Y(_2928_),
    .B1(_2729_));
 sg13g2_nor2_1 _7373_ (.A(_1623_),
    .B(net1871),
    .Y(_2929_));
 sg13g2_o21ai_1 _7374_ (.B1(net1889),
    .Y(_2930_),
    .A1(_2731_),
    .A2(_2929_));
 sg13g2_nor2_1 _7375_ (.A(_2928_),
    .B(_2930_),
    .Y(_2931_));
 sg13g2_a21oi_2 _7376_ (.B1(_2725_),
    .Y(_2932_),
    .A2(_1896_),
    .A1(net1855));
 sg13g2_nand2_1 _7377_ (.Y(_2933_),
    .A(_1863_),
    .B(_2932_));
 sg13g2_nand2_1 _7378_ (.Y(_2934_),
    .A(_1748_),
    .B(_1771_));
 sg13g2_nand2_1 _7379_ (.Y(_2935_),
    .A(net2261),
    .B(_1770_));
 sg13g2_o21ai_1 _7380_ (.B1(_2935_),
    .Y(_2936_),
    .A1(net2261),
    .A2(_1679_));
 sg13g2_a221oi_1 _7381_ (.B2(_1834_),
    .C1(net1981),
    .B1(_2934_),
    .A1(net2015),
    .Y(_2937_),
    .A2(_2933_));
 sg13g2_a221oi_1 _7382_ (.B2(_2936_),
    .C1(_2931_),
    .B1(_1890_),
    .A1(net1950),
    .Y(_2938_),
    .A2(_1839_));
 sg13g2_a22oi_1 _7383_ (.Y(_2939_),
    .B1(_2937_),
    .B2(_2938_),
    .A2(net1817),
    .A1(net1876));
 sg13g2_a21oi_2 _7384_ (.B1(_1936_),
    .Y(_2940_),
    .A2(_2939_),
    .A1(_2927_));
 sg13g2_a21oi_1 _7385_ (.A1(net2284),
    .A2(net2008),
    .Y(_2941_),
    .B1(_1728_));
 sg13g2_a21oi_1 _7386_ (.A1(_2779_),
    .A2(_2941_),
    .Y(_2942_),
    .B1(net1942));
 sg13g2_o21ai_1 _7387_ (.B1(net1848),
    .Y(_2943_),
    .A1(net2284),
    .A2(net1871));
 sg13g2_a221oi_1 _7388_ (.B2(net2221),
    .C1(net2209),
    .B1(_2047_),
    .A1(_1437_),
    .Y(_2944_),
    .A2(net2009));
 sg13g2_a221oi_1 _7389_ (.B2(_2944_),
    .C1(net2192),
    .B1(_2943_),
    .A1(net2206),
    .Y(_2945_),
    .A2(_1584_));
 sg13g2_a21oi_2 _7390_ (.B1(net1987),
    .Y(_2946_),
    .A2(_1712_),
    .A1(_1578_));
 sg13g2_nor4_1 _7391_ (.A(net1934),
    .B(_2942_),
    .C(_2945_),
    .D(_2946_),
    .Y(_2947_));
 sg13g2_nand2_1 _7392_ (.Y(_2948_),
    .A(net2104),
    .B(net1850));
 sg13g2_o21ai_1 _7393_ (.B1(_2948_),
    .Y(_2949_),
    .A1(net2008),
    .A2(_2104_));
 sg13g2_o21ai_1 _7394_ (.B1(_2949_),
    .Y(_2950_),
    .A1(_1899_),
    .A2(_2712_));
 sg13g2_and2_1 _7395_ (.A(net1884),
    .B(_2950_),
    .X(_2951_));
 sg13g2_a22oi_1 _7396_ (.Y(_2952_),
    .B1(_2136_),
    .B2(net1924),
    .A2(_2017_),
    .A1(net2104));
 sg13g2_nor3_1 _7397_ (.A(net2087),
    .B(_1710_),
    .C(_2952_),
    .Y(_2953_));
 sg13g2_nor2_1 _7398_ (.A(net2225),
    .B(_2692_),
    .Y(_2954_));
 sg13g2_nor3_1 _7399_ (.A(net2006),
    .B(net1985),
    .C(net1854),
    .Y(_2955_));
 sg13g2_a221oi_1 _7400_ (.B2(_2954_),
    .C1(_2955_),
    .B1(_2677_),
    .A1(net1890),
    .Y(_2956_),
    .A2(_2017_));
 sg13g2_o21ai_1 _7401_ (.B1(net1983),
    .Y(_2957_),
    .A1(_2951_),
    .A2(_2953_));
 sg13g2_o21ai_1 _7402_ (.B1(_2957_),
    .Y(_2958_),
    .A1(_1992_),
    .A2(_2956_));
 sg13g2_o21ai_1 _7403_ (.B1(net1770),
    .Y(_2959_),
    .A1(_2947_),
    .A2(_2958_));
 sg13g2_nand3_1 _7404_ (.B(net1813),
    .C(_2321_),
    .A(net1861),
    .Y(_2960_));
 sg13g2_a21o_1 _7405_ (.A2(_2960_),
    .A1(_1937_),
    .B1(_2763_),
    .X(_2961_));
 sg13g2_nor3_1 _7406_ (.A(_0091_),
    .B(net1933),
    .C(_1572_),
    .Y(_2962_));
 sg13g2_o21ai_1 _7407_ (.B1(net1813),
    .Y(_2963_),
    .A1(net1817),
    .A2(_2962_));
 sg13g2_a21oi_1 _7408_ (.A1(_2961_),
    .A2(_2963_),
    .Y(_2964_),
    .B1(_1861_));
 sg13g2_nand2_1 _7409_ (.Y(_2965_),
    .A(net1938),
    .B(_2665_));
 sg13g2_nor2_1 _7410_ (.A(net2250),
    .B(_1982_),
    .Y(_2966_));
 sg13g2_o21ai_1 _7411_ (.B1(net2086),
    .Y(_2967_),
    .A1(net1909),
    .A2(net1897));
 sg13g2_a21oi_1 _7412_ (.A1(net1909),
    .A2(_2966_),
    .Y(_2968_),
    .B1(_2967_));
 sg13g2_a22oi_1 _7413_ (.Y(_2969_),
    .B1(_2081_),
    .B2(_1761_),
    .A2(_1993_),
    .A1(_1921_));
 sg13g2_o21ai_1 _7414_ (.B1(_2969_),
    .Y(_2970_),
    .A1(_2965_),
    .A2(_2968_));
 sg13g2_nand2_1 _7415_ (.Y(_2971_),
    .A(_1829_),
    .B(_2970_));
 sg13g2_a21oi_1 _7416_ (.A1(_2623_),
    .A2(_2870_),
    .Y(_2972_),
    .B1(_2940_));
 sg13g2_o21ai_1 _7417_ (.B1(_2972_),
    .Y(_2973_),
    .A1(net1933),
    .A2(_2836_));
 sg13g2_nor4_2 _7418_ (.A(_1538_),
    .B(_2901_),
    .C(_2918_),
    .Y(_2974_),
    .D(_2964_));
 sg13g2_nand3_1 _7419_ (.B(_2971_),
    .C(_2974_),
    .A(_2959_),
    .Y(_2975_));
 sg13g2_nor4_2 _7420_ (.A(_2854_),
    .B(_2896_),
    .C(_2973_),
    .Y(_2976_),
    .D(_2975_));
 sg13g2_o21ai_1 _7421_ (.B1(_1565_),
    .Y(_2977_),
    .A1(net1929),
    .A2(_1594_));
 sg13g2_a221oi_1 _7422_ (.B2(net2187),
    .C1(_2977_),
    .B1(_2810_),
    .A1(net1949),
    .Y(_2978_),
    .A2(_1589_));
 sg13g2_nor2_1 _7423_ (.A(net2184),
    .B(_2978_),
    .Y(_2979_));
 sg13g2_nor3_1 _7424_ (.A(net1929),
    .B(_1588_),
    .C(_1921_),
    .Y(_2980_));
 sg13g2_nand2b_1 _7425_ (.Y(_2981_),
    .B(_2818_),
    .A_N(_2980_));
 sg13g2_o21ai_1 _7426_ (.B1(_2981_),
    .Y(_2982_),
    .A1(_2808_),
    .A2(_2979_));
 sg13g2_o21ai_1 _7427_ (.B1(\draw_game_inst.board_x[0] ),
    .Y(_2983_),
    .A1(net1756),
    .A2(_2982_));
 sg13g2_nor2_1 _7428_ (.A(\draw_game_inst.board_x[1] ),
    .B(_2822_),
    .Y(_2984_));
 sg13g2_o21ai_1 _7429_ (.B1(_2984_),
    .Y(_2985_),
    .A1(_2976_),
    .A2(_2983_));
 sg13g2_a21oi_1 _7430_ (.A1(_1654_),
    .A2(_1915_),
    .Y(_2986_),
    .B1(net1935));
 sg13g2_o21ai_1 _7431_ (.B1(_2986_),
    .Y(_2987_),
    .A1(_1685_),
    .A2(_2168_));
 sg13g2_nand2_1 _7432_ (.Y(_2988_),
    .A(_1918_),
    .B(_2987_));
 sg13g2_o21ai_1 _7433_ (.B1(net2189),
    .Y(_2989_),
    .A1(net2204),
    .A2(_2274_));
 sg13g2_o21ai_1 _7434_ (.B1(_2989_),
    .Y(_2990_),
    .A1(net2189),
    .A2(_2073_));
 sg13g2_nor3_1 _7435_ (.A(_1568_),
    .B(_2988_),
    .C(_2990_),
    .Y(_2991_));
 sg13g2_nor2_1 _7436_ (.A(net1893),
    .B(_1769_),
    .Y(_2992_));
 sg13g2_o21ai_1 _7437_ (.B1(_2154_),
    .Y(_2993_),
    .A1(net1892),
    .A2(_1769_));
 sg13g2_a221oi_1 _7438_ (.B2(net2083),
    .C1(_2133_),
    .B1(_2993_),
    .A1(net1814),
    .Y(_2994_),
    .A2(net1852));
 sg13g2_a21oi_1 _7439_ (.A1(net1886),
    .A2(_2406_),
    .Y(_2995_),
    .B1(_2142_));
 sg13g2_o21ai_1 _7440_ (.B1(_2995_),
    .Y(_2996_),
    .A1(net2197),
    .A2(_2994_));
 sg13g2_nand2b_1 _7441_ (.Y(_2997_),
    .B(_2935_),
    .A_N(_2131_));
 sg13g2_nand2_1 _7442_ (.Y(_2998_),
    .A(net2072),
    .B(_2997_));
 sg13g2_nand2_1 _7443_ (.Y(_2999_),
    .A(net2243),
    .B(_1770_));
 sg13g2_a21oi_1 _7444_ (.A1(net2238),
    .A2(_1770_),
    .Y(_3000_),
    .B1(net2082));
 sg13g2_a221oi_1 _7445_ (.B2(_3000_),
    .C1(net2197),
    .B1(_2998_),
    .A1(_1949_),
    .Y(_3001_),
    .A2(_2311_));
 sg13g2_a221oi_1 _7446_ (.B2(_1771_),
    .C1(net1946),
    .B1(_2356_),
    .A1(net2238),
    .Y(_3002_),
    .A2(net1813));
 sg13g2_nand4_1 _7447_ (.B(net1888),
    .C(net1870),
    .A(net1893),
    .Y(_3003_),
    .D(net1821));
 sg13g2_o21ai_1 _7448_ (.B1(_3003_),
    .Y(_3004_),
    .A1(_2109_),
    .A2(_2862_));
 sg13g2_nor4_1 _7449_ (.A(net2183),
    .B(_3001_),
    .C(_3002_),
    .D(_3004_),
    .Y(_3005_));
 sg13g2_a221oi_1 _7450_ (.B2(net1940),
    .C1(_1936_),
    .B1(_2996_),
    .A1(_1575_),
    .Y(_3006_),
    .A2(_2159_));
 sg13g2_o21ai_1 _7451_ (.B1(_3006_),
    .Y(_3007_),
    .A1(net2181),
    .A2(_3005_));
 sg13g2_nand2_1 _7452_ (.Y(_3008_),
    .A(_1765_),
    .B(_1999_));
 sg13g2_inv_1 _7453_ (.Y(_3009_),
    .A(_3008_));
 sg13g2_nand2b_1 _7454_ (.Y(_3010_),
    .B(_2919_),
    .A_N(_1750_));
 sg13g2_a221oi_1 _7455_ (.B2(net2231),
    .C1(net2080),
    .B1(_2649_),
    .A1(net1914),
    .Y(_3011_),
    .A2(_1705_));
 sg13g2_a221oi_1 _7456_ (.B2(net1996),
    .C1(_3011_),
    .B1(_3010_),
    .A1(net1867),
    .Y(_3012_),
    .A2(_3009_));
 sg13g2_nand3_1 _7457_ (.B(_1856_),
    .C(_3012_),
    .A(_1702_),
    .Y(_3013_));
 sg13g2_nand3_1 _7458_ (.B(_1722_),
    .C(net1861),
    .A(_1706_),
    .Y(_3014_));
 sg13g2_nor3_1 _7459_ (.A(net1825),
    .B(_1810_),
    .C(_2353_),
    .Y(_3015_));
 sg13g2_nor3_1 _7460_ (.A(net2008),
    .B(net1891),
    .C(net1850),
    .Y(_3016_));
 sg13g2_or3_1 _7461_ (.A(_1794_),
    .B(_3015_),
    .C(_3016_),
    .X(_3017_));
 sg13g2_nand2_2 _7462_ (.Y(_3018_),
    .A(net1914),
    .B(_2191_));
 sg13g2_nand3_1 _7463_ (.B(_1983_),
    .C(_3018_),
    .A(net2229),
    .Y(_3019_));
 sg13g2_a221oi_1 _7464_ (.B2(net1922),
    .C1(net1987),
    .B1(net1848),
    .A1(net2012),
    .Y(_3020_),
    .A2(net1836));
 sg13g2_a22oi_1 _7465_ (.Y(_3021_),
    .B1(_3019_),
    .B2(_3020_),
    .A2(_3014_),
    .A1(net1863));
 sg13g2_nand2_1 _7466_ (.Y(_3022_),
    .A(net1868),
    .B(_2049_));
 sg13g2_nand3_1 _7467_ (.B(_2948_),
    .C(_3018_),
    .A(net1997),
    .Y(_3023_));
 sg13g2_o21ai_1 _7468_ (.B1(_2165_),
    .Y(_3024_),
    .A1(_1545_),
    .A2(_1640_));
 sg13g2_nand4_1 _7469_ (.B(_3022_),
    .C(_3023_),
    .A(net2191),
    .Y(_3025_),
    .D(_3024_));
 sg13g2_a22oi_1 _7470_ (.Y(_3026_),
    .B1(net1848),
    .B2(net2284),
    .A2(_1790_),
    .A1(net2229));
 sg13g2_a21oi_1 _7471_ (.A1(_1729_),
    .A2(_3026_),
    .Y(_3027_),
    .B1(net1930));
 sg13g2_o21ai_1 _7472_ (.B1(net1906),
    .Y(_3028_),
    .A1(net2229),
    .A2(_1790_));
 sg13g2_a21oi_1 _7473_ (.A1(net2229),
    .A2(_2032_),
    .Y(_3029_),
    .B1(_3028_));
 sg13g2_nor3_1 _7474_ (.A(net1934),
    .B(_3027_),
    .C(_3029_),
    .Y(_3030_));
 sg13g2_a22oi_1 _7475_ (.Y(_3031_),
    .B1(_3025_),
    .B2(_3030_),
    .A2(_3021_),
    .A1(_3017_));
 sg13g2_nand2b_1 _7476_ (.Y(_3032_),
    .B(_1981_),
    .A_N(_3031_));
 sg13g2_o21ai_1 _7477_ (.B1(net1856),
    .Y(_3033_),
    .A1(_1683_),
    .A2(_1740_));
 sg13g2_a21oi_1 _7478_ (.A1(net1895),
    .A2(_2018_),
    .Y(_3034_),
    .B1(net2203));
 sg13g2_a21oi_2 _7479_ (.B1(net2199),
    .Y(_3035_),
    .A2(_3034_),
    .A1(_3033_));
 sg13g2_o21ai_1 _7480_ (.B1(net1883),
    .Y(_3036_),
    .A1(net2227),
    .A2(net1850));
 sg13g2_a21oi_1 _7481_ (.A1(net2227),
    .A2(net1922),
    .Y(_3037_),
    .B1(_3036_));
 sg13g2_a21oi_1 _7482_ (.A1(_1749_),
    .A2(_2238_),
    .Y(_3038_),
    .B1(_1556_));
 sg13g2_a21oi_1 _7483_ (.A1(net2017),
    .A2(net2008),
    .Y(_3039_),
    .B1(_2224_));
 sg13g2_nor4_1 _7484_ (.A(_3035_),
    .B(_3037_),
    .C(_3038_),
    .D(_3039_),
    .Y(_3040_));
 sg13g2_nand3_1 _7485_ (.B(net1983),
    .C(_3040_),
    .A(net1770),
    .Y(_3041_));
 sg13g2_nand4_1 _7486_ (.B(_3013_),
    .C(_3032_),
    .A(_3007_),
    .Y(_3042_),
    .D(_3041_));
 sg13g2_nor2_1 _7487_ (.A(_2991_),
    .B(_3042_),
    .Y(_3043_));
 sg13g2_a21o_1 _7488_ (.A2(_1882_),
    .A1(net2075),
    .B1(net2084),
    .X(_3044_));
 sg13g2_o21ai_1 _7489_ (.B1(net1894),
    .Y(_3045_),
    .A1(net1919),
    .A2(_2178_));
 sg13g2_o21ai_1 _7490_ (.B1(_3045_),
    .Y(_3046_),
    .A1(_1801_),
    .A2(_2109_));
 sg13g2_nor3_1 _7491_ (.A(net2199),
    .B(_3044_),
    .C(_3046_),
    .Y(_3047_));
 sg13g2_a221oi_1 _7492_ (.B2(_1788_),
    .C1(_2195_),
    .B1(net1879),
    .A1(net2265),
    .Y(_3048_),
    .A2(net2030));
 sg13g2_nand3_1 _7493_ (.B(net1875),
    .C(_2037_),
    .A(net2108),
    .Y(_3049_));
 sg13g2_o21ai_1 _7494_ (.B1(net1840),
    .Y(_3050_),
    .A1(_1715_),
    .A2(_1787_));
 sg13g2_nor2b_1 _7495_ (.A(_3050_),
    .B_N(_3049_),
    .Y(_3051_));
 sg13g2_nor3_1 _7496_ (.A(_3047_),
    .B(_3048_),
    .C(_3051_),
    .Y(_3052_));
 sg13g2_o21ai_1 _7497_ (.B1(_3052_),
    .Y(_3053_),
    .A1(_2120_),
    .A2(_2253_));
 sg13g2_o21ai_1 _7498_ (.B1(net2240),
    .Y(_3054_),
    .A1(net1882),
    .A2(_1788_));
 sg13g2_nand3_1 _7499_ (.B(_1742_),
    .C(net1849),
    .A(net2005),
    .Y(_3055_));
 sg13g2_nand3_1 _7500_ (.B(_3054_),
    .C(_3055_),
    .A(_1657_),
    .Y(_3056_));
 sg13g2_a21oi_1 _7501_ (.A1(net2010),
    .A2(_2495_),
    .Y(_3057_),
    .B1(_3056_));
 sg13g2_o21ai_1 _7502_ (.B1(_3049_),
    .Y(_3058_),
    .A1(_1457_),
    .A2(_1965_));
 sg13g2_a21oi_1 _7503_ (.A1(_1862_),
    .A2(_2681_),
    .Y(_3059_),
    .B1(net2084));
 sg13g2_nand3_1 _7504_ (.B(_1790_),
    .C(_2283_),
    .A(net2241),
    .Y(_3060_));
 sg13g2_a22oi_1 _7505_ (.Y(_3061_),
    .B1(_3059_),
    .B2(_3060_),
    .A2(_2831_),
    .A1(net1867));
 sg13g2_o21ai_1 _7506_ (.B1(_3061_),
    .Y(_3062_),
    .A1(_1582_),
    .A2(_3058_));
 sg13g2_a21o_1 _7507_ (.A2(_3062_),
    .A1(net2088),
    .B1(_3057_),
    .X(_3063_));
 sg13g2_a22oi_1 _7508_ (.Y(_3064_),
    .B1(_3063_),
    .B2(net1771),
    .A2(_3053_),
    .A1(_1702_));
 sg13g2_nor2_1 _7509_ (.A(net1935),
    .B(_3064_),
    .Y(_3065_));
 sg13g2_nand3_1 _7510_ (.B(_2154_),
    .C(_2310_),
    .A(_1627_),
    .Y(_3066_));
 sg13g2_a21oi_2 _7511_ (.B1(_2290_),
    .Y(_3067_),
    .A2(_1786_),
    .A1(net1869));
 sg13g2_nor2_1 _7512_ (.A(_1562_),
    .B(net1988),
    .Y(_3068_));
 sg13g2_o21ai_1 _7513_ (.B1(_2866_),
    .Y(_3069_),
    .A1(net2235),
    .A2(_2385_));
 sg13g2_a221oi_1 _7514_ (.B2(_3068_),
    .C1(net2185),
    .B1(_2254_),
    .A1(net1950),
    .Y(_3070_),
    .A2(net1819));
 sg13g2_o21ai_1 _7515_ (.B1(_3070_),
    .Y(_3071_),
    .A1(_1884_),
    .A2(_3067_));
 sg13g2_a221oi_1 _7516_ (.B2(net1907),
    .C1(_3071_),
    .B1(_3069_),
    .A1(net2015),
    .Y(_3072_),
    .A2(_3066_));
 sg13g2_and2_1 _7517_ (.A(_1962_),
    .B(_2826_),
    .X(_3073_));
 sg13g2_o21ai_1 _7518_ (.B1(_1615_),
    .Y(_3074_),
    .A1(_3072_),
    .A2(_3073_));
 sg13g2_nor2_1 _7519_ (.A(net2188),
    .B(_2631_),
    .Y(_3075_));
 sg13g2_nand2b_1 _7520_ (.Y(_3076_),
    .B(_3075_),
    .A_N(_1588_));
 sg13g2_nor3_1 _7521_ (.A(_1430_),
    .B(net1839),
    .C(_1649_),
    .Y(_3077_));
 sg13g2_nor2_2 _7522_ (.A(net2017),
    .B(net1824),
    .Y(_3078_));
 sg13g2_nor4_1 _7523_ (.A(net2184),
    .B(_2946_),
    .C(_3077_),
    .D(_3078_),
    .Y(_3079_));
 sg13g2_o21ai_1 _7524_ (.B1(_2034_),
    .Y(_3080_),
    .A1(net2253),
    .A2(_2046_));
 sg13g2_a21oi_1 _7525_ (.A1(_1810_),
    .A2(_2871_),
    .Y(_3081_),
    .B1(_1558_));
 sg13g2_a21oi_1 _7526_ (.A1(_2194_),
    .A2(_3080_),
    .Y(_3082_),
    .B1(_3081_));
 sg13g2_nand4_1 _7527_ (.B(_3076_),
    .C(_3079_),
    .A(net1770),
    .Y(_3083_),
    .D(_3082_));
 sg13g2_nand3_1 _7528_ (.B(_3074_),
    .C(_3083_),
    .A(_2988_),
    .Y(_3084_));
 sg13g2_and2_1 _7529_ (.A(net2180),
    .B(_3084_),
    .X(_3085_));
 sg13g2_o21ai_1 _7530_ (.B1(_3018_),
    .Y(_3086_),
    .A1(net2256),
    .A2(_2046_));
 sg13g2_a22oi_1 _7531_ (.Y(_3087_),
    .B1(_3086_),
    .B2(net2228),
    .A2(_1735_),
    .A1(net1920));
 sg13g2_nand2_1 _7532_ (.Y(_3088_),
    .A(net1861),
    .B(_3087_));
 sg13g2_o21ai_1 _7533_ (.B1(net1883),
    .Y(_3089_),
    .A1(net2223),
    .A2(_1790_));
 sg13g2_a221oi_1 _7534_ (.B2(_3089_),
    .C1(_1545_),
    .B1(_2523_),
    .A1(_1436_),
    .Y(_3090_),
    .A2(_1665_));
 sg13g2_a221oi_1 _7535_ (.B2(net1863),
    .C1(_3090_),
    .B1(_3088_),
    .A1(net1914),
    .Y(_3091_),
    .A2(_3078_));
 sg13g2_nor2_1 _7536_ (.A(_1547_),
    .B(_2883_),
    .Y(_3092_));
 sg13g2_nor2_1 _7537_ (.A(_1695_),
    .B(_2544_),
    .Y(_3093_));
 sg13g2_nor2_1 _7538_ (.A(net1930),
    .B(_3093_),
    .Y(_3094_));
 sg13g2_a221oi_1 _7539_ (.B2(net2223),
    .C1(net1904),
    .B1(net1820),
    .A1(net2066),
    .Y(_3095_),
    .A2(net2286));
 sg13g2_nor4_1 _7540_ (.A(_2881_),
    .B(_3092_),
    .C(_3094_),
    .D(_3095_),
    .Y(_3096_));
 sg13g2_nor2_1 _7541_ (.A(_3091_),
    .B(_3096_),
    .Y(_3097_));
 sg13g2_o21ai_1 _7542_ (.B1(net1756),
    .Y(_3098_),
    .A1(_1782_),
    .A2(_3097_));
 sg13g2_nand3_1 _7543_ (.B(net1839),
    .C(net1861),
    .A(net1924),
    .Y(_3099_));
 sg13g2_nand2_1 _7544_ (.Y(_3100_),
    .A(_2965_),
    .B(_3099_));
 sg13g2_nor3_1 _7545_ (.A(net2251),
    .B(_1982_),
    .C(_2172_),
    .Y(_3101_));
 sg13g2_a21oi_1 _7546_ (.A1(net1839),
    .A2(_1654_),
    .Y(_3102_),
    .B1(_3101_));
 sg13g2_o21ai_1 _7547_ (.B1(net2086),
    .Y(_3103_),
    .A1(net1932),
    .A2(_3102_));
 sg13g2_nand2_1 _7548_ (.Y(_3104_),
    .A(_3100_),
    .B(_3103_));
 sg13g2_a21oi_1 _7549_ (.A1(net2079),
    .A2(_0093_),
    .Y(_3105_),
    .B1(net1913));
 sg13g2_o21ai_1 _7550_ (.B1(_3105_),
    .Y(_3106_),
    .A1(net2250),
    .A2(net2003));
 sg13g2_o21ai_1 _7551_ (.B1(_3104_),
    .Y(_3107_),
    .A1(_1937_),
    .A2(_3106_));
 sg13g2_o21ai_1 _7552_ (.B1(net2071),
    .Y(_3108_),
    .A1(net1827),
    .A2(_1748_));
 sg13g2_a221oi_1 _7553_ (.B2(_1908_),
    .C1(net2196),
    .B1(_3108_),
    .A1(_2719_),
    .Y(_3109_),
    .A2(_2998_));
 sg13g2_a21oi_1 _7554_ (.A1(net2237),
    .A2(_1946_),
    .Y(_3110_),
    .B1(_2074_));
 sg13g2_o21ai_1 _7555_ (.B1(net2195),
    .Y(_3111_),
    .A1(net1926),
    .A2(net1902));
 sg13g2_nor3_1 _7556_ (.A(_1675_),
    .B(_2070_),
    .C(_3111_),
    .Y(_3112_));
 sg13g2_nor4_2 _7557_ (.A(net1981),
    .B(_3109_),
    .C(_3110_),
    .Y(_3113_),
    .D(_3112_));
 sg13g2_a221oi_1 _7558_ (.B2(net1772),
    .C1(_3098_),
    .B1(_3113_),
    .A1(_1829_),
    .Y(_3114_),
    .A2(_3107_));
 sg13g2_a21oi_1 _7559_ (.A1(_2038_),
    .A2(_2847_),
    .Y(_3115_),
    .B1(net2229));
 sg13g2_a21oi_1 _7560_ (.A1(_1684_),
    .A2(_1721_),
    .Y(_3116_),
    .B1(net1991));
 sg13g2_a21oi_1 _7561_ (.A1(_1721_),
    .A2(_2036_),
    .Y(_3117_),
    .B1(net1854));
 sg13g2_nor4_1 _7562_ (.A(net2209),
    .B(_3115_),
    .C(_3116_),
    .D(_3117_),
    .Y(_3118_));
 sg13g2_a221oi_1 _7563_ (.B2(net1853),
    .C1(_3118_),
    .B1(_3009_),
    .A1(net2215),
    .Y(_3119_),
    .A2(_2687_));
 sg13g2_or2_1 _7564_ (.X(_3120_),
    .B(_3119_),
    .A(_1858_));
 sg13g2_a21oi_1 _7565_ (.A1(_1627_),
    .A2(_2102_),
    .Y(_3121_),
    .B1(net1988));
 sg13g2_a22oi_1 _7566_ (.Y(_3122_),
    .B1(_2343_),
    .B2(net2015),
    .A2(net1822),
    .A1(net1907));
 sg13g2_nand2_1 _7567_ (.Y(_3123_),
    .A(_2118_),
    .B(_3122_));
 sg13g2_o21ai_1 _7568_ (.B1(net1939),
    .Y(_3124_),
    .A1(_3121_),
    .A2(_3123_));
 sg13g2_o21ai_1 _7569_ (.B1(net1998),
    .Y(_3125_),
    .A1(net1827),
    .A2(_1748_));
 sg13g2_nand2_1 _7570_ (.Y(_3126_),
    .A(_2111_),
    .B(_3125_));
 sg13g2_a221oi_1 _7571_ (.B2(net1910),
    .C1(_3126_),
    .B1(_2114_),
    .A1(net1852),
    .Y(_3127_),
    .A2(_2112_));
 sg13g2_nor2_1 _7572_ (.A(net2236),
    .B(_2113_),
    .Y(_3128_));
 sg13g2_a22oi_1 _7573_ (.Y(_3129_),
    .B1(_1850_),
    .B2(_3128_),
    .A2(net1822),
    .A1(net2236));
 sg13g2_nor2_1 _7574_ (.A(net1946),
    .B(_3129_),
    .Y(_3130_));
 sg13g2_o21ai_1 _7575_ (.B1(_2124_),
    .Y(_3131_),
    .A1(net2195),
    .A2(_3127_));
 sg13g2_o21ai_1 _7576_ (.B1(net2092),
    .Y(_3132_),
    .A1(_3130_),
    .A2(_3131_));
 sg13g2_nand3_1 _7577_ (.B(_3124_),
    .C(_3132_),
    .A(_2100_),
    .Y(_3133_));
 sg13g2_nand3_1 _7578_ (.B(_3120_),
    .C(_3133_),
    .A(_3114_),
    .Y(_3134_));
 sg13g2_nor3_2 _7579_ (.A(_3065_),
    .B(_3085_),
    .C(_3134_),
    .Y(_3135_));
 sg13g2_o21ai_1 _7580_ (.B1(net2079),
    .Y(_3136_),
    .A1(net1913),
    .A2(net2000));
 sg13g2_a221oi_1 _7581_ (.B2(_2278_),
    .C1(net2184),
    .B1(_3136_),
    .A1(_2441_),
    .Y(_3137_),
    .A2(_2811_));
 sg13g2_nor2_1 _7582_ (.A(_2808_),
    .B(_3137_),
    .Y(_3138_));
 sg13g2_a21oi_1 _7583_ (.A1(net2205),
    .A2(_1930_),
    .Y(_3139_),
    .B1(_1937_));
 sg13g2_o21ai_1 _7584_ (.B1(_3139_),
    .Y(_3140_),
    .A1(_1675_),
    .A2(_1921_));
 sg13g2_nor2_1 _7585_ (.A(net1757),
    .B(_3138_),
    .Y(_3141_));
 sg13g2_a22oi_1 _7586_ (.Y(_3142_),
    .B1(_3140_),
    .B2(_3141_),
    .A2(_3135_),
    .A1(_3043_));
 sg13g2_nand2b_1 _7587_ (.Y(_3143_),
    .B(_1440_),
    .A_N(_3142_));
 sg13g2_a22oi_1 _7588_ (.Y(_3144_),
    .B1(_1949_),
    .B2(_2932_),
    .A2(_1769_),
    .A1(net2212));
 sg13g2_nand2_1 _7589_ (.Y(_3145_),
    .A(net1994),
    .B(net1825));
 sg13g2_a21oi_1 _7590_ (.A1(net1893),
    .A2(_2422_),
    .Y(_3146_),
    .B1(net1989));
 sg13g2_a21oi_1 _7591_ (.A1(net2243),
    .A2(_1938_),
    .Y(_3147_),
    .B1(_2406_));
 sg13g2_o21ai_1 _7592_ (.B1(net1984),
    .Y(_3148_),
    .A1(net1945),
    .A2(_3147_));
 sg13g2_a221oi_1 _7593_ (.B2(_3146_),
    .C1(_3148_),
    .B1(_3145_),
    .A1(net2090),
    .Y(_3149_),
    .A2(_3144_));
 sg13g2_o21ai_1 _7594_ (.B1(net1817),
    .Y(_3150_),
    .A1(net1837),
    .A2(net1877));
 sg13g2_o21ai_1 _7595_ (.B1(net1889),
    .Y(_3151_),
    .A1(_2140_),
    .A2(_2992_));
 sg13g2_a21oi_1 _7596_ (.A1(_2422_),
    .A2(_2999_),
    .Y(_3152_),
    .B1(net1931));
 sg13g2_a21oi_1 _7597_ (.A1(net1893),
    .A2(net1985),
    .Y(_3153_),
    .B1(_2992_));
 sg13g2_a21oi_1 _7598_ (.A1(_2550_),
    .A2(_2999_),
    .Y(_3154_),
    .B1(net1944));
 sg13g2_o21ai_1 _7599_ (.B1(_3151_),
    .Y(_3155_),
    .A1(net1904),
    .A2(_3153_));
 sg13g2_nor4_1 _7600_ (.A(net1936),
    .B(_3152_),
    .C(_3154_),
    .D(_3155_),
    .Y(_3156_));
 sg13g2_nor2_1 _7601_ (.A(_3149_),
    .B(_3156_),
    .Y(_3157_));
 sg13g2_a21oi_2 _7602_ (.B1(_1936_),
    .Y(_3158_),
    .A2(_3157_),
    .A1(_3150_));
 sg13g2_o21ai_1 _7603_ (.B1(net2217),
    .Y(_3159_),
    .A1(net1814),
    .A2(_1944_));
 sg13g2_nor2b_1 _7604_ (.A(_1628_),
    .B_N(_3159_),
    .Y(_3160_));
 sg13g2_a21oi_1 _7605_ (.A1(_2640_),
    .A2(_3160_),
    .Y(_3161_),
    .B1(net2201));
 sg13g2_nand3_1 _7606_ (.B(_1745_),
    .C(_1748_),
    .A(net2075),
    .Y(_3162_));
 sg13g2_and3_1 _7607_ (.X(_3163_),
    .A(net1888),
    .B(_2458_),
    .C(_3162_));
 sg13g2_a21oi_1 _7608_ (.A1(net1893),
    .A2(_1743_),
    .Y(_3164_),
    .B1(_2072_));
 sg13g2_nor4_2 _7609_ (.A(net1936),
    .B(_3161_),
    .C(_3163_),
    .Y(_3165_),
    .D(_3164_));
 sg13g2_nand3_1 _7610_ (.B(_1704_),
    .C(net1817),
    .A(net1825),
    .Y(_3166_));
 sg13g2_nand3_1 _7611_ (.B(_2809_),
    .C(_2906_),
    .A(_1761_),
    .Y(_3167_));
 sg13g2_nand2_1 _7612_ (.Y(_3168_),
    .A(net1852),
    .B(_2423_));
 sg13g2_nand2b_1 _7613_ (.Y(_3169_),
    .B(_3126_),
    .A_N(_1587_));
 sg13g2_a21oi_1 _7614_ (.A1(net1902),
    .A2(_2899_),
    .Y(_3170_),
    .B1(_1937_));
 sg13g2_nand3_1 _7615_ (.B(_3169_),
    .C(_3170_),
    .A(_3168_),
    .Y(_3171_));
 sg13g2_nand3_1 _7616_ (.B(_3167_),
    .C(_3171_),
    .A(_3166_),
    .Y(_3172_));
 sg13g2_o21ai_1 _7617_ (.B1(net1772),
    .Y(_3173_),
    .A1(_3165_),
    .A2(_3172_));
 sg13g2_a22oi_1 _7618_ (.Y(_3174_),
    .B1(net1857),
    .B2(_2033_),
    .A2(_1790_),
    .A1(net1891));
 sg13g2_a21oi_1 _7619_ (.A1(_1729_),
    .A2(_3174_),
    .Y(_3175_),
    .B1(net1930));
 sg13g2_a21oi_1 _7620_ (.A1(_2031_),
    .A2(_2135_),
    .Y(_3176_),
    .B1(net1990));
 sg13g2_a221oi_1 _7621_ (.B2(_1750_),
    .C1(net2070),
    .B1(_1713_),
    .A1(net2257),
    .Y(_3177_),
    .A2(_1458_));
 sg13g2_o21ai_1 _7622_ (.B1(net1948),
    .Y(_3178_),
    .A1(_1728_),
    .A2(_3177_));
 sg13g2_nor2_1 _7623_ (.A(net2070),
    .B(_2191_),
    .Y(_3179_));
 sg13g2_o21ai_1 _7624_ (.B1(_3179_),
    .Y(_3180_),
    .A1(net2258),
    .A2(_1789_));
 sg13g2_nor2b_1 _7625_ (.A(_3028_),
    .B_N(_3180_),
    .Y(_3181_));
 sg13g2_nand3_1 _7626_ (.B(_1655_),
    .C(_2114_),
    .A(_1461_),
    .Y(_3182_));
 sg13g2_nor2b_1 _7627_ (.A(net2240),
    .B_N(net2295),
    .Y(_3183_));
 sg13g2_a21oi_1 _7628_ (.A1(net1856),
    .A2(_2018_),
    .Y(_3184_),
    .B1(_3183_));
 sg13g2_o21ai_1 _7629_ (.B1(_3182_),
    .Y(_3185_),
    .A1(net2215),
    .A2(_3184_));
 sg13g2_nor2_1 _7630_ (.A(net1851),
    .B(_2530_),
    .Y(_3186_));
 sg13g2_or4_1 _7631_ (.A(net2086),
    .B(_1968_),
    .C(_2856_),
    .D(_3186_),
    .X(_3187_));
 sg13g2_o21ai_1 _7632_ (.B1(_1567_),
    .Y(_3188_),
    .A1(net1913),
    .A2(net1891));
 sg13g2_a21oi_1 _7633_ (.A1(_1635_),
    .A2(_3188_),
    .Y(_3189_),
    .B1(net1932));
 sg13g2_nand2b_1 _7634_ (.Y(_3190_),
    .B(_2560_),
    .A_N(_1427_));
 sg13g2_o21ai_1 _7635_ (.B1(_3190_),
    .Y(_3191_),
    .A1(net2189),
    .A2(_2815_));
 sg13g2_nor2_1 _7636_ (.A(_2809_),
    .B(_3191_),
    .Y(_3192_));
 sg13g2_nor3_1 _7637_ (.A(net2182),
    .B(_2855_),
    .C(_3192_),
    .Y(_3193_));
 sg13g2_a21oi_1 _7638_ (.A1(_2861_),
    .A2(_3193_),
    .Y(_3194_),
    .B1(net2179));
 sg13g2_a21oi_1 _7639_ (.A1(_3187_),
    .A2(_3189_),
    .Y(_3195_),
    .B1(_3194_));
 sg13g2_nand2_1 _7640_ (.Y(_3196_),
    .A(net2066),
    .B(_2091_));
 sg13g2_a21oi_1 _7641_ (.A1(net1853),
    .A2(_2345_),
    .Y(_3197_),
    .B1(_3196_));
 sg13g2_or2_1 _7642_ (.X(_3198_),
    .B(_3197_),
    .A(net2188));
 sg13g2_nor3_1 _7643_ (.A(net2223),
    .B(_1977_),
    .C(_2119_),
    .Y(_3199_));
 sg13g2_nor2_1 _7644_ (.A(_2883_),
    .B(_3199_),
    .Y(_3200_));
 sg13g2_nor2_1 _7645_ (.A(_2881_),
    .B(_3200_),
    .Y(_3201_));
 sg13g2_a21oi_1 _7646_ (.A1(_2238_),
    .A2(_2677_),
    .Y(_3202_),
    .B1(_1556_));
 sg13g2_a22oi_1 _7647_ (.Y(_3203_),
    .B1(_2047_),
    .B2(net2224),
    .A2(_1812_),
    .A1(_1735_));
 sg13g2_a221oi_1 _7648_ (.B2(net1914),
    .C1(net1980),
    .B1(_3078_),
    .A1(_2047_),
    .Y(_3204_),
    .A2(_2414_));
 sg13g2_o21ai_1 _7649_ (.B1(_3204_),
    .Y(_3205_),
    .A1(net1986),
    .A2(_3203_));
 sg13g2_nor2_1 _7650_ (.A(_3202_),
    .B(_3205_),
    .Y(_3206_));
 sg13g2_a22oi_1 _7651_ (.Y(_3207_),
    .B1(_3206_),
    .B2(_2874_),
    .A2(_3201_),
    .A1(_3198_));
 sg13g2_o21ai_1 _7652_ (.B1(net1756),
    .Y(_3208_),
    .A1(_1782_),
    .A2(_3207_));
 sg13g2_a21oi_1 _7653_ (.A1(net1813),
    .A2(_1961_),
    .Y(_3209_),
    .B1(net1939));
 sg13g2_a22oi_1 _7654_ (.Y(_3210_),
    .B1(net1996),
    .B2(_2781_),
    .A2(_1565_),
    .A1(_1558_));
 sg13g2_a21o_1 _7655_ (.A2(_1584_),
    .A1(net2079),
    .B1(net2085),
    .X(_3211_));
 sg13g2_nor2_1 _7656_ (.A(_1620_),
    .B(_2172_),
    .Y(_3212_));
 sg13g2_a21oi_1 _7657_ (.A1(net1813),
    .A2(_3212_),
    .Y(_3213_),
    .B1(_3211_));
 sg13g2_nor2_1 _7658_ (.A(_3210_),
    .B(_3213_),
    .Y(_3214_));
 sg13g2_nor2_1 _7659_ (.A(net2185),
    .B(_3214_),
    .Y(_3215_));
 sg13g2_nor2_1 _7660_ (.A(_3209_),
    .B(_3215_),
    .Y(_3216_));
 sg13g2_a22oi_1 _7661_ (.Y(_3217_),
    .B1(_1682_),
    .B2(_2899_),
    .A2(net1830),
    .A1(net1998));
 sg13g2_a21oi_1 _7662_ (.A1(_2300_),
    .A2(_3217_),
    .Y(_3218_),
    .B1(net1864));
 sg13g2_a21oi_1 _7663_ (.A1(_1623_),
    .A2(_1966_),
    .Y(_3219_),
    .B1(net1851));
 sg13g2_nor4_1 _7664_ (.A(_1937_),
    .B(_1970_),
    .C(_3126_),
    .D(_3219_),
    .Y(_3220_));
 sg13g2_nor3_1 _7665_ (.A(_3216_),
    .B(_3218_),
    .C(_3220_),
    .Y(_3221_));
 sg13g2_a21oi_1 _7666_ (.A1(net2221),
    .A2(_2966_),
    .Y(_3222_),
    .B1(_2073_));
 sg13g2_o21ai_1 _7667_ (.B1(net2085),
    .Y(_3223_),
    .A1(_1567_),
    .A2(_3222_));
 sg13g2_nor2b_1 _7668_ (.A(_2965_),
    .B_N(_3223_),
    .Y(_3224_));
 sg13g2_a21oi_1 _7669_ (.A1(net2205),
    .A2(_1588_),
    .Y(_3225_),
    .B1(_3211_));
 sg13g2_nor3_1 _7670_ (.A(net1980),
    .B(_2977_),
    .C(_3225_),
    .Y(_3226_));
 sg13g2_o21ai_1 _7671_ (.B1(_1829_),
    .Y(_3227_),
    .A1(_3224_),
    .A2(_3226_));
 sg13g2_a21oi_1 _7672_ (.A1(net2246),
    .A2(_2110_),
    .Y(_3228_),
    .B1(_3044_));
 sg13g2_o21ai_1 _7673_ (.B1(net1829),
    .Y(_3229_),
    .A1(_1648_),
    .A2(_2031_));
 sg13g2_inv_1 _7674_ (.Y(_3230_),
    .A(_3229_));
 sg13g2_nor2_1 _7675_ (.A(_1621_),
    .B(_2069_),
    .Y(_3231_));
 sg13g2_a21oi_1 _7676_ (.A1(_2037_),
    .A2(_3231_),
    .Y(_3232_),
    .B1(net2215));
 sg13g2_a22oi_1 _7677_ (.Y(_3233_),
    .B1(_3230_),
    .B2(net2241),
    .A2(_2182_),
    .A1(net2010));
 sg13g2_a21oi_1 _7678_ (.A1(_3232_),
    .A2(_3233_),
    .Y(_3234_),
    .B1(_3228_));
 sg13g2_nor2_1 _7679_ (.A(net2199),
    .B(_3234_),
    .Y(_3235_));
 sg13g2_nand3_1 _7680_ (.B(_1546_),
    .C(_1691_),
    .A(net2010),
    .Y(_3236_));
 sg13g2_nand3_1 _7681_ (.B(net1875),
    .C(_2036_),
    .A(net1926),
    .Y(_3237_));
 sg13g2_a21oi_1 _7682_ (.A1(_3236_),
    .A2(_3237_),
    .Y(_3238_),
    .B1(net1824));
 sg13g2_o21ai_1 _7683_ (.B1(net1940),
    .Y(_3239_),
    .A1(_3235_),
    .A2(_3238_));
 sg13g2_a21oi_1 _7684_ (.A1(net1856),
    .A2(_2184_),
    .Y(_3240_),
    .B1(_3183_));
 sg13g2_nor2_1 _7685_ (.A(net2215),
    .B(_3240_),
    .Y(_3241_));
 sg13g2_nand3_1 _7686_ (.B(net1895),
    .C(_2182_),
    .A(net2215),
    .Y(_3242_));
 sg13g2_a21oi_2 _7687_ (.B1(_2466_),
    .Y(_3243_),
    .A2(net1868),
    .A1(net2259));
 sg13g2_o21ai_1 _7688_ (.B1(_3242_),
    .Y(_3244_),
    .A1(_2109_),
    .A2(_3243_));
 sg13g2_or3_1 _7689_ (.A(_1857_),
    .B(_3241_),
    .C(_3244_),
    .X(_3245_));
 sg13g2_a21oi_2 _7690_ (.B1(_1703_),
    .Y(_3246_),
    .A2(_3245_),
    .A1(_3239_));
 sg13g2_o21ai_1 _7691_ (.B1(_3232_),
    .Y(_3247_),
    .A1(net1926),
    .A2(_2687_));
 sg13g2_a21o_1 _7692_ (.A2(_3058_),
    .A1(net2240),
    .B1(_3247_),
    .X(_3248_));
 sg13g2_o21ai_1 _7693_ (.B1(_3059_),
    .Y(_3249_),
    .A1(_1637_),
    .A2(_1789_));
 sg13g2_nand3_1 _7694_ (.B(_3248_),
    .C(_3249_),
    .A(net2088),
    .Y(_3250_));
 sg13g2_a21oi_1 _7695_ (.A1(net1927),
    .A2(net2006),
    .Y(_3251_),
    .B1(_2017_));
 sg13g2_o21ai_1 _7696_ (.B1(net2199),
    .Y(_3252_),
    .A1(_1655_),
    .A2(_3251_));
 sg13g2_nand4_1 _7697_ (.B(net1771),
    .C(_3250_),
    .A(net1940),
    .Y(_3253_),
    .D(_3252_));
 sg13g2_nand2_2 _7698_ (.Y(_3254_),
    .A(net2264),
    .B(_2840_));
 sg13g2_a21oi_1 _7699_ (.A1(_1810_),
    .A2(_3254_),
    .Y(_3255_),
    .B1(_1556_));
 sg13g2_nor2_1 _7700_ (.A(_1648_),
    .B(_2712_),
    .Y(_3256_));
 sg13g2_o21ai_1 _7701_ (.B1(net1983),
    .Y(_3257_),
    .A1(_3036_),
    .A2(_3256_));
 sg13g2_nor3_1 _7702_ (.A(_3035_),
    .B(_3255_),
    .C(_3257_),
    .Y(_3258_));
 sg13g2_o21ai_1 _7703_ (.B1(_3258_),
    .Y(_3259_),
    .A1(net1942),
    .A2(net2017));
 sg13g2_a21oi_1 _7704_ (.A1(_2388_),
    .A2(_2414_),
    .Y(_3260_),
    .B1(_3075_));
 sg13g2_o21ai_1 _7705_ (.B1(_3260_),
    .Y(_3261_),
    .A1(_2046_),
    .A2(_2195_));
 sg13g2_or4_1 _7706_ (.A(net1934),
    .B(_2946_),
    .C(_3081_),
    .D(_3261_),
    .X(_3262_));
 sg13g2_a21oi_2 _7707_ (.B1(_3078_),
    .Y(_3263_),
    .A2(_3262_),
    .A1(_3259_));
 sg13g2_o21ai_1 _7708_ (.B1(_3254_),
    .Y(_3264_),
    .A1(net2258),
    .A2(_1640_));
 sg13g2_a21oi_1 _7709_ (.A1(net2069),
    .A2(_3264_),
    .Y(_3265_),
    .B1(net2203));
 sg13g2_a21oi_1 _7710_ (.A1(_2193_),
    .A2(_3265_),
    .Y(_3266_),
    .B1(net2192));
 sg13g2_a221oi_1 _7711_ (.B2(net1914),
    .C1(net2230),
    .B1(_2705_),
    .A1(net1900),
    .Y(_3267_),
    .A2(_1648_));
 sg13g2_nand2_1 _7712_ (.Y(_3268_),
    .A(net2104),
    .B(_2388_));
 sg13g2_a21o_1 _7713_ (.A2(_3268_),
    .A1(_3179_),
    .B1(net1986),
    .X(_3269_));
 sg13g2_a21oi_1 _7714_ (.A1(_1681_),
    .A2(_2179_),
    .Y(_3270_),
    .B1(net1824));
 sg13g2_nor3_1 _7715_ (.A(net1942),
    .B(net2022),
    .C(net1991),
    .Y(_3271_));
 sg13g2_o21ai_1 _7716_ (.B1(net1983),
    .Y(_3272_),
    .A1(_3267_),
    .A2(_3269_));
 sg13g2_nor4_1 _7717_ (.A(_3266_),
    .B(_3270_),
    .C(_3271_),
    .D(_3272_),
    .Y(_3273_));
 sg13g2_nand2_1 _7718_ (.Y(_3274_),
    .A(net1937),
    .B(_3178_));
 sg13g2_nor4_1 _7719_ (.A(_3175_),
    .B(_3176_),
    .C(_3181_),
    .D(_3274_),
    .Y(_3275_));
 sg13g2_o21ai_1 _7720_ (.B1(_1981_),
    .Y(_3276_),
    .A1(_3273_),
    .A2(_3275_));
 sg13g2_o21ai_1 _7721_ (.B1(_3276_),
    .Y(_3277_),
    .A1(_1858_),
    .A2(_3185_));
 sg13g2_o21ai_1 _7722_ (.B1(_3253_),
    .Y(_3278_),
    .A1(_1861_),
    .A2(_3221_));
 sg13g2_or2_1 _7723_ (.X(_3279_),
    .B(_3278_),
    .A(_3208_));
 sg13g2_nor4_2 _7724_ (.A(_3158_),
    .B(_3246_),
    .C(_3277_),
    .Y(_3280_),
    .D(_3279_));
 sg13g2_a22oi_1 _7725_ (.Y(_3281_),
    .B1(_3263_),
    .B2(net1770),
    .A2(_3195_),
    .A1(_1918_));
 sg13g2_nand4_1 _7726_ (.B(_3227_),
    .C(_3280_),
    .A(_3173_),
    .Y(_3282_),
    .D(_3281_));
 sg13g2_a221oi_1 _7727_ (.B2(net2085),
    .C1(net2184),
    .B1(_3105_),
    .A1(_1675_),
    .Y(_3283_),
    .A2(_2811_));
 sg13g2_a221oi_1 _7728_ (.B2(net1819),
    .C1(_2817_),
    .B1(_1834_),
    .A1(net2221),
    .Y(_3284_),
    .A2(net1885));
 sg13g2_a221oi_1 _7729_ (.B2(net1949),
    .C1(_2855_),
    .B1(_2867_),
    .A1(_1890_),
    .Y(_3285_),
    .A2(_2865_));
 sg13g2_a21oi_1 _7730_ (.A1(_3284_),
    .A2(_3285_),
    .Y(_3286_),
    .B1(net1756));
 sg13g2_o21ai_1 _7731_ (.B1(_3286_),
    .Y(_3287_),
    .A1(_2808_),
    .A2(_3283_));
 sg13g2_nand2_1 _7732_ (.Y(_3288_),
    .A(_3282_),
    .B(_3287_));
 sg13g2_a21oi_1 _7733_ (.A1(_1450_),
    .A2(_3288_),
    .Y(_3289_),
    .B1(\draw_game_inst.board_x[2] ));
 sg13g2_nand3_1 _7734_ (.B(_3143_),
    .C(_3289_),
    .A(_2985_),
    .Y(_3290_));
 sg13g2_a21oi_1 _7735_ (.A1(_1532_),
    .A2(_1614_),
    .Y(_3291_),
    .B1(net1756));
 sg13g2_a21o_2 _7736_ (.A2(_3290_),
    .A1(_2622_),
    .B1(_3291_),
    .X(_3292_));
 sg13g2_nor2_1 _7737_ (.A(_1485_),
    .B(_3292_),
    .Y(_3293_));
 sg13g2_a22oi_1 _7738_ (.Y(_3294_),
    .B1(\draw_game_inst.new_tiles[11] ),
    .B2(net2276),
    .A2(\draw_game_inst.new_tiles[10] ),
    .A1(net2280));
 sg13g2_a22oi_1 _7739_ (.Y(_3295_),
    .B1(net2021),
    .B2(\draw_game_inst.new_tiles[9] ),
    .A2(net2023),
    .A1(\draw_game_inst.new_tiles[8] ));
 sg13g2_o21ai_1 _7740_ (.B1(_3295_),
    .Y(_3296_),
    .A1(net2023),
    .A2(_3294_));
 sg13g2_nand2_1 _7741_ (.Y(_3297_),
    .A(_1486_),
    .B(_3296_));
 sg13g2_a22oi_1 _7742_ (.Y(_3298_),
    .B1(\draw_game_inst.new_tiles[7] ),
    .B2(net2276),
    .A2(\draw_game_inst.new_tiles[6] ),
    .A1(net2280));
 sg13g2_a22oi_1 _7743_ (.Y(_3299_),
    .B1(net2021),
    .B2(\draw_game_inst.new_tiles[5] ),
    .A2(net2023),
    .A1(\draw_game_inst.new_tiles[4] ));
 sg13g2_o21ai_1 _7744_ (.B1(_3299_),
    .Y(_3300_),
    .A1(net2023),
    .A2(_3298_));
 sg13g2_a22oi_1 _7745_ (.Y(_3301_),
    .B1(\draw_game_inst.new_tiles[3] ),
    .B2(net2276),
    .A2(\draw_game_inst.new_tiles[2] ),
    .A1(net2280));
 sg13g2_a22oi_1 _7746_ (.Y(_3302_),
    .B1(net2021),
    .B2(\draw_game_inst.new_tiles[1] ),
    .A2(net2023),
    .A1(\draw_game_inst.new_tiles[0] ));
 sg13g2_o21ai_1 _7747_ (.B1(_3302_),
    .Y(_3303_),
    .A1(net2023),
    .A2(_3301_));
 sg13g2_nand2b_1 _7748_ (.Y(_3304_),
    .B(_3303_),
    .A_N(_1480_));
 sg13g2_a22oi_1 _7749_ (.Y(_3305_),
    .B1(\draw_game_inst.new_tiles[15] ),
    .B2(net2276),
    .A2(\draw_game_inst.new_tiles[14] ),
    .A1(net2280));
 sg13g2_a22oi_1 _7750_ (.Y(_3306_),
    .B1(net2021),
    .B2(\draw_game_inst.new_tiles[13] ),
    .A2(net2023),
    .A1(\draw_game_inst.new_tiles[12] ));
 sg13g2_o21ai_1 _7751_ (.B1(_3306_),
    .Y(_3307_),
    .A1(net2023),
    .A2(_3305_));
 sg13g2_a22oi_1 _7752_ (.Y(_3308_),
    .B1(_3307_),
    .B2(_1490_),
    .A2(_3300_),
    .A1(net2031));
 sg13g2_nand3_1 _7753_ (.B(_3304_),
    .C(_3308_),
    .A(_3297_),
    .Y(_3309_));
 sg13g2_inv_1 _7754_ (.Y(_3310_),
    .A(_3309_));
 sg13g2_nor2_1 _7755_ (.A(\draw_game_inst.new_tiles_counter[0] ),
    .B(\draw_game_inst.new_tiles_counter[1] ),
    .Y(_3311_));
 sg13g2_a21oi_2 _7756_ (.B1(_3310_),
    .Y(_3312_),
    .A2(_3311_),
    .A1(net451));
 sg13g2_a21oi_2 _7757_ (.B1(_4008_),
    .Y(_3313_),
    .A2(net5),
    .A1(net6));
 sg13g2_mux2_1 _7758_ (.A0(_3313_),
    .A1(net479),
    .S(_3312_),
    .X(_3314_));
 sg13g2_nand2_1 _7759_ (.Y(_3315_),
    .A(net8),
    .B(\draw_game_inst.board_y[4] ));
 sg13g2_nor3_1 _7760_ (.A(\draw_game_inst.x[9] ),
    .B(net2179),
    .C(_3315_),
    .Y(_3316_));
 sg13g2_nand4_1 _7761_ (.B(_1482_),
    .C(_1486_),
    .A(_1470_),
    .Y(_3317_),
    .D(_3316_));
 sg13g2_nor2b_2 _7762_ (.A(_3317_),
    .B_N(_1485_),
    .Y(_3318_));
 sg13g2_nor2b_1 _7763_ (.A(_1485_),
    .B_N(_3292_),
    .Y(_3319_));
 sg13g2_inv_1 _7764_ (.Y(_3320_),
    .A(_3319_));
 sg13g2_nand3_1 _7765_ (.B(net1890),
    .C(net1883),
    .A(_1575_),
    .Y(_3321_));
 sg13g2_nor4_2 _7766_ (.A(\draw_game_inst.board_x[0] ),
    .B(\draw_game_inst.board_x[1] ),
    .C(\draw_game_inst.board_x[2] ),
    .Y(_3322_),
    .D(_1721_));
 sg13g2_nand2_1 _7767_ (.Y(_3323_),
    .A(_1479_),
    .B(_3321_));
 sg13g2_or3_1 _7768_ (.A(_1462_),
    .B(_3322_),
    .C(_3323_),
    .X(_3324_));
 sg13g2_and3_1 _7769_ (.X(_3325_),
    .A(_3313_),
    .B(_3319_),
    .C(_3324_));
 sg13g2_inv_1 _7770_ (.Y(_3326_),
    .A(_3325_));
 sg13g2_a22oi_1 _7771_ (.Y(_3327_),
    .B1(_3318_),
    .B2(net2296),
    .A2(_3314_),
    .A1(_3293_));
 sg13g2_a21oi_1 _7772_ (.A1(_3326_),
    .A2(_3327_),
    .Y(_0186_),
    .B1(_1473_));
 sg13g2_o21ai_1 _7773_ (.B1(_3293_),
    .Y(_3328_),
    .A1(_4054_),
    .A2(_3310_));
 sg13g2_a21oi_1 _7774_ (.A1(net2291),
    .A2(_3318_),
    .Y(_3329_),
    .B1(_3325_));
 sg13g2_a21oi_1 _7775_ (.A1(_3328_),
    .A2(_3329_),
    .Y(_0187_),
    .B1(_1473_));
 sg13g2_nor2_1 _7776_ (.A(_3320_),
    .B(_3324_),
    .Y(_3330_));
 sg13g2_nand3b_1 _7777_ (.B(_3330_),
    .C(\draw_game_inst.board_x[0] ),
    .Y(_3331_),
    .A_N(_3313_));
 sg13g2_nand2_1 _7778_ (.Y(_3332_),
    .A(net1009),
    .B(_3312_));
 sg13g2_a221oi_1 _7779_ (.B2(_3293_),
    .C1(_3325_),
    .B1(_3332_),
    .A1(net2286),
    .Y(_3333_),
    .A2(_3318_));
 sg13g2_a21oi_1 _7780_ (.A1(_3331_),
    .A2(_3333_),
    .Y(_0188_),
    .B1(net985));
 sg13g2_or2_1 _7781_ (.X(_3334_),
    .B(_3317_),
    .A(_4049_));
 sg13g2_a21oi_1 _7782_ (.A1(_1485_),
    .A2(_3334_),
    .Y(_3335_),
    .B1(_1473_));
 sg13g2_nor2b_1 _7783_ (.A(_3330_),
    .B_N(_3335_),
    .Y(_0189_));
 sg13g2_a21oi_1 _7784_ (.A1(net2278),
    .A2(_3318_),
    .Y(_3336_),
    .B1(_3325_));
 sg13g2_nor2_1 _7785_ (.A(_1473_),
    .B(_3336_),
    .Y(_0190_));
 sg13g2_or4_1 _7786_ (.A(_1485_),
    .B(_3292_),
    .C(_3312_),
    .D(_3313_),
    .X(_3337_));
 sg13g2_a21oi_1 _7787_ (.A1(net972),
    .A2(_3318_),
    .Y(_3338_),
    .B1(_3325_));
 sg13g2_a21oi_1 _7788_ (.A1(_3337_),
    .A2(_3338_),
    .Y(_0191_),
    .B1(_1473_));
 sg13g2_nor2b_2 _7789_ (.A(vsync_prev),
    .B_N(\vga_sync_gen.vsync ),
    .Y(_3339_));
 sg13g2_nand2b_1 _7790_ (.Y(_3340_),
    .B(\vga_sync_gen.vsync ),
    .A_N(vsync_prev));
 sg13g2_o21ai_1 _7791_ (.B1(net1971),
    .Y(_3341_),
    .A1(_3990_),
    .A2(net2115));
 sg13g2_a21oi_1 _7792_ (.A1(net2115),
    .A2(\debug_controller_inst.grid_in[0] ),
    .Y(_3342_),
    .B1(_3341_));
 sg13g2_o21ai_1 _7793_ (.B1(net2333),
    .Y(_3343_),
    .A1(net703),
    .A2(net1971));
 sg13g2_nor2_1 _7794_ (.A(_3342_),
    .B(_3343_),
    .Y(_0192_));
 sg13g2_a21oi_1 _7795_ (.A1(net2115),
    .A2(\debug_controller_inst.grid_in[1] ),
    .Y(_3344_),
    .B1(_3341_));
 sg13g2_o21ai_1 _7796_ (.B1(net2327),
    .Y(_3345_),
    .A1(net746),
    .A2(net1971));
 sg13g2_nor2_1 _7797_ (.A(_3344_),
    .B(_3345_),
    .Y(_0193_));
 sg13g2_a21oi_1 _7798_ (.A1(net2118),
    .A2(\debug_controller_inst.grid_in[2] ),
    .Y(_3346_),
    .B1(net1964));
 sg13g2_o21ai_1 _7799_ (.B1(net2317),
    .Y(_3347_),
    .A1(net727),
    .A2(net1975));
 sg13g2_nor2_1 _7800_ (.A(_3346_),
    .B(_3347_),
    .Y(_0194_));
 sg13g2_a21oi_1 _7801_ (.A1(net2121),
    .A2(\debug_controller_inst.grid_in[3] ),
    .Y(_3348_),
    .B1(_3341_));
 sg13g2_o21ai_1 _7802_ (.B1(net2333),
    .Y(_3349_),
    .A1(net653),
    .A2(net1973));
 sg13g2_nor2_1 _7803_ (.A(_3348_),
    .B(_3349_),
    .Y(_0195_));
 sg13g2_a21o_2 _7804_ (.A2(net2274),
    .A1(net642),
    .B1(net1961),
    .X(_3350_));
 sg13g2_a21oi_1 _7805_ (.A1(net2115),
    .A2(\debug_controller_inst.grid_in[4] ),
    .Y(_3351_),
    .B1(_3350_));
 sg13g2_o21ai_1 _7806_ (.B1(net2333),
    .Y(_3352_),
    .A1(net694),
    .A2(net1973));
 sg13g2_nor2_1 _7807_ (.A(_3351_),
    .B(_3352_),
    .Y(_0196_));
 sg13g2_a21oi_1 _7808_ (.A1(net2115),
    .A2(\debug_controller_inst.grid_in[5] ),
    .Y(_3353_),
    .B1(_3350_));
 sg13g2_o21ai_1 _7809_ (.B1(net2333),
    .Y(_3354_),
    .A1(net781),
    .A2(net1971));
 sg13g2_nor2_1 _7810_ (.A(_3353_),
    .B(_3354_),
    .Y(_0197_));
 sg13g2_a21oi_1 _7811_ (.A1(net2117),
    .A2(\debug_controller_inst.grid_in[6] ),
    .Y(_3355_),
    .B1(net1964));
 sg13g2_o21ai_1 _7812_ (.B1(net2317),
    .Y(_3356_),
    .A1(net705),
    .A2(net1974));
 sg13g2_nor2_1 _7813_ (.A(_3355_),
    .B(_3356_),
    .Y(_0198_));
 sg13g2_a21oi_1 _7814_ (.A1(net2121),
    .A2(\debug_controller_inst.grid_in[7] ),
    .Y(_3357_),
    .B1(_3350_));
 sg13g2_o21ai_1 _7815_ (.B1(net2333),
    .Y(_3358_),
    .A1(net707),
    .A2(net1972));
 sg13g2_nor2_1 _7816_ (.A(_3357_),
    .B(_3358_),
    .Y(_0199_));
 sg13g2_a21o_2 _7817_ (.A2(net2275),
    .A1(net789),
    .B1(net1963),
    .X(_3359_));
 sg13g2_a21oi_1 _7818_ (.A1(net2116),
    .A2(\debug_controller_inst.grid_in[8] ),
    .Y(_3360_),
    .B1(_3359_));
 sg13g2_o21ai_1 _7819_ (.B1(net2327),
    .Y(_3361_),
    .A1(net766),
    .A2(net1972));
 sg13g2_nor2_1 _7820_ (.A(_3360_),
    .B(_3361_),
    .Y(_0200_));
 sg13g2_a21oi_1 _7821_ (.A1(net2114),
    .A2(\debug_controller_inst.grid_in[9] ),
    .Y(_3362_),
    .B1(_3359_));
 sg13g2_o21ai_1 _7822_ (.B1(net2327),
    .Y(_3363_),
    .A1(net853),
    .A2(net1972));
 sg13g2_nor2_1 _7823_ (.A(_3362_),
    .B(_3363_),
    .Y(_0201_));
 sg13g2_a21oi_1 _7824_ (.A1(net2117),
    .A2(\debug_controller_inst.grid_in[10] ),
    .Y(_3364_),
    .B1(net1964));
 sg13g2_o21ai_1 _7825_ (.B1(net2318),
    .Y(_3365_),
    .A1(net852),
    .A2(net1975));
 sg13g2_nor2_1 _7826_ (.A(_3364_),
    .B(_3365_),
    .Y(_0202_));
 sg13g2_a21oi_1 _7827_ (.A1(net2116),
    .A2(\debug_controller_inst.grid_in[11] ),
    .Y(_3366_),
    .B1(_3359_));
 sg13g2_o21ai_1 _7828_ (.B1(net2333),
    .Y(_3367_),
    .A1(net661),
    .A2(net1972));
 sg13g2_nor2_1 _7829_ (.A(_3366_),
    .B(_3367_),
    .Y(_0203_));
 sg13g2_a21o_2 _7830_ (.A2(net2275),
    .A1(net812),
    .B1(net1963),
    .X(_3368_));
 sg13g2_a21oi_1 _7831_ (.A1(net2116),
    .A2(\debug_controller_inst.grid_in[12] ),
    .Y(_3369_),
    .B1(_3368_));
 sg13g2_o21ai_1 _7832_ (.B1(net2316),
    .Y(_3370_),
    .A1(net748),
    .A2(net1972));
 sg13g2_nor2_1 _7833_ (.A(_3369_),
    .B(_3370_),
    .Y(_0204_));
 sg13g2_a21oi_1 _7834_ (.A1(net2116),
    .A2(\debug_controller_inst.grid_in[13] ),
    .Y(_3371_),
    .B1(_3368_));
 sg13g2_o21ai_1 _7835_ (.B1(net2327),
    .Y(_3372_),
    .A1(net814),
    .A2(net1972));
 sg13g2_nor2_1 _7836_ (.A(_3371_),
    .B(_3372_),
    .Y(_0205_));
 sg13g2_a21oi_1 _7837_ (.A1(net2117),
    .A2(\debug_controller_inst.grid_in[14] ),
    .Y(_3373_),
    .B1(net1965));
 sg13g2_o21ai_1 _7838_ (.B1(net2318),
    .Y(_3374_),
    .A1(net721),
    .A2(net1975));
 sg13g2_nor2_1 _7839_ (.A(_3373_),
    .B(_3374_),
    .Y(_0206_));
 sg13g2_a21oi_1 _7840_ (.A1(net2116),
    .A2(\debug_controller_inst.grid_in[15] ),
    .Y(_3375_),
    .B1(_3368_));
 sg13g2_o21ai_1 _7841_ (.B1(net2320),
    .Y(_3376_),
    .A1(net669),
    .A2(net1972));
 sg13g2_nor2_1 _7842_ (.A(_3375_),
    .B(_3376_),
    .Y(_0207_));
 sg13g2_a21o_2 _7843_ (.A2(net2273),
    .A1(net656),
    .B1(net1961),
    .X(_3377_));
 sg13g2_a21oi_1 _7844_ (.A1(net2121),
    .A2(\debug_controller_inst.grid_in[16] ),
    .Y(_3378_),
    .B1(_3377_));
 sg13g2_o21ai_1 _7845_ (.B1(net2320),
    .Y(_3379_),
    .A1(net795),
    .A2(net1978));
 sg13g2_nor2_1 _7846_ (.A(_3378_),
    .B(_3379_),
    .Y(_0208_));
 sg13g2_a21oi_1 _7847_ (.A1(net2121),
    .A2(\debug_controller_inst.grid_in[17] ),
    .Y(_3380_),
    .B1(_3377_));
 sg13g2_o21ai_1 _7848_ (.B1(net2333),
    .Y(_3381_),
    .A1(net762),
    .A2(net1978));
 sg13g2_nor2_1 _7849_ (.A(_3380_),
    .B(_3381_),
    .Y(_0209_));
 sg13g2_a21oi_1 _7850_ (.A1(net2119),
    .A2(\debug_controller_inst.grid_in[18] ),
    .Y(_3382_),
    .B1(net1966));
 sg13g2_o21ai_1 _7851_ (.B1(net2322),
    .Y(_3383_),
    .A1(net734),
    .A2(net1976));
 sg13g2_nor2_1 _7852_ (.A(_3382_),
    .B(_3383_),
    .Y(_0210_));
 sg13g2_a21oi_1 _7853_ (.A1(net2120),
    .A2(\debug_controller_inst.grid_in[19] ),
    .Y(_3384_),
    .B1(_3377_));
 sg13g2_o21ai_1 _7854_ (.B1(net2320),
    .Y(_3385_),
    .A1(net685),
    .A2(net1977));
 sg13g2_nor2_1 _7855_ (.A(_3384_),
    .B(_3385_),
    .Y(_0211_));
 sg13g2_a21o_2 _7856_ (.A2(net2273),
    .A1(\welcome_screen_grid[20] ),
    .B1(net1962),
    .X(_3386_));
 sg13g2_a21oi_1 _7857_ (.A1(net2120),
    .A2(\debug_controller_inst.grid_in[20] ),
    .Y(_3387_),
    .B1(_3386_));
 sg13g2_o21ai_1 _7858_ (.B1(net2320),
    .Y(_3388_),
    .A1(net759),
    .A2(net1978));
 sg13g2_nor2_1 _7859_ (.A(_3387_),
    .B(_3388_),
    .Y(_0212_));
 sg13g2_a21oi_1 _7860_ (.A1(net2120),
    .A2(\debug_controller_inst.grid_in[21] ),
    .Y(_3389_),
    .B1(_3386_));
 sg13g2_o21ai_1 _7861_ (.B1(net2334),
    .Y(_3390_),
    .A1(net775),
    .A2(net1978));
 sg13g2_nor2_1 _7862_ (.A(_3389_),
    .B(_3390_),
    .Y(_0213_));
 sg13g2_a21oi_1 _7863_ (.A1(net2119),
    .A2(\debug_controller_inst.grid_in[22] ),
    .Y(_3391_),
    .B1(net1966));
 sg13g2_o21ai_1 _7864_ (.B1(net2322),
    .Y(_3392_),
    .A1(net683),
    .A2(net1976));
 sg13g2_nor2_1 _7865_ (.A(_3391_),
    .B(_3392_),
    .Y(_0214_));
 sg13g2_a21oi_1 _7866_ (.A1(net2120),
    .A2(\debug_controller_inst.grid_in[23] ),
    .Y(_3393_),
    .B1(_3386_));
 sg13g2_o21ai_1 _7867_ (.B1(net2320),
    .Y(_3394_),
    .A1(net785),
    .A2(net1977));
 sg13g2_nor2_1 _7868_ (.A(_3393_),
    .B(_3394_),
    .Y(_0215_));
 sg13g2_a21o_2 _7869_ (.A2(net2273),
    .A1(\welcome_screen_grid[24] ),
    .B1(net1962),
    .X(_3395_));
 sg13g2_a21oi_1 _7870_ (.A1(net2120),
    .A2(\debug_controller_inst.grid_in[24] ),
    .Y(_3396_),
    .B1(_3395_));
 sg13g2_o21ai_1 _7871_ (.B1(net2324),
    .Y(_3397_),
    .A1(net701),
    .A2(net1977));
 sg13g2_nor2_1 _7872_ (.A(_3396_),
    .B(_3397_),
    .Y(_0216_));
 sg13g2_a21oi_1 _7873_ (.A1(net2121),
    .A2(\debug_controller_inst.grid_in[25] ),
    .Y(_3398_),
    .B1(_3395_));
 sg13g2_o21ai_1 _7874_ (.B1(net2334),
    .Y(_3399_),
    .A1(net779),
    .A2(net1977));
 sg13g2_nor2_1 _7875_ (.A(_3398_),
    .B(_3399_),
    .Y(_0217_));
 sg13g2_a21oi_1 _7876_ (.A1(net2119),
    .A2(\debug_controller_inst.grid_in[26] ),
    .Y(_3400_),
    .B1(net1967));
 sg13g2_o21ai_1 _7877_ (.B1(net2322),
    .Y(_3401_),
    .A1(net719),
    .A2(net1979));
 sg13g2_nor2_1 _7878_ (.A(_3400_),
    .B(_3401_),
    .Y(_0218_));
 sg13g2_a21oi_1 _7879_ (.A1(net2121),
    .A2(\debug_controller_inst.grid_in[27] ),
    .Y(_3402_),
    .B1(_3395_));
 sg13g2_o21ai_1 _7880_ (.B1(net2320),
    .Y(_3403_),
    .A1(net750),
    .A2(net1977));
 sg13g2_nor2_1 _7881_ (.A(_3402_),
    .B(_3403_),
    .Y(_0219_));
 sg13g2_a21o_2 _7882_ (.A2(net2273),
    .A1(\welcome_screen_grid[28] ),
    .B1(net1962),
    .X(_3404_));
 sg13g2_a21oi_1 _7883_ (.A1(net2120),
    .A2(\debug_controller_inst.grid_in[28] ),
    .Y(_3405_),
    .B1(_3404_));
 sg13g2_o21ai_1 _7884_ (.B1(net2320),
    .Y(_3406_),
    .A1(net699),
    .A2(net1977));
 sg13g2_nor2_1 _7885_ (.A(_3405_),
    .B(_3406_),
    .Y(_0220_));
 sg13g2_a21oi_1 _7886_ (.A1(net2120),
    .A2(\debug_controller_inst.grid_in[29] ),
    .Y(_3407_),
    .B1(_3404_));
 sg13g2_o21ai_1 _7887_ (.B1(net2334),
    .Y(_3408_),
    .A1(net768),
    .A2(net1977));
 sg13g2_nor2_1 _7888_ (.A(_3407_),
    .B(_3408_),
    .Y(_0221_));
 sg13g2_a21oi_1 _7889_ (.A1(net2119),
    .A2(\debug_controller_inst.grid_in[30] ),
    .Y(_3409_),
    .B1(net1967));
 sg13g2_o21ai_1 _7890_ (.B1(net2321),
    .Y(_3410_),
    .A1(net831),
    .A2(net1979));
 sg13g2_nor2_1 _7891_ (.A(_3409_),
    .B(_3410_),
    .Y(_0222_));
 sg13g2_a21oi_1 _7892_ (.A1(net2120),
    .A2(\debug_controller_inst.grid_in[31] ),
    .Y(_3411_),
    .B1(_3404_));
 sg13g2_o21ai_1 _7893_ (.B1(net2320),
    .Y(_3412_),
    .A1(net692),
    .A2(net1977));
 sg13g2_nor2_1 _7894_ (.A(_3411_),
    .B(_3412_),
    .Y(_0223_));
 sg13g2_o21ai_1 _7895_ (.B1(net1968),
    .Y(_3413_),
    .A1(_3989_),
    .A2(net2111));
 sg13g2_a21oi_1 _7896_ (.A1(net2111),
    .A2(\debug_controller_inst.grid_in[32] ),
    .Y(_3414_),
    .B1(_3413_));
 sg13g2_o21ai_1 _7897_ (.B1(net2328),
    .Y(_3415_),
    .A1(net824),
    .A2(net1968));
 sg13g2_nor2_1 _7898_ (.A(_3414_),
    .B(_3415_),
    .Y(_0224_));
 sg13g2_a21oi_1 _7899_ (.A1(net2111),
    .A2(\debug_controller_inst.grid_in[33] ),
    .Y(_3416_),
    .B1(_3413_));
 sg13g2_o21ai_1 _7900_ (.B1(net2329),
    .Y(_3417_),
    .A1(net761),
    .A2(net1970));
 sg13g2_nor2_1 _7901_ (.A(_3416_),
    .B(_3417_),
    .Y(_0225_));
 sg13g2_a21oi_1 _7902_ (.A1(net2117),
    .A2(\debug_controller_inst.grid_in[34] ),
    .Y(_3418_),
    .B1(net1964));
 sg13g2_o21ai_1 _7903_ (.B1(net2317),
    .Y(_3419_),
    .A1(net709),
    .A2(net1974));
 sg13g2_nor2_1 _7904_ (.A(_3418_),
    .B(_3419_),
    .Y(_0226_));
 sg13g2_a21oi_1 _7905_ (.A1(net2111),
    .A2(\debug_controller_inst.grid_in[35] ),
    .Y(_3420_),
    .B1(_3413_));
 sg13g2_o21ai_1 _7906_ (.B1(net2328),
    .Y(_3421_),
    .A1(net744),
    .A2(net1968));
 sg13g2_nor2_1 _7907_ (.A(_3420_),
    .B(_3421_),
    .Y(_0227_));
 sg13g2_a21o_1 _7908_ (.A2(net2274),
    .A1(net733),
    .B1(net1961),
    .X(_3422_));
 sg13g2_a21oi_1 _7909_ (.A1(net2113),
    .A2(\debug_controller_inst.grid_in[36] ),
    .Y(_3423_),
    .B1(_3422_));
 sg13g2_o21ai_1 _7910_ (.B1(net2328),
    .Y(_3424_),
    .A1(net752),
    .A2(net1968));
 sg13g2_nor2_1 _7911_ (.A(_3423_),
    .B(_3424_),
    .Y(_0228_));
 sg13g2_a21oi_1 _7912_ (.A1(net2112),
    .A2(\debug_controller_inst.grid_in[37] ),
    .Y(_3425_),
    .B1(_3422_));
 sg13g2_o21ai_1 _7913_ (.B1(net2328),
    .Y(_3426_),
    .A1(net777),
    .A2(net1969));
 sg13g2_nor2_1 _7914_ (.A(_3425_),
    .B(_3426_),
    .Y(_0229_));
 sg13g2_a21oi_1 _7915_ (.A1(net2117),
    .A2(\debug_controller_inst.grid_in[38] ),
    .Y(_3427_),
    .B1(net1964));
 sg13g2_o21ai_1 _7916_ (.B1(net2317),
    .Y(_3428_),
    .A1(net834),
    .A2(net1974));
 sg13g2_nor2_1 _7917_ (.A(_3427_),
    .B(_3428_),
    .Y(_0230_));
 sg13g2_a21oi_1 _7918_ (.A1(net2114),
    .A2(\debug_controller_inst.grid_in[39] ),
    .Y(_3429_),
    .B1(_3422_));
 sg13g2_o21ai_1 _7919_ (.B1(net2328),
    .Y(_3430_),
    .A1(net729),
    .A2(net1973));
 sg13g2_nor2_1 _7920_ (.A(_3429_),
    .B(_3430_),
    .Y(_0231_));
 sg13g2_a21o_1 _7921_ (.A2(net2275),
    .A1(net758),
    .B1(net1961),
    .X(_3431_));
 sg13g2_a21oi_1 _7922_ (.A1(net2113),
    .A2(\debug_controller_inst.grid_in[40] ),
    .Y(_3432_),
    .B1(_3431_));
 sg13g2_o21ai_1 _7923_ (.B1(net2314),
    .Y(_3433_),
    .A1(net798),
    .A2(net1968));
 sg13g2_nor2_1 _7924_ (.A(_3432_),
    .B(_3433_),
    .Y(_0232_));
 sg13g2_a21oi_1 _7925_ (.A1(net2111),
    .A2(\debug_controller_inst.grid_in[41] ),
    .Y(_3434_),
    .B1(_3431_));
 sg13g2_o21ai_1 _7926_ (.B1(net2328),
    .Y(_3435_),
    .A1(net805),
    .A2(net1970));
 sg13g2_nor2_1 _7927_ (.A(_3434_),
    .B(_3435_),
    .Y(_0233_));
 sg13g2_a21oi_1 _7928_ (.A1(net2117),
    .A2(\debug_controller_inst.grid_in[42] ),
    .Y(_3436_),
    .B1(net1964));
 sg13g2_o21ai_1 _7929_ (.B1(net2317),
    .Y(_3437_),
    .A1(net674),
    .A2(net1975));
 sg13g2_nor2_1 _7930_ (.A(_3436_),
    .B(_3437_),
    .Y(_0234_));
 sg13g2_a21oi_1 _7931_ (.A1(net2113),
    .A2(\debug_controller_inst.grid_in[43] ),
    .Y(_3438_),
    .B1(_3431_));
 sg13g2_o21ai_1 _7932_ (.B1(net2314),
    .Y(_3439_),
    .A1(net821),
    .A2(net1968));
 sg13g2_nor2_1 _7933_ (.A(_3438_),
    .B(_3439_),
    .Y(_0235_));
 sg13g2_a21o_1 _7934_ (.A2(net2273),
    .A1(net647),
    .B1(net1961),
    .X(_3440_));
 sg13g2_a21oi_1 _7935_ (.A1(net2113),
    .A2(\debug_controller_inst.grid_in[44] ),
    .Y(_3441_),
    .B1(_3440_));
 sg13g2_o21ai_1 _7936_ (.B1(net2316),
    .Y(_3442_),
    .A1(net793),
    .A2(net1968));
 sg13g2_nor2_1 _7937_ (.A(_3441_),
    .B(_3442_),
    .Y(_0236_));
 sg13g2_a21oi_1 _7938_ (.A1(net2111),
    .A2(\debug_controller_inst.grid_in[45] ),
    .Y(_3443_),
    .B1(_3440_));
 sg13g2_o21ai_1 _7939_ (.B1(net2328),
    .Y(_3444_),
    .A1(net808),
    .A2(net1970));
 sg13g2_nor2_1 _7940_ (.A(_3443_),
    .B(_3444_),
    .Y(_0237_));
 sg13g2_a21oi_1 _7941_ (.A1(net2117),
    .A2(\debug_controller_inst.grid_in[46] ),
    .Y(_3445_),
    .B1(net1964));
 sg13g2_o21ai_1 _7942_ (.B1(net2317),
    .Y(_3446_),
    .A1(net696),
    .A2(net1974));
 sg13g2_nor2_1 _7943_ (.A(_3445_),
    .B(_3446_),
    .Y(_0238_));
 sg13g2_a21oi_1 _7944_ (.A1(net2113),
    .A2(\debug_controller_inst.grid_in[47] ),
    .Y(_3447_),
    .B1(_3440_));
 sg13g2_o21ai_1 _7945_ (.B1(net2316),
    .Y(_3448_),
    .A1(net764),
    .A2(net1968));
 sg13g2_nor2_1 _7946_ (.A(_3447_),
    .B(_3448_),
    .Y(_0239_));
 sg13g2_a21o_1 _7947_ (.A2(net2273),
    .A1(net621),
    .B1(net1961),
    .X(_3449_));
 sg13g2_a21oi_1 _7948_ (.A1(net2114),
    .A2(\debug_controller_inst.grid_in[48] ),
    .Y(_3450_),
    .B1(_3449_));
 sg13g2_o21ai_1 _7949_ (.B1(net2330),
    .Y(_3451_),
    .A1(net688),
    .A2(net1969));
 sg13g2_nor2_1 _7950_ (.A(_3450_),
    .B(_3451_),
    .Y(_0240_));
 sg13g2_a21oi_1 _7951_ (.A1(net2114),
    .A2(\debug_controller_inst.grid_in[49] ),
    .Y(_3452_),
    .B1(_3449_));
 sg13g2_o21ai_1 _7952_ (.B1(net2330),
    .Y(_3453_),
    .A1(net826),
    .A2(net1971));
 sg13g2_nor2_1 _7953_ (.A(_3452_),
    .B(_3453_),
    .Y(_0241_));
 sg13g2_a21oi_1 _7954_ (.A1(net2118),
    .A2(\debug_controller_inst.grid_in[50] ),
    .Y(_3454_),
    .B1(net1965));
 sg13g2_o21ai_1 _7955_ (.B1(net2322),
    .Y(_3455_),
    .A1(net783),
    .A2(net1974));
 sg13g2_nor2_1 _7956_ (.A(_3454_),
    .B(_3455_),
    .Y(_0242_));
 sg13g2_a21oi_1 _7957_ (.A1(net2114),
    .A2(\debug_controller_inst.grid_in[51] ),
    .Y(_3456_),
    .B1(_3449_));
 sg13g2_o21ai_1 _7958_ (.B1(net2327),
    .Y(_3457_),
    .A1(net651),
    .A2(net1971));
 sg13g2_nor2_1 _7959_ (.A(_3456_),
    .B(_3457_),
    .Y(_0243_));
 sg13g2_a21o_1 _7960_ (.A2(net2273),
    .A1(net636),
    .B1(net1962),
    .X(_3458_));
 sg13g2_a21oi_1 _7961_ (.A1(net2114),
    .A2(\debug_controller_inst.grid_in[52] ),
    .Y(_3459_),
    .B1(_3458_));
 sg13g2_o21ai_1 _7962_ (.B1(net2327),
    .Y(_3460_),
    .A1(net754),
    .A2(net1969));
 sg13g2_nor2_1 _7963_ (.A(_3459_),
    .B(_3460_),
    .Y(_0244_));
 sg13g2_a21oi_1 _7964_ (.A1(net2114),
    .A2(\debug_controller_inst.grid_in[53] ),
    .Y(_3461_),
    .B1(_3458_));
 sg13g2_o21ai_1 _7965_ (.B1(net2329),
    .Y(_3462_),
    .A1(net680),
    .A2(net1971));
 sg13g2_nor2_1 _7966_ (.A(_3461_),
    .B(_3462_),
    .Y(_0245_));
 sg13g2_a21oi_1 _7967_ (.A1(net2119),
    .A2(\debug_controller_inst.grid_in[54] ),
    .Y(_3463_),
    .B1(net1965));
 sg13g2_o21ai_1 _7968_ (.B1(net2322),
    .Y(_3464_),
    .A1(net818),
    .A2(net1974));
 sg13g2_nor2_1 _7969_ (.A(_3463_),
    .B(_3464_),
    .Y(_0246_));
 sg13g2_a21oi_1 _7970_ (.A1(net2114),
    .A2(\debug_controller_inst.grid_in[55] ),
    .Y(_3465_),
    .B1(_3458_));
 sg13g2_o21ai_1 _7971_ (.B1(net2327),
    .Y(_3466_),
    .A1(net773),
    .A2(net1971));
 sg13g2_nor2_1 _7972_ (.A(_3465_),
    .B(_3466_),
    .Y(_0247_));
 sg13g2_a21o_1 _7973_ (.A2(net2273),
    .A1(net613),
    .B1(net1961),
    .X(_3467_));
 sg13g2_a21oi_1 _7974_ (.A1(net2112),
    .A2(\debug_controller_inst.grid_in[56] ),
    .Y(_3468_),
    .B1(_3467_));
 sg13g2_o21ai_1 _7975_ (.B1(net2327),
    .Y(_3469_),
    .A1(net717),
    .A2(net1969));
 sg13g2_nor2_1 _7976_ (.A(_3468_),
    .B(_3469_),
    .Y(_0248_));
 sg13g2_a21oi_1 _7977_ (.A1(net2112),
    .A2(\debug_controller_inst.grid_in[57] ),
    .Y(_3470_),
    .B1(_3467_));
 sg13g2_o21ai_1 _7978_ (.B1(net2329),
    .Y(_3471_),
    .A1(net677),
    .A2(net1969));
 sg13g2_nor2_1 _7979_ (.A(_3470_),
    .B(_3471_),
    .Y(_0249_));
 sg13g2_a21oi_1 _7980_ (.A1(net2118),
    .A2(\debug_controller_inst.grid_in[58] ),
    .Y(_3472_),
    .B1(net1964));
 sg13g2_o21ai_1 _7981_ (.B1(net2317),
    .Y(_3473_),
    .A1(net756),
    .A2(net1974));
 sg13g2_nor2_1 _7982_ (.A(_3472_),
    .B(_3473_),
    .Y(_0250_));
 sg13g2_a21oi_1 _7983_ (.A1(net2112),
    .A2(\debug_controller_inst.grid_in[59] ),
    .Y(_3474_),
    .B1(_3467_));
 sg13g2_o21ai_1 _7984_ (.B1(net2329),
    .Y(_3475_),
    .A1(net731),
    .A2(net1969));
 sg13g2_nor2_1 _7985_ (.A(_3474_),
    .B(_3475_),
    .Y(_0251_));
 sg13g2_a21o_1 _7986_ (.A2(net2274),
    .A1(net711),
    .B1(net1962),
    .X(_3476_));
 sg13g2_a21oi_1 _7987_ (.A1(net2112),
    .A2(\debug_controller_inst.grid_in[60] ),
    .Y(_3477_),
    .B1(_3476_));
 sg13g2_o21ai_1 _7988_ (.B1(net2328),
    .Y(_3478_),
    .A1(net637),
    .A2(net1969));
 sg13g2_nor2_1 _7989_ (.A(_3477_),
    .B(_3478_),
    .Y(_0252_));
 sg13g2_a21oi_1 _7990_ (.A1(net2111),
    .A2(\debug_controller_inst.grid_in[61] ),
    .Y(_3479_),
    .B1(_3476_));
 sg13g2_o21ai_1 _7991_ (.B1(net2329),
    .Y(_3480_),
    .A1(net723),
    .A2(net1969));
 sg13g2_nor2_1 _7992_ (.A(_3479_),
    .B(_3480_),
    .Y(_0253_));
 sg13g2_a21oi_1 _7993_ (.A1(net2117),
    .A2(\debug_controller_inst.grid_in[62] ),
    .Y(_3481_),
    .B1(net1965));
 sg13g2_o21ai_1 _7994_ (.B1(net2322),
    .Y(_3482_),
    .A1(net740),
    .A2(net1974));
 sg13g2_nor2_1 _7995_ (.A(_3481_),
    .B(_3482_),
    .Y(_0254_));
 sg13g2_a21oi_1 _7996_ (.A1(net2111),
    .A2(\debug_controller_inst.grid_in[63] ),
    .Y(_3483_),
    .B1(_3476_));
 sg13g2_o21ai_1 _7997_ (.B1(net2329),
    .Y(_3484_),
    .A1(net715),
    .A2(net1970));
 sg13g2_nor2_1 _7998_ (.A(_3483_),
    .B(_3484_),
    .Y(_0255_));
 sg13g2_nand2_2 _7999_ (.Y(_3485_),
    .A(\gamepad_pmod.decoder.data_reg[8] ),
    .B(_0496_));
 sg13g2_nand2b_1 _8000_ (.Y(_3486_),
    .B(_3485_),
    .A_N(_0497_));
 sg13g2_nor4_1 _8001_ (.A(_0499_),
    .B(_0501_),
    .C(_0503_),
    .D(_3486_),
    .Y(_3487_));
 sg13g2_o21ai_1 _8002_ (.B1(net2275),
    .Y(_3488_),
    .A1(net1963),
    .A2(_3487_));
 sg13g2_nand2_1 _8003_ (.Y(_0256_),
    .A(net2315),
    .B(net962));
 sg13g2_nand2_1 _8004_ (.Y(_3489_),
    .A(net559),
    .B(_0496_));
 sg13g2_nor2_1 _8005_ (.A(net2305),
    .B(_3489_),
    .Y(_0257_));
 sg13g2_nor3_1 _8006_ (.A(\draw_game_inst.new_tiles_counter[0] ),
    .B(\new_tiles_counter[0] ),
    .C(\draw_game_inst.new_tiles_counter[1] ),
    .Y(_3490_));
 sg13g2_nand2b_1 _8007_ (.Y(_3491_),
    .B(_3490_),
    .A_N(\draw_game_inst.new_tiles_counter[2] ));
 sg13g2_or2_1 _8008_ (.X(_3492_),
    .B(_3491_),
    .A(\new_tiles_counter[4] ));
 sg13g2_o21ai_1 _8009_ (.B1(net2317),
    .Y(_3493_),
    .A1(net1966),
    .A2(_3492_));
 sg13g2_nor2_1 _8010_ (.A(_4053_),
    .B(net1812),
    .Y(_0258_));
 sg13g2_nor3_1 _8011_ (.A(net2159),
    .B(\game_logic_inst.added_tile_index[1] ),
    .C(_4052_),
    .Y(_3494_));
 sg13g2_nand2_1 _8012_ (.Y(_3495_),
    .A(_4050_),
    .B(_3494_));
 sg13g2_a21oi_1 _8013_ (.A1(net424),
    .A2(_3495_),
    .Y(_0259_),
    .B1(net1811));
 sg13g2_nor3_1 _8014_ (.A(\game_logic_inst.added_tile_index[2] ),
    .B(_4051_),
    .C(\game_logic_inst.added_tile_index[0] ),
    .Y(_3496_));
 sg13g2_nand2_1 _8015_ (.Y(_3497_),
    .A(_4050_),
    .B(_3496_));
 sg13g2_a21oi_1 _8016_ (.A1(net425),
    .A2(_3497_),
    .Y(_0260_),
    .B1(net1811));
 sg13g2_nand2_1 _8017_ (.Y(_3498_),
    .A(\game_logic_inst.added_tile_index[1] ),
    .B(\game_logic_inst.added_tile_index[0] ));
 sg13g2_or3_1 _8018_ (.A(net2158),
    .B(net2159),
    .C(_3498_),
    .X(_3499_));
 sg13g2_a21oi_1 _8019_ (.A1(net437),
    .A2(_3499_),
    .Y(_0261_),
    .B1(net1811));
 sg13g2_nor2_1 _8020_ (.A(\game_logic_inst.added_tile_index[1] ),
    .B(\game_logic_inst.added_tile_index[0] ),
    .Y(_3500_));
 sg13g2_nand3_1 _8021_ (.B(net2159),
    .C(_3500_),
    .A(_4050_),
    .Y(_3501_));
 sg13g2_a21oi_1 _8022_ (.A1(net429),
    .A2(_3501_),
    .Y(_0262_),
    .B1(net1811));
 sg13g2_nand3_1 _8023_ (.B(_4051_),
    .C(\game_logic_inst.added_tile_index[0] ),
    .A(net2159),
    .Y(_3502_));
 sg13g2_o21ai_1 _8024_ (.B1(net481),
    .Y(_3503_),
    .A1(net2158),
    .A2(_3502_));
 sg13g2_nor2b_1 _8025_ (.A(net1812),
    .B_N(_3503_),
    .Y(_0263_));
 sg13g2_nand3_1 _8026_ (.B(\game_logic_inst.added_tile_index[1] ),
    .C(_4052_),
    .A(net2159),
    .Y(_3504_));
 sg13g2_o21ai_1 _8027_ (.B1(net474),
    .Y(_3505_),
    .A1(net2158),
    .A2(_3504_));
 sg13g2_nor2b_1 _8028_ (.A(net1811),
    .B_N(net475),
    .Y(_0264_));
 sg13g2_nand4_1 _8029_ (.B(\game_logic_inst.added_tile_index[2] ),
    .C(\game_logic_inst.added_tile_index[1] ),
    .A(_4050_),
    .Y(_3506_),
    .D(\game_logic_inst.added_tile_index[0] ));
 sg13g2_a21oi_1 _8030_ (.A1(net431),
    .A2(_3506_),
    .Y(_0265_),
    .B1(net1811));
 sg13g2_nor3_1 _8031_ (.A(net2159),
    .B(\game_logic_inst.added_tile_index[1] ),
    .C(\game_logic_inst.added_tile_index[0] ),
    .Y(_3507_));
 sg13g2_nand2_1 _8032_ (.Y(_3508_),
    .A(net2158),
    .B(_3507_));
 sg13g2_a21oi_1 _8033_ (.A1(net418),
    .A2(_3508_),
    .Y(_0266_),
    .B1(net1812));
 sg13g2_nand2_1 _8034_ (.Y(_3509_),
    .A(net2158),
    .B(_3494_));
 sg13g2_a21oi_1 _8035_ (.A1(net427),
    .A2(_3509_),
    .Y(_0267_),
    .B1(net1812));
 sg13g2_nand2_1 _8036_ (.Y(_3510_),
    .A(net2158),
    .B(_3496_));
 sg13g2_a21oi_1 _8037_ (.A1(net420),
    .A2(_3510_),
    .Y(_0268_),
    .B1(net1812));
 sg13g2_or3_1 _8038_ (.A(_4050_),
    .B(net2159),
    .C(_3498_),
    .X(_3511_));
 sg13g2_a21oi_1 _8039_ (.A1(net422),
    .A2(_3511_),
    .Y(_0269_),
    .B1(net1812));
 sg13g2_nand3_1 _8040_ (.B(net2159),
    .C(_3500_),
    .A(net2158),
    .Y(_3512_));
 sg13g2_a21oi_1 _8041_ (.A1(net435),
    .A2(_3512_),
    .Y(_0270_),
    .B1(net1811));
 sg13g2_o21ai_1 _8042_ (.B1(net458),
    .Y(_3513_),
    .A1(_4050_),
    .A2(_3502_));
 sg13g2_nor2b_1 _8043_ (.A(net1811),
    .B_N(_3513_),
    .Y(_0271_));
 sg13g2_o21ai_1 _8044_ (.B1(net463),
    .Y(_3514_),
    .A1(_4050_),
    .A2(_3504_));
 sg13g2_nor2b_1 _8045_ (.A(net1812),
    .B_N(_3514_),
    .Y(_0272_));
 sg13g2_nand4_1 _8046_ (.B(\game_logic_inst.added_tile_index[2] ),
    .C(\game_logic_inst.added_tile_index[1] ),
    .A(\game_logic_inst.added_tile_index[3] ),
    .Y(_3515_),
    .D(\game_logic_inst.added_tile_index[0] ));
 sg13g2_a21oi_1 _8047_ (.A1(net433),
    .A2(_3515_),
    .Y(_0273_),
    .B1(_3493_));
 sg13g2_nand2_1 _8048_ (.Y(_3516_),
    .A(net1976),
    .B(_3492_));
 sg13g2_and2_1 _8049_ (.A(_4050_),
    .B(_3507_),
    .X(_3517_));
 sg13g2_and2_1 _8050_ (.A(_3516_),
    .B(_3517_),
    .X(_3518_));
 sg13g2_o21ai_1 _8051_ (.B1(net2323),
    .Y(_3519_),
    .A1(net445),
    .A2(_3516_));
 sg13g2_a21oi_1 _8052_ (.A1(net445),
    .A2(_3518_),
    .Y(_0274_),
    .B1(_3519_));
 sg13g2_nand2b_1 _8053_ (.Y(_3520_),
    .B(_3518_),
    .A_N(net479));
 sg13g2_xnor2_1 _8054_ (.Y(_3521_),
    .A(\draw_game_inst.new_tiles_counter[0] ),
    .B(\new_tiles_counter[0] ));
 sg13g2_nand3_1 _8055_ (.B(_3492_),
    .C(_3521_),
    .A(net1976),
    .Y(_3522_));
 sg13g2_a21oi_1 _8056_ (.A1(_3520_),
    .A2(_3522_),
    .Y(_0275_),
    .B1(net2307));
 sg13g2_o21ai_1 _8057_ (.B1(\draw_game_inst.new_tiles_counter[1] ),
    .Y(_3523_),
    .A1(\draw_game_inst.new_tiles_counter[0] ),
    .A2(\new_tiles_counter[0] ));
 sg13g2_nor2b_1 _8058_ (.A(_3490_),
    .B_N(_3523_),
    .Y(_3524_));
 sg13g2_nand3_1 _8059_ (.B(net1966),
    .C(_3517_),
    .A(net982),
    .Y(_3525_));
 sg13g2_o21ai_1 _8060_ (.B1(_3525_),
    .Y(_3526_),
    .A1(_3516_),
    .A2(_3524_));
 sg13g2_and2_1 _8061_ (.A(net2323),
    .B(_3526_),
    .X(_0276_));
 sg13g2_nand2b_1 _8062_ (.Y(_3527_),
    .B(\draw_game_inst.new_tiles_counter[2] ),
    .A_N(_3490_));
 sg13g2_and2_1 _8063_ (.A(net1976),
    .B(_3491_),
    .X(_3528_));
 sg13g2_a221oi_1 _8064_ (.B2(_3528_),
    .C1(net2307),
    .B1(_3527_),
    .A1(net451),
    .Y(_0277_),
    .A2(_3518_));
 sg13g2_a21oi_1 _8065_ (.A1(net578),
    .A2(_3491_),
    .Y(_3529_),
    .B1(_3516_));
 sg13g2_nor2b_1 _8066_ (.A(net578),
    .B_N(_3517_),
    .Y(_3530_));
 sg13g2_nor3_1 _8067_ (.A(net2302),
    .B(_3529_),
    .C(_3530_),
    .Y(_0278_));
 sg13g2_nor2_2 _8068_ (.A(btn_select_prev),
    .B(_3489_),
    .Y(_3531_));
 sg13g2_o21ai_1 _8069_ (.B1(net2333),
    .Y(_3532_),
    .A1(retro_colors),
    .A2(_3531_));
 sg13g2_a21oi_1 _8070_ (.A1(_4008_),
    .A2(_3531_),
    .Y(_0279_),
    .B1(_3532_));
 sg13g2_and2_1 _8071_ (.A(net2335),
    .B(net1),
    .X(_0280_));
 sg13g2_xor2_1 _8072_ (.B(\btn_up_debounce.button_sync_1 ),
    .A(net616),
    .X(_3533_));
 sg13g2_nor4_1 _8073_ (.A(\btn_up_debounce.debounce_counter[1] ),
    .B(\btn_up_debounce.debounce_counter[0] ),
    .C(\btn_up_debounce.debounce_counter[3] ),
    .D(\btn_up_debounce.debounce_counter[2] ),
    .Y(_3534_));
 sg13g2_nand3_1 _8074_ (.B(\btn_up_debounce.debounce_counter[16] ),
    .C(_3534_),
    .A(\btn_up_debounce.debounce_counter[15] ),
    .Y(_3535_));
 sg13g2_nand4_1 _8075_ (.B(\btn_up_debounce.debounce_counter[12] ),
    .C(\btn_up_debounce.debounce_counter[14] ),
    .A(_4035_),
    .Y(_3536_),
    .D(\btn_up_debounce.debounce_counter[17] ));
 sg13g2_nor4_1 _8076_ (.A(\btn_up_debounce.debounce_counter[9] ),
    .B(\btn_up_debounce.debounce_counter[8] ),
    .C(\btn_up_debounce.debounce_counter[11] ),
    .D(net544),
    .Y(_3537_));
 sg13g2_nor4_1 _8077_ (.A(\btn_up_debounce.debounce_counter[5] ),
    .B(\btn_up_debounce.debounce_counter[6] ),
    .C(_3535_),
    .D(_3536_),
    .Y(_3538_));
 sg13g2_and4_1 _8078_ (.A(\btn_up_debounce.debounce_counter[4] ),
    .B(net597),
    .C(_3537_),
    .D(_3538_),
    .X(_3539_));
 sg13g2_inv_1 _8079_ (.Y(_3540_),
    .A(_3539_));
 sg13g2_nand3_1 _8080_ (.B(_3533_),
    .C(_3540_),
    .A(net2331),
    .Y(_3541_));
 sg13g2_nor2_1 _8081_ (.A(_4075_),
    .B(net1807),
    .Y(_0281_));
 sg13g2_xnor2_1 _8082_ (.Y(_3542_),
    .A(\btn_up_debounce.debounce_counter[1] ),
    .B(net713));
 sg13g2_nor2_1 _8083_ (.A(net1807),
    .B(net714),
    .Y(_0282_));
 sg13g2_and3_1 _8084_ (.X(_3543_),
    .A(\btn_up_debounce.debounce_counter[1] ),
    .B(\btn_up_debounce.debounce_counter[0] ),
    .C(net487));
 sg13g2_a21oi_1 _8085_ (.A1(\btn_up_debounce.debounce_counter[1] ),
    .A2(\btn_up_debounce.debounce_counter[0] ),
    .Y(_3544_),
    .B1(net487));
 sg13g2_nor3_1 _8086_ (.A(net1807),
    .B(_3543_),
    .C(net488),
    .Y(_0283_));
 sg13g2_and2_1 _8087_ (.A(net649),
    .B(_3543_),
    .X(_3545_));
 sg13g2_nor2_1 _8088_ (.A(net649),
    .B(_3543_),
    .Y(_3546_));
 sg13g2_nor3_1 _8089_ (.A(net1807),
    .B(_3545_),
    .C(net650),
    .Y(_0284_));
 sg13g2_and2_1 _8090_ (.A(net624),
    .B(_3545_),
    .X(_3547_));
 sg13g2_nor2_1 _8091_ (.A(net624),
    .B(_3545_),
    .Y(_3548_));
 sg13g2_nor3_1 _8092_ (.A(net1807),
    .B(_3547_),
    .C(net625),
    .Y(_0285_));
 sg13g2_and2_1 _8093_ (.A(net619),
    .B(_3547_),
    .X(_3549_));
 sg13g2_nor2_1 _8094_ (.A(net619),
    .B(_3547_),
    .Y(_3550_));
 sg13g2_nor3_1 _8095_ (.A(net1807),
    .B(_3549_),
    .C(net620),
    .Y(_0286_));
 sg13g2_nor2_1 _8096_ (.A(net641),
    .B(_3549_),
    .Y(_3551_));
 sg13g2_and2_1 _8097_ (.A(net641),
    .B(_3549_),
    .X(_3552_));
 sg13g2_nor3_1 _8098_ (.A(net1807),
    .B(_3551_),
    .C(_3552_),
    .Y(_0287_));
 sg13g2_nor2_1 _8099_ (.A(net597),
    .B(_3552_),
    .Y(_3553_));
 sg13g2_and2_1 _8100_ (.A(net597),
    .B(_3552_),
    .X(_3554_));
 sg13g2_nor3_1 _8101_ (.A(_3541_),
    .B(net598),
    .C(_3554_),
    .Y(_0288_));
 sg13g2_nor2_1 _8102_ (.A(net788),
    .B(_3554_),
    .Y(_3555_));
 sg13g2_and2_1 _8103_ (.A(net788),
    .B(_3554_),
    .X(_3556_));
 sg13g2_nor3_1 _8104_ (.A(net1806),
    .B(_3555_),
    .C(_3556_),
    .Y(_0289_));
 sg13g2_xnor2_1 _8105_ (.Y(_3557_),
    .A(net843),
    .B(_3556_));
 sg13g2_nor2_1 _8106_ (.A(net1806),
    .B(_3557_),
    .Y(_0290_));
 sg13g2_a21oi_1 _8107_ (.A1(\btn_up_debounce.debounce_counter[9] ),
    .A2(_3556_),
    .Y(_3558_),
    .B1(net544));
 sg13g2_and3_1 _8108_ (.X(_3559_),
    .A(\btn_up_debounce.debounce_counter[9] ),
    .B(net544),
    .C(_3556_));
 sg13g2_nor3_1 _8109_ (.A(net1806),
    .B(net545),
    .C(_3559_),
    .Y(_0291_));
 sg13g2_xnor2_1 _8110_ (.Y(_3560_),
    .A(net800),
    .B(_3559_));
 sg13g2_nor2_1 _8111_ (.A(_3541_),
    .B(net801),
    .Y(_0292_));
 sg13g2_a21oi_1 _8112_ (.A1(\btn_up_debounce.debounce_counter[11] ),
    .A2(_3559_),
    .Y(_3561_),
    .B1(net562));
 sg13g2_and3_1 _8113_ (.X(_3562_),
    .A(\btn_up_debounce.debounce_counter[11] ),
    .B(net562),
    .C(_3559_));
 sg13g2_nor3_1 _8114_ (.A(_3541_),
    .B(net563),
    .C(_3562_),
    .Y(_0293_));
 sg13g2_nor2_1 _8115_ (.A(net643),
    .B(_3562_),
    .Y(_3563_));
 sg13g2_and2_1 _8116_ (.A(net643),
    .B(_3562_),
    .X(_3564_));
 sg13g2_nor3_1 _8117_ (.A(net1806),
    .B(net644),
    .C(_3564_),
    .Y(_0294_));
 sg13g2_nor2_1 _8118_ (.A(net609),
    .B(_3564_),
    .Y(_3565_));
 sg13g2_and2_1 _8119_ (.A(net609),
    .B(_3564_),
    .X(_3566_));
 sg13g2_nor3_1 _8120_ (.A(net1806),
    .B(net610),
    .C(_3566_),
    .Y(_0295_));
 sg13g2_nor2_1 _8121_ (.A(net618),
    .B(_3566_),
    .Y(_3567_));
 sg13g2_and2_1 _8122_ (.A(net618),
    .B(_3566_),
    .X(_3568_));
 sg13g2_nor3_1 _8123_ (.A(net1806),
    .B(_3567_),
    .C(_3568_),
    .Y(_0296_));
 sg13g2_nor2_1 _8124_ (.A(net623),
    .B(_3568_),
    .Y(_3569_));
 sg13g2_and2_1 _8125_ (.A(net623),
    .B(_3568_),
    .X(_3570_));
 sg13g2_nor3_1 _8126_ (.A(net1806),
    .B(_3569_),
    .C(_3570_),
    .Y(_0297_));
 sg13g2_nor2_1 _8127_ (.A(net552),
    .B(_3570_),
    .Y(_3571_));
 sg13g2_a21oi_1 _8128_ (.A1(net552),
    .A2(_3570_),
    .Y(_3572_),
    .B1(net1806));
 sg13g2_nor2b_1 _8129_ (.A(net553),
    .B_N(_3572_),
    .Y(_0298_));
 sg13g2_and2_1 _8130_ (.A(net2325),
    .B(net977),
    .X(_0299_));
 sg13g2_o21ai_1 _8131_ (.B1(net2331),
    .Y(_3573_),
    .A1(\btn_up_debounce.button_sync_1 ),
    .A2(_3540_));
 sg13g2_a21oi_1 _8132_ (.A1(_4007_),
    .A2(_3540_),
    .Y(_0300_),
    .B1(_3573_));
 sg13g2_and2_1 _8133_ (.A(net2335),
    .B(net2),
    .X(_0301_));
 sg13g2_xor2_1 _8134_ (.B(net459),
    .A(\btn_down_debounce.debounced ),
    .X(_3574_));
 sg13g2_nor2_1 _8135_ (.A(net496),
    .B(\btn_down_debounce.debounce_counter[1] ),
    .Y(_3575_));
 sg13g2_nor3_1 _8136_ (.A(\btn_down_debounce.debounce_counter[3] ),
    .B(\btn_down_debounce.debounce_counter[2] ),
    .C(\btn_down_debounce.debounce_counter[5] ),
    .Y(_3576_));
 sg13g2_nand4_1 _8137_ (.B(\btn_down_debounce.debounce_counter[14] ),
    .C(net484),
    .A(\btn_down_debounce.debounce_counter[15] ),
    .Y(_3577_),
    .D(\btn_down_debounce.debounce_counter[16] ));
 sg13g2_nor3_1 _8138_ (.A(\btn_down_debounce.debounce_counter[11] ),
    .B(\btn_down_debounce.debounce_counter[10] ),
    .C(\btn_down_debounce.debounce_counter[13] ),
    .Y(_3578_));
 sg13g2_nand2_1 _8139_ (.Y(_3579_),
    .A(\btn_down_debounce.debounce_counter[12] ),
    .B(_3578_));
 sg13g2_nor4_1 _8140_ (.A(\btn_down_debounce.debounce_counter[6] ),
    .B(_4038_),
    .C(\btn_down_debounce.debounce_counter[9] ),
    .D(_3577_),
    .Y(_3580_));
 sg13g2_nand4_1 _8141_ (.B(_3575_),
    .C(_3576_),
    .A(\btn_down_debounce.debounce_counter[4] ),
    .Y(_3581_),
    .D(_3580_));
 sg13g2_nor3_1 _8142_ (.A(\btn_down_debounce.debounce_counter[8] ),
    .B(_3579_),
    .C(_3581_),
    .Y(_3582_));
 sg13g2_inv_1 _8143_ (.Y(_3583_),
    .A(_3582_));
 sg13g2_nand3_1 _8144_ (.B(_3574_),
    .C(_3583_),
    .A(net2331),
    .Y(_3584_));
 sg13g2_inv_1 _8145_ (.Y(_3585_),
    .A(net1805));
 sg13g2_and2_1 _8146_ (.A(net440),
    .B(_3585_),
    .X(_0302_));
 sg13g2_and2_1 _8147_ (.A(net496),
    .B(\btn_down_debounce.debounce_counter[1] ),
    .X(_3586_));
 sg13g2_nor3_1 _8148_ (.A(net497),
    .B(net1805),
    .C(_3586_),
    .Y(_0303_));
 sg13g2_and2_1 _8149_ (.A(net667),
    .B(_3586_),
    .X(_3587_));
 sg13g2_nor2_1 _8150_ (.A(net667),
    .B(_3586_),
    .Y(_3588_));
 sg13g2_nor3_1 _8151_ (.A(net1805),
    .B(_3587_),
    .C(net668),
    .Y(_0304_));
 sg13g2_and2_1 _8152_ (.A(net580),
    .B(_3587_),
    .X(_3589_));
 sg13g2_nor2_1 _8153_ (.A(net580),
    .B(_3587_),
    .Y(_3590_));
 sg13g2_nor3_1 _8154_ (.A(net1805),
    .B(_3589_),
    .C(net581),
    .Y(_0305_));
 sg13g2_and2_1 _8155_ (.A(net565),
    .B(_3589_),
    .X(_3591_));
 sg13g2_nor2_1 _8156_ (.A(net565),
    .B(_3589_),
    .Y(_3592_));
 sg13g2_nor3_1 _8157_ (.A(net1805),
    .B(_3591_),
    .C(net566),
    .Y(_0306_));
 sg13g2_and2_1 _8158_ (.A(net604),
    .B(_3591_),
    .X(_3593_));
 sg13g2_nor2_1 _8159_ (.A(net604),
    .B(_3591_),
    .Y(_3594_));
 sg13g2_nor3_1 _8160_ (.A(net1805),
    .B(_3593_),
    .C(_3594_),
    .Y(_0307_));
 sg13g2_nor2_1 _8161_ (.A(net787),
    .B(_3593_),
    .Y(_3595_));
 sg13g2_and2_1 _8162_ (.A(net787),
    .B(_3593_),
    .X(_3596_));
 sg13g2_nor3_1 _8163_ (.A(net1804),
    .B(_3595_),
    .C(_3596_),
    .Y(_0308_));
 sg13g2_nor2_1 _8164_ (.A(net663),
    .B(_3596_),
    .Y(_3597_));
 sg13g2_and2_1 _8165_ (.A(net663),
    .B(_3596_),
    .X(_3598_));
 sg13g2_nor3_1 _8166_ (.A(net1804),
    .B(net664),
    .C(_3598_),
    .Y(_0309_));
 sg13g2_nor2_1 _8167_ (.A(net679),
    .B(_3598_),
    .Y(_3599_));
 sg13g2_and2_1 _8168_ (.A(net679),
    .B(_3598_),
    .X(_3600_));
 sg13g2_nor3_1 _8169_ (.A(net1804),
    .B(_3599_),
    .C(_3600_),
    .Y(_0310_));
 sg13g2_xnor2_1 _8170_ (.Y(_3601_),
    .A(net807),
    .B(_3600_));
 sg13g2_nor2_1 _8171_ (.A(net1804),
    .B(_3601_),
    .Y(_0311_));
 sg13g2_a21oi_1 _8172_ (.A1(\btn_down_debounce.debounce_counter[9] ),
    .A2(_3600_),
    .Y(_3602_),
    .B1(net547));
 sg13g2_and3_1 _8173_ (.X(_3603_),
    .A(net807),
    .B(net547),
    .C(_3600_));
 sg13g2_nor3_1 _8174_ (.A(net1804),
    .B(net548),
    .C(_3603_),
    .Y(_0312_));
 sg13g2_xnor2_1 _8175_ (.Y(_3604_),
    .A(net811),
    .B(_3603_));
 sg13g2_nor2_1 _8176_ (.A(net1804),
    .B(_3604_),
    .Y(_0313_));
 sg13g2_a21oi_1 _8177_ (.A1(\btn_down_debounce.debounce_counter[11] ),
    .A2(_3603_),
    .Y(_3605_),
    .B1(net525));
 sg13g2_and3_1 _8178_ (.X(_3606_),
    .A(net1028),
    .B(net525),
    .C(_3603_));
 sg13g2_nor3_1 _8179_ (.A(net1804),
    .B(net526),
    .C(_3606_),
    .Y(_0314_));
 sg13g2_nor2_1 _8180_ (.A(net665),
    .B(_3606_),
    .Y(_3607_));
 sg13g2_and2_1 _8181_ (.A(net665),
    .B(_3606_),
    .X(_3608_));
 sg13g2_nor3_1 _8182_ (.A(net1804),
    .B(_3607_),
    .C(_3608_),
    .Y(_0315_));
 sg13g2_and2_1 _8183_ (.A(net833),
    .B(_3608_),
    .X(_3609_));
 sg13g2_o21ai_1 _8184_ (.B1(_3585_),
    .Y(_3610_),
    .A1(net833),
    .A2(_3608_));
 sg13g2_nor2_1 _8185_ (.A(_3609_),
    .B(_3610_),
    .Y(_0316_));
 sg13g2_and2_1 _8186_ (.A(net847),
    .B(_3609_),
    .X(_3611_));
 sg13g2_o21ai_1 _8187_ (.B1(_3585_),
    .Y(_3612_),
    .A1(net847),
    .A2(_3609_));
 sg13g2_nor2_1 _8188_ (.A(_3611_),
    .B(_3612_),
    .Y(_0317_));
 sg13g2_o21ai_1 _8189_ (.B1(_3585_),
    .Y(_3613_),
    .A1(net514),
    .A2(_3611_));
 sg13g2_a21oi_1 _8190_ (.A1(net514),
    .A2(_3611_),
    .Y(_0318_),
    .B1(_3613_));
 sg13g2_a21oi_1 _8191_ (.A1(\btn_down_debounce.debounce_counter[16] ),
    .A2(_3611_),
    .Y(_3614_),
    .B1(net484));
 sg13g2_nor2b_1 _8192_ (.A(_3577_),
    .B_N(_3608_),
    .Y(_3615_));
 sg13g2_nor3_1 _8193_ (.A(net1805),
    .B(net485),
    .C(_3615_),
    .Y(_0319_));
 sg13g2_o21ai_1 _8194_ (.B1(net2331),
    .Y(_3616_),
    .A1(net459),
    .A2(_3583_));
 sg13g2_a21oi_1 _8195_ (.A1(_4006_),
    .A2(_3583_),
    .Y(_0320_),
    .B1(net460));
 sg13g2_and2_1 _8196_ (.A(net2335),
    .B(net3),
    .X(_0321_));
 sg13g2_xor2_1 _8197_ (.B(net502),
    .A(\btn_left_debounce.debounced ),
    .X(_3617_));
 sg13g2_nor4_1 _8198_ (.A(\btn_left_debounce.debounce_counter[1] ),
    .B(\btn_left_debounce.debounce_counter[0] ),
    .C(\btn_left_debounce.debounce_counter[3] ),
    .D(\btn_left_debounce.debounce_counter[2] ),
    .Y(_3618_));
 sg13g2_nand2_1 _8199_ (.Y(_3619_),
    .A(\btn_left_debounce.debounce_counter[12] ),
    .B(\btn_left_debounce.debounce_counter[17] ));
 sg13g2_or4_1 _8200_ (.A(\btn_left_debounce.debounce_counter[9] ),
    .B(\btn_left_debounce.debounce_counter[8] ),
    .C(\btn_left_debounce.debounce_counter[11] ),
    .D(\btn_left_debounce.debounce_counter[10] ),
    .X(_3620_));
 sg13g2_nand2_1 _8201_ (.Y(_3621_),
    .A(\btn_left_debounce.debounce_counter[4] ),
    .B(\btn_left_debounce.debounce_counter[7] ));
 sg13g2_nor4_1 _8202_ (.A(\btn_left_debounce.debounce_counter[13] ),
    .B(_4037_),
    .C(_3619_),
    .D(_3621_),
    .Y(_3622_));
 sg13g2_nand4_1 _8203_ (.B(\btn_left_debounce.debounce_counter[16] ),
    .C(_3618_),
    .A(\btn_left_debounce.debounce_counter[15] ),
    .Y(_3623_),
    .D(_3622_));
 sg13g2_nor4_1 _8204_ (.A(\btn_left_debounce.debounce_counter[5] ),
    .B(\btn_left_debounce.debounce_counter[6] ),
    .C(_3620_),
    .D(_3623_),
    .Y(_3624_));
 sg13g2_inv_1 _8205_ (.Y(_3625_),
    .A(_3624_));
 sg13g2_nand3_1 _8206_ (.B(_3617_),
    .C(_3625_),
    .A(net2331),
    .Y(_3626_));
 sg13g2_nor2_1 _8207_ (.A(_4076_),
    .B(net1802),
    .Y(_0322_));
 sg13g2_xnor2_1 _8208_ (.Y(_3627_),
    .A(net828),
    .B(\btn_left_debounce.debounce_counter[0] ));
 sg13g2_nor2_1 _8209_ (.A(net1802),
    .B(net829),
    .Y(_0323_));
 sg13g2_and3_1 _8210_ (.X(_3628_),
    .A(\btn_left_debounce.debounce_counter[1] ),
    .B(\btn_left_debounce.debounce_counter[0] ),
    .C(net531));
 sg13g2_a21oi_1 _8211_ (.A1(\btn_left_debounce.debounce_counter[1] ),
    .A2(\btn_left_debounce.debounce_counter[0] ),
    .Y(_3629_),
    .B1(net531));
 sg13g2_nor3_1 _8212_ (.A(net1802),
    .B(_3628_),
    .C(net532),
    .Y(_0324_));
 sg13g2_and2_1 _8213_ (.A(net639),
    .B(_3628_),
    .X(_3630_));
 sg13g2_nor2_1 _8214_ (.A(net639),
    .B(_3628_),
    .Y(_3631_));
 sg13g2_nor3_1 _8215_ (.A(net1802),
    .B(_3630_),
    .C(net640),
    .Y(_0325_));
 sg13g2_and2_1 _8216_ (.A(net572),
    .B(_3630_),
    .X(_3632_));
 sg13g2_nor2_1 _8217_ (.A(net572),
    .B(_3630_),
    .Y(_3633_));
 sg13g2_nor3_1 _8218_ (.A(net1802),
    .B(_3632_),
    .C(net573),
    .Y(_0326_));
 sg13g2_and2_1 _8219_ (.A(net626),
    .B(_3632_),
    .X(_3634_));
 sg13g2_nor2_1 _8220_ (.A(net626),
    .B(_3632_),
    .Y(_3635_));
 sg13g2_nor3_1 _8221_ (.A(net1803),
    .B(_3634_),
    .C(_3635_),
    .Y(_0327_));
 sg13g2_nor2_1 _8222_ (.A(net635),
    .B(_3634_),
    .Y(_3636_));
 sg13g2_and2_1 _8223_ (.A(net635),
    .B(_3634_),
    .X(_3637_));
 sg13g2_nor3_1 _8224_ (.A(net1803),
    .B(_3636_),
    .C(_3637_),
    .Y(_0328_));
 sg13g2_nor2_1 _8225_ (.A(net658),
    .B(_3637_),
    .Y(_3638_));
 sg13g2_and2_1 _8226_ (.A(net658),
    .B(_3637_),
    .X(_3639_));
 sg13g2_nor3_1 _8227_ (.A(net1802),
    .B(_3638_),
    .C(_3639_),
    .Y(_0329_));
 sg13g2_nor2_1 _8228_ (.A(net687),
    .B(_3639_),
    .Y(_3640_));
 sg13g2_and2_1 _8229_ (.A(net687),
    .B(_3639_),
    .X(_3641_));
 sg13g2_nor3_1 _8230_ (.A(net1802),
    .B(_3640_),
    .C(_3641_),
    .Y(_0330_));
 sg13g2_xnor2_1 _8231_ (.Y(_3642_),
    .A(net803),
    .B(_3641_));
 sg13g2_nor2_1 _8232_ (.A(net1802),
    .B(_3642_),
    .Y(_0331_));
 sg13g2_a21oi_1 _8233_ (.A1(\btn_left_debounce.debounce_counter[9] ),
    .A2(_3641_),
    .Y(_3643_),
    .B1(net520));
 sg13g2_and3_1 _8234_ (.X(_3644_),
    .A(\btn_left_debounce.debounce_counter[9] ),
    .B(net520),
    .C(_3641_));
 sg13g2_nor3_1 _8235_ (.A(_3626_),
    .B(net521),
    .C(_3644_),
    .Y(_0332_));
 sg13g2_xnor2_1 _8236_ (.Y(_3645_),
    .A(net767),
    .B(_3644_));
 sg13g2_nor2_1 _8237_ (.A(_3626_),
    .B(_3645_),
    .Y(_0333_));
 sg13g2_a21oi_1 _8238_ (.A1(\btn_left_debounce.debounce_counter[11] ),
    .A2(_3644_),
    .Y(_3646_),
    .B1(net536));
 sg13g2_and3_1 _8239_ (.X(_3647_),
    .A(\btn_left_debounce.debounce_counter[11] ),
    .B(net536),
    .C(_3644_));
 sg13g2_nor3_1 _8240_ (.A(net1803),
    .B(net537),
    .C(_3647_),
    .Y(_0334_));
 sg13g2_nor2_1 _8241_ (.A(net659),
    .B(_3647_),
    .Y(_3648_));
 sg13g2_and2_1 _8242_ (.A(net659),
    .B(_3647_),
    .X(_3649_));
 sg13g2_nor3_1 _8243_ (.A(net1803),
    .B(net660),
    .C(_3649_),
    .Y(_0335_));
 sg13g2_nor2_1 _8244_ (.A(net671),
    .B(_3649_),
    .Y(_3650_));
 sg13g2_and2_1 _8245_ (.A(net671),
    .B(_3649_),
    .X(_3651_));
 sg13g2_nor3_1 _8246_ (.A(_3626_),
    .B(_3650_),
    .C(_3651_),
    .Y(_0336_));
 sg13g2_nor2_1 _8247_ (.A(net630),
    .B(_3651_),
    .Y(_3652_));
 sg13g2_and2_1 _8248_ (.A(net630),
    .B(_3651_),
    .X(_3653_));
 sg13g2_nor3_1 _8249_ (.A(net1803),
    .B(net631),
    .C(_3653_),
    .Y(_0337_));
 sg13g2_nor2_1 _8250_ (.A(net698),
    .B(_3653_),
    .Y(_3654_));
 sg13g2_and2_1 _8251_ (.A(net698),
    .B(_3653_),
    .X(_3655_));
 sg13g2_nor3_1 _8252_ (.A(net1803),
    .B(_3654_),
    .C(_3655_),
    .Y(_0338_));
 sg13g2_nor2_1 _8253_ (.A(net588),
    .B(_3655_),
    .Y(_3656_));
 sg13g2_a21oi_1 _8254_ (.A1(net588),
    .A2(_3655_),
    .Y(_3657_),
    .B1(net1803));
 sg13g2_nor2b_1 _8255_ (.A(net589),
    .B_N(_3657_),
    .Y(_0339_));
 sg13g2_and2_1 _8256_ (.A(net2331),
    .B(net943),
    .X(_0340_));
 sg13g2_o21ai_1 _8257_ (.B1(net2331),
    .Y(_3658_),
    .A1(net502),
    .A2(_3625_));
 sg13g2_a21oi_1 _8258_ (.A1(_4005_),
    .A2(_3625_),
    .Y(_0341_),
    .B1(net503));
 sg13g2_and2_1 _8259_ (.A(net2323),
    .B(net4),
    .X(_0342_));
 sg13g2_xor2_1 _8260_ (.B(\btn_right_debounce.button_sync_1 ),
    .A(\btn_right_debounce.debounced ),
    .X(_3659_));
 sg13g2_nor4_1 _8261_ (.A(\btn_right_debounce.debounce_counter[1] ),
    .B(\btn_right_debounce.debounce_counter[0] ),
    .C(\btn_right_debounce.debounce_counter[3] ),
    .D(\btn_right_debounce.debounce_counter[2] ),
    .Y(_3660_));
 sg13g2_nand3_1 _8262_ (.B(\btn_right_debounce.debounce_counter[16] ),
    .C(_3660_),
    .A(\btn_right_debounce.debounce_counter[15] ),
    .Y(_3661_));
 sg13g2_nand4_1 _8263_ (.B(\btn_right_debounce.debounce_counter[12] ),
    .C(\btn_right_debounce.debounce_counter[14] ),
    .A(_4036_),
    .Y(_3662_),
    .D(\btn_right_debounce.debounce_counter[17] ));
 sg13g2_nor4_1 _8264_ (.A(\btn_right_debounce.debounce_counter[9] ),
    .B(\btn_right_debounce.debounce_counter[8] ),
    .C(\btn_right_debounce.debounce_counter[11] ),
    .D(net522),
    .Y(_3663_));
 sg13g2_nor4_1 _8265_ (.A(\btn_right_debounce.debounce_counter[5] ),
    .B(\btn_right_debounce.debounce_counter[6] ),
    .C(_3661_),
    .D(_3662_),
    .Y(_3664_));
 sg13g2_and4_1 _8266_ (.A(net570),
    .B(net611),
    .C(_3663_),
    .D(_3664_),
    .X(_3665_));
 sg13g2_inv_1 _8267_ (.Y(_3666_),
    .A(_3665_));
 sg13g2_nand3_1 _8268_ (.B(_3659_),
    .C(_3666_),
    .A(net2326),
    .Y(_3667_));
 sg13g2_inv_1 _8269_ (.Y(_3668_),
    .A(net1800));
 sg13g2_and2_1 _8270_ (.A(net442),
    .B(_3668_),
    .X(_0343_));
 sg13g2_xnor2_1 _8271_ (.Y(_3669_),
    .A(net839),
    .B(\btn_right_debounce.debounce_counter[0] ));
 sg13g2_nor2_1 _8272_ (.A(net1800),
    .B(net840),
    .Y(_0344_));
 sg13g2_and3_1 _8273_ (.X(_3670_),
    .A(\btn_right_debounce.debounce_counter[1] ),
    .B(\btn_right_debounce.debounce_counter[0] ),
    .C(net492));
 sg13g2_a21oi_1 _8274_ (.A1(\btn_right_debounce.debounce_counter[1] ),
    .A2(\btn_right_debounce.debounce_counter[0] ),
    .Y(_3671_),
    .B1(net492));
 sg13g2_nor3_1 _8275_ (.A(net1801),
    .B(_3670_),
    .C(net493),
    .Y(_0345_));
 sg13g2_and2_1 _8276_ (.A(net672),
    .B(_3670_),
    .X(_3672_));
 sg13g2_nor2_1 _8277_ (.A(net672),
    .B(_3670_),
    .Y(_3673_));
 sg13g2_nor3_1 _8278_ (.A(net1801),
    .B(_3672_),
    .C(net673),
    .Y(_0346_));
 sg13g2_and2_1 _8279_ (.A(net570),
    .B(_3672_),
    .X(_3674_));
 sg13g2_nor2_1 _8280_ (.A(net570),
    .B(_3672_),
    .Y(_3675_));
 sg13g2_nor3_1 _8281_ (.A(net1800),
    .B(_3674_),
    .C(net571),
    .Y(_0347_));
 sg13g2_and2_1 _8282_ (.A(net629),
    .B(_3674_),
    .X(_3676_));
 sg13g2_nor2_1 _8283_ (.A(net629),
    .B(_3674_),
    .Y(_3677_));
 sg13g2_nor3_1 _8284_ (.A(net1800),
    .B(_3676_),
    .C(_3677_),
    .Y(_0348_));
 sg13g2_nor2_1 _8285_ (.A(net666),
    .B(_3676_),
    .Y(_3678_));
 sg13g2_and2_1 _8286_ (.A(net666),
    .B(_3676_),
    .X(_3679_));
 sg13g2_nor3_1 _8287_ (.A(net1800),
    .B(_3678_),
    .C(_3679_),
    .Y(_0349_));
 sg13g2_nor2_1 _8288_ (.A(net611),
    .B(_3679_),
    .Y(_3680_));
 sg13g2_and2_1 _8289_ (.A(net611),
    .B(_3679_),
    .X(_3681_));
 sg13g2_nor3_1 _8290_ (.A(net1801),
    .B(net612),
    .C(_3681_),
    .Y(_0350_));
 sg13g2_nor2_1 _8291_ (.A(net600),
    .B(_3681_),
    .Y(_3682_));
 sg13g2_and2_1 _8292_ (.A(net600),
    .B(_3681_),
    .X(_3683_));
 sg13g2_nor3_1 _8293_ (.A(net1801),
    .B(net601),
    .C(_3683_),
    .Y(_0351_));
 sg13g2_xnor2_1 _8294_ (.Y(_3684_),
    .A(net820),
    .B(_3683_));
 sg13g2_nor2_1 _8295_ (.A(net1801),
    .B(_3684_),
    .Y(_0352_));
 sg13g2_a21oi_1 _8296_ (.A1(\btn_right_debounce.debounce_counter[9] ),
    .A2(_3683_),
    .Y(_3685_),
    .B1(net522));
 sg13g2_and3_1 _8297_ (.X(_3686_),
    .A(net820),
    .B(net522),
    .C(_3683_));
 sg13g2_nor3_1 _8298_ (.A(net1801),
    .B(net523),
    .C(_3686_),
    .Y(_0353_));
 sg13g2_xnor2_1 _8299_ (.Y(_3687_),
    .A(net841),
    .B(_3686_));
 sg13g2_nor2_1 _8300_ (.A(net1801),
    .B(_3687_),
    .Y(_0354_));
 sg13g2_a21oi_1 _8301_ (.A1(\btn_right_debounce.debounce_counter[11] ),
    .A2(_3686_),
    .Y(_3688_),
    .B1(net574));
 sg13g2_and3_1 _8302_ (.X(_3689_),
    .A(\btn_right_debounce.debounce_counter[11] ),
    .B(net574),
    .C(_3686_));
 sg13g2_nor3_1 _8303_ (.A(net1800),
    .B(net575),
    .C(_3689_),
    .Y(_0355_));
 sg13g2_nor2_1 _8304_ (.A(net632),
    .B(_3689_),
    .Y(_3690_));
 sg13g2_and2_1 _8305_ (.A(net632),
    .B(_3689_),
    .X(_3691_));
 sg13g2_nor3_1 _8306_ (.A(net1800),
    .B(net633),
    .C(_3691_),
    .Y(_0356_));
 sg13g2_and2_1 _8307_ (.A(net836),
    .B(_3691_),
    .X(_3692_));
 sg13g2_o21ai_1 _8308_ (.B1(_3668_),
    .Y(_3693_),
    .A1(net836),
    .A2(_3691_));
 sg13g2_nor2_1 _8309_ (.A(_3692_),
    .B(_3693_),
    .Y(_0357_));
 sg13g2_o21ai_1 _8310_ (.B1(_3668_),
    .Y(_3694_),
    .A1(net584),
    .A2(_3692_));
 sg13g2_a21oi_1 _8311_ (.A1(net584),
    .A2(_3692_),
    .Y(_0358_),
    .B1(_3694_));
 sg13g2_a21oi_1 _8312_ (.A1(\btn_right_debounce.debounce_counter[15] ),
    .A2(_3692_),
    .Y(_3695_),
    .B1(net528));
 sg13g2_and3_1 _8313_ (.X(_3696_),
    .A(\btn_right_debounce.debounce_counter[15] ),
    .B(net528),
    .C(_3692_));
 sg13g2_nor3_1 _8314_ (.A(net1800),
    .B(net529),
    .C(_3696_),
    .Y(_0359_));
 sg13g2_o21ai_1 _8315_ (.B1(_3668_),
    .Y(_3697_),
    .A1(net500),
    .A2(_3696_));
 sg13g2_a21oi_1 _8316_ (.A1(net500),
    .A2(_3696_),
    .Y(_0360_),
    .B1(_3697_));
 sg13g2_and2_1 _8317_ (.A(net2332),
    .B(net944),
    .X(_0361_));
 sg13g2_o21ai_1 _8318_ (.B1(net2326),
    .Y(_3698_),
    .A1(\btn_right_debounce.button_sync_1 ),
    .A2(_3666_));
 sg13g2_a21oi_1 _8319_ (.A1(_4004_),
    .A2(_3666_),
    .Y(_0362_),
    .B1(_3698_));
 sg13g2_and2_1 _8320_ (.A(net2314),
    .B(_0506_),
    .X(_0363_));
 sg13g2_nor2b_1 _8321_ (.A(net634),
    .B_N(net417),
    .Y(_3699_));
 sg13g2_nor2_1 _8322_ (.A(net2304),
    .B(net1960),
    .Y(_3700_));
 sg13g2_a22oi_1 _8323_ (.Y(_0364_),
    .B1(net1847),
    .B2(_4002_),
    .A2(net1960),
    .A1(_4003_));
 sg13g2_a22oi_1 _8324_ (.Y(_0365_),
    .B1(net1847),
    .B2(_4001_),
    .A2(net1959),
    .A1(_4002_));
 sg13g2_a22oi_1 _8325_ (.Y(_0366_),
    .B1(net1846),
    .B2(_4000_),
    .A2(net1959),
    .A1(_4001_));
 sg13g2_a22oi_1 _8326_ (.Y(_0367_),
    .B1(net1846),
    .B2(_3999_),
    .A2(net1959),
    .A1(_4000_));
 sg13g2_a22oi_1 _8327_ (.Y(_0368_),
    .B1(net1846),
    .B2(_3998_),
    .A2(net1959),
    .A1(_3999_));
 sg13g2_a22oi_1 _8328_ (.Y(_0369_),
    .B1(net1846),
    .B2(_3997_),
    .A2(net1959),
    .A1(_3998_));
 sg13g2_a22oi_1 _8329_ (.Y(_0370_),
    .B1(net1846),
    .B2(_3996_),
    .A2(net1959),
    .A1(_3997_));
 sg13g2_a22oi_1 _8330_ (.Y(_0371_),
    .B1(net1846),
    .B2(_3995_),
    .A2(net1959),
    .A1(_3996_));
 sg13g2_a22oi_1 _8331_ (.Y(_0372_),
    .B1(net1847),
    .B2(_3994_),
    .A2(net1960),
    .A1(_3995_));
 sg13g2_a22oi_1 _8332_ (.Y(_0373_),
    .B1(net1847),
    .B2(_3993_),
    .A2(net1960),
    .A1(_3994_));
 sg13g2_a22oi_1 _8333_ (.Y(_0374_),
    .B1(net1846),
    .B2(_3992_),
    .A2(net1959),
    .A1(_3993_));
 sg13g2_a22oi_1 _8334_ (.Y(_0375_),
    .B1(net1846),
    .B2(_3991_),
    .A2(net1960),
    .A1(_3992_));
 sg13g2_and2_1 _8335_ (.A(net2323),
    .B(net7),
    .X(_0376_));
 sg13g2_and2_2 _8336_ (.A(net2335),
    .B(net804),
    .X(_0377_));
 sg13g2_and2_1 _8337_ (.A(net2335),
    .B(net6),
    .X(_0378_));
 sg13g2_and2_1 _8338_ (.A(net2329),
    .B(net797),
    .X(_0379_));
 sg13g2_xor2_1 _8339_ (.B(net473),
    .A(net517),
    .X(_3701_));
 sg13g2_xor2_1 _8340_ (.B(net790),
    .A(net882),
    .X(_3702_));
 sg13g2_o21ai_1 _8341_ (.B1(net2313),
    .Y(_3703_),
    .A1(_3701_),
    .A2(_3702_));
 sg13g2_a21oi_1 _8342_ (.A1(_3701_),
    .A2(_3702_),
    .Y(_0380_),
    .B1(_3703_));
 sg13g2_nand2b_1 _8343_ (.Y(_0381_),
    .B(net2312),
    .A_N(net790));
 sg13g2_and2_1 _8344_ (.A(net2308),
    .B(net517),
    .X(_0382_));
 sg13g2_nand2b_1 _8345_ (.Y(_0383_),
    .B(net2309),
    .A_N(net539));
 sg13g2_nand2b_1 _8346_ (.Y(_0384_),
    .B(net2308),
    .A_N(net462));
 sg13g2_nand2b_1 _8347_ (.Y(_0385_),
    .B(net2308),
    .A_N(net505));
 sg13g2_nand2b_1 _8348_ (.Y(_0386_),
    .B(net2308),
    .A_N(net483));
 sg13g2_nand2b_1 _8349_ (.Y(_0387_),
    .B(net2308),
    .A_N(net495));
 sg13g2_and2_1 _8350_ (.A(net2308),
    .B(net516),
    .X(_0388_));
 sg13g2_nand2b_1 _8351_ (.Y(_0389_),
    .B(net2308),
    .A_N(net478));
 sg13g2_and2_1 _8352_ (.A(net2309),
    .B(net464),
    .X(_0390_));
 sg13g2_nand2b_1 _8353_ (.Y(_0391_),
    .B(net2311),
    .A_N(net542));
 sg13g2_nand2b_1 _8354_ (.Y(_0392_),
    .B(net2310),
    .A_N(net482));
 sg13g2_nand2b_1 _8355_ (.Y(_0393_),
    .B(net2310),
    .A_N(net499));
 sg13g2_nand2b_1 _8356_ (.Y(_0394_),
    .B(net2310),
    .A_N(net476));
 sg13g2_nand2b_1 _8357_ (.Y(_0395_),
    .B(net2310),
    .A_N(net577));
 sg13g2_and2_1 _8358_ (.A(net2310),
    .B(net477),
    .X(_0396_));
 sg13g2_and2_1 _8359_ (.A(net2310),
    .B(net447),
    .X(_0397_));
 sg13g2_and2_1 _8360_ (.A(net2312),
    .B(net454),
    .X(_0398_));
 sg13g2_nand2b_1 _8361_ (.Y(_0399_),
    .B(net2312),
    .A_N(net457));
 sg13g2_and2_1 _8362_ (.A(net2312),
    .B(net449),
    .X(_0400_));
 sg13g2_and2_1 _8363_ (.A(net2312),
    .B(net472),
    .X(_0401_));
 sg13g2_nand2b_1 _8364_ (.Y(_0402_),
    .B(net2312),
    .A_N(net473));
 sg13g2_and2_1 _8365_ (.A(net2314),
    .B(net471),
    .X(_0403_));
 sg13g2_and2_1 _8366_ (.A(net2314),
    .B(net455),
    .X(_0404_));
 sg13g2_and2_1 _8367_ (.A(net2314),
    .B(net453),
    .X(_0405_));
 sg13g2_and2_1 _8368_ (.A(net2314),
    .B(net448),
    .X(_0406_));
 sg13g2_and2_1 _8369_ (.A(net2325),
    .B(net446),
    .X(_0407_));
 sg13g2_and2_1 _8370_ (.A(net2325),
    .B(net450),
    .X(_0408_));
 sg13g2_nand2b_1 _8371_ (.Y(_0409_),
    .B(net2326),
    .A_N(net2272));
 sg13g2_and2_1 _8372_ (.A(net2325),
    .B(net2270),
    .X(_0410_));
 sg13g2_nor2_1 _8373_ (.A(net2305),
    .B(_4025_),
    .Y(_0411_));
 sg13g2_nand2_1 _8374_ (.Y(_3704_),
    .A(\draw_game_inst.y[9] ),
    .B(net1883));
 sg13g2_nor4_1 _8375_ (.A(\draw_game_inst.y[8] ),
    .B(\draw_game_inst.y[7] ),
    .C(\draw_game_inst.board_y[6] ),
    .D(_3704_),
    .Y(_3705_));
 sg13g2_a21oi_2 _8376_ (.B1(net2306),
    .Y(_3706_),
    .A2(_3705_),
    .A1(_1478_));
 sg13g2_nand2_2 _8377_ (.Y(_3707_),
    .A(_1446_),
    .B(_3706_));
 sg13g2_inv_1 _8378_ (.Y(_3708_),
    .A(_3707_));
 sg13g2_a22oi_1 _8379_ (.Y(_3709_),
    .B1(_3708_),
    .B2(net2251),
    .A2(net1815),
    .A1(net2256));
 sg13g2_inv_1 _8380_ (.Y(_0412_),
    .A(_3709_));
 sg13g2_o21ai_1 _8381_ (.B1(_3708_),
    .Y(_3710_),
    .A1(net1857),
    .A2(net1848));
 sg13g2_o21ai_1 _8382_ (.B1(_3710_),
    .Y(_0413_),
    .A1(net2069),
    .A2(_1448_));
 sg13g2_nand2_1 _8383_ (.Y(_3711_),
    .A(net2209),
    .B(net1815));
 sg13g2_o21ai_1 _8384_ (.B1(_3711_),
    .Y(_0414_),
    .A1(_3243_),
    .A2(_3707_));
 sg13g2_or3_1 _8385_ (.A(net2203),
    .B(net1991),
    .C(_3707_),
    .X(_3712_));
 sg13g2_nor2_1 _8386_ (.A(net1815),
    .B(_3706_),
    .Y(_3713_));
 sg13g2_nor3_1 _8387_ (.A(net2087),
    .B(net2203),
    .C(net1991),
    .Y(_3714_));
 sg13g2_a221oi_1 _8388_ (.B2(_1448_),
    .C1(_3713_),
    .B1(_3714_),
    .A1(net2087),
    .Y(_0415_),
    .A2(_3712_));
 sg13g2_nand3_1 _8389_ (.B(net1890),
    .C(net1883),
    .A(_1448_),
    .Y(_3715_));
 sg13g2_xor2_1 _8390_ (.B(_3715_),
    .A(net2184),
    .X(_3716_));
 sg13g2_nor2_1 _8391_ (.A(_3713_),
    .B(_3716_),
    .Y(_0416_));
 sg13g2_nand2_1 _8392_ (.Y(_3717_),
    .A(net2181),
    .B(_1447_));
 sg13g2_nor3_1 _8393_ (.A(net2183),
    .B(net1991),
    .C(net1986),
    .Y(_3718_));
 sg13g2_xnor2_1 _8394_ (.Y(_3719_),
    .A(net2181),
    .B(_3718_));
 sg13g2_o21ai_1 _8395_ (.B1(_3717_),
    .Y(_0417_),
    .A1(_3707_),
    .A2(_3719_));
 sg13g2_nor2_1 _8396_ (.A(net1815),
    .B(_3321_),
    .Y(_3720_));
 sg13g2_xnor2_1 _8397_ (.Y(_3721_),
    .A(net910),
    .B(_3720_));
 sg13g2_nor2_1 _8398_ (.A(_3713_),
    .B(_3721_),
    .Y(_0418_));
 sg13g2_nand2_1 _8399_ (.Y(_3722_),
    .A(\draw_game_inst.y[7] ),
    .B(net1815));
 sg13g2_nor2_1 _8400_ (.A(net770),
    .B(_3321_),
    .Y(_3723_));
 sg13g2_xnor2_1 _8401_ (.Y(_3724_),
    .A(\draw_game_inst.y[7] ),
    .B(_3723_));
 sg13g2_o21ai_1 _8402_ (.B1(_3722_),
    .Y(_0419_),
    .A1(_3707_),
    .A2(net771));
 sg13g2_a21oi_1 _8403_ (.A1(net2031),
    .A2(_3720_),
    .Y(_3725_),
    .B1(net858));
 sg13g2_or2_1 _8404_ (.X(_3726_),
    .B(_3321_),
    .A(_1426_));
 sg13g2_a21oi_1 _8405_ (.A1(_3706_),
    .A2(_3726_),
    .Y(_3727_),
    .B1(net1815));
 sg13g2_nor2_1 _8406_ (.A(_3725_),
    .B(_3727_),
    .Y(_0420_));
 sg13g2_nand4_1 _8407_ (.B(net2031),
    .C(_1472_),
    .A(net858),
    .Y(_3728_),
    .D(_3720_));
 sg13g2_o21ai_1 _8408_ (.B1(net859),
    .Y(_0421_),
    .A1(_4040_),
    .A2(_3727_));
 sg13g2_and2_1 _8409_ (.A(net2335),
    .B(net5),
    .X(_0422_));
 sg13g2_and2_1 _8410_ (.A(net2329),
    .B(net848),
    .X(_0423_));
 sg13g2_nor2b_1 _8411_ (.A(\gamepad_pmod.driver.pmod_latch_prev ),
    .B_N(net416),
    .Y(_3729_));
 sg13g2_nor2_1 _8412_ (.A(net2304),
    .B(net1957),
    .Y(_3730_));
 sg13g2_a22oi_1 _8413_ (.Y(_0424_),
    .B1(net1845),
    .B2(_4011_),
    .A2(net1958),
    .A1(_4002_));
 sg13g2_a22oi_1 _8414_ (.Y(_0425_),
    .B1(net1845),
    .B2(_4010_),
    .A2(net1958),
    .A1(_4001_));
 sg13g2_a22oi_1 _8415_ (.Y(_0426_),
    .B1(net1845),
    .B2(_4013_),
    .A2(net1958),
    .A1(_4000_));
 sg13g2_a22oi_1 _8416_ (.Y(_0427_),
    .B1(net1845),
    .B2(_4012_),
    .A2(net1958),
    .A1(_3999_));
 sg13g2_a22oi_1 _8417_ (.Y(_0428_),
    .B1(net1844),
    .B2(_4015_),
    .A2(net1957),
    .A1(_3998_));
 sg13g2_a22oi_1 _8418_ (.Y(_0429_),
    .B1(net1844),
    .B2(_4014_),
    .A2(net1957),
    .A1(_3997_));
 sg13g2_a22oi_1 _8419_ (.Y(_0430_),
    .B1(net1844),
    .B2(_4017_),
    .A2(net1957),
    .A1(_3996_));
 sg13g2_a22oi_1 _8420_ (.Y(_0431_),
    .B1(net1844),
    .B2(_4016_),
    .A2(net1957),
    .A1(_3995_));
 sg13g2_a22oi_1 _8421_ (.Y(_0432_),
    .B1(net1844),
    .B2(_4019_),
    .A2(net1957),
    .A1(_3994_));
 sg13g2_a22oi_1 _8422_ (.Y(_0433_),
    .B1(net1844),
    .B2(_4018_),
    .A2(net1957),
    .A1(_3993_));
 sg13g2_a22oi_1 _8423_ (.Y(_0434_),
    .B1(net1844),
    .B2(_4021_),
    .A2(net1958),
    .A1(_3992_));
 sg13g2_a22oi_1 _8424_ (.Y(_0435_),
    .B1(net1844),
    .B2(_4020_),
    .A2(net1957),
    .A1(_3991_));
 sg13g2_nor2b_2 _8425_ (.A(\lfsr_inst.lfsr[29] ),
    .B_N(net2271),
    .Y(_3731_));
 sg13g2_nand2b_1 _8426_ (.Y(_3732_),
    .B(net2272),
    .A_N(net2270));
 sg13g2_and2_1 _8427_ (.A(net2271),
    .B(net2270),
    .X(_3733_));
 sg13g2_nand2_1 _8428_ (.Y(_3734_),
    .A(net2271),
    .B(\lfsr_inst.lfsr[29] ));
 sg13g2_nor2_2 _8429_ (.A(net2271),
    .B(net2270),
    .Y(_3735_));
 sg13g2_nor2b_2 _8430_ (.A(net2271),
    .B_N(net2270),
    .Y(_3736_));
 sg13g2_nand2b_1 _8431_ (.Y(_3737_),
    .B(net2270),
    .A_N(net2272));
 sg13g2_a22oi_1 _8432_ (.Y(_3738_),
    .B1(_3733_),
    .B2(\welcome_screen_grid[60] ),
    .A2(_3731_),
    .A1(\welcome_screen_grid[52] ));
 sg13g2_a221oi_1 _8433_ (.B2(\welcome_screen_grid[56] ),
    .C1(_4025_),
    .B1(_3736_),
    .A1(\welcome_screen_grid[48] ),
    .Y(_3739_),
    .A2(_3735_));
 sg13g2_nand2_1 _8434_ (.Y(_3740_),
    .A(_3738_),
    .B(_3739_));
 sg13g2_a21oi_1 _8435_ (.A1(\welcome_screen_grid[40] ),
    .A2(_3736_),
    .Y(_3741_),
    .B1(\lfsr_inst.lfsr[30] ));
 sg13g2_nand2_1 _8436_ (.Y(_3742_),
    .A(\welcome_screen_grid[32] ),
    .B(_3735_));
 sg13g2_a22oi_1 _8437_ (.Y(_3743_),
    .B1(_3733_),
    .B2(\welcome_screen_grid[44] ),
    .A2(_3731_),
    .A1(\welcome_screen_grid[36] ));
 sg13g2_nand3_1 _8438_ (.B(_3742_),
    .C(_3743_),
    .A(_3741_),
    .Y(_3744_));
 sg13g2_nand3_1 _8439_ (.B(_3740_),
    .C(_3744_),
    .A(\lfsr_inst.lfsr[31] ),
    .Y(_3745_));
 sg13g2_nand4_1 _8440_ (.B(\welcome_screen_inst.welcome_counter[3] ),
    .C(net676),
    .A(net736),
    .Y(_3746_),
    .D(\welcome_screen_inst.welcome_counter[1] ));
 sg13g2_nor2_2 _8441_ (.A(\welcome_screen_inst.welcome_counter[0] ),
    .B(_3746_),
    .Y(_3747_));
 sg13g2_and2_1 _8442_ (.A(\welcome_screen_grid[0] ),
    .B(_3735_),
    .X(_3748_));
 sg13g2_a21oi_1 _8443_ (.A1(\welcome_screen_grid[11] ),
    .A2(_3736_),
    .Y(_3749_),
    .B1(\lfsr_inst.lfsr[30] ));
 sg13g2_a221oi_1 _8444_ (.B2(\welcome_screen_grid[12] ),
    .C1(_3748_),
    .B1(_3733_),
    .A1(\welcome_screen_grid[4] ),
    .Y(_3750_),
    .A2(_3731_));
 sg13g2_a22oi_1 _8445_ (.Y(_3751_),
    .B1(_3736_),
    .B2(\welcome_screen_grid[24] ),
    .A2(_3733_),
    .A1(\welcome_screen_grid[28] ));
 sg13g2_a221oi_1 _8446_ (.B2(\welcome_screen_grid[16] ),
    .C1(_4025_),
    .B1(_3735_),
    .A1(\welcome_screen_grid[20] ),
    .Y(_3752_),
    .A2(_3731_));
 sg13g2_a221oi_1 _8447_ (.B2(_3752_),
    .C1(\lfsr_inst.lfsr[31] ),
    .B1(_3751_),
    .A1(_3749_),
    .Y(_3753_),
    .A2(_3750_));
 sg13g2_nand2b_1 _8448_ (.Y(_3754_),
    .B(_3747_),
    .A_N(_3753_));
 sg13g2_nand2b_1 _8449_ (.Y(_3755_),
    .B(_3745_),
    .A_N(_3754_));
 sg13g2_nor4_1 _8450_ (.A(net2271),
    .B(net2270),
    .C(\lfsr_inst.lfsr[30] ),
    .D(\lfsr_inst.lfsr[31] ),
    .Y(_3756_));
 sg13g2_o21ai_1 _8451_ (.B1(net2325),
    .Y(_3757_),
    .A1(net1797),
    .A2(_3756_));
 sg13g2_a21oi_1 _8452_ (.A1(_3990_),
    .A2(net1797),
    .Y(_0436_),
    .B1(_3757_));
 sg13g2_nand2b_1 _8453_ (.Y(_3758_),
    .B(_4025_),
    .A_N(_3754_));
 sg13g2_nor2_1 _8454_ (.A(_3732_),
    .B(_3758_),
    .Y(_3759_));
 sg13g2_a22oi_1 _8455_ (.Y(_3760_),
    .B1(_3759_),
    .B2(net2094),
    .A2(net1797),
    .A1(net642));
 sg13g2_nor2_1 _8456_ (.A(net2305),
    .B(_3760_),
    .Y(_0437_));
 sg13g2_nor2_1 _8457_ (.A(_3737_),
    .B(_3758_),
    .Y(_3761_));
 sg13g2_a22oi_1 _8458_ (.Y(_3762_),
    .B1(_3761_),
    .B2(net2094),
    .A2(net1797),
    .A1(net789));
 sg13g2_nor2_1 _8459_ (.A(net2305),
    .B(_3762_),
    .Y(_0438_));
 sg13g2_nor2_1 _8460_ (.A(_3734_),
    .B(_3758_),
    .Y(_3763_));
 sg13g2_a22oi_1 _8461_ (.Y(_3764_),
    .B1(_3763_),
    .B2(_4026_),
    .A2(net1798),
    .A1(net812));
 sg13g2_nor2_1 _8462_ (.A(net2303),
    .B(net813),
    .Y(_0439_));
 sg13g2_or2_1 _8463_ (.X(_3765_),
    .B(_3754_),
    .A(_4025_));
 sg13g2_nor3_1 _8464_ (.A(net2271),
    .B(\lfsr_inst.lfsr[29] ),
    .C(_3765_),
    .Y(_3766_));
 sg13g2_a22oi_1 _8465_ (.Y(_3767_),
    .B1(_3766_),
    .B2(net2094),
    .A2(net1798),
    .A1(net656));
 sg13g2_nor2_1 _8466_ (.A(net2304),
    .B(net657),
    .Y(_0440_));
 sg13g2_nor2_1 _8467_ (.A(_3732_),
    .B(_3765_),
    .Y(_3768_));
 sg13g2_a22oi_1 _8468_ (.Y(_3769_),
    .B1(_3768_),
    .B2(net2094),
    .A2(net1799),
    .A1(net823));
 sg13g2_nor2_1 _8469_ (.A(net2304),
    .B(_3769_),
    .Y(_0441_));
 sg13g2_nor2_1 _8470_ (.A(_3737_),
    .B(_3765_),
    .Y(_3770_));
 sg13g2_a22oi_1 _8471_ (.Y(_3771_),
    .B1(_3770_),
    .B2(net2094),
    .A2(net1799),
    .A1(net739));
 sg13g2_nor2_1 _8472_ (.A(net2303),
    .B(_3771_),
    .Y(_0442_));
 sg13g2_nor2_1 _8473_ (.A(_3734_),
    .B(_3765_),
    .Y(_3772_));
 sg13g2_a22oi_1 _8474_ (.Y(_3773_),
    .B1(_3772_),
    .B2(net2094),
    .A2(net1797),
    .A1(net593));
 sg13g2_nor2_1 _8475_ (.A(net2305),
    .B(net594),
    .Y(_0443_));
 sg13g2_a21oi_2 _8476_ (.B1(net2094),
    .Y(_3774_),
    .A2(_3744_),
    .A1(_3740_));
 sg13g2_nor4_1 _8477_ (.A(net2271),
    .B(net2270),
    .C(\lfsr_inst.lfsr[30] ),
    .D(net2094),
    .Y(_3775_));
 sg13g2_o21ai_1 _8478_ (.B1(net2325),
    .Y(_3776_),
    .A1(net1797),
    .A2(_3775_));
 sg13g2_a21oi_1 _8479_ (.A1(_3989_),
    .A2(net1797),
    .Y(_0444_),
    .B1(_3776_));
 sg13g2_a22oi_1 _8480_ (.Y(_3777_),
    .B1(_3759_),
    .B2(_3774_),
    .A2(net1799),
    .A1(net733));
 sg13g2_nor2_1 _8481_ (.A(net2305),
    .B(_3777_),
    .Y(_0445_));
 sg13g2_a22oi_1 _8482_ (.Y(_3778_),
    .B1(_3761_),
    .B2(_3774_),
    .A2(net1797),
    .A1(net758));
 sg13g2_nor2_1 _8483_ (.A(net2305),
    .B(_3778_),
    .Y(_0446_));
 sg13g2_a22oi_1 _8484_ (.Y(_3779_),
    .B1(_3763_),
    .B2(_3774_),
    .A2(net1798),
    .A1(net647));
 sg13g2_nor2_1 _8485_ (.A(net2303),
    .B(net648),
    .Y(_0447_));
 sg13g2_a22oi_1 _8486_ (.Y(_3780_),
    .B1(_3766_),
    .B2(_3774_),
    .A2(net1798),
    .A1(net621));
 sg13g2_nor2_1 _8487_ (.A(net2303),
    .B(net622),
    .Y(_0448_));
 sg13g2_a22oi_1 _8488_ (.Y(_3781_),
    .B1(_3768_),
    .B2(_3774_),
    .A2(net1798),
    .A1(net636));
 sg13g2_nor2_1 _8489_ (.A(net2303),
    .B(_3781_),
    .Y(_0449_));
 sg13g2_a22oi_1 _8490_ (.Y(_3782_),
    .B1(_3770_),
    .B2(_3774_),
    .A2(net1799),
    .A1(net613));
 sg13g2_nor2_1 _8491_ (.A(net2303),
    .B(_3782_),
    .Y(_0450_));
 sg13g2_a22oi_1 _8492_ (.Y(_3783_),
    .B1(_3772_),
    .B2(_3774_),
    .A2(net1798),
    .A1(net711));
 sg13g2_nor2_1 _8493_ (.A(net2303),
    .B(net712),
    .Y(_0451_));
 sg13g2_o21ai_1 _8494_ (.B1(net1798),
    .Y(_3784_),
    .A1(net1961),
    .A2(_3747_));
 sg13g2_nor2b_1 _8495_ (.A(_3746_),
    .B_N(_3784_),
    .Y(_3785_));
 sg13g2_nand2_1 _8496_ (.Y(_3786_),
    .A(\welcome_screen_inst.welcome_counter[0] ),
    .B(_3784_));
 sg13g2_nor2b_1 _8497_ (.A(_3785_),
    .B_N(_3786_),
    .Y(_3787_));
 sg13g2_or2_1 _8498_ (.X(_3788_),
    .B(_3784_),
    .A(net997));
 sg13g2_and3_1 _8499_ (.X(_0452_),
    .A(net2325),
    .B(_3787_),
    .C(_3788_));
 sg13g2_a21oi_1 _8500_ (.A1(net627),
    .A2(_3787_),
    .Y(_3789_),
    .B1(net2304));
 sg13g2_o21ai_1 _8501_ (.B1(_3789_),
    .Y(_0453_),
    .A1(net627),
    .A2(_3786_));
 sg13g2_and3_1 _8502_ (.X(_3790_),
    .A(net676),
    .B(\welcome_screen_inst.welcome_counter[1] ),
    .C(\welcome_screen_inst.welcome_counter[0] ));
 sg13g2_a21oi_1 _8503_ (.A1(net627),
    .A2(\welcome_screen_inst.welcome_counter[0] ),
    .Y(_3791_),
    .B1(net676));
 sg13g2_nor3_1 _8504_ (.A(_3747_),
    .B(_3790_),
    .C(_3791_),
    .Y(_3792_));
 sg13g2_a21oi_1 _8505_ (.A1(_3784_),
    .A2(_3792_),
    .Y(_3793_),
    .B1(net2303));
 sg13g2_o21ai_1 _8506_ (.B1(_3793_),
    .Y(_0454_),
    .A1(_3988_),
    .A2(_3784_));
 sg13g2_nand3_1 _8507_ (.B(_3784_),
    .C(_3790_),
    .A(net791),
    .Y(_3794_));
 sg13g2_a21oi_1 _8508_ (.A1(_3784_),
    .A2(_3790_),
    .Y(_3795_),
    .B1(net791));
 sg13g2_nand2_1 _8509_ (.Y(_3796_),
    .A(net1798),
    .B(_3794_));
 sg13g2_o21ai_1 _8510_ (.B1(net2325),
    .Y(_0455_),
    .A1(net792),
    .A2(_3796_));
 sg13g2_nor2b_1 _8511_ (.A(net736),
    .B_N(_3794_),
    .Y(_3797_));
 sg13g2_o21ai_1 _8512_ (.B1(net2331),
    .Y(_0456_),
    .A1(_3785_),
    .A2(net737));
 sg13g2_nor2_1 _8513_ (.A(net2160),
    .B(_0508_),
    .Y(_3798_));
 sg13g2_nor4_1 _8514_ (.A(debug_btn_right),
    .B(net844),
    .C(debug_btn_down),
    .D(debug_btn_left),
    .Y(_3799_));
 sg13g2_o21ai_1 _8515_ (.B1(net2315),
    .Y(_3800_),
    .A1(net849),
    .A2(_3798_));
 sg13g2_a21oi_1 _8516_ (.A1(_3798_),
    .A2(_3799_),
    .Y(_0457_),
    .B1(_3800_));
 sg13g2_nand3_1 _8517_ (.B(_0800_),
    .C(_0802_),
    .A(_0557_),
    .Y(_3801_));
 sg13g2_xor2_1 _8518_ (.B(_0902_),
    .A(_0544_),
    .X(_3802_));
 sg13g2_nand2b_1 _8519_ (.Y(_3803_),
    .B(_0538_),
    .A_N(_0856_));
 sg13g2_or2_1 _8520_ (.X(_3804_),
    .B(_0800_),
    .A(_0557_));
 sg13g2_o21ai_1 _8521_ (.B1(_0561_),
    .Y(_3805_),
    .A1(_0772_),
    .A2(_0773_));
 sg13g2_o21ai_1 _8522_ (.B1(_0562_),
    .Y(_3806_),
    .A1(_0987_),
    .A2(_0988_));
 sg13g2_nand2_1 _8523_ (.Y(_3807_),
    .A(_0540_),
    .B(_0925_));
 sg13g2_o21ai_1 _8524_ (.B1(_0531_),
    .Y(_3808_),
    .A1(_0974_),
    .A2(_0975_));
 sg13g2_a21oi_1 _8525_ (.A1(_0784_),
    .A2(_0785_),
    .Y(_3809_),
    .B1(_0555_));
 sg13g2_o21ai_1 _8526_ (.B1(_0529_),
    .Y(_3810_),
    .A1(_0692_),
    .A2(_0693_));
 sg13g2_xor2_1 _8527_ (.B(_0953_),
    .A(_0546_),
    .X(_3811_));
 sg13g2_nand2_1 _8528_ (.Y(_3812_),
    .A(_0535_),
    .B(_0942_));
 sg13g2_nand2b_1 _8529_ (.Y(_3813_),
    .B(_1006_),
    .A_N(_0556_));
 sg13g2_or2_1 _8530_ (.X(_3814_),
    .B(_0963_),
    .A(_0550_));
 sg13g2_a22oi_1 _8531_ (.Y(_3815_),
    .B1(_0771_),
    .B2(_0564_),
    .A2(_0691_),
    .A1(_0560_));
 sg13g2_nand4_1 _8532_ (.B(_3808_),
    .C(_3810_),
    .A(_3801_),
    .Y(_3816_),
    .D(_3815_));
 sg13g2_a21o_1 _8533_ (.A2(_1007_),
    .A1(_0556_),
    .B1(_3809_),
    .X(_3817_));
 sg13g2_a22oi_1 _8534_ (.Y(_3818_),
    .B1(_0963_),
    .B2(_0550_),
    .A2(_0856_),
    .A1(_0537_));
 sg13g2_nand3_1 _8535_ (.B(_3805_),
    .C(_3818_),
    .A(_3804_),
    .Y(_3819_));
 sg13g2_nand3_1 _8536_ (.B(_3813_),
    .C(_3814_),
    .A(_3802_),
    .Y(_3820_));
 sg13g2_nor4_2 _8537_ (.A(_3816_),
    .B(_3817_),
    .C(_3819_),
    .Y(_3821_),
    .D(_3820_));
 sg13g2_o21ai_1 _8538_ (.B1(_3803_),
    .Y(_3822_),
    .A1(_0535_),
    .A2(_0942_));
 sg13g2_o21ai_1 _8539_ (.B1(_3812_),
    .Y(_3823_),
    .A1(_0540_),
    .A2(_0925_));
 sg13g2_nand3_1 _8540_ (.B(_3807_),
    .C(_3811_),
    .A(_3806_),
    .Y(_3824_));
 sg13g2_nor4_2 _8541_ (.A(\game_logic_inst.valid_move ),
    .B(_3822_),
    .C(_3823_),
    .Y(_3825_),
    .D(_3824_));
 sg13g2_and2_1 _8542_ (.A(_3821_),
    .B(_3825_),
    .X(_3826_));
 sg13g2_or3_1 _8543_ (.A(net2160),
    .B(net1790),
    .C(_0888_),
    .X(_3827_));
 sg13g2_o21ai_1 _8544_ (.B1(net2310),
    .Y(_3828_),
    .A1(net2160),
    .A2(net1808));
 sg13g2_a221oi_1 _8545_ (.B2(_3987_),
    .C1(_3828_),
    .B1(_3827_),
    .A1(net1768),
    .Y(_0458_),
    .A2(_3826_));
 sg13g2_nand3b_1 _8546_ (.B(net2041),
    .C(net2172),
    .Y(_3829_),
    .A_N(net1790));
 sg13g2_a22oi_1 _8547_ (.Y(_3830_),
    .B1(_3829_),
    .B2(net2176),
    .A2(net1809),
    .A1(net2172));
 sg13g2_nor2_1 _8548_ (.A(net2301),
    .B(net966),
    .Y(_0459_));
 sg13g2_and2_1 _8549_ (.A(net2308),
    .B(net444),
    .X(_0460_));
 sg13g2_xor2_1 _8550_ (.B(net967),
    .A(\game_logic_inst.lfsr_shift[0] ),
    .X(_3831_));
 sg13g2_nor2_1 _8551_ (.A(net2301),
    .B(net968),
    .Y(_0461_));
 sg13g2_o21ai_1 _8552_ (.B1(net1808),
    .Y(_3832_),
    .A1(net2275),
    .A2(_3485_));
 sg13g2_a21o_1 _8553_ (.A2(_3832_),
    .A1(net2313),
    .B1(_0511_),
    .X(_0462_));
 sg13g2_or4_1 _8554_ (.A(net2160),
    .B(_0747_),
    .C(_0748_),
    .D(net2033),
    .X(_3833_));
 sg13g2_nand4_1 _8555_ (.B(net2170),
    .C(_0069_),
    .A(_3986_),
    .Y(_3834_),
    .D(_0747_));
 sg13g2_a21oi_1 _8556_ (.A1(_3833_),
    .A2(_3834_),
    .Y(_3835_),
    .B1(net1809));
 sg13g2_nor3_1 _8557_ (.A(net2099),
    .B(net2041),
    .C(net1759),
    .Y(_3836_));
 sg13g2_nor2_1 _8558_ (.A(net2170),
    .B(_3832_),
    .Y(_3837_));
 sg13g2_nor2_1 _8559_ (.A(net2160),
    .B(net1794),
    .Y(_3838_));
 sg13g2_nor4_2 _8560_ (.A(_3835_),
    .B(_3836_),
    .C(_3837_),
    .Y(_3839_),
    .D(_3838_));
 sg13g2_a21oi_1 _8561_ (.A1(_3821_),
    .A2(_3825_),
    .Y(_3840_),
    .B1(net849));
 sg13g2_a21oi_1 _8562_ (.A1(net896),
    .A2(_3986_),
    .Y(_3841_),
    .B1(net2099));
 sg13g2_o21ai_1 _8563_ (.B1(_3841_),
    .Y(_3842_),
    .A1(_3986_),
    .A2(_3840_));
 sg13g2_o21ai_1 _8564_ (.B1(net2312),
    .Y(_3843_),
    .A1(net896),
    .A2(_3839_));
 sg13g2_a21oi_1 _8565_ (.A1(_3839_),
    .A2(_3842_),
    .Y(_0463_),
    .B1(_3843_));
 sg13g2_xnor2_1 _8566_ (.Y(_3844_),
    .A(\game_logic_inst.add_new_tiles[1] ),
    .B(\game_logic_inst.add_new_tiles[0] ));
 sg13g2_a21oi_1 _8567_ (.A1(net567),
    .A2(_3844_),
    .Y(_3845_),
    .B1(net2160));
 sg13g2_o21ai_1 _8568_ (.B1(net2312),
    .Y(_3846_),
    .A1(\game_logic_inst.add_new_tiles[1] ),
    .A2(_3839_));
 sg13g2_a21oi_1 _8569_ (.A1(_3839_),
    .A2(net568),
    .Y(_0464_),
    .B1(_3846_));
 sg13g2_nand3_1 _8570_ (.B(_0750_),
    .C(_0888_),
    .A(_0511_),
    .Y(_3847_));
 sg13g2_nor2b_2 _8571_ (.A(_3847_),
    .B_N(_0704_),
    .Y(_0465_));
 sg13g2_nor2b_2 _8572_ (.A(_3847_),
    .B_N(_0703_),
    .Y(_0466_));
 sg13g2_nor2_2 _8573_ (.A(_0702_),
    .B(_3847_),
    .Y(_0467_));
 sg13g2_nor2_2 _8574_ (.A(_0700_),
    .B(_3847_),
    .Y(_0468_));
 sg13g2_nand2_1 _8575_ (.Y(_3848_),
    .A(net8),
    .B(net11));
 sg13g2_nand2b_2 _8576_ (.Y(_3849_),
    .B(_3848_),
    .A_N(net12));
 sg13g2_nand2_1 _8577_ (.Y(_3850_),
    .A(net9),
    .B(net8));
 sg13g2_nor3_2 _8578_ (.A(net10),
    .B(_3849_),
    .C(_3850_),
    .Y(_3851_));
 sg13g2_and2_1 _8579_ (.A(net2319),
    .B(net1843),
    .X(_0469_));
 sg13g2_nand3_1 _8580_ (.B(_0500_),
    .C(net1809),
    .A(_0498_),
    .Y(_3852_));
 sg13g2_a21oi_1 _8581_ (.A1(net2170),
    .A2(_3852_),
    .Y(_3853_),
    .B1(net856));
 sg13g2_nor2_1 _8582_ (.A(\game_logic_inst.current_direction[3] ),
    .B(net555),
    .Y(_3854_));
 sg13g2_nand3b_1 _8583_ (.B(net2043),
    .C(_0069_),
    .Y(_3855_),
    .A_N(net567));
 sg13g2_o21ai_1 _8584_ (.B1(net2170),
    .Y(_3856_),
    .A1(_3854_),
    .A2(_3855_));
 sg13g2_o21ai_1 _8585_ (.B1(net2313),
    .Y(_3857_),
    .A1(net1809),
    .A2(_3856_));
 sg13g2_nor2_1 _8586_ (.A(_3853_),
    .B(_3857_),
    .Y(_0470_));
 sg13g2_nor2_1 _8587_ (.A(net2160),
    .B(net1760),
    .Y(_3858_));
 sg13g2_a22oi_1 _8588_ (.Y(_3859_),
    .B1(_3858_),
    .B2(net582),
    .A2(_3827_),
    .A1(net2157));
 sg13g2_nor2_1 _8589_ (.A(net2301),
    .B(net583),
    .Y(_0471_));
 sg13g2_nor4_1 _8590_ (.A(net2160),
    .B(net2060),
    .C(net2041),
    .D(net1760),
    .Y(_3860_));
 sg13g2_a21oi_1 _8591_ (.A1(net2153),
    .A2(_3827_),
    .Y(_3861_),
    .B1(_3860_));
 sg13g2_nor2_1 _8592_ (.A(net2301),
    .B(_3861_),
    .Y(_0472_));
 sg13g2_mux4_1 _8593_ (.S0(net2132),
    .A0(\debug_controller_inst.grid_in[32] ),
    .A1(\debug_controller_inst.grid_in[36] ),
    .A2(\debug_controller_inst.grid_in[40] ),
    .A3(\debug_controller_inst.grid_in[44] ),
    .S1(net2128),
    .X(_3862_));
 sg13g2_nor2_1 _8594_ (.A(net2125),
    .B(_3862_),
    .Y(_3863_));
 sg13g2_o21ai_1 _8595_ (.B1(net2124),
    .Y(_3864_),
    .A1(net2131),
    .A2(\debug_controller_inst.grid_in[48] ));
 sg13g2_a21oi_1 _8596_ (.A1(net2131),
    .A2(_4028_),
    .Y(_3865_),
    .B1(_3864_));
 sg13g2_nor2_1 _8597_ (.A(net2131),
    .B(\debug_controller_inst.grid_in[56] ),
    .Y(_3866_));
 sg13g2_o21ai_1 _8598_ (.B1(net2128),
    .Y(_3867_),
    .A1(net2123),
    .A2(\debug_controller_inst.grid_in[60] ));
 sg13g2_o21ai_1 _8599_ (.B1(net2126),
    .Y(_3868_),
    .A1(_3866_),
    .A2(_3867_));
 sg13g2_o21ai_1 _8600_ (.B1(\debug_controller_inst.grid_addr[3] ),
    .Y(_3869_),
    .A1(_3865_),
    .A2(_3868_));
 sg13g2_mux4_1 _8601_ (.S0(net2131),
    .A0(\debug_controller_inst.grid_in[0] ),
    .A1(\debug_controller_inst.grid_in[4] ),
    .A2(\debug_controller_inst.grid_in[8] ),
    .A3(\debug_controller_inst.grid_in[12] ),
    .S1(net2129),
    .X(_3870_));
 sg13g2_nor2_1 _8602_ (.A(net2125),
    .B(_3870_),
    .Y(_3871_));
 sg13g2_o21ai_1 _8603_ (.B1(net2124),
    .Y(_3872_),
    .A1(net2131),
    .A2(\debug_controller_inst.grid_in[16] ));
 sg13g2_a21oi_1 _8604_ (.A1(net2133),
    .A2(_4027_),
    .Y(_3873_),
    .B1(_3872_));
 sg13g2_nor2_1 _8605_ (.A(net2123),
    .B(\debug_controller_inst.grid_in[28] ),
    .Y(_3874_));
 sg13g2_o21ai_1 _8606_ (.B1(net2128),
    .Y(_3875_),
    .A1(net2131),
    .A2(\debug_controller_inst.grid_in[24] ));
 sg13g2_o21ai_1 _8607_ (.B1(net2125),
    .Y(_3876_),
    .A1(_3874_),
    .A2(_3875_));
 sg13g2_o21ai_1 _8608_ (.B1(_3975_),
    .Y(_3877_),
    .A1(_3873_),
    .A2(_3876_));
 sg13g2_nor2_1 _8609_ (.A(_3871_),
    .B(_3877_),
    .Y(_3878_));
 sg13g2_o21ai_1 _8610_ (.B1(_3851_),
    .Y(_3879_),
    .A1(_3863_),
    .A2(_3869_));
 sg13g2_nor2_2 _8611_ (.A(_3878_),
    .B(_3879_),
    .Y(_3880_));
 sg13g2_o21ai_1 _8612_ (.B1(net2318),
    .Y(_3881_),
    .A1(net855),
    .A2(net1843));
 sg13g2_nor2_1 _8613_ (.A(_3880_),
    .B(_3881_),
    .Y(_0473_));
 sg13g2_mux4_1 _8614_ (.S0(net2132),
    .A0(\debug_controller_inst.grid_in[33] ),
    .A1(\debug_controller_inst.grid_in[37] ),
    .A2(\debug_controller_inst.grid_in[41] ),
    .A3(\debug_controller_inst.grid_in[45] ),
    .S1(net2128),
    .X(_3882_));
 sg13g2_nor2_1 _8615_ (.A(net2125),
    .B(_3882_),
    .Y(_3883_));
 sg13g2_o21ai_1 _8616_ (.B1(net2124),
    .Y(_3884_),
    .A1(net2132),
    .A2(\debug_controller_inst.grid_in[49] ));
 sg13g2_a21oi_1 _8617_ (.A1(net2132),
    .A2(_4030_),
    .Y(_3885_),
    .B1(_3884_));
 sg13g2_nor2_1 _8618_ (.A(net2132),
    .B(\debug_controller_inst.grid_in[57] ),
    .Y(_3886_));
 sg13g2_o21ai_1 _8619_ (.B1(net2129),
    .Y(_3887_),
    .A1(net2123),
    .A2(\debug_controller_inst.grid_in[61] ));
 sg13g2_o21ai_1 _8620_ (.B1(net2125),
    .Y(_3888_),
    .A1(_3886_),
    .A2(_3887_));
 sg13g2_o21ai_1 _8621_ (.B1(\debug_controller_inst.grid_addr[3] ),
    .Y(_3889_),
    .A1(_3885_),
    .A2(_3888_));
 sg13g2_mux4_1 _8622_ (.S0(net2132),
    .A0(\debug_controller_inst.grid_in[1] ),
    .A1(\debug_controller_inst.grid_in[5] ),
    .A2(\debug_controller_inst.grid_in[9] ),
    .A3(\debug_controller_inst.grid_in[13] ),
    .S1(net2128),
    .X(_3890_));
 sg13g2_nor2_1 _8623_ (.A(net2125),
    .B(_3890_),
    .Y(_3891_));
 sg13g2_o21ai_1 _8624_ (.B1(net2124),
    .Y(_3892_),
    .A1(net2133),
    .A2(\debug_controller_inst.grid_in[17] ));
 sg13g2_a21oi_1 _8625_ (.A1(net2133),
    .A2(_4029_),
    .Y(_3893_),
    .B1(_3892_));
 sg13g2_nor2_1 _8626_ (.A(net2123),
    .B(\debug_controller_inst.grid_in[29] ),
    .Y(_3894_));
 sg13g2_o21ai_1 _8627_ (.B1(net2129),
    .Y(_3895_),
    .A1(net2132),
    .A2(\debug_controller_inst.grid_in[25] ));
 sg13g2_o21ai_1 _8628_ (.B1(net2125),
    .Y(_3896_),
    .A1(_3894_),
    .A2(_3895_));
 sg13g2_o21ai_1 _8629_ (.B1(_3975_),
    .Y(_3897_),
    .A1(_3893_),
    .A2(_3896_));
 sg13g2_nor2_1 _8630_ (.A(_3891_),
    .B(_3897_),
    .Y(_3898_));
 sg13g2_o21ai_1 _8631_ (.B1(net1843),
    .Y(_3899_),
    .A1(_3883_),
    .A2(_3889_));
 sg13g2_nor2_2 _8632_ (.A(_3898_),
    .B(_3899_),
    .Y(_3900_));
 sg13g2_o21ai_1 _8633_ (.B1(net2318),
    .Y(_3901_),
    .A1(net919),
    .A2(net1843));
 sg13g2_nor2_1 _8634_ (.A(_3900_),
    .B(_3901_),
    .Y(_0474_));
 sg13g2_mux4_1 _8635_ (.S0(net2135),
    .A0(\debug_controller_inst.grid_in[34] ),
    .A1(\debug_controller_inst.grid_in[38] ),
    .A2(\debug_controller_inst.grid_in[42] ),
    .A3(\debug_controller_inst.grid_in[46] ),
    .S1(net2130),
    .X(_3902_));
 sg13g2_nor2_1 _8636_ (.A(net2127),
    .B(_3902_),
    .Y(_3903_));
 sg13g2_o21ai_1 _8637_ (.B1(net2124),
    .Y(_3904_),
    .A1(net2135),
    .A2(\debug_controller_inst.grid_in[50] ));
 sg13g2_a21oi_1 _8638_ (.A1(net2135),
    .A2(_4032_),
    .Y(_3905_),
    .B1(_3904_));
 sg13g2_nor2_1 _8639_ (.A(net2135),
    .B(\debug_controller_inst.grid_in[58] ),
    .Y(_3906_));
 sg13g2_o21ai_1 _8640_ (.B1(net2130),
    .Y(_3907_),
    .A1(_3978_),
    .A2(\debug_controller_inst.grid_in[62] ));
 sg13g2_o21ai_1 _8641_ (.B1(net2127),
    .Y(_3908_),
    .A1(_3906_),
    .A2(_3907_));
 sg13g2_o21ai_1 _8642_ (.B1(\debug_controller_inst.grid_addr[3] ),
    .Y(_3909_),
    .A1(_3905_),
    .A2(_3908_));
 sg13g2_mux4_1 _8643_ (.S0(net2135),
    .A0(\debug_controller_inst.grid_in[2] ),
    .A1(\debug_controller_inst.grid_in[6] ),
    .A2(\debug_controller_inst.grid_in[10] ),
    .A3(\debug_controller_inst.grid_in[14] ),
    .S1(net2130),
    .X(_3910_));
 sg13g2_nor2_1 _8644_ (.A(net2127),
    .B(_3910_),
    .Y(_3911_));
 sg13g2_o21ai_1 _8645_ (.B1(_3977_),
    .Y(_3912_),
    .A1(net2135),
    .A2(\debug_controller_inst.grid_in[18] ));
 sg13g2_a21oi_1 _8646_ (.A1(net2135),
    .A2(_4031_),
    .Y(_3913_),
    .B1(_3912_));
 sg13g2_nor2_1 _8647_ (.A(net2123),
    .B(\debug_controller_inst.grid_in[30] ),
    .Y(_3914_));
 sg13g2_o21ai_1 _8648_ (.B1(net2130),
    .Y(_3915_),
    .A1(net2135),
    .A2(\debug_controller_inst.grid_in[26] ));
 sg13g2_o21ai_1 _8649_ (.B1(net2127),
    .Y(_3916_),
    .A1(_3914_),
    .A2(_3915_));
 sg13g2_o21ai_1 _8650_ (.B1(_3975_),
    .Y(_3917_),
    .A1(_3913_),
    .A2(_3916_));
 sg13g2_nor2_1 _8651_ (.A(_3911_),
    .B(_3917_),
    .Y(_3918_));
 sg13g2_o21ai_1 _8652_ (.B1(net1843),
    .Y(_3919_),
    .A1(_3903_),
    .A2(_3909_));
 sg13g2_nor2_1 _8653_ (.A(_3918_),
    .B(_3919_),
    .Y(_3920_));
 sg13g2_o21ai_1 _8654_ (.B1(net2319),
    .Y(_3921_),
    .A1(net830),
    .A2(net1843));
 sg13g2_nor2_1 _8655_ (.A(_3920_),
    .B(_3921_),
    .Y(_0475_));
 sg13g2_mux4_1 _8656_ (.S0(net2134),
    .A0(\debug_controller_inst.grid_in[35] ),
    .A1(\debug_controller_inst.grid_in[39] ),
    .A2(\debug_controller_inst.grid_in[43] ),
    .A3(\debug_controller_inst.grid_in[47] ),
    .S1(net2128),
    .X(_3922_));
 sg13g2_nor2_1 _8657_ (.A(net2126),
    .B(_3922_),
    .Y(_3923_));
 sg13g2_o21ai_1 _8658_ (.B1(net2124),
    .Y(_3924_),
    .A1(net2134),
    .A2(\debug_controller_inst.grid_in[51] ));
 sg13g2_a21oi_1 _8659_ (.A1(net2134),
    .A2(_4034_),
    .Y(_3925_),
    .B1(_3924_));
 sg13g2_nor2_1 _8660_ (.A(net2134),
    .B(\debug_controller_inst.grid_in[59] ),
    .Y(_3926_));
 sg13g2_o21ai_1 _8661_ (.B1(net2128),
    .Y(_3927_),
    .A1(net2123),
    .A2(\debug_controller_inst.grid_in[63] ));
 sg13g2_o21ai_1 _8662_ (.B1(net2126),
    .Y(_3928_),
    .A1(_3926_),
    .A2(_3927_));
 sg13g2_o21ai_1 _8663_ (.B1(\debug_controller_inst.grid_addr[3] ),
    .Y(_3929_),
    .A1(_3925_),
    .A2(_3928_));
 sg13g2_mux4_1 _8664_ (.S0(net2132),
    .A0(\debug_controller_inst.grid_in[3] ),
    .A1(\debug_controller_inst.grid_in[7] ),
    .A2(\debug_controller_inst.grid_in[11] ),
    .A3(\debug_controller_inst.grid_in[15] ),
    .S1(net2129),
    .X(_3930_));
 sg13g2_nor2_1 _8665_ (.A(net2125),
    .B(_3930_),
    .Y(_3931_));
 sg13g2_o21ai_1 _8666_ (.B1(net2124),
    .Y(_3932_),
    .A1(net2131),
    .A2(\debug_controller_inst.grid_in[19] ));
 sg13g2_a21oi_1 _8667_ (.A1(net2131),
    .A2(_4033_),
    .Y(_3933_),
    .B1(_3932_));
 sg13g2_nor2_1 _8668_ (.A(net2123),
    .B(\debug_controller_inst.grid_in[31] ),
    .Y(_3934_));
 sg13g2_o21ai_1 _8669_ (.B1(net2128),
    .Y(_3935_),
    .A1(net2134),
    .A2(\debug_controller_inst.grid_in[27] ));
 sg13g2_o21ai_1 _8670_ (.B1(net2126),
    .Y(_3936_),
    .A1(_3934_),
    .A2(_3935_));
 sg13g2_o21ai_1 _8671_ (.B1(_3975_),
    .Y(_3937_),
    .A1(_3933_),
    .A2(_3936_));
 sg13g2_nor2_1 _8672_ (.A(_3931_),
    .B(_3937_),
    .Y(_3938_));
 sg13g2_o21ai_1 _8673_ (.B1(net1843),
    .Y(_3939_),
    .A1(_3923_),
    .A2(_3929_));
 sg13g2_nor2_2 _8674_ (.A(_3938_),
    .B(_3939_),
    .Y(_3940_));
 sg13g2_o21ai_1 _8675_ (.B1(net2319),
    .Y(_3941_),
    .A1(net890),
    .A2(net1843));
 sg13g2_nor2_1 _8676_ (.A(_3940_),
    .B(_3941_),
    .Y(_0476_));
 sg13g2_nand2_1 _8677_ (.Y(_3942_),
    .A(net8),
    .B(net10));
 sg13g2_nand2_1 _8678_ (.Y(_3943_),
    .A(_3850_),
    .B(_3942_));
 sg13g2_nor4_2 _8679_ (.A(net12),
    .B(net2302),
    .C(_3848_),
    .Y(_3944_),
    .D(_3943_));
 sg13g2_and2_2 _8680_ (.A(net13),
    .B(_3944_),
    .X(_0477_));
 sg13g2_and2_1 _8681_ (.A(net14),
    .B(_3944_),
    .X(_0478_));
 sg13g2_and2_2 _8682_ (.A(net15),
    .B(_3944_),
    .X(_0479_));
 sg13g2_and2_1 _8683_ (.A(net16),
    .B(_3944_),
    .X(_0480_));
 sg13g2_nor3_2 _8684_ (.A(net9),
    .B(_3849_),
    .C(_3942_),
    .Y(_3945_));
 sg13g2_and2_1 _8685_ (.A(net2321),
    .B(net1841),
    .X(_0481_));
 sg13g2_o21ai_1 _8686_ (.B1(net2323),
    .Y(_3946_),
    .A1(net937),
    .A2(_3945_));
 sg13g2_a21oi_1 _8687_ (.A1(_3985_),
    .A2(_3945_),
    .Y(_0482_),
    .B1(_3946_));
 sg13g2_o21ai_1 _8688_ (.B1(net2322),
    .Y(_3947_),
    .A1(net2147),
    .A2(net1842));
 sg13g2_a21oi_1 _8689_ (.A1(_3983_),
    .A2(net1842),
    .Y(_0483_),
    .B1(_3947_));
 sg13g2_o21ai_1 _8690_ (.B1(net2323),
    .Y(_3948_),
    .A1(net2144),
    .A2(net1842));
 sg13g2_a21oi_1 _8691_ (.A1(_3981_),
    .A2(net1842),
    .Y(_0484_),
    .B1(_3948_));
 sg13g2_o21ai_1 _8692_ (.B1(net2321),
    .Y(_3949_),
    .A1(net2142),
    .A2(net1841));
 sg13g2_a21oi_1 _8693_ (.A1(_3980_),
    .A2(net1842),
    .Y(_0485_),
    .B1(_3949_));
 sg13g2_o21ai_1 _8694_ (.B1(net2321),
    .Y(_3950_),
    .A1(net725),
    .A2(net1841));
 sg13g2_a21oi_1 _8695_ (.A1(_3978_),
    .A2(net1841),
    .Y(_0486_),
    .B1(_3950_));
 sg13g2_o21ai_1 _8696_ (.B1(net2321),
    .Y(_3951_),
    .A1(net690),
    .A2(net1841));
 sg13g2_a21oi_1 _8697_ (.A1(_3977_),
    .A2(net1841),
    .Y(_0487_),
    .B1(_3951_));
 sg13g2_o21ai_1 _8698_ (.B1(net2321),
    .Y(_3952_),
    .A1(net816),
    .A2(net1842));
 sg13g2_a21oi_1 _8699_ (.A1(_3976_),
    .A2(net1842),
    .Y(_0488_),
    .B1(_3952_));
 sg13g2_o21ai_1 _8700_ (.B1(net2321),
    .Y(_3953_),
    .A1(net988),
    .A2(net1841));
 sg13g2_a21oi_1 _8701_ (.A1(_3975_),
    .A2(net1841),
    .Y(_0489_),
    .B1(_3953_));
 sg13g2_and2_1 _8702_ (.A(net2326),
    .B(net990),
    .X(_0490_));
 sg13g2_nor2b_2 _8703_ (.A(_3849_),
    .B_N(_3943_),
    .Y(_3954_));
 sg13g2_nand2b_1 _8704_ (.Y(_3955_),
    .B(_3943_),
    .A_N(_3849_));
 sg13g2_and3_2 _8705_ (.X(_3956_),
    .A(net9),
    .B(net8),
    .C(net10));
 sg13g2_nand2b_2 _8706_ (.Y(_3957_),
    .B(_3956_),
    .A_N(_3849_));
 sg13g2_inv_1 _8707_ (.Y(_3958_),
    .A(_3957_));
 sg13g2_nor2_1 _8708_ (.A(net13),
    .B(_3957_),
    .Y(_3959_));
 sg13g2_nor2_1 _8709_ (.A(net893),
    .B(_3956_),
    .Y(_3960_));
 sg13g2_o21ai_1 _8710_ (.B1(_3954_),
    .Y(_3961_),
    .A1(_3959_),
    .A2(_3960_));
 sg13g2_o21ai_1 _8711_ (.B1(_3961_),
    .Y(_3962_),
    .A1(net2136),
    .A2(_3954_));
 sg13g2_nor2_1 _8712_ (.A(net2302),
    .B(net894),
    .Y(_0491_));
 sg13g2_nor2_1 _8713_ (.A(_3977_),
    .B(net2123),
    .Y(_3963_));
 sg13g2_o21ai_1 _8714_ (.B1(_3954_),
    .Y(_3964_),
    .A1(_3956_),
    .A2(_3963_));
 sg13g2_nor2_1 _8715_ (.A(_3983_),
    .B(_3957_),
    .Y(_3965_));
 sg13g2_o21ai_1 _8716_ (.B1(_3954_),
    .Y(_3966_),
    .A1(net2136),
    .A2(_3956_));
 sg13g2_o21ai_1 _8717_ (.B1(net2323),
    .Y(_3967_),
    .A1(_3964_),
    .A2(_3965_));
 sg13g2_a21oi_1 _8718_ (.A1(net2124),
    .A2(_3966_),
    .Y(_0492_),
    .B1(_3967_));
 sg13g2_a21o_1 _8719_ (.A2(_3963_),
    .A1(net2127),
    .B1(_3958_),
    .X(_3968_));
 sg13g2_a21oi_1 _8720_ (.A1(net15),
    .A2(_3956_),
    .Y(_3969_),
    .B1(_3955_));
 sg13g2_a221oi_1 _8721_ (.B2(_3969_),
    .C1(net2302),
    .B1(_3968_),
    .A1(_3976_),
    .Y(_0493_),
    .A2(_3964_));
 sg13g2_nand2_1 _8722_ (.Y(_3970_),
    .A(net955),
    .B(_3955_));
 sg13g2_nand2b_1 _8723_ (.Y(_3971_),
    .B(_3963_),
    .A_N(_0164_));
 sg13g2_xnor2_1 _8724_ (.Y(_3972_),
    .A(_3975_),
    .B(_3971_));
 sg13g2_a22oi_1 _8725_ (.Y(_3973_),
    .B1(_3957_),
    .B2(_3972_),
    .A2(_3956_),
    .A1(_3980_));
 sg13g2_nand2_1 _8726_ (.Y(_3974_),
    .A(_3954_),
    .B(_3973_));
 sg13g2_a21oi_1 _8727_ (.A1(_3970_),
    .A2(_3974_),
    .Y(_0494_),
    .B1(net2302));
 sg13g2_dfrbp_1 _8728_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net214),
    .D(_0175_),
    .Q_N(_4355_),
    .Q(vsync_prev));
 sg13g2_dfrbp_1 _8729_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net173),
    .D(_0176_),
    .Q_N(_0174_),
    .Q(\draw_game_inst.board_x[0] ));
 sg13g2_dfrbp_1 _8730_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net172),
    .D(_0177_),
    .Q_N(_4354_),
    .Q(\draw_game_inst.board_x[1] ));
 sg13g2_dfrbp_1 _8731_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net171),
    .D(_0178_),
    .Q_N(_4353_),
    .Q(\draw_game_inst.board_x[2] ));
 sg13g2_dfrbp_1 _8732_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net170),
    .D(_0179_),
    .Q_N(_0095_),
    .Q(\draw_game_inst.board_x[3] ));
 sg13g2_dfrbp_1 _8733_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net169),
    .D(_0180_),
    .Q_N(_0096_),
    .Q(\draw_game_inst.board_x[4] ));
 sg13g2_dfrbp_1 _8734_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net168),
    .D(_0181_),
    .Q_N(_0094_),
    .Q(\draw_game_inst.board_x[5] ));
 sg13g2_dfrbp_1 _8735_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net167),
    .D(_0182_),
    .Q_N(_4352_),
    .Q(\draw_game_inst.x[6] ));
 sg13g2_dfrbp_1 _8736_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net166),
    .D(_0183_),
    .Q_N(_4351_),
    .Q(\draw_game_inst.x[7] ));
 sg13g2_dfrbp_1 _8737_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net165),
    .D(_0184_),
    .Q_N(_4350_),
    .Q(\draw_game_inst.x[8] ));
 sg13g2_dfrbp_1 _8738_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net164),
    .D(_0185_),
    .Q_N(_4349_),
    .Q(\draw_game_inst.x[9] ));
 sg13g2_dfrbp_1 _8739_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net163),
    .D(_0186_),
    .Q_N(_4348_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _8740_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net162),
    .D(_0187_),
    .Q_N(_4347_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _8741_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net161),
    .D(net1010),
    .Q_N(_4346_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _8742_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net160),
    .D(_0189_),
    .Q_N(_4345_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _8743_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net159),
    .D(_0190_),
    .Q_N(_4344_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _8744_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net158),
    .D(_0191_),
    .Q_N(_4343_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _8745_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net157),
    .D(net704),
    .Q_N(_4342_),
    .Q(\draw_game_inst.grid[0] ));
 sg13g2_dfrbp_1 _8746_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net155),
    .D(net747),
    .Q_N(_4341_),
    .Q(\draw_game_inst.grid[1] ));
 sg13g2_dfrbp_1 _8747_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net153),
    .D(net728),
    .Q_N(_4340_),
    .Q(\draw_game_inst.grid[2] ));
 sg13g2_dfrbp_1 _8748_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net151),
    .D(net654),
    .Q_N(_4339_),
    .Q(\draw_game_inst.grid[3] ));
 sg13g2_dfrbp_1 _8749_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net149),
    .D(net695),
    .Q_N(_4338_),
    .Q(\draw_game_inst.grid[4] ));
 sg13g2_dfrbp_1 _8750_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net147),
    .D(net782),
    .Q_N(_4337_),
    .Q(\draw_game_inst.grid[5] ));
 sg13g2_dfrbp_1 _8751_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net145),
    .D(net706),
    .Q_N(_4336_),
    .Q(\draw_game_inst.grid[6] ));
 sg13g2_dfrbp_1 _8752_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net143),
    .D(net708),
    .Q_N(_4335_),
    .Q(\draw_game_inst.grid[7] ));
 sg13g2_dfrbp_1 _8753_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net141),
    .D(_0200_),
    .Q_N(_4334_),
    .Q(\draw_game_inst.grid[8] ));
 sg13g2_dfrbp_1 _8754_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net139),
    .D(net854),
    .Q_N(_4333_),
    .Q(\draw_game_inst.grid[9] ));
 sg13g2_dfrbp_1 _8755_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net137),
    .D(_0202_),
    .Q_N(_4332_),
    .Q(\draw_game_inst.grid[10] ));
 sg13g2_dfrbp_1 _8756_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net135),
    .D(net662),
    .Q_N(_4331_),
    .Q(\draw_game_inst.grid[11] ));
 sg13g2_dfrbp_1 _8757_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net133),
    .D(net749),
    .Q_N(_4330_),
    .Q(\draw_game_inst.grid[12] ));
 sg13g2_dfrbp_1 _8758_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net131),
    .D(net815),
    .Q_N(_4329_),
    .Q(\draw_game_inst.grid[13] ));
 sg13g2_dfrbp_1 _8759_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net129),
    .D(net722),
    .Q_N(_4328_),
    .Q(\draw_game_inst.grid[14] ));
 sg13g2_dfrbp_1 _8760_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net127),
    .D(net670),
    .Q_N(_4327_),
    .Q(\draw_game_inst.grid[15] ));
 sg13g2_dfrbp_1 _8761_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net125),
    .D(net796),
    .Q_N(_4326_),
    .Q(\draw_game_inst.grid[16] ));
 sg13g2_dfrbp_1 _8762_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net123),
    .D(net763),
    .Q_N(_4325_),
    .Q(\draw_game_inst.grid[17] ));
 sg13g2_dfrbp_1 _8763_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net121),
    .D(net735),
    .Q_N(_4324_),
    .Q(\draw_game_inst.grid[18] ));
 sg13g2_dfrbp_1 _8764_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net119),
    .D(net686),
    .Q_N(_4323_),
    .Q(\draw_game_inst.grid[19] ));
 sg13g2_dfrbp_1 _8765_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net117),
    .D(net760),
    .Q_N(_4322_),
    .Q(\draw_game_inst.grid[20] ));
 sg13g2_dfrbp_1 _8766_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net115),
    .D(net776),
    .Q_N(_4321_),
    .Q(\draw_game_inst.grid[21] ));
 sg13g2_dfrbp_1 _8767_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net113),
    .D(net684),
    .Q_N(_4320_),
    .Q(\draw_game_inst.grid[22] ));
 sg13g2_dfrbp_1 _8768_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net111),
    .D(net786),
    .Q_N(_4319_),
    .Q(\draw_game_inst.grid[23] ));
 sg13g2_dfrbp_1 _8769_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net109),
    .D(net702),
    .Q_N(_4318_),
    .Q(\draw_game_inst.grid[24] ));
 sg13g2_dfrbp_1 _8770_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net107),
    .D(net780),
    .Q_N(_4317_),
    .Q(\draw_game_inst.grid[25] ));
 sg13g2_dfrbp_1 _8771_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net105),
    .D(net720),
    .Q_N(_4316_),
    .Q(\draw_game_inst.grid[26] ));
 sg13g2_dfrbp_1 _8772_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net103),
    .D(net751),
    .Q_N(_4315_),
    .Q(\draw_game_inst.grid[27] ));
 sg13g2_dfrbp_1 _8773_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net101),
    .D(net700),
    .Q_N(_4314_),
    .Q(\draw_game_inst.grid[28] ));
 sg13g2_dfrbp_1 _8774_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net99),
    .D(net769),
    .Q_N(_4313_),
    .Q(\draw_game_inst.grid[29] ));
 sg13g2_dfrbp_1 _8775_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net97),
    .D(net832),
    .Q_N(_4312_),
    .Q(\draw_game_inst.grid[30] ));
 sg13g2_dfrbp_1 _8776_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net95),
    .D(net693),
    .Q_N(_4311_),
    .Q(\draw_game_inst.grid[31] ));
 sg13g2_dfrbp_1 _8777_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net93),
    .D(net825),
    .Q_N(_4310_),
    .Q(\draw_game_inst.grid[32] ));
 sg13g2_dfrbp_1 _8778_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net91),
    .D(_0225_),
    .Q_N(_4309_),
    .Q(\draw_game_inst.grid[33] ));
 sg13g2_dfrbp_1 _8779_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net89),
    .D(net710),
    .Q_N(_4308_),
    .Q(\draw_game_inst.grid[34] ));
 sg13g2_dfrbp_1 _8780_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net87),
    .D(net745),
    .Q_N(_4307_),
    .Q(\draw_game_inst.grid[35] ));
 sg13g2_dfrbp_1 _8781_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net85),
    .D(net753),
    .Q_N(_4306_),
    .Q(\draw_game_inst.grid[36] ));
 sg13g2_dfrbp_1 _8782_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net83),
    .D(net778),
    .Q_N(_4305_),
    .Q(\draw_game_inst.grid[37] ));
 sg13g2_dfrbp_1 _8783_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net81),
    .D(net835),
    .Q_N(_4304_),
    .Q(\draw_game_inst.grid[38] ));
 sg13g2_dfrbp_1 _8784_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net79),
    .D(net730),
    .Q_N(_4303_),
    .Q(\draw_game_inst.grid[39] ));
 sg13g2_dfrbp_1 _8785_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net77),
    .D(net799),
    .Q_N(_4302_),
    .Q(\draw_game_inst.grid[40] ));
 sg13g2_dfrbp_1 _8786_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net75),
    .D(net806),
    .Q_N(_4301_),
    .Q(\draw_game_inst.grid[41] ));
 sg13g2_dfrbp_1 _8787_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net73),
    .D(net675),
    .Q_N(_4300_),
    .Q(\draw_game_inst.grid[42] ));
 sg13g2_dfrbp_1 _8788_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net71),
    .D(net822),
    .Q_N(_4299_),
    .Q(\draw_game_inst.grid[43] ));
 sg13g2_dfrbp_1 _8789_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net69),
    .D(net794),
    .Q_N(_4298_),
    .Q(\draw_game_inst.grid[44] ));
 sg13g2_dfrbp_1 _8790_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net67),
    .D(net809),
    .Q_N(_4297_),
    .Q(\draw_game_inst.grid[45] ));
 sg13g2_dfrbp_1 _8791_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net65),
    .D(net697),
    .Q_N(_4296_),
    .Q(\draw_game_inst.grid[46] ));
 sg13g2_dfrbp_1 _8792_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net63),
    .D(net765),
    .Q_N(_4295_),
    .Q(\draw_game_inst.grid[47] ));
 sg13g2_dfrbp_1 _8793_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net61),
    .D(net689),
    .Q_N(_4294_),
    .Q(\draw_game_inst.grid[48] ));
 sg13g2_dfrbp_1 _8794_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net59),
    .D(net827),
    .Q_N(_4293_),
    .Q(\draw_game_inst.grid[49] ));
 sg13g2_dfrbp_1 _8795_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net57),
    .D(net784),
    .Q_N(_4292_),
    .Q(\draw_game_inst.grid[50] ));
 sg13g2_dfrbp_1 _8796_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net55),
    .D(net652),
    .Q_N(_4291_),
    .Q(\draw_game_inst.grid[51] ));
 sg13g2_dfrbp_1 _8797_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net53),
    .D(net755),
    .Q_N(_4290_),
    .Q(\draw_game_inst.grid[52] ));
 sg13g2_dfrbp_1 _8798_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net51),
    .D(net681),
    .Q_N(_4289_),
    .Q(\draw_game_inst.grid[53] ));
 sg13g2_dfrbp_1 _8799_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net49),
    .D(net819),
    .Q_N(_4288_),
    .Q(\draw_game_inst.grid[54] ));
 sg13g2_dfrbp_1 _8800_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net47),
    .D(net774),
    .Q_N(_4287_),
    .Q(\draw_game_inst.grid[55] ));
 sg13g2_dfrbp_1 _8801_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net45),
    .D(net718),
    .Q_N(_4286_),
    .Q(\draw_game_inst.grid[56] ));
 sg13g2_dfrbp_1 _8802_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net43),
    .D(net678),
    .Q_N(_4285_),
    .Q(\draw_game_inst.grid[57] ));
 sg13g2_dfrbp_1 _8803_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net41),
    .D(net757),
    .Q_N(_4284_),
    .Q(\draw_game_inst.grid[58] ));
 sg13g2_dfrbp_1 _8804_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net39),
    .D(net732),
    .Q_N(_4283_),
    .Q(\draw_game_inst.grid[59] ));
 sg13g2_dfrbp_1 _8805_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net37),
    .D(net638),
    .Q_N(_4282_),
    .Q(\draw_game_inst.grid[60] ));
 sg13g2_dfrbp_1 _8806_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net35),
    .D(net724),
    .Q_N(_4281_),
    .Q(\draw_game_inst.grid[61] ));
 sg13g2_dfrbp_1 _8807_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net33),
    .D(net741),
    .Q_N(_4280_),
    .Q(\draw_game_inst.grid[62] ));
 sg13g2_dfrbp_1 _8808_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net31),
    .D(net716),
    .Q_N(_4279_),
    .Q(\draw_game_inst.grid[63] ));
 sg13g2_dfrbp_1 _8809_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net29),
    .D(_0256_),
    .Q_N(_0165_),
    .Q(show_welcome_screen));
 sg13g2_dfrbp_1 _8810_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net27),
    .D(_0257_),
    .Q_N(_4278_),
    .Q(btn_select_prev));
 sg13g2_dfrbp_1 _8811_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net26),
    .D(_0258_),
    .Q_N(_4277_),
    .Q(\draw_game_inst.new_tiles[0] ));
 sg13g2_dfrbp_1 _8812_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net25),
    .D(_0259_),
    .Q_N(_0070_),
    .Q(\draw_game_inst.new_tiles[1] ));
 sg13g2_dfrbp_1 _8813_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net415),
    .D(net426),
    .Q_N(_0071_),
    .Q(\draw_game_inst.new_tiles[2] ));
 sg13g2_dfrbp_1 _8814_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net414),
    .D(net438),
    .Q_N(_0072_),
    .Q(\draw_game_inst.new_tiles[3] ));
 sg13g2_dfrbp_1 _8815_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net413),
    .D(net430),
    .Q_N(_0073_),
    .Q(\draw_game_inst.new_tiles[4] ));
 sg13g2_dfrbp_1 _8816_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net412),
    .D(_0263_),
    .Q_N(_0074_),
    .Q(\draw_game_inst.new_tiles[5] ));
 sg13g2_dfrbp_1 _8817_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net411),
    .D(_0264_),
    .Q_N(_0075_),
    .Q(\draw_game_inst.new_tiles[6] ));
 sg13g2_dfrbp_1 _8818_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net410),
    .D(net432),
    .Q_N(_0076_),
    .Q(\draw_game_inst.new_tiles[7] ));
 sg13g2_dfrbp_1 _8819_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net409),
    .D(net419),
    .Q_N(_0077_),
    .Q(\draw_game_inst.new_tiles[8] ));
 sg13g2_dfrbp_1 _8820_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net408),
    .D(net428),
    .Q_N(_0078_),
    .Q(\draw_game_inst.new_tiles[9] ));
 sg13g2_dfrbp_1 _8821_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net407),
    .D(net421),
    .Q_N(_0079_),
    .Q(\draw_game_inst.new_tiles[10] ));
 sg13g2_dfrbp_1 _8822_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net406),
    .D(net423),
    .Q_N(_0080_),
    .Q(\draw_game_inst.new_tiles[11] ));
 sg13g2_dfrbp_1 _8823_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net405),
    .D(net436),
    .Q_N(_0081_),
    .Q(\draw_game_inst.new_tiles[12] ));
 sg13g2_dfrbp_1 _8824_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net404),
    .D(_0271_),
    .Q_N(_0082_),
    .Q(\draw_game_inst.new_tiles[13] ));
 sg13g2_dfrbp_1 _8825_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net403),
    .D(_0272_),
    .Q_N(_0083_),
    .Q(\draw_game_inst.new_tiles[14] ));
 sg13g2_dfrbp_1 _8826_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net402),
    .D(net434),
    .Q_N(_0084_),
    .Q(\draw_game_inst.new_tiles[15] ));
 sg13g2_dfrbp_1 _8827_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net401),
    .D(_0274_),
    .Q_N(_0085_),
    .Q(\new_tiles_counter[0] ));
 sg13g2_dfrbp_1 _8828_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net400),
    .D(net480),
    .Q_N(_0086_),
    .Q(\draw_game_inst.new_tiles_counter[0] ));
 sg13g2_dfrbp_1 _8829_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net399),
    .D(_0276_),
    .Q_N(_4276_),
    .Q(\draw_game_inst.new_tiles_counter[1] ));
 sg13g2_dfrbp_1 _8830_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net398),
    .D(net452),
    .Q_N(_0087_),
    .Q(\draw_game_inst.new_tiles_counter[2] ));
 sg13g2_dfrbp_1 _8831_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net397),
    .D(net579),
    .Q_N(_4275_),
    .Q(\new_tiles_counter[4] ));
 sg13g2_dfrbp_1 _8832_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net396),
    .D(net466),
    .Q_N(_0167_),
    .Q(retro_colors));
 sg13g2_dfrbp_1 _8833_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net394),
    .D(_0280_),
    .Q_N(_4274_),
    .Q(\btn_up_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 _8834_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net393),
    .D(_0281_),
    .Q_N(_0173_),
    .Q(\btn_up_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 _8835_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net392),
    .D(_0282_),
    .Q_N(_4273_),
    .Q(\btn_up_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 _8836_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net391),
    .D(net489),
    .Q_N(_4272_),
    .Q(\btn_up_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 _8837_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net326),
    .D(_0284_),
    .Q_N(_4271_),
    .Q(\btn_up_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 _8838_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net325),
    .D(_0285_),
    .Q_N(_4270_),
    .Q(\btn_up_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 _8839_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net324),
    .D(_0286_),
    .Q_N(_4269_),
    .Q(\btn_up_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 _8840_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net323),
    .D(_0287_),
    .Q_N(_4268_),
    .Q(\btn_up_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 _8841_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net322),
    .D(net599),
    .Q_N(_4267_),
    .Q(\btn_up_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 _8842_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net321),
    .D(_0289_),
    .Q_N(_4266_),
    .Q(\btn_up_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 _8843_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net320),
    .D(_0290_),
    .Q_N(_4265_),
    .Q(\btn_up_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 _8844_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net319),
    .D(net546),
    .Q_N(_4264_),
    .Q(\btn_up_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 _8845_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net318),
    .D(net802),
    .Q_N(_4263_),
    .Q(\btn_up_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 _8846_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net317),
    .D(net564),
    .Q_N(_4262_),
    .Q(\btn_up_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 _8847_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net316),
    .D(_0294_),
    .Q_N(_4261_),
    .Q(\btn_up_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 _8848_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net315),
    .D(_0295_),
    .Q_N(_4260_),
    .Q(\btn_up_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 _8849_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net314),
    .D(_0296_),
    .Q_N(_4259_),
    .Q(\btn_up_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 _8850_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net310),
    .D(_0297_),
    .Q_N(_4258_),
    .Q(\btn_up_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 _8851_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net309),
    .D(net554),
    .Q_N(_4257_),
    .Q(\btn_up_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 _8852_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net308),
    .D(_0299_),
    .Q_N(_4256_),
    .Q(\btn_right_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 _8853_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net307),
    .D(net617),
    .Q_N(_4255_),
    .Q(\btn_up_debounce.debounced ));
 sg13g2_dfrbp_1 _8854_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net305),
    .D(_0301_),
    .Q_N(_4254_),
    .Q(\btn_down_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 _8855_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net304),
    .D(_0302_),
    .Q_N(_0172_),
    .Q(\btn_down_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 _8856_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net303),
    .D(net498),
    .Q_N(_4253_),
    .Q(\btn_down_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 _8857_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net302),
    .D(_0304_),
    .Q_N(_4252_),
    .Q(\btn_down_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 _8858_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net301),
    .D(_0305_),
    .Q_N(_4251_),
    .Q(\btn_down_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 _8859_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net300),
    .D(_0306_),
    .Q_N(_4250_),
    .Q(\btn_down_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 _8860_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net299),
    .D(_0307_),
    .Q_N(_4249_),
    .Q(\btn_down_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 _8861_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net298),
    .D(_0308_),
    .Q_N(_4248_),
    .Q(\btn_down_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 _8862_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net297),
    .D(_0309_),
    .Q_N(_4247_),
    .Q(\btn_down_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 _8863_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net296),
    .D(_0310_),
    .Q_N(_4246_),
    .Q(\btn_down_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 _8864_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net295),
    .D(_0311_),
    .Q_N(_4245_),
    .Q(\btn_down_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 _8865_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net294),
    .D(net549),
    .Q_N(_4244_),
    .Q(\btn_down_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 _8866_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net293),
    .D(_0313_),
    .Q_N(_4243_),
    .Q(\btn_down_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 _8867_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net292),
    .D(net527),
    .Q_N(_4242_),
    .Q(\btn_down_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 _8868_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net291),
    .D(_0315_),
    .Q_N(_4241_),
    .Q(\btn_down_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 _8869_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net290),
    .D(_0316_),
    .Q_N(_4240_),
    .Q(\btn_down_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 _8870_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net289),
    .D(_0317_),
    .Q_N(_4239_),
    .Q(\btn_down_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 _8871_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net288),
    .D(net515),
    .Q_N(_4238_),
    .Q(\btn_down_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 _8872_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net287),
    .D(net486),
    .Q_N(_4237_),
    .Q(\btn_down_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 _8873_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net286),
    .D(net461),
    .Q_N(_4236_),
    .Q(\btn_down_debounce.debounced ));
 sg13g2_dfrbp_1 _8874_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net284),
    .D(_0321_),
    .Q_N(_4235_),
    .Q(\btn_left_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 _8875_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net283),
    .D(_0322_),
    .Q_N(_0171_),
    .Q(\btn_left_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 _8876_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net282),
    .D(_0323_),
    .Q_N(_4234_),
    .Q(\btn_left_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 _8877_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net281),
    .D(net533),
    .Q_N(_4233_),
    .Q(\btn_left_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 _8878_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net280),
    .D(_0325_),
    .Q_N(_4232_),
    .Q(\btn_left_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 _8879_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net279),
    .D(_0326_),
    .Q_N(_4231_),
    .Q(\btn_left_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 _8880_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net278),
    .D(_0327_),
    .Q_N(_4230_),
    .Q(\btn_left_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 _8881_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net277),
    .D(_0328_),
    .Q_N(_4229_),
    .Q(\btn_left_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 _8882_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net276),
    .D(_0329_),
    .Q_N(_4228_),
    .Q(\btn_left_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 _8883_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net274),
    .D(_0330_),
    .Q_N(_4227_),
    .Q(\btn_left_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 _8884_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net273),
    .D(_0331_),
    .Q_N(_4226_),
    .Q(\btn_left_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 _8885_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net272),
    .D(_0332_),
    .Q_N(_4225_),
    .Q(\btn_left_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 _8886_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net271),
    .D(_0333_),
    .Q_N(_4224_),
    .Q(\btn_left_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 _8887_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net270),
    .D(net538),
    .Q_N(_4223_),
    .Q(\btn_left_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 _8888_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net269),
    .D(_0335_),
    .Q_N(_4222_),
    .Q(\btn_left_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 _8889_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net268),
    .D(_0336_),
    .Q_N(_4221_),
    .Q(\btn_left_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 _8890_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net267),
    .D(_0337_),
    .Q_N(_4220_),
    .Q(\btn_left_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 _8891_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net266),
    .D(_0338_),
    .Q_N(_4219_),
    .Q(\btn_left_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 _8892_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net265),
    .D(net590),
    .Q_N(_4218_),
    .Q(\btn_left_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 _8893_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net263),
    .D(_0340_),
    .Q_N(_4217_),
    .Q(\btn_down_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 _8894_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net262),
    .D(net504),
    .Q_N(_4216_),
    .Q(\btn_left_debounce.debounced ));
 sg13g2_dfrbp_1 _8895_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net260),
    .D(_0342_),
    .Q_N(_4215_),
    .Q(\btn_right_debounce.button_sync_0 ));
 sg13g2_dfrbp_1 _8896_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net259),
    .D(_0343_),
    .Q_N(_0170_),
    .Q(\btn_right_debounce.debounce_counter[0] ));
 sg13g2_dfrbp_1 _8897_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net258),
    .D(_0344_),
    .Q_N(_4214_),
    .Q(\btn_right_debounce.debounce_counter[1] ));
 sg13g2_dfrbp_1 _8898_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net257),
    .D(net494),
    .Q_N(_4213_),
    .Q(\btn_right_debounce.debounce_counter[2] ));
 sg13g2_dfrbp_1 _8899_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net256),
    .D(_0346_),
    .Q_N(_4212_),
    .Q(\btn_right_debounce.debounce_counter[3] ));
 sg13g2_dfrbp_1 _8900_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net255),
    .D(_0347_),
    .Q_N(_4211_),
    .Q(\btn_right_debounce.debounce_counter[4] ));
 sg13g2_dfrbp_1 _8901_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net254),
    .D(_0348_),
    .Q_N(_4210_),
    .Q(\btn_right_debounce.debounce_counter[5] ));
 sg13g2_dfrbp_1 _8902_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net253),
    .D(_0349_),
    .Q_N(_4209_),
    .Q(\btn_right_debounce.debounce_counter[6] ));
 sg13g2_dfrbp_1 _8903_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net252),
    .D(_0350_),
    .Q_N(_4208_),
    .Q(\btn_right_debounce.debounce_counter[7] ));
 sg13g2_dfrbp_1 _8904_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net251),
    .D(_0351_),
    .Q_N(_4207_),
    .Q(\btn_right_debounce.debounce_counter[8] ));
 sg13g2_dfrbp_1 _8905_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net250),
    .D(_0352_),
    .Q_N(_4206_),
    .Q(\btn_right_debounce.debounce_counter[9] ));
 sg13g2_dfrbp_1 _8906_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net249),
    .D(net524),
    .Q_N(_4205_),
    .Q(\btn_right_debounce.debounce_counter[10] ));
 sg13g2_dfrbp_1 _8907_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net248),
    .D(net842),
    .Q_N(_4204_),
    .Q(\btn_right_debounce.debounce_counter[11] ));
 sg13g2_dfrbp_1 _8908_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net247),
    .D(net576),
    .Q_N(_4203_),
    .Q(\btn_right_debounce.debounce_counter[12] ));
 sg13g2_dfrbp_1 _8909_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net246),
    .D(_0356_),
    .Q_N(_4202_),
    .Q(\btn_right_debounce.debounce_counter[13] ));
 sg13g2_dfrbp_1 _8910_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net245),
    .D(_0357_),
    .Q_N(_4201_),
    .Q(\btn_right_debounce.debounce_counter[14] ));
 sg13g2_dfrbp_1 _8911_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net244),
    .D(net585),
    .Q_N(_4200_),
    .Q(\btn_right_debounce.debounce_counter[15] ));
 sg13g2_dfrbp_1 _8912_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net243),
    .D(net530),
    .Q_N(_4199_),
    .Q(\btn_right_debounce.debounce_counter[16] ));
 sg13g2_dfrbp_1 _8913_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net242),
    .D(net501),
    .Q_N(_4198_),
    .Q(\btn_right_debounce.debounce_counter[17] ));
 sg13g2_dfrbp_1 _8914_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net241),
    .D(_0361_),
    .Q_N(_4197_),
    .Q(\btn_left_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 _8915_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net240),
    .D(net646),
    .Q_N(_4196_),
    .Q(\btn_right_debounce.debounced ));
 sg13g2_dfrbp_1 _8916_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net215),
    .D(_0363_),
    .Q_N(_4356_),
    .Q(\game_logic_inst.prev_any_button_pressed ));
 sg13g2_dfrbp_1 _8917_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net264),
    .D(net417),
    .Q_N(_4357_),
    .Q(\gamepad_pmod.driver.pmod_clk_prev ));
 sg13g2_dfrbp_1 _8918_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net238),
    .D(net416),
    .Q_N(_4195_),
    .Q(\gamepad_pmod.driver.pmod_latch_prev ));
 sg13g2_dfrbp_1 _8919_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net237),
    .D(net513),
    .Q_N(_4194_),
    .Q(\gamepad_pmod.driver.shift_reg[0] ));
 sg13g2_dfrbp_1 _8920_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net235),
    .D(net587),
    .Q_N(_4193_),
    .Q(\gamepad_pmod.driver.shift_reg[1] ));
 sg13g2_dfrbp_1 _8921_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net233),
    .D(net470),
    .Q_N(_4192_),
    .Q(\gamepad_pmod.driver.shift_reg[2] ));
 sg13g2_dfrbp_1 _8922_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net231),
    .D(net606),
    .Q_N(_4191_),
    .Q(\gamepad_pmod.driver.shift_reg[3] ));
 sg13g2_dfrbp_1 _8923_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net229),
    .D(_0368_),
    .Q_N(_4190_),
    .Q(\gamepad_pmod.driver.shift_reg[4] ));
 sg13g2_dfrbp_1 _8924_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net227),
    .D(net615),
    .Q_N(_4189_),
    .Q(\gamepad_pmod.driver.shift_reg[5] ));
 sg13g2_dfrbp_1 _8925_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net225),
    .D(net608),
    .Q_N(_4188_),
    .Q(\gamepad_pmod.driver.shift_reg[6] ));
 sg13g2_dfrbp_1 _8926_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net223),
    .D(net596),
    .Q_N(_4187_),
    .Q(\gamepad_pmod.driver.shift_reg[7] ));
 sg13g2_dfrbp_1 _8927_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net221),
    .D(net592),
    .Q_N(_4186_),
    .Q(\gamepad_pmod.driver.shift_reg[8] ));
 sg13g2_dfrbp_1 _8928_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net219),
    .D(_0373_),
    .Q_N(_4185_),
    .Q(\gamepad_pmod.driver.shift_reg[9] ));
 sg13g2_dfrbp_1 _8929_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net217),
    .D(net468),
    .Q_N(_4184_),
    .Q(\gamepad_pmod.driver.shift_reg[10] ));
 sg13g2_dfrbp_1 _8930_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net213),
    .D(net541),
    .Q_N(_4183_),
    .Q(\gamepad_pmod.driver.shift_reg[11] ));
 sg13g2_dfrbp_1 _8931_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net211),
    .D(_0376_),
    .Q_N(_4182_),
    .Q(\gamepad_pmod.driver.pmod_data_sync[0] ));
 sg13g2_dfrbp_1 _8932_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net210),
    .D(_0377_),
    .Q_N(_4181_),
    .Q(\gamepad_pmod.driver.pmod_data_sync[1] ));
 sg13g2_dfrbp_1 _8933_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net209),
    .D(_0378_),
    .Q_N(_4180_),
    .Q(\gamepad_pmod.driver.pmod_clk_sync[0] ));
 sg13g2_dfrbp_1 _8934_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net208),
    .D(_0379_),
    .Q_N(_4179_),
    .Q(\gamepad_pmod.driver.pmod_clk_sync[1] ));
 sg13g2_dfrbp_1 _8935_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net207),
    .D(_0380_),
    .Q_N(_4178_),
    .Q(\game_logic_inst.lfsr_value[0] ));
 sg13g2_dfrbp_1 _8936_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net206),
    .D(_0381_),
    .Q_N(_4177_),
    .Q(\game_logic_inst.lfsr_value[1] ));
 sg13g2_dfrbp_1 _8937_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net205),
    .D(_0382_),
    .Q_N(_4176_),
    .Q(\game_logic_inst.lfsr_value[2] ));
 sg13g2_dfrbp_1 _8938_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net204),
    .D(_0383_),
    .Q_N(_4175_),
    .Q(\game_logic_inst.lfsr_value[3] ));
 sg13g2_dfrbp_1 _8939_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net203),
    .D(_0384_),
    .Q_N(_4174_),
    .Q(\game_logic_inst.lfsr_value[4] ));
 sg13g2_dfrbp_1 _8940_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net202),
    .D(_0385_),
    .Q_N(_4173_),
    .Q(\game_logic_inst.lfsr_value[5] ));
 sg13g2_dfrbp_1 _8941_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net201),
    .D(_0386_),
    .Q_N(_4172_),
    .Q(\game_logic_inst.lfsr_value[6] ));
 sg13g2_dfrbp_1 _8942_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net200),
    .D(_0387_),
    .Q_N(_4171_),
    .Q(\game_logic_inst.lfsr_value[7] ));
 sg13g2_dfrbp_1 _8943_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net199),
    .D(_0388_),
    .Q_N(_4170_),
    .Q(\game_logic_inst.lfsr_value[8] ));
 sg13g2_dfrbp_1 _8944_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net198),
    .D(_0389_),
    .Q_N(_4169_),
    .Q(\game_logic_inst.lfsr_value[9] ));
 sg13g2_dfrbp_1 _8945_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net197),
    .D(_0390_),
    .Q_N(_4168_),
    .Q(\game_logic_inst.lfsr_value[10] ));
 sg13g2_dfrbp_1 _8946_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net196),
    .D(_0391_),
    .Q_N(_4167_),
    .Q(\game_logic_inst.lfsr_value[11] ));
 sg13g2_dfrbp_1 _8947_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net195),
    .D(_0392_),
    .Q_N(_4166_),
    .Q(\game_logic_inst.lfsr_value[12] ));
 sg13g2_dfrbp_1 _8948_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net194),
    .D(_0393_),
    .Q_N(_4165_),
    .Q(\game_logic_inst.lfsr_value[13] ));
 sg13g2_dfrbp_1 _8949_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net193),
    .D(_0394_),
    .Q_N(_4164_),
    .Q(\game_logic_inst.lfsr_value[14] ));
 sg13g2_dfrbp_1 _8950_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net192),
    .D(_0395_),
    .Q_N(_4163_),
    .Q(\game_logic_inst.lfsr_value[15] ));
 sg13g2_dfrbp_1 _8951_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net191),
    .D(_0396_),
    .Q_N(_4162_),
    .Q(\lfsr_inst.lfsr[16] ));
 sg13g2_dfrbp_1 _8952_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net190),
    .D(_0397_),
    .Q_N(_4161_),
    .Q(\lfsr_inst.lfsr[17] ));
 sg13g2_dfrbp_1 _8953_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net189),
    .D(_0398_),
    .Q_N(_4160_),
    .Q(\lfsr_inst.lfsr[18] ));
 sg13g2_dfrbp_1 _8954_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net188),
    .D(_0399_),
    .Q_N(_4159_),
    .Q(\lfsr_inst.lfsr[19] ));
 sg13g2_dfrbp_1 _8955_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net187),
    .D(_0400_),
    .Q_N(_4158_),
    .Q(\lfsr_inst.lfsr[20] ));
 sg13g2_dfrbp_1 _8956_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net186),
    .D(_0401_),
    .Q_N(_4157_),
    .Q(\lfsr_inst.lfsr[21] ));
 sg13g2_dfrbp_1 _8957_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net185),
    .D(_0402_),
    .Q_N(_4156_),
    .Q(\lfsr_inst.lfsr[22] ));
 sg13g2_dfrbp_1 _8958_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net184),
    .D(_0403_),
    .Q_N(_4155_),
    .Q(\lfsr_inst.lfsr[23] ));
 sg13g2_dfrbp_1 _8959_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net183),
    .D(_0404_),
    .Q_N(_4154_),
    .Q(\lfsr_inst.lfsr[24] ));
 sg13g2_dfrbp_1 _8960_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net182),
    .D(_0405_),
    .Q_N(_4153_),
    .Q(\lfsr_inst.lfsr[25] ));
 sg13g2_dfrbp_1 _8961_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net181),
    .D(_0406_),
    .Q_N(_4152_),
    .Q(\lfsr_inst.lfsr[26] ));
 sg13g2_dfrbp_1 _8962_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net180),
    .D(_0407_),
    .Q_N(_4151_),
    .Q(\lfsr_inst.lfsr[27] ));
 sg13g2_dfrbp_1 _8963_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net179),
    .D(_0408_),
    .Q_N(_4150_),
    .Q(\lfsr_inst.lfsr[28] ));
 sg13g2_dfrbp_1 _8964_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net178),
    .D(_0409_),
    .Q_N(_4149_),
    .Q(\lfsr_inst.lfsr[29] ));
 sg13g2_dfrbp_1 _8965_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net177),
    .D(_0410_),
    .Q_N(_4148_),
    .Q(\lfsr_inst.lfsr[30] ));
 sg13g2_dfrbp_1 _8966_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net275),
    .D(_0411_),
    .Q_N(_4358_),
    .Q(\lfsr_inst.lfsr[31] ));
 sg13g2_dfrbp_1 _8967_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net176),
    .D(net921),
    .Q_N(_4147_),
    .Q(hsync));
 sg13g2_dfrbp_1 _8968_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net175),
    .D(_0412_),
    .Q_N(_0169_),
    .Q(\draw_game_inst.board_y[0] ));
 sg13g2_dfrbp_1 _8969_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net156),
    .D(_0413_),
    .Q_N(_0093_),
    .Q(\draw_game_inst.board_y[1] ));
 sg13g2_dfrbp_1 _8970_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net152),
    .D(_0414_),
    .Q_N(_0092_),
    .Q(\draw_game_inst.board_y[2] ));
 sg13g2_dfrbp_1 _8971_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net148),
    .D(_0415_),
    .Q_N(_0091_),
    .Q(\draw_game_inst.board_y[3] ));
 sg13g2_dfrbp_1 _8972_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net144),
    .D(_0416_),
    .Q_N(_0090_),
    .Q(\draw_game_inst.board_y[4] ));
 sg13g2_dfrbp_1 _8973_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net140),
    .D(net979),
    .Q_N(_4146_),
    .Q(\draw_game_inst.board_y[5] ));
 sg13g2_dfrbp_1 _8974_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net136),
    .D(_0418_),
    .Q_N(_0089_),
    .Q(\draw_game_inst.board_y[6] ));
 sg13g2_dfrbp_1 _8975_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net132),
    .D(net772),
    .Q_N(_0088_),
    .Q(\draw_game_inst.y[7] ));
 sg13g2_dfrbp_1 _8976_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net128),
    .D(_0420_),
    .Q_N(_4145_),
    .Q(\draw_game_inst.y[8] ));
 sg13g2_dfrbp_1 _8977_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net311),
    .D(net860),
    .Q_N(_4359_),
    .Q(\draw_game_inst.y[9] ));
 sg13g2_dfrbp_1 _8978_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net124),
    .D(_0068_),
    .Q_N(_4144_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_dfrbp_1 _8979_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net120),
    .D(_0422_),
    .Q_N(_4143_),
    .Q(\gamepad_pmod.driver.pmod_latch_sync[0] ));
 sg13g2_dfrbp_1 _8980_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net118),
    .D(_0423_),
    .Q_N(_4142_),
    .Q(\gamepad_pmod.driver.pmod_latch_sync[1] ));
 sg13g2_dfrbp_1 _8981_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net116),
    .D(net511),
    .Q_N(_4141_),
    .Q(\gamepad_pmod.decoder.data_reg[0] ));
 sg13g2_dfrbp_1 _8982_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net112),
    .D(net491),
    .Q_N(_4140_),
    .Q(\gamepad_pmod.decoder.data_reg[1] ));
 sg13g2_dfrbp_1 _8983_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net108),
    .D(net507),
    .Q_N(_4139_),
    .Q(\gamepad_pmod.decoder.data_reg[2] ));
 sg13g2_dfrbp_1 _8984_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net104),
    .D(net519),
    .Q_N(_4138_),
    .Q(\gamepad_pmod.decoder.data_reg[3] ));
 sg13g2_dfrbp_1 _8985_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net100),
    .D(net561),
    .Q_N(_4137_),
    .Q(\gamepad_pmod.decoder.data_reg[4] ));
 sg13g2_dfrbp_1 _8986_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net96),
    .D(net603),
    .Q_N(_4136_),
    .Q(\gamepad_pmod.decoder.data_reg[5] ));
 sg13g2_dfrbp_1 _8987_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net92),
    .D(net558),
    .Q_N(_4135_),
    .Q(\gamepad_pmod.decoder.data_reg[6] ));
 sg13g2_dfrbp_1 _8988_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net88),
    .D(net551),
    .Q_N(_4134_),
    .Q(\gamepad_pmod.decoder.data_reg[7] ));
 sg13g2_dfrbp_1 _8989_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net84),
    .D(_0432_),
    .Q_N(_4133_),
    .Q(\gamepad_pmod.decoder.data_reg[8] ));
 sg13g2_dfrbp_1 _8990_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net80),
    .D(_0433_),
    .Q_N(_4132_),
    .Q(\gamepad_pmod.decoder.data_reg[9] ));
 sg13g2_dfrbp_1 _8991_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net76),
    .D(net535),
    .Q_N(_4131_),
    .Q(\gamepad_pmod.decoder.data_reg[10] ));
 sg13g2_dfrbp_1 _8992_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net72),
    .D(net509),
    .Q_N(_4130_),
    .Q(\gamepad_pmod.decoder.data_reg[11] ));
 sg13g2_dfrbp_1 _8993_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net68),
    .D(net838),
    .Q_N(_4129_),
    .Q(\welcome_screen_grid[0] ));
 sg13g2_dfrbp_1 _8994_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net64),
    .D(_0437_),
    .Q_N(_4128_),
    .Q(\welcome_screen_grid[4] ));
 sg13g2_dfrbp_1 _8995_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net60),
    .D(_0438_),
    .Q_N(_4127_),
    .Q(\welcome_screen_grid[11] ));
 sg13g2_dfrbp_1 _8996_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net56),
    .D(_0439_),
    .Q_N(_4126_),
    .Q(\welcome_screen_grid[12] ));
 sg13g2_dfrbp_1 _8997_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net52),
    .D(_0440_),
    .Q_N(_4125_),
    .Q(\welcome_screen_grid[16] ));
 sg13g2_dfrbp_1 _8998_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net48),
    .D(_0441_),
    .Q_N(_4124_),
    .Q(\welcome_screen_grid[20] ));
 sg13g2_dfrbp_1 _8999_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net44),
    .D(_0442_),
    .Q_N(_4123_),
    .Q(\welcome_screen_grid[24] ));
 sg13g2_dfrbp_1 _9000_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net40),
    .D(_0443_),
    .Q_N(_4122_),
    .Q(\welcome_screen_grid[28] ));
 sg13g2_dfrbp_1 _9001_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net36),
    .D(net743),
    .Q_N(_4121_),
    .Q(\welcome_screen_grid[32] ));
 sg13g2_dfrbp_1 _9002_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net32),
    .D(_0445_),
    .Q_N(_4120_),
    .Q(\welcome_screen_grid[36] ));
 sg13g2_dfrbp_1 _9003_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net28),
    .D(_0446_),
    .Q_N(_4119_),
    .Q(\welcome_screen_grid[40] ));
 sg13g2_dfrbp_1 _9004_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net306),
    .D(_0447_),
    .Q_N(_4118_),
    .Q(\welcome_screen_grid[44] ));
 sg13g2_dfrbp_1 _9005_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net261),
    .D(_0448_),
    .Q_N(_4117_),
    .Q(\welcome_screen_grid[48] ));
 sg13g2_dfrbp_1 _9006_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net236),
    .D(_0449_),
    .Q_N(_4116_),
    .Q(\welcome_screen_grid[52] ));
 sg13g2_dfrbp_1 _9007_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net232),
    .D(_0450_),
    .Q_N(_4115_),
    .Q(\welcome_screen_grid[56] ));
 sg13g2_dfrbp_1 _9008_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net228),
    .D(_0451_),
    .Q_N(_4114_),
    .Q(\welcome_screen_grid[60] ));
 sg13g2_dfrbp_1 _9009_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net224),
    .D(_0452_),
    .Q_N(_4113_),
    .Q(\welcome_screen_inst.welcome_counter[0] ));
 sg13g2_dfrbp_1 _9010_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net220),
    .D(net628),
    .Q_N(_4112_),
    .Q(\welcome_screen_inst.welcome_counter[1] ));
 sg13g2_dfrbp_1 _9011_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net216),
    .D(_0454_),
    .Q_N(_4111_),
    .Q(\welcome_screen_inst.welcome_counter[2] ));
 sg13g2_dfrbp_1 _9012_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net174),
    .D(_0455_),
    .Q_N(_4110_),
    .Q(\welcome_screen_inst.welcome_counter[3] ));
 sg13g2_dfrbp_1 _9013_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net312),
    .D(net738),
    .Q_N(_4360_),
    .Q(\welcome_screen_inst.welcome_counter[4] ));
 sg13g2_dfrbp_1 _9014_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net313),
    .D(net556),
    .Q_N(_4361_),
    .Q(\game_logic_inst.current_direction[1] ));
 sg13g2_dfrbp_1 _9015_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net327),
    .D(net864),
    .Q_N(_4362_),
    .Q(\game_logic_inst.current_direction[2] ));
 sg13g2_dfrbp_1 _9016_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net150),
    .D(_0002_),
    .Q_N(_4109_),
    .Q(\game_logic_inst.current_direction[3] ));
 sg13g2_dfrbp_1 _9017_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net142),
    .D(net850),
    .Q_N(_4108_),
    .Q(\game_logic_inst.debug_move_reg ));
 sg13g2_dfrbp_1 _9018_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net134),
    .D(_0458_),
    .Q_N(_4107_),
    .Q(\game_logic_inst.valid_move ));
 sg13g2_dfrbp_1 _9019_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net126),
    .D(_0459_),
    .Q_N(_0097_),
    .Q(\game_logic_inst.calculate_move ));
 sg13g2_dfrbp_1 _9020_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net114),
    .D(_0460_),
    .Q_N(_0168_),
    .Q(\game_logic_inst.lfsr_shift[0] ));
 sg13g2_dfrbp_1 _9021_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net110),
    .D(_0461_),
    .Q_N(_4106_),
    .Q(\game_logic_inst.lfsr_shift[1] ));
 sg13g2_dfrbp_1 _9022_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net106),
    .D(_0462_),
    .Q_N(_0166_),
    .Q(\game_logic_inst.game_started ));
 sg13g2_dfrbp_1 _9023_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net102),
    .D(_0463_),
    .Q_N(_4105_),
    .Q(\game_logic_inst.add_new_tiles[0] ));
 sg13g2_dfrbp_1 _9024_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net94),
    .D(net569),
    .Q_N(_4104_),
    .Q(\game_logic_inst.add_new_tiles[1] ));
 sg13g2_dfrbp_1 _9025_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net86),
    .D(_0465_),
    .Q_N(_4103_),
    .Q(\game_logic_inst.added_tile_index[0] ));
 sg13g2_dfrbp_1 _9026_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net82),
    .D(_0466_),
    .Q_N(_4102_),
    .Q(\game_logic_inst.added_tile_index[1] ));
 sg13g2_dfrbp_1 _9027_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net78),
    .D(_0467_),
    .Q_N(_4101_),
    .Q(\game_logic_inst.added_tile_index[2] ));
 sg13g2_dfrbp_1 _9028_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net74),
    .D(_0468_),
    .Q_N(_4100_),
    .Q(\game_logic_inst.added_tile_index[3] ));
 sg13g2_dfrbp_1 _9029_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net328),
    .D(_0469_),
    .Q_N(_4363_),
    .Q(\debug_controller_inst.data_out_en ));
 sg13g2_dfrbp_1 _9030_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net329),
    .D(_0003_),
    .Q_N(_0099_),
    .Q(\debug_controller_inst.grid_in[0] ));
 sg13g2_dfrbp_1 _9031_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net330),
    .D(_0014_),
    .Q_N(_0100_),
    .Q(\debug_controller_inst.grid_in[1] ));
 sg13g2_dfrbp_1 _9032_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net331),
    .D(_0025_),
    .Q_N(_0101_),
    .Q(\debug_controller_inst.grid_in[2] ));
 sg13g2_dfrbp_1 _9033_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net332),
    .D(net907),
    .Q_N(_0102_),
    .Q(\debug_controller_inst.grid_in[3] ));
 sg13g2_dfrbp_1 _9034_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net333),
    .D(_0047_),
    .Q_N(_0103_),
    .Q(\debug_controller_inst.grid_in[4] ));
 sg13g2_dfrbp_1 _9035_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net334),
    .D(_0058_),
    .Q_N(_0105_),
    .Q(\debug_controller_inst.grid_in[5] ));
 sg13g2_dfrbp_1 _9036_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net335),
    .D(_0063_),
    .Q_N(_0107_),
    .Q(\debug_controller_inst.grid_in[6] ));
 sg13g2_dfrbp_1 _9037_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net336),
    .D(_0064_),
    .Q_N(_0109_),
    .Q(\debug_controller_inst.grid_in[7] ));
 sg13g2_dfrbp_1 _9038_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net337),
    .D(_0065_),
    .Q_N(_0111_),
    .Q(\debug_controller_inst.grid_in[8] ));
 sg13g2_dfrbp_1 _9039_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net338),
    .D(_0066_),
    .Q_N(_0113_),
    .Q(\debug_controller_inst.grid_in[9] ));
 sg13g2_dfrbp_1 _9040_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net339),
    .D(_0004_),
    .Q_N(_0115_),
    .Q(\debug_controller_inst.grid_in[10] ));
 sg13g2_dfrbp_1 _9041_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net340),
    .D(net899),
    .Q_N(_0117_),
    .Q(\debug_controller_inst.grid_in[11] ));
 sg13g2_dfrbp_1 _9042_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net341),
    .D(_0006_),
    .Q_N(_0119_),
    .Q(\debug_controller_inst.grid_in[12] ));
 sg13g2_dfrbp_1 _9043_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net342),
    .D(_0007_),
    .Q_N(_0121_),
    .Q(\debug_controller_inst.grid_in[13] ));
 sg13g2_dfrbp_1 _9044_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net343),
    .D(_0008_),
    .Q_N(_0123_),
    .Q(\debug_controller_inst.grid_in[14] ));
 sg13g2_dfrbp_1 _9045_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net344),
    .D(_0009_),
    .Q_N(_0125_),
    .Q(\debug_controller_inst.grid_in[15] ));
 sg13g2_dfrbp_1 _9046_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net345),
    .D(_0010_),
    .Q_N(_0104_),
    .Q(\debug_controller_inst.grid_in[16] ));
 sg13g2_dfrbp_1 _9047_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net346),
    .D(_0011_),
    .Q_N(_0106_),
    .Q(\debug_controller_inst.grid_in[17] ));
 sg13g2_dfrbp_1 _9048_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net347),
    .D(_0012_),
    .Q_N(_0108_),
    .Q(\debug_controller_inst.grid_in[18] ));
 sg13g2_dfrbp_1 _9049_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net348),
    .D(_0013_),
    .Q_N(_0110_),
    .Q(\debug_controller_inst.grid_in[19] ));
 sg13g2_dfrbp_1 _9050_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net349),
    .D(_0015_),
    .Q_N(_0127_),
    .Q(\debug_controller_inst.grid_in[20] ));
 sg13g2_dfrbp_1 _9051_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net350),
    .D(_0016_),
    .Q_N(_0128_),
    .Q(\debug_controller_inst.grid_in[21] ));
 sg13g2_dfrbp_1 _9052_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net351),
    .D(net904),
    .Q_N(_0129_),
    .Q(\debug_controller_inst.grid_in[22] ));
 sg13g2_dfrbp_1 _9053_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net352),
    .D(net975),
    .Q_N(_0130_),
    .Q(\debug_controller_inst.grid_in[23] ));
 sg13g2_dfrbp_1 _9054_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net353),
    .D(_0019_),
    .Q_N(_0131_),
    .Q(\debug_controller_inst.grid_in[24] ));
 sg13g2_dfrbp_1 _9055_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net354),
    .D(_0020_),
    .Q_N(_0133_),
    .Q(\debug_controller_inst.grid_in[25] ));
 sg13g2_dfrbp_1 _9056_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net355),
    .D(_0021_),
    .Q_N(_0135_),
    .Q(\debug_controller_inst.grid_in[26] ));
 sg13g2_dfrbp_1 _9057_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net356),
    .D(net964),
    .Q_N(_0137_),
    .Q(\debug_controller_inst.grid_in[27] ));
 sg13g2_dfrbp_1 _9058_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net357),
    .D(_0023_),
    .Q_N(_0139_),
    .Q(\debug_controller_inst.grid_in[28] ));
 sg13g2_dfrbp_1 _9059_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net358),
    .D(_0024_),
    .Q_N(_0141_),
    .Q(\debug_controller_inst.grid_in[29] ));
 sg13g2_dfrbp_1 _9060_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net359),
    .D(_0026_),
    .Q_N(_0143_),
    .Q(\debug_controller_inst.grid_in[30] ));
 sg13g2_dfrbp_1 _9061_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net360),
    .D(_0027_),
    .Q_N(_0145_),
    .Q(\debug_controller_inst.grid_in[31] ));
 sg13g2_dfrbp_1 _9062_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net361),
    .D(net953),
    .Q_N(_0112_),
    .Q(\debug_controller_inst.grid_in[32] ));
 sg13g2_dfrbp_1 _9063_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net362),
    .D(_0029_),
    .Q_N(_0114_),
    .Q(\debug_controller_inst.grid_in[33] ));
 sg13g2_dfrbp_1 _9064_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net363),
    .D(_0030_),
    .Q_N(_0116_),
    .Q(\debug_controller_inst.grid_in[34] ));
 sg13g2_dfrbp_1 _9065_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net364),
    .D(net996),
    .Q_N(_0118_),
    .Q(\debug_controller_inst.grid_in[35] ));
 sg13g2_dfrbp_1 _9066_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net365),
    .D(_0032_),
    .Q_N(_0132_),
    .Q(\debug_controller_inst.grid_in[36] ));
 sg13g2_dfrbp_1 _9067_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net366),
    .D(_0033_),
    .Q_N(_0134_),
    .Q(\debug_controller_inst.grid_in[37] ));
 sg13g2_dfrbp_1 _9068_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net367),
    .D(_0034_),
    .Q_N(_0136_),
    .Q(\debug_controller_inst.grid_in[38] ));
 sg13g2_dfrbp_1 _9069_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net368),
    .D(_0035_),
    .Q_N(_0138_),
    .Q(\debug_controller_inst.grid_in[39] ));
 sg13g2_dfrbp_1 _9070_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net369),
    .D(_0037_),
    .Q_N(_0147_),
    .Q(\debug_controller_inst.grid_in[40] ));
 sg13g2_dfrbp_1 _9071_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net370),
    .D(_0038_),
    .Q_N(_0148_),
    .Q(\debug_controller_inst.grid_in[41] ));
 sg13g2_dfrbp_1 _9072_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net371),
    .D(_0039_),
    .Q_N(_0149_),
    .Q(\debug_controller_inst.grid_in[42] ));
 sg13g2_dfrbp_1 _9073_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net372),
    .D(net909),
    .Q_N(_0150_),
    .Q(\debug_controller_inst.grid_in[43] ));
 sg13g2_dfrbp_1 _9074_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net373),
    .D(_0041_),
    .Q_N(_0151_),
    .Q(\debug_controller_inst.grid_in[44] ));
 sg13g2_dfrbp_1 _9075_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net374),
    .D(_0042_),
    .Q_N(_0153_),
    .Q(\debug_controller_inst.grid_in[45] ));
 sg13g2_dfrbp_1 _9076_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net375),
    .D(_0043_),
    .Q_N(_0155_),
    .Q(\debug_controller_inst.grid_in[46] ));
 sg13g2_dfrbp_1 _9077_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net376),
    .D(_0044_),
    .Q_N(_0157_),
    .Q(\debug_controller_inst.grid_in[47] ));
 sg13g2_dfrbp_1 _9078_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net377),
    .D(net1003),
    .Q_N(_0120_),
    .Q(\debug_controller_inst.grid_in[48] ));
 sg13g2_dfrbp_1 _9079_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net378),
    .D(_0046_),
    .Q_N(_0122_),
    .Q(\debug_controller_inst.grid_in[49] ));
 sg13g2_dfrbp_1 _9080_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net379),
    .D(_0048_),
    .Q_N(_0124_),
    .Q(\debug_controller_inst.grid_in[50] ));
 sg13g2_dfrbp_1 _9081_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net380),
    .D(_0049_),
    .Q_N(_0126_),
    .Q(\debug_controller_inst.grid_in[51] ));
 sg13g2_dfrbp_1 _9082_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net381),
    .D(_0050_),
    .Q_N(_0140_),
    .Q(\debug_controller_inst.grid_in[52] ));
 sg13g2_dfrbp_1 _9083_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net382),
    .D(_0051_),
    .Q_N(_0142_),
    .Q(\debug_controller_inst.grid_in[53] ));
 sg13g2_dfrbp_1 _9084_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net383),
    .D(net981),
    .Q_N(_0144_),
    .Q(\debug_controller_inst.grid_in[54] ));
 sg13g2_dfrbp_1 _9085_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net384),
    .D(net951),
    .Q_N(_0146_),
    .Q(\debug_controller_inst.grid_in[55] ));
 sg13g2_dfrbp_1 _9086_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net385),
    .D(_0054_),
    .Q_N(_0152_),
    .Q(\debug_controller_inst.grid_in[56] ));
 sg13g2_dfrbp_1 _9087_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net386),
    .D(_0055_),
    .Q_N(_0154_),
    .Q(\debug_controller_inst.grid_in[57] ));
 sg13g2_dfrbp_1 _9088_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net387),
    .D(_0056_),
    .Q_N(_0156_),
    .Q(\debug_controller_inst.grid_in[58] ));
 sg13g2_dfrbp_1 _9089_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net388),
    .D(_0057_),
    .Q_N(_0158_),
    .Q(\debug_controller_inst.grid_in[59] ));
 sg13g2_dfrbp_1 _9090_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net389),
    .D(_0059_),
    .Q_N(_0159_),
    .Q(\debug_controller_inst.grid_in[60] ));
 sg13g2_dfrbp_1 _9091_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net390),
    .D(_0060_),
    .Q_N(_0160_),
    .Q(\debug_controller_inst.grid_in[61] ));
 sg13g2_dfrbp_1 _9092_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net46),
    .D(_0061_),
    .Q_N(_0161_),
    .Q(\debug_controller_inst.grid_in[62] ));
 sg13g2_dfrbp_1 _9093_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net70),
    .D(net971),
    .Q_N(_0162_),
    .Q(\debug_controller_inst.grid_in[63] ));
 sg13g2_dfrbp_1 _9094_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net66),
    .D(net857),
    .Q_N(_0069_),
    .Q(\game_logic_inst.should_transpose ));
 sg13g2_dfrbp_1 _9095_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net58),
    .D(_0471_),
    .Q_N(_0098_),
    .Q(\game_logic_inst.current_row_index[0] ));
 sg13g2_dfrbp_1 _9096_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net50),
    .D(_0472_),
    .Q_N(_4099_),
    .Q(\game_logic_inst.current_row_index[1] ));
 sg13g2_dfrbp_1 _9097_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net42),
    .D(_0473_),
    .Q_N(_4098_),
    .Q(uio_out[4]));
 sg13g2_dfrbp_1 _9098_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net34),
    .D(_0474_),
    .Q_N(_4097_),
    .Q(uio_out[5]));
 sg13g2_dfrbp_1 _9099_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net395),
    .D(_0475_),
    .Q_N(_4096_),
    .Q(uio_out[6]));
 sg13g2_dfrbp_1 _9100_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net239),
    .D(_0476_),
    .Q_N(_4095_),
    .Q(uio_out[7]));
 sg13g2_dfrbp_1 _9101_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net230),
    .D(_0477_),
    .Q_N(_4094_),
    .Q(debug_btn_up));
 sg13g2_dfrbp_1 _9102_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net226),
    .D(_0478_),
    .Q_N(_4093_),
    .Q(debug_btn_down));
 sg13g2_dfrbp_1 _9103_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net222),
    .D(_0479_),
    .Q_N(_4092_),
    .Q(debug_btn_left));
 sg13g2_dfrbp_1 _9104_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net218),
    .D(_0480_),
    .Q_N(_4091_),
    .Q(debug_btn_right));
 sg13g2_dfrbp_1 _9105_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net212),
    .D(_0481_),
    .Q_N(_4090_),
    .Q(\debug_controller_inst.grid_out_valid ));
 sg13g2_dfrbp_1 _9106_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net154),
    .D(_0482_),
    .Q_N(_4089_),
    .Q(\debug_controller_inst.grid_out_data[0] ));
 sg13g2_dfrbp_1 _9107_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net138),
    .D(_0483_),
    .Q_N(_4088_),
    .Q(\debug_controller_inst.grid_out_data[1] ));
 sg13g2_dfrbp_1 _9108_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net122),
    .D(_0484_),
    .Q_N(_4087_),
    .Q(\debug_controller_inst.grid_out_data[2] ));
 sg13g2_dfrbp_1 _9109_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net90),
    .D(_0485_),
    .Q_N(_4086_),
    .Q(\debug_controller_inst.grid_out_data[3] ));
 sg13g2_dfrbp_1 _9110_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net54),
    .D(net726),
    .Q_N(_4085_),
    .Q(\debug_controller_inst.grid_out_addr[0] ));
 sg13g2_dfrbp_1 _9111_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net38),
    .D(net691),
    .Q_N(_4084_),
    .Q(\debug_controller_inst.grid_out_addr[1] ));
 sg13g2_dfrbp_1 _9112_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net285),
    .D(net817),
    .Q_N(_4083_),
    .Q(\debug_controller_inst.grid_out_addr[2] ));
 sg13g2_dfrbp_1 _9113_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net146),
    .D(_0489_),
    .Q_N(_4082_),
    .Q(\debug_controller_inst.grid_out_addr[3] ));
 sg13g2_dfrbp_1 _9114_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net98),
    .D(_0490_),
    .Q_N(_4081_),
    .Q(\btn_up_debounce.button_sync_1 ));
 sg13g2_dfrbp_1 _9115_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net62),
    .D(_0491_),
    .Q_N(_0163_),
    .Q(\debug_controller_inst.grid_addr[0] ));
 sg13g2_dfrbp_1 _9116_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net30),
    .D(_0492_),
    .Q_N(_4080_),
    .Q(\debug_controller_inst.grid_addr[1] ));
 sg13g2_dfrbp_1 _9117_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net130),
    .D(_0493_),
    .Q_N(_0164_),
    .Q(\debug_controller_inst.grid_addr[2] ));
 sg13g2_dfrbp_1 _9118_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net234),
    .D(net956),
    .Q_N(_4079_),
    .Q(\debug_controller_inst.grid_addr[3] ));
 sg13g2_tiehi _8811__26 (.L_HI(net26));
 sg13g2_tiehi _8810__27 (.L_HI(net27));
 sg13g2_tiehi _9003__28 (.L_HI(net28));
 sg13g2_tiehi _8809__29 (.L_HI(net29));
 sg13g2_tiehi _9116__30 (.L_HI(net30));
 sg13g2_tiehi _8808__31 (.L_HI(net31));
 sg13g2_tiehi _9002__32 (.L_HI(net32));
 sg13g2_tiehi _8807__33 (.L_HI(net33));
 sg13g2_tiehi _9098__34 (.L_HI(net34));
 sg13g2_tiehi _8806__35 (.L_HI(net35));
 sg13g2_tiehi _9001__36 (.L_HI(net36));
 sg13g2_tiehi _8805__37 (.L_HI(net37));
 sg13g2_tiehi _9111__38 (.L_HI(net38));
 sg13g2_tiehi _8804__39 (.L_HI(net39));
 sg13g2_tiehi _9000__40 (.L_HI(net40));
 sg13g2_tiehi _8803__41 (.L_HI(net41));
 sg13g2_tiehi _9097__42 (.L_HI(net42));
 sg13g2_tiehi _8802__43 (.L_HI(net43));
 sg13g2_tiehi _8999__44 (.L_HI(net44));
 sg13g2_tiehi _8801__45 (.L_HI(net45));
 sg13g2_tiehi _9092__46 (.L_HI(net46));
 sg13g2_tiehi _8800__47 (.L_HI(net47));
 sg13g2_tiehi _8998__48 (.L_HI(net48));
 sg13g2_tiehi _8799__49 (.L_HI(net49));
 sg13g2_tiehi _9096__50 (.L_HI(net50));
 sg13g2_tiehi _8798__51 (.L_HI(net51));
 sg13g2_tiehi _8997__52 (.L_HI(net52));
 sg13g2_tiehi _8797__53 (.L_HI(net53));
 sg13g2_tiehi _9110__54 (.L_HI(net54));
 sg13g2_tiehi _8796__55 (.L_HI(net55));
 sg13g2_tiehi _8996__56 (.L_HI(net56));
 sg13g2_tiehi _8795__57 (.L_HI(net57));
 sg13g2_tiehi _9095__58 (.L_HI(net58));
 sg13g2_tiehi _8794__59 (.L_HI(net59));
 sg13g2_tiehi _8995__60 (.L_HI(net60));
 sg13g2_tiehi _8793__61 (.L_HI(net61));
 sg13g2_tiehi _9115__62 (.L_HI(net62));
 sg13g2_tiehi _8792__63 (.L_HI(net63));
 sg13g2_tiehi _8994__64 (.L_HI(net64));
 sg13g2_tiehi _8791__65 (.L_HI(net65));
 sg13g2_tiehi _9094__66 (.L_HI(net66));
 sg13g2_tiehi _8790__67 (.L_HI(net67));
 sg13g2_tiehi _8993__68 (.L_HI(net68));
 sg13g2_tiehi _8789__69 (.L_HI(net69));
 sg13g2_tiehi _9093__70 (.L_HI(net70));
 sg13g2_tiehi _8788__71 (.L_HI(net71));
 sg13g2_tiehi _8992__72 (.L_HI(net72));
 sg13g2_tiehi _8787__73 (.L_HI(net73));
 sg13g2_tiehi _9028__74 (.L_HI(net74));
 sg13g2_tiehi _8786__75 (.L_HI(net75));
 sg13g2_tiehi _8991__76 (.L_HI(net76));
 sg13g2_tiehi _8785__77 (.L_HI(net77));
 sg13g2_tiehi _9027__78 (.L_HI(net78));
 sg13g2_tiehi _8784__79 (.L_HI(net79));
 sg13g2_tiehi _8990__80 (.L_HI(net80));
 sg13g2_tiehi _8783__81 (.L_HI(net81));
 sg13g2_tiehi _9026__82 (.L_HI(net82));
 sg13g2_tiehi _8782__83 (.L_HI(net83));
 sg13g2_tiehi _8989__84 (.L_HI(net84));
 sg13g2_tiehi _8781__85 (.L_HI(net85));
 sg13g2_tiehi _9025__86 (.L_HI(net86));
 sg13g2_tiehi _8780__87 (.L_HI(net87));
 sg13g2_tiehi _8988__88 (.L_HI(net88));
 sg13g2_tiehi _8779__89 (.L_HI(net89));
 sg13g2_tiehi _9109__90 (.L_HI(net90));
 sg13g2_tiehi _8778__91 (.L_HI(net91));
 sg13g2_tiehi _8987__92 (.L_HI(net92));
 sg13g2_tiehi _8777__93 (.L_HI(net93));
 sg13g2_tiehi _9024__94 (.L_HI(net94));
 sg13g2_tiehi _8776__95 (.L_HI(net95));
 sg13g2_tiehi _8986__96 (.L_HI(net96));
 sg13g2_tiehi _8775__97 (.L_HI(net97));
 sg13g2_tiehi _9114__98 (.L_HI(net98));
 sg13g2_tiehi _8774__99 (.L_HI(net99));
 sg13g2_tiehi _8985__100 (.L_HI(net100));
 sg13g2_tiehi _8773__101 (.L_HI(net101));
 sg13g2_tiehi _9023__102 (.L_HI(net102));
 sg13g2_tiehi _8772__103 (.L_HI(net103));
 sg13g2_tiehi _8984__104 (.L_HI(net104));
 sg13g2_tiehi _8771__105 (.L_HI(net105));
 sg13g2_tiehi _9022__106 (.L_HI(net106));
 sg13g2_tiehi _8770__107 (.L_HI(net107));
 sg13g2_tiehi _8983__108 (.L_HI(net108));
 sg13g2_tiehi _8769__109 (.L_HI(net109));
 sg13g2_tiehi _9021__110 (.L_HI(net110));
 sg13g2_tiehi _8768__111 (.L_HI(net111));
 sg13g2_tiehi _8982__112 (.L_HI(net112));
 sg13g2_tiehi _8767__113 (.L_HI(net113));
 sg13g2_tiehi _9020__114 (.L_HI(net114));
 sg13g2_tiehi _8766__115 (.L_HI(net115));
 sg13g2_tiehi _8981__116 (.L_HI(net116));
 sg13g2_tiehi _8765__117 (.L_HI(net117));
 sg13g2_tiehi _8980__118 (.L_HI(net118));
 sg13g2_tiehi _8764__119 (.L_HI(net119));
 sg13g2_tiehi _8979__120 (.L_HI(net120));
 sg13g2_tiehi _8763__121 (.L_HI(net121));
 sg13g2_tiehi _9108__122 (.L_HI(net122));
 sg13g2_tiehi _8762__123 (.L_HI(net123));
 sg13g2_tiehi _8978__124 (.L_HI(net124));
 sg13g2_tiehi _8761__125 (.L_HI(net125));
 sg13g2_tiehi _9019__126 (.L_HI(net126));
 sg13g2_tiehi _8760__127 (.L_HI(net127));
 sg13g2_tiehi _8976__128 (.L_HI(net128));
 sg13g2_tiehi _8759__129 (.L_HI(net129));
 sg13g2_tiehi _9117__130 (.L_HI(net130));
 sg13g2_tiehi _8758__131 (.L_HI(net131));
 sg13g2_tiehi _8975__132 (.L_HI(net132));
 sg13g2_tiehi _8757__133 (.L_HI(net133));
 sg13g2_tiehi _9018__134 (.L_HI(net134));
 sg13g2_tiehi _8756__135 (.L_HI(net135));
 sg13g2_tiehi _8974__136 (.L_HI(net136));
 sg13g2_tiehi _8755__137 (.L_HI(net137));
 sg13g2_tiehi _9107__138 (.L_HI(net138));
 sg13g2_tiehi _8754__139 (.L_HI(net139));
 sg13g2_tiehi _8973__140 (.L_HI(net140));
 sg13g2_tiehi _8753__141 (.L_HI(net141));
 sg13g2_tiehi _9017__142 (.L_HI(net142));
 sg13g2_tiehi _8752__143 (.L_HI(net143));
 sg13g2_tiehi _8972__144 (.L_HI(net144));
 sg13g2_tiehi _8751__145 (.L_HI(net145));
 sg13g2_tiehi _9113__146 (.L_HI(net146));
 sg13g2_tiehi _8750__147 (.L_HI(net147));
 sg13g2_tiehi _8971__148 (.L_HI(net148));
 sg13g2_tiehi _8749__149 (.L_HI(net149));
 sg13g2_tiehi _9016__150 (.L_HI(net150));
 sg13g2_tiehi _8748__151 (.L_HI(net151));
 sg13g2_tiehi _8970__152 (.L_HI(net152));
 sg13g2_tiehi _8747__153 (.L_HI(net153));
 sg13g2_tiehi _9106__154 (.L_HI(net154));
 sg13g2_tiehi _8746__155 (.L_HI(net155));
 sg13g2_tiehi _8969__156 (.L_HI(net156));
 sg13g2_tiehi _8745__157 (.L_HI(net157));
 sg13g2_tiehi _8744__158 (.L_HI(net158));
 sg13g2_tiehi _8743__159 (.L_HI(net159));
 sg13g2_tiehi _8742__160 (.L_HI(net160));
 sg13g2_tiehi _8741__161 (.L_HI(net161));
 sg13g2_tiehi _8740__162 (.L_HI(net162));
 sg13g2_tiehi _8739__163 (.L_HI(net163));
 sg13g2_tiehi _8738__164 (.L_HI(net164));
 sg13g2_tiehi _8737__165 (.L_HI(net165));
 sg13g2_tiehi _8736__166 (.L_HI(net166));
 sg13g2_tiehi _8735__167 (.L_HI(net167));
 sg13g2_tiehi _8734__168 (.L_HI(net168));
 sg13g2_tiehi _8733__169 (.L_HI(net169));
 sg13g2_tiehi _8732__170 (.L_HI(net170));
 sg13g2_tiehi _8731__171 (.L_HI(net171));
 sg13g2_tiehi _8730__172 (.L_HI(net172));
 sg13g2_tiehi _8729__173 (.L_HI(net173));
 sg13g2_tiehi _9012__174 (.L_HI(net174));
 sg13g2_tiehi _8968__175 (.L_HI(net175));
 sg13g2_tiehi _8967__176 (.L_HI(net176));
 sg13g2_tiehi _8965__177 (.L_HI(net177));
 sg13g2_tiehi _8964__178 (.L_HI(net178));
 sg13g2_tiehi _8963__179 (.L_HI(net179));
 sg13g2_tiehi _8962__180 (.L_HI(net180));
 sg13g2_tiehi _8961__181 (.L_HI(net181));
 sg13g2_tiehi _8960__182 (.L_HI(net182));
 sg13g2_tiehi _8959__183 (.L_HI(net183));
 sg13g2_tiehi _8958__184 (.L_HI(net184));
 sg13g2_tiehi _8957__185 (.L_HI(net185));
 sg13g2_tiehi _8956__186 (.L_HI(net186));
 sg13g2_tiehi _8955__187 (.L_HI(net187));
 sg13g2_tiehi _8954__188 (.L_HI(net188));
 sg13g2_tiehi _8953__189 (.L_HI(net189));
 sg13g2_tiehi _8952__190 (.L_HI(net190));
 sg13g2_tiehi _8951__191 (.L_HI(net191));
 sg13g2_tiehi _8950__192 (.L_HI(net192));
 sg13g2_tiehi _8949__193 (.L_HI(net193));
 sg13g2_tiehi _8948__194 (.L_HI(net194));
 sg13g2_tiehi _8947__195 (.L_HI(net195));
 sg13g2_tiehi _8946__196 (.L_HI(net196));
 sg13g2_tiehi _8945__197 (.L_HI(net197));
 sg13g2_tiehi _8944__198 (.L_HI(net198));
 sg13g2_tiehi _8943__199 (.L_HI(net199));
 sg13g2_tiehi _8942__200 (.L_HI(net200));
 sg13g2_tiehi _8941__201 (.L_HI(net201));
 sg13g2_tiehi _8940__202 (.L_HI(net202));
 sg13g2_tiehi _8939__203 (.L_HI(net203));
 sg13g2_tiehi _8938__204 (.L_HI(net204));
 sg13g2_tiehi _8937__205 (.L_HI(net205));
 sg13g2_tiehi _8936__206 (.L_HI(net206));
 sg13g2_tiehi _8935__207 (.L_HI(net207));
 sg13g2_tiehi _8934__208 (.L_HI(net208));
 sg13g2_tiehi _8933__209 (.L_HI(net209));
 sg13g2_tiehi _8932__210 (.L_HI(net210));
 sg13g2_tiehi _8931__211 (.L_HI(net211));
 sg13g2_tiehi _9105__212 (.L_HI(net212));
 sg13g2_tiehi _8930__213 (.L_HI(net213));
 sg13g2_tiehi _8728__214 (.L_HI(net214));
 sg13g2_tiehi _8916__215 (.L_HI(net215));
 sg13g2_tiehi _9011__216 (.L_HI(net216));
 sg13g2_tiehi _8929__217 (.L_HI(net217));
 sg13g2_tiehi _9104__218 (.L_HI(net218));
 sg13g2_tiehi _8928__219 (.L_HI(net219));
 sg13g2_tiehi _9010__220 (.L_HI(net220));
 sg13g2_tiehi _8927__221 (.L_HI(net221));
 sg13g2_tiehi _9103__222 (.L_HI(net222));
 sg13g2_tiehi _8926__223 (.L_HI(net223));
 sg13g2_tiehi _9009__224 (.L_HI(net224));
 sg13g2_tiehi _8925__225 (.L_HI(net225));
 sg13g2_tiehi _9102__226 (.L_HI(net226));
 sg13g2_tiehi _8924__227 (.L_HI(net227));
 sg13g2_tiehi _9008__228 (.L_HI(net228));
 sg13g2_tiehi _8923__229 (.L_HI(net229));
 sg13g2_tiehi _9101__230 (.L_HI(net230));
 sg13g2_tiehi _8922__231 (.L_HI(net231));
 sg13g2_tiehi _9007__232 (.L_HI(net232));
 sg13g2_tiehi _8921__233 (.L_HI(net233));
 sg13g2_tiehi _9118__234 (.L_HI(net234));
 sg13g2_tiehi _8920__235 (.L_HI(net235));
 sg13g2_tiehi _9006__236 (.L_HI(net236));
 sg13g2_tiehi _8919__237 (.L_HI(net237));
 sg13g2_tiehi _8918__238 (.L_HI(net238));
 sg13g2_tiehi _9100__239 (.L_HI(net239));
 sg13g2_tiehi _8915__240 (.L_HI(net240));
 sg13g2_tiehi _8914__241 (.L_HI(net241));
 sg13g2_tiehi _8913__242 (.L_HI(net242));
 sg13g2_tiehi _8912__243 (.L_HI(net243));
 sg13g2_tiehi _8911__244 (.L_HI(net244));
 sg13g2_tiehi _8910__245 (.L_HI(net245));
 sg13g2_tiehi _8909__246 (.L_HI(net246));
 sg13g2_tiehi _8908__247 (.L_HI(net247));
 sg13g2_tiehi _8907__248 (.L_HI(net248));
 sg13g2_tiehi _8906__249 (.L_HI(net249));
 sg13g2_tiehi _8905__250 (.L_HI(net250));
 sg13g2_tiehi _8904__251 (.L_HI(net251));
 sg13g2_tiehi _8903__252 (.L_HI(net252));
 sg13g2_tiehi _8902__253 (.L_HI(net253));
 sg13g2_tiehi _8901__254 (.L_HI(net254));
 sg13g2_tiehi _8900__255 (.L_HI(net255));
 sg13g2_tiehi _8899__256 (.L_HI(net256));
 sg13g2_tiehi _8898__257 (.L_HI(net257));
 sg13g2_tiehi _8897__258 (.L_HI(net258));
 sg13g2_tiehi _8896__259 (.L_HI(net259));
 sg13g2_tiehi _8895__260 (.L_HI(net260));
 sg13g2_tiehi _9005__261 (.L_HI(net261));
 sg13g2_tiehi _8894__262 (.L_HI(net262));
 sg13g2_tiehi _8893__263 (.L_HI(net263));
 sg13g2_tiehi _8917__264 (.L_HI(net264));
 sg13g2_tiehi _8892__265 (.L_HI(net265));
 sg13g2_tiehi _8891__266 (.L_HI(net266));
 sg13g2_tiehi _8890__267 (.L_HI(net267));
 sg13g2_tiehi _8889__268 (.L_HI(net268));
 sg13g2_tiehi _8888__269 (.L_HI(net269));
 sg13g2_tiehi _8887__270 (.L_HI(net270));
 sg13g2_tiehi _8886__271 (.L_HI(net271));
 sg13g2_tiehi _8885__272 (.L_HI(net272));
 sg13g2_tiehi _8884__273 (.L_HI(net273));
 sg13g2_tiehi _8883__274 (.L_HI(net274));
 sg13g2_tiehi _8966__275 (.L_HI(net275));
 sg13g2_tiehi _8882__276 (.L_HI(net276));
 sg13g2_tiehi _8881__277 (.L_HI(net277));
 sg13g2_tiehi _8880__278 (.L_HI(net278));
 sg13g2_tiehi _8879__279 (.L_HI(net279));
 sg13g2_tiehi _8878__280 (.L_HI(net280));
 sg13g2_tiehi _8877__281 (.L_HI(net281));
 sg13g2_tiehi _8876__282 (.L_HI(net282));
 sg13g2_tiehi _8875__283 (.L_HI(net283));
 sg13g2_tiehi _8874__284 (.L_HI(net284));
 sg13g2_tiehi _9112__285 (.L_HI(net285));
 sg13g2_tiehi _8873__286 (.L_HI(net286));
 sg13g2_tiehi _8872__287 (.L_HI(net287));
 sg13g2_tiehi _8871__288 (.L_HI(net288));
 sg13g2_tiehi _8870__289 (.L_HI(net289));
 sg13g2_tiehi _8869__290 (.L_HI(net290));
 sg13g2_tiehi _8868__291 (.L_HI(net291));
 sg13g2_tiehi _8867__292 (.L_HI(net292));
 sg13g2_tiehi _8866__293 (.L_HI(net293));
 sg13g2_tiehi _8865__294 (.L_HI(net294));
 sg13g2_tiehi _8864__295 (.L_HI(net295));
 sg13g2_tiehi _8863__296 (.L_HI(net296));
 sg13g2_tiehi _8862__297 (.L_HI(net297));
 sg13g2_tiehi _8861__298 (.L_HI(net298));
 sg13g2_tiehi _8860__299 (.L_HI(net299));
 sg13g2_tiehi _8859__300 (.L_HI(net300));
 sg13g2_tiehi _8858__301 (.L_HI(net301));
 sg13g2_tiehi _8857__302 (.L_HI(net302));
 sg13g2_tiehi _8856__303 (.L_HI(net303));
 sg13g2_tiehi _8855__304 (.L_HI(net304));
 sg13g2_tiehi _8854__305 (.L_HI(net305));
 sg13g2_tiehi _9004__306 (.L_HI(net306));
 sg13g2_tiehi _8853__307 (.L_HI(net307));
 sg13g2_tiehi _8852__308 (.L_HI(net308));
 sg13g2_tiehi _8851__309 (.L_HI(net309));
 sg13g2_tiehi _8850__310 (.L_HI(net310));
 sg13g2_tiehi _8977__311 (.L_HI(net311));
 sg13g2_tiehi _9013__312 (.L_HI(net312));
 sg13g2_tiehi _9014__313 (.L_HI(net313));
 sg13g2_tiehi _8849__314 (.L_HI(net314));
 sg13g2_tiehi _8848__315 (.L_HI(net315));
 sg13g2_tiehi _8847__316 (.L_HI(net316));
 sg13g2_tiehi _8846__317 (.L_HI(net317));
 sg13g2_tiehi _8845__318 (.L_HI(net318));
 sg13g2_tiehi _8844__319 (.L_HI(net319));
 sg13g2_tiehi _8843__320 (.L_HI(net320));
 sg13g2_tiehi _8842__321 (.L_HI(net321));
 sg13g2_tiehi _8841__322 (.L_HI(net322));
 sg13g2_tiehi _8840__323 (.L_HI(net323));
 sg13g2_tiehi _8839__324 (.L_HI(net324));
 sg13g2_tiehi _8838__325 (.L_HI(net325));
 sg13g2_tiehi _8837__326 (.L_HI(net326));
 sg13g2_tiehi _9015__327 (.L_HI(net327));
 sg13g2_tiehi _9029__328 (.L_HI(net328));
 sg13g2_tiehi _9030__329 (.L_HI(net329));
 sg13g2_tiehi _9031__330 (.L_HI(net330));
 sg13g2_tiehi _9032__331 (.L_HI(net331));
 sg13g2_tiehi _9033__332 (.L_HI(net332));
 sg13g2_tiehi _9034__333 (.L_HI(net333));
 sg13g2_tiehi _9035__334 (.L_HI(net334));
 sg13g2_tiehi _9036__335 (.L_HI(net335));
 sg13g2_tiehi _9037__336 (.L_HI(net336));
 sg13g2_tiehi _9038__337 (.L_HI(net337));
 sg13g2_tiehi _9039__338 (.L_HI(net338));
 sg13g2_tiehi _9040__339 (.L_HI(net339));
 sg13g2_tiehi _9041__340 (.L_HI(net340));
 sg13g2_tiehi _9042__341 (.L_HI(net341));
 sg13g2_tiehi _9043__342 (.L_HI(net342));
 sg13g2_tiehi _9044__343 (.L_HI(net343));
 sg13g2_tiehi _9045__344 (.L_HI(net344));
 sg13g2_tiehi _9046__345 (.L_HI(net345));
 sg13g2_tiehi _9047__346 (.L_HI(net346));
 sg13g2_tiehi _9048__347 (.L_HI(net347));
 sg13g2_tiehi _9049__348 (.L_HI(net348));
 sg13g2_tiehi _9050__349 (.L_HI(net349));
 sg13g2_tiehi _9051__350 (.L_HI(net350));
 sg13g2_tiehi _9052__351 (.L_HI(net351));
 sg13g2_tiehi _9053__352 (.L_HI(net352));
 sg13g2_tiehi _9054__353 (.L_HI(net353));
 sg13g2_tiehi _9055__354 (.L_HI(net354));
 sg13g2_tiehi _9056__355 (.L_HI(net355));
 sg13g2_tiehi _9057__356 (.L_HI(net356));
 sg13g2_tiehi _9058__357 (.L_HI(net357));
 sg13g2_tiehi _9059__358 (.L_HI(net358));
 sg13g2_tiehi _9060__359 (.L_HI(net359));
 sg13g2_tiehi _9061__360 (.L_HI(net360));
 sg13g2_tiehi _9062__361 (.L_HI(net361));
 sg13g2_tiehi _9063__362 (.L_HI(net362));
 sg13g2_tiehi _9064__363 (.L_HI(net363));
 sg13g2_tiehi _9065__364 (.L_HI(net364));
 sg13g2_tiehi _9066__365 (.L_HI(net365));
 sg13g2_tiehi _9067__366 (.L_HI(net366));
 sg13g2_tiehi _9068__367 (.L_HI(net367));
 sg13g2_tiehi _9069__368 (.L_HI(net368));
 sg13g2_tiehi _9070__369 (.L_HI(net369));
 sg13g2_tiehi _9071__370 (.L_HI(net370));
 sg13g2_tiehi _9072__371 (.L_HI(net371));
 sg13g2_tiehi _9073__372 (.L_HI(net372));
 sg13g2_tiehi _9074__373 (.L_HI(net373));
 sg13g2_tiehi _9075__374 (.L_HI(net374));
 sg13g2_tiehi _9076__375 (.L_HI(net375));
 sg13g2_tiehi _9077__376 (.L_HI(net376));
 sg13g2_tiehi _9078__377 (.L_HI(net377));
 sg13g2_tiehi _9079__378 (.L_HI(net378));
 sg13g2_tiehi _9080__379 (.L_HI(net379));
 sg13g2_tiehi _9081__380 (.L_HI(net380));
 sg13g2_tiehi _9082__381 (.L_HI(net381));
 sg13g2_tiehi _9083__382 (.L_HI(net382));
 sg13g2_tiehi _9084__383 (.L_HI(net383));
 sg13g2_tiehi _9085__384 (.L_HI(net384));
 sg13g2_tiehi _9086__385 (.L_HI(net385));
 sg13g2_tiehi _9087__386 (.L_HI(net386));
 sg13g2_tiehi _9088__387 (.L_HI(net387));
 sg13g2_tiehi _9089__388 (.L_HI(net388));
 sg13g2_tiehi _9090__389 (.L_HI(net389));
 sg13g2_tiehi _9091__390 (.L_HI(net390));
 sg13g2_tiehi _8836__391 (.L_HI(net391));
 sg13g2_tiehi _8835__392 (.L_HI(net392));
 sg13g2_tiehi _8834__393 (.L_HI(net393));
 sg13g2_tiehi _8833__394 (.L_HI(net394));
 sg13g2_tiehi _9099__395 (.L_HI(net395));
 sg13g2_tiehi _8832__396 (.L_HI(net396));
 sg13g2_tiehi _8831__397 (.L_HI(net397));
 sg13g2_tiehi _8830__398 (.L_HI(net398));
 sg13g2_tiehi _8829__399 (.L_HI(net399));
 sg13g2_tiehi _8828__400 (.L_HI(net400));
 sg13g2_tiehi _8827__401 (.L_HI(net401));
 sg13g2_tiehi _8826__402 (.L_HI(net402));
 sg13g2_tiehi _8825__403 (.L_HI(net403));
 sg13g2_tiehi _8824__404 (.L_HI(net404));
 sg13g2_tiehi _8823__405 (.L_HI(net405));
 sg13g2_tiehi _8822__406 (.L_HI(net406));
 sg13g2_tiehi _8821__407 (.L_HI(net407));
 sg13g2_tiehi _8820__408 (.L_HI(net408));
 sg13g2_tiehi _8819__409 (.L_HI(net409));
 sg13g2_tiehi _8818__410 (.L_HI(net410));
 sg13g2_tiehi _8817__411 (.L_HI(net411));
 sg13g2_tiehi _8816__412 (.L_HI(net412));
 sg13g2_tiehi _8815__413 (.L_HI(net413));
 sg13g2_tiehi _8814__414 (.L_HI(net414));
 sg13g2_tiehi _8813__415 (.L_HI(net415));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_2048_vga_game_18 (.L_LO(net18));
 sg13g2_tielo tt_um_2048_vga_game_19 (.L_LO(net19));
 sg13g2_tielo tt_um_2048_vga_game_20 (.L_LO(net20));
 sg13g2_tielo tt_um_2048_vga_game_21 (.L_LO(net21));
 sg13g2_tielo tt_um_2048_vga_game_22 (.L_LO(net22));
 sg13g2_tielo tt_um_2048_vga_game_23 (.L_LO(net23));
 sg13g2_tielo tt_um_2048_vga_game_24 (.L_LO(net24));
 sg13g2_tiehi _8812__25 (.L_HI(net25));
 sg13g2_buf_1 _9518_ (.A(\debug_controller_inst.data_out_en ),
    .X(uio_oe[4]));
 sg13g2_buf_1 _9519_ (.A(\debug_controller_inst.data_out_en ),
    .X(uio_oe[5]));
 sg13g2_buf_1 _9520_ (.A(\debug_controller_inst.data_out_en ),
    .X(uio_oe[6]));
 sg13g2_buf_1 _9521_ (.A(\debug_controller_inst.data_out_en ),
    .X(uio_oe[7]));
 sg13g2_buf_2 _9522_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _9523_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout1756 (.A(_1537_),
    .X(net1756));
 sg13g2_buf_2 fanout1757 (.A(_1537_),
    .X(net1757));
 sg13g2_buf_4 fanout1758 (.X(net1758),
    .A(_0861_));
 sg13g2_buf_4 fanout1759 (.X(net1759),
    .A(net1760));
 sg13g2_buf_4 fanout1760 (.X(net1760),
    .A(_0761_));
 sg13g2_buf_2 fanout1761 (.A(net1763),
    .X(net1761));
 sg13g2_buf_1 fanout1762 (.A(net1763),
    .X(net1762));
 sg13g2_buf_2 fanout1763 (.A(net1769),
    .X(net1763));
 sg13g2_buf_2 fanout1764 (.A(net1766),
    .X(net1764));
 sg13g2_buf_2 fanout1765 (.A(net1766),
    .X(net1765));
 sg13g2_buf_2 fanout1766 (.A(net1769),
    .X(net1766));
 sg13g2_buf_2 fanout1767 (.A(net1768),
    .X(net1767));
 sg13g2_buf_2 fanout1768 (.A(net1769),
    .X(net1768));
 sg13g2_buf_1 fanout1769 (.A(_0760_),
    .X(net1769));
 sg13g2_buf_4 fanout1770 (.X(net1770),
    .A(_1733_));
 sg13g2_buf_4 fanout1771 (.X(net1771),
    .A(_1663_));
 sg13g2_buf_4 fanout1772 (.X(net1772),
    .A(_1615_));
 sg13g2_buf_4 fanout1773 (.X(net1773),
    .A(net1774));
 sg13g2_buf_2 fanout1774 (.A(_1165_),
    .X(net1774));
 sg13g2_buf_4 fanout1775 (.X(net1775),
    .A(net1776));
 sg13g2_buf_4 fanout1776 (.X(net1776),
    .A(net1779));
 sg13g2_buf_4 fanout1777 (.X(net1777),
    .A(net1778));
 sg13g2_buf_4 fanout1778 (.X(net1778),
    .A(net1779));
 sg13g2_buf_2 fanout1779 (.A(net1781),
    .X(net1779));
 sg13g2_buf_4 fanout1780 (.X(net1780),
    .A(net1781));
 sg13g2_buf_2 fanout1781 (.A(_0865_),
    .X(net1781));
 sg13g2_buf_2 fanout1782 (.A(net1787),
    .X(net1782));
 sg13g2_buf_1 fanout1783 (.A(net1787),
    .X(net1783));
 sg13g2_buf_2 fanout1784 (.A(net1786),
    .X(net1784));
 sg13g2_buf_2 fanout1785 (.A(net1786),
    .X(net1785));
 sg13g2_buf_2 fanout1786 (.A(net1787),
    .X(net1786));
 sg13g2_buf_2 fanout1787 (.A(_0859_),
    .X(net1787));
 sg13g2_buf_2 fanout1788 (.A(net1790),
    .X(net1788));
 sg13g2_buf_1 fanout1789 (.A(net1790),
    .X(net1789));
 sg13g2_buf_2 fanout1790 (.A(_0859_),
    .X(net1790));
 sg13g2_buf_2 fanout1791 (.A(net1792),
    .X(net1791));
 sg13g2_buf_4 fanout1792 (.X(net1792),
    .A(_0698_));
 sg13g2_buf_2 fanout1793 (.A(net1794),
    .X(net1793));
 sg13g2_buf_2 fanout1794 (.A(net1795),
    .X(net1794));
 sg13g2_buf_2 fanout1795 (.A(_0697_),
    .X(net1795));
 sg13g2_buf_2 fanout1796 (.A(_0618_),
    .X(net1796));
 sg13g2_buf_2 fanout1797 (.A(net1799),
    .X(net1797));
 sg13g2_buf_2 fanout1798 (.A(net1799),
    .X(net1798));
 sg13g2_buf_2 fanout1799 (.A(_3755_),
    .X(net1799));
 sg13g2_buf_2 fanout1800 (.A(_3667_),
    .X(net1800));
 sg13g2_buf_2 fanout1801 (.A(_3667_),
    .X(net1801));
 sg13g2_buf_2 fanout1802 (.A(net1803),
    .X(net1802));
 sg13g2_buf_2 fanout1803 (.A(_3626_),
    .X(net1803));
 sg13g2_buf_2 fanout1804 (.A(_3584_),
    .X(net1804));
 sg13g2_buf_2 fanout1805 (.A(_3584_),
    .X(net1805));
 sg13g2_buf_2 fanout1806 (.A(net1807),
    .X(net1806));
 sg13g2_buf_2 fanout1807 (.A(_3541_),
    .X(net1807));
 sg13g2_buf_4 fanout1808 (.X(net1808),
    .A(_0508_));
 sg13g2_buf_2 fanout1809 (.A(_0507_),
    .X(net1809));
 sg13g2_buf_2 fanout1810 (.A(_0580_),
    .X(net1810));
 sg13g2_buf_2 fanout1811 (.A(net1812),
    .X(net1811));
 sg13g2_buf_2 fanout1812 (.A(_3493_),
    .X(net1812));
 sg13g2_buf_4 fanout1813 (.X(net1813),
    .A(_1940_));
 sg13g2_buf_4 fanout1814 (.X(net1814),
    .A(_1678_));
 sg13g2_buf_4 fanout1815 (.X(net1815),
    .A(_1447_));
 sg13g2_buf_2 fanout1816 (.A(_0579_),
    .X(net1816));
 sg13g2_buf_4 fanout1817 (.X(net1817),
    .A(_1964_));
 sg13g2_buf_4 fanout1818 (.X(net1818),
    .A(_1865_));
 sg13g2_buf_4 fanout1819 (.X(net1819),
    .A(_1854_));
 sg13g2_buf_4 fanout1820 (.X(net1820),
    .A(_1783_));
 sg13g2_buf_4 fanout1821 (.X(net1821),
    .A(_1677_));
 sg13g2_buf_4 fanout1822 (.X(net1822),
    .A(net1823));
 sg13g2_buf_4 fanout1823 (.X(net1823),
    .A(_1669_));
 sg13g2_buf_4 fanout1824 (.X(net1824),
    .A(_1658_));
 sg13g2_buf_4 fanout1825 (.X(net1825),
    .A(_1646_));
 sg13g2_buf_2 fanout1826 (.A(_1646_),
    .X(net1826));
 sg13g2_buf_4 fanout1827 (.X(net1827),
    .A(net1828));
 sg13g2_buf_4 fanout1828 (.X(net1828),
    .A(net1829));
 sg13g2_buf_2 fanout1829 (.A(_1645_),
    .X(net1829));
 sg13g2_buf_4 fanout1830 (.X(net1830),
    .A(net1831));
 sg13g2_buf_4 fanout1831 (.X(net1831),
    .A(_1641_));
 sg13g2_buf_4 fanout1832 (.X(net1832),
    .A(_1633_));
 sg13g2_buf_2 fanout1833 (.A(_1633_),
    .X(net1833));
 sg13g2_buf_2 fanout1834 (.A(_1632_),
    .X(net1834));
 sg13g2_buf_4 fanout1835 (.X(net1835),
    .A(_1619_));
 sg13g2_buf_4 fanout1836 (.X(net1836),
    .A(net1837));
 sg13g2_buf_4 fanout1837 (.X(net1837),
    .A(_1618_));
 sg13g2_buf_4 fanout1838 (.X(net1838),
    .A(net1839));
 sg13g2_buf_4 fanout1839 (.X(net1839),
    .A(_1562_));
 sg13g2_buf_4 fanout1840 (.X(net1840),
    .A(_1557_));
 sg13g2_buf_2 fanout1841 (.A(net1842),
    .X(net1841));
 sg13g2_buf_2 fanout1842 (.A(_3945_),
    .X(net1842));
 sg13g2_buf_4 fanout1843 (.X(net1843),
    .A(_3851_));
 sg13g2_buf_4 fanout1844 (.X(net1844),
    .A(_3730_));
 sg13g2_buf_2 fanout1845 (.A(_3730_),
    .X(net1845));
 sg13g2_buf_4 fanout1846 (.X(net1846),
    .A(_3700_));
 sg13g2_buf_2 fanout1847 (.A(_3700_),
    .X(net1847));
 sg13g2_buf_4 fanout1848 (.X(net1848),
    .A(_2068_));
 sg13g2_buf_2 fanout1849 (.A(_2068_),
    .X(net1849));
 sg13g2_buf_4 fanout1850 (.X(net1850),
    .A(_2033_));
 sg13g2_buf_4 fanout1851 (.X(net1851),
    .A(_1879_));
 sg13g2_buf_4 fanout1852 (.X(net1852),
    .A(net1853));
 sg13g2_buf_4 fanout1853 (.X(net1853),
    .A(_1878_));
 sg13g2_buf_4 fanout1854 (.X(net1854),
    .A(_1801_));
 sg13g2_buf_4 fanout1855 (.X(net1855),
    .A(net1857));
 sg13g2_buf_2 fanout1856 (.A(net1857),
    .X(net1856));
 sg13g2_buf_4 fanout1857 (.X(net1857),
    .A(_1800_));
 sg13g2_buf_4 fanout1858 (.X(net1858),
    .A(_1785_));
 sg13g2_buf_4 fanout1859 (.X(net1859),
    .A(_1784_));
 sg13g2_buf_2 fanout1860 (.A(_1784_),
    .X(net1860));
 sg13g2_buf_4 fanout1861 (.X(net1861),
    .A(net1862));
 sg13g2_buf_2 fanout1862 (.A(_1773_),
    .X(net1862));
 sg13g2_buf_4 fanout1863 (.X(net1863),
    .A(_1762_));
 sg13g2_buf_2 fanout1864 (.A(_1762_),
    .X(net1864));
 sg13g2_buf_2 fanout1865 (.A(net1867),
    .X(net1865));
 sg13g2_buf_1 fanout1866 (.A(net1867),
    .X(net1866));
 sg13g2_buf_2 fanout1867 (.A(_1636_),
    .X(net1867));
 sg13g2_buf_4 fanout1868 (.X(net1868),
    .A(_1636_));
 sg13g2_buf_4 fanout1869 (.X(net1869),
    .A(_1630_));
 sg13g2_buf_4 fanout1870 (.X(net1870),
    .A(_1630_));
 sg13g2_buf_4 fanout1871 (.X(net1871),
    .A(_1629_));
 sg13g2_buf_2 fanout1872 (.A(_1629_),
    .X(net1872));
 sg13g2_buf_4 fanout1873 (.X(net1873),
    .A(net1874));
 sg13g2_buf_2 fanout1874 (.A(net1875),
    .X(net1874));
 sg13g2_buf_4 fanout1875 (.X(net1875),
    .A(_1622_));
 sg13g2_buf_4 fanout1876 (.X(net1876),
    .A(net1877));
 sg13g2_buf_4 fanout1877 (.X(net1877),
    .A(net1878));
 sg13g2_buf_4 fanout1878 (.X(net1878),
    .A(_1621_));
 sg13g2_buf_4 fanout1879 (.X(net1879),
    .A(net1880));
 sg13g2_buf_4 fanout1880 (.X(net1880),
    .A(_1617_));
 sg13g2_buf_4 fanout1881 (.X(net1881),
    .A(net1882));
 sg13g2_buf_4 fanout1882 (.X(net1882),
    .A(_1616_));
 sg13g2_buf_4 fanout1883 (.X(net1883),
    .A(net1885));
 sg13g2_buf_2 fanout1884 (.A(net1885),
    .X(net1884));
 sg13g2_buf_4 fanout1885 (.X(net1885),
    .A(_1592_));
 sg13g2_buf_4 fanout1886 (.X(net1886),
    .A(net1889));
 sg13g2_buf_2 fanout1887 (.A(net1889),
    .X(net1887));
 sg13g2_buf_4 fanout1888 (.X(net1888),
    .A(net1889));
 sg13g2_buf_4 fanout1889 (.X(net1889),
    .A(_1592_));
 sg13g2_buf_4 fanout1890 (.X(net1890),
    .A(net1891));
 sg13g2_buf_8 fanout1891 (.A(_1585_),
    .X(net1891));
 sg13g2_buf_4 fanout1892 (.X(net1892),
    .A(net1896));
 sg13g2_buf_2 fanout1893 (.A(net1895),
    .X(net1893));
 sg13g2_buf_2 fanout1894 (.A(net1895),
    .X(net1894));
 sg13g2_buf_2 fanout1895 (.A(net1896),
    .X(net1895));
 sg13g2_buf_2 fanout1896 (.A(_1585_),
    .X(net1896));
 sg13g2_buf_4 fanout1897 (.X(net1897),
    .A(net1898));
 sg13g2_buf_4 fanout1898 (.X(net1898),
    .A(net1899));
 sg13g2_buf_2 fanout1899 (.A(net1900),
    .X(net1899));
 sg13g2_buf_4 fanout1900 (.X(net1900),
    .A(_1563_));
 sg13g2_buf_4 fanout1901 (.X(net1901),
    .A(net1902));
 sg13g2_buf_4 fanout1902 (.X(net1902),
    .A(_1561_));
 sg13g2_buf_4 fanout1903 (.X(net1903),
    .A(_1560_));
 sg13g2_buf_8 fanout1904 (.A(_1552_),
    .X(net1904));
 sg13g2_buf_4 fanout1905 (.X(net1905),
    .A(net1908));
 sg13g2_buf_2 fanout1906 (.A(net1908),
    .X(net1906));
 sg13g2_buf_4 fanout1907 (.X(net1907),
    .A(net1908));
 sg13g2_buf_4 fanout1908 (.X(net1908),
    .A(_1551_));
 sg13g2_buf_4 fanout1909 (.X(net1909),
    .A(_1549_));
 sg13g2_buf_2 fanout1910 (.A(_1549_),
    .X(net1910));
 sg13g2_buf_4 fanout1911 (.X(net1911),
    .A(_1546_));
 sg13g2_buf_4 fanout1912 (.X(net1912),
    .A(net1915));
 sg13g2_buf_4 fanout1913 (.X(net1913),
    .A(net1915));
 sg13g2_buf_4 fanout1914 (.X(net1914),
    .A(net1915));
 sg13g2_buf_8 fanout1915 (.A(_1544_),
    .X(net1915));
 sg13g2_buf_4 fanout1916 (.X(net1916),
    .A(net1917));
 sg13g2_buf_2 fanout1917 (.A(_1543_),
    .X(net1917));
 sg13g2_buf_4 fanout1918 (.X(net1918),
    .A(_1543_));
 sg13g2_buf_4 fanout1919 (.X(net1919),
    .A(_1543_));
 sg13g2_buf_4 fanout1920 (.X(net1920),
    .A(net1921));
 sg13g2_buf_4 fanout1921 (.X(net1921),
    .A(_1542_));
 sg13g2_buf_4 fanout1922 (.X(net1922),
    .A(_1541_));
 sg13g2_buf_2 fanout1923 (.A(_1541_),
    .X(net1923));
 sg13g2_buf_4 fanout1924 (.X(net1924),
    .A(net1928));
 sg13g2_buf_2 fanout1925 (.A(net1928),
    .X(net1925));
 sg13g2_buf_4 fanout1926 (.X(net1926),
    .A(net1928));
 sg13g2_buf_2 fanout1927 (.A(net1928),
    .X(net1927));
 sg13g2_buf_2 fanout1928 (.A(_1477_),
    .X(net1928));
 sg13g2_buf_4 fanout1929 (.X(net1929),
    .A(net1931));
 sg13g2_buf_2 fanout1930 (.A(net1931),
    .X(net1930));
 sg13g2_buf_4 fanout1931 (.X(net1931),
    .A(_1475_));
 sg13g2_buf_2 fanout1932 (.A(net1933),
    .X(net1932));
 sg13g2_buf_2 fanout1933 (.A(net1934),
    .X(net1933));
 sg13g2_buf_4 fanout1934 (.X(net1934),
    .A(_1433_));
 sg13g2_buf_4 fanout1935 (.X(net1935),
    .A(_1433_));
 sg13g2_buf_4 fanout1936 (.X(net1936),
    .A(_1433_));
 sg13g2_buf_4 fanout1937 (.X(net1937),
    .A(net1938));
 sg13g2_buf_4 fanout1938 (.X(net1938),
    .A(net1941));
 sg13g2_buf_4 fanout1939 (.X(net1939),
    .A(net1941));
 sg13g2_buf_4 fanout1940 (.X(net1940),
    .A(net1941));
 sg13g2_buf_2 fanout1941 (.A(_1432_),
    .X(net1941));
 sg13g2_buf_4 fanout1942 (.X(net1942),
    .A(net1943));
 sg13g2_buf_4 fanout1943 (.X(net1943),
    .A(_1429_));
 sg13g2_buf_4 fanout1944 (.X(net1944),
    .A(net1946));
 sg13g2_buf_1 fanout1945 (.A(net1946),
    .X(net1945));
 sg13g2_buf_4 fanout1946 (.X(net1946),
    .A(_1429_));
 sg13g2_buf_4 fanout1947 (.X(net1947),
    .A(net1948));
 sg13g2_buf_4 fanout1948 (.X(net1948),
    .A(net1949));
 sg13g2_buf_4 fanout1949 (.X(net1949),
    .A(_1428_));
 sg13g2_buf_4 fanout1950 (.X(net1950),
    .A(_1428_));
 sg13g2_buf_4 fanout1951 (.X(net1951),
    .A(_1019_));
 sg13g2_buf_2 fanout1952 (.A(_1019_),
    .X(net1952));
 sg13g2_buf_4 fanout1953 (.X(net1953),
    .A(_1018_));
 sg13g2_buf_4 fanout1954 (.X(net1954),
    .A(_0630_));
 sg13g2_buf_4 fanout1955 (.X(net1955),
    .A(_0551_));
 sg13g2_buf_4 fanout1956 (.X(net1956),
    .A(_0536_));
 sg13g2_buf_2 fanout1957 (.A(net1958),
    .X(net1957));
 sg13g2_buf_2 fanout1958 (.A(_3729_),
    .X(net1958));
 sg13g2_buf_2 fanout1959 (.A(_3699_),
    .X(net1959));
 sg13g2_buf_1 fanout1960 (.A(_3699_),
    .X(net1960));
 sg13g2_buf_2 fanout1961 (.A(net1963),
    .X(net1961));
 sg13g2_buf_1 fanout1962 (.A(net1963),
    .X(net1962));
 sg13g2_buf_2 fanout1963 (.A(net1967),
    .X(net1963));
 sg13g2_buf_2 fanout1964 (.A(net1965),
    .X(net1964));
 sg13g2_buf_1 fanout1965 (.A(net1966),
    .X(net1965));
 sg13g2_buf_2 fanout1966 (.A(net1967),
    .X(net1966));
 sg13g2_buf_4 fanout1967 (.X(net1967),
    .A(_3340_));
 sg13g2_buf_2 fanout1968 (.A(net1973),
    .X(net1968));
 sg13g2_buf_2 fanout1969 (.A(net1970),
    .X(net1969));
 sg13g2_buf_2 fanout1970 (.A(net1973),
    .X(net1970));
 sg13g2_buf_2 fanout1971 (.A(net1972),
    .X(net1971));
 sg13g2_buf_2 fanout1972 (.A(net1973),
    .X(net1972));
 sg13g2_buf_2 fanout1973 (.A(_3339_),
    .X(net1973));
 sg13g2_buf_2 fanout1974 (.A(net1976),
    .X(net1974));
 sg13g2_buf_1 fanout1975 (.A(net1976),
    .X(net1975));
 sg13g2_buf_2 fanout1976 (.A(net1979),
    .X(net1976));
 sg13g2_buf_2 fanout1977 (.A(net1979),
    .X(net1977));
 sg13g2_buf_1 fanout1978 (.A(net1979),
    .X(net1978));
 sg13g2_buf_2 fanout1979 (.A(_3339_),
    .X(net1979));
 sg13g2_buf_4 fanout1980 (.X(net1980),
    .A(net1981));
 sg13g2_buf_8 fanout1981 (.A(_1760_),
    .X(net1981));
 sg13g2_buf_2 fanout1982 (.A(_1760_),
    .X(net1982));
 sg13g2_buf_4 fanout1983 (.X(net1983),
    .A(_1759_));
 sg13g2_buf_4 fanout1984 (.X(net1984),
    .A(_1759_));
 sg13g2_buf_4 fanout1985 (.X(net1985),
    .A(_1690_));
 sg13g2_buf_4 fanout1986 (.X(net1986),
    .A(net1987));
 sg13g2_buf_2 fanout1987 (.A(_1593_),
    .X(net1987));
 sg13g2_buf_4 fanout1988 (.X(net1988),
    .A(net1990));
 sg13g2_buf_1 fanout1989 (.A(net1990),
    .X(net1989));
 sg13g2_buf_4 fanout1990 (.X(net1990),
    .A(_1593_));
 sg13g2_buf_4 fanout1991 (.X(net1991),
    .A(net1993));
 sg13g2_buf_1 fanout1992 (.A(net1993),
    .X(net1992));
 sg13g2_buf_4 fanout1993 (.X(net1993),
    .A(_1586_));
 sg13g2_buf_4 fanout1994 (.X(net1994),
    .A(_1586_));
 sg13g2_buf_4 fanout1995 (.X(net1995),
    .A(_1586_));
 sg13g2_buf_4 fanout1996 (.X(net1996),
    .A(net1999));
 sg13g2_buf_4 fanout1997 (.X(net1997),
    .A(net1999));
 sg13g2_buf_4 fanout1998 (.X(net1998),
    .A(net1999));
 sg13g2_buf_4 fanout1999 (.X(net1999),
    .A(_1581_));
 sg13g2_buf_4 fanout2000 (.X(net2000),
    .A(net2001));
 sg13g2_buf_8 fanout2001 (.A(_1553_),
    .X(net2001));
 sg13g2_buf_4 fanout2002 (.X(net2002),
    .A(net2003));
 sg13g2_buf_4 fanout2003 (.X(net2003),
    .A(_1550_));
 sg13g2_buf_4 fanout2004 (.X(net2004),
    .A(_1540_));
 sg13g2_buf_4 fanout2005 (.X(net2005),
    .A(_1540_));
 sg13g2_buf_4 fanout2006 (.X(net2006),
    .A(_1539_));
 sg13g2_buf_4 fanout2007 (.X(net2007),
    .A(_1539_));
 sg13g2_buf_4 fanout2008 (.X(net2008),
    .A(net2009));
 sg13g2_buf_4 fanout2009 (.X(net2009),
    .A(net2012));
 sg13g2_buf_2 fanout2010 (.A(net2011),
    .X(net2010));
 sg13g2_buf_4 fanout2011 (.X(net2011),
    .A(net2012));
 sg13g2_buf_2 fanout2012 (.A(_1476_),
    .X(net2012));
 sg13g2_buf_4 fanout2013 (.X(net2013),
    .A(net2016));
 sg13g2_buf_4 fanout2014 (.X(net2014),
    .A(net2016));
 sg13g2_buf_4 fanout2015 (.X(net2015),
    .A(net2016));
 sg13g2_buf_4 fanout2016 (.X(net2016),
    .A(_1474_));
 sg13g2_buf_4 fanout2017 (.X(net2017),
    .A(_1459_));
 sg13g2_buf_2 fanout2018 (.A(_1459_),
    .X(net2018));
 sg13g2_buf_4 fanout2019 (.X(net2019),
    .A(_1444_));
 sg13g2_buf_2 fanout2020 (.A(net2021),
    .X(net2020));
 sg13g2_buf_4 fanout2021 (.X(net2021),
    .A(_1444_));
 sg13g2_buf_4 fanout2022 (.X(net2022),
    .A(_1442_));
 sg13g2_buf_4 fanout2023 (.X(net2023),
    .A(_1438_));
 sg13g2_buf_2 fanout2024 (.A(_1438_),
    .X(net2024));
 sg13g2_buf_2 fanout2025 (.A(net2028),
    .X(net2025));
 sg13g2_buf_2 fanout2026 (.A(net2028),
    .X(net2026));
 sg13g2_buf_4 fanout2027 (.X(net2027),
    .A(net2028));
 sg13g2_buf_2 fanout2028 (.A(_1438_),
    .X(net2028));
 sg13g2_buf_4 fanout2029 (.X(net2029),
    .A(_1434_));
 sg13g2_buf_4 fanout2030 (.X(net2030),
    .A(_1434_));
 sg13g2_buf_4 fanout2031 (.X(net2031),
    .A(_1425_));
 sg13g2_buf_4 fanout2032 (.X(net2032),
    .A(net2033));
 sg13g2_buf_4 fanout2033 (.X(net2033),
    .A(_0864_));
 sg13g2_buf_4 fanout2034 (.X(net2034),
    .A(_0863_));
 sg13g2_buf_4 fanout2035 (.X(net2035),
    .A(_0701_));
 sg13g2_buf_2 fanout2036 (.A(net2038),
    .X(net2036));
 sg13g2_buf_4 fanout2037 (.X(net2037),
    .A(net2038));
 sg13g2_buf_2 fanout2038 (.A(_0528_),
    .X(net2038));
 sg13g2_buf_2 fanout2039 (.A(net2040),
    .X(net2039));
 sg13g2_buf_2 fanout2040 (.A(_0527_),
    .X(net2040));
 sg13g2_buf_2 fanout2041 (.A(net2043),
    .X(net2041));
 sg13g2_buf_2 fanout2042 (.A(net2043),
    .X(net2042));
 sg13g2_buf_2 fanout2043 (.A(_0527_),
    .X(net2043));
 sg13g2_buf_2 fanout2044 (.A(net2045),
    .X(net2044));
 sg13g2_buf_2 fanout2045 (.A(_0525_),
    .X(net2045));
 sg13g2_buf_2 fanout2046 (.A(_0525_),
    .X(net2046));
 sg13g2_buf_1 fanout2047 (.A(_0525_),
    .X(net2047));
 sg13g2_buf_4 fanout2048 (.X(net2048),
    .A(_0524_));
 sg13g2_buf_2 fanout2049 (.A(_0524_),
    .X(net2049));
 sg13g2_buf_2 fanout2050 (.A(net2053),
    .X(net2050));
 sg13g2_buf_4 fanout2051 (.X(net2051),
    .A(net2053));
 sg13g2_buf_2 fanout2052 (.A(net2053),
    .X(net2052));
 sg13g2_buf_2 fanout2053 (.A(_0523_),
    .X(net2053));
 sg13g2_buf_2 fanout2054 (.A(net2056),
    .X(net2054));
 sg13g2_buf_2 fanout2055 (.A(net2056),
    .X(net2055));
 sg13g2_buf_4 fanout2056 (.X(net2056),
    .A(_0522_));
 sg13g2_buf_2 fanout2057 (.A(net2061),
    .X(net2057));
 sg13g2_buf_2 fanout2058 (.A(net2061),
    .X(net2058));
 sg13g2_buf_2 fanout2059 (.A(net2060),
    .X(net2059));
 sg13g2_buf_4 fanout2060 (.X(net2060),
    .A(net2061));
 sg13g2_buf_4 fanout2061 (.X(net2061),
    .A(_0521_));
 sg13g2_buf_4 fanout2062 (.X(net2062),
    .A(_4048_));
 sg13g2_buf_4 fanout2063 (.X(net2063),
    .A(net2064));
 sg13g2_buf_4 fanout2064 (.X(net2064),
    .A(_4047_));
 sg13g2_buf_2 fanout2065 (.A(net2066),
    .X(net2065));
 sg13g2_buf_4 fanout2066 (.X(net2066),
    .A(_4046_));
 sg13g2_buf_4 fanout2067 (.X(net2067),
    .A(net2068));
 sg13g2_buf_4 fanout2068 (.X(net2068),
    .A(net2078));
 sg13g2_buf_4 fanout2069 (.X(net2069),
    .A(net2078));
 sg13g2_buf_2 fanout2070 (.A(net2078),
    .X(net2070));
 sg13g2_buf_4 fanout2071 (.X(net2071),
    .A(net2073));
 sg13g2_buf_2 fanout2072 (.A(net2073),
    .X(net2072));
 sg13g2_buf_4 fanout2073 (.X(net2073),
    .A(net2078));
 sg13g2_buf_4 fanout2074 (.X(net2074),
    .A(net2077));
 sg13g2_buf_4 fanout2075 (.X(net2075),
    .A(net2077));
 sg13g2_buf_2 fanout2076 (.A(net2077),
    .X(net2076));
 sg13g2_buf_2 fanout2077 (.A(net2078),
    .X(net2077));
 sg13g2_buf_4 fanout2078 (.X(net2078),
    .A(_4045_));
 sg13g2_buf_4 fanout2079 (.X(net2079),
    .A(net2080));
 sg13g2_buf_4 fanout2080 (.X(net2080),
    .A(_4044_));
 sg13g2_buf_2 fanout2081 (.A(_4044_),
    .X(net2081));
 sg13g2_buf_4 fanout2082 (.X(net2082),
    .A(net2083));
 sg13g2_buf_2 fanout2083 (.A(net2084),
    .X(net2083));
 sg13g2_buf_4 fanout2084 (.X(net2084),
    .A(_4044_));
 sg13g2_buf_2 fanout2085 (.A(net2087),
    .X(net2085));
 sg13g2_buf_2 fanout2086 (.A(net2087),
    .X(net2086));
 sg13g2_buf_4 fanout2087 (.X(net2087),
    .A(net2090));
 sg13g2_buf_4 fanout2088 (.X(net2088),
    .A(net2089));
 sg13g2_buf_4 fanout2089 (.X(net2089),
    .A(net2090));
 sg13g2_buf_4 fanout2090 (.X(net2090),
    .A(_4043_));
 sg13g2_buf_4 fanout2091 (.X(net2091),
    .A(net2092));
 sg13g2_buf_4 fanout2092 (.X(net2092),
    .A(_4041_));
 sg13g2_buf_1 fanout2093 (.A(_4041_),
    .X(net2093));
 sg13g2_buf_4 fanout2094 (.X(net2094),
    .A(_4026_));
 sg13g2_buf_4 fanout2095 (.X(net2095),
    .A(net2096));
 sg13g2_buf_4 fanout2096 (.X(net2096),
    .A(net2103));
 sg13g2_buf_2 fanout2097 (.A(net2098),
    .X(net2097));
 sg13g2_buf_4 fanout2098 (.X(net2098),
    .A(net2103));
 sg13g2_buf_2 fanout2099 (.A(net2102),
    .X(net2099));
 sg13g2_buf_2 fanout2100 (.A(net2101),
    .X(net2100));
 sg13g2_buf_2 fanout2101 (.A(net2102),
    .X(net2101));
 sg13g2_buf_2 fanout2102 (.A(net2103),
    .X(net2102));
 sg13g2_buf_2 fanout2103 (.A(_4023_),
    .X(net2103));
 sg13g2_buf_4 fanout2104 (.X(net2104),
    .A(net2105));
 sg13g2_buf_4 fanout2105 (.X(net2105),
    .A(net2106));
 sg13g2_buf_4 fanout2106 (.X(net2106),
    .A(_4022_));
 sg13g2_buf_4 fanout2107 (.X(net2107),
    .A(net2109));
 sg13g2_buf_2 fanout2108 (.A(net2109),
    .X(net2108));
 sg13g2_buf_2 fanout2109 (.A(net2110),
    .X(net2109));
 sg13g2_buf_4 fanout2110 (.X(net2110),
    .A(_4022_));
 sg13g2_buf_2 fanout2111 (.A(net2113),
    .X(net2111));
 sg13g2_buf_1 fanout2112 (.A(net2113),
    .X(net2112));
 sg13g2_buf_2 fanout2113 (.A(net2122),
    .X(net2113));
 sg13g2_buf_2 fanout2114 (.A(net2116),
    .X(net2114));
 sg13g2_buf_1 fanout2115 (.A(net2116),
    .X(net2115));
 sg13g2_buf_2 fanout2116 (.A(net2122),
    .X(net2116));
 sg13g2_buf_2 fanout2117 (.A(net2118),
    .X(net2117));
 sg13g2_buf_1 fanout2118 (.A(net2119),
    .X(net2118));
 sg13g2_buf_2 fanout2119 (.A(net2122),
    .X(net2119));
 sg13g2_buf_2 fanout2120 (.A(net2121),
    .X(net2120));
 sg13g2_buf_2 fanout2121 (.A(net2122),
    .X(net2121));
 sg13g2_buf_2 fanout2122 (.A(_4009_),
    .X(net2122));
 sg13g2_buf_2 fanout2123 (.A(_3978_),
    .X(net2123));
 sg13g2_buf_4 fanout2124 (.X(net2124),
    .A(_3977_));
 sg13g2_buf_2 fanout2125 (.A(net2126),
    .X(net2125));
 sg13g2_buf_1 fanout2126 (.A(net2127),
    .X(net2126));
 sg13g2_buf_2 fanout2127 (.A(net998),
    .X(net2127));
 sg13g2_buf_4 fanout2128 (.X(net2128),
    .A(net2130));
 sg13g2_buf_2 fanout2129 (.A(net2130),
    .X(net2129));
 sg13g2_buf_2 fanout2130 (.A(\debug_controller_inst.grid_addr[1] ),
    .X(net2130));
 sg13g2_buf_2 fanout2131 (.A(net2133),
    .X(net2131));
 sg13g2_buf_4 fanout2132 (.X(net2132),
    .A(net2133));
 sg13g2_buf_1 fanout2133 (.A(net2134),
    .X(net2133));
 sg13g2_buf_2 fanout2134 (.A(net2136),
    .X(net2134));
 sg13g2_buf_4 fanout2135 (.X(net2135),
    .A(net2136));
 sg13g2_buf_2 fanout2136 (.A(net1020),
    .X(net2136));
 sg13g2_buf_4 fanout2137 (.X(net2137),
    .A(net2138));
 sg13g2_buf_4 fanout2138 (.X(net2138),
    .A(net816));
 sg13g2_buf_4 fanout2139 (.X(net2139),
    .A(\debug_controller_inst.grid_out_addr[1] ));
 sg13g2_buf_4 fanout2140 (.X(net2140),
    .A(\debug_controller_inst.grid_out_addr[0] ));
 sg13g2_buf_4 fanout2141 (.X(net2141),
    .A(net995));
 sg13g2_buf_4 fanout2142 (.X(net2142),
    .A(net995));
 sg13g2_buf_4 fanout2143 (.X(net2143),
    .A(net2144));
 sg13g2_buf_4 fanout2144 (.X(net2144),
    .A(net989));
 sg13g2_buf_4 fanout2145 (.X(net2145),
    .A(net2147));
 sg13g2_buf_2 fanout2146 (.A(net2147),
    .X(net2146));
 sg13g2_buf_4 fanout2147 (.X(net2147),
    .A(net986));
 sg13g2_buf_4 fanout2148 (.X(net2148),
    .A(net1027));
 sg13g2_buf_2 fanout2149 (.A(net937),
    .X(net2149));
 sg13g2_buf_4 fanout2150 (.X(net2150),
    .A(net2151));
 sg13g2_buf_2 fanout2151 (.A(net2152),
    .X(net2151));
 sg13g2_buf_2 fanout2152 (.A(net2153),
    .X(net2152));
 sg13g2_buf_4 fanout2153 (.X(net2153),
    .A(net983));
 sg13g2_buf_8 fanout2154 (.A(net2155),
    .X(net2154));
 sg13g2_buf_4 fanout2155 (.X(net2155),
    .A(net2156));
 sg13g2_buf_2 fanout2156 (.A(net2157),
    .X(net2156));
 sg13g2_buf_4 fanout2157 (.X(net2157),
    .A(\game_logic_inst.current_row_index[0] ));
 sg13g2_buf_2 fanout2158 (.A(\game_logic_inst.added_tile_index[3] ),
    .X(net2158));
 sg13g2_buf_2 fanout2159 (.A(\game_logic_inst.added_tile_index[2] ),
    .X(net2159));
 sg13g2_buf_2 fanout2160 (.A(net851),
    .X(net2160));
 sg13g2_buf_2 fanout2161 (.A(net2162),
    .X(net2161));
 sg13g2_buf_4 fanout2162 (.X(net2162),
    .A(net2163));
 sg13g2_buf_4 fanout2163 (.X(net2163),
    .A(net2169));
 sg13g2_buf_2 fanout2164 (.A(net2165),
    .X(net2164));
 sg13g2_buf_2 fanout2165 (.A(net2166),
    .X(net2165));
 sg13g2_buf_2 fanout2166 (.A(net2169),
    .X(net2166));
 sg13g2_buf_2 fanout2167 (.A(net2169),
    .X(net2167));
 sg13g2_buf_1 fanout2168 (.A(net2169),
    .X(net2168));
 sg13g2_buf_2 fanout2169 (.A(\game_logic_inst.game_started ),
    .X(net2169));
 sg13g2_buf_2 fanout2170 (.A(net2172),
    .X(net2170));
 sg13g2_buf_1 fanout2171 (.A(net2172),
    .X(net2171));
 sg13g2_buf_2 fanout2172 (.A(\game_logic_inst.game_started ),
    .X(net2172));
 sg13g2_buf_2 fanout2173 (.A(net2175),
    .X(net2173));
 sg13g2_buf_2 fanout2174 (.A(net2175),
    .X(net2174));
 sg13g2_buf_2 fanout2175 (.A(\game_logic_inst.game_started ),
    .X(net2175));
 sg13g2_buf_4 fanout2176 (.X(net2176),
    .A(net965));
 sg13g2_buf_2 fanout2177 (.A(net2178),
    .X(net2177));
 sg13g2_buf_4 fanout2178 (.X(net2178),
    .A(\game_logic_inst.calculate_move ));
 sg13g2_buf_4 fanout2179 (.X(net2179),
    .A(net2181));
 sg13g2_buf_4 fanout2180 (.X(net2180),
    .A(net2181));
 sg13g2_buf_4 fanout2181 (.X(net2181),
    .A(net978));
 sg13g2_buf_4 fanout2182 (.X(net2182),
    .A(net2183));
 sg13g2_buf_8 fanout2183 (.A(_0090_),
    .X(net2183));
 sg13g2_buf_4 fanout2184 (.X(net2184),
    .A(\draw_game_inst.board_y[4] ));
 sg13g2_buf_4 fanout2185 (.X(net2185),
    .A(net2186));
 sg13g2_buf_4 fanout2186 (.X(net2186),
    .A(\draw_game_inst.board_y[4] ));
 sg13g2_buf_2 fanout2187 (.A(net2190),
    .X(net2187));
 sg13g2_buf_2 fanout2188 (.A(net2190),
    .X(net2188));
 sg13g2_buf_2 fanout2189 (.A(net2190),
    .X(net2189));
 sg13g2_buf_4 fanout2190 (.X(net2190),
    .A(\draw_game_inst.board_y[3] ));
 sg13g2_buf_4 fanout2191 (.X(net2191),
    .A(net2192));
 sg13g2_buf_4 fanout2192 (.X(net2192),
    .A(\draw_game_inst.board_y[3] ));
 sg13g2_buf_2 fanout2193 (.A(net2202),
    .X(net2193));
 sg13g2_buf_1 fanout2194 (.A(net2202),
    .X(net2194));
 sg13g2_buf_4 fanout2195 (.X(net2195),
    .A(net2198));
 sg13g2_buf_2 fanout2196 (.A(net2198),
    .X(net2196));
 sg13g2_buf_2 fanout2197 (.A(net2198),
    .X(net2197));
 sg13g2_buf_1 fanout2198 (.A(net2202),
    .X(net2198));
 sg13g2_buf_4 fanout2199 (.X(net2199),
    .A(net2202));
 sg13g2_buf_4 fanout2200 (.X(net2200),
    .A(net2201));
 sg13g2_buf_2 fanout2201 (.A(net2202),
    .X(net2201));
 sg13g2_buf_4 fanout2202 (.X(net2202),
    .A(\draw_game_inst.board_y[3] ));
 sg13g2_buf_4 fanout2203 (.X(net2203),
    .A(net2204));
 sg13g2_buf_4 fanout2204 (.X(net2204),
    .A(_0092_));
 sg13g2_buf_2 fanout2205 (.A(net2207),
    .X(net2205));
 sg13g2_buf_2 fanout2206 (.A(net2207),
    .X(net2206));
 sg13g2_buf_2 fanout2207 (.A(net2208),
    .X(net2207));
 sg13g2_buf_4 fanout2208 (.X(net2208),
    .A(net2220));
 sg13g2_buf_4 fanout2209 (.X(net2209),
    .A(net2220));
 sg13g2_buf_4 fanout2210 (.X(net2210),
    .A(net2213));
 sg13g2_buf_2 fanout2211 (.A(net2213),
    .X(net2211));
 sg13g2_buf_4 fanout2212 (.X(net2212),
    .A(net2213));
 sg13g2_buf_2 fanout2213 (.A(net2214),
    .X(net2213));
 sg13g2_buf_4 fanout2214 (.X(net2214),
    .A(net2219));
 sg13g2_buf_2 fanout2215 (.A(net2216),
    .X(net2215));
 sg13g2_buf_2 fanout2216 (.A(net2219),
    .X(net2216));
 sg13g2_buf_2 fanout2217 (.A(net2219),
    .X(net2217));
 sg13g2_buf_1 fanout2218 (.A(net2219),
    .X(net2218));
 sg13g2_buf_2 fanout2219 (.A(net2220),
    .X(net2219));
 sg13g2_buf_2 fanout2220 (.A(\draw_game_inst.board_y[2] ),
    .X(net2220));
 sg13g2_buf_4 fanout2221 (.X(net2221),
    .A(net2222));
 sg13g2_buf_4 fanout2222 (.X(net2222),
    .A(net2232));
 sg13g2_buf_2 fanout2223 (.A(net2226),
    .X(net2223));
 sg13g2_buf_2 fanout2224 (.A(net2226),
    .X(net2224));
 sg13g2_buf_2 fanout2225 (.A(net2226),
    .X(net2225));
 sg13g2_buf_1 fanout2226 (.A(net2232),
    .X(net2226));
 sg13g2_buf_4 fanout2227 (.X(net2227),
    .A(net2228));
 sg13g2_buf_2 fanout2228 (.A(net2232),
    .X(net2228));
 sg13g2_buf_2 fanout2229 (.A(net2231),
    .X(net2229));
 sg13g2_buf_1 fanout2230 (.A(net2231),
    .X(net2230));
 sg13g2_buf_4 fanout2231 (.X(net2231),
    .A(net2232));
 sg13g2_buf_4 fanout2232 (.X(net2232),
    .A(net2249));
 sg13g2_buf_2 fanout2233 (.A(net2234),
    .X(net2233));
 sg13g2_buf_2 fanout2234 (.A(net2235),
    .X(net2234));
 sg13g2_buf_2 fanout2235 (.A(net2249),
    .X(net2235));
 sg13g2_buf_4 fanout2236 (.X(net2236),
    .A(net2239));
 sg13g2_buf_2 fanout2237 (.A(net2239),
    .X(net2237));
 sg13g2_buf_2 fanout2238 (.A(net2239),
    .X(net2238));
 sg13g2_buf_2 fanout2239 (.A(net2249),
    .X(net2239));
 sg13g2_buf_2 fanout2240 (.A(net2241),
    .X(net2240));
 sg13g2_buf_2 fanout2241 (.A(net2242),
    .X(net2241));
 sg13g2_buf_2 fanout2242 (.A(net2248),
    .X(net2242));
 sg13g2_buf_2 fanout2243 (.A(net2245),
    .X(net2243));
 sg13g2_buf_1 fanout2244 (.A(net2245),
    .X(net2244));
 sg13g2_buf_2 fanout2245 (.A(net2248),
    .X(net2245));
 sg13g2_buf_4 fanout2246 (.X(net2246),
    .A(net2248));
 sg13g2_buf_2 fanout2247 (.A(net2248),
    .X(net2247));
 sg13g2_buf_1 fanout2248 (.A(net2249),
    .X(net2248));
 sg13g2_buf_4 fanout2249 (.X(net2249),
    .A(\draw_game_inst.board_y[1] ));
 sg13g2_buf_2 fanout2250 (.A(net2251),
    .X(net2250));
 sg13g2_buf_4 fanout2251 (.X(net2251),
    .A(net2252));
 sg13g2_buf_4 fanout2252 (.X(net2252),
    .A(_0169_));
 sg13g2_buf_4 fanout2253 (.X(net2253),
    .A(net2254));
 sg13g2_buf_2 fanout2254 (.A(net2255),
    .X(net2254));
 sg13g2_buf_4 fanout2255 (.X(net2255),
    .A(net2269));
 sg13g2_buf_4 fanout2256 (.X(net2256),
    .A(net2259));
 sg13g2_buf_2 fanout2257 (.A(net2259),
    .X(net2257));
 sg13g2_buf_2 fanout2258 (.A(net2259),
    .X(net2258));
 sg13g2_buf_2 fanout2259 (.A(net2269),
    .X(net2259));
 sg13g2_buf_4 fanout2260 (.X(net2260),
    .A(net2263));
 sg13g2_buf_4 fanout2261 (.X(net2261),
    .A(net2263));
 sg13g2_buf_2 fanout2262 (.A(net2263),
    .X(net2262));
 sg13g2_buf_2 fanout2263 (.A(net2269),
    .X(net2263));
 sg13g2_buf_4 fanout2264 (.X(net2264),
    .A(net2265));
 sg13g2_buf_2 fanout2265 (.A(net2268),
    .X(net2265));
 sg13g2_buf_4 fanout2266 (.X(net2266),
    .A(net2268));
 sg13g2_buf_4 fanout2267 (.X(net2267),
    .A(net2268));
 sg13g2_buf_2 fanout2268 (.A(net2269),
    .X(net2268));
 sg13g2_buf_4 fanout2269 (.X(net2269),
    .A(\draw_game_inst.board_y[0] ));
 sg13g2_buf_2 fanout2270 (.A(net1021),
    .X(net2270));
 sg13g2_buf_2 fanout2271 (.A(net2272),
    .X(net2271));
 sg13g2_buf_1 fanout2272 (.A(net902),
    .X(net2272));
 sg13g2_buf_2 fanout2273 (.A(net2274),
    .X(net2273));
 sg13g2_buf_1 fanout2274 (.A(net2275),
    .X(net2274));
 sg13g2_buf_2 fanout2275 (.A(net961),
    .X(net2275));
 sg13g2_buf_4 fanout2276 (.X(net2276),
    .A(net2279));
 sg13g2_buf_4 fanout2277 (.X(net2277),
    .A(net2278));
 sg13g2_buf_4 fanout2278 (.X(net2278),
    .A(net2279));
 sg13g2_buf_4 fanout2279 (.X(net2279),
    .A(\draw_game_inst.x[7] ));
 sg13g2_buf_4 fanout2280 (.X(net2280),
    .A(net2283));
 sg13g2_buf_4 fanout2281 (.X(net2281),
    .A(net2282));
 sg13g2_buf_4 fanout2282 (.X(net2282),
    .A(net2283));
 sg13g2_buf_2 fanout2283 (.A(\draw_game_inst.x[6] ),
    .X(net2283));
 sg13g2_buf_4 fanout2284 (.X(net2284),
    .A(net2285));
 sg13g2_buf_4 fanout2285 (.X(net2285),
    .A(_0094_));
 sg13g2_buf_4 fanout2286 (.X(net2286),
    .A(net1011));
 sg13g2_buf_4 fanout2287 (.X(net2287),
    .A(net2288));
 sg13g2_buf_4 fanout2288 (.X(net2288),
    .A(net2289));
 sg13g2_buf_4 fanout2289 (.X(net2289),
    .A(\draw_game_inst.board_x[5] ));
 sg13g2_buf_4 fanout2290 (.X(net2290),
    .A(net2291));
 sg13g2_buf_2 fanout2291 (.A(\draw_game_inst.board_x[4] ),
    .X(net2291));
 sg13g2_buf_4 fanout2292 (.X(net2292),
    .A(net2294));
 sg13g2_buf_2 fanout2293 (.A(net2294),
    .X(net2293));
 sg13g2_buf_4 fanout2294 (.X(net2294),
    .A(\draw_game_inst.board_x[4] ));
 sg13g2_buf_4 fanout2295 (.X(net2295),
    .A(_0095_));
 sg13g2_buf_4 fanout2296 (.X(net2296),
    .A(net2300));
 sg13g2_buf_4 fanout2297 (.X(net2297),
    .A(net2299));
 sg13g2_buf_2 fanout2298 (.A(net2299),
    .X(net2298));
 sg13g2_buf_2 fanout2299 (.A(net2300),
    .X(net2299));
 sg13g2_buf_2 fanout2300 (.A(\draw_game_inst.board_x[3] ),
    .X(net2300));
 sg13g2_buf_4 fanout2301 (.X(net2301),
    .A(net2302));
 sg13g2_buf_4 fanout2302 (.X(net2302),
    .A(net2307));
 sg13g2_buf_2 fanout2303 (.A(net2304),
    .X(net2303));
 sg13g2_buf_2 fanout2304 (.A(net2305),
    .X(net2304));
 sg13g2_buf_4 fanout2305 (.X(net2305),
    .A(net2306));
 sg13g2_buf_4 fanout2306 (.X(net2306),
    .A(net2307));
 sg13g2_buf_4 fanout2307 (.X(net2307),
    .A(_4024_));
 sg13g2_buf_2 fanout2308 (.A(net2309),
    .X(net2308));
 sg13g2_buf_2 fanout2309 (.A(net2310),
    .X(net2309));
 sg13g2_buf_2 fanout2310 (.A(net2311),
    .X(net2310));
 sg13g2_buf_4 fanout2311 (.X(net2311),
    .A(net2337));
 sg13g2_buf_2 fanout2312 (.A(net2313),
    .X(net2312));
 sg13g2_buf_1 fanout2313 (.A(net2315),
    .X(net2313));
 sg13g2_buf_2 fanout2314 (.A(net2315),
    .X(net2314));
 sg13g2_buf_1 fanout2315 (.A(net2316),
    .X(net2315));
 sg13g2_buf_4 fanout2316 (.X(net2316),
    .A(net2337));
 sg13g2_buf_2 fanout2317 (.A(net2319),
    .X(net2317));
 sg13g2_buf_1 fanout2318 (.A(net2319),
    .X(net2318));
 sg13g2_buf_2 fanout2319 (.A(net2324),
    .X(net2319));
 sg13g2_buf_2 fanout2320 (.A(net2321),
    .X(net2320));
 sg13g2_buf_2 fanout2321 (.A(net2324),
    .X(net2321));
 sg13g2_buf_2 fanout2322 (.A(net2323),
    .X(net2322));
 sg13g2_buf_4 fanout2323 (.X(net2323),
    .A(net2324));
 sg13g2_buf_2 fanout2324 (.A(net2337),
    .X(net2324));
 sg13g2_buf_2 fanout2325 (.A(net2332),
    .X(net2325));
 sg13g2_buf_2 fanout2326 (.A(net2332),
    .X(net2326));
 sg13g2_buf_2 fanout2327 (.A(net2330),
    .X(net2327));
 sg13g2_buf_2 fanout2328 (.A(net2330),
    .X(net2328));
 sg13g2_buf_2 fanout2329 (.A(net2330),
    .X(net2329));
 sg13g2_buf_2 fanout2330 (.A(net2332),
    .X(net2330));
 sg13g2_buf_4 fanout2331 (.X(net2331),
    .A(net2332));
 sg13g2_buf_2 fanout2332 (.A(net2336),
    .X(net2332));
 sg13g2_buf_4 fanout2333 (.X(net2333),
    .A(net2334));
 sg13g2_buf_1 fanout2334 (.A(net2336),
    .X(net2334));
 sg13g2_buf_2 fanout2335 (.A(net2336),
    .X(net2335));
 sg13g2_buf_2 fanout2336 (.A(net2337),
    .X(net2336));
 sg13g2_buf_2 fanout2337 (.A(rst_n),
    .X(net2337));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_2 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_tielo tt_um_2048_vga_game_17 (.L_LO(net17));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_4_15_0_clk));
 sg13g2_inv_4 clkload2 (.A(clknet_leaf_3_clk));
 sg13g2_inv_4 clkload3 (.A(clknet_leaf_60_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_61_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_4_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_57_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_6_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_11_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_20_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_16_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_17_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_10_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_25_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_23_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_42_clk));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_39_clk));
 sg13g2_inv_8 clkload18 (.A(clknet_leaf_30_clk));
 sg13g2_inv_8 clkload19 (.A(clknet_leaf_45_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_49_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_8_clk));
 sg13g2_inv_4 clkload22 (.A(clknet_leaf_28_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_31_clk));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_7_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\gamepad_pmod.driver.pmod_latch_sync[1] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold2 (.A(\gamepad_pmod.driver.pmod_clk_sync[1] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0077_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0266_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0079_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0268_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0080_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0269_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0070_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0071_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0260_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0078_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0267_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0073_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0262_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0076_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0265_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0084_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0273_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0081_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0270_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0072_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0261_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0174_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0172_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0171_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0170_),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0173_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0168_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0085_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold31 (.A(\lfsr_inst.lfsr[26] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold32 (.A(\lfsr_inst.lfsr[16] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold33 (.A(\lfsr_inst.lfsr[25] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold34 (.A(\lfsr_inst.lfsr[19] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold35 (.A(\lfsr_inst.lfsr[27] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0087_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0277_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold38 (.A(\lfsr_inst.lfsr[24] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold39 (.A(\lfsr_inst.lfsr[17] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold40 (.A(\lfsr_inst.lfsr[23] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold41 (.A(\draw_game_inst.new_tiles[0] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold42 (.A(\lfsr_inst.lfsr[18] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0082_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold44 (.A(\btn_down_debounce.button_sync_1 ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold45 (.A(_3616_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0320_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold47 (.A(\game_logic_inst.lfsr_value[3] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0083_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold49 (.A(\game_logic_inst.lfsr_value[9] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0167_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0279_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold52 (.A(\gamepad_pmod.driver.shift_reg[9] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0374_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold54 (.A(\gamepad_pmod.driver.shift_reg[1] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0366_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold56 (.A(\lfsr_inst.lfsr[22] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold57 (.A(\lfsr_inst.lfsr[20] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold58 (.A(\lfsr_inst.lfsr[21] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0075_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold60 (.A(_3505_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold61 (.A(\game_logic_inst.lfsr_value[13] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold62 (.A(\game_logic_inst.lfsr_value[15] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold63 (.A(\game_logic_inst.lfsr_value[8] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0086_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0275_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0074_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold67 (.A(\game_logic_inst.lfsr_value[11] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold68 (.A(\game_logic_inst.lfsr_value[5] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold69 (.A(\btn_down_debounce.debounce_counter[17] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold70 (.A(_3614_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0319_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold72 (.A(\btn_up_debounce.debounce_counter[2] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold73 (.A(_3544_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0283_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold75 (.A(\gamepad_pmod.decoder.data_reg[1] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0425_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold77 (.A(\btn_right_debounce.debounce_counter[2] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold78 (.A(_3671_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0345_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold80 (.A(\game_logic_inst.lfsr_value[6] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold81 (.A(\btn_down_debounce.debounce_counter[0] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold82 (.A(_3575_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0303_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold84 (.A(\game_logic_inst.lfsr_value[12] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold85 (.A(\btn_right_debounce.debounce_counter[17] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0360_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold87 (.A(\btn_left_debounce.button_sync_1 ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold88 (.A(_3658_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0341_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold90 (.A(\game_logic_inst.lfsr_value[4] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold91 (.A(\gamepad_pmod.decoder.data_reg[2] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0426_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold93 (.A(\gamepad_pmod.decoder.data_reg[11] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0435_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold95 (.A(\gamepad_pmod.decoder.data_reg[0] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0424_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold97 (.A(\gamepad_pmod.driver.pmod_data_sync[1] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0364_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold99 (.A(\btn_down_debounce.debounce_counter[16] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0318_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold101 (.A(\game_logic_inst.lfsr_value[7] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold102 (.A(\game_logic_inst.lfsr_value[1] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold103 (.A(\gamepad_pmod.decoder.data_reg[3] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0427_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold105 (.A(\btn_left_debounce.debounce_counter[10] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold106 (.A(_3643_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold107 (.A(\btn_right_debounce.debounce_counter[10] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold108 (.A(_3685_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0353_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold110 (.A(\btn_down_debounce.debounce_counter[12] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold111 (.A(_3605_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0314_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold113 (.A(\btn_right_debounce.debounce_counter[16] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold114 (.A(_3695_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0359_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold116 (.A(\btn_left_debounce.debounce_counter[2] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold117 (.A(_3629_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0324_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold119 (.A(\gamepad_pmod.decoder.data_reg[10] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0434_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold121 (.A(\btn_left_debounce.debounce_counter[12] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold122 (.A(_3646_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0334_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold124 (.A(\game_logic_inst.lfsr_value[2] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold125 (.A(\gamepad_pmod.driver.shift_reg[11] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0375_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold127 (.A(\game_logic_inst.lfsr_value[10] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold128 (.A(\vga_sync_gen.vsync ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold129 (.A(\btn_up_debounce.debounce_counter[10] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold130 (.A(_3558_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0291_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold132 (.A(\btn_down_debounce.debounce_counter[10] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold133 (.A(_3602_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0312_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold135 (.A(\gamepad_pmod.decoder.data_reg[7] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0431_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold137 (.A(\btn_up_debounce.debounce_counter[17] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold138 (.A(_3571_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0298_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold140 (.A(\game_logic_inst.current_direction[1] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0000_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold142 (.A(\gamepad_pmod.decoder.data_reg[6] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0430_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold144 (.A(\gamepad_pmod.decoder.data_reg[9] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold145 (.A(\gamepad_pmod.decoder.data_reg[4] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0428_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold147 (.A(\btn_up_debounce.debounce_counter[12] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold148 (.A(_3561_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0293_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold150 (.A(\btn_down_debounce.debounce_counter[4] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold151 (.A(_3592_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0097_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold153 (.A(_3845_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0464_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold155 (.A(\btn_right_debounce.debounce_counter[4] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold156 (.A(_3675_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold157 (.A(\btn_left_debounce.debounce_counter[4] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold158 (.A(_3633_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold159 (.A(\btn_right_debounce.debounce_counter[12] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold160 (.A(_3688_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0355_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold162 (.A(\game_logic_inst.lfsr_value[14] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold163 (.A(\new_tiles_counter[4] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0278_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold165 (.A(\btn_down_debounce.debounce_counter[3] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold166 (.A(_3590_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0098_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold168 (.A(_3859_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold169 (.A(\btn_right_debounce.debounce_counter[15] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0358_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold171 (.A(\gamepad_pmod.driver.shift_reg[0] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0365_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold173 (.A(\btn_left_debounce.debounce_counter[17] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold174 (.A(_3656_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0339_),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold176 (.A(\gamepad_pmod.driver.shift_reg[8] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0372_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold178 (.A(\welcome_screen_grid[28] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold179 (.A(_3773_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold180 (.A(\gamepad_pmod.driver.shift_reg[7] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0371_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold182 (.A(\btn_up_debounce.debounce_counter[7] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold183 (.A(_3553_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0288_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold185 (.A(\btn_right_debounce.debounce_counter[8] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold186 (.A(_3682_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold187 (.A(\gamepad_pmod.decoder.data_reg[5] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0429_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold189 (.A(\btn_down_debounce.debounce_counter[5] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold190 (.A(\gamepad_pmod.driver.shift_reg[3] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0367_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold192 (.A(\gamepad_pmod.driver.shift_reg[6] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0370_),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold194 (.A(\btn_up_debounce.debounce_counter[14] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold195 (.A(_3565_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold196 (.A(\btn_right_debounce.debounce_counter[7] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold197 (.A(_3680_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold198 (.A(\welcome_screen_grid[56] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold199 (.A(\gamepad_pmod.driver.shift_reg[5] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0369_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold201 (.A(\btn_up_debounce.debounced ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0300_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold203 (.A(\btn_up_debounce.debounce_counter[15] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold204 (.A(\btn_up_debounce.debounce_counter[5] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold205 (.A(_3550_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold206 (.A(\welcome_screen_grid[48] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold207 (.A(_3780_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold208 (.A(\btn_up_debounce.debounce_counter[16] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold209 (.A(\btn_up_debounce.debounce_counter[4] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold210 (.A(_3548_),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold211 (.A(\btn_left_debounce.debounce_counter[5] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold212 (.A(\welcome_screen_inst.welcome_counter[1] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0453_),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold214 (.A(\btn_right_debounce.debounce_counter[5] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold215 (.A(\btn_left_debounce.debounce_counter[15] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold216 (.A(_3652_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold217 (.A(\btn_right_debounce.debounce_counter[13] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold218 (.A(_3690_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold219 (.A(\gamepad_pmod.driver.pmod_clk_prev ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold220 (.A(\btn_left_debounce.debounce_counter[6] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold221 (.A(\welcome_screen_grid[52] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold222 (.A(\draw_game_inst.grid[60] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0252_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold224 (.A(\btn_left_debounce.debounce_counter[3] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold225 (.A(_3631_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold226 (.A(\btn_up_debounce.debounce_counter[6] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold227 (.A(\welcome_screen_grid[4] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold228 (.A(\btn_up_debounce.debounce_counter[13] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold229 (.A(_3563_),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold230 (.A(\btn_right_debounce.debounced ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0362_),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold232 (.A(\welcome_screen_grid[44] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold233 (.A(_3779_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold234 (.A(\btn_up_debounce.debounce_counter[3] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold235 (.A(_3546_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold236 (.A(\draw_game_inst.grid[51] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0243_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold238 (.A(\draw_game_inst.grid[3] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0195_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold240 (.A(\gamepad_pmod.driver.shift_reg[4] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold241 (.A(\welcome_screen_grid[16] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold242 (.A(_3767_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold243 (.A(\btn_left_debounce.debounce_counter[7] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold244 (.A(\btn_left_debounce.debounce_counter[13] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold245 (.A(_3648_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold246 (.A(\draw_game_inst.grid[11] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0203_),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold248 (.A(\btn_down_debounce.debounce_counter[7] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold249 (.A(_3597_),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold250 (.A(\btn_down_debounce.debounce_counter[13] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold251 (.A(\btn_right_debounce.debounce_counter[6] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold252 (.A(\btn_down_debounce.debounce_counter[2] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold253 (.A(_3588_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold254 (.A(\draw_game_inst.grid[15] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0207_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold256 (.A(\btn_left_debounce.debounce_counter[14] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold257 (.A(\btn_right_debounce.debounce_counter[3] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold258 (.A(_3673_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold259 (.A(\draw_game_inst.grid[42] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0234_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold261 (.A(\welcome_screen_inst.welcome_counter[2] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold262 (.A(\draw_game_inst.grid[57] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0249_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold264 (.A(\btn_down_debounce.debounce_counter[8] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold265 (.A(\draw_game_inst.grid[53] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0245_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold267 (.A(\gamepad_pmod.decoder.data_reg[8] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold268 (.A(\draw_game_inst.grid[22] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0214_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold270 (.A(\draw_game_inst.grid[19] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0211_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold272 (.A(\btn_left_debounce.debounce_counter[8] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold273 (.A(\draw_game_inst.grid[48] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0240_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold275 (.A(\debug_controller_inst.grid_out_addr[1] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0487_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold277 (.A(\draw_game_inst.grid[31] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0223_),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold279 (.A(\draw_game_inst.grid[4] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0196_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold281 (.A(\draw_game_inst.grid[46] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0238_),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold283 (.A(\btn_left_debounce.debounce_counter[16] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold284 (.A(\draw_game_inst.grid[28] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0220_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold286 (.A(\draw_game_inst.grid[24] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0216_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold288 (.A(\draw_game_inst.grid[0] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0192_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold290 (.A(\draw_game_inst.grid[6] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0198_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold292 (.A(\draw_game_inst.grid[7] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0199_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold294 (.A(\draw_game_inst.grid[34] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0226_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold296 (.A(\welcome_screen_grid[60] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold297 (.A(_3783_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold298 (.A(\btn_up_debounce.debounce_counter[0] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold299 (.A(_3542_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold300 (.A(\draw_game_inst.grid[63] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0255_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold302 (.A(\draw_game_inst.grid[56] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0248_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold304 (.A(\draw_game_inst.grid[26] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0218_),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold306 (.A(\draw_game_inst.grid[14] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0206_),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold308 (.A(\draw_game_inst.grid[61] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0253_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold310 (.A(\debug_controller_inst.grid_out_addr[0] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0486_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold312 (.A(\draw_game_inst.grid[2] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0194_),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold314 (.A(\draw_game_inst.grid[39] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0231_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold316 (.A(\draw_game_inst.grid[59] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0251_),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold318 (.A(\welcome_screen_grid[36] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold319 (.A(\draw_game_inst.grid[18] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0210_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold321 (.A(\welcome_screen_inst.welcome_counter[4] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold322 (.A(_3797_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0456_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold324 (.A(\welcome_screen_grid[24] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold325 (.A(\draw_game_inst.grid[62] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0254_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold327 (.A(\welcome_screen_grid[32] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0444_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold329 (.A(\draw_game_inst.grid[35] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0227_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold331 (.A(\draw_game_inst.grid[1] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0193_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold333 (.A(\draw_game_inst.grid[12] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0204_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold335 (.A(\draw_game_inst.grid[27] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0219_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold337 (.A(\draw_game_inst.grid[36] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0228_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold339 (.A(\draw_game_inst.grid[52] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0244_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold341 (.A(\draw_game_inst.grid[58] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0250_),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold343 (.A(\welcome_screen_grid[40] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold344 (.A(\draw_game_inst.grid[20] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0212_),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold346 (.A(\draw_game_inst.grid[33] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold347 (.A(\draw_game_inst.grid[17] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0209_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold349 (.A(\draw_game_inst.grid[47] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0239_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold351 (.A(\draw_game_inst.grid[8] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold352 (.A(\btn_left_debounce.debounce_counter[11] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold353 (.A(\draw_game_inst.grid[29] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0221_),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0089_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold356 (.A(_3724_),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0419_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold358 (.A(\draw_game_inst.grid[55] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0247_),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold360 (.A(\draw_game_inst.grid[21] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0213_),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold362 (.A(\draw_game_inst.grid[37] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0229_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold364 (.A(\draw_game_inst.grid[25] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0217_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold366 (.A(\draw_game_inst.grid[5] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0197_),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold368 (.A(\draw_game_inst.grid[50] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0242_),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold370 (.A(\draw_game_inst.grid[23] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0215_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold372 (.A(\btn_down_debounce.debounce_counter[6] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold373 (.A(\btn_up_debounce.debounce_counter[8] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold374 (.A(\welcome_screen_grid[11] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold375 (.A(\game_logic_inst.lfsr_value[0] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold376 (.A(\welcome_screen_inst.welcome_counter[3] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold377 (.A(_3795_),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold378 (.A(\draw_game_inst.grid[44] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0236_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold380 (.A(\draw_game_inst.grid[16] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0208_),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold382 (.A(\gamepad_pmod.driver.pmod_clk_sync[0] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold383 (.A(\draw_game_inst.grid[40] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0232_),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold385 (.A(\btn_up_debounce.debounce_counter[11] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold386 (.A(_3560_),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0292_),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold388 (.A(\btn_left_debounce.debounce_counter[9] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold389 (.A(\gamepad_pmod.driver.pmod_data_sync[0] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold390 (.A(\draw_game_inst.grid[41] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0233_),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold392 (.A(\btn_down_debounce.debounce_counter[9] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold393 (.A(\draw_game_inst.grid[45] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0237_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0132_),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold396 (.A(\btn_down_debounce.debounce_counter[11] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold397 (.A(\welcome_screen_grid[12] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold398 (.A(_3764_),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold399 (.A(\draw_game_inst.grid[13] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0205_),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold401 (.A(\debug_controller_inst.grid_out_addr[2] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0488_),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold403 (.A(\draw_game_inst.grid[54] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0246_),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold405 (.A(\btn_right_debounce.debounce_counter[9] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold406 (.A(\draw_game_inst.grid[43] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0235_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold408 (.A(\welcome_screen_grid[20] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold409 (.A(\draw_game_inst.grid[32] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0224_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold411 (.A(\draw_game_inst.grid[49] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0241_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold413 (.A(\btn_left_debounce.debounce_counter[1] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold414 (.A(_3627_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold415 (.A(uio_out[6]),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold416 (.A(\draw_game_inst.grid[30] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0222_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold418 (.A(\btn_down_debounce.debounce_counter[14] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold419 (.A(\draw_game_inst.grid[38] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0230_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold421 (.A(\btn_right_debounce.debounce_counter[14] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold422 (.A(\welcome_screen_grid[0] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0436_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold424 (.A(\btn_right_debounce.debounce_counter[1] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold425 (.A(_3669_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold426 (.A(\btn_right_debounce.debounce_counter[11] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0354_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold428 (.A(\btn_up_debounce.debounce_counter[9] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold429 (.A(debug_btn_up),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0500_),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold431 (.A(_0514_),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold432 (.A(\btn_down_debounce.debounce_counter[15] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold433 (.A(\gamepad_pmod.driver.pmod_latch_sync[0] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold434 (.A(\game_logic_inst.debug_move_reg ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0457_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0166_),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold437 (.A(\draw_game_inst.grid[10] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold438 (.A(\draw_game_inst.grid[9] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0201_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold440 (.A(uio_out[4]),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold441 (.A(\game_logic_inst.should_transpose ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold442 (.A(_0470_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold443 (.A(\draw_game_inst.y[8] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold444 (.A(_3728_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold445 (.A(_0421_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0151_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold447 (.A(_1270_),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold448 (.A(\game_logic_inst.current_direction[2] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold449 (.A(_0001_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0109_),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold451 (.A(_0924_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0155_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold453 (.A(_0157_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold454 (.A(_1292_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold455 (.A(_0101_),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0161_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold457 (.A(_0149_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0100_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold459 (.A(\draw_game_inst.y[8] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0148_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0152_),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold462 (.A(_1368_),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0103_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0872_),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold465 (.A(_0119_),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0986_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold467 (.A(\lfsr_inst.lfsr[31] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0138_),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold469 (.A(_1228_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold470 (.A(_0125_),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold471 (.A(_1015_),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0131_),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold473 (.A(_1101_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold474 (.A(_0159_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold475 (.A(uio_out[7]),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0156_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold477 (.A(_1383_),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0163_),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold479 (.A(_3962_),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0147_),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold481 (.A(\game_logic_inst.add_new_tiles[0] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0117_),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0971_),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0005_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold485 (.A(_0105_),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold486 (.A(_0892_),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold487 (.A(\lfsr_inst.lfsr[28] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold488 (.A(_0129_),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold489 (.A(_0017_),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold490 (.A(_0102_),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold491 (.A(_0808_),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold492 (.A(_0036_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0150_),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold494 (.A(_0040_),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold495 (.A(\draw_game_inst.board_y[6] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold496 (.A(_0154_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold497 (.A(_1376_),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0127_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0153_),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold500 (.A(_1278_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold501 (.A(\lfsr_inst.lfsr[30] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold502 (.A(_0158_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold503 (.A(_1390_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold504 (.A(uio_out[5]),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold505 (.A(\draw_game_inst.x[9] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold506 (.A(_0067_),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold507 (.A(_0134_),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold508 (.A(_1214_),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold509 (.A(_0121_),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold510 (.A(_0997_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold511 (.A(_0140_),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold512 (.A(_0136_),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold513 (.A(_1221_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold514 (.A(_0111_),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold515 (.A(_0939_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0135_),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold517 (.A(_1118_),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold518 (.A(_0123_),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold519 (.A(_1005_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold520 (.A(_0115_),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold521 (.A(_0961_),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold522 (.A(\debug_controller_inst.grid_out_data[0] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0160_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold524 (.A(\draw_game_inst.board_x[2] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold525 (.A(_0142_),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold526 (.A(_1343_),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold527 (.A(_0099_),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold528 (.A(\btn_down_debounce.button_sync_0 ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold529 (.A(\btn_left_debounce.button_sync_0 ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold530 (.A(_0133_),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold531 (.A(_1110_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold532 (.A(_0107_),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0910_),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold534 (.A(_0146_),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold535 (.A(_1358_),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold536 (.A(_0053_),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0112_),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold538 (.A(_0028_),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold539 (.A(\game_logic_inst.valid_move ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold540 (.A(\debug_controller_inst.grid_addr[3] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold541 (.A(_0494_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold542 (.A(_0113_),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold543 (.A(_0951_),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0143_),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold545 (.A(_1153_),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold546 (.A(show_welcome_screen),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold547 (.A(_3488_),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0137_),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold549 (.A(_0022_),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold550 (.A(\game_logic_inst.calculate_move ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold551 (.A(_3830_),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold552 (.A(\game_logic_inst.lfsr_shift[1] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold553 (.A(_3831_),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold554 (.A(_0162_),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold555 (.A(_1424_),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold556 (.A(_0062_),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold557 (.A(\draw_game_inst.x[8] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold558 (.A(_0130_),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold559 (.A(_1089_),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold560 (.A(_0018_),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold561 (.A(_0128_),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold562 (.A(\btn_right_debounce.button_sync_0 ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold563 (.A(\draw_game_inst.board_y[5] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold564 (.A(_0417_),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold565 (.A(_0144_),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold566 (.A(_0052_),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold567 (.A(\draw_game_inst.new_tiles_counter[1] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold568 (.A(\game_logic_inst.current_row_index[1] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold569 (.A(\draw_game_inst.x[9] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold570 (.A(_1473_),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold571 (.A(\debug_controller_inst.grid_out_data[1] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold572 (.A(\draw_game_inst.board_x[1] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold573 (.A(\debug_controller_inst.grid_out_addr[3] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold574 (.A(\debug_controller_inst.grid_out_data[2] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold575 (.A(\btn_up_debounce.button_sync_0 ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold576 (.A(_0106_),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold577 (.A(_1037_),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold578 (.A(_0108_),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold579 (.A(\draw_game_inst.y[9] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold580 (.A(\debug_controller_inst.grid_out_data[3] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold581 (.A(_0031_),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold582 (.A(\welcome_screen_inst.welcome_counter[0] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold583 (.A(\debug_controller_inst.grid_addr[2] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold584 (.A(_0145_),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold585 (.A(_1161_),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold586 (.A(_0126_),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold587 (.A(_0120_),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold588 (.A(_0045_),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold589 (.A(_0104_),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold590 (.A(_1029_),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold591 (.A(_0109_),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold592 (.A(_1048_),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold593 (.A(_1051_),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold594 (.A(\draw_game_inst.new_tiles_counter[2] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold595 (.A(_0188_),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold596 (.A(\draw_game_inst.board_x[5] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold597 (.A(_0122_),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold598 (.A(_1310_),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold599 (.A(_0116_),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold600 (.A(_1186_),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold601 (.A(_0114_),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold602 (.A(_1180_),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold603 (.A(_0141_),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold604 (.A(_1145_),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold605 (.A(\debug_controller_inst.grid_addr[0] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold606 (.A(\lfsr_inst.lfsr[29] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold607 (.A(_0139_),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold608 (.A(_1137_),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold609 (.A(_0124_),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold610 (.A(debug_btn_left),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold611 (.A(_0156_),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold612 (.A(\debug_controller_inst.grid_out_data[0] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold613 (.A(\btn_down_debounce.debounce_counter[11] ),
    .X(net1028));
 sg13g2_antennanp ANTENNA_1 (.A(_0468_));
 sg13g2_antennanp ANTENNA_2 (.A(_0468_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_fill_2 FILLER_8_532 ();
 sg13g2_fill_1 FILLER_8_534 ();
 sg13g2_fill_2 FILLER_8_547 ();
 sg13g2_fill_1 FILLER_8_549 ();
 sg13g2_decap_8 FILLER_8_554 ();
 sg13g2_decap_8 FILLER_8_561 ();
 sg13g2_decap_8 FILLER_8_568 ();
 sg13g2_decap_8 FILLER_8_575 ();
 sg13g2_decap_8 FILLER_8_582 ();
 sg13g2_decap_8 FILLER_8_589 ();
 sg13g2_decap_8 FILLER_8_596 ();
 sg13g2_decap_8 FILLER_8_603 ();
 sg13g2_decap_8 FILLER_8_610 ();
 sg13g2_decap_8 FILLER_8_617 ();
 sg13g2_decap_8 FILLER_8_624 ();
 sg13g2_decap_8 FILLER_8_631 ();
 sg13g2_decap_8 FILLER_8_638 ();
 sg13g2_decap_8 FILLER_8_645 ();
 sg13g2_decap_8 FILLER_8_652 ();
 sg13g2_decap_8 FILLER_8_659 ();
 sg13g2_decap_8 FILLER_8_666 ();
 sg13g2_decap_8 FILLER_8_673 ();
 sg13g2_decap_8 FILLER_8_680 ();
 sg13g2_decap_8 FILLER_8_687 ();
 sg13g2_decap_8 FILLER_8_694 ();
 sg13g2_decap_8 FILLER_8_701 ();
 sg13g2_decap_8 FILLER_8_708 ();
 sg13g2_decap_8 FILLER_8_715 ();
 sg13g2_decap_8 FILLER_8_722 ();
 sg13g2_decap_8 FILLER_8_729 ();
 sg13g2_decap_8 FILLER_8_736 ();
 sg13g2_decap_8 FILLER_8_743 ();
 sg13g2_decap_8 FILLER_8_750 ();
 sg13g2_decap_8 FILLER_8_757 ();
 sg13g2_decap_8 FILLER_8_764 ();
 sg13g2_decap_8 FILLER_8_771 ();
 sg13g2_decap_8 FILLER_8_778 ();
 sg13g2_decap_8 FILLER_8_785 ();
 sg13g2_decap_8 FILLER_8_792 ();
 sg13g2_decap_8 FILLER_8_799 ();
 sg13g2_decap_8 FILLER_8_806 ();
 sg13g2_decap_8 FILLER_8_813 ();
 sg13g2_decap_8 FILLER_8_820 ();
 sg13g2_decap_8 FILLER_8_827 ();
 sg13g2_decap_8 FILLER_8_834 ();
 sg13g2_decap_8 FILLER_8_841 ();
 sg13g2_decap_8 FILLER_8_848 ();
 sg13g2_decap_8 FILLER_8_855 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_fill_2 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_4 FILLER_9_476 ();
 sg13g2_fill_2 FILLER_9_489 ();
 sg13g2_fill_1 FILLER_9_491 ();
 sg13g2_fill_2 FILLER_9_510 ();
 sg13g2_fill_2 FILLER_9_542 ();
 sg13g2_decap_8 FILLER_9_562 ();
 sg13g2_decap_8 FILLER_9_569 ();
 sg13g2_decap_8 FILLER_9_576 ();
 sg13g2_decap_8 FILLER_9_583 ();
 sg13g2_decap_8 FILLER_9_590 ();
 sg13g2_decap_8 FILLER_9_597 ();
 sg13g2_decap_8 FILLER_9_604 ();
 sg13g2_decap_8 FILLER_9_611 ();
 sg13g2_decap_8 FILLER_9_618 ();
 sg13g2_decap_8 FILLER_9_625 ();
 sg13g2_decap_8 FILLER_9_632 ();
 sg13g2_decap_8 FILLER_9_639 ();
 sg13g2_decap_8 FILLER_9_646 ();
 sg13g2_decap_8 FILLER_9_653 ();
 sg13g2_decap_8 FILLER_9_660 ();
 sg13g2_decap_8 FILLER_9_667 ();
 sg13g2_decap_8 FILLER_9_674 ();
 sg13g2_decap_8 FILLER_9_681 ();
 sg13g2_decap_8 FILLER_9_688 ();
 sg13g2_decap_8 FILLER_9_695 ();
 sg13g2_decap_8 FILLER_9_702 ();
 sg13g2_decap_8 FILLER_9_709 ();
 sg13g2_decap_8 FILLER_9_716 ();
 sg13g2_decap_8 FILLER_9_723 ();
 sg13g2_decap_8 FILLER_9_730 ();
 sg13g2_decap_8 FILLER_9_737 ();
 sg13g2_decap_8 FILLER_9_744 ();
 sg13g2_decap_8 FILLER_9_751 ();
 sg13g2_decap_8 FILLER_9_758 ();
 sg13g2_decap_8 FILLER_9_765 ();
 sg13g2_decap_8 FILLER_9_772 ();
 sg13g2_decap_8 FILLER_9_779 ();
 sg13g2_decap_8 FILLER_9_786 ();
 sg13g2_decap_8 FILLER_9_793 ();
 sg13g2_decap_8 FILLER_9_800 ();
 sg13g2_decap_8 FILLER_9_807 ();
 sg13g2_decap_8 FILLER_9_814 ();
 sg13g2_decap_8 FILLER_9_821 ();
 sg13g2_decap_8 FILLER_9_828 ();
 sg13g2_decap_8 FILLER_9_835 ();
 sg13g2_decap_8 FILLER_9_842 ();
 sg13g2_decap_8 FILLER_9_849 ();
 sg13g2_decap_4 FILLER_9_856 ();
 sg13g2_fill_2 FILLER_9_860 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_102 ();
 sg13g2_decap_4 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_118 ();
 sg13g2_fill_2 FILLER_10_177 ();
 sg13g2_fill_1 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_198 ();
 sg13g2_decap_4 FILLER_10_205 ();
 sg13g2_decap_8 FILLER_10_223 ();
 sg13g2_decap_8 FILLER_10_230 ();
 sg13g2_decap_8 FILLER_10_237 ();
 sg13g2_decap_8 FILLER_10_244 ();
 sg13g2_decap_8 FILLER_10_251 ();
 sg13g2_decap_8 FILLER_10_258 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_fill_2 FILLER_10_462 ();
 sg13g2_fill_1 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_573 ();
 sg13g2_decap_8 FILLER_10_580 ();
 sg13g2_decap_8 FILLER_10_587 ();
 sg13g2_decap_8 FILLER_10_594 ();
 sg13g2_decap_8 FILLER_10_601 ();
 sg13g2_decap_8 FILLER_10_608 ();
 sg13g2_decap_8 FILLER_10_615 ();
 sg13g2_decap_8 FILLER_10_622 ();
 sg13g2_decap_8 FILLER_10_629 ();
 sg13g2_decap_8 FILLER_10_636 ();
 sg13g2_decap_8 FILLER_10_643 ();
 sg13g2_decap_8 FILLER_10_650 ();
 sg13g2_decap_8 FILLER_10_657 ();
 sg13g2_decap_8 FILLER_10_664 ();
 sg13g2_decap_8 FILLER_10_671 ();
 sg13g2_decap_8 FILLER_10_678 ();
 sg13g2_decap_8 FILLER_10_685 ();
 sg13g2_decap_8 FILLER_10_692 ();
 sg13g2_decap_8 FILLER_10_699 ();
 sg13g2_decap_8 FILLER_10_706 ();
 sg13g2_decap_8 FILLER_10_713 ();
 sg13g2_decap_8 FILLER_10_720 ();
 sg13g2_decap_8 FILLER_10_727 ();
 sg13g2_decap_8 FILLER_10_734 ();
 sg13g2_decap_8 FILLER_10_741 ();
 sg13g2_decap_8 FILLER_10_748 ();
 sg13g2_decap_8 FILLER_10_755 ();
 sg13g2_decap_8 FILLER_10_762 ();
 sg13g2_decap_8 FILLER_10_769 ();
 sg13g2_decap_8 FILLER_10_776 ();
 sg13g2_decap_8 FILLER_10_783 ();
 sg13g2_decap_8 FILLER_10_790 ();
 sg13g2_decap_8 FILLER_10_797 ();
 sg13g2_decap_8 FILLER_10_804 ();
 sg13g2_decap_8 FILLER_10_811 ();
 sg13g2_decap_8 FILLER_10_818 ();
 sg13g2_decap_8 FILLER_10_825 ();
 sg13g2_decap_8 FILLER_10_832 ();
 sg13g2_decap_8 FILLER_10_839 ();
 sg13g2_decap_8 FILLER_10_846 ();
 sg13g2_decap_8 FILLER_10_853 ();
 sg13g2_fill_2 FILLER_10_860 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_4 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_81 ();
 sg13g2_fill_1 FILLER_11_131 ();
 sg13g2_fill_1 FILLER_11_141 ();
 sg13g2_decap_8 FILLER_11_150 ();
 sg13g2_fill_1 FILLER_11_157 ();
 sg13g2_decap_8 FILLER_11_292 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_4 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_8 FILLER_11_424 ();
 sg13g2_decap_8 FILLER_11_431 ();
 sg13g2_decap_8 FILLER_11_438 ();
 sg13g2_decap_8 FILLER_11_445 ();
 sg13g2_decap_8 FILLER_11_452 ();
 sg13g2_decap_8 FILLER_11_459 ();
 sg13g2_decap_8 FILLER_11_466 ();
 sg13g2_fill_2 FILLER_11_473 ();
 sg13g2_decap_8 FILLER_11_479 ();
 sg13g2_fill_2 FILLER_11_486 ();
 sg13g2_fill_1 FILLER_11_488 ();
 sg13g2_fill_2 FILLER_11_556 ();
 sg13g2_decap_8 FILLER_11_584 ();
 sg13g2_decap_8 FILLER_11_591 ();
 sg13g2_decap_8 FILLER_11_598 ();
 sg13g2_decap_8 FILLER_11_605 ();
 sg13g2_decap_8 FILLER_11_612 ();
 sg13g2_decap_8 FILLER_11_619 ();
 sg13g2_decap_8 FILLER_11_626 ();
 sg13g2_decap_8 FILLER_11_633 ();
 sg13g2_decap_8 FILLER_11_640 ();
 sg13g2_decap_8 FILLER_11_647 ();
 sg13g2_decap_8 FILLER_11_654 ();
 sg13g2_decap_8 FILLER_11_661 ();
 sg13g2_decap_8 FILLER_11_668 ();
 sg13g2_decap_8 FILLER_11_675 ();
 sg13g2_decap_8 FILLER_11_682 ();
 sg13g2_decap_8 FILLER_11_689 ();
 sg13g2_decap_8 FILLER_11_696 ();
 sg13g2_decap_8 FILLER_11_703 ();
 sg13g2_decap_8 FILLER_11_710 ();
 sg13g2_decap_8 FILLER_11_717 ();
 sg13g2_decap_8 FILLER_11_724 ();
 sg13g2_decap_8 FILLER_11_731 ();
 sg13g2_decap_8 FILLER_11_738 ();
 sg13g2_decap_8 FILLER_11_745 ();
 sg13g2_decap_8 FILLER_11_752 ();
 sg13g2_decap_8 FILLER_11_759 ();
 sg13g2_decap_8 FILLER_11_766 ();
 sg13g2_decap_8 FILLER_11_773 ();
 sg13g2_decap_8 FILLER_11_780 ();
 sg13g2_decap_8 FILLER_11_787 ();
 sg13g2_decap_8 FILLER_11_794 ();
 sg13g2_decap_8 FILLER_11_801 ();
 sg13g2_decap_8 FILLER_11_808 ();
 sg13g2_decap_8 FILLER_11_815 ();
 sg13g2_decap_8 FILLER_11_822 ();
 sg13g2_decap_8 FILLER_11_829 ();
 sg13g2_decap_8 FILLER_11_836 ();
 sg13g2_decap_8 FILLER_11_843 ();
 sg13g2_decap_8 FILLER_11_850 ();
 sg13g2_decap_4 FILLER_11_857 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_fill_2 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_72 ();
 sg13g2_decap_4 FILLER_12_87 ();
 sg13g2_decap_4 FILLER_12_96 ();
 sg13g2_decap_4 FILLER_12_104 ();
 sg13g2_fill_2 FILLER_12_108 ();
 sg13g2_decap_8 FILLER_12_160 ();
 sg13g2_fill_2 FILLER_12_172 ();
 sg13g2_fill_1 FILLER_12_183 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_fill_2 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_206 ();
 sg13g2_decap_8 FILLER_12_213 ();
 sg13g2_decap_8 FILLER_12_220 ();
 sg13g2_fill_1 FILLER_12_227 ();
 sg13g2_decap_8 FILLER_12_232 ();
 sg13g2_fill_2 FILLER_12_239 ();
 sg13g2_fill_1 FILLER_12_241 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_decap_8 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_274 ();
 sg13g2_fill_1 FILLER_12_276 ();
 sg13g2_fill_2 FILLER_12_281 ();
 sg13g2_fill_1 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_decap_8 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_8 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_12_412 ();
 sg13g2_decap_8 FILLER_12_419 ();
 sg13g2_decap_8 FILLER_12_426 ();
 sg13g2_decap_8 FILLER_12_433 ();
 sg13g2_decap_8 FILLER_12_440 ();
 sg13g2_decap_8 FILLER_12_447 ();
 sg13g2_decap_4 FILLER_12_454 ();
 sg13g2_fill_2 FILLER_12_458 ();
 sg13g2_fill_1 FILLER_12_504 ();
 sg13g2_fill_1 FILLER_12_594 ();
 sg13g2_decap_8 FILLER_12_599 ();
 sg13g2_decap_8 FILLER_12_606 ();
 sg13g2_decap_8 FILLER_12_613 ();
 sg13g2_decap_8 FILLER_12_620 ();
 sg13g2_decap_8 FILLER_12_627 ();
 sg13g2_decap_8 FILLER_12_634 ();
 sg13g2_decap_8 FILLER_12_641 ();
 sg13g2_decap_8 FILLER_12_648 ();
 sg13g2_decap_8 FILLER_12_655 ();
 sg13g2_decap_8 FILLER_12_662 ();
 sg13g2_decap_8 FILLER_12_669 ();
 sg13g2_decap_8 FILLER_12_676 ();
 sg13g2_decap_8 FILLER_12_683 ();
 sg13g2_decap_8 FILLER_12_690 ();
 sg13g2_decap_8 FILLER_12_697 ();
 sg13g2_decap_8 FILLER_12_704 ();
 sg13g2_decap_8 FILLER_12_711 ();
 sg13g2_decap_8 FILLER_12_718 ();
 sg13g2_decap_8 FILLER_12_725 ();
 sg13g2_decap_8 FILLER_12_732 ();
 sg13g2_decap_8 FILLER_12_739 ();
 sg13g2_decap_8 FILLER_12_746 ();
 sg13g2_decap_8 FILLER_12_753 ();
 sg13g2_decap_8 FILLER_12_760 ();
 sg13g2_decap_8 FILLER_12_767 ();
 sg13g2_decap_8 FILLER_12_774 ();
 sg13g2_decap_8 FILLER_12_781 ();
 sg13g2_decap_8 FILLER_12_788 ();
 sg13g2_decap_8 FILLER_12_795 ();
 sg13g2_decap_8 FILLER_12_802 ();
 sg13g2_decap_8 FILLER_12_809 ();
 sg13g2_decap_8 FILLER_12_816 ();
 sg13g2_decap_8 FILLER_12_823 ();
 sg13g2_decap_8 FILLER_12_830 ();
 sg13g2_decap_8 FILLER_12_837 ();
 sg13g2_decap_8 FILLER_12_844 ();
 sg13g2_decap_8 FILLER_12_851 ();
 sg13g2_decap_4 FILLER_12_858 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_115 ();
 sg13g2_decap_8 FILLER_13_202 ();
 sg13g2_fill_2 FILLER_13_209 ();
 sg13g2_decap_8 FILLER_13_237 ();
 sg13g2_decap_8 FILLER_13_244 ();
 sg13g2_decap_8 FILLER_13_251 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_4 FILLER_13_284 ();
 sg13g2_fill_2 FILLER_13_302 ();
 sg13g2_fill_1 FILLER_13_304 ();
 sg13g2_fill_1 FILLER_13_309 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_4 FILLER_13_462 ();
 sg13g2_fill_1 FILLER_13_466 ();
 sg13g2_fill_1 FILLER_13_512 ();
 sg13g2_fill_2 FILLER_13_538 ();
 sg13g2_fill_2 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_613 ();
 sg13g2_decap_8 FILLER_13_620 ();
 sg13g2_decap_8 FILLER_13_627 ();
 sg13g2_decap_8 FILLER_13_634 ();
 sg13g2_decap_8 FILLER_13_641 ();
 sg13g2_decap_8 FILLER_13_648 ();
 sg13g2_decap_8 FILLER_13_655 ();
 sg13g2_decap_8 FILLER_13_662 ();
 sg13g2_decap_8 FILLER_13_669 ();
 sg13g2_decap_8 FILLER_13_676 ();
 sg13g2_decap_8 FILLER_13_683 ();
 sg13g2_decap_8 FILLER_13_690 ();
 sg13g2_decap_8 FILLER_13_697 ();
 sg13g2_decap_8 FILLER_13_704 ();
 sg13g2_decap_8 FILLER_13_711 ();
 sg13g2_decap_8 FILLER_13_718 ();
 sg13g2_decap_8 FILLER_13_725 ();
 sg13g2_decap_8 FILLER_13_732 ();
 sg13g2_decap_8 FILLER_13_739 ();
 sg13g2_decap_8 FILLER_13_746 ();
 sg13g2_decap_8 FILLER_13_753 ();
 sg13g2_decap_8 FILLER_13_760 ();
 sg13g2_decap_8 FILLER_13_767 ();
 sg13g2_decap_8 FILLER_13_774 ();
 sg13g2_decap_8 FILLER_13_781 ();
 sg13g2_decap_8 FILLER_13_788 ();
 sg13g2_decap_8 FILLER_13_795 ();
 sg13g2_decap_8 FILLER_13_802 ();
 sg13g2_decap_8 FILLER_13_809 ();
 sg13g2_decap_8 FILLER_13_816 ();
 sg13g2_decap_8 FILLER_13_823 ();
 sg13g2_decap_8 FILLER_13_830 ();
 sg13g2_decap_8 FILLER_13_837 ();
 sg13g2_decap_8 FILLER_13_844 ();
 sg13g2_decap_8 FILLER_13_851 ();
 sg13g2_decap_4 FILLER_13_858 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_fill_2 FILLER_14_70 ();
 sg13g2_fill_1 FILLER_14_72 ();
 sg13g2_fill_1 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_97 ();
 sg13g2_decap_4 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_107 ();
 sg13g2_fill_2 FILLER_14_117 ();
 sg13g2_fill_2 FILLER_14_145 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_4 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_decap_8 FILLER_14_233 ();
 sg13g2_decap_8 FILLER_14_240 ();
 sg13g2_decap_4 FILLER_14_247 ();
 sg13g2_fill_2 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_344 ();
 sg13g2_fill_2 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_4 FILLER_14_469 ();
 sg13g2_fill_1 FILLER_14_473 ();
 sg13g2_fill_1 FILLER_14_500 ();
 sg13g2_fill_2 FILLER_14_536 ();
 sg13g2_fill_2 FILLER_14_572 ();
 sg13g2_fill_1 FILLER_14_589 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_4 FILLER_15_63 ();
 sg13g2_fill_2 FILLER_15_67 ();
 sg13g2_fill_1 FILLER_15_121 ();
 sg13g2_fill_1 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_161 ();
 sg13g2_fill_1 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_190 ();
 sg13g2_fill_1 FILLER_15_204 ();
 sg13g2_fill_1 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_220 ();
 sg13g2_fill_2 FILLER_15_227 ();
 sg13g2_fill_1 FILLER_15_229 ();
 sg13g2_decap_8 FILLER_15_239 ();
 sg13g2_fill_1 FILLER_15_246 ();
 sg13g2_decap_8 FILLER_15_250 ();
 sg13g2_decap_8 FILLER_15_257 ();
 sg13g2_decap_4 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_4 FILLER_15_280 ();
 sg13g2_fill_1 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_299 ();
 sg13g2_fill_1 FILLER_15_313 ();
 sg13g2_fill_1 FILLER_15_328 ();
 sg13g2_fill_2 FILLER_15_333 ();
 sg13g2_decap_8 FILLER_15_387 ();
 sg13g2_fill_1 FILLER_15_394 ();
 sg13g2_decap_4 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_decap_8 FILLER_15_431 ();
 sg13g2_decap_8 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_decap_8 FILLER_15_459 ();
 sg13g2_fill_2 FILLER_15_466 ();
 sg13g2_fill_1 FILLER_15_468 ();
 sg13g2_fill_1 FILLER_15_495 ();
 sg13g2_fill_2 FILLER_15_509 ();
 sg13g2_fill_1 FILLER_15_511 ();
 sg13g2_fill_2 FILLER_15_517 ();
 sg13g2_fill_1 FILLER_15_533 ();
 sg13g2_fill_2 FILLER_15_553 ();
 sg13g2_fill_1 FILLER_15_555 ();
 sg13g2_fill_2 FILLER_15_565 ();
 sg13g2_fill_1 FILLER_15_567 ();
 sg13g2_fill_2 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_618 ();
 sg13g2_decap_8 FILLER_15_625 ();
 sg13g2_decap_8 FILLER_15_632 ();
 sg13g2_decap_8 FILLER_15_639 ();
 sg13g2_decap_4 FILLER_15_646 ();
 sg13g2_fill_1 FILLER_15_650 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_4 FILLER_16_35 ();
 sg13g2_fill_2 FILLER_16_39 ();
 sg13g2_decap_4 FILLER_16_50 ();
 sg13g2_fill_2 FILLER_16_54 ();
 sg13g2_fill_2 FILLER_16_61 ();
 sg13g2_decap_4 FILLER_16_67 ();
 sg13g2_fill_1 FILLER_16_71 ();
 sg13g2_decap_8 FILLER_16_87 ();
 sg13g2_decap_8 FILLER_16_94 ();
 sg13g2_decap_4 FILLER_16_101 ();
 sg13g2_fill_1 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_110 ();
 sg13g2_decap_4 FILLER_16_117 ();
 sg13g2_fill_1 FILLER_16_121 ();
 sg13g2_decap_4 FILLER_16_131 ();
 sg13g2_fill_2 FILLER_16_135 ();
 sg13g2_fill_2 FILLER_16_145 ();
 sg13g2_decap_4 FILLER_16_269 ();
 sg13g2_fill_2 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_decap_8 FILLER_16_325 ();
 sg13g2_decap_4 FILLER_16_332 ();
 sg13g2_fill_1 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_fill_2 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_447 ();
 sg13g2_decap_4 FILLER_16_454 ();
 sg13g2_fill_2 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_4 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_484 ();
 sg13g2_decap_4 FILLER_16_491 ();
 sg13g2_fill_1 FILLER_16_504 ();
 sg13g2_decap_4 FILLER_16_515 ();
 sg13g2_fill_1 FILLER_16_519 ();
 sg13g2_fill_2 FILLER_16_581 ();
 sg13g2_fill_1 FILLER_16_583 ();
 sg13g2_decap_8 FILLER_16_610 ();
 sg13g2_decap_4 FILLER_16_617 ();
 sg13g2_fill_2 FILLER_16_625 ();
 sg13g2_decap_8 FILLER_16_634 ();
 sg13g2_fill_2 FILLER_16_641 ();
 sg13g2_fill_1 FILLER_16_643 ();
 sg13g2_decap_8 FILLER_16_670 ();
 sg13g2_fill_1 FILLER_16_677 ();
 sg13g2_decap_8 FILLER_16_682 ();
 sg13g2_decap_8 FILLER_16_689 ();
 sg13g2_decap_8 FILLER_16_696 ();
 sg13g2_decap_8 FILLER_16_703 ();
 sg13g2_decap_8 FILLER_16_710 ();
 sg13g2_decap_8 FILLER_16_717 ();
 sg13g2_decap_8 FILLER_16_724 ();
 sg13g2_decap_8 FILLER_16_731 ();
 sg13g2_decap_8 FILLER_16_738 ();
 sg13g2_decap_8 FILLER_16_745 ();
 sg13g2_decap_8 FILLER_16_752 ();
 sg13g2_decap_8 FILLER_16_759 ();
 sg13g2_decap_8 FILLER_16_766 ();
 sg13g2_decap_8 FILLER_16_773 ();
 sg13g2_decap_8 FILLER_16_780 ();
 sg13g2_decap_8 FILLER_16_787 ();
 sg13g2_decap_8 FILLER_16_794 ();
 sg13g2_decap_8 FILLER_16_801 ();
 sg13g2_decap_8 FILLER_16_808 ();
 sg13g2_decap_8 FILLER_16_815 ();
 sg13g2_decap_8 FILLER_16_822 ();
 sg13g2_decap_8 FILLER_16_829 ();
 sg13g2_decap_8 FILLER_16_836 ();
 sg13g2_decap_8 FILLER_16_843 ();
 sg13g2_decap_8 FILLER_16_850 ();
 sg13g2_decap_4 FILLER_16_857 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_95 ();
 sg13g2_decap_8 FILLER_17_102 ();
 sg13g2_decap_4 FILLER_17_109 ();
 sg13g2_decap_4 FILLER_17_117 ();
 sg13g2_decap_8 FILLER_17_166 ();
 sg13g2_decap_4 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_194 ();
 sg13g2_fill_2 FILLER_17_213 ();
 sg13g2_decap_8 FILLER_17_219 ();
 sg13g2_fill_2 FILLER_17_226 ();
 sg13g2_fill_2 FILLER_17_261 ();
 sg13g2_fill_1 FILLER_17_263 ();
 sg13g2_fill_2 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_4 FILLER_17_343 ();
 sg13g2_fill_2 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_fill_1 FILLER_17_382 ();
 sg13g2_decap_4 FILLER_17_392 ();
 sg13g2_fill_2 FILLER_17_396 ();
 sg13g2_decap_8 FILLER_17_407 ();
 sg13g2_decap_4 FILLER_17_414 ();
 sg13g2_fill_1 FILLER_17_418 ();
 sg13g2_decap_4 FILLER_17_423 ();
 sg13g2_fill_2 FILLER_17_467 ();
 sg13g2_fill_1 FILLER_17_469 ();
 sg13g2_fill_2 FILLER_17_496 ();
 sg13g2_fill_1 FILLER_17_508 ();
 sg13g2_fill_1 FILLER_17_527 ();
 sg13g2_fill_2 FILLER_17_538 ();
 sg13g2_fill_2 FILLER_17_554 ();
 sg13g2_decap_8 FILLER_17_604 ();
 sg13g2_decap_4 FILLER_17_611 ();
 sg13g2_fill_1 FILLER_17_615 ();
 sg13g2_decap_4 FILLER_17_663 ();
 sg13g2_decap_8 FILLER_17_697 ();
 sg13g2_decap_8 FILLER_17_704 ();
 sg13g2_decap_8 FILLER_17_711 ();
 sg13g2_decap_8 FILLER_17_718 ();
 sg13g2_decap_8 FILLER_17_725 ();
 sg13g2_decap_8 FILLER_17_732 ();
 sg13g2_decap_8 FILLER_17_739 ();
 sg13g2_decap_8 FILLER_17_746 ();
 sg13g2_decap_8 FILLER_17_753 ();
 sg13g2_decap_8 FILLER_17_760 ();
 sg13g2_decap_8 FILLER_17_767 ();
 sg13g2_decap_8 FILLER_17_774 ();
 sg13g2_decap_8 FILLER_17_781 ();
 sg13g2_decap_8 FILLER_17_788 ();
 sg13g2_decap_8 FILLER_17_795 ();
 sg13g2_decap_8 FILLER_17_802 ();
 sg13g2_decap_8 FILLER_17_809 ();
 sg13g2_decap_8 FILLER_17_816 ();
 sg13g2_decap_8 FILLER_17_823 ();
 sg13g2_decap_8 FILLER_17_830 ();
 sg13g2_decap_8 FILLER_17_837 ();
 sg13g2_decap_8 FILLER_17_844 ();
 sg13g2_decap_8 FILLER_17_851 ();
 sg13g2_decap_4 FILLER_17_858 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_fill_1 FILLER_18_128 ();
 sg13g2_fill_1 FILLER_18_143 ();
 sg13g2_fill_2 FILLER_18_149 ();
 sg13g2_fill_2 FILLER_18_255 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_fill_2 FILLER_18_291 ();
 sg13g2_fill_1 FILLER_18_293 ();
 sg13g2_fill_2 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_414 ();
 sg13g2_fill_2 FILLER_18_421 ();
 sg13g2_fill_2 FILLER_18_445 ();
 sg13g2_fill_1 FILLER_18_447 ();
 sg13g2_decap_4 FILLER_18_474 ();
 sg13g2_fill_2 FILLER_18_478 ();
 sg13g2_fill_2 FILLER_18_506 ();
 sg13g2_fill_2 FILLER_18_522 ();
 sg13g2_fill_1 FILLER_18_539 ();
 sg13g2_fill_1 FILLER_18_549 ();
 sg13g2_fill_1 FILLER_18_559 ();
 sg13g2_decap_8 FILLER_18_587 ();
 sg13g2_decap_8 FILLER_18_594 ();
 sg13g2_decap_8 FILLER_18_601 ();
 sg13g2_fill_2 FILLER_18_608 ();
 sg13g2_fill_1 FILLER_18_610 ();
 sg13g2_fill_1 FILLER_18_624 ();
 sg13g2_decap_8 FILLER_18_703 ();
 sg13g2_decap_8 FILLER_18_710 ();
 sg13g2_decap_8 FILLER_18_717 ();
 sg13g2_decap_8 FILLER_18_724 ();
 sg13g2_decap_8 FILLER_18_731 ();
 sg13g2_decap_8 FILLER_18_738 ();
 sg13g2_decap_8 FILLER_18_745 ();
 sg13g2_decap_8 FILLER_18_752 ();
 sg13g2_decap_8 FILLER_18_759 ();
 sg13g2_decap_8 FILLER_18_766 ();
 sg13g2_decap_8 FILLER_18_773 ();
 sg13g2_decap_8 FILLER_18_780 ();
 sg13g2_decap_8 FILLER_18_787 ();
 sg13g2_decap_8 FILLER_18_794 ();
 sg13g2_decap_8 FILLER_18_801 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_829 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_decap_8 FILLER_18_843 ();
 sg13g2_decap_8 FILLER_18_850 ();
 sg13g2_decap_4 FILLER_18_857 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_4 FILLER_19_18 ();
 sg13g2_fill_2 FILLER_19_22 ();
 sg13g2_fill_2 FILLER_19_29 ();
 sg13g2_fill_2 FILLER_19_54 ();
 sg13g2_fill_2 FILLER_19_75 ();
 sg13g2_decap_8 FILLER_19_96 ();
 sg13g2_decap_4 FILLER_19_115 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_fill_1 FILLER_19_163 ();
 sg13g2_decap_4 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_185 ();
 sg13g2_fill_2 FILLER_19_190 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_229 ();
 sg13g2_decap_4 FILLER_19_236 ();
 sg13g2_fill_2 FILLER_19_244 ();
 sg13g2_fill_2 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_304 ();
 sg13g2_decap_4 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_351 ();
 sg13g2_fill_2 FILLER_19_358 ();
 sg13g2_fill_1 FILLER_19_360 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_fill_2 FILLER_19_396 ();
 sg13g2_fill_2 FILLER_19_402 ();
 sg13g2_fill_1 FILLER_19_404 ();
 sg13g2_fill_2 FILLER_19_450 ();
 sg13g2_fill_1 FILLER_19_452 ();
 sg13g2_fill_2 FILLER_19_458 ();
 sg13g2_fill_2 FILLER_19_473 ();
 sg13g2_fill_1 FILLER_19_475 ();
 sg13g2_decap_8 FILLER_19_480 ();
 sg13g2_decap_8 FILLER_19_487 ();
 sg13g2_fill_2 FILLER_19_499 ();
 sg13g2_fill_1 FILLER_19_501 ();
 sg13g2_fill_1 FILLER_19_536 ();
 sg13g2_fill_1 FILLER_19_571 ();
 sg13g2_decap_8 FILLER_19_576 ();
 sg13g2_decap_8 FILLER_19_583 ();
 sg13g2_decap_8 FILLER_19_590 ();
 sg13g2_decap_4 FILLER_19_597 ();
 sg13g2_fill_1 FILLER_19_601 ();
 sg13g2_decap_8 FILLER_19_718 ();
 sg13g2_decap_8 FILLER_19_725 ();
 sg13g2_decap_8 FILLER_19_732 ();
 sg13g2_decap_8 FILLER_19_739 ();
 sg13g2_decap_8 FILLER_19_746 ();
 sg13g2_decap_8 FILLER_19_753 ();
 sg13g2_decap_8 FILLER_19_760 ();
 sg13g2_decap_8 FILLER_19_767 ();
 sg13g2_decap_8 FILLER_19_774 ();
 sg13g2_decap_8 FILLER_19_781 ();
 sg13g2_decap_8 FILLER_19_788 ();
 sg13g2_decap_8 FILLER_19_795 ();
 sg13g2_decap_8 FILLER_19_802 ();
 sg13g2_decap_8 FILLER_19_809 ();
 sg13g2_decap_8 FILLER_19_816 ();
 sg13g2_decap_8 FILLER_19_823 ();
 sg13g2_decap_8 FILLER_19_830 ();
 sg13g2_decap_8 FILLER_19_837 ();
 sg13g2_decap_8 FILLER_19_844 ();
 sg13g2_decap_8 FILLER_19_851 ();
 sg13g2_decap_4 FILLER_19_858 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_2 FILLER_20_42 ();
 sg13g2_fill_2 FILLER_20_106 ();
 sg13g2_fill_1 FILLER_20_108 ();
 sg13g2_decap_4 FILLER_20_144 ();
 sg13g2_decap_4 FILLER_20_163 ();
 sg13g2_fill_2 FILLER_20_193 ();
 sg13g2_fill_1 FILLER_20_195 ();
 sg13g2_fill_2 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_225 ();
 sg13g2_fill_1 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_324 ();
 sg13g2_fill_2 FILLER_20_331 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_fill_1 FILLER_20_380 ();
 sg13g2_fill_2 FILLER_20_386 ();
 sg13g2_fill_2 FILLER_20_402 ();
 sg13g2_fill_1 FILLER_20_404 ();
 sg13g2_fill_2 FILLER_20_425 ();
 sg13g2_fill_2 FILLER_20_453 ();
 sg13g2_fill_1 FILLER_20_455 ();
 sg13g2_decap_4 FILLER_20_491 ();
 sg13g2_fill_1 FILLER_20_495 ();
 sg13g2_fill_1 FILLER_20_505 ();
 sg13g2_fill_2 FILLER_20_519 ();
 sg13g2_fill_1 FILLER_20_521 ();
 sg13g2_fill_2 FILLER_20_542 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_4 FILLER_20_588 ();
 sg13g2_fill_1 FILLER_20_592 ();
 sg13g2_fill_2 FILLER_20_596 ();
 sg13g2_fill_1 FILLER_20_611 ();
 sg13g2_fill_1 FILLER_20_659 ();
 sg13g2_fill_1 FILLER_20_669 ();
 sg13g2_fill_2 FILLER_20_690 ();
 sg13g2_decap_8 FILLER_20_727 ();
 sg13g2_decap_8 FILLER_20_734 ();
 sg13g2_decap_8 FILLER_20_741 ();
 sg13g2_decap_8 FILLER_20_748 ();
 sg13g2_decap_8 FILLER_20_755 ();
 sg13g2_decap_8 FILLER_20_762 ();
 sg13g2_decap_8 FILLER_20_769 ();
 sg13g2_decap_8 FILLER_20_776 ();
 sg13g2_decap_8 FILLER_20_783 ();
 sg13g2_decap_8 FILLER_20_790 ();
 sg13g2_decap_8 FILLER_20_797 ();
 sg13g2_decap_8 FILLER_20_804 ();
 sg13g2_decap_8 FILLER_20_811 ();
 sg13g2_decap_8 FILLER_20_818 ();
 sg13g2_decap_8 FILLER_20_825 ();
 sg13g2_decap_8 FILLER_20_832 ();
 sg13g2_decap_8 FILLER_20_839 ();
 sg13g2_decap_8 FILLER_20_846 ();
 sg13g2_decap_8 FILLER_20_853 ();
 sg13g2_fill_2 FILLER_20_860 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_4 FILLER_21_14 ();
 sg13g2_fill_2 FILLER_21_18 ();
 sg13g2_fill_2 FILLER_21_36 ();
 sg13g2_fill_1 FILLER_21_38 ();
 sg13g2_fill_2 FILLER_21_63 ();
 sg13g2_fill_1 FILLER_21_65 ();
 sg13g2_decap_4 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_74 ();
 sg13g2_fill_1 FILLER_21_93 ();
 sg13g2_fill_2 FILLER_21_102 ();
 sg13g2_fill_1 FILLER_21_104 ();
 sg13g2_fill_2 FILLER_21_125 ();
 sg13g2_fill_2 FILLER_21_148 ();
 sg13g2_fill_1 FILLER_21_155 ();
 sg13g2_decap_4 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_178 ();
 sg13g2_fill_1 FILLER_21_185 ();
 sg13g2_decap_4 FILLER_21_197 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_252 ();
 sg13g2_fill_1 FILLER_21_254 ();
 sg13g2_fill_1 FILLER_21_279 ();
 sg13g2_fill_1 FILLER_21_302 ();
 sg13g2_fill_2 FILLER_21_319 ();
 sg13g2_fill_1 FILLER_21_321 ();
 sg13g2_decap_4 FILLER_21_357 ();
 sg13g2_fill_1 FILLER_21_370 ();
 sg13g2_fill_2 FILLER_21_479 ();
 sg13g2_decap_8 FILLER_21_488 ();
 sg13g2_fill_1 FILLER_21_495 ();
 sg13g2_fill_2 FILLER_21_570 ();
 sg13g2_decap_8 FILLER_21_576 ();
 sg13g2_decap_4 FILLER_21_583 ();
 sg13g2_fill_1 FILLER_21_587 ();
 sg13g2_fill_2 FILLER_21_614 ();
 sg13g2_fill_2 FILLER_21_666 ();
 sg13g2_fill_2 FILLER_21_677 ();
 sg13g2_fill_1 FILLER_21_679 ();
 sg13g2_fill_1 FILLER_21_716 ();
 sg13g2_decap_8 FILLER_21_726 ();
 sg13g2_decap_8 FILLER_21_733 ();
 sg13g2_decap_8 FILLER_21_740 ();
 sg13g2_decap_8 FILLER_21_747 ();
 sg13g2_decap_8 FILLER_21_754 ();
 sg13g2_decap_8 FILLER_21_761 ();
 sg13g2_decap_8 FILLER_21_768 ();
 sg13g2_decap_8 FILLER_21_775 ();
 sg13g2_decap_8 FILLER_21_782 ();
 sg13g2_decap_8 FILLER_21_789 ();
 sg13g2_decap_8 FILLER_21_796 ();
 sg13g2_decap_8 FILLER_21_803 ();
 sg13g2_decap_8 FILLER_21_810 ();
 sg13g2_decap_8 FILLER_21_817 ();
 sg13g2_decap_8 FILLER_21_824 ();
 sg13g2_decap_8 FILLER_21_831 ();
 sg13g2_decap_8 FILLER_21_838 ();
 sg13g2_decap_8 FILLER_21_845 ();
 sg13g2_decap_8 FILLER_21_852 ();
 sg13g2_fill_2 FILLER_21_859 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_fill_1 FILLER_22_36 ();
 sg13g2_fill_2 FILLER_22_80 ();
 sg13g2_decap_8 FILLER_22_87 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_fill_1 FILLER_22_145 ();
 sg13g2_decap_4 FILLER_22_172 ();
 sg13g2_fill_2 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_200 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_decap_8 FILLER_22_215 ();
 sg13g2_decap_8 FILLER_22_222 ();
 sg13g2_fill_2 FILLER_22_229 ();
 sg13g2_fill_1 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_4 FILLER_22_252 ();
 sg13g2_fill_2 FILLER_22_273 ();
 sg13g2_fill_1 FILLER_22_279 ();
 sg13g2_fill_2 FILLER_22_332 ();
 sg13g2_fill_2 FILLER_22_356 ();
 sg13g2_fill_1 FILLER_22_384 ();
 sg13g2_fill_1 FILLER_22_394 ();
 sg13g2_fill_2 FILLER_22_400 ();
 sg13g2_fill_1 FILLER_22_402 ();
 sg13g2_fill_2 FILLER_22_425 ();
 sg13g2_fill_1 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_4 FILLER_22_441 ();
 sg13g2_fill_1 FILLER_22_445 ();
 sg13g2_fill_1 FILLER_22_457 ();
 sg13g2_fill_2 FILLER_22_496 ();
 sg13g2_fill_1 FILLER_22_498 ();
 sg13g2_decap_8 FILLER_22_503 ();
 sg13g2_fill_2 FILLER_22_510 ();
 sg13g2_fill_1 FILLER_22_512 ();
 sg13g2_fill_2 FILLER_22_551 ();
 sg13g2_fill_1 FILLER_22_598 ();
 sg13g2_fill_1 FILLER_22_603 ();
 sg13g2_fill_2 FILLER_22_617 ();
 sg13g2_fill_1 FILLER_22_619 ();
 sg13g2_fill_1 FILLER_22_630 ();
 sg13g2_fill_1 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_731 ();
 sg13g2_decap_8 FILLER_22_738 ();
 sg13g2_decap_8 FILLER_22_745 ();
 sg13g2_decap_8 FILLER_22_752 ();
 sg13g2_decap_8 FILLER_22_759 ();
 sg13g2_decap_8 FILLER_22_766 ();
 sg13g2_decap_8 FILLER_22_773 ();
 sg13g2_decap_8 FILLER_22_780 ();
 sg13g2_decap_8 FILLER_22_787 ();
 sg13g2_decap_8 FILLER_22_794 ();
 sg13g2_decap_8 FILLER_22_801 ();
 sg13g2_decap_8 FILLER_22_808 ();
 sg13g2_decap_8 FILLER_22_815 ();
 sg13g2_decap_8 FILLER_22_822 ();
 sg13g2_decap_8 FILLER_22_829 ();
 sg13g2_decap_8 FILLER_22_836 ();
 sg13g2_decap_8 FILLER_22_843 ();
 sg13g2_decap_8 FILLER_22_850 ();
 sg13g2_decap_4 FILLER_22_857 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_4 FILLER_23_70 ();
 sg13g2_decap_4 FILLER_23_85 ();
 sg13g2_fill_2 FILLER_23_89 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_1 FILLER_23_118 ();
 sg13g2_fill_1 FILLER_23_124 ();
 sg13g2_decap_4 FILLER_23_134 ();
 sg13g2_decap_4 FILLER_23_152 ();
 sg13g2_fill_1 FILLER_23_156 ();
 sg13g2_decap_4 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_173 ();
 sg13g2_fill_1 FILLER_23_180 ();
 sg13g2_fill_2 FILLER_23_190 ();
 sg13g2_fill_1 FILLER_23_192 ();
 sg13g2_fill_1 FILLER_23_210 ();
 sg13g2_fill_2 FILLER_23_229 ();
 sg13g2_fill_1 FILLER_23_231 ();
 sg13g2_fill_2 FILLER_23_244 ();
 sg13g2_fill_1 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_278 ();
 sg13g2_decap_4 FILLER_23_285 ();
 sg13g2_fill_2 FILLER_23_289 ();
 sg13g2_decap_8 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_302 ();
 sg13g2_fill_1 FILLER_23_384 ();
 sg13g2_fill_1 FILLER_23_424 ();
 sg13g2_fill_1 FILLER_23_430 ();
 sg13g2_fill_1 FILLER_23_495 ();
 sg13g2_decap_8 FILLER_23_505 ();
 sg13g2_fill_1 FILLER_23_512 ();
 sg13g2_decap_4 FILLER_23_539 ();
 sg13g2_fill_2 FILLER_23_587 ();
 sg13g2_fill_1 FILLER_23_654 ();
 sg13g2_fill_2 FILLER_23_669 ();
 sg13g2_decap_4 FILLER_23_724 ();
 sg13g2_fill_1 FILLER_23_728 ();
 sg13g2_fill_1 FILLER_23_740 ();
 sg13g2_fill_2 FILLER_23_745 ();
 sg13g2_decap_8 FILLER_23_751 ();
 sg13g2_decap_8 FILLER_23_758 ();
 sg13g2_decap_8 FILLER_23_765 ();
 sg13g2_decap_8 FILLER_23_772 ();
 sg13g2_decap_8 FILLER_23_779 ();
 sg13g2_decap_8 FILLER_23_786 ();
 sg13g2_decap_8 FILLER_23_793 ();
 sg13g2_decap_8 FILLER_23_800 ();
 sg13g2_decap_8 FILLER_23_807 ();
 sg13g2_decap_8 FILLER_23_814 ();
 sg13g2_decap_8 FILLER_23_821 ();
 sg13g2_decap_8 FILLER_23_828 ();
 sg13g2_decap_8 FILLER_23_835 ();
 sg13g2_decap_8 FILLER_23_842 ();
 sg13g2_decap_8 FILLER_23_849 ();
 sg13g2_decap_4 FILLER_23_856 ();
 sg13g2_fill_2 FILLER_23_860 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_fill_1 FILLER_24_33 ();
 sg13g2_fill_1 FILLER_24_79 ();
 sg13g2_fill_2 FILLER_24_108 ();
 sg13g2_decap_8 FILLER_24_115 ();
 sg13g2_decap_4 FILLER_24_122 ();
 sg13g2_fill_1 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_fill_2 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_4 FILLER_24_154 ();
 sg13g2_fill_1 FILLER_24_158 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_4 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_decap_4 FILLER_24_193 ();
 sg13g2_fill_2 FILLER_24_197 ();
 sg13g2_decap_4 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_decap_4 FILLER_24_213 ();
 sg13g2_decap_8 FILLER_24_227 ();
 sg13g2_fill_2 FILLER_24_234 ();
 sg13g2_fill_1 FILLER_24_236 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_decap_4 FILLER_24_268 ();
 sg13g2_decap_4 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_300 ();
 sg13g2_fill_2 FILLER_24_307 ();
 sg13g2_decap_4 FILLER_24_321 ();
 sg13g2_fill_1 FILLER_24_325 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_fill_2 FILLER_24_372 ();
 sg13g2_fill_2 FILLER_24_400 ();
 sg13g2_fill_1 FILLER_24_402 ();
 sg13g2_decap_4 FILLER_24_417 ();
 sg13g2_decap_8 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_24_436 ();
 sg13g2_decap_4 FILLER_24_503 ();
 sg13g2_decap_4 FILLER_24_522 ();
 sg13g2_decap_4 FILLER_24_540 ();
 sg13g2_decap_4 FILLER_24_575 ();
 sg13g2_fill_2 FILLER_24_579 ();
 sg13g2_fill_2 FILLER_24_599 ();
 sg13g2_fill_1 FILLER_24_601 ();
 sg13g2_fill_1 FILLER_24_689 ();
 sg13g2_decap_4 FILLER_24_716 ();
 sg13g2_decap_8 FILLER_24_724 ();
 sg13g2_decap_4 FILLER_24_731 ();
 sg13g2_fill_2 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_759 ();
 sg13g2_decap_8 FILLER_24_766 ();
 sg13g2_decap_8 FILLER_24_773 ();
 sg13g2_decap_8 FILLER_24_780 ();
 sg13g2_decap_8 FILLER_24_787 ();
 sg13g2_decap_8 FILLER_24_794 ();
 sg13g2_decap_8 FILLER_24_801 ();
 sg13g2_decap_8 FILLER_24_808 ();
 sg13g2_decap_8 FILLER_24_815 ();
 sg13g2_decap_8 FILLER_24_822 ();
 sg13g2_decap_8 FILLER_24_829 ();
 sg13g2_decap_8 FILLER_24_836 ();
 sg13g2_decap_8 FILLER_24_843 ();
 sg13g2_decap_8 FILLER_24_850 ();
 sg13g2_decap_4 FILLER_24_857 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_fill_1 FILLER_25_26 ();
 sg13g2_fill_1 FILLER_25_34 ();
 sg13g2_fill_2 FILLER_25_67 ();
 sg13g2_fill_1 FILLER_25_91 ();
 sg13g2_fill_2 FILLER_25_130 ();
 sg13g2_fill_1 FILLER_25_140 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_fill_2 FILLER_25_172 ();
 sg13g2_decap_4 FILLER_25_180 ();
 sg13g2_fill_2 FILLER_25_184 ();
 sg13g2_fill_1 FILLER_25_193 ();
 sg13g2_decap_4 FILLER_25_198 ();
 sg13g2_fill_1 FILLER_25_230 ();
 sg13g2_fill_2 FILLER_25_234 ();
 sg13g2_fill_1 FILLER_25_253 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_353 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_fill_2 FILLER_25_371 ();
 sg13g2_fill_1 FILLER_25_373 ();
 sg13g2_fill_2 FILLER_25_409 ();
 sg13g2_decap_4 FILLER_25_429 ();
 sg13g2_fill_1 FILLER_25_433 ();
 sg13g2_fill_2 FILLER_25_446 ();
 sg13g2_decap_8 FILLER_25_515 ();
 sg13g2_decap_4 FILLER_25_522 ();
 sg13g2_fill_2 FILLER_25_526 ();
 sg13g2_fill_2 FILLER_25_665 ();
 sg13g2_fill_1 FILLER_25_667 ();
 sg13g2_fill_2 FILLER_25_703 ();
 sg13g2_decap_8 FILLER_25_774 ();
 sg13g2_decap_8 FILLER_25_781 ();
 sg13g2_decap_8 FILLER_25_788 ();
 sg13g2_decap_8 FILLER_25_795 ();
 sg13g2_decap_8 FILLER_25_802 ();
 sg13g2_decap_8 FILLER_25_809 ();
 sg13g2_decap_8 FILLER_25_816 ();
 sg13g2_decap_8 FILLER_25_823 ();
 sg13g2_decap_8 FILLER_25_830 ();
 sg13g2_decap_8 FILLER_25_837 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_decap_8 FILLER_25_851 ();
 sg13g2_decap_4 FILLER_25_858 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_fill_2 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_23 ();
 sg13g2_decap_4 FILLER_26_50 ();
 sg13g2_fill_2 FILLER_26_54 ();
 sg13g2_fill_2 FILLER_26_60 ();
 sg13g2_fill_2 FILLER_26_80 ();
 sg13g2_fill_1 FILLER_26_82 ();
 sg13g2_decap_4 FILLER_26_94 ();
 sg13g2_fill_1 FILLER_26_102 ();
 sg13g2_fill_1 FILLER_26_107 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_4 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_fill_2 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_209 ();
 sg13g2_fill_1 FILLER_26_236 ();
 sg13g2_fill_2 FILLER_26_260 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_4 FILLER_26_319 ();
 sg13g2_fill_2 FILLER_26_334 ();
 sg13g2_fill_1 FILLER_26_336 ();
 sg13g2_decap_4 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_decap_4 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_26_416 ();
 sg13g2_fill_2 FILLER_26_423 ();
 sg13g2_fill_2 FILLER_26_464 ();
 sg13g2_decap_8 FILLER_26_505 ();
 sg13g2_decap_4 FILLER_26_517 ();
 sg13g2_fill_2 FILLER_26_521 ();
 sg13g2_decap_4 FILLER_26_554 ();
 sg13g2_decap_4 FILLER_26_567 ();
 sg13g2_fill_1 FILLER_26_571 ();
 sg13g2_fill_2 FILLER_26_607 ();
 sg13g2_fill_1 FILLER_26_640 ();
 sg13g2_fill_2 FILLER_26_667 ();
 sg13g2_decap_4 FILLER_26_687 ();
 sg13g2_fill_1 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_695 ();
 sg13g2_decap_8 FILLER_26_702 ();
 sg13g2_fill_1 FILLER_26_709 ();
 sg13g2_fill_2 FILLER_26_753 ();
 sg13g2_fill_1 FILLER_26_755 ();
 sg13g2_decap_8 FILLER_26_780 ();
 sg13g2_decap_8 FILLER_26_787 ();
 sg13g2_decap_8 FILLER_26_794 ();
 sg13g2_decap_8 FILLER_26_801 ();
 sg13g2_decap_8 FILLER_26_808 ();
 sg13g2_decap_8 FILLER_26_815 ();
 sg13g2_decap_8 FILLER_26_822 ();
 sg13g2_decap_8 FILLER_26_829 ();
 sg13g2_decap_8 FILLER_26_836 ();
 sg13g2_decap_8 FILLER_26_843 ();
 sg13g2_decap_8 FILLER_26_850 ();
 sg13g2_decap_4 FILLER_26_857 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_fill_1 FILLER_27_44 ();
 sg13g2_fill_2 FILLER_27_80 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_157 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_fill_2 FILLER_27_186 ();
 sg13g2_decap_4 FILLER_27_193 ();
 sg13g2_decap_4 FILLER_27_202 ();
 sg13g2_fill_2 FILLER_27_206 ();
 sg13g2_decap_8 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_decap_8 FILLER_27_237 ();
 sg13g2_decap_8 FILLER_27_244 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_258 ();
 sg13g2_fill_2 FILLER_27_264 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_fill_1 FILLER_27_330 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_fill_2 FILLER_27_385 ();
 sg13g2_fill_1 FILLER_27_392 ();
 sg13g2_fill_2 FILLER_27_422 ();
 sg13g2_fill_2 FILLER_27_502 ();
 sg13g2_decap_4 FILLER_27_510 ();
 sg13g2_fill_2 FILLER_27_521 ();
 sg13g2_decap_4 FILLER_27_604 ();
 sg13g2_fill_1 FILLER_27_608 ();
 sg13g2_fill_1 FILLER_27_617 ();
 sg13g2_decap_4 FILLER_27_663 ();
 sg13g2_fill_1 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_790 ();
 sg13g2_decap_8 FILLER_27_797 ();
 sg13g2_decap_8 FILLER_27_804 ();
 sg13g2_decap_8 FILLER_27_811 ();
 sg13g2_decap_8 FILLER_27_818 ();
 sg13g2_decap_8 FILLER_27_825 ();
 sg13g2_decap_8 FILLER_27_832 ();
 sg13g2_decap_8 FILLER_27_839 ();
 sg13g2_decap_8 FILLER_27_846 ();
 sg13g2_decap_8 FILLER_27_853 ();
 sg13g2_fill_2 FILLER_27_860 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_fill_2 FILLER_28_63 ();
 sg13g2_fill_1 FILLER_28_65 ();
 sg13g2_fill_2 FILLER_28_116 ();
 sg13g2_fill_1 FILLER_28_118 ();
 sg13g2_fill_2 FILLER_28_124 ();
 sg13g2_fill_1 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_decap_8 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_198 ();
 sg13g2_fill_1 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_fill_2 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_4 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_235 ();
 sg13g2_decap_4 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_265 ();
 sg13g2_decap_8 FILLER_28_306 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_345 ();
 sg13g2_fill_1 FILLER_28_351 ();
 sg13g2_fill_1 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_374 ();
 sg13g2_fill_2 FILLER_28_387 ();
 sg13g2_fill_1 FILLER_28_389 ();
 sg13g2_decap_4 FILLER_28_398 ();
 sg13g2_fill_1 FILLER_28_402 ();
 sg13g2_fill_1 FILLER_28_422 ();
 sg13g2_fill_1 FILLER_28_475 ();
 sg13g2_fill_2 FILLER_28_485 ();
 sg13g2_fill_1 FILLER_28_487 ();
 sg13g2_fill_1 FILLER_28_558 ();
 sg13g2_fill_2 FILLER_28_571 ();
 sg13g2_decap_8 FILLER_28_649 ();
 sg13g2_decap_8 FILLER_28_656 ();
 sg13g2_fill_2 FILLER_28_663 ();
 sg13g2_fill_1 FILLER_28_665 ();
 sg13g2_decap_8 FILLER_28_670 ();
 sg13g2_fill_1 FILLER_28_677 ();
 sg13g2_fill_1 FILLER_28_702 ();
 sg13g2_fill_2 FILLER_28_734 ();
 sg13g2_fill_1 FILLER_28_760 ();
 sg13g2_decap_8 FILLER_28_804 ();
 sg13g2_decap_8 FILLER_28_811 ();
 sg13g2_decap_8 FILLER_28_818 ();
 sg13g2_decap_8 FILLER_28_825 ();
 sg13g2_decap_8 FILLER_28_832 ();
 sg13g2_decap_8 FILLER_28_839 ();
 sg13g2_decap_8 FILLER_28_846 ();
 sg13g2_decap_8 FILLER_28_853 ();
 sg13g2_fill_2 FILLER_28_860 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_15 ();
 sg13g2_fill_1 FILLER_29_17 ();
 sg13g2_fill_1 FILLER_29_42 ();
 sg13g2_decap_4 FILLER_29_53 ();
 sg13g2_decap_4 FILLER_29_90 ();
 sg13g2_fill_2 FILLER_29_94 ();
 sg13g2_fill_2 FILLER_29_100 ();
 sg13g2_fill_1 FILLER_29_110 ();
 sg13g2_decap_4 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_decap_4 FILLER_29_136 ();
 sg13g2_fill_1 FILLER_29_140 ();
 sg13g2_decap_4 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_165 ();
 sg13g2_fill_2 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_194 ();
 sg13g2_decap_4 FILLER_29_199 ();
 sg13g2_fill_1 FILLER_29_203 ();
 sg13g2_fill_1 FILLER_29_217 ();
 sg13g2_fill_2 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_230 ();
 sg13g2_fill_2 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_248 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_323 ();
 sg13g2_fill_2 FILLER_29_329 ();
 sg13g2_fill_1 FILLER_29_339 ();
 sg13g2_fill_2 FILLER_29_353 ();
 sg13g2_decap_4 FILLER_29_378 ();
 sg13g2_fill_2 FILLER_29_395 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_decap_8 FILLER_29_421 ();
 sg13g2_decap_4 FILLER_29_428 ();
 sg13g2_fill_1 FILLER_29_432 ();
 sg13g2_decap_8 FILLER_29_489 ();
 sg13g2_fill_2 FILLER_29_496 ();
 sg13g2_fill_1 FILLER_29_498 ();
 sg13g2_fill_2 FILLER_29_503 ();
 sg13g2_fill_1 FILLER_29_505 ();
 sg13g2_fill_2 FILLER_29_515 ();
 sg13g2_fill_2 FILLER_29_550 ();
 sg13g2_fill_1 FILLER_29_563 ();
 sg13g2_fill_2 FILLER_29_614 ();
 sg13g2_fill_1 FILLER_29_616 ();
 sg13g2_decap_4 FILLER_29_651 ();
 sg13g2_fill_1 FILLER_29_700 ();
 sg13g2_fill_1 FILLER_29_710 ();
 sg13g2_fill_2 FILLER_29_754 ();
 sg13g2_fill_2 FILLER_29_774 ();
 sg13g2_fill_1 FILLER_29_776 ();
 sg13g2_decap_8 FILLER_29_808 ();
 sg13g2_decap_8 FILLER_29_815 ();
 sg13g2_decap_8 FILLER_29_822 ();
 sg13g2_decap_8 FILLER_29_829 ();
 sg13g2_decap_8 FILLER_29_836 ();
 sg13g2_decap_8 FILLER_29_843 ();
 sg13g2_decap_8 FILLER_29_850 ();
 sg13g2_decap_4 FILLER_29_857 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_30_50 ();
 sg13g2_fill_1 FILLER_30_57 ();
 sg13g2_decap_8 FILLER_30_66 ();
 sg13g2_decap_4 FILLER_30_73 ();
 sg13g2_decap_4 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_100 ();
 sg13g2_decap_4 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_116 ();
 sg13g2_fill_1 FILLER_30_127 ();
 sg13g2_fill_1 FILLER_30_160 ();
 sg13g2_fill_2 FILLER_30_166 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_1 FILLER_30_190 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_decap_8 FILLER_30_232 ();
 sg13g2_fill_1 FILLER_30_239 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_335 ();
 sg13g2_fill_2 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_369 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_fill_2 FILLER_30_403 ();
 sg13g2_fill_1 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_30_410 ();
 sg13g2_decap_4 FILLER_30_417 ();
 sg13g2_decap_8 FILLER_30_434 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_fill_1 FILLER_30_448 ();
 sg13g2_decap_4 FILLER_30_466 ();
 sg13g2_fill_2 FILLER_30_470 ();
 sg13g2_decap_4 FILLER_30_476 ();
 sg13g2_fill_1 FILLER_30_480 ();
 sg13g2_fill_2 FILLER_30_507 ();
 sg13g2_fill_1 FILLER_30_538 ();
 sg13g2_fill_2 FILLER_30_578 ();
 sg13g2_fill_1 FILLER_30_580 ();
 sg13g2_decap_4 FILLER_30_585 ();
 sg13g2_decap_4 FILLER_30_592 ();
 sg13g2_fill_2 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_620 ();
 sg13g2_fill_1 FILLER_30_646 ();
 sg13g2_fill_2 FILLER_30_673 ();
 sg13g2_fill_1 FILLER_30_694 ();
 sg13g2_fill_1 FILLER_30_700 ();
 sg13g2_fill_2 FILLER_30_737 ();
 sg13g2_fill_2 FILLER_30_743 ();
 sg13g2_fill_2 FILLER_30_765 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_decap_8 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_828 ();
 sg13g2_decap_8 FILLER_30_835 ();
 sg13g2_decap_8 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_849 ();
 sg13g2_decap_4 FILLER_30_856 ();
 sg13g2_fill_2 FILLER_30_860 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_9 ();
 sg13g2_fill_1 FILLER_31_20 ();
 sg13g2_decap_4 FILLER_31_54 ();
 sg13g2_fill_1 FILLER_31_72 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_90 ();
 sg13g2_decap_4 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_130 ();
 sg13g2_fill_2 FILLER_31_137 ();
 sg13g2_fill_2 FILLER_31_153 ();
 sg13g2_decap_8 FILLER_31_169 ();
 sg13g2_fill_1 FILLER_31_182 ();
 sg13g2_fill_2 FILLER_31_193 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_199 ();
 sg13g2_fill_2 FILLER_31_211 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_fill_1 FILLER_31_219 ();
 sg13g2_decap_4 FILLER_31_224 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_fill_2 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_282 ();
 sg13g2_decap_4 FILLER_31_320 ();
 sg13g2_fill_2 FILLER_31_324 ();
 sg13g2_fill_2 FILLER_31_349 ();
 sg13g2_fill_1 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_381 ();
 sg13g2_fill_2 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_481 ();
 sg13g2_fill_1 FILLER_31_488 ();
 sg13g2_fill_1 FILLER_31_534 ();
 sg13g2_fill_1 FILLER_31_560 ();
 sg13g2_fill_1 FILLER_31_590 ();
 sg13g2_decap_4 FILLER_31_632 ();
 sg13g2_fill_2 FILLER_31_636 ();
 sg13g2_decap_8 FILLER_31_641 ();
 sg13g2_fill_2 FILLER_31_648 ();
 sg13g2_fill_1 FILLER_31_650 ();
 sg13g2_fill_2 FILLER_31_655 ();
 sg13g2_decap_8 FILLER_31_661 ();
 sg13g2_fill_1 FILLER_31_702 ();
 sg13g2_fill_2 FILLER_31_739 ();
 sg13g2_fill_2 FILLER_31_753 ();
 sg13g2_fill_1 FILLER_31_774 ();
 sg13g2_decap_8 FILLER_31_801 ();
 sg13g2_decap_8 FILLER_31_808 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_decap_8 FILLER_31_822 ();
 sg13g2_decap_8 FILLER_31_829 ();
 sg13g2_decap_8 FILLER_31_836 ();
 sg13g2_decap_8 FILLER_31_843 ();
 sg13g2_decap_8 FILLER_31_850 ();
 sg13g2_decap_4 FILLER_31_857 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_fill_2 FILLER_32_67 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_fill_2 FILLER_32_103 ();
 sg13g2_fill_1 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_131 ();
 sg13g2_decap_8 FILLER_32_167 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_fill_2 FILLER_32_188 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_fill_2 FILLER_32_207 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_258 ();
 sg13g2_decap_8 FILLER_32_264 ();
 sg13g2_decap_4 FILLER_32_271 ();
 sg13g2_fill_1 FILLER_32_278 ();
 sg13g2_fill_2 FILLER_32_283 ();
 sg13g2_fill_1 FILLER_32_285 ();
 sg13g2_fill_1 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_316 ();
 sg13g2_decap_4 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_327 ();
 sg13g2_fill_2 FILLER_32_360 ();
 sg13g2_fill_1 FILLER_32_377 ();
 sg13g2_fill_2 FILLER_32_392 ();
 sg13g2_fill_1 FILLER_32_413 ();
 sg13g2_fill_1 FILLER_32_418 ();
 sg13g2_fill_1 FILLER_32_438 ();
 sg13g2_fill_2 FILLER_32_448 ();
 sg13g2_fill_1 FILLER_32_481 ();
 sg13g2_fill_2 FILLER_32_522 ();
 sg13g2_fill_2 FILLER_32_541 ();
 sg13g2_fill_2 FILLER_32_560 ();
 sg13g2_fill_2 FILLER_32_571 ();
 sg13g2_fill_2 FILLER_32_583 ();
 sg13g2_fill_1 FILLER_32_624 ();
 sg13g2_fill_1 FILLER_32_640 ();
 sg13g2_fill_2 FILLER_32_667 ();
 sg13g2_fill_1 FILLER_32_669 ();
 sg13g2_fill_1 FILLER_32_684 ();
 sg13g2_fill_2 FILLER_32_699 ();
 sg13g2_fill_2 FILLER_32_714 ();
 sg13g2_decap_8 FILLER_32_797 ();
 sg13g2_decap_8 FILLER_32_804 ();
 sg13g2_decap_8 FILLER_32_811 ();
 sg13g2_decap_8 FILLER_32_818 ();
 sg13g2_decap_8 FILLER_32_825 ();
 sg13g2_decap_8 FILLER_32_832 ();
 sg13g2_decap_8 FILLER_32_839 ();
 sg13g2_decap_8 FILLER_32_846 ();
 sg13g2_decap_8 FILLER_32_853 ();
 sg13g2_fill_2 FILLER_32_860 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_9 ();
 sg13g2_fill_2 FILLER_33_19 ();
 sg13g2_fill_2 FILLER_33_39 ();
 sg13g2_fill_1 FILLER_33_71 ();
 sg13g2_fill_2 FILLER_33_101 ();
 sg13g2_fill_1 FILLER_33_103 ();
 sg13g2_fill_1 FILLER_33_110 ();
 sg13g2_fill_1 FILLER_33_124 ();
 sg13g2_decap_4 FILLER_33_135 ();
 sg13g2_fill_1 FILLER_33_139 ();
 sg13g2_decap_4 FILLER_33_148 ();
 sg13g2_fill_2 FILLER_33_156 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_fill_2 FILLER_33_193 ();
 sg13g2_fill_1 FILLER_33_195 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_decap_8 FILLER_33_214 ();
 sg13g2_decap_8 FILLER_33_221 ();
 sg13g2_decap_4 FILLER_33_228 ();
 sg13g2_fill_2 FILLER_33_240 ();
 sg13g2_decap_4 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_decap_8 FILLER_33_323 ();
 sg13g2_decap_4 FILLER_33_330 ();
 sg13g2_decap_4 FILLER_33_339 ();
 sg13g2_fill_2 FILLER_33_343 ();
 sg13g2_fill_2 FILLER_33_349 ();
 sg13g2_fill_2 FILLER_33_370 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_2 FILLER_33_413 ();
 sg13g2_fill_1 FILLER_33_415 ();
 sg13g2_fill_1 FILLER_33_421 ();
 sg13g2_fill_2 FILLER_33_431 ();
 sg13g2_fill_1 FILLER_33_433 ();
 sg13g2_fill_2 FILLER_33_448 ();
 sg13g2_decap_4 FILLER_33_480 ();
 sg13g2_fill_1 FILLER_33_484 ();
 sg13g2_fill_2 FILLER_33_511 ();
 sg13g2_fill_1 FILLER_33_540 ();
 sg13g2_fill_2 FILLER_33_596 ();
 sg13g2_fill_2 FILLER_33_619 ();
 sg13g2_decap_8 FILLER_33_647 ();
 sg13g2_decap_8 FILLER_33_654 ();
 sg13g2_decap_8 FILLER_33_661 ();
 sg13g2_fill_1 FILLER_33_668 ();
 sg13g2_fill_1 FILLER_33_673 ();
 sg13g2_fill_2 FILLER_33_700 ();
 sg13g2_fill_1 FILLER_33_702 ();
 sg13g2_decap_8 FILLER_33_785 ();
 sg13g2_decap_8 FILLER_33_792 ();
 sg13g2_decap_8 FILLER_33_799 ();
 sg13g2_decap_8 FILLER_33_806 ();
 sg13g2_decap_8 FILLER_33_813 ();
 sg13g2_decap_8 FILLER_33_820 ();
 sg13g2_decap_8 FILLER_33_827 ();
 sg13g2_decap_8 FILLER_33_834 ();
 sg13g2_decap_8 FILLER_33_841 ();
 sg13g2_decap_8 FILLER_33_848 ();
 sg13g2_decap_8 FILLER_33_855 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_15 ();
 sg13g2_fill_1 FILLER_34_19 ();
 sg13g2_fill_2 FILLER_34_45 ();
 sg13g2_fill_2 FILLER_34_87 ();
 sg13g2_fill_1 FILLER_34_94 ();
 sg13g2_fill_1 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_178 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_214 ();
 sg13g2_decap_8 FILLER_34_225 ();
 sg13g2_decap_4 FILLER_34_232 ();
 sg13g2_decap_8 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_248 ();
 sg13g2_decap_8 FILLER_34_264 ();
 sg13g2_fill_1 FILLER_34_271 ();
 sg13g2_fill_2 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_fill_2 FILLER_34_396 ();
 sg13g2_fill_1 FILLER_34_451 ();
 sg13g2_decap_4 FILLER_34_487 ();
 sg13g2_fill_1 FILLER_34_491 ();
 sg13g2_fill_2 FILLER_34_500 ();
 sg13g2_fill_1 FILLER_34_502 ();
 sg13g2_fill_2 FILLER_34_530 ();
 sg13g2_fill_2 FILLER_34_566 ();
 sg13g2_fill_1 FILLER_34_568 ();
 sg13g2_decap_8 FILLER_34_573 ();
 sg13g2_fill_2 FILLER_34_580 ();
 sg13g2_fill_1 FILLER_34_582 ();
 sg13g2_fill_2 FILLER_34_652 ();
 sg13g2_fill_1 FILLER_34_693 ();
 sg13g2_fill_1 FILLER_34_699 ();
 sg13g2_fill_2 FILLER_34_725 ();
 sg13g2_fill_1 FILLER_34_727 ();
 sg13g2_fill_2 FILLER_34_750 ();
 sg13g2_fill_1 FILLER_34_752 ();
 sg13g2_decap_8 FILLER_34_792 ();
 sg13g2_decap_8 FILLER_34_799 ();
 sg13g2_decap_8 FILLER_34_806 ();
 sg13g2_decap_8 FILLER_34_813 ();
 sg13g2_decap_8 FILLER_34_820 ();
 sg13g2_decap_8 FILLER_34_827 ();
 sg13g2_decap_8 FILLER_34_834 ();
 sg13g2_decap_8 FILLER_34_841 ();
 sg13g2_decap_8 FILLER_34_848 ();
 sg13g2_decap_8 FILLER_34_855 ();
 sg13g2_fill_2 FILLER_35_44 ();
 sg13g2_fill_1 FILLER_35_46 ();
 sg13g2_decap_8 FILLER_35_73 ();
 sg13g2_decap_8 FILLER_35_80 ();
 sg13g2_decap_8 FILLER_35_87 ();
 sg13g2_fill_2 FILLER_35_94 ();
 sg13g2_decap_4 FILLER_35_122 ();
 sg13g2_fill_2 FILLER_35_126 ();
 sg13g2_decap_4 FILLER_35_133 ();
 sg13g2_fill_2 FILLER_35_159 ();
 sg13g2_fill_1 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_166 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_fill_2 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_decap_4 FILLER_35_230 ();
 sg13g2_fill_1 FILLER_35_234 ();
 sg13g2_fill_2 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_fill_2 FILLER_35_269 ();
 sg13g2_fill_1 FILLER_35_298 ();
 sg13g2_fill_2 FILLER_35_317 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_decap_4 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_334 ();
 sg13g2_decap_8 FILLER_35_352 ();
 sg13g2_decap_4 FILLER_35_359 ();
 sg13g2_fill_1 FILLER_35_393 ();
 sg13g2_decap_4 FILLER_35_409 ();
 sg13g2_decap_4 FILLER_35_489 ();
 sg13g2_fill_2 FILLER_35_493 ();
 sg13g2_fill_2 FILLER_35_547 ();
 sg13g2_fill_1 FILLER_35_584 ();
 sg13g2_fill_1 FILLER_35_593 ();
 sg13g2_decap_8 FILLER_35_647 ();
 sg13g2_fill_1 FILLER_35_663 ();
 sg13g2_fill_2 FILLER_35_780 ();
 sg13g2_fill_1 FILLER_35_782 ();
 sg13g2_decap_8 FILLER_35_796 ();
 sg13g2_decap_8 FILLER_35_803 ();
 sg13g2_decap_8 FILLER_35_810 ();
 sg13g2_decap_8 FILLER_35_817 ();
 sg13g2_decap_8 FILLER_35_824 ();
 sg13g2_decap_8 FILLER_35_831 ();
 sg13g2_decap_8 FILLER_35_838 ();
 sg13g2_decap_8 FILLER_35_845 ();
 sg13g2_decap_8 FILLER_35_852 ();
 sg13g2_fill_2 FILLER_35_859 ();
 sg13g2_fill_1 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_4 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_18 ();
 sg13g2_fill_2 FILLER_36_54 ();
 sg13g2_fill_1 FILLER_36_56 ();
 sg13g2_fill_1 FILLER_36_62 ();
 sg13g2_fill_2 FILLER_36_68 ();
 sg13g2_fill_1 FILLER_36_70 ();
 sg13g2_fill_1 FILLER_36_85 ();
 sg13g2_decap_8 FILLER_36_109 ();
 sg13g2_decap_8 FILLER_36_116 ();
 sg13g2_decap_8 FILLER_36_123 ();
 sg13g2_decap_4 FILLER_36_130 ();
 sg13g2_decap_8 FILLER_36_143 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_decap_4 FILLER_36_174 ();
 sg13g2_fill_2 FILLER_36_178 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_fill_1 FILLER_36_189 ();
 sg13g2_decap_4 FILLER_36_195 ();
 sg13g2_fill_2 FILLER_36_199 ();
 sg13g2_decap_4 FILLER_36_209 ();
 sg13g2_fill_2 FILLER_36_213 ();
 sg13g2_fill_2 FILLER_36_225 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_247 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_fill_2 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_decap_4 FILLER_36_352 ();
 sg13g2_fill_2 FILLER_36_402 ();
 sg13g2_fill_2 FILLER_36_439 ();
 sg13g2_fill_2 FILLER_36_476 ();
 sg13g2_fill_1 FILLER_36_510 ();
 sg13g2_fill_2 FILLER_36_519 ();
 sg13g2_fill_1 FILLER_36_521 ();
 sg13g2_fill_1 FILLER_36_525 ();
 sg13g2_fill_2 FILLER_36_540 ();
 sg13g2_decap_4 FILLER_36_570 ();
 sg13g2_fill_2 FILLER_36_630 ();
 sg13g2_fill_1 FILLER_36_645 ();
 sg13g2_fill_1 FILLER_36_690 ();
 sg13g2_fill_2 FILLER_36_724 ();
 sg13g2_decap_8 FILLER_36_798 ();
 sg13g2_decap_8 FILLER_36_805 ();
 sg13g2_decap_8 FILLER_36_812 ();
 sg13g2_decap_8 FILLER_36_819 ();
 sg13g2_decap_8 FILLER_36_826 ();
 sg13g2_decap_8 FILLER_36_833 ();
 sg13g2_decap_8 FILLER_36_840 ();
 sg13g2_decap_8 FILLER_36_847 ();
 sg13g2_decap_8 FILLER_36_854 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_34 ();
 sg13g2_fill_1 FILLER_37_46 ();
 sg13g2_fill_2 FILLER_37_71 ();
 sg13g2_fill_1 FILLER_37_73 ();
 sg13g2_fill_1 FILLER_37_80 ();
 sg13g2_decap_8 FILLER_37_101 ();
 sg13g2_fill_2 FILLER_37_113 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_decap_8 FILLER_37_177 ();
 sg13g2_fill_1 FILLER_37_184 ();
 sg13g2_fill_2 FILLER_37_193 ();
 sg13g2_fill_1 FILLER_37_206 ();
 sg13g2_fill_2 FILLER_37_213 ();
 sg13g2_fill_1 FILLER_37_215 ();
 sg13g2_fill_2 FILLER_37_230 ();
 sg13g2_fill_1 FILLER_37_232 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_fill_2 FILLER_37_245 ();
 sg13g2_fill_1 FILLER_37_247 ();
 sg13g2_decap_4 FILLER_37_258 ();
 sg13g2_fill_2 FILLER_37_262 ();
 sg13g2_decap_4 FILLER_37_269 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_decap_8 FILLER_37_323 ();
 sg13g2_fill_1 FILLER_37_330 ();
 sg13g2_fill_1 FILLER_37_362 ();
 sg13g2_fill_2 FILLER_37_393 ();
 sg13g2_fill_1 FILLER_37_395 ();
 sg13g2_fill_1 FILLER_37_410 ();
 sg13g2_fill_1 FILLER_37_428 ();
 sg13g2_decap_8 FILLER_37_442 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_4 FILLER_37_483 ();
 sg13g2_fill_2 FILLER_37_487 ();
 sg13g2_decap_8 FILLER_37_493 ();
 sg13g2_decap_8 FILLER_37_500 ();
 sg13g2_fill_2 FILLER_37_507 ();
 sg13g2_fill_1 FILLER_37_535 ();
 sg13g2_fill_2 FILLER_37_545 ();
 sg13g2_fill_1 FILLER_37_547 ();
 sg13g2_fill_1 FILLER_37_577 ();
 sg13g2_fill_1 FILLER_37_617 ();
 sg13g2_fill_1 FILLER_37_627 ();
 sg13g2_decap_8 FILLER_37_639 ();
 sg13g2_decap_4 FILLER_37_646 ();
 sg13g2_fill_1 FILLER_37_681 ();
 sg13g2_fill_1 FILLER_37_762 ();
 sg13g2_fill_2 FILLER_37_773 ();
 sg13g2_fill_1 FILLER_37_775 ();
 sg13g2_fill_2 FILLER_37_785 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_fill_1 FILLER_37_861 ();
 sg13g2_fill_1 FILLER_38_46 ();
 sg13g2_fill_1 FILLER_38_60 ();
 sg13g2_decap_8 FILLER_38_85 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_fill_1 FILLER_38_94 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_8 FILLER_38_144 ();
 sg13g2_decap_4 FILLER_38_151 ();
 sg13g2_fill_2 FILLER_38_163 ();
 sg13g2_fill_1 FILLER_38_170 ();
 sg13g2_fill_2 FILLER_38_176 ();
 sg13g2_fill_1 FILLER_38_178 ();
 sg13g2_decap_8 FILLER_38_185 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_decap_4 FILLER_38_221 ();
 sg13g2_decap_4 FILLER_38_230 ();
 sg13g2_fill_1 FILLER_38_234 ();
 sg13g2_fill_2 FILLER_38_251 ();
 sg13g2_fill_1 FILLER_38_258 ();
 sg13g2_decap_8 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_291 ();
 sg13g2_fill_1 FILLER_38_293 ();
 sg13g2_fill_2 FILLER_38_298 ();
 sg13g2_fill_2 FILLER_38_308 ();
 sg13g2_fill_1 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_337 ();
 sg13g2_fill_1 FILLER_38_339 ();
 sg13g2_fill_2 FILLER_38_345 ();
 sg13g2_fill_1 FILLER_38_356 ();
 sg13g2_fill_1 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_fill_2 FILLER_38_400 ();
 sg13g2_fill_1 FILLER_38_402 ();
 sg13g2_fill_1 FILLER_38_480 ();
 sg13g2_fill_1 FILLER_38_507 ();
 sg13g2_fill_2 FILLER_38_524 ();
 sg13g2_fill_2 FILLER_38_535 ();
 sg13g2_fill_2 FILLER_38_567 ();
 sg13g2_fill_2 FILLER_38_583 ();
 sg13g2_decap_8 FILLER_38_589 ();
 sg13g2_decap_8 FILLER_38_596 ();
 sg13g2_decap_4 FILLER_38_603 ();
 sg13g2_decap_4 FILLER_38_610 ();
 sg13g2_fill_2 FILLER_38_614 ();
 sg13g2_decap_8 FILLER_38_650 ();
 sg13g2_decap_4 FILLER_38_657 ();
 sg13g2_fill_2 FILLER_38_709 ();
 sg13g2_decap_4 FILLER_38_724 ();
 sg13g2_fill_2 FILLER_38_728 ();
 sg13g2_fill_2 FILLER_38_736 ();
 sg13g2_decap_8 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_749 ();
 sg13g2_fill_2 FILLER_38_790 ();
 sg13g2_decap_8 FILLER_38_818 ();
 sg13g2_decap_8 FILLER_38_825 ();
 sg13g2_decap_8 FILLER_38_832 ();
 sg13g2_decap_8 FILLER_38_839 ();
 sg13g2_decap_8 FILLER_38_846 ();
 sg13g2_decap_8 FILLER_38_853 ();
 sg13g2_fill_2 FILLER_38_860 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_7 ();
 sg13g2_fill_1 FILLER_39_29 ();
 sg13g2_fill_2 FILLER_39_39 ();
 sg13g2_fill_1 FILLER_39_41 ();
 sg13g2_decap_8 FILLER_39_73 ();
 sg13g2_decap_8 FILLER_39_80 ();
 sg13g2_decap_4 FILLER_39_97 ();
 sg13g2_fill_2 FILLER_39_101 ();
 sg13g2_fill_1 FILLER_39_111 ();
 sg13g2_decap_8 FILLER_39_115 ();
 sg13g2_fill_2 FILLER_39_122 ();
 sg13g2_fill_1 FILLER_39_124 ();
 sg13g2_fill_1 FILLER_39_132 ();
 sg13g2_fill_1 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_186 ();
 sg13g2_fill_2 FILLER_39_193 ();
 sg13g2_fill_2 FILLER_39_199 ();
 sg13g2_decap_8 FILLER_39_205 ();
 sg13g2_decap_4 FILLER_39_212 ();
 sg13g2_fill_2 FILLER_39_221 ();
 sg13g2_decap_8 FILLER_39_228 ();
 sg13g2_fill_2 FILLER_39_235 ();
 sg13g2_fill_1 FILLER_39_237 ();
 sg13g2_fill_2 FILLER_39_266 ();
 sg13g2_fill_1 FILLER_39_268 ();
 sg13g2_fill_2 FILLER_39_274 ();
 sg13g2_fill_1 FILLER_39_276 ();
 sg13g2_fill_1 FILLER_39_286 ();
 sg13g2_decap_8 FILLER_39_306 ();
 sg13g2_fill_2 FILLER_39_313 ();
 sg13g2_fill_2 FILLER_39_333 ();
 sg13g2_fill_1 FILLER_39_423 ();
 sg13g2_decap_8 FILLER_39_429 ();
 sg13g2_fill_1 FILLER_39_451 ();
 sg13g2_decap_8 FILLER_39_470 ();
 sg13g2_decap_8 FILLER_39_477 ();
 sg13g2_decap_8 FILLER_39_484 ();
 sg13g2_fill_2 FILLER_39_571 ();
 sg13g2_fill_1 FILLER_39_573 ();
 sg13g2_fill_2 FILLER_39_626 ();
 sg13g2_fill_1 FILLER_39_647 ();
 sg13g2_decap_4 FILLER_39_707 ();
 sg13g2_decap_8 FILLER_39_716 ();
 sg13g2_decap_8 FILLER_39_735 ();
 sg13g2_fill_2 FILLER_39_742 ();
 sg13g2_fill_1 FILLER_39_744 ();
 sg13g2_fill_2 FILLER_39_777 ();
 sg13g2_decap_8 FILLER_39_821 ();
 sg13g2_decap_8 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_842 ();
 sg13g2_decap_8 FILLER_39_849 ();
 sg13g2_decap_4 FILLER_39_856 ();
 sg13g2_fill_2 FILLER_39_860 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_fill_1 FILLER_40_29 ();
 sg13g2_decap_4 FILLER_40_46 ();
 sg13g2_fill_1 FILLER_40_50 ();
 sg13g2_fill_2 FILLER_40_56 ();
 sg13g2_decap_4 FILLER_40_62 ();
 sg13g2_fill_2 FILLER_40_66 ();
 sg13g2_decap_4 FILLER_40_73 ();
 sg13g2_fill_2 FILLER_40_77 ();
 sg13g2_fill_2 FILLER_40_84 ();
 sg13g2_fill_2 FILLER_40_96 ();
 sg13g2_decap_4 FILLER_40_124 ();
 sg13g2_fill_2 FILLER_40_142 ();
 sg13g2_decap_8 FILLER_40_148 ();
 sg13g2_decap_4 FILLER_40_155 ();
 sg13g2_fill_1 FILLER_40_167 ();
 sg13g2_decap_8 FILLER_40_178 ();
 sg13g2_fill_2 FILLER_40_185 ();
 sg13g2_fill_1 FILLER_40_187 ();
 sg13g2_decap_4 FILLER_40_234 ();
 sg13g2_decap_4 FILLER_40_248 ();
 sg13g2_fill_1 FILLER_40_280 ();
 sg13g2_fill_1 FILLER_40_333 ();
 sg13g2_decap_8 FILLER_40_365 ();
 sg13g2_fill_2 FILLER_40_372 ();
 sg13g2_fill_1 FILLER_40_382 ();
 sg13g2_fill_2 FILLER_40_396 ();
 sg13g2_fill_1 FILLER_40_398 ();
 sg13g2_fill_1 FILLER_40_417 ();
 sg13g2_decap_8 FILLER_40_431 ();
 sg13g2_fill_2 FILLER_40_464 ();
 sg13g2_fill_1 FILLER_40_466 ();
 sg13g2_fill_2 FILLER_40_503 ();
 sg13g2_fill_1 FILLER_40_505 ();
 sg13g2_decap_8 FILLER_40_510 ();
 sg13g2_decap_8 FILLER_40_517 ();
 sg13g2_decap_4 FILLER_40_524 ();
 sg13g2_decap_8 FILLER_40_532 ();
 sg13g2_fill_1 FILLER_40_539 ();
 sg13g2_fill_2 FILLER_40_544 ();
 sg13g2_fill_1 FILLER_40_546 ();
 sg13g2_decap_8 FILLER_40_557 ();
 sg13g2_decap_8 FILLER_40_564 ();
 sg13g2_decap_4 FILLER_40_571 ();
 sg13g2_fill_2 FILLER_40_575 ();
 sg13g2_decap_8 FILLER_40_585 ();
 sg13g2_decap_8 FILLER_40_592 ();
 sg13g2_decap_8 FILLER_40_599 ();
 sg13g2_fill_1 FILLER_40_606 ();
 sg13g2_fill_2 FILLER_40_611 ();
 sg13g2_fill_1 FILLER_40_613 ();
 sg13g2_fill_2 FILLER_40_623 ();
 sg13g2_decap_8 FILLER_40_650 ();
 sg13g2_fill_2 FILLER_40_657 ();
 sg13g2_decap_8 FILLER_40_663 ();
 sg13g2_decap_8 FILLER_40_670 ();
 sg13g2_fill_2 FILLER_40_677 ();
 sg13g2_fill_2 FILLER_40_684 ();
 sg13g2_fill_2 FILLER_40_762 ();
 sg13g2_fill_1 FILLER_40_764 ();
 sg13g2_decap_8 FILLER_40_823 ();
 sg13g2_decap_8 FILLER_40_830 ();
 sg13g2_decap_8 FILLER_40_837 ();
 sg13g2_decap_8 FILLER_40_844 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_4 FILLER_40_858 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_33 ();
 sg13g2_decap_8 FILLER_41_39 ();
 sg13g2_fill_1 FILLER_41_46 ();
 sg13g2_decap_8 FILLER_41_52 ();
 sg13g2_decap_8 FILLER_41_59 ();
 sg13g2_fill_2 FILLER_41_129 ();
 sg13g2_decap_8 FILLER_41_146 ();
 sg13g2_fill_1 FILLER_41_153 ();
 sg13g2_fill_1 FILLER_41_166 ();
 sg13g2_decap_8 FILLER_41_186 ();
 sg13g2_decap_8 FILLER_41_193 ();
 sg13g2_decap_4 FILLER_41_200 ();
 sg13g2_fill_1 FILLER_41_204 ();
 sg13g2_decap_8 FILLER_41_212 ();
 sg13g2_decap_4 FILLER_41_280 ();
 sg13g2_fill_2 FILLER_41_284 ();
 sg13g2_decap_4 FILLER_41_326 ();
 sg13g2_fill_1 FILLER_41_330 ();
 sg13g2_decap_4 FILLER_41_336 ();
 sg13g2_fill_1 FILLER_41_340 ();
 sg13g2_decap_8 FILLER_41_354 ();
 sg13g2_fill_1 FILLER_41_361 ();
 sg13g2_fill_2 FILLER_41_381 ();
 sg13g2_fill_2 FILLER_41_388 ();
 sg13g2_fill_2 FILLER_41_405 ();
 sg13g2_fill_1 FILLER_41_407 ();
 sg13g2_fill_2 FILLER_41_434 ();
 sg13g2_fill_1 FILLER_41_436 ();
 sg13g2_fill_1 FILLER_41_450 ();
 sg13g2_decap_8 FILLER_41_493 ();
 sg13g2_decap_4 FILLER_41_500 ();
 sg13g2_decap_8 FILLER_41_512 ();
 sg13g2_decap_8 FILLER_41_524 ();
 sg13g2_decap_8 FILLER_41_531 ();
 sg13g2_decap_4 FILLER_41_538 ();
 sg13g2_fill_2 FILLER_41_542 ();
 sg13g2_fill_2 FILLER_41_556 ();
 sg13g2_decap_8 FILLER_41_566 ();
 sg13g2_decap_8 FILLER_41_589 ();
 sg13g2_decap_4 FILLER_41_615 ();
 sg13g2_decap_8 FILLER_41_643 ();
 sg13g2_decap_4 FILLER_41_650 ();
 sg13g2_fill_1 FILLER_41_654 ();
 sg13g2_decap_4 FILLER_41_660 ();
 sg13g2_fill_1 FILLER_41_664 ();
 sg13g2_fill_2 FILLER_41_671 ();
 sg13g2_fill_2 FILLER_41_681 ();
 sg13g2_fill_1 FILLER_41_691 ();
 sg13g2_fill_1 FILLER_41_705 ();
 sg13g2_decap_8 FILLER_41_720 ();
 sg13g2_fill_2 FILLER_41_727 ();
 sg13g2_fill_2 FILLER_41_733 ();
 sg13g2_fill_1 FILLER_41_735 ();
 sg13g2_fill_2 FILLER_41_745 ();
 sg13g2_fill_1 FILLER_41_747 ();
 sg13g2_fill_2 FILLER_41_806 ();
 sg13g2_fill_1 FILLER_41_808 ();
 sg13g2_decap_8 FILLER_41_822 ();
 sg13g2_decap_8 FILLER_41_829 ();
 sg13g2_decap_8 FILLER_41_836 ();
 sg13g2_decap_8 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_850 ();
 sg13g2_decap_4 FILLER_41_857 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_fill_1 FILLER_42_26 ();
 sg13g2_fill_2 FILLER_42_36 ();
 sg13g2_fill_1 FILLER_42_38 ();
 sg13g2_decap_4 FILLER_42_65 ();
 sg13g2_decap_4 FILLER_42_74 ();
 sg13g2_decap_8 FILLER_42_82 ();
 sg13g2_fill_1 FILLER_42_89 ();
 sg13g2_fill_2 FILLER_42_133 ();
 sg13g2_fill_1 FILLER_42_135 ();
 sg13g2_decap_8 FILLER_42_148 ();
 sg13g2_decap_4 FILLER_42_209 ();
 sg13g2_fill_1 FILLER_42_213 ();
 sg13g2_fill_2 FILLER_42_233 ();
 sg13g2_fill_1 FILLER_42_235 ();
 sg13g2_fill_2 FILLER_42_241 ();
 sg13g2_fill_1 FILLER_42_243 ();
 sg13g2_fill_1 FILLER_42_267 ();
 sg13g2_fill_2 FILLER_42_289 ();
 sg13g2_decap_4 FILLER_42_294 ();
 sg13g2_fill_2 FILLER_42_324 ();
 sg13g2_fill_1 FILLER_42_326 ();
 sg13g2_fill_1 FILLER_42_337 ();
 sg13g2_fill_2 FILLER_42_343 ();
 sg13g2_fill_1 FILLER_42_345 ();
 sg13g2_decap_4 FILLER_42_350 ();
 sg13g2_fill_2 FILLER_42_359 ();
 sg13g2_fill_1 FILLER_42_361 ();
 sg13g2_fill_1 FILLER_42_398 ();
 sg13g2_fill_1 FILLER_42_410 ();
 sg13g2_decap_4 FILLER_42_443 ();
 sg13g2_fill_2 FILLER_42_447 ();
 sg13g2_decap_4 FILLER_42_483 ();
 sg13g2_decap_4 FILLER_42_497 ();
 sg13g2_fill_2 FILLER_42_501 ();
 sg13g2_fill_2 FILLER_42_519 ();
 sg13g2_fill_2 FILLER_42_541 ();
 sg13g2_decap_8 FILLER_42_557 ();
 sg13g2_decap_4 FILLER_42_564 ();
 sg13g2_fill_2 FILLER_42_586 ();
 sg13g2_fill_2 FILLER_42_618 ();
 sg13g2_fill_1 FILLER_42_620 ();
 sg13g2_fill_1 FILLER_42_630 ();
 sg13g2_decap_8 FILLER_42_635 ();
 sg13g2_fill_1 FILLER_42_642 ();
 sg13g2_fill_2 FILLER_42_677 ();
 sg13g2_decap_8 FILLER_42_688 ();
 sg13g2_fill_1 FILLER_42_695 ();
 sg13g2_fill_2 FILLER_42_702 ();
 sg13g2_fill_1 FILLER_42_704 ();
 sg13g2_decap_4 FILLER_42_726 ();
 sg13g2_fill_2 FILLER_42_750 ();
 sg13g2_fill_1 FILLER_42_752 ();
 sg13g2_decap_4 FILLER_42_757 ();
 sg13g2_fill_2 FILLER_42_761 ();
 sg13g2_fill_2 FILLER_42_784 ();
 sg13g2_fill_1 FILLER_42_786 ();
 sg13g2_decap_8 FILLER_42_817 ();
 sg13g2_decap_8 FILLER_42_824 ();
 sg13g2_decap_8 FILLER_42_831 ();
 sg13g2_decap_8 FILLER_42_838 ();
 sg13g2_decap_8 FILLER_42_845 ();
 sg13g2_decap_8 FILLER_42_852 ();
 sg13g2_fill_2 FILLER_42_859 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_15 ();
 sg13g2_fill_1 FILLER_43_48 ();
 sg13g2_decap_4 FILLER_43_54 ();
 sg13g2_fill_1 FILLER_43_58 ();
 sg13g2_decap_4 FILLER_43_64 ();
 sg13g2_fill_2 FILLER_43_68 ();
 sg13g2_fill_1 FILLER_43_80 ();
 sg13g2_decap_4 FILLER_43_86 ();
 sg13g2_fill_2 FILLER_43_90 ();
 sg13g2_fill_2 FILLER_43_125 ();
 sg13g2_fill_1 FILLER_43_127 ();
 sg13g2_fill_2 FILLER_43_143 ();
 sg13g2_fill_2 FILLER_43_155 ();
 sg13g2_fill_1 FILLER_43_186 ();
 sg13g2_fill_2 FILLER_43_218 ();
 sg13g2_fill_1 FILLER_43_220 ();
 sg13g2_fill_2 FILLER_43_286 ();
 sg13g2_decap_4 FILLER_43_296 ();
 sg13g2_fill_1 FILLER_43_317 ();
 sg13g2_fill_1 FILLER_43_322 ();
 sg13g2_fill_2 FILLER_43_333 ();
 sg13g2_fill_1 FILLER_43_380 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_fill_1 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_fill_2 FILLER_43_468 ();
 sg13g2_fill_2 FILLER_43_486 ();
 sg13g2_fill_2 FILLER_43_493 ();
 sg13g2_fill_1 FILLER_43_495 ();
 sg13g2_fill_1 FILLER_43_504 ();
 sg13g2_decap_8 FILLER_43_520 ();
 sg13g2_decap_4 FILLER_43_527 ();
 sg13g2_fill_2 FILLER_43_536 ();
 sg13g2_fill_1 FILLER_43_538 ();
 sg13g2_decap_8 FILLER_43_562 ();
 sg13g2_fill_2 FILLER_43_569 ();
 sg13g2_fill_1 FILLER_43_571 ();
 sg13g2_decap_4 FILLER_43_597 ();
 sg13g2_fill_2 FILLER_43_601 ();
 sg13g2_decap_4 FILLER_43_637 ();
 sg13g2_fill_1 FILLER_43_641 ();
 sg13g2_decap_4 FILLER_43_652 ();
 sg13g2_fill_1 FILLER_43_656 ();
 sg13g2_decap_8 FILLER_43_661 ();
 sg13g2_fill_2 FILLER_43_668 ();
 sg13g2_fill_1 FILLER_43_670 ();
 sg13g2_decap_8 FILLER_43_704 ();
 sg13g2_decap_4 FILLER_43_711 ();
 sg13g2_fill_2 FILLER_43_715 ();
 sg13g2_decap_8 FILLER_43_725 ();
 sg13g2_fill_1 FILLER_43_732 ();
 sg13g2_decap_4 FILLER_43_741 ();
 sg13g2_fill_1 FILLER_43_745 ();
 sg13g2_decap_8 FILLER_43_762 ();
 sg13g2_fill_2 FILLER_43_769 ();
 sg13g2_fill_1 FILLER_43_771 ();
 sg13g2_fill_2 FILLER_43_780 ();
 sg13g2_fill_1 FILLER_43_782 ();
 sg13g2_decap_4 FILLER_43_789 ();
 sg13g2_decap_8 FILLER_43_822 ();
 sg13g2_decap_8 FILLER_43_829 ();
 sg13g2_decap_8 FILLER_43_836 ();
 sg13g2_decap_8 FILLER_43_843 ();
 sg13g2_decap_8 FILLER_43_850 ();
 sg13g2_decap_4 FILLER_43_857 ();
 sg13g2_fill_1 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_4 FILLER_44_46 ();
 sg13g2_decap_4 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_93 ();
 sg13g2_decap_8 FILLER_44_100 ();
 sg13g2_decap_4 FILLER_44_107 ();
 sg13g2_fill_2 FILLER_44_137 ();
 sg13g2_fill_1 FILLER_44_148 ();
 sg13g2_fill_2 FILLER_44_211 ();
 sg13g2_fill_1 FILLER_44_255 ();
 sg13g2_fill_1 FILLER_44_305 ();
 sg13g2_fill_2 FILLER_44_311 ();
 sg13g2_fill_1 FILLER_44_313 ();
 sg13g2_fill_1 FILLER_44_336 ();
 sg13g2_fill_2 FILLER_44_346 ();
 sg13g2_fill_1 FILLER_44_368 ();
 sg13g2_fill_2 FILLER_44_379 ();
 sg13g2_fill_1 FILLER_44_394 ();
 sg13g2_decap_8 FILLER_44_423 ();
 sg13g2_decap_8 FILLER_44_430 ();
 sg13g2_decap_8 FILLER_44_437 ();
 sg13g2_fill_2 FILLER_44_444 ();
 sg13g2_decap_4 FILLER_44_460 ();
 sg13g2_fill_1 FILLER_44_464 ();
 sg13g2_fill_1 FILLER_44_474 ();
 sg13g2_decap_8 FILLER_44_481 ();
 sg13g2_decap_8 FILLER_44_488 ();
 sg13g2_decap_4 FILLER_44_495 ();
 sg13g2_fill_2 FILLER_44_499 ();
 sg13g2_decap_8 FILLER_44_510 ();
 sg13g2_fill_2 FILLER_44_517 ();
 sg13g2_fill_1 FILLER_44_519 ();
 sg13g2_decap_4 FILLER_44_530 ();
 sg13g2_fill_1 FILLER_44_556 ();
 sg13g2_decap_8 FILLER_44_566 ();
 sg13g2_decap_4 FILLER_44_578 ();
 sg13g2_fill_1 FILLER_44_582 ();
 sg13g2_fill_2 FILLER_44_596 ();
 sg13g2_fill_1 FILLER_44_598 ();
 sg13g2_decap_8 FILLER_44_614 ();
 sg13g2_decap_4 FILLER_44_621 ();
 sg13g2_fill_1 FILLER_44_625 ();
 sg13g2_fill_2 FILLER_44_651 ();
 sg13g2_fill_2 FILLER_44_678 ();
 sg13g2_decap_8 FILLER_44_697 ();
 sg13g2_decap_4 FILLER_44_704 ();
 sg13g2_fill_1 FILLER_44_708 ();
 sg13g2_decap_8 FILLER_44_721 ();
 sg13g2_fill_2 FILLER_44_728 ();
 sg13g2_decap_4 FILLER_44_742 ();
 sg13g2_fill_2 FILLER_44_754 ();
 sg13g2_fill_1 FILLER_44_756 ();
 sg13g2_fill_2 FILLER_44_769 ();
 sg13g2_fill_1 FILLER_44_771 ();
 sg13g2_fill_2 FILLER_44_778 ();
 sg13g2_fill_1 FILLER_44_780 ();
 sg13g2_decap_4 FILLER_44_813 ();
 sg13g2_fill_1 FILLER_44_817 ();
 sg13g2_decap_8 FILLER_44_826 ();
 sg13g2_decap_8 FILLER_44_833 ();
 sg13g2_decap_8 FILLER_44_840 ();
 sg13g2_decap_8 FILLER_44_847 ();
 sg13g2_decap_8 FILLER_44_854 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_45 ();
 sg13g2_decap_4 FILLER_45_68 ();
 sg13g2_fill_2 FILLER_45_90 ();
 sg13g2_decap_4 FILLER_45_104 ();
 sg13g2_fill_2 FILLER_45_125 ();
 sg13g2_fill_1 FILLER_45_127 ();
 sg13g2_fill_1 FILLER_45_189 ();
 sg13g2_decap_4 FILLER_45_219 ();
 sg13g2_fill_1 FILLER_45_223 ();
 sg13g2_decap_8 FILLER_45_298 ();
 sg13g2_fill_2 FILLER_45_305 ();
 sg13g2_fill_1 FILLER_45_333 ();
 sg13g2_fill_2 FILLER_45_343 ();
 sg13g2_fill_2 FILLER_45_418 ();
 sg13g2_fill_1 FILLER_45_420 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_decap_4 FILLER_45_462 ();
 sg13g2_decap_8 FILLER_45_482 ();
 sg13g2_fill_2 FILLER_45_489 ();
 sg13g2_fill_1 FILLER_45_491 ();
 sg13g2_fill_2 FILLER_45_512 ();
 sg13g2_decap_4 FILLER_45_528 ();
 sg13g2_fill_2 FILLER_45_532 ();
 sg13g2_fill_2 FILLER_45_544 ();
 sg13g2_decap_4 FILLER_45_550 ();
 sg13g2_fill_1 FILLER_45_554 ();
 sg13g2_decap_4 FILLER_45_560 ();
 sg13g2_fill_1 FILLER_45_564 ();
 sg13g2_decap_8 FILLER_45_570 ();
 sg13g2_fill_2 FILLER_45_577 ();
 sg13g2_fill_1 FILLER_45_579 ();
 sg13g2_decap_8 FILLER_45_585 ();
 sg13g2_decap_8 FILLER_45_592 ();
 sg13g2_decap_8 FILLER_45_604 ();
 sg13g2_decap_4 FILLER_45_611 ();
 sg13g2_fill_2 FILLER_45_625 ();
 sg13g2_fill_1 FILLER_45_627 ();
 sg13g2_decap_8 FILLER_45_636 ();
 sg13g2_decap_8 FILLER_45_643 ();
 sg13g2_decap_8 FILLER_45_650 ();
 sg13g2_decap_4 FILLER_45_657 ();
 sg13g2_decap_8 FILLER_45_666 ();
 sg13g2_decap_8 FILLER_45_673 ();
 sg13g2_fill_2 FILLER_45_680 ();
 sg13g2_fill_1 FILLER_45_682 ();
 sg13g2_decap_4 FILLER_45_693 ();
 sg13g2_fill_2 FILLER_45_697 ();
 sg13g2_decap_4 FILLER_45_719 ();
 sg13g2_decap_8 FILLER_45_739 ();
 sg13g2_fill_2 FILLER_45_746 ();
 sg13g2_fill_1 FILLER_45_753 ();
 sg13g2_fill_2 FILLER_45_770 ();
 sg13g2_fill_1 FILLER_45_772 ();
 sg13g2_decap_8 FILLER_45_779 ();
 sg13g2_decap_8 FILLER_45_786 ();
 sg13g2_decap_4 FILLER_45_793 ();
 sg13g2_fill_2 FILLER_45_797 ();
 sg13g2_decap_8 FILLER_45_805 ();
 sg13g2_fill_1 FILLER_45_812 ();
 sg13g2_fill_1 FILLER_45_841 ();
 sg13g2_decap_8 FILLER_45_853 ();
 sg13g2_fill_2 FILLER_45_860 ();
 sg13g2_fill_1 FILLER_46_51 ();
 sg13g2_fill_2 FILLER_46_61 ();
 sg13g2_decap_4 FILLER_46_97 ();
 sg13g2_fill_2 FILLER_46_101 ();
 sg13g2_decap_8 FILLER_46_109 ();
 sg13g2_decap_4 FILLER_46_116 ();
 sg13g2_fill_1 FILLER_46_120 ();
 sg13g2_decap_8 FILLER_46_151 ();
 sg13g2_decap_4 FILLER_46_161 ();
 sg13g2_decap_4 FILLER_46_182 ();
 sg13g2_decap_4 FILLER_46_190 ();
 sg13g2_fill_1 FILLER_46_194 ();
 sg13g2_fill_2 FILLER_46_216 ();
 sg13g2_fill_1 FILLER_46_218 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_fill_2 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_258 ();
 sg13g2_decap_4 FILLER_46_265 ();
 sg13g2_decap_8 FILLER_46_278 ();
 sg13g2_decap_8 FILLER_46_285 ();
 sg13g2_decap_8 FILLER_46_292 ();
 sg13g2_fill_1 FILLER_46_348 ();
 sg13g2_fill_2 FILLER_46_358 ();
 sg13g2_fill_2 FILLER_46_374 ();
 sg13g2_fill_1 FILLER_46_376 ();
 sg13g2_decap_8 FILLER_46_421 ();
 sg13g2_fill_2 FILLER_46_428 ();
 sg13g2_fill_1 FILLER_46_430 ();
 sg13g2_fill_2 FILLER_46_440 ();
 sg13g2_fill_1 FILLER_46_442 ();
 sg13g2_fill_1 FILLER_46_455 ();
 sg13g2_fill_2 FILLER_46_482 ();
 sg13g2_decap_8 FILLER_46_507 ();
 sg13g2_fill_1 FILLER_46_514 ();
 sg13g2_fill_1 FILLER_46_520 ();
 sg13g2_fill_1 FILLER_46_535 ();
 sg13g2_decap_4 FILLER_46_563 ();
 sg13g2_fill_2 FILLER_46_590 ();
 sg13g2_fill_1 FILLER_46_597 ();
 sg13g2_fill_2 FILLER_46_613 ();
 sg13g2_decap_4 FILLER_46_642 ();
 sg13g2_fill_2 FILLER_46_655 ();
 sg13g2_fill_1 FILLER_46_657 ();
 sg13g2_fill_2 FILLER_46_691 ();
 sg13g2_fill_1 FILLER_46_693 ();
 sg13g2_decap_8 FILLER_46_717 ();
 sg13g2_decap_8 FILLER_46_736 ();
 sg13g2_decap_4 FILLER_46_743 ();
 sg13g2_fill_2 FILLER_46_747 ();
 sg13g2_decap_8 FILLER_46_759 ();
 sg13g2_decap_8 FILLER_46_766 ();
 sg13g2_decap_4 FILLER_46_789 ();
 sg13g2_fill_1 FILLER_46_793 ();
 sg13g2_decap_8 FILLER_46_802 ();
 sg13g2_decap_4 FILLER_46_809 ();
 sg13g2_decap_8 FILLER_46_832 ();
 sg13g2_decap_4 FILLER_46_839 ();
 sg13g2_fill_1 FILLER_46_843 ();
 sg13g2_decap_8 FILLER_46_853 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_11 ();
 sg13g2_fill_1 FILLER_47_17 ();
 sg13g2_fill_2 FILLER_47_36 ();
 sg13g2_fill_1 FILLER_47_52 ();
 sg13g2_decap_8 FILLER_47_58 ();
 sg13g2_fill_2 FILLER_47_86 ();
 sg13g2_fill_1 FILLER_47_88 ();
 sg13g2_fill_2 FILLER_47_115 ();
 sg13g2_decap_4 FILLER_47_126 ();
 sg13g2_fill_2 FILLER_47_130 ();
 sg13g2_decap_8 FILLER_47_136 ();
 sg13g2_decap_8 FILLER_47_143 ();
 sg13g2_decap_8 FILLER_47_150 ();
 sg13g2_fill_1 FILLER_47_178 ();
 sg13g2_decap_4 FILLER_47_191 ();
 sg13g2_fill_1 FILLER_47_195 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_4 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_249 ();
 sg13g2_fill_2 FILLER_47_256 ();
 sg13g2_fill_1 FILLER_47_258 ();
 sg13g2_fill_2 FILLER_47_280 ();
 sg13g2_fill_1 FILLER_47_282 ();
 sg13g2_fill_1 FILLER_47_291 ();
 sg13g2_fill_1 FILLER_47_297 ();
 sg13g2_fill_2 FILLER_47_315 ();
 sg13g2_fill_2 FILLER_47_326 ();
 sg13g2_fill_2 FILLER_47_349 ();
 sg13g2_decap_8 FILLER_47_355 ();
 sg13g2_decap_8 FILLER_47_411 ();
 sg13g2_fill_2 FILLER_47_418 ();
 sg13g2_decap_8 FILLER_47_428 ();
 sg13g2_decap_8 FILLER_47_435 ();
 sg13g2_fill_1 FILLER_47_447 ();
 sg13g2_fill_1 FILLER_47_476 ();
 sg13g2_fill_1 FILLER_47_489 ();
 sg13g2_decap_4 FILLER_47_495 ();
 sg13g2_fill_1 FILLER_47_519 ();
 sg13g2_fill_2 FILLER_47_536 ();
 sg13g2_fill_1 FILLER_47_538 ();
 sg13g2_decap_8 FILLER_47_554 ();
 sg13g2_decap_4 FILLER_47_566 ();
 sg13g2_fill_1 FILLER_47_570 ();
 sg13g2_decap_8 FILLER_47_591 ();
 sg13g2_fill_1 FILLER_47_598 ();
 sg13g2_fill_1 FILLER_47_607 ();
 sg13g2_decap_4 FILLER_47_615 ();
 sg13g2_decap_4 FILLER_47_627 ();
 sg13g2_decap_4 FILLER_47_635 ();
 sg13g2_fill_1 FILLER_47_657 ();
 sg13g2_decap_4 FILLER_47_668 ();
 sg13g2_fill_2 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_703 ();
 sg13g2_decap_4 FILLER_47_721 ();
 sg13g2_fill_2 FILLER_47_754 ();
 sg13g2_fill_1 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_775 ();
 sg13g2_decap_8 FILLER_47_782 ();
 sg13g2_fill_1 FILLER_47_789 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_827 ();
 sg13g2_fill_2 FILLER_47_834 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_28 ();
 sg13g2_decap_4 FILLER_48_67 ();
 sg13g2_fill_1 FILLER_48_106 ();
 sg13g2_decap_8 FILLER_48_150 ();
 sg13g2_decap_8 FILLER_48_165 ();
 sg13g2_fill_2 FILLER_48_172 ();
 sg13g2_fill_2 FILLER_48_179 ();
 sg13g2_fill_1 FILLER_48_181 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_fill_2 FILLER_48_217 ();
 sg13g2_fill_1 FILLER_48_219 ();
 sg13g2_decap_4 FILLER_48_227 ();
 sg13g2_fill_1 FILLER_48_231 ();
 sg13g2_fill_2 FILLER_48_253 ();
 sg13g2_fill_2 FILLER_48_259 ();
 sg13g2_fill_1 FILLER_48_261 ();
 sg13g2_decap_8 FILLER_48_283 ();
 sg13g2_decap_4 FILLER_48_290 ();
 sg13g2_fill_1 FILLER_48_304 ();
 sg13g2_fill_2 FILLER_48_366 ();
 sg13g2_fill_1 FILLER_48_368 ();
 sg13g2_fill_2 FILLER_48_387 ();
 sg13g2_fill_2 FILLER_48_403 ();
 sg13g2_fill_1 FILLER_48_405 ();
 sg13g2_fill_1 FILLER_48_412 ();
 sg13g2_fill_2 FILLER_48_421 ();
 sg13g2_fill_1 FILLER_48_423 ();
 sg13g2_fill_1 FILLER_48_430 ();
 sg13g2_decap_8 FILLER_48_458 ();
 sg13g2_decap_4 FILLER_48_465 ();
 sg13g2_decap_4 FILLER_48_486 ();
 sg13g2_decap_8 FILLER_48_499 ();
 sg13g2_decap_8 FILLER_48_506 ();
 sg13g2_decap_8 FILLER_48_513 ();
 sg13g2_decap_4 FILLER_48_541 ();
 sg13g2_fill_1 FILLER_48_545 ();
 sg13g2_fill_2 FILLER_48_551 ();
 sg13g2_fill_1 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_559 ();
 sg13g2_decap_8 FILLER_48_566 ();
 sg13g2_decap_4 FILLER_48_573 ();
 sg13g2_fill_2 FILLER_48_587 ();
 sg13g2_fill_1 FILLER_48_589 ();
 sg13g2_fill_1 FILLER_48_596 ();
 sg13g2_fill_1 FILLER_48_605 ();
 sg13g2_fill_2 FILLER_48_614 ();
 sg13g2_decap_8 FILLER_48_650 ();
 sg13g2_decap_4 FILLER_48_666 ();
 sg13g2_fill_1 FILLER_48_670 ();
 sg13g2_decap_4 FILLER_48_677 ();
 sg13g2_fill_2 FILLER_48_681 ();
 sg13g2_decap_4 FILLER_48_698 ();
 sg13g2_fill_2 FILLER_48_702 ();
 sg13g2_decap_8 FILLER_48_709 ();
 sg13g2_fill_2 FILLER_48_716 ();
 sg13g2_decap_4 FILLER_48_727 ();
 sg13g2_fill_2 FILLER_48_731 ();
 sg13g2_fill_2 FILLER_48_738 ();
 sg13g2_decap_8 FILLER_48_745 ();
 sg13g2_decap_8 FILLER_48_752 ();
 sg13g2_fill_2 FILLER_48_759 ();
 sg13g2_fill_1 FILLER_48_761 ();
 sg13g2_decap_8 FILLER_48_780 ();
 sg13g2_fill_1 FILLER_48_787 ();
 sg13g2_fill_2 FILLER_48_809 ();
 sg13g2_fill_1 FILLER_48_811 ();
 sg13g2_fill_1 FILLER_48_818 ();
 sg13g2_fill_1 FILLER_48_824 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_fill_2 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_853 ();
 sg13g2_fill_2 FILLER_48_860 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_73 ();
 sg13g2_fill_2 FILLER_49_80 ();
 sg13g2_decap_4 FILLER_49_92 ();
 sg13g2_fill_1 FILLER_49_96 ();
 sg13g2_decap_4 FILLER_49_106 ();
 sg13g2_decap_4 FILLER_49_124 ();
 sg13g2_fill_2 FILLER_49_128 ();
 sg13g2_fill_2 FILLER_49_151 ();
 sg13g2_fill_1 FILLER_49_153 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_4 FILLER_49_182 ();
 sg13g2_fill_2 FILLER_49_186 ();
 sg13g2_decap_4 FILLER_49_209 ();
 sg13g2_fill_2 FILLER_49_213 ();
 sg13g2_fill_1 FILLER_49_253 ();
 sg13g2_fill_2 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_274 ();
 sg13g2_fill_2 FILLER_49_281 ();
 sg13g2_fill_1 FILLER_49_283 ();
 sg13g2_fill_2 FILLER_49_342 ();
 sg13g2_fill_2 FILLER_49_353 ();
 sg13g2_fill_1 FILLER_49_355 ();
 sg13g2_fill_1 FILLER_49_373 ();
 sg13g2_fill_1 FILLER_49_379 ();
 sg13g2_fill_2 FILLER_49_411 ();
 sg13g2_fill_1 FILLER_49_413 ();
 sg13g2_fill_2 FILLER_49_418 ();
 sg13g2_decap_8 FILLER_49_428 ();
 sg13g2_fill_2 FILLER_49_435 ();
 sg13g2_fill_1 FILLER_49_437 ();
 sg13g2_decap_8 FILLER_49_452 ();
 sg13g2_decap_8 FILLER_49_459 ();
 sg13g2_fill_1 FILLER_49_466 ();
 sg13g2_decap_8 FILLER_49_484 ();
 sg13g2_decap_4 FILLER_49_491 ();
 sg13g2_fill_2 FILLER_49_495 ();
 sg13g2_fill_2 FILLER_49_526 ();
 sg13g2_fill_1 FILLER_49_528 ();
 sg13g2_fill_2 FILLER_49_567 ();
 sg13g2_decap_4 FILLER_49_577 ();
 sg13g2_fill_1 FILLER_49_591 ();
 sg13g2_fill_2 FILLER_49_596 ();
 sg13g2_decap_4 FILLER_49_602 ();
 sg13g2_fill_1 FILLER_49_606 ();
 sg13g2_decap_8 FILLER_49_613 ();
 sg13g2_fill_1 FILLER_49_620 ();
 sg13g2_decap_8 FILLER_49_625 ();
 sg13g2_decap_4 FILLER_49_632 ();
 sg13g2_fill_2 FILLER_49_644 ();
 sg13g2_fill_1 FILLER_49_646 ();
 sg13g2_fill_1 FILLER_49_654 ();
 sg13g2_fill_1 FILLER_49_660 ();
 sg13g2_decap_4 FILLER_49_671 ();
 sg13g2_fill_1 FILLER_49_675 ();
 sg13g2_fill_1 FILLER_49_681 ();
 sg13g2_fill_2 FILLER_49_693 ();
 sg13g2_decap_4 FILLER_49_701 ();
 sg13g2_fill_1 FILLER_49_705 ();
 sg13g2_decap_4 FILLER_49_749 ();
 sg13g2_fill_1 FILLER_49_753 ();
 sg13g2_fill_1 FILLER_49_774 ();
 sg13g2_fill_2 FILLER_49_804 ();
 sg13g2_fill_1 FILLER_49_812 ();
 sg13g2_decap_4 FILLER_49_834 ();
 sg13g2_fill_1 FILLER_49_838 ();
 sg13g2_decap_4 FILLER_49_858 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_9 ();
 sg13g2_fill_1 FILLER_50_36 ();
 sg13g2_fill_1 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_74 ();
 sg13g2_decap_4 FILLER_50_81 ();
 sg13g2_fill_1 FILLER_50_85 ();
 sg13g2_decap_4 FILLER_50_102 ();
 sg13g2_decap_8 FILLER_50_118 ();
 sg13g2_fill_2 FILLER_50_125 ();
 sg13g2_decap_8 FILLER_50_148 ();
 sg13g2_decap_8 FILLER_50_155 ();
 sg13g2_decap_8 FILLER_50_162 ();
 sg13g2_fill_2 FILLER_50_169 ();
 sg13g2_decap_8 FILLER_50_192 ();
 sg13g2_decap_4 FILLER_50_199 ();
 sg13g2_decap_4 FILLER_50_211 ();
 sg13g2_fill_1 FILLER_50_219 ();
 sg13g2_decap_4 FILLER_50_225 ();
 sg13g2_decap_4 FILLER_50_250 ();
 sg13g2_fill_2 FILLER_50_254 ();
 sg13g2_fill_1 FILLER_50_260 ();
 sg13g2_decap_8 FILLER_50_274 ();
 sg13g2_decap_4 FILLER_50_281 ();
 sg13g2_fill_1 FILLER_50_285 ();
 sg13g2_decap_4 FILLER_50_299 ();
 sg13g2_fill_1 FILLER_50_303 ();
 sg13g2_fill_1 FILLER_50_353 ();
 sg13g2_fill_2 FILLER_50_392 ();
 sg13g2_fill_1 FILLER_50_394 ();
 sg13g2_fill_1 FILLER_50_421 ();
 sg13g2_decap_4 FILLER_50_436 ();
 sg13g2_decap_4 FILLER_50_460 ();
 sg13g2_fill_2 FILLER_50_487 ();
 sg13g2_decap_8 FILLER_50_508 ();
 sg13g2_fill_2 FILLER_50_515 ();
 sg13g2_fill_1 FILLER_50_517 ();
 sg13g2_decap_8 FILLER_50_523 ();
 sg13g2_decap_4 FILLER_50_530 ();
 sg13g2_fill_1 FILLER_50_534 ();
 sg13g2_decap_4 FILLER_50_540 ();
 sg13g2_fill_1 FILLER_50_544 ();
 sg13g2_decap_8 FILLER_50_560 ();
 sg13g2_fill_2 FILLER_50_567 ();
 sg13g2_fill_1 FILLER_50_569 ();
 sg13g2_decap_4 FILLER_50_575 ();
 sg13g2_fill_2 FILLER_50_579 ();
 sg13g2_decap_8 FILLER_50_589 ();
 sg13g2_decap_8 FILLER_50_596 ();
 sg13g2_fill_2 FILLER_50_603 ();
 sg13g2_fill_1 FILLER_50_621 ();
 sg13g2_decap_4 FILLER_50_627 ();
 sg13g2_decap_8 FILLER_50_644 ();
 sg13g2_fill_2 FILLER_50_651 ();
 sg13g2_fill_1 FILLER_50_658 ();
 sg13g2_fill_1 FILLER_50_669 ();
 sg13g2_decap_4 FILLER_50_678 ();
 sg13g2_fill_1 FILLER_50_682 ();
 sg13g2_decap_4 FILLER_50_695 ();
 sg13g2_fill_1 FILLER_50_699 ();
 sg13g2_decap_8 FILLER_50_708 ();
 sg13g2_decap_8 FILLER_50_715 ();
 sg13g2_fill_1 FILLER_50_722 ();
 sg13g2_decap_8 FILLER_50_732 ();
 sg13g2_fill_2 FILLER_50_747 ();
 sg13g2_decap_4 FILLER_50_759 ();
 sg13g2_fill_2 FILLER_50_763 ();
 sg13g2_fill_2 FILLER_50_769 ();
 sg13g2_fill_2 FILLER_50_776 ();
 sg13g2_fill_1 FILLER_50_778 ();
 sg13g2_decap_8 FILLER_50_790 ();
 sg13g2_fill_2 FILLER_50_802 ();
 sg13g2_decap_8 FILLER_50_815 ();
 sg13g2_decap_8 FILLER_50_831 ();
 sg13g2_decap_4 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_35 ();
 sg13g2_fill_2 FILLER_51_48 ();
 sg13g2_fill_1 FILLER_51_50 ();
 sg13g2_decap_8 FILLER_51_62 ();
 sg13g2_decap_8 FILLER_51_69 ();
 sg13g2_fill_1 FILLER_51_85 ();
 sg13g2_decap_8 FILLER_51_101 ();
 sg13g2_decap_8 FILLER_51_108 ();
 sg13g2_fill_1 FILLER_51_120 ();
 sg13g2_fill_2 FILLER_51_132 ();
 sg13g2_decap_4 FILLER_51_176 ();
 sg13g2_fill_2 FILLER_51_180 ();
 sg13g2_decap_4 FILLER_51_194 ();
 sg13g2_fill_2 FILLER_51_229 ();
 sg13g2_fill_2 FILLER_51_241 ();
 sg13g2_fill_1 FILLER_51_251 ();
 sg13g2_fill_1 FILLER_51_262 ();
 sg13g2_decap_8 FILLER_51_276 ();
 sg13g2_fill_2 FILLER_51_283 ();
 sg13g2_decap_4 FILLER_51_310 ();
 sg13g2_fill_1 FILLER_51_314 ();
 sg13g2_decap_4 FILLER_51_319 ();
 sg13g2_fill_1 FILLER_51_344 ();
 sg13g2_fill_1 FILLER_51_363 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_fill_1 FILLER_51_415 ();
 sg13g2_fill_1 FILLER_51_449 ();
 sg13g2_fill_2 FILLER_51_464 ();
 sg13g2_fill_1 FILLER_51_466 ();
 sg13g2_decap_8 FILLER_51_475 ();
 sg13g2_decap_8 FILLER_51_482 ();
 sg13g2_decap_4 FILLER_51_489 ();
 sg13g2_fill_2 FILLER_51_493 ();
 sg13g2_fill_2 FILLER_51_511 ();
 sg13g2_fill_1 FILLER_51_513 ();
 sg13g2_decap_4 FILLER_51_519 ();
 sg13g2_fill_1 FILLER_51_541 ();
 sg13g2_decap_4 FILLER_51_560 ();
 sg13g2_fill_2 FILLER_51_564 ();
 sg13g2_fill_1 FILLER_51_593 ();
 sg13g2_decap_8 FILLER_51_605 ();
 sg13g2_decap_4 FILLER_51_612 ();
 sg13g2_fill_1 FILLER_51_621 ();
 sg13g2_decap_8 FILLER_51_638 ();
 sg13g2_fill_2 FILLER_51_655 ();
 sg13g2_decap_8 FILLER_51_673 ();
 sg13g2_fill_2 FILLER_51_680 ();
 sg13g2_decap_4 FILLER_51_686 ();
 sg13g2_fill_2 FILLER_51_690 ();
 sg13g2_fill_2 FILLER_51_729 ();
 sg13g2_fill_2 FILLER_51_737 ();
 sg13g2_decap_4 FILLER_51_743 ();
 sg13g2_decap_8 FILLER_51_764 ();
 sg13g2_fill_2 FILLER_51_771 ();
 sg13g2_fill_2 FILLER_51_785 ();
 sg13g2_decap_8 FILLER_51_799 ();
 sg13g2_fill_1 FILLER_51_806 ();
 sg13g2_decap_8 FILLER_51_817 ();
 sg13g2_fill_2 FILLER_51_824 ();
 sg13g2_fill_1 FILLER_51_836 ();
 sg13g2_decap_8 FILLER_51_855 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_4 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_42 ();
 sg13g2_decap_4 FILLER_52_65 ();
 sg13g2_fill_2 FILLER_52_74 ();
 sg13g2_fill_1 FILLER_52_76 ();
 sg13g2_decap_4 FILLER_52_97 ();
 sg13g2_fill_1 FILLER_52_111 ();
 sg13g2_fill_2 FILLER_52_123 ();
 sg13g2_decap_4 FILLER_52_137 ();
 sg13g2_fill_1 FILLER_52_141 ();
 sg13g2_decap_8 FILLER_52_150 ();
 sg13g2_decap_8 FILLER_52_157 ();
 sg13g2_fill_2 FILLER_52_164 ();
 sg13g2_decap_8 FILLER_52_179 ();
 sg13g2_decap_8 FILLER_52_186 ();
 sg13g2_decap_8 FILLER_52_193 ();
 sg13g2_decap_4 FILLER_52_200 ();
 sg13g2_fill_2 FILLER_52_204 ();
 sg13g2_fill_1 FILLER_52_211 ();
 sg13g2_fill_1 FILLER_52_221 ();
 sg13g2_decap_8 FILLER_52_225 ();
 sg13g2_decap_4 FILLER_52_232 ();
 sg13g2_fill_1 FILLER_52_236 ();
 sg13g2_decap_8 FILLER_52_251 ();
 sg13g2_fill_2 FILLER_52_258 ();
 sg13g2_decap_4 FILLER_52_273 ();
 sg13g2_fill_1 FILLER_52_277 ();
 sg13g2_fill_2 FILLER_52_298 ();
 sg13g2_fill_1 FILLER_52_300 ();
 sg13g2_fill_1 FILLER_52_314 ();
 sg13g2_fill_1 FILLER_52_320 ();
 sg13g2_decap_4 FILLER_52_366 ();
 sg13g2_fill_1 FILLER_52_370 ();
 sg13g2_fill_2 FILLER_52_380 ();
 sg13g2_fill_1 FILLER_52_390 ();
 sg13g2_fill_1 FILLER_52_404 ();
 sg13g2_fill_1 FILLER_52_420 ();
 sg13g2_fill_2 FILLER_52_429 ();
 sg13g2_decap_4 FILLER_52_436 ();
 sg13g2_decap_4 FILLER_52_444 ();
 sg13g2_fill_2 FILLER_52_448 ();
 sg13g2_decap_8 FILLER_52_455 ();
 sg13g2_decap_4 FILLER_52_462 ();
 sg13g2_fill_2 FILLER_52_466 ();
 sg13g2_fill_2 FILLER_52_492 ();
 sg13g2_fill_1 FILLER_52_494 ();
 sg13g2_decap_4 FILLER_52_523 ();
 sg13g2_fill_2 FILLER_52_527 ();
 sg13g2_decap_8 FILLER_52_535 ();
 sg13g2_fill_2 FILLER_52_542 ();
 sg13g2_fill_2 FILLER_52_556 ();
 sg13g2_fill_1 FILLER_52_558 ();
 sg13g2_decap_8 FILLER_52_567 ();
 sg13g2_decap_8 FILLER_52_574 ();
 sg13g2_fill_2 FILLER_52_581 ();
 sg13g2_fill_1 FILLER_52_595 ();
 sg13g2_decap_8 FILLER_52_606 ();
 sg13g2_fill_2 FILLER_52_613 ();
 sg13g2_fill_1 FILLER_52_615 ();
 sg13g2_decap_8 FILLER_52_630 ();
 sg13g2_decap_4 FILLER_52_637 ();
 sg13g2_fill_2 FILLER_52_641 ();
 sg13g2_decap_4 FILLER_52_649 ();
 sg13g2_fill_2 FILLER_52_653 ();
 sg13g2_decap_4 FILLER_52_670 ();
 sg13g2_decap_4 FILLER_52_679 ();
 sg13g2_fill_1 FILLER_52_707 ();
 sg13g2_decap_8 FILLER_52_714 ();
 sg13g2_decap_8 FILLER_52_735 ();
 sg13g2_fill_1 FILLER_52_742 ();
 sg13g2_fill_1 FILLER_52_761 ();
 sg13g2_decap_8 FILLER_52_768 ();
 sg13g2_fill_2 FILLER_52_775 ();
 sg13g2_fill_1 FILLER_52_777 ();
 sg13g2_decap_4 FILLER_52_787 ();
 sg13g2_fill_2 FILLER_52_796 ();
 sg13g2_fill_1 FILLER_52_798 ();
 sg13g2_fill_2 FILLER_52_817 ();
 sg13g2_fill_1 FILLER_52_832 ();
 sg13g2_fill_2 FILLER_52_837 ();
 sg13g2_fill_1 FILLER_52_839 ();
 sg13g2_fill_1 FILLER_52_846 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_4 FILLER_53_7 ();
 sg13g2_fill_2 FILLER_53_11 ();
 sg13g2_fill_1 FILLER_53_16 ();
 sg13g2_fill_1 FILLER_53_38 ();
 sg13g2_decap_8 FILLER_53_48 ();
 sg13g2_decap_8 FILLER_53_55 ();
 sg13g2_decap_8 FILLER_53_62 ();
 sg13g2_decap_8 FILLER_53_69 ();
 sg13g2_decap_4 FILLER_53_76 ();
 sg13g2_decap_8 FILLER_53_99 ();
 sg13g2_fill_2 FILLER_53_106 ();
 sg13g2_decap_4 FILLER_53_114 ();
 sg13g2_fill_1 FILLER_53_123 ();
 sg13g2_fill_1 FILLER_53_141 ();
 sg13g2_decap_8 FILLER_53_153 ();
 sg13g2_fill_1 FILLER_53_202 ();
 sg13g2_fill_1 FILLER_53_222 ();
 sg13g2_decap_8 FILLER_53_228 ();
 sg13g2_fill_2 FILLER_53_235 ();
 sg13g2_fill_2 FILLER_53_249 ();
 sg13g2_fill_1 FILLER_53_251 ();
 sg13g2_decap_4 FILLER_53_257 ();
 sg13g2_decap_4 FILLER_53_276 ();
 sg13g2_fill_1 FILLER_53_280 ();
 sg13g2_decap_8 FILLER_53_294 ();
 sg13g2_fill_2 FILLER_53_301 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_357 ();
 sg13g2_decap_8 FILLER_53_391 ();
 sg13g2_decap_4 FILLER_53_398 ();
 sg13g2_decap_4 FILLER_53_416 ();
 sg13g2_fill_2 FILLER_53_420 ();
 sg13g2_decap_8 FILLER_53_433 ();
 sg13g2_decap_4 FILLER_53_440 ();
 sg13g2_fill_2 FILLER_53_444 ();
 sg13g2_decap_4 FILLER_53_466 ();
 sg13g2_decap_4 FILLER_53_487 ();
 sg13g2_decap_4 FILLER_53_501 ();
 sg13g2_fill_2 FILLER_53_505 ();
 sg13g2_fill_2 FILLER_53_521 ();
 sg13g2_decap_8 FILLER_53_533 ();
 sg13g2_decap_4 FILLER_53_540 ();
 sg13g2_fill_1 FILLER_53_544 ();
 sg13g2_fill_2 FILLER_53_571 ();
 sg13g2_fill_1 FILLER_53_573 ();
 sg13g2_fill_1 FILLER_53_578 ();
 sg13g2_decap_4 FILLER_53_584 ();
 sg13g2_fill_1 FILLER_53_588 ();
 sg13g2_decap_8 FILLER_53_594 ();
 sg13g2_fill_2 FILLER_53_601 ();
 sg13g2_decap_4 FILLER_53_608 ();
 sg13g2_decap_4 FILLER_53_620 ();
 sg13g2_fill_2 FILLER_53_624 ();
 sg13g2_fill_1 FILLER_53_647 ();
 sg13g2_fill_2 FILLER_53_652 ();
 sg13g2_decap_4 FILLER_53_673 ();
 sg13g2_fill_1 FILLER_53_677 ();
 sg13g2_decap_8 FILLER_53_694 ();
 sg13g2_decap_4 FILLER_53_701 ();
 sg13g2_decap_8 FILLER_53_710 ();
 sg13g2_decap_8 FILLER_53_717 ();
 sg13g2_fill_1 FILLER_53_724 ();
 sg13g2_decap_4 FILLER_53_746 ();
 sg13g2_fill_2 FILLER_53_750 ();
 sg13g2_decap_8 FILLER_53_767 ();
 sg13g2_fill_2 FILLER_53_774 ();
 sg13g2_fill_1 FILLER_53_776 ();
 sg13g2_decap_4 FILLER_53_800 ();
 sg13g2_fill_2 FILLER_53_804 ();
 sg13g2_decap_8 FILLER_53_820 ();
 sg13g2_fill_1 FILLER_53_827 ();
 sg13g2_decap_8 FILLER_53_853 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_27 ();
 sg13g2_fill_2 FILLER_54_45 ();
 sg13g2_fill_1 FILLER_54_47 ();
 sg13g2_decap_8 FILLER_54_53 ();
 sg13g2_decap_8 FILLER_54_60 ();
 sg13g2_fill_1 FILLER_54_87 ();
 sg13g2_fill_2 FILLER_54_98 ();
 sg13g2_fill_2 FILLER_54_111 ();
 sg13g2_decap_4 FILLER_54_141 ();
 sg13g2_decap_8 FILLER_54_161 ();
 sg13g2_decap_8 FILLER_54_168 ();
 sg13g2_decap_8 FILLER_54_175 ();
 sg13g2_decap_4 FILLER_54_182 ();
 sg13g2_fill_1 FILLER_54_186 ();
 sg13g2_decap_8 FILLER_54_195 ();
 sg13g2_decap_8 FILLER_54_202 ();
 sg13g2_fill_2 FILLER_54_209 ();
 sg13g2_fill_2 FILLER_54_216 ();
 sg13g2_fill_1 FILLER_54_218 ();
 sg13g2_fill_2 FILLER_54_228 ();
 sg13g2_fill_1 FILLER_54_230 ();
 sg13g2_decap_8 FILLER_54_249 ();
 sg13g2_fill_2 FILLER_54_256 ();
 sg13g2_fill_1 FILLER_54_258 ();
 sg13g2_decap_8 FILLER_54_267 ();
 sg13g2_decap_8 FILLER_54_318 ();
 sg13g2_fill_1 FILLER_54_325 ();
 sg13g2_fill_2 FILLER_54_346 ();
 sg13g2_fill_1 FILLER_54_348 ();
 sg13g2_decap_8 FILLER_54_367 ();
 sg13g2_fill_1 FILLER_54_374 ();
 sg13g2_decap_4 FILLER_54_382 ();
 sg13g2_decap_4 FILLER_54_404 ();
 sg13g2_fill_1 FILLER_54_419 ();
 sg13g2_decap_8 FILLER_54_445 ();
 sg13g2_decap_4 FILLER_54_472 ();
 sg13g2_decap_4 FILLER_54_481 ();
 sg13g2_fill_2 FILLER_54_490 ();
 sg13g2_fill_1 FILLER_54_492 ();
 sg13g2_decap_8 FILLER_54_503 ();
 sg13g2_fill_2 FILLER_54_510 ();
 sg13g2_fill_2 FILLER_54_522 ();
 sg13g2_fill_1 FILLER_54_524 ();
 sg13g2_fill_2 FILLER_54_539 ();
 sg13g2_decap_4 FILLER_54_547 ();
 sg13g2_decap_4 FILLER_54_562 ();
 sg13g2_fill_2 FILLER_54_566 ();
 sg13g2_decap_4 FILLER_54_573 ();
 sg13g2_fill_2 FILLER_54_577 ();
 sg13g2_decap_4 FILLER_54_591 ();
 sg13g2_decap_4 FILLER_54_601 ();
 sg13g2_fill_1 FILLER_54_605 ();
 sg13g2_fill_2 FILLER_54_624 ();
 sg13g2_decap_4 FILLER_54_631 ();
 sg13g2_fill_2 FILLER_54_635 ();
 sg13g2_fill_1 FILLER_54_643 ();
 sg13g2_fill_1 FILLER_54_695 ();
 sg13g2_decap_4 FILLER_54_705 ();
 sg13g2_fill_1 FILLER_54_709 ();
 sg13g2_decap_4 FILLER_54_718 ();
 sg13g2_fill_1 FILLER_54_722 ();
 sg13g2_decap_8 FILLER_54_737 ();
 sg13g2_decap_4 FILLER_54_744 ();
 sg13g2_decap_8 FILLER_54_766 ();
 sg13g2_fill_1 FILLER_54_773 ();
 sg13g2_fill_2 FILLER_54_779 ();
 sg13g2_decap_4 FILLER_54_789 ();
 sg13g2_decap_8 FILLER_54_801 ();
 sg13g2_fill_1 FILLER_54_808 ();
 sg13g2_decap_4 FILLER_54_821 ();
 sg13g2_decap_4 FILLER_54_846 ();
 sg13g2_decap_8 FILLER_54_855 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_9 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_fill_2 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_4 FILLER_55_77 ();
 sg13g2_fill_1 FILLER_55_81 ();
 sg13g2_decap_8 FILLER_55_88 ();
 sg13g2_decap_8 FILLER_55_95 ();
 sg13g2_decap_4 FILLER_55_102 ();
 sg13g2_fill_1 FILLER_55_106 ();
 sg13g2_decap_4 FILLER_55_110 ();
 sg13g2_fill_1 FILLER_55_114 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_4 FILLER_55_140 ();
 sg13g2_fill_1 FILLER_55_144 ();
 sg13g2_fill_1 FILLER_55_153 ();
 sg13g2_decap_8 FILLER_55_196 ();
 sg13g2_fill_1 FILLER_55_203 ();
 sg13g2_decap_4 FILLER_55_213 ();
 sg13g2_fill_2 FILLER_55_221 ();
 sg13g2_fill_2 FILLER_55_227 ();
 sg13g2_fill_1 FILLER_55_229 ();
 sg13g2_fill_2 FILLER_55_236 ();
 sg13g2_fill_1 FILLER_55_238 ();
 sg13g2_decap_8 FILLER_55_245 ();
 sg13g2_decap_4 FILLER_55_252 ();
 sg13g2_fill_2 FILLER_55_291 ();
 sg13g2_fill_1 FILLER_55_299 ();
 sg13g2_decap_8 FILLER_55_365 ();
 sg13g2_decap_8 FILLER_55_372 ();
 sg13g2_fill_2 FILLER_55_379 ();
 sg13g2_fill_1 FILLER_55_381 ();
 sg13g2_fill_2 FILLER_55_387 ();
 sg13g2_fill_1 FILLER_55_389 ();
 sg13g2_decap_8 FILLER_55_396 ();
 sg13g2_decap_4 FILLER_55_403 ();
 sg13g2_fill_1 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_55_413 ();
 sg13g2_decap_8 FILLER_55_420 ();
 sg13g2_decap_8 FILLER_55_427 ();
 sg13g2_decap_8 FILLER_55_438 ();
 sg13g2_decap_4 FILLER_55_445 ();
 sg13g2_fill_2 FILLER_55_449 ();
 sg13g2_fill_2 FILLER_55_492 ();
 sg13g2_fill_2 FILLER_55_502 ();
 sg13g2_fill_2 FILLER_55_530 ();
 sg13g2_fill_1 FILLER_55_532 ();
 sg13g2_fill_2 FILLER_55_558 ();
 sg13g2_fill_1 FILLER_55_560 ();
 sg13g2_fill_1 FILLER_55_567 ();
 sg13g2_fill_1 FILLER_55_587 ();
 sg13g2_decap_4 FILLER_55_593 ();
 sg13g2_fill_2 FILLER_55_597 ();
 sg13g2_fill_2 FILLER_55_611 ();
 sg13g2_fill_1 FILLER_55_613 ();
 sg13g2_fill_2 FILLER_55_620 ();
 sg13g2_decap_8 FILLER_55_633 ();
 sg13g2_decap_8 FILLER_55_640 ();
 sg13g2_fill_1 FILLER_55_647 ();
 sg13g2_decap_8 FILLER_55_652 ();
 sg13g2_fill_2 FILLER_55_659 ();
 sg13g2_decap_8 FILLER_55_668 ();
 sg13g2_decap_8 FILLER_55_675 ();
 sg13g2_decap_4 FILLER_55_682 ();
 sg13g2_fill_1 FILLER_55_686 ();
 sg13g2_decap_8 FILLER_55_696 ();
 sg13g2_decap_4 FILLER_55_708 ();
 sg13g2_fill_1 FILLER_55_712 ();
 sg13g2_decap_4 FILLER_55_718 ();
 sg13g2_fill_1 FILLER_55_733 ();
 sg13g2_decap_4 FILLER_55_760 ();
 sg13g2_fill_2 FILLER_55_764 ();
 sg13g2_decap_4 FILLER_55_774 ();
 sg13g2_fill_2 FILLER_55_786 ();
 sg13g2_fill_1 FILLER_55_793 ();
 sg13g2_decap_4 FILLER_55_799 ();
 sg13g2_fill_2 FILLER_55_803 ();
 sg13g2_decap_8 FILLER_55_822 ();
 sg13g2_fill_2 FILLER_55_829 ();
 sg13g2_fill_2 FILLER_55_835 ();
 sg13g2_decap_8 FILLER_55_855 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_7 ();
 sg13g2_decap_4 FILLER_56_32 ();
 sg13g2_fill_2 FILLER_56_36 ();
 sg13g2_fill_1 FILLER_56_43 ();
 sg13g2_decap_8 FILLER_56_104 ();
 sg13g2_fill_2 FILLER_56_121 ();
 sg13g2_fill_1 FILLER_56_123 ();
 sg13g2_fill_1 FILLER_56_133 ();
 sg13g2_decap_4 FILLER_56_167 ();
 sg13g2_fill_2 FILLER_56_171 ();
 sg13g2_decap_8 FILLER_56_177 ();
 sg13g2_fill_1 FILLER_56_184 ();
 sg13g2_decap_8 FILLER_56_190 ();
 sg13g2_fill_1 FILLER_56_197 ();
 sg13g2_fill_2 FILLER_56_224 ();
 sg13g2_decap_4 FILLER_56_258 ();
 sg13g2_fill_1 FILLER_56_262 ();
 sg13g2_fill_1 FILLER_56_280 ();
 sg13g2_fill_1 FILLER_56_313 ();
 sg13g2_fill_1 FILLER_56_318 ();
 sg13g2_fill_1 FILLER_56_338 ();
 sg13g2_decap_8 FILLER_56_356 ();
 sg13g2_decap_4 FILLER_56_363 ();
 sg13g2_fill_1 FILLER_56_367 ();
 sg13g2_fill_2 FILLER_56_388 ();
 sg13g2_fill_1 FILLER_56_390 ();
 sg13g2_fill_2 FILLER_56_397 ();
 sg13g2_fill_1 FILLER_56_399 ();
 sg13g2_fill_2 FILLER_56_426 ();
 sg13g2_decap_4 FILLER_56_459 ();
 sg13g2_fill_2 FILLER_56_463 ();
 sg13g2_decap_8 FILLER_56_475 ();
 sg13g2_decap_8 FILLER_56_482 ();
 sg13g2_decap_8 FILLER_56_489 ();
 sg13g2_fill_2 FILLER_56_496 ();
 sg13g2_fill_1 FILLER_56_498 ();
 sg13g2_decap_4 FILLER_56_509 ();
 sg13g2_fill_2 FILLER_56_513 ();
 sg13g2_fill_1 FILLER_56_524 ();
 sg13g2_fill_2 FILLER_56_533 ();
 sg13g2_decap_8 FILLER_56_541 ();
 sg13g2_decap_8 FILLER_56_552 ();
 sg13g2_decap_8 FILLER_56_567 ();
 sg13g2_fill_2 FILLER_56_574 ();
 sg13g2_decap_8 FILLER_56_601 ();
 sg13g2_decap_4 FILLER_56_608 ();
 sg13g2_fill_1 FILLER_56_620 ();
 sg13g2_decap_4 FILLER_56_625 ();
 sg13g2_fill_1 FILLER_56_633 ();
 sg13g2_fill_1 FILLER_56_645 ();
 sg13g2_fill_1 FILLER_56_657 ();
 sg13g2_fill_1 FILLER_56_663 ();
 sg13g2_fill_1 FILLER_56_679 ();
 sg13g2_fill_1 FILLER_56_700 ();
 sg13g2_fill_2 FILLER_56_719 ();
 sg13g2_decap_4 FILLER_56_737 ();
 sg13g2_fill_1 FILLER_56_741 ();
 sg13g2_decap_8 FILLER_56_754 ();
 sg13g2_decap_4 FILLER_56_770 ();
 sg13g2_decap_4 FILLER_56_780 ();
 sg13g2_fill_1 FILLER_56_784 ();
 sg13g2_fill_2 FILLER_56_789 ();
 sg13g2_decap_4 FILLER_56_798 ();
 sg13g2_fill_2 FILLER_56_802 ();
 sg13g2_fill_1 FILLER_56_814 ();
 sg13g2_fill_2 FILLER_56_828 ();
 sg13g2_fill_1 FILLER_56_847 ();
 sg13g2_decap_4 FILLER_56_856 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_20 ();
 sg13g2_fill_2 FILLER_57_28 ();
 sg13g2_fill_2 FILLER_57_36 ();
 sg13g2_fill_1 FILLER_57_38 ();
 sg13g2_decap_8 FILLER_57_47 ();
 sg13g2_fill_2 FILLER_57_65 ();
 sg13g2_fill_1 FILLER_57_67 ();
 sg13g2_decap_4 FILLER_57_73 ();
 sg13g2_fill_1 FILLER_57_77 ();
 sg13g2_decap_4 FILLER_57_88 ();
 sg13g2_decap_4 FILLER_57_96 ();
 sg13g2_fill_2 FILLER_57_116 ();
 sg13g2_decap_8 FILLER_57_130 ();
 sg13g2_decap_8 FILLER_57_137 ();
 sg13g2_fill_2 FILLER_57_144 ();
 sg13g2_decap_4 FILLER_57_156 ();
 sg13g2_fill_2 FILLER_57_160 ();
 sg13g2_fill_2 FILLER_57_193 ();
 sg13g2_fill_1 FILLER_57_195 ();
 sg13g2_decap_8 FILLER_57_201 ();
 sg13g2_fill_2 FILLER_57_208 ();
 sg13g2_fill_2 FILLER_57_218 ();
 sg13g2_fill_1 FILLER_57_220 ();
 sg13g2_decap_8 FILLER_57_224 ();
 sg13g2_fill_2 FILLER_57_236 ();
 sg13g2_fill_1 FILLER_57_238 ();
 sg13g2_fill_1 FILLER_57_253 ();
 sg13g2_fill_1 FILLER_57_327 ();
 sg13g2_decap_8 FILLER_57_368 ();
 sg13g2_fill_1 FILLER_57_375 ();
 sg13g2_decap_8 FILLER_57_393 ();
 sg13g2_decap_4 FILLER_57_400 ();
 sg13g2_decap_8 FILLER_57_415 ();
 sg13g2_decap_8 FILLER_57_422 ();
 sg13g2_fill_2 FILLER_57_429 ();
 sg13g2_fill_2 FILLER_57_439 ();
 sg13g2_fill_1 FILLER_57_441 ();
 sg13g2_fill_2 FILLER_57_452 ();
 sg13g2_fill_2 FILLER_57_471 ();
 sg13g2_fill_1 FILLER_57_473 ();
 sg13g2_fill_1 FILLER_57_483 ();
 sg13g2_fill_2 FILLER_57_514 ();
 sg13g2_fill_1 FILLER_57_516 ();
 sg13g2_decap_4 FILLER_57_536 ();
 sg13g2_fill_2 FILLER_57_540 ();
 sg13g2_fill_2 FILLER_57_569 ();
 sg13g2_fill_1 FILLER_57_571 ();
 sg13g2_decap_8 FILLER_57_586 ();
 sg13g2_fill_2 FILLER_57_593 ();
 sg13g2_fill_2 FILLER_57_600 ();
 sg13g2_fill_1 FILLER_57_602 ();
 sg13g2_decap_8 FILLER_57_613 ();
 sg13g2_fill_2 FILLER_57_643 ();
 sg13g2_fill_1 FILLER_57_645 ();
 sg13g2_decap_4 FILLER_57_659 ();
 sg13g2_fill_2 FILLER_57_663 ();
 sg13g2_decap_4 FILLER_57_670 ();
 sg13g2_fill_1 FILLER_57_674 ();
 sg13g2_fill_2 FILLER_57_681 ();
 sg13g2_decap_8 FILLER_57_691 ();
 sg13g2_decap_4 FILLER_57_698 ();
 sg13g2_fill_1 FILLER_57_702 ();
 sg13g2_decap_8 FILLER_57_707 ();
 sg13g2_fill_2 FILLER_57_714 ();
 sg13g2_decap_4 FILLER_57_722 ();
 sg13g2_fill_2 FILLER_57_726 ();
 sg13g2_decap_4 FILLER_57_736 ();
 sg13g2_fill_2 FILLER_57_740 ();
 sg13g2_decap_4 FILLER_57_748 ();
 sg13g2_fill_1 FILLER_57_752 ();
 sg13g2_decap_8 FILLER_57_764 ();
 sg13g2_fill_2 FILLER_57_771 ();
 sg13g2_decap_4 FILLER_57_789 ();
 sg13g2_fill_2 FILLER_57_793 ();
 sg13g2_decap_4 FILLER_57_805 ();
 sg13g2_fill_2 FILLER_57_809 ();
 sg13g2_decap_8 FILLER_57_821 ();
 sg13g2_decap_8 FILLER_57_828 ();
 sg13g2_fill_2 FILLER_57_835 ();
 sg13g2_decap_8 FILLER_57_854 ();
 sg13g2_fill_1 FILLER_57_861 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_7 ();
 sg13g2_decap_4 FILLER_58_48 ();
 sg13g2_decap_4 FILLER_58_57 ();
 sg13g2_decap_8 FILLER_58_66 ();
 sg13g2_fill_1 FILLER_58_73 ();
 sg13g2_fill_1 FILLER_58_80 ();
 sg13g2_decap_8 FILLER_58_97 ();
 sg13g2_fill_1 FILLER_58_104 ();
 sg13g2_decap_4 FILLER_58_109 ();
 sg13g2_fill_2 FILLER_58_113 ();
 sg13g2_decap_8 FILLER_58_124 ();
 sg13g2_decap_8 FILLER_58_131 ();
 sg13g2_fill_1 FILLER_58_138 ();
 sg13g2_fill_1 FILLER_58_144 ();
 sg13g2_decap_8 FILLER_58_156 ();
 sg13g2_decap_4 FILLER_58_163 ();
 sg13g2_fill_1 FILLER_58_167 ();
 sg13g2_fill_1 FILLER_58_185 ();
 sg13g2_fill_2 FILLER_58_269 ();
 sg13g2_fill_2 FILLER_58_290 ();
 sg13g2_fill_2 FILLER_58_319 ();
 sg13g2_fill_1 FILLER_58_321 ();
 sg13g2_fill_2 FILLER_58_337 ();
 sg13g2_fill_1 FILLER_58_339 ();
 sg13g2_fill_1 FILLER_58_353 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_decap_8 FILLER_58_382 ();
 sg13g2_fill_2 FILLER_58_389 ();
 sg13g2_decap_4 FILLER_58_423 ();
 sg13g2_fill_2 FILLER_58_427 ();
 sg13g2_fill_1 FILLER_58_437 ();
 sg13g2_decap_8 FILLER_58_444 ();
 sg13g2_decap_4 FILLER_58_471 ();
 sg13g2_decap_4 FILLER_58_480 ();
 sg13g2_fill_2 FILLER_58_489 ();
 sg13g2_fill_1 FILLER_58_491 ();
 sg13g2_decap_4 FILLER_58_512 ();
 sg13g2_fill_1 FILLER_58_516 ();
 sg13g2_decap_4 FILLER_58_526 ();
 sg13g2_decap_4 FILLER_58_535 ();
 sg13g2_fill_1 FILLER_58_539 ();
 sg13g2_fill_1 FILLER_58_548 ();
 sg13g2_decap_4 FILLER_58_558 ();
 sg13g2_fill_2 FILLER_58_562 ();
 sg13g2_fill_1 FILLER_58_569 ();
 sg13g2_fill_2 FILLER_58_575 ();
 sg13g2_fill_1 FILLER_58_577 ();
 sg13g2_fill_2 FILLER_58_593 ();
 sg13g2_decap_8 FILLER_58_609 ();
 sg13g2_decap_8 FILLER_58_616 ();
 sg13g2_decap_4 FILLER_58_623 ();
 sg13g2_fill_2 FILLER_58_627 ();
 sg13g2_decap_4 FILLER_58_648 ();
 sg13g2_fill_2 FILLER_58_652 ();
 sg13g2_fill_2 FILLER_58_660 ();
 sg13g2_fill_1 FILLER_58_662 ();
 sg13g2_decap_8 FILLER_58_668 ();
 sg13g2_decap_4 FILLER_58_680 ();
 sg13g2_fill_1 FILLER_58_684 ();
 sg13g2_fill_2 FILLER_58_697 ();
 sg13g2_fill_1 FILLER_58_699 ();
 sg13g2_decap_8 FILLER_58_724 ();
 sg13g2_fill_2 FILLER_58_731 ();
 sg13g2_fill_2 FILLER_58_743 ();
 sg13g2_fill_2 FILLER_58_766 ();
 sg13g2_fill_1 FILLER_58_768 ();
 sg13g2_decap_4 FILLER_58_788 ();
 sg13g2_fill_1 FILLER_58_828 ();
 sg13g2_fill_2 FILLER_58_848 ();
 sg13g2_decap_4 FILLER_58_858 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_32 ();
 sg13g2_fill_1 FILLER_59_39 ();
 sg13g2_fill_2 FILLER_59_45 ();
 sg13g2_decap_8 FILLER_59_66 ();
 sg13g2_fill_2 FILLER_59_73 ();
 sg13g2_fill_1 FILLER_59_75 ();
 sg13g2_decap_8 FILLER_59_118 ();
 sg13g2_fill_2 FILLER_59_125 ();
 sg13g2_decap_8 FILLER_59_148 ();
 sg13g2_fill_2 FILLER_59_155 ();
 sg13g2_fill_2 FILLER_59_183 ();
 sg13g2_fill_2 FILLER_59_241 ();
 sg13g2_fill_1 FILLER_59_243 ();
 sg13g2_decap_8 FILLER_59_254 ();
 sg13g2_decap_4 FILLER_59_261 ();
 sg13g2_fill_1 FILLER_59_265 ();
 sg13g2_fill_1 FILLER_59_302 ();
 sg13g2_fill_2 FILLER_59_388 ();
 sg13g2_fill_1 FILLER_59_404 ();
 sg13g2_decap_4 FILLER_59_415 ();
 sg13g2_fill_2 FILLER_59_429 ();
 sg13g2_decap_8 FILLER_59_437 ();
 sg13g2_decap_8 FILLER_59_444 ();
 sg13g2_fill_2 FILLER_59_451 ();
 sg13g2_fill_1 FILLER_59_459 ();
 sg13g2_decap_4 FILLER_59_483 ();
 sg13g2_fill_2 FILLER_59_493 ();
 sg13g2_decap_4 FILLER_59_503 ();
 sg13g2_fill_1 FILLER_59_507 ();
 sg13g2_decap_4 FILLER_59_533 ();
 sg13g2_fill_2 FILLER_59_549 ();
 sg13g2_decap_8 FILLER_59_559 ();
 sg13g2_decap_8 FILLER_59_566 ();
 sg13g2_fill_1 FILLER_59_573 ();
 sg13g2_decap_8 FILLER_59_582 ();
 sg13g2_decap_8 FILLER_59_589 ();
 sg13g2_decap_4 FILLER_59_596 ();
 sg13g2_fill_2 FILLER_59_620 ();
 sg13g2_fill_1 FILLER_59_622 ();
 sg13g2_decap_8 FILLER_59_631 ();
 sg13g2_fill_1 FILLER_59_638 ();
 sg13g2_fill_2 FILLER_59_647 ();
 sg13g2_decap_4 FILLER_59_658 ();
 sg13g2_decap_8 FILLER_59_678 ();
 sg13g2_decap_8 FILLER_59_696 ();
 sg13g2_decap_4 FILLER_59_703 ();
 sg13g2_fill_1 FILLER_59_707 ();
 sg13g2_fill_2 FILLER_59_719 ();
 sg13g2_fill_2 FILLER_59_729 ();
 sg13g2_fill_2 FILLER_59_744 ();
 sg13g2_fill_1 FILLER_59_746 ();
 sg13g2_fill_2 FILLER_59_751 ();
 sg13g2_decap_8 FILLER_59_763 ();
 sg13g2_fill_2 FILLER_59_770 ();
 sg13g2_fill_1 FILLER_59_772 ();
 sg13g2_decap_8 FILLER_59_786 ();
 sg13g2_decap_4 FILLER_59_793 ();
 sg13g2_fill_1 FILLER_59_797 ();
 sg13g2_fill_2 FILLER_59_808 ();
 sg13g2_fill_1 FILLER_59_810 ();
 sg13g2_decap_8 FILLER_59_820 ();
 sg13g2_fill_2 FILLER_59_827 ();
 sg13g2_decap_4 FILLER_59_846 ();
 sg13g2_decap_4 FILLER_59_858 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_fill_1 FILLER_60_31 ();
 sg13g2_decap_4 FILLER_60_61 ();
 sg13g2_decap_8 FILLER_60_92 ();
 sg13g2_fill_2 FILLER_60_99 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_fill_2 FILLER_60_112 ();
 sg13g2_fill_1 FILLER_60_114 ();
 sg13g2_fill_2 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_153 ();
 sg13g2_decap_4 FILLER_60_160 ();
 sg13g2_fill_1 FILLER_60_180 ();
 sg13g2_fill_1 FILLER_60_195 ();
 sg13g2_fill_2 FILLER_60_314 ();
 sg13g2_fill_1 FILLER_60_316 ();
 sg13g2_fill_2 FILLER_60_360 ();
 sg13g2_fill_1 FILLER_60_376 ();
 sg13g2_decap_8 FILLER_60_381 ();
 sg13g2_decap_8 FILLER_60_388 ();
 sg13g2_fill_1 FILLER_60_395 ();
 sg13g2_decap_4 FILLER_60_409 ();
 sg13g2_fill_2 FILLER_60_413 ();
 sg13g2_fill_2 FILLER_60_444 ();
 sg13g2_fill_1 FILLER_60_446 ();
 sg13g2_fill_1 FILLER_60_460 ();
 sg13g2_decap_4 FILLER_60_492 ();
 sg13g2_fill_2 FILLER_60_507 ();
 sg13g2_fill_1 FILLER_60_509 ();
 sg13g2_fill_2 FILLER_60_515 ();
 sg13g2_fill_1 FILLER_60_517 ();
 sg13g2_fill_2 FILLER_60_524 ();
 sg13g2_decap_4 FILLER_60_539 ();
 sg13g2_fill_2 FILLER_60_543 ();
 sg13g2_decap_8 FILLER_60_550 ();
 sg13g2_fill_2 FILLER_60_557 ();
 sg13g2_fill_1 FILLER_60_559 ();
 sg13g2_fill_2 FILLER_60_567 ();
 sg13g2_fill_1 FILLER_60_569 ();
 sg13g2_decap_4 FILLER_60_599 ();
 sg13g2_fill_1 FILLER_60_614 ();
 sg13g2_decap_8 FILLER_60_624 ();
 sg13g2_fill_2 FILLER_60_631 ();
 sg13g2_fill_1 FILLER_60_633 ();
 sg13g2_fill_2 FILLER_60_639 ();
 sg13g2_fill_1 FILLER_60_641 ();
 sg13g2_decap_8 FILLER_60_653 ();
 sg13g2_decap_8 FILLER_60_660 ();
 sg13g2_fill_1 FILLER_60_667 ();
 sg13g2_fill_1 FILLER_60_678 ();
 sg13g2_decap_4 FILLER_60_688 ();
 sg13g2_decap_8 FILLER_60_697 ();
 sg13g2_fill_2 FILLER_60_704 ();
 sg13g2_fill_2 FILLER_60_724 ();
 sg13g2_decap_4 FILLER_60_742 ();
 sg13g2_fill_2 FILLER_60_746 ();
 sg13g2_decap_4 FILLER_60_753 ();
 sg13g2_fill_2 FILLER_60_757 ();
 sg13g2_decap_4 FILLER_60_763 ();
 sg13g2_fill_2 FILLER_60_767 ();
 sg13g2_fill_2 FILLER_60_775 ();
 sg13g2_fill_1 FILLER_60_777 ();
 sg13g2_decap_8 FILLER_60_803 ();
 sg13g2_decap_4 FILLER_60_810 ();
 sg13g2_fill_1 FILLER_60_814 ();
 sg13g2_decap_8 FILLER_60_825 ();
 sg13g2_fill_1 FILLER_60_832 ();
 sg13g2_fill_1 FILLER_60_837 ();
 sg13g2_decap_8 FILLER_60_850 ();
 sg13g2_decap_4 FILLER_60_857 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_decap_4 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_4 ();
 sg13g2_decap_8 FILLER_61_26 ();
 sg13g2_fill_2 FILLER_61_33 ();
 sg13g2_decap_8 FILLER_61_55 ();
 sg13g2_decap_4 FILLER_61_62 ();
 sg13g2_fill_2 FILLER_61_66 ();
 sg13g2_fill_2 FILLER_61_86 ();
 sg13g2_fill_1 FILLER_61_88 ();
 sg13g2_fill_1 FILLER_61_114 ();
 sg13g2_decap_8 FILLER_61_127 ();
 sg13g2_decap_4 FILLER_61_134 ();
 sg13g2_fill_1 FILLER_61_138 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_fill_2 FILLER_61_168 ();
 sg13g2_fill_2 FILLER_61_186 ();
 sg13g2_decap_8 FILLER_61_206 ();
 sg13g2_fill_2 FILLER_61_213 ();
 sg13g2_fill_1 FILLER_61_224 ();
 sg13g2_fill_1 FILLER_61_230 ();
 sg13g2_fill_1 FILLER_61_239 ();
 sg13g2_fill_1 FILLER_61_258 ();
 sg13g2_decap_8 FILLER_61_336 ();
 sg13g2_fill_1 FILLER_61_343 ();
 sg13g2_decap_4 FILLER_61_392 ();
 sg13g2_fill_2 FILLER_61_396 ();
 sg13g2_decap_8 FILLER_61_406 ();
 sg13g2_decap_8 FILLER_61_413 ();
 sg13g2_fill_2 FILLER_61_420 ();
 sg13g2_fill_1 FILLER_61_422 ();
 sg13g2_decap_4 FILLER_61_437 ();
 sg13g2_fill_1 FILLER_61_441 ();
 sg13g2_decap_8 FILLER_61_464 ();
 sg13g2_decap_8 FILLER_61_471 ();
 sg13g2_decap_4 FILLER_61_478 ();
 sg13g2_fill_1 FILLER_61_482 ();
 sg13g2_fill_2 FILLER_61_487 ();
 sg13g2_decap_8 FILLER_61_495 ();
 sg13g2_decap_8 FILLER_61_502 ();
 sg13g2_fill_2 FILLER_61_513 ();
 sg13g2_decap_8 FILLER_61_521 ();
 sg13g2_fill_2 FILLER_61_528 ();
 sg13g2_decap_4 FILLER_61_549 ();
 sg13g2_fill_2 FILLER_61_553 ();
 sg13g2_decap_4 FILLER_61_559 ();
 sg13g2_fill_2 FILLER_61_563 ();
 sg13g2_decap_4 FILLER_61_573 ();
 sg13g2_fill_2 FILLER_61_577 ();
 sg13g2_decap_4 FILLER_61_588 ();
 sg13g2_fill_1 FILLER_61_592 ();
 sg13g2_decap_8 FILLER_61_605 ();
 sg13g2_fill_1 FILLER_61_612 ();
 sg13g2_fill_2 FILLER_61_626 ();
 sg13g2_fill_1 FILLER_61_628 ();
 sg13g2_fill_1 FILLER_61_648 ();
 sg13g2_decap_4 FILLER_61_653 ();
 sg13g2_fill_1 FILLER_61_667 ();
 sg13g2_decap_4 FILLER_61_680 ();
 sg13g2_fill_1 FILLER_61_684 ();
 sg13g2_decap_4 FILLER_61_696 ();
 sg13g2_decap_4 FILLER_61_713 ();
 sg13g2_fill_2 FILLER_61_717 ();
 sg13g2_fill_1 FILLER_61_734 ();
 sg13g2_decap_4 FILLER_61_752 ();
 sg13g2_decap_4 FILLER_61_783 ();
 sg13g2_fill_1 FILLER_61_791 ();
 sg13g2_decap_8 FILLER_61_802 ();
 sg13g2_fill_1 FILLER_61_809 ();
 sg13g2_fill_2 FILLER_61_833 ();
 sg13g2_fill_1 FILLER_61_835 ();
 sg13g2_fill_2 FILLER_61_859 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_11 ();
 sg13g2_decap_8 FILLER_62_30 ();
 sg13g2_fill_2 FILLER_62_37 ();
 sg13g2_decap_8 FILLER_62_44 ();
 sg13g2_fill_2 FILLER_62_51 ();
 sg13g2_decap_8 FILLER_62_62 ();
 sg13g2_decap_8 FILLER_62_69 ();
 sg13g2_decap_4 FILLER_62_76 ();
 sg13g2_fill_1 FILLER_62_80 ();
 sg13g2_decap_4 FILLER_62_89 ();
 sg13g2_decap_4 FILLER_62_105 ();
 sg13g2_fill_2 FILLER_62_109 ();
 sg13g2_decap_8 FILLER_62_117 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_4 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_152 ();
 sg13g2_decap_4 FILLER_62_159 ();
 sg13g2_decap_8 FILLER_62_202 ();
 sg13g2_decap_4 FILLER_62_209 ();
 sg13g2_fill_1 FILLER_62_233 ();
 sg13g2_decap_4 FILLER_62_253 ();
 sg13g2_decap_4 FILLER_62_261 ();
 sg13g2_fill_2 FILLER_62_268 ();
 sg13g2_decap_8 FILLER_62_275 ();
 sg13g2_fill_1 FILLER_62_282 ();
 sg13g2_decap_4 FILLER_62_287 ();
 sg13g2_fill_1 FILLER_62_291 ();
 sg13g2_decap_8 FILLER_62_327 ();
 sg13g2_decap_8 FILLER_62_334 ();
 sg13g2_fill_2 FILLER_62_341 ();
 sg13g2_fill_1 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_62_375 ();
 sg13g2_decap_4 FILLER_62_382 ();
 sg13g2_fill_2 FILLER_62_386 ();
 sg13g2_decap_8 FILLER_62_404 ();
 sg13g2_fill_2 FILLER_62_419 ();
 sg13g2_fill_2 FILLER_62_442 ();
 sg13g2_decap_8 FILLER_62_448 ();
 sg13g2_decap_4 FILLER_62_455 ();
 sg13g2_decap_4 FILLER_62_469 ();
 sg13g2_fill_2 FILLER_62_473 ();
 sg13g2_fill_2 FILLER_62_489 ();
 sg13g2_decap_8 FILLER_62_497 ();
 sg13g2_fill_1 FILLER_62_504 ();
 sg13g2_decap_4 FILLER_62_521 ();
 sg13g2_fill_2 FILLER_62_543 ();
 sg13g2_fill_1 FILLER_62_545 ();
 sg13g2_fill_2 FILLER_62_567 ();
 sg13g2_fill_1 FILLER_62_569 ();
 sg13g2_decap_4 FILLER_62_586 ();
 sg13g2_decap_4 FILLER_62_607 ();
 sg13g2_decap_8 FILLER_62_616 ();
 sg13g2_decap_4 FILLER_62_650 ();
 sg13g2_fill_2 FILLER_62_654 ();
 sg13g2_decap_4 FILLER_62_678 ();
 sg13g2_fill_1 FILLER_62_682 ();
 sg13g2_fill_2 FILLER_62_687 ();
 sg13g2_fill_2 FILLER_62_695 ();
 sg13g2_decap_8 FILLER_62_702 ();
 sg13g2_decap_8 FILLER_62_709 ();
 sg13g2_decap_8 FILLER_62_716 ();
 sg13g2_decap_4 FILLER_62_723 ();
 sg13g2_fill_2 FILLER_62_732 ();
 sg13g2_fill_1 FILLER_62_734 ();
 sg13g2_decap_8 FILLER_62_739 ();
 sg13g2_fill_2 FILLER_62_746 ();
 sg13g2_decap_4 FILLER_62_753 ();
 sg13g2_fill_1 FILLER_62_757 ();
 sg13g2_decap_8 FILLER_62_767 ();
 sg13g2_fill_1 FILLER_62_774 ();
 sg13g2_fill_2 FILLER_62_786 ();
 sg13g2_decap_4 FILLER_62_804 ();
 sg13g2_fill_2 FILLER_62_808 ();
 sg13g2_decap_8 FILLER_62_823 ();
 sg13g2_decap_4 FILLER_62_830 ();
 sg13g2_decap_8 FILLER_62_855 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_7 ();
 sg13g2_fill_2 FILLER_63_39 ();
 sg13g2_fill_1 FILLER_63_41 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_fill_2 FILLER_63_70 ();
 sg13g2_fill_1 FILLER_63_72 ();
 sg13g2_decap_8 FILLER_63_97 ();
 sg13g2_decap_4 FILLER_63_104 ();
 sg13g2_fill_1 FILLER_63_120 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_decap_4 FILLER_63_161 ();
 sg13g2_fill_2 FILLER_63_165 ();
 sg13g2_decap_8 FILLER_63_208 ();
 sg13g2_fill_2 FILLER_63_215 ();
 sg13g2_fill_1 FILLER_63_217 ();
 sg13g2_fill_1 FILLER_63_221 ();
 sg13g2_decap_4 FILLER_63_236 ();
 sg13g2_fill_1 FILLER_63_240 ();
 sg13g2_decap_4 FILLER_63_277 ();
 sg13g2_fill_1 FILLER_63_300 ();
 sg13g2_fill_2 FILLER_63_310 ();
 sg13g2_fill_1 FILLER_63_312 ();
 sg13g2_decap_8 FILLER_63_339 ();
 sg13g2_decap_4 FILLER_63_346 ();
 sg13g2_fill_2 FILLER_63_350 ();
 sg13g2_decap_4 FILLER_63_356 ();
 sg13g2_decap_4 FILLER_63_364 ();
 sg13g2_decap_4 FILLER_63_373 ();
 sg13g2_decap_4 FILLER_63_395 ();
 sg13g2_fill_1 FILLER_63_399 ();
 sg13g2_decap_4 FILLER_63_408 ();
 sg13g2_fill_1 FILLER_63_412 ();
 sg13g2_fill_2 FILLER_63_417 ();
 sg13g2_decap_8 FILLER_63_434 ();
 sg13g2_decap_4 FILLER_63_441 ();
 sg13g2_fill_2 FILLER_63_445 ();
 sg13g2_fill_1 FILLER_63_451 ();
 sg13g2_decap_8 FILLER_63_466 ();
 sg13g2_decap_4 FILLER_63_473 ();
 sg13g2_fill_1 FILLER_63_487 ();
 sg13g2_decap_8 FILLER_63_507 ();
 sg13g2_decap_4 FILLER_63_522 ();
 sg13g2_fill_2 FILLER_63_526 ();
 sg13g2_decap_8 FILLER_63_546 ();
 sg13g2_fill_2 FILLER_63_553 ();
 sg13g2_fill_1 FILLER_63_563 ();
 sg13g2_fill_1 FILLER_63_581 ();
 sg13g2_decap_8 FILLER_63_596 ();
 sg13g2_fill_2 FILLER_63_603 ();
 sg13g2_fill_1 FILLER_63_605 ();
 sg13g2_decap_8 FILLER_63_626 ();
 sg13g2_fill_2 FILLER_63_638 ();
 sg13g2_fill_1 FILLER_63_640 ();
 sg13g2_decap_8 FILLER_63_646 ();
 sg13g2_decap_4 FILLER_63_653 ();
 sg13g2_fill_1 FILLER_63_657 ();
 sg13g2_fill_2 FILLER_63_664 ();
 sg13g2_fill_2 FILLER_63_689 ();
 sg13g2_decap_4 FILLER_63_721 ();
 sg13g2_fill_2 FILLER_63_729 ();
 sg13g2_fill_2 FILLER_63_746 ();
 sg13g2_fill_1 FILLER_63_748 ();
 sg13g2_fill_2 FILLER_63_768 ();
 sg13g2_fill_1 FILLER_63_770 ();
 sg13g2_decap_8 FILLER_63_782 ();
 sg13g2_decap_4 FILLER_63_789 ();
 sg13g2_fill_2 FILLER_63_802 ();
 sg13g2_fill_1 FILLER_63_809 ();
 sg13g2_decap_8 FILLER_63_820 ();
 sg13g2_fill_1 FILLER_63_827 ();
 sg13g2_fill_1 FILLER_63_837 ();
 sg13g2_decap_8 FILLER_63_846 ();
 sg13g2_decap_8 FILLER_63_853 ();
 sg13g2_fill_2 FILLER_63_860 ();
 sg13g2_decap_4 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_4 ();
 sg13g2_fill_2 FILLER_64_28 ();
 sg13g2_fill_2 FILLER_64_38 ();
 sg13g2_fill_2 FILLER_64_58 ();
 sg13g2_fill_1 FILLER_64_60 ();
 sg13g2_decap_4 FILLER_64_71 ();
 sg13g2_decap_8 FILLER_64_88 ();
 sg13g2_fill_1 FILLER_64_95 ();
 sg13g2_decap_4 FILLER_64_116 ();
 sg13g2_fill_1 FILLER_64_120 ();
 sg13g2_fill_2 FILLER_64_135 ();
 sg13g2_decap_4 FILLER_64_141 ();
 sg13g2_fill_1 FILLER_64_145 ();
 sg13g2_decap_8 FILLER_64_160 ();
 sg13g2_fill_2 FILLER_64_200 ();
 sg13g2_decap_8 FILLER_64_206 ();
 sg13g2_fill_2 FILLER_64_213 ();
 sg13g2_fill_2 FILLER_64_233 ();
 sg13g2_fill_1 FILLER_64_235 ();
 sg13g2_decap_8 FILLER_64_255 ();
 sg13g2_decap_4 FILLER_64_262 ();
 sg13g2_fill_1 FILLER_64_283 ();
 sg13g2_decap_4 FILLER_64_320 ();
 sg13g2_decap_4 FILLER_64_328 ();
 sg13g2_fill_2 FILLER_64_332 ();
 sg13g2_decap_4 FILLER_64_368 ();
 sg13g2_decap_8 FILLER_64_388 ();
 sg13g2_decap_8 FILLER_64_395 ();
 sg13g2_fill_2 FILLER_64_402 ();
 sg13g2_fill_2 FILLER_64_420 ();
 sg13g2_fill_1 FILLER_64_422 ();
 sg13g2_decap_8 FILLER_64_428 ();
 sg13g2_decap_4 FILLER_64_435 ();
 sg13g2_fill_1 FILLER_64_439 ();
 sg13g2_decap_8 FILLER_64_466 ();
 sg13g2_fill_2 FILLER_64_473 ();
 sg13g2_fill_1 FILLER_64_480 ();
 sg13g2_fill_2 FILLER_64_490 ();
 sg13g2_fill_2 FILLER_64_497 ();
 sg13g2_fill_1 FILLER_64_499 ();
 sg13g2_decap_8 FILLER_64_518 ();
 sg13g2_decap_4 FILLER_64_525 ();
 sg13g2_fill_1 FILLER_64_529 ();
 sg13g2_decap_8 FILLER_64_553 ();
 sg13g2_fill_1 FILLER_64_560 ();
 sg13g2_decap_4 FILLER_64_566 ();
 sg13g2_fill_1 FILLER_64_590 ();
 sg13g2_decap_8 FILLER_64_610 ();
 sg13g2_fill_2 FILLER_64_617 ();
 sg13g2_fill_1 FILLER_64_619 ();
 sg13g2_decap_4 FILLER_64_629 ();
 sg13g2_decap_8 FILLER_64_659 ();
 sg13g2_fill_2 FILLER_64_666 ();
 sg13g2_fill_2 FILLER_64_673 ();
 sg13g2_decap_8 FILLER_64_680 ();
 sg13g2_decap_8 FILLER_64_687 ();
 sg13g2_fill_2 FILLER_64_694 ();
 sg13g2_fill_2 FILLER_64_709 ();
 sg13g2_fill_2 FILLER_64_715 ();
 sg13g2_fill_1 FILLER_64_717 ();
 sg13g2_decap_8 FILLER_64_733 ();
 sg13g2_decap_8 FILLER_64_740 ();
 sg13g2_fill_2 FILLER_64_747 ();
 sg13g2_decap_4 FILLER_64_767 ();
 sg13g2_fill_1 FILLER_64_771 ();
 sg13g2_decap_8 FILLER_64_790 ();
 sg13g2_fill_1 FILLER_64_797 ();
 sg13g2_fill_1 FILLER_64_806 ();
 sg13g2_fill_1 FILLER_64_820 ();
 sg13g2_fill_2 FILLER_64_829 ();
 sg13g2_decap_4 FILLER_64_858 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_11 ();
 sg13g2_decap_4 FILLER_65_24 ();
 sg13g2_fill_2 FILLER_65_34 ();
 sg13g2_fill_2 FILLER_65_44 ();
 sg13g2_fill_1 FILLER_65_46 ();
 sg13g2_fill_2 FILLER_65_61 ();
 sg13g2_fill_1 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_74 ();
 sg13g2_fill_2 FILLER_65_87 ();
 sg13g2_decap_8 FILLER_65_162 ();
 sg13g2_decap_8 FILLER_65_169 ();
 sg13g2_fill_1 FILLER_65_176 ();
 sg13g2_decap_8 FILLER_65_181 ();
 sg13g2_decap_8 FILLER_65_188 ();
 sg13g2_fill_2 FILLER_65_195 ();
 sg13g2_fill_1 FILLER_65_197 ();
 sg13g2_fill_1 FILLER_65_224 ();
 sg13g2_fill_2 FILLER_65_257 ();
 sg13g2_fill_1 FILLER_65_259 ();
 sg13g2_fill_2 FILLER_65_277 ();
 sg13g2_decap_4 FILLER_65_285 ();
 sg13g2_fill_1 FILLER_65_294 ();
 sg13g2_fill_2 FILLER_65_312 ();
 sg13g2_decap_4 FILLER_65_331 ();
 sg13g2_fill_1 FILLER_65_335 ();
 sg13g2_decap_4 FILLER_65_340 ();
 sg13g2_fill_1 FILLER_65_344 ();
 sg13g2_fill_2 FILLER_65_358 ();
 sg13g2_fill_2 FILLER_65_408 ();
 sg13g2_fill_1 FILLER_65_410 ();
 sg13g2_fill_1 FILLER_65_423 ();
 sg13g2_fill_2 FILLER_65_434 ();
 sg13g2_fill_1 FILLER_65_436 ();
 sg13g2_fill_1 FILLER_65_441 ();
 sg13g2_fill_2 FILLER_65_450 ();
 sg13g2_fill_2 FILLER_65_463 ();
 sg13g2_fill_1 FILLER_65_486 ();
 sg13g2_fill_2 FILLER_65_499 ();
 sg13g2_fill_1 FILLER_65_501 ();
 sg13g2_decap_8 FILLER_65_512 ();
 sg13g2_decap_4 FILLER_65_519 ();
 sg13g2_fill_1 FILLER_65_523 ();
 sg13g2_fill_1 FILLER_65_529 ();
 sg13g2_fill_1 FILLER_65_535 ();
 sg13g2_decap_4 FILLER_65_563 ();
 sg13g2_fill_1 FILLER_65_567 ();
 sg13g2_decap_8 FILLER_65_586 ();
 sg13g2_decap_4 FILLER_65_593 ();
 sg13g2_fill_2 FILLER_65_597 ();
 sg13g2_fill_2 FILLER_65_604 ();
 sg13g2_fill_1 FILLER_65_606 ();
 sg13g2_decap_8 FILLER_65_612 ();
 sg13g2_decap_4 FILLER_65_619 ();
 sg13g2_decap_4 FILLER_65_636 ();
 sg13g2_fill_1 FILLER_65_640 ();
 sg13g2_decap_4 FILLER_65_651 ();
 sg13g2_fill_2 FILLER_65_655 ();
 sg13g2_decap_8 FILLER_65_684 ();
 sg13g2_decap_4 FILLER_65_696 ();
 sg13g2_fill_2 FILLER_65_705 ();
 sg13g2_decap_4 FILLER_65_727 ();
 sg13g2_fill_2 FILLER_65_731 ();
 sg13g2_decap_8 FILLER_65_760 ();
 sg13g2_decap_4 FILLER_65_767 ();
 sg13g2_fill_1 FILLER_65_771 ();
 sg13g2_fill_2 FILLER_65_785 ();
 sg13g2_fill_1 FILLER_65_787 ();
 sg13g2_fill_2 FILLER_65_795 ();
 sg13g2_decap_4 FILLER_65_802 ();
 sg13g2_decap_4 FILLER_65_815 ();
 sg13g2_decap_4 FILLER_65_838 ();
 sg13g2_fill_1 FILLER_65_842 ();
 sg13g2_decap_8 FILLER_65_854 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_7 ();
 sg13g2_fill_1 FILLER_66_11 ();
 sg13g2_decap_4 FILLER_66_20 ();
 sg13g2_fill_2 FILLER_66_45 ();
 sg13g2_fill_1 FILLER_66_47 ();
 sg13g2_fill_2 FILLER_66_56 ();
 sg13g2_fill_1 FILLER_66_58 ();
 sg13g2_fill_2 FILLER_66_75 ();
 sg13g2_fill_1 FILLER_66_77 ();
 sg13g2_decap_4 FILLER_66_99 ();
 sg13g2_fill_2 FILLER_66_103 ();
 sg13g2_decap_8 FILLER_66_111 ();
 sg13g2_fill_2 FILLER_66_128 ();
 sg13g2_fill_1 FILLER_66_130 ();
 sg13g2_decap_8 FILLER_66_136 ();
 sg13g2_fill_1 FILLER_66_143 ();
 sg13g2_fill_1 FILLER_66_149 ();
 sg13g2_decap_8 FILLER_66_155 ();
 sg13g2_decap_4 FILLER_66_162 ();
 sg13g2_fill_1 FILLER_66_166 ();
 sg13g2_fill_1 FILLER_66_171 ();
 sg13g2_fill_1 FILLER_66_177 ();
 sg13g2_decap_8 FILLER_66_191 ();
 sg13g2_decap_8 FILLER_66_198 ();
 sg13g2_decap_4 FILLER_66_205 ();
 sg13g2_decap_4 FILLER_66_213 ();
 sg13g2_fill_2 FILLER_66_240 ();
 sg13g2_fill_1 FILLER_66_242 ();
 sg13g2_decap_8 FILLER_66_258 ();
 sg13g2_fill_2 FILLER_66_265 ();
 sg13g2_fill_1 FILLER_66_267 ();
 sg13g2_fill_2 FILLER_66_308 ();
 sg13g2_fill_2 FILLER_66_336 ();
 sg13g2_fill_1 FILLER_66_343 ();
 sg13g2_decap_8 FILLER_66_348 ();
 sg13g2_decap_8 FILLER_66_355 ();
 sg13g2_fill_2 FILLER_66_362 ();
 sg13g2_decap_8 FILLER_66_369 ();
 sg13g2_fill_1 FILLER_66_376 ();
 sg13g2_fill_1 FILLER_66_381 ();
 sg13g2_decap_8 FILLER_66_391 ();
 sg13g2_decap_4 FILLER_66_398 ();
 sg13g2_fill_1 FILLER_66_402 ();
 sg13g2_decap_8 FILLER_66_407 ();
 sg13g2_fill_2 FILLER_66_414 ();
 sg13g2_fill_1 FILLER_66_416 ();
 sg13g2_fill_2 FILLER_66_426 ();
 sg13g2_fill_1 FILLER_66_428 ();
 sg13g2_fill_2 FILLER_66_438 ();
 sg13g2_decap_8 FILLER_66_472 ();
 sg13g2_decap_8 FILLER_66_496 ();
 sg13g2_fill_2 FILLER_66_503 ();
 sg13g2_fill_1 FILLER_66_505 ();
 sg13g2_fill_2 FILLER_66_510 ();
 sg13g2_fill_1 FILLER_66_517 ();
 sg13g2_fill_2 FILLER_66_529 ();
 sg13g2_fill_1 FILLER_66_531 ();
 sg13g2_fill_1 FILLER_66_541 ();
 sg13g2_decap_8 FILLER_66_552 ();
 sg13g2_fill_2 FILLER_66_564 ();
 sg13g2_fill_1 FILLER_66_566 ();
 sg13g2_decap_4 FILLER_66_578 ();
 sg13g2_fill_2 FILLER_66_602 ();
 sg13g2_decap_8 FILLER_66_618 ();
 sg13g2_decap_8 FILLER_66_631 ();
 sg13g2_decap_8 FILLER_66_638 ();
 sg13g2_fill_1 FILLER_66_645 ();
 sg13g2_fill_2 FILLER_66_651 ();
 sg13g2_decap_4 FILLER_66_679 ();
 sg13g2_fill_2 FILLER_66_683 ();
 sg13g2_decap_8 FILLER_66_702 ();
 sg13g2_fill_2 FILLER_66_709 ();
 sg13g2_fill_1 FILLER_66_711 ();
 sg13g2_fill_1 FILLER_66_716 ();
 sg13g2_decap_8 FILLER_66_727 ();
 sg13g2_decap_8 FILLER_66_734 ();
 sg13g2_fill_1 FILLER_66_741 ();
 sg13g2_decap_8 FILLER_66_756 ();
 sg13g2_decap_4 FILLER_66_763 ();
 sg13g2_fill_1 FILLER_66_767 ();
 sg13g2_decap_8 FILLER_66_773 ();
 sg13g2_fill_1 FILLER_66_780 ();
 sg13g2_fill_1 FILLER_66_794 ();
 sg13g2_fill_2 FILLER_66_800 ();
 sg13g2_decap_8 FILLER_66_808 ();
 sg13g2_fill_2 FILLER_66_815 ();
 sg13g2_decap_8 FILLER_66_826 ();
 sg13g2_decap_8 FILLER_66_833 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_7 ();
 sg13g2_decap_4 FILLER_67_69 ();
 sg13g2_decap_4 FILLER_67_110 ();
 sg13g2_decap_8 FILLER_67_118 ();
 sg13g2_decap_4 FILLER_67_135 ();
 sg13g2_fill_2 FILLER_67_139 ();
 sg13g2_fill_2 FILLER_67_215 ();
 sg13g2_fill_1 FILLER_67_217 ();
 sg13g2_fill_2 FILLER_67_228 ();
 sg13g2_fill_1 FILLER_67_230 ();
 sg13g2_fill_2 FILLER_67_277 ();
 sg13g2_decap_8 FILLER_67_288 ();
 sg13g2_decap_4 FILLER_67_295 ();
 sg13g2_fill_1 FILLER_67_299 ();
 sg13g2_fill_2 FILLER_67_309 ();
 sg13g2_fill_1 FILLER_67_311 ();
 sg13g2_fill_2 FILLER_67_330 ();
 sg13g2_fill_1 FILLER_67_332 ();
 sg13g2_decap_8 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_67_371 ();
 sg13g2_decap_4 FILLER_67_378 ();
 sg13g2_decap_4 FILLER_67_390 ();
 sg13g2_decap_8 FILLER_67_399 ();
 sg13g2_fill_2 FILLER_67_406 ();
 sg13g2_fill_1 FILLER_67_424 ();
 sg13g2_decap_8 FILLER_67_430 ();
 sg13g2_fill_2 FILLER_67_437 ();
 sg13g2_fill_1 FILLER_67_439 ();
 sg13g2_fill_2 FILLER_67_453 ();
 sg13g2_decap_8 FILLER_67_464 ();
 sg13g2_fill_2 FILLER_67_471 ();
 sg13g2_fill_1 FILLER_67_473 ();
 sg13g2_fill_2 FILLER_67_484 ();
 sg13g2_decap_4 FILLER_67_498 ();
 sg13g2_fill_1 FILLER_67_507 ();
 sg13g2_fill_2 FILLER_67_521 ();
 sg13g2_fill_1 FILLER_67_523 ();
 sg13g2_decap_4 FILLER_67_535 ();
 sg13g2_fill_1 FILLER_67_539 ();
 sg13g2_fill_2 FILLER_67_567 ();
 sg13g2_decap_8 FILLER_67_595 ();
 sg13g2_decap_4 FILLER_67_602 ();
 sg13g2_fill_1 FILLER_67_606 ();
 sg13g2_fill_1 FILLER_67_611 ();
 sg13g2_decap_8 FILLER_67_620 ();
 sg13g2_fill_1 FILLER_67_627 ();
 sg13g2_fill_1 FILLER_67_642 ();
 sg13g2_decap_4 FILLER_67_649 ();
 sg13g2_fill_1 FILLER_67_653 ();
 sg13g2_decap_4 FILLER_67_660 ();
 sg13g2_decap_8 FILLER_67_676 ();
 sg13g2_fill_2 FILLER_67_683 ();
 sg13g2_decap_8 FILLER_67_690 ();
 sg13g2_fill_2 FILLER_67_697 ();
 sg13g2_decap_8 FILLER_67_717 ();
 sg13g2_decap_4 FILLER_67_724 ();
 sg13g2_fill_1 FILLER_67_734 ();
 sg13g2_decap_4 FILLER_67_753 ();
 sg13g2_fill_1 FILLER_67_774 ();
 sg13g2_fill_2 FILLER_67_789 ();
 sg13g2_decap_8 FILLER_67_797 ();
 sg13g2_fill_2 FILLER_67_804 ();
 sg13g2_decap_4 FILLER_67_816 ();
 sg13g2_fill_2 FILLER_67_820 ();
 sg13g2_fill_2 FILLER_67_832 ();
 sg13g2_fill_1 FILLER_67_834 ();
 sg13g2_decap_4 FILLER_67_858 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_27 ();
 sg13g2_decap_8 FILLER_68_34 ();
 sg13g2_decap_4 FILLER_68_41 ();
 sg13g2_fill_1 FILLER_68_45 ();
 sg13g2_decap_8 FILLER_68_52 ();
 sg13g2_fill_2 FILLER_68_59 ();
 sg13g2_fill_1 FILLER_68_61 ();
 sg13g2_decap_4 FILLER_68_96 ();
 sg13g2_fill_2 FILLER_68_100 ();
 sg13g2_fill_2 FILLER_68_111 ();
 sg13g2_fill_1 FILLER_68_113 ();
 sg13g2_fill_1 FILLER_68_129 ();
 sg13g2_decap_4 FILLER_68_139 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_fill_2 FILLER_68_154 ();
 sg13g2_fill_1 FILLER_68_156 ();
 sg13g2_fill_1 FILLER_68_193 ();
 sg13g2_fill_2 FILLER_68_203 ();
 sg13g2_fill_1 FILLER_68_205 ();
 sg13g2_fill_1 FILLER_68_232 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_decap_8 FILLER_68_277 ();
 sg13g2_decap_4 FILLER_68_284 ();
 sg13g2_fill_2 FILLER_68_288 ();
 sg13g2_fill_1 FILLER_68_321 ();
 sg13g2_fill_2 FILLER_68_391 ();
 sg13g2_fill_1 FILLER_68_393 ();
 sg13g2_fill_2 FILLER_68_410 ();
 sg13g2_fill_2 FILLER_68_423 ();
 sg13g2_fill_1 FILLER_68_425 ();
 sg13g2_decap_8 FILLER_68_441 ();
 sg13g2_fill_2 FILLER_68_448 ();
 sg13g2_fill_1 FILLER_68_450 ();
 sg13g2_decap_4 FILLER_68_455 ();
 sg13g2_fill_2 FILLER_68_459 ();
 sg13g2_decap_4 FILLER_68_470 ();
 sg13g2_fill_2 FILLER_68_474 ();
 sg13g2_fill_2 FILLER_68_481 ();
 sg13g2_fill_1 FILLER_68_483 ();
 sg13g2_decap_8 FILLER_68_494 ();
 sg13g2_decap_8 FILLER_68_501 ();
 sg13g2_decap_4 FILLER_68_508 ();
 sg13g2_fill_2 FILLER_68_512 ();
 sg13g2_fill_1 FILLER_68_519 ();
 sg13g2_decap_4 FILLER_68_525 ();
 sg13g2_fill_1 FILLER_68_529 ();
 sg13g2_fill_2 FILLER_68_535 ();
 sg13g2_decap_4 FILLER_68_542 ();
 sg13g2_decap_8 FILLER_68_551 ();
 sg13g2_decap_4 FILLER_68_558 ();
 sg13g2_fill_2 FILLER_68_562 ();
 sg13g2_fill_1 FILLER_68_568 ();
 sg13g2_decap_8 FILLER_68_572 ();
 sg13g2_decap_8 FILLER_68_584 ();
 sg13g2_decap_4 FILLER_68_591 ();
 sg13g2_fill_2 FILLER_68_595 ();
 sg13g2_fill_2 FILLER_68_615 ();
 sg13g2_fill_1 FILLER_68_617 ();
 sg13g2_decap_4 FILLER_68_628 ();
 sg13g2_fill_2 FILLER_68_637 ();
 sg13g2_fill_1 FILLER_68_639 ();
 sg13g2_decap_8 FILLER_68_657 ();
 sg13g2_fill_2 FILLER_68_664 ();
 sg13g2_decap_4 FILLER_68_676 ();
 sg13g2_fill_1 FILLER_68_685 ();
 sg13g2_fill_2 FILLER_68_710 ();
 sg13g2_fill_1 FILLER_68_712 ();
 sg13g2_fill_2 FILLER_68_719 ();
 sg13g2_decap_4 FILLER_68_734 ();
 sg13g2_fill_1 FILLER_68_738 ();
 sg13g2_decap_8 FILLER_68_744 ();
 sg13g2_decap_8 FILLER_68_751 ();
 sg13g2_fill_2 FILLER_68_758 ();
 sg13g2_fill_2 FILLER_68_765 ();
 sg13g2_fill_1 FILLER_68_777 ();
 sg13g2_fill_1 FILLER_68_789 ();
 sg13g2_decap_4 FILLER_68_806 ();
 sg13g2_decap_4 FILLER_68_834 ();
 sg13g2_decap_4 FILLER_68_856 ();
 sg13g2_fill_2 FILLER_68_860 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_33 ();
 sg13g2_fill_2 FILLER_69_40 ();
 sg13g2_decap_8 FILLER_69_72 ();
 sg13g2_decap_8 FILLER_69_79 ();
 sg13g2_fill_1 FILLER_69_86 ();
 sg13g2_fill_2 FILLER_69_122 ();
 sg13g2_fill_2 FILLER_69_206 ();
 sg13g2_decap_8 FILLER_69_294 ();
 sg13g2_decap_4 FILLER_69_305 ();
 sg13g2_decap_4 FILLER_69_313 ();
 sg13g2_fill_2 FILLER_69_343 ();
 sg13g2_decap_8 FILLER_69_349 ();
 sg13g2_decap_8 FILLER_69_356 ();
 sg13g2_decap_4 FILLER_69_367 ();
 sg13g2_fill_1 FILLER_69_371 ();
 sg13g2_fill_2 FILLER_69_376 ();
 sg13g2_decap_8 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_69_398 ();
 sg13g2_decap_8 FILLER_69_417 ();
 sg13g2_fill_2 FILLER_69_424 ();
 sg13g2_fill_1 FILLER_69_432 ();
 sg13g2_fill_2 FILLER_69_466 ();
 sg13g2_fill_1 FILLER_69_468 ();
 sg13g2_fill_2 FILLER_69_495 ();
 sg13g2_fill_2 FILLER_69_546 ();
 sg13g2_fill_1 FILLER_69_548 ();
 sg13g2_fill_1 FILLER_69_555 ();
 sg13g2_fill_2 FILLER_69_579 ();
 sg13g2_decap_4 FILLER_69_587 ();
 sg13g2_fill_1 FILLER_69_591 ();
 sg13g2_decap_8 FILLER_69_617 ();
 sg13g2_decap_4 FILLER_69_624 ();
 sg13g2_fill_1 FILLER_69_628 ();
 sg13g2_fill_2 FILLER_69_637 ();
 sg13g2_fill_1 FILLER_69_639 ();
 sg13g2_decap_8 FILLER_69_645 ();
 sg13g2_fill_2 FILLER_69_652 ();
 sg13g2_decap_4 FILLER_69_658 ();
 sg13g2_fill_1 FILLER_69_667 ();
 sg13g2_decap_4 FILLER_69_680 ();
 sg13g2_decap_8 FILLER_69_695 ();
 sg13g2_decap_4 FILLER_69_702 ();
 sg13g2_fill_2 FILLER_69_712 ();
 sg13g2_fill_1 FILLER_69_714 ();
 sg13g2_fill_1 FILLER_69_751 ();
 sg13g2_fill_2 FILLER_69_775 ();
 sg13g2_decap_8 FILLER_69_792 ();
 sg13g2_decap_4 FILLER_69_799 ();
 sg13g2_fill_1 FILLER_69_821 ();
 sg13g2_decap_8 FILLER_69_826 ();
 sg13g2_decap_4 FILLER_69_833 ();
 sg13g2_fill_1 FILLER_69_837 ();
 sg13g2_decap_8 FILLER_69_843 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_11 ();
 sg13g2_fill_2 FILLER_70_16 ();
 sg13g2_fill_2 FILLER_70_22 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_fill_1 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_66 ();
 sg13g2_decap_8 FILLER_70_73 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_fill_1 FILLER_70_91 ();
 sg13g2_fill_2 FILLER_70_105 ();
 sg13g2_fill_1 FILLER_70_107 ();
 sg13g2_fill_1 FILLER_70_128 ();
 sg13g2_fill_2 FILLER_70_143 ();
 sg13g2_fill_1 FILLER_70_145 ();
 sg13g2_fill_1 FILLER_70_161 ();
 sg13g2_fill_2 FILLER_70_185 ();
 sg13g2_fill_1 FILLER_70_187 ();
 sg13g2_fill_2 FILLER_70_208 ();
 sg13g2_decap_8 FILLER_70_275 ();
 sg13g2_decap_8 FILLER_70_290 ();
 sg13g2_fill_1 FILLER_70_297 ();
 sg13g2_fill_1 FILLER_70_324 ();
 sg13g2_fill_2 FILLER_70_347 ();
 sg13g2_decap_8 FILLER_70_363 ();
 sg13g2_fill_2 FILLER_70_370 ();
 sg13g2_fill_1 FILLER_70_380 ();
 sg13g2_decap_8 FILLER_70_386 ();
 sg13g2_decap_8 FILLER_70_393 ();
 sg13g2_fill_2 FILLER_70_400 ();
 sg13g2_fill_2 FILLER_70_422 ();
 sg13g2_decap_4 FILLER_70_438 ();
 sg13g2_fill_1 FILLER_70_442 ();
 sg13g2_decap_8 FILLER_70_447 ();
 sg13g2_fill_1 FILLER_70_454 ();
 sg13g2_decap_8 FILLER_70_472 ();
 sg13g2_decap_4 FILLER_70_484 ();
 sg13g2_decap_8 FILLER_70_509 ();
 sg13g2_fill_1 FILLER_70_516 ();
 sg13g2_decap_8 FILLER_70_531 ();
 sg13g2_fill_2 FILLER_70_538 ();
 sg13g2_decap_8 FILLER_70_551 ();
 sg13g2_decap_8 FILLER_70_558 ();
 sg13g2_decap_4 FILLER_70_565 ();
 sg13g2_fill_2 FILLER_70_569 ();
 sg13g2_fill_1 FILLER_70_587 ();
 sg13g2_decap_8 FILLER_70_593 ();
 sg13g2_fill_2 FILLER_70_600 ();
 sg13g2_decap_8 FILLER_70_608 ();
 sg13g2_fill_1 FILLER_70_615 ();
 sg13g2_fill_2 FILLER_70_639 ();
 sg13g2_fill_1 FILLER_70_641 ();
 sg13g2_fill_1 FILLER_70_648 ();
 sg13g2_decap_8 FILLER_70_682 ();
 sg13g2_fill_2 FILLER_70_689 ();
 sg13g2_decap_8 FILLER_70_706 ();
 sg13g2_decap_8 FILLER_70_713 ();
 sg13g2_decap_4 FILLER_70_725 ();
 sg13g2_decap_4 FILLER_70_737 ();
 sg13g2_fill_1 FILLER_70_741 ();
 sg13g2_decap_8 FILLER_70_748 ();
 sg13g2_fill_2 FILLER_70_755 ();
 sg13g2_fill_1 FILLER_70_757 ();
 sg13g2_decap_4 FILLER_70_764 ();
 sg13g2_fill_1 FILLER_70_768 ();
 sg13g2_fill_2 FILLER_70_778 ();
 sg13g2_fill_1 FILLER_70_780 ();
 sg13g2_fill_2 FILLER_70_786 ();
 sg13g2_fill_1 FILLER_70_788 ();
 sg13g2_fill_1 FILLER_70_801 ();
 sg13g2_fill_2 FILLER_70_807 ();
 sg13g2_fill_1 FILLER_70_809 ();
 sg13g2_fill_2 FILLER_70_838 ();
 sg13g2_fill_1 FILLER_70_840 ();
 sg13g2_decap_4 FILLER_70_857 ();
 sg13g2_fill_1 FILLER_70_861 ();
 sg13g2_fill_1 FILLER_71_26 ();
 sg13g2_decap_4 FILLER_71_53 ();
 sg13g2_fill_2 FILLER_71_68 ();
 sg13g2_decap_8 FILLER_71_74 ();
 sg13g2_decap_4 FILLER_71_81 ();
 sg13g2_fill_2 FILLER_71_111 ();
 sg13g2_fill_1 FILLER_71_127 ();
 sg13g2_fill_1 FILLER_71_141 ();
 sg13g2_fill_1 FILLER_71_151 ();
 sg13g2_fill_1 FILLER_71_182 ();
 sg13g2_fill_2 FILLER_71_204 ();
 sg13g2_decap_4 FILLER_71_218 ();
 sg13g2_fill_1 FILLER_71_222 ();
 sg13g2_fill_1 FILLER_71_236 ();
 sg13g2_decap_4 FILLER_71_254 ();
 sg13g2_fill_2 FILLER_71_274 ();
 sg13g2_decap_8 FILLER_71_307 ();
 sg13g2_fill_1 FILLER_71_314 ();
 sg13g2_fill_2 FILLER_71_355 ();
 sg13g2_fill_2 FILLER_71_390 ();
 sg13g2_fill_1 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_408 ();
 sg13g2_fill_2 FILLER_71_415 ();
 sg13g2_fill_1 FILLER_71_417 ();
 sg13g2_fill_2 FILLER_71_440 ();
 sg13g2_fill_1 FILLER_71_442 ();
 sg13g2_fill_1 FILLER_71_455 ();
 sg13g2_decap_8 FILLER_71_461 ();
 sg13g2_decap_4 FILLER_71_468 ();
 sg13g2_fill_1 FILLER_71_472 ();
 sg13g2_decap_4 FILLER_71_478 ();
 sg13g2_fill_2 FILLER_71_482 ();
 sg13g2_decap_8 FILLER_71_498 ();
 sg13g2_decap_4 FILLER_71_505 ();
 sg13g2_fill_2 FILLER_71_530 ();
 sg13g2_decap_8 FILLER_71_544 ();
 sg13g2_fill_1 FILLER_71_551 ();
 sg13g2_fill_1 FILLER_71_557 ();
 sg13g2_decap_8 FILLER_71_564 ();
 sg13g2_decap_4 FILLER_71_571 ();
 sg13g2_fill_2 FILLER_71_575 ();
 sg13g2_decap_4 FILLER_71_600 ();
 sg13g2_fill_2 FILLER_71_604 ();
 sg13g2_fill_2 FILLER_71_618 ();
 sg13g2_fill_2 FILLER_71_637 ();
 sg13g2_fill_1 FILLER_71_639 ();
 sg13g2_decap_8 FILLER_71_645 ();
 sg13g2_decap_8 FILLER_71_657 ();
 sg13g2_decap_8 FILLER_71_680 ();
 sg13g2_fill_2 FILLER_71_687 ();
 sg13g2_fill_1 FILLER_71_689 ();
 sg13g2_fill_2 FILLER_71_698 ();
 sg13g2_decap_4 FILLER_71_716 ();
 sg13g2_fill_1 FILLER_71_720 ();
 sg13g2_fill_2 FILLER_71_726 ();
 sg13g2_fill_1 FILLER_71_738 ();
 sg13g2_fill_2 FILLER_71_745 ();
 sg13g2_fill_1 FILLER_71_747 ();
 sg13g2_decap_8 FILLER_71_764 ();
 sg13g2_fill_2 FILLER_71_771 ();
 sg13g2_decap_4 FILLER_71_792 ();
 sg13g2_fill_1 FILLER_71_796 ();
 sg13g2_fill_1 FILLER_71_802 ();
 sg13g2_decap_4 FILLER_71_813 ();
 sg13g2_fill_1 FILLER_71_817 ();
 sg13g2_decap_8 FILLER_71_827 ();
 sg13g2_fill_2 FILLER_71_834 ();
 sg13g2_fill_1 FILLER_71_836 ();
 sg13g2_decap_4 FILLER_71_845 ();
 sg13g2_fill_1 FILLER_71_849 ();
 sg13g2_decap_4 FILLER_71_858 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_19 ();
 sg13g2_fill_2 FILLER_72_38 ();
 sg13g2_fill_2 FILLER_72_96 ();
 sg13g2_fill_1 FILLER_72_98 ();
 sg13g2_fill_1 FILLER_72_127 ();
 sg13g2_fill_2 FILLER_72_163 ();
 sg13g2_decap_4 FILLER_72_183 ();
 sg13g2_fill_2 FILLER_72_187 ();
 sg13g2_decap_8 FILLER_72_211 ();
 sg13g2_fill_2 FILLER_72_218 ();
 sg13g2_fill_1 FILLER_72_220 ();
 sg13g2_decap_8 FILLER_72_257 ();
 sg13g2_decap_8 FILLER_72_272 ();
 sg13g2_decap_8 FILLER_72_279 ();
 sg13g2_fill_1 FILLER_72_286 ();
 sg13g2_fill_2 FILLER_72_291 ();
 sg13g2_fill_1 FILLER_72_301 ();
 sg13g2_fill_2 FILLER_72_316 ();
 sg13g2_fill_1 FILLER_72_318 ();
 sg13g2_decap_4 FILLER_72_349 ();
 sg13g2_fill_1 FILLER_72_353 ();
 sg13g2_fill_2 FILLER_72_364 ();
 sg13g2_fill_2 FILLER_72_371 ();
 sg13g2_fill_2 FILLER_72_395 ();
 sg13g2_fill_1 FILLER_72_397 ();
 sg13g2_fill_1 FILLER_72_403 ();
 sg13g2_decap_4 FILLER_72_409 ();
 sg13g2_decap_8 FILLER_72_426 ();
 sg13g2_decap_8 FILLER_72_433 ();
 sg13g2_decap_8 FILLER_72_440 ();
 sg13g2_fill_2 FILLER_72_447 ();
 sg13g2_fill_1 FILLER_72_449 ();
 sg13g2_decap_4 FILLER_72_462 ();
 sg13g2_fill_1 FILLER_72_466 ();
 sg13g2_fill_1 FILLER_72_487 ();
 sg13g2_fill_2 FILLER_72_496 ();
 sg13g2_fill_2 FILLER_72_504 ();
 sg13g2_fill_1 FILLER_72_506 ();
 sg13g2_decap_4 FILLER_72_531 ();
 sg13g2_fill_1 FILLER_72_535 ();
 sg13g2_fill_2 FILLER_72_553 ();
 sg13g2_decap_4 FILLER_72_572 ();
 sg13g2_fill_2 FILLER_72_576 ();
 sg13g2_decap_4 FILLER_72_583 ();
 sg13g2_fill_2 FILLER_72_596 ();
 sg13g2_decap_8 FILLER_72_613 ();
 sg13g2_decap_4 FILLER_72_620 ();
 sg13g2_fill_2 FILLER_72_624 ();
 sg13g2_fill_2 FILLER_72_635 ();
 sg13g2_fill_1 FILLER_72_637 ();
 sg13g2_decap_8 FILLER_72_655 ();
 sg13g2_decap_4 FILLER_72_662 ();
 sg13g2_fill_2 FILLER_72_682 ();
 sg13g2_fill_1 FILLER_72_700 ();
 sg13g2_fill_1 FILLER_72_716 ();
 sg13g2_decap_8 FILLER_72_738 ();
 sg13g2_decap_4 FILLER_72_750 ();
 sg13g2_fill_1 FILLER_72_754 ();
 sg13g2_fill_2 FILLER_72_761 ();
 sg13g2_fill_1 FILLER_72_763 ();
 sg13g2_fill_2 FILLER_72_770 ();
 sg13g2_fill_1 FILLER_72_772 ();
 sg13g2_decap_8 FILLER_72_783 ();
 sg13g2_fill_2 FILLER_72_808 ();
 sg13g2_fill_1 FILLER_72_810 ();
 sg13g2_fill_2 FILLER_72_817 ();
 sg13g2_decap_8 FILLER_72_825 ();
 sg13g2_fill_1 FILLER_72_832 ();
 sg13g2_decap_8 FILLER_72_838 ();
 sg13g2_decap_4 FILLER_72_845 ();
 sg13g2_fill_1 FILLER_72_849 ();
 sg13g2_decap_8 FILLER_72_855 ();
 sg13g2_fill_2 FILLER_73_26 ();
 sg13g2_decap_8 FILLER_73_85 ();
 sg13g2_fill_2 FILLER_73_131 ();
 sg13g2_fill_2 FILLER_73_138 ();
 sg13g2_fill_1 FILLER_73_140 ();
 sg13g2_fill_2 FILLER_73_149 ();
 sg13g2_decap_4 FILLER_73_165 ();
 sg13g2_fill_1 FILLER_73_169 ();
 sg13g2_fill_1 FILLER_73_209 ();
 sg13g2_decap_8 FILLER_73_216 ();
 sg13g2_decap_8 FILLER_73_223 ();
 sg13g2_fill_2 FILLER_73_230 ();
 sg13g2_fill_1 FILLER_73_236 ();
 sg13g2_decap_8 FILLER_73_240 ();
 sg13g2_fill_1 FILLER_73_256 ();
 sg13g2_fill_1 FILLER_73_293 ();
 sg13g2_fill_2 FILLER_73_311 ();
 sg13g2_fill_1 FILLER_73_313 ();
 sg13g2_decap_4 FILLER_73_322 ();
 sg13g2_fill_2 FILLER_73_342 ();
 sg13g2_decap_4 FILLER_73_362 ();
 sg13g2_fill_2 FILLER_73_366 ();
 sg13g2_fill_2 FILLER_73_382 ();
 sg13g2_fill_1 FILLER_73_384 ();
 sg13g2_fill_2 FILLER_73_389 ();
 sg13g2_fill_1 FILLER_73_391 ();
 sg13g2_fill_2 FILLER_73_398 ();
 sg13g2_fill_2 FILLER_73_426 ();
 sg13g2_fill_1 FILLER_73_428 ();
 sg13g2_decap_8 FILLER_73_437 ();
 sg13g2_fill_1 FILLER_73_460 ();
 sg13g2_decap_4 FILLER_73_467 ();
 sg13g2_fill_2 FILLER_73_471 ();
 sg13g2_decap_8 FILLER_73_478 ();
 sg13g2_fill_1 FILLER_73_485 ();
 sg13g2_decap_8 FILLER_73_496 ();
 sg13g2_decap_8 FILLER_73_511 ();
 sg13g2_fill_2 FILLER_73_518 ();
 sg13g2_fill_1 FILLER_73_520 ();
 sg13g2_decap_8 FILLER_73_526 ();
 sg13g2_decap_4 FILLER_73_533 ();
 sg13g2_fill_2 FILLER_73_537 ();
 sg13g2_decap_4 FILLER_73_552 ();
 sg13g2_fill_2 FILLER_73_556 ();
 sg13g2_fill_2 FILLER_73_563 ();
 sg13g2_fill_1 FILLER_73_565 ();
 sg13g2_fill_2 FILLER_73_580 ();
 sg13g2_decap_8 FILLER_73_606 ();
 sg13g2_decap_8 FILLER_73_613 ();
 sg13g2_fill_1 FILLER_73_625 ();
 sg13g2_decap_4 FILLER_73_637 ();
 sg13g2_fill_2 FILLER_73_641 ();
 sg13g2_decap_4 FILLER_73_648 ();
 sg13g2_decap_4 FILLER_73_657 ();
 sg13g2_fill_1 FILLER_73_667 ();
 sg13g2_decap_8 FILLER_73_691 ();
 sg13g2_decap_8 FILLER_73_698 ();
 sg13g2_fill_2 FILLER_73_705 ();
 sg13g2_fill_1 FILLER_73_707 ();
 sg13g2_decap_4 FILLER_73_711 ();
 sg13g2_decap_4 FILLER_73_728 ();
 sg13g2_fill_2 FILLER_73_738 ();
 sg13g2_fill_1 FILLER_73_740 ();
 sg13g2_fill_2 FILLER_73_750 ();
 sg13g2_fill_1 FILLER_73_752 ();
 sg13g2_fill_2 FILLER_73_759 ();
 sg13g2_fill_1 FILLER_73_767 ();
 sg13g2_decap_8 FILLER_73_790 ();
 sg13g2_fill_2 FILLER_73_797 ();
 sg13g2_decap_4 FILLER_73_810 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_91 ();
 sg13g2_fill_1 FILLER_74_93 ();
 sg13g2_fill_2 FILLER_74_99 ();
 sg13g2_fill_2 FILLER_74_119 ();
 sg13g2_fill_1 FILLER_74_138 ();
 sg13g2_fill_2 FILLER_74_143 ();
 sg13g2_fill_1 FILLER_74_183 ();
 sg13g2_decap_4 FILLER_74_192 ();
 sg13g2_decap_8 FILLER_74_223 ();
 sg13g2_decap_4 FILLER_74_230 ();
 sg13g2_fill_1 FILLER_74_234 ();
 sg13g2_fill_2 FILLER_74_243 ();
 sg13g2_decap_8 FILLER_74_258 ();
 sg13g2_decap_8 FILLER_74_265 ();
 sg13g2_fill_1 FILLER_74_272 ();
 sg13g2_decap_8 FILLER_74_277 ();
 sg13g2_decap_8 FILLER_74_284 ();
 sg13g2_decap_4 FILLER_74_291 ();
 sg13g2_fill_1 FILLER_74_295 ();
 sg13g2_decap_8 FILLER_74_308 ();
 sg13g2_decap_8 FILLER_74_315 ();
 sg13g2_fill_1 FILLER_74_322 ();
 sg13g2_fill_2 FILLER_74_342 ();
 sg13g2_fill_2 FILLER_74_388 ();
 sg13g2_decap_4 FILLER_74_395 ();
 sg13g2_fill_2 FILLER_74_399 ();
 sg13g2_fill_1 FILLER_74_410 ();
 sg13g2_decap_8 FILLER_74_415 ();
 sg13g2_decap_8 FILLER_74_422 ();
 sg13g2_decap_4 FILLER_74_429 ();
 sg13g2_fill_1 FILLER_74_433 ();
 sg13g2_fill_1 FILLER_74_446 ();
 sg13g2_fill_2 FILLER_74_452 ();
 sg13g2_fill_1 FILLER_74_454 ();
 sg13g2_decap_8 FILLER_74_463 ();
 sg13g2_decap_4 FILLER_74_470 ();
 sg13g2_fill_1 FILLER_74_474 ();
 sg13g2_decap_4 FILLER_74_492 ();
 sg13g2_fill_1 FILLER_74_496 ();
 sg13g2_fill_1 FILLER_74_513 ();
 sg13g2_decap_8 FILLER_74_534 ();
 sg13g2_fill_2 FILLER_74_541 ();
 sg13g2_decap_4 FILLER_74_564 ();
 sg13g2_fill_2 FILLER_74_568 ();
 sg13g2_decap_4 FILLER_74_582 ();
 sg13g2_fill_2 FILLER_74_590 ();
 sg13g2_decap_4 FILLER_74_600 ();
 sg13g2_fill_2 FILLER_74_622 ();
 sg13g2_fill_1 FILLER_74_624 ();
 sg13g2_decap_4 FILLER_74_646 ();
 sg13g2_decap_4 FILLER_74_671 ();
 sg13g2_fill_1 FILLER_74_684 ();
 sg13g2_decap_4 FILLER_74_690 ();
 sg13g2_fill_2 FILLER_74_694 ();
 sg13g2_fill_1 FILLER_74_723 ();
 sg13g2_fill_2 FILLER_74_734 ();
 sg13g2_decap_4 FILLER_74_748 ();
 sg13g2_fill_1 FILLER_74_752 ();
 sg13g2_decap_4 FILLER_74_767 ();
 sg13g2_fill_2 FILLER_74_771 ();
 sg13g2_fill_1 FILLER_74_778 ();
 sg13g2_fill_1 FILLER_74_785 ();
 sg13g2_decap_8 FILLER_74_792 ();
 sg13g2_decap_8 FILLER_74_799 ();
 sg13g2_fill_2 FILLER_74_806 ();
 sg13g2_decap_4 FILLER_74_812 ();
 sg13g2_fill_2 FILLER_74_816 ();
 sg13g2_fill_2 FILLER_74_831 ();
 sg13g2_decap_4 FILLER_74_837 ();
 sg13g2_fill_1 FILLER_74_841 ();
 sg13g2_decap_8 FILLER_74_850 ();
 sg13g2_decap_4 FILLER_74_857 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_30 ();
 sg13g2_fill_1 FILLER_75_40 ();
 sg13g2_fill_2 FILLER_75_52 ();
 sg13g2_fill_1 FILLER_75_54 ();
 sg13g2_fill_2 FILLER_75_102 ();
 sg13g2_fill_1 FILLER_75_104 ();
 sg13g2_decap_8 FILLER_75_114 ();
 sg13g2_fill_2 FILLER_75_173 ();
 sg13g2_fill_1 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_180 ();
 sg13g2_fill_1 FILLER_75_187 ();
 sg13g2_fill_2 FILLER_75_202 ();
 sg13g2_fill_1 FILLER_75_204 ();
 sg13g2_fill_1 FILLER_75_210 ();
 sg13g2_fill_2 FILLER_75_224 ();
 sg13g2_fill_1 FILLER_75_226 ();
 sg13g2_decap_4 FILLER_75_273 ();
 sg13g2_fill_1 FILLER_75_287 ();
 sg13g2_decap_4 FILLER_75_331 ();
 sg13g2_fill_2 FILLER_75_340 ();
 sg13g2_fill_1 FILLER_75_342 ();
 sg13g2_fill_1 FILLER_75_348 ();
 sg13g2_fill_2 FILLER_75_376 ();
 sg13g2_fill_1 FILLER_75_390 ();
 sg13g2_fill_2 FILLER_75_408 ();
 sg13g2_fill_2 FILLER_75_413 ();
 sg13g2_fill_2 FILLER_75_423 ();
 sg13g2_decap_8 FILLER_75_437 ();
 sg13g2_decap_4 FILLER_75_444 ();
 sg13g2_fill_1 FILLER_75_448 ();
 sg13g2_decap_4 FILLER_75_455 ();
 sg13g2_fill_1 FILLER_75_463 ();
 sg13g2_fill_2 FILLER_75_484 ();
 sg13g2_fill_1 FILLER_75_486 ();
 sg13g2_decap_8 FILLER_75_509 ();
 sg13g2_fill_1 FILLER_75_516 ();
 sg13g2_decap_8 FILLER_75_554 ();
 sg13g2_fill_1 FILLER_75_561 ();
 sg13g2_decap_8 FILLER_75_606 ();
 sg13g2_decap_8 FILLER_75_613 ();
 sg13g2_decap_4 FILLER_75_635 ();
 sg13g2_decap_8 FILLER_75_659 ();
 sg13g2_fill_1 FILLER_75_666 ();
 sg13g2_fill_1 FILLER_75_672 ();
 sg13g2_fill_2 FILLER_75_688 ();
 sg13g2_fill_1 FILLER_75_695 ();
 sg13g2_decap_4 FILLER_75_709 ();
 sg13g2_fill_2 FILLER_75_713 ();
 sg13g2_fill_2 FILLER_75_721 ();
 sg13g2_fill_1 FILLER_75_723 ();
 sg13g2_decap_8 FILLER_75_730 ();
 sg13g2_decap_4 FILLER_75_737 ();
 sg13g2_fill_2 FILLER_75_741 ();
 sg13g2_decap_8 FILLER_75_755 ();
 sg13g2_fill_1 FILLER_75_762 ();
 sg13g2_fill_2 FILLER_75_767 ();
 sg13g2_decap_4 FILLER_75_774 ();
 sg13g2_fill_2 FILLER_75_778 ();
 sg13g2_fill_2 FILLER_75_804 ();
 sg13g2_fill_1 FILLER_75_806 ();
 sg13g2_decap_8 FILLER_75_835 ();
 sg13g2_decap_8 FILLER_75_842 ();
 sg13g2_decap_8 FILLER_75_849 ();
 sg13g2_decap_4 FILLER_75_856 ();
 sg13g2_fill_2 FILLER_75_860 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_42 ();
 sg13g2_fill_2 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_131 ();
 sg13g2_decap_4 FILLER_76_138 ();
 sg13g2_fill_1 FILLER_76_151 ();
 sg13g2_decap_4 FILLER_76_200 ();
 sg13g2_fill_1 FILLER_76_268 ();
 sg13g2_decap_4 FILLER_76_297 ();
 sg13g2_decap_4 FILLER_76_306 ();
 sg13g2_fill_2 FILLER_76_310 ();
 sg13g2_fill_2 FILLER_76_321 ();
 sg13g2_decap_4 FILLER_76_328 ();
 sg13g2_fill_1 FILLER_76_332 ();
 sg13g2_decap_8 FILLER_76_380 ();
 sg13g2_fill_2 FILLER_76_387 ();
 sg13g2_fill_2 FILLER_76_432 ();
 sg13g2_fill_1 FILLER_76_434 ();
 sg13g2_fill_2 FILLER_76_447 ();
 sg13g2_fill_1 FILLER_76_449 ();
 sg13g2_fill_2 FILLER_76_458 ();
 sg13g2_fill_1 FILLER_76_460 ();
 sg13g2_decap_8 FILLER_76_469 ();
 sg13g2_fill_2 FILLER_76_476 ();
 sg13g2_fill_1 FILLER_76_478 ();
 sg13g2_decap_8 FILLER_76_484 ();
 sg13g2_fill_2 FILLER_76_491 ();
 sg13g2_fill_1 FILLER_76_493 ();
 sg13g2_decap_4 FILLER_76_504 ();
 sg13g2_fill_2 FILLER_76_508 ();
 sg13g2_decap_8 FILLER_76_526 ();
 sg13g2_decap_8 FILLER_76_533 ();
 sg13g2_decap_4 FILLER_76_560 ();
 sg13g2_fill_1 FILLER_76_564 ();
 sg13g2_decap_8 FILLER_76_570 ();
 sg13g2_fill_1 FILLER_76_577 ();
 sg13g2_decap_8 FILLER_76_583 ();
 sg13g2_fill_1 FILLER_76_590 ();
 sg13g2_decap_4 FILLER_76_595 ();
 sg13g2_fill_1 FILLER_76_599 ();
 sg13g2_decap_4 FILLER_76_608 ();
 sg13g2_fill_1 FILLER_76_612 ();
 sg13g2_decap_4 FILLER_76_619 ();
 sg13g2_fill_1 FILLER_76_623 ();
 sg13g2_fill_1 FILLER_76_634 ();
 sg13g2_decap_4 FILLER_76_640 ();
 sg13g2_fill_1 FILLER_76_644 ();
 sg13g2_decap_4 FILLER_76_653 ();
 sg13g2_decap_8 FILLER_76_663 ();
 sg13g2_fill_2 FILLER_76_670 ();
 sg13g2_fill_1 FILLER_76_682 ();
 sg13g2_decap_8 FILLER_76_694 ();
 sg13g2_fill_1 FILLER_76_701 ();
 sg13g2_decap_4 FILLER_76_712 ();
 sg13g2_fill_1 FILLER_76_716 ();
 sg13g2_fill_1 FILLER_76_723 ();
 sg13g2_decap_8 FILLER_76_729 ();
 sg13g2_fill_2 FILLER_76_736 ();
 sg13g2_fill_2 FILLER_76_744 ();
 sg13g2_fill_1 FILLER_76_766 ();
 sg13g2_fill_2 FILLER_76_779 ();
 sg13g2_decap_8 FILLER_76_793 ();
 sg13g2_fill_2 FILLER_76_800 ();
 sg13g2_fill_1 FILLER_76_802 ();
 sg13g2_decap_4 FILLER_76_807 ();
 sg13g2_decap_4 FILLER_76_824 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_8 FILLER_76_849 ();
 sg13g2_decap_4 FILLER_76_856 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_4 FILLER_77_7 ();
 sg13g2_fill_2 FILLER_77_11 ();
 sg13g2_fill_2 FILLER_77_17 ();
 sg13g2_fill_1 FILLER_77_19 ();
 sg13g2_fill_1 FILLER_77_33 ();
 sg13g2_fill_1 FILLER_77_52 ();
 sg13g2_fill_2 FILLER_77_58 ();
 sg13g2_fill_1 FILLER_77_60 ();
 sg13g2_fill_2 FILLER_77_74 ();
 sg13g2_fill_2 FILLER_77_107 ();
 sg13g2_fill_1 FILLER_77_109 ();
 sg13g2_fill_1 FILLER_77_123 ();
 sg13g2_decap_4 FILLER_77_188 ();
 sg13g2_decap_4 FILLER_77_221 ();
 sg13g2_fill_1 FILLER_77_230 ();
 sg13g2_fill_2 FILLER_77_261 ();
 sg13g2_fill_2 FILLER_77_277 ();
 sg13g2_fill_1 FILLER_77_296 ();
 sg13g2_fill_1 FILLER_77_307 ();
 sg13g2_fill_2 FILLER_77_357 ();
 sg13g2_fill_1 FILLER_77_364 ();
 sg13g2_fill_2 FILLER_77_373 ();
 sg13g2_fill_1 FILLER_77_375 ();
 sg13g2_fill_1 FILLER_77_380 ();
 sg13g2_fill_2 FILLER_77_392 ();
 sg13g2_fill_1 FILLER_77_394 ();
 sg13g2_fill_2 FILLER_77_405 ();
 sg13g2_decap_8 FILLER_77_411 ();
 sg13g2_decap_8 FILLER_77_418 ();
 sg13g2_fill_2 FILLER_77_425 ();
 sg13g2_fill_1 FILLER_77_427 ();
 sg13g2_fill_2 FILLER_77_433 ();
 sg13g2_fill_1 FILLER_77_435 ();
 sg13g2_decap_4 FILLER_77_445 ();
 sg13g2_fill_1 FILLER_77_449 ();
 sg13g2_fill_2 FILLER_77_478 ();
 sg13g2_fill_2 FILLER_77_494 ();
 sg13g2_decap_8 FILLER_77_510 ();
 sg13g2_decap_4 FILLER_77_517 ();
 sg13g2_fill_1 FILLER_77_527 ();
 sg13g2_fill_1 FILLER_77_541 ();
 sg13g2_fill_2 FILLER_77_550 ();
 sg13g2_fill_1 FILLER_77_552 ();
 sg13g2_fill_2 FILLER_77_561 ();
 sg13g2_fill_1 FILLER_77_563 ();
 sg13g2_fill_2 FILLER_77_580 ();
 sg13g2_fill_1 FILLER_77_582 ();
 sg13g2_decap_4 FILLER_77_612 ();
 sg13g2_decap_4 FILLER_77_634 ();
 sg13g2_decap_4 FILLER_77_656 ();
 sg13g2_fill_2 FILLER_77_660 ();
 sg13g2_fill_2 FILLER_77_676 ();
 sg13g2_fill_1 FILLER_77_678 ();
 sg13g2_decap_4 FILLER_77_682 ();
 sg13g2_fill_2 FILLER_77_690 ();
 sg13g2_fill_2 FILLER_77_697 ();
 sg13g2_fill_1 FILLER_77_699 ();
 sg13g2_fill_2 FILLER_77_715 ();
 sg13g2_fill_1 FILLER_77_717 ();
 sg13g2_decap_8 FILLER_77_732 ();
 sg13g2_decap_8 FILLER_77_739 ();
 sg13g2_fill_1 FILLER_77_746 ();
 sg13g2_decap_8 FILLER_77_755 ();
 sg13g2_decap_8 FILLER_77_762 ();
 sg13g2_fill_2 FILLER_77_769 ();
 sg13g2_fill_2 FILLER_77_790 ();
 sg13g2_fill_2 FILLER_77_816 ();
 sg13g2_fill_1 FILLER_77_818 ();
 sg13g2_decap_4 FILLER_77_824 ();
 sg13g2_decap_8 FILLER_77_831 ();
 sg13g2_decap_8 FILLER_77_838 ();
 sg13g2_fill_2 FILLER_77_845 ();
 sg13g2_decap_4 FILLER_77_858 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_48 ();
 sg13g2_fill_2 FILLER_78_99 ();
 sg13g2_fill_1 FILLER_78_101 ();
 sg13g2_decap_8 FILLER_78_138 ();
 sg13g2_decap_4 FILLER_78_145 ();
 sg13g2_fill_1 FILLER_78_158 ();
 sg13g2_fill_2 FILLER_78_185 ();
 sg13g2_decap_4 FILLER_78_222 ();
 sg13g2_fill_1 FILLER_78_235 ();
 sg13g2_fill_2 FILLER_78_253 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_fill_1 FILLER_78_335 ();
 sg13g2_fill_2 FILLER_78_349 ();
 sg13g2_fill_1 FILLER_78_355 ();
 sg13g2_fill_2 FILLER_78_391 ();
 sg13g2_fill_1 FILLER_78_401 ();
 sg13g2_fill_1 FILLER_78_436 ();
 sg13g2_fill_1 FILLER_78_453 ();
 sg13g2_decap_8 FILLER_78_462 ();
 sg13g2_fill_2 FILLER_78_469 ();
 sg13g2_fill_2 FILLER_78_477 ();
 sg13g2_decap_8 FILLER_78_484 ();
 sg13g2_decap_4 FILLER_78_491 ();
 sg13g2_fill_2 FILLER_78_495 ();
 sg13g2_fill_2 FILLER_78_502 ();
 sg13g2_fill_1 FILLER_78_504 ();
 sg13g2_fill_2 FILLER_78_513 ();
 sg13g2_fill_1 FILLER_78_515 ();
 sg13g2_decap_4 FILLER_78_530 ();
 sg13g2_fill_1 FILLER_78_534 ();
 sg13g2_fill_2 FILLER_78_544 ();
 sg13g2_fill_1 FILLER_78_546 ();
 sg13g2_decap_8 FILLER_78_555 ();
 sg13g2_decap_4 FILLER_78_562 ();
 sg13g2_fill_1 FILLER_78_566 ();
 sg13g2_fill_1 FILLER_78_571 ();
 sg13g2_decap_4 FILLER_78_577 ();
 sg13g2_fill_1 FILLER_78_581 ();
 sg13g2_decap_8 FILLER_78_587 ();
 sg13g2_decap_8 FILLER_78_598 ();
 sg13g2_fill_1 FILLER_78_605 ();
 sg13g2_decap_8 FILLER_78_612 ();
 sg13g2_fill_1 FILLER_78_619 ();
 sg13g2_fill_2 FILLER_78_632 ();
 sg13g2_decap_8 FILLER_78_651 ();
 sg13g2_fill_1 FILLER_78_658 ();
 sg13g2_decap_8 FILLER_78_675 ();
 sg13g2_fill_1 FILLER_78_682 ();
 sg13g2_decap_8 FILLER_78_699 ();
 sg13g2_decap_8 FILLER_78_706 ();
 sg13g2_fill_1 FILLER_78_744 ();
 sg13g2_fill_1 FILLER_78_771 ();
 sg13g2_decap_8 FILLER_78_780 ();
 sg13g2_decap_4 FILLER_78_787 ();
 sg13g2_fill_2 FILLER_78_791 ();
 sg13g2_fill_2 FILLER_78_799 ();
 sg13g2_fill_1 FILLER_78_801 ();
 sg13g2_fill_1 FILLER_78_822 ();
 sg13g2_decap_8 FILLER_78_839 ();
 sg13g2_decap_8 FILLER_78_846 ();
 sg13g2_decap_8 FILLER_78_853 ();
 sg13g2_fill_2 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_9 ();
 sg13g2_fill_2 FILLER_79_129 ();
 sg13g2_decap_8 FILLER_79_162 ();
 sg13g2_fill_1 FILLER_79_169 ();
 sg13g2_decap_8 FILLER_79_174 ();
 sg13g2_fill_2 FILLER_79_181 ();
 sg13g2_fill_1 FILLER_79_183 ();
 sg13g2_decap_8 FILLER_79_192 ();
 sg13g2_decap_4 FILLER_79_199 ();
 sg13g2_decap_4 FILLER_79_207 ();
 sg13g2_fill_2 FILLER_79_211 ();
 sg13g2_decap_4 FILLER_79_223 ();
 sg13g2_fill_1 FILLER_79_227 ();
 sg13g2_fill_1 FILLER_79_232 ();
 sg13g2_fill_2 FILLER_79_272 ();
 sg13g2_fill_1 FILLER_79_287 ();
 sg13g2_fill_1 FILLER_79_301 ();
 sg13g2_fill_1 FILLER_79_315 ();
 sg13g2_fill_2 FILLER_79_334 ();
 sg13g2_fill_1 FILLER_79_367 ();
 sg13g2_decap_8 FILLER_79_376 ();
 sg13g2_decap_4 FILLER_79_383 ();
 sg13g2_decap_8 FILLER_79_398 ();
 sg13g2_fill_2 FILLER_79_405 ();
 sg13g2_decap_8 FILLER_79_411 ();
 sg13g2_fill_2 FILLER_79_418 ();
 sg13g2_decap_8 FILLER_79_424 ();
 sg13g2_fill_1 FILLER_79_431 ();
 sg13g2_decap_8 FILLER_79_437 ();
 sg13g2_decap_4 FILLER_79_444 ();
 sg13g2_fill_2 FILLER_79_448 ();
 sg13g2_fill_1 FILLER_79_458 ();
 sg13g2_decap_8 FILLER_79_529 ();
 sg13g2_decap_4 FILLER_79_536 ();
 sg13g2_fill_1 FILLER_79_540 ();
 sg13g2_decap_8 FILLER_79_545 ();
 sg13g2_decap_4 FILLER_79_552 ();
 sg13g2_fill_2 FILLER_79_556 ();
 sg13g2_decap_4 FILLER_79_598 ();
 sg13g2_fill_2 FILLER_79_602 ();
 sg13g2_decap_8 FILLER_79_608 ();
 sg13g2_decap_4 FILLER_79_633 ();
 sg13g2_decap_8 FILLER_79_641 ();
 sg13g2_fill_1 FILLER_79_648 ();
 sg13g2_fill_2 FILLER_79_653 ();
 sg13g2_decap_4 FILLER_79_671 ();
 sg13g2_fill_1 FILLER_79_675 ();
 sg13g2_decap_8 FILLER_79_697 ();
 sg13g2_decap_8 FILLER_79_704 ();
 sg13g2_decap_8 FILLER_79_721 ();
 sg13g2_fill_2 FILLER_79_728 ();
 sg13g2_decap_8 FILLER_79_742 ();
 sg13g2_decap_4 FILLER_79_753 ();
 sg13g2_fill_2 FILLER_79_757 ();
 sg13g2_fill_2 FILLER_79_766 ();
 sg13g2_decap_8 FILLER_79_776 ();
 sg13g2_decap_8 FILLER_79_783 ();
 sg13g2_decap_8 FILLER_79_790 ();
 sg13g2_decap_8 FILLER_79_797 ();
 sg13g2_decap_8 FILLER_79_804 ();
 sg13g2_decap_8 FILLER_79_811 ();
 sg13g2_decap_8 FILLER_79_818 ();
 sg13g2_decap_8 FILLER_79_825 ();
 sg13g2_decap_8 FILLER_79_832 ();
 sg13g2_decap_8 FILLER_79_839 ();
 sg13g2_decap_8 FILLER_79_846 ();
 sg13g2_decap_8 FILLER_79_853 ();
 sg13g2_fill_2 FILLER_79_860 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_fill_2 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_16 ();
 sg13g2_fill_2 FILLER_80_34 ();
 sg13g2_fill_1 FILLER_80_87 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_4 FILLER_80_187 ();
 sg13g2_fill_1 FILLER_80_243 ();
 sg13g2_fill_2 FILLER_80_284 ();
 sg13g2_fill_2 FILLER_80_317 ();
 sg13g2_fill_2 FILLER_80_350 ();
 sg13g2_fill_1 FILLER_80_356 ();
 sg13g2_decap_4 FILLER_80_422 ();
 sg13g2_fill_1 FILLER_80_426 ();
 sg13g2_decap_4 FILLER_80_463 ();
 sg13g2_fill_2 FILLER_80_467 ();
 sg13g2_decap_8 FILLER_80_478 ();
 sg13g2_decap_8 FILLER_80_485 ();
 sg13g2_fill_2 FILLER_80_492 ();
 sg13g2_decap_8 FILLER_80_498 ();
 sg13g2_decap_4 FILLER_80_505 ();
 sg13g2_fill_2 FILLER_80_509 ();
 sg13g2_fill_2 FILLER_80_528 ();
 sg13g2_decap_8 FILLER_80_564 ();
 sg13g2_decap_8 FILLER_80_571 ();
 sg13g2_decap_8 FILLER_80_578 ();
 sg13g2_decap_8 FILLER_80_585 ();
 sg13g2_fill_1 FILLER_80_592 ();
 sg13g2_fill_1 FILLER_80_619 ();
 sg13g2_fill_2 FILLER_80_635 ();
 sg13g2_fill_1 FILLER_80_637 ();
 sg13g2_decap_8 FILLER_80_664 ();
 sg13g2_decap_8 FILLER_80_671 ();
 sg13g2_decap_8 FILLER_80_678 ();
 sg13g2_fill_1 FILLER_80_685 ();
 sg13g2_fill_1 FILLER_80_694 ();
 sg13g2_fill_1 FILLER_80_714 ();
 sg13g2_decap_8 FILLER_80_723 ();
 sg13g2_fill_2 FILLER_80_730 ();
 sg13g2_decap_8 FILLER_80_740 ();
 sg13g2_fill_2 FILLER_80_747 ();
 sg13g2_decap_8 FILLER_80_757 ();
 sg13g2_decap_8 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_776 ();
 sg13g2_decap_8 FILLER_80_783 ();
 sg13g2_decap_8 FILLER_80_790 ();
 sg13g2_decap_8 FILLER_80_797 ();
 sg13g2_decap_8 FILLER_80_804 ();
 sg13g2_decap_8 FILLER_80_811 ();
 sg13g2_decap_8 FILLER_80_818 ();
 sg13g2_decap_8 FILLER_80_825 ();
 sg13g2_decap_8 FILLER_80_832 ();
 sg13g2_decap_8 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_846 ();
 sg13g2_decap_8 FILLER_80_853 ();
 sg13g2_fill_2 FILLER_80_860 ();
 assign uio_oe[0] = net17;
 assign uio_oe[1] = net18;
 assign uio_oe[2] = net19;
 assign uio_oe[3] = net20;
 assign uio_out[0] = net21;
 assign uio_out[1] = net22;
 assign uio_out[2] = net23;
 assign uio_out[3] = net24;
endmodule
