module tt_um_iz_neuron (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire params_ready_internal;
 wire spike_out_internal;
 wire \system_inst.internal_param_a[0] ;
 wire \system_inst.internal_param_a[1] ;
 wire \system_inst.internal_param_a[2] ;
 wire \system_inst.internal_param_a[3] ;
 wire \system_inst.internal_param_a[4] ;
 wire \system_inst.internal_param_a[5] ;
 wire \system_inst.internal_param_a[6] ;
 wire \system_inst.internal_param_a[7] ;
 wire \system_inst.internal_param_b[0] ;
 wire \system_inst.internal_param_b[1] ;
 wire \system_inst.internal_param_b[2] ;
 wire \system_inst.internal_param_b[3] ;
 wire \system_inst.internal_param_b[4] ;
 wire \system_inst.internal_param_b[5] ;
 wire \system_inst.internal_param_b[6] ;
 wire \system_inst.internal_param_b[7] ;
 wire \system_inst.internal_param_c[0] ;
 wire \system_inst.internal_param_c[1] ;
 wire \system_inst.internal_param_c[2] ;
 wire \system_inst.internal_param_c[3] ;
 wire \system_inst.internal_param_c[4] ;
 wire \system_inst.internal_param_c[5] ;
 wire \system_inst.internal_param_c[6] ;
 wire \system_inst.internal_param_d[0] ;
 wire \system_inst.internal_param_d[1] ;
 wire \system_inst.internal_param_d[2] ;
 wire \system_inst.internal_param_d[3] ;
 wire \system_inst.internal_param_d[4] ;
 wire \system_inst.internal_param_d[5] ;
 wire \system_inst.internal_param_d[6] ;
 wire \system_inst.internal_param_d[7] ;
 wire \system_inst.loader.bit_count[0] ;
 wire \system_inst.loader.bit_count[1] ;
 wire \system_inst.loader.bit_count[2] ;
 wire \system_inst.loader.load_enable_prev ;
 wire \system_inst.loader.shift_reg[0] ;
 wire \system_inst.loader.shift_reg[1] ;
 wire \system_inst.loader.shift_reg[2] ;
 wire \system_inst.loader.shift_reg[3] ;
 wire \system_inst.loader.shift_reg[4] ;
 wire \system_inst.loader.shift_reg[5] ;
 wire \system_inst.loader.shift_reg[6] ;
 wire \system_inst.loader.state[0] ;
 wire \system_inst.loader.state[1] ;
 wire \system_inst.loader.state[2] ;
 wire \system_inst.loader.state[3] ;
 wire \system_inst.loader.state[4] ;
 wire \system_inst.loader.state[5] ;
 wire \system_inst.neuron.membrane_scaled[1] ;
 wire \system_inst.neuron.membrane_scaled[2] ;
 wire \system_inst.neuron.membrane_scaled[3] ;
 wire \system_inst.neuron.membrane_scaled[4] ;
 wire \system_inst.neuron.membrane_scaled[5] ;
 wire \system_inst.neuron.membrane_scaled[6] ;
 wire \system_inst.neuron.membrane_scaled[7] ;
 wire \system_inst.neuron.membrane_scaled[8] ;
 wire \system_inst.neuron.u[0] ;
 wire \system_inst.neuron.u[10] ;
 wire \system_inst.neuron.u[11] ;
 wire \system_inst.neuron.u[12] ;
 wire \system_inst.neuron.u[13] ;
 wire \system_inst.neuron.u[1] ;
 wire \system_inst.neuron.u[2] ;
 wire \system_inst.neuron.u[3] ;
 wire \system_inst.neuron.u[4] ;
 wire \system_inst.neuron.u[5] ;
 wire \system_inst.neuron.u[6] ;
 wire \system_inst.neuron.u[7] ;
 wire \system_inst.neuron.u[8] ;
 wire \system_inst.neuron.u[9] ;
 wire \system_inst.neuron.v[10] ;
 wire \system_inst.neuron.v[11] ;
 wire \system_inst.neuron.v[12] ;
 wire \system_inst.neuron.v[13] ;
 wire \system_inst.neuron.v[8] ;
 wire \system_inst.neuron.v[9] ;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire clknet_0_clk;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;

 sg13g2_inv_1 _3028_ (.Y(_1164_),
    .A(\system_inst.neuron.u[12] ));
 sg13g2_inv_1 _3029_ (.Y(_1175_),
    .A(net181));
 sg13g2_inv_1 _3030_ (.Y(_1186_),
    .A(\system_inst.neuron.u[5] ));
 sg13g2_inv_2 _3031_ (.Y(_1197_),
    .A(net142));
 sg13g2_inv_2 _3032_ (.Y(_1208_),
    .A(net119));
 sg13g2_inv_2 _3033_ (.Y(_1219_),
    .A(net121));
 sg13g2_inv_2 _3034_ (.Y(_1230_),
    .A(net137));
 sg13g2_inv_2 _3035_ (.Y(_1241_),
    .A(net139));
 sg13g2_inv_2 _3036_ (.Y(_1252_),
    .A(net128));
 sg13g2_inv_1 _3037_ (.Y(_1263_),
    .A(net122));
 sg13g2_inv_1 _3038_ (.Y(_1274_),
    .A(net124));
 sg13g2_inv_1 _3039_ (.Y(_1285_),
    .A(net112));
 sg13g2_inv_1 _3040_ (.Y(_1296_),
    .A(net160));
 sg13g2_inv_1 _3041_ (.Y(_1307_),
    .A(net768));
 sg13g2_inv_1 _3042_ (.Y(_1318_),
    .A(net775));
 sg13g2_inv_1 _3043_ (.Y(_1329_),
    .A(net778));
 sg13g2_inv_1 _3044_ (.Y(_1340_),
    .A(net786));
 sg13g2_inv_2 _3045_ (.Y(_1351_),
    .A(\system_inst.neuron.u[1] ));
 sg13g2_inv_2 _3046_ (.Y(_1362_),
    .A(\system_inst.neuron.u[0] ));
 sg13g2_inv_4 _3047_ (.A(net798),
    .Y(_1373_));
 sg13g2_inv_2 _3048_ (.Y(_1384_),
    .A(net803));
 sg13g2_inv_2 _3049_ (.Y(_1395_),
    .A(net848));
 sg13g2_inv_4 _3050_ (.A(net856),
    .Y(_1406_));
 sg13g2_inv_4 _3051_ (.A(net870),
    .Y(_1417_));
 sg13g2_inv_1 _3052_ (.Y(_1428_),
    .A(_0033_));
 sg13g2_inv_1 _3053_ (.Y(_1439_),
    .A(net4));
 sg13g2_inv_1 _3054_ (.Y(_1450_),
    .A(_0026_));
 sg13g2_inv_1 _3055_ (.Y(_1461_),
    .A(_0015_));
 sg13g2_inv_4 _3056_ (.A(_0019_),
    .Y(_1472_));
 sg13g2_inv_1 _3057_ (.Y(_1483_),
    .A(net157));
 sg13g2_inv_1 _3058_ (.Y(_1494_),
    .A(_0034_));
 sg13g2_inv_1 _3059_ (.Y(_1505_),
    .A(\system_inst.loader.state[1] ));
 sg13g2_inv_1 _3060_ (.Y(_1516_),
    .A(net882));
 sg13g2_inv_1 _3061_ (.Y(_1527_),
    .A(_0006_));
 sg13g2_nand2_2 _3062_ (.Y(_1538_),
    .A(net805),
    .B(net810));
 sg13g2_and2_2 _3063_ (.A(net816),
    .B(net820),
    .X(_1549_));
 sg13g2_nand2_2 _3064_ (.Y(_1560_),
    .A(net816),
    .B(net820));
 sg13g2_o21ai_1 _3065_ (.B1(_1384_),
    .Y(_1571_),
    .A1(_1538_),
    .A2(_1560_));
 sg13g2_nand2_1 _3066_ (.Y(_1582_),
    .A(_1373_),
    .B(_1571_));
 sg13g2_nor2_1 _3067_ (.A(net814),
    .B(net819),
    .Y(_1593_));
 sg13g2_nor3_1 _3068_ (.A(_0024_),
    .B(_1538_),
    .C(_1593_),
    .Y(_1604_));
 sg13g2_xnor2_1 _3069_ (.Y(_1615_),
    .A(net801),
    .B(_1604_));
 sg13g2_nor2_2 _3070_ (.A(net815),
    .B(net826),
    .Y(_1626_));
 sg13g2_nand3b_1 _3071_ (.B(_1626_),
    .C(net819),
    .Y(_1637_),
    .A_N(_0025_));
 sg13g2_nor2_1 _3072_ (.A(net808),
    .B(net811),
    .Y(_1648_));
 sg13g2_nor2b_1 _3073_ (.A(_1538_),
    .B_N(_1593_),
    .Y(_1659_));
 sg13g2_o21ai_1 _3074_ (.B1(_0024_),
    .Y(_1670_),
    .A1(_1648_),
    .A2(_1659_));
 sg13g2_a21oi_1 _3075_ (.A1(net801),
    .A2(_1670_),
    .Y(_1681_),
    .B1(_1637_));
 sg13g2_or2_1 _3076_ (.X(_1692_),
    .B(_1681_),
    .A(_1615_));
 sg13g2_and2_2 _3077_ (.A(net722),
    .B(_1692_),
    .X(_1703_));
 sg13g2_inv_1 _3078_ (.Y(uo_out[0]),
    .A(_1703_));
 sg13g2_o21ai_1 _3079_ (.B1(_1703_),
    .Y(uo_out[1]),
    .A1(_0033_),
    .A2(_1615_));
 sg13g2_o21ai_1 _3080_ (.B1(_1703_),
    .Y(uo_out[2]),
    .A1(_0032_),
    .A2(_1615_));
 sg13g2_o21ai_1 _3081_ (.B1(_1703_),
    .Y(uo_out[3]),
    .A1(_0031_),
    .A2(_1615_));
 sg13g2_o21ai_1 _3082_ (.B1(_1703_),
    .Y(uo_out[4]),
    .A1(_0030_),
    .A2(_1615_));
 sg13g2_o21ai_1 _3083_ (.B1(_1703_),
    .Y(uo_out[5]),
    .A1(_0029_),
    .A2(_1615_));
 sg13g2_o21ai_1 _3084_ (.B1(_1703_),
    .Y(uo_out[6]),
    .A1(_0028_),
    .A2(_1615_));
 sg13g2_o21ai_1 _3085_ (.B1(_1703_),
    .Y(uo_out[7]),
    .A1(_0027_),
    .A2(_1615_));
 sg13g2_nand2b_1 _3086_ (.Y(_1794_),
    .B(net11),
    .A_N(\system_inst.loader.load_enable_prev ));
 sg13g2_nor2_1 _3087_ (.A(net1),
    .B(net871),
    .Y(_1805_));
 sg13g2_o21ai_1 _3088_ (.B1(net166),
    .Y(_1816_),
    .A1(_1794_),
    .A2(_1805_));
 sg13g2_nand3b_1 _3089_ (.B(net1),
    .C(net133),
    .Y(_1827_),
    .A_N(net11));
 sg13g2_nand3_1 _3090_ (.B(_1816_),
    .C(_1827_),
    .A(net884),
    .Y(_0000_));
 sg13g2_nand2_2 _3091_ (.Y(_1848_),
    .A(net105),
    .B(net111));
 sg13g2_nand2_2 _3092_ (.Y(_1859_),
    .A(net11),
    .B(net1));
 sg13g2_nor3_2 _3093_ (.A(net159),
    .B(_1848_),
    .C(_1859_),
    .Y(_1870_));
 sg13g2_or3_2 _3094_ (.A(_0016_),
    .B(_1848_),
    .C(_1859_),
    .X(_1881_));
 sg13g2_nor2_2 _3095_ (.A(net133),
    .B(\system_inst.loader.state[0] ),
    .Y(_1892_));
 sg13g2_nor3_1 _3096_ (.A(\system_inst.loader.load_enable_prev ),
    .B(_1859_),
    .C(_1892_),
    .Y(_1903_));
 sg13g2_a21oi_1 _3097_ (.A1(net115),
    .A2(_1881_),
    .Y(_1914_),
    .B1(_1903_));
 sg13g2_nor2_1 _3098_ (.A(net872),
    .B(net116),
    .Y(_0003_));
 sg13g2_and2_1 _3099_ (.A(net11),
    .B(net882),
    .X(_0050_));
 sg13g2_a21o_1 _3100_ (.A2(_0050_),
    .A1(\system_inst.loader.load_enable_prev ),
    .B1(_1805_),
    .X(_1945_));
 sg13g2_nor2_1 _3101_ (.A(_1505_),
    .B(_1881_),
    .Y(_1956_));
 sg13g2_a22oi_1 _3102_ (.Y(_1967_),
    .B1(net719),
    .B2(net882),
    .A2(_1945_),
    .A1(net133));
 sg13g2_inv_1 _3103_ (.Y(_0004_),
    .A(net134));
 sg13g2_and2_2 _3104_ (.A(net108),
    .B(_1870_),
    .X(_1988_));
 sg13g2_nand2_1 _3105_ (.Y(_1999_),
    .A(net108),
    .B(_1870_));
 sg13g2_nand2_1 _3106_ (.Y(_2008_),
    .A(net127),
    .B(_1881_));
 sg13g2_a21oi_1 _3107_ (.A1(net716),
    .A2(_2008_),
    .Y(_0001_),
    .B1(net871));
 sg13g2_and2_2 _3108_ (.A(\system_inst.loader.state[2] ),
    .B(_1870_),
    .X(_2027_));
 sg13g2_nand2_2 _3109_ (.Y(_2034_),
    .A(net135),
    .B(_1870_));
 sg13g2_nand2_1 _3110_ (.Y(_2040_),
    .A(net108),
    .B(_1881_));
 sg13g2_a21oi_1 _3111_ (.A1(_2034_),
    .A2(_2040_),
    .Y(_0005_),
    .B1(net871));
 sg13g2_and2_1 _3112_ (.A(net115),
    .B(_1870_),
    .X(_2051_));
 sg13g2_a21oi_1 _3113_ (.A1(net135),
    .A2(_1881_),
    .Y(_2057_),
    .B1(net713));
 sg13g2_nor2_1 _3114_ (.A(net871),
    .B(_2057_),
    .Y(_0002_));
 sg13g2_and3_1 _3115_ (.X(_2070_),
    .A(net146),
    .B(net1),
    .C(net10));
 sg13g2_nand3_1 _3116_ (.B(net1),
    .C(net10),
    .A(net146),
    .Y(_2079_));
 sg13g2_nor2_2 _3117_ (.A(net720),
    .B(net725),
    .Y(_2087_));
 sg13g2_o21ai_1 _3118_ (.B1(net883),
    .Y(_2095_),
    .A1(net722),
    .A2(_2079_));
 sg13g2_inv_1 _3119_ (.Y(_2104_),
    .A(_2095_));
 sg13g2_and2_1 _3120_ (.A(net811),
    .B(net7),
    .X(_2114_));
 sg13g2_nand2_1 _3121_ (.Y(_2124_),
    .A(net806),
    .B(net8));
 sg13g2_xor2_1 _3122_ (.B(net8),
    .A(net806),
    .X(_2135_));
 sg13g2_xnor2_1 _3123_ (.Y(_2145_),
    .A(\system_inst.neuron.u[13] ),
    .B(net801));
 sg13g2_xor2_1 _3124_ (.B(_2135_),
    .A(_2114_),
    .X(_2155_));
 sg13g2_and2_1 _3125_ (.A(_2145_),
    .B(_2155_),
    .X(_2165_));
 sg13g2_a21oi_1 _3126_ (.A1(_2114_),
    .A2(_2135_),
    .Y(_2175_),
    .B1(_2165_));
 sg13g2_nand2_2 _3127_ (.Y(_2186_),
    .A(net798),
    .B(net802));
 sg13g2_xor2_1 _3128_ (.B(net803),
    .A(net799),
    .X(_2196_));
 sg13g2_nor2_1 _3129_ (.A(net9),
    .B(_2124_),
    .Y(_2205_));
 sg13g2_xor2_1 _3130_ (.B(_2124_),
    .A(net9),
    .X(_2211_));
 sg13g2_xor2_1 _3131_ (.B(_2211_),
    .A(_2196_),
    .X(_2212_));
 sg13g2_nand2b_1 _3132_ (.Y(_2213_),
    .B(_2212_),
    .A_N(_2175_));
 sg13g2_and2_1 _3133_ (.A(net802),
    .B(net864),
    .X(_2214_));
 sg13g2_nand2_2 _3134_ (.Y(_2215_),
    .A(net805),
    .B(net869));
 sg13g2_and3_2 _3135_ (.X(_2216_),
    .A(net805),
    .B(net869),
    .C(_2214_));
 sg13g2_nand2_2 _3136_ (.Y(_2217_),
    .A(net806),
    .B(net857));
 sg13g2_nor2b_1 _3137_ (.A(net869),
    .B_N(net798),
    .Y(_2218_));
 sg13g2_nand2_1 _3138_ (.Y(_2219_),
    .A(_2214_),
    .B(_2218_));
 sg13g2_xnor2_1 _3139_ (.Y(_2220_),
    .A(_2214_),
    .B(_2218_));
 sg13g2_xor2_1 _3140_ (.B(_2220_),
    .A(_2217_),
    .X(_2221_));
 sg13g2_nand2_1 _3141_ (.Y(_2222_),
    .A(_2216_),
    .B(_2221_));
 sg13g2_xnor2_1 _3142_ (.Y(_2223_),
    .A(_2216_),
    .B(_2221_));
 sg13g2_a22oi_1 _3143_ (.Y(_2224_),
    .B1(net849),
    .B2(net810),
    .A2(net844),
    .A1(net814));
 sg13g2_nand2_2 _3144_ (.Y(_2225_),
    .A(net811),
    .B(net843));
 sg13g2_nand4_1 _3145_ (.B(net814),
    .C(net843),
    .A(net810),
    .Y(_2226_),
    .D(net849));
 sg13g2_nor2b_2 _3146_ (.A(_2224_),
    .B_N(_2226_),
    .Y(_2227_));
 sg13g2_nand2_2 _3147_ (.Y(_2228_),
    .A(net818),
    .B(net837));
 sg13g2_nand3_1 _3148_ (.B(net838),
    .C(_2227_),
    .A(net818),
    .Y(_2229_));
 sg13g2_xor2_1 _3149_ (.B(_2228_),
    .A(_2227_),
    .X(_2230_));
 sg13g2_o21ai_1 _3150_ (.B1(_2222_),
    .Y(_2231_),
    .A1(_2223_),
    .A2(_2230_));
 sg13g2_nand2_2 _3151_ (.Y(_2232_),
    .A(net818),
    .B(net830));
 sg13g2_nand2_1 _3152_ (.Y(_2233_),
    .A(net810),
    .B(net837));
 sg13g2_nand2_2 _3153_ (.Y(_2234_),
    .A(net814),
    .B(net837));
 sg13g2_xor2_1 _3154_ (.B(_2234_),
    .A(_2225_),
    .X(_2235_));
 sg13g2_nand2b_1 _3155_ (.Y(_2236_),
    .B(_2235_),
    .A_N(_2232_));
 sg13g2_xnor2_1 _3156_ (.Y(_2237_),
    .A(_2232_),
    .B(_2235_));
 sg13g2_o21ai_1 _3157_ (.B1(_2219_),
    .Y(_2238_),
    .A1(_2217_),
    .A2(_2220_));
 sg13g2_and2_1 _3158_ (.A(net805),
    .B(net849),
    .X(_2239_));
 sg13g2_nand2_1 _3159_ (.Y(_2240_),
    .A(net806),
    .B(net850));
 sg13g2_nand2_2 _3160_ (.Y(_2241_),
    .A(net803),
    .B(net857));
 sg13g2_nor2b_1 _3161_ (.A(net864),
    .B_N(net799),
    .Y(_2242_));
 sg13g2_nor2b_1 _3162_ (.A(_2241_),
    .B_N(_2242_),
    .Y(_2243_));
 sg13g2_xnor2_1 _3163_ (.Y(_2244_),
    .A(_2241_),
    .B(_2242_));
 sg13g2_xnor2_1 _3164_ (.Y(_2245_),
    .A(_2240_),
    .B(_2244_));
 sg13g2_and2_1 _3165_ (.A(_2238_),
    .B(_2245_),
    .X(_2246_));
 sg13g2_or2_1 _3166_ (.X(_2247_),
    .B(_2245_),
    .A(_2238_));
 sg13g2_xnor2_1 _3167_ (.Y(_2248_),
    .A(_2238_),
    .B(_2245_));
 sg13g2_xnor2_1 _3168_ (.Y(_2249_),
    .A(_2237_),
    .B(_2248_));
 sg13g2_nand2_1 _3169_ (.Y(_2250_),
    .A(_2231_),
    .B(_2249_));
 sg13g2_and2_2 _3170_ (.A(net824),
    .B(net829),
    .X(_2251_));
 sg13g2_nand2_2 _3171_ (.Y(_2252_),
    .A(net824),
    .B(net829));
 sg13g2_and2_1 _3172_ (.A(_2226_),
    .B(_2229_),
    .X(_2253_));
 sg13g2_and2_2 _3173_ (.A(net820),
    .B(net824),
    .X(_2254_));
 sg13g2_xor2_1 _3174_ (.B(_2232_),
    .A(net825),
    .X(_2255_));
 sg13g2_nor2_1 _3175_ (.A(_2234_),
    .B(_2255_),
    .Y(_2256_));
 sg13g2_xor2_1 _3176_ (.B(_2255_),
    .A(_2234_),
    .X(_2257_));
 sg13g2_nor2b_1 _3177_ (.A(_2253_),
    .B_N(_2257_),
    .Y(_2258_));
 sg13g2_xnor2_1 _3178_ (.Y(_2259_),
    .A(_2253_),
    .B(_2257_));
 sg13g2_xnor2_1 _3179_ (.Y(_2260_),
    .A(_2251_),
    .B(_2259_));
 sg13g2_xnor2_1 _3180_ (.Y(_2261_),
    .A(_2231_),
    .B(_2249_));
 sg13g2_o21ai_1 _3181_ (.B1(_2250_),
    .Y(_2262_),
    .A1(_2260_),
    .A2(_2261_));
 sg13g2_a21oi_1 _3182_ (.A1(net830),
    .A2(_2254_),
    .Y(_2263_),
    .B1(_2256_));
 sg13g2_o21ai_1 _3183_ (.B1(_2236_),
    .Y(_2264_),
    .A1(_2225_),
    .A2(_2234_));
 sg13g2_nand2_1 _3184_ (.Y(_2265_),
    .A(net814),
    .B(net830));
 sg13g2_xnor2_1 _3185_ (.Y(_2266_),
    .A(_2254_),
    .B(_2265_));
 sg13g2_nand2b_1 _3186_ (.Y(_2267_),
    .B(_2266_),
    .A_N(_2233_));
 sg13g2_xnor2_1 _3187_ (.Y(_2268_),
    .A(_2233_),
    .B(_2266_));
 sg13g2_nand2_1 _3188_ (.Y(_2269_),
    .A(_2264_),
    .B(_2268_));
 sg13g2_xnor2_1 _3189_ (.Y(_2270_),
    .A(_2264_),
    .B(_2268_));
 sg13g2_xnor2_1 _3190_ (.Y(_2271_),
    .A(_2263_),
    .B(_2270_));
 sg13g2_a21oi_2 _3191_ (.B1(_2246_),
    .Y(_2272_),
    .A2(_2247_),
    .A1(_2237_));
 sg13g2_a21oi_2 _3192_ (.B1(_2243_),
    .Y(_2273_),
    .A2(_2244_),
    .A1(_2239_));
 sg13g2_nand2_2 _3193_ (.Y(_2274_),
    .A(net806),
    .B(net843));
 sg13g2_nor2_1 _3194_ (.A(_1395_),
    .B(net855),
    .Y(_2275_));
 sg13g2_nand2_2 _3195_ (.Y(_2276_),
    .A(net802),
    .B(net850));
 sg13g2_nor2b_2 _3196_ (.A(net856),
    .B_N(net799),
    .Y(_2277_));
 sg13g2_nand2b_1 _3197_ (.Y(_2278_),
    .B(_2277_),
    .A_N(_2276_));
 sg13g2_xnor2_1 _3198_ (.Y(_2279_),
    .A(_2276_),
    .B(_2277_));
 sg13g2_nand2b_1 _3199_ (.Y(_2280_),
    .B(_2279_),
    .A_N(_2274_));
 sg13g2_xnor2_1 _3200_ (.Y(_2281_),
    .A(_2274_),
    .B(_2279_));
 sg13g2_nor2b_1 _3201_ (.A(_2273_),
    .B_N(_2281_),
    .Y(_2282_));
 sg13g2_xnor2_1 _3202_ (.Y(_2283_),
    .A(_2273_),
    .B(_2281_));
 sg13g2_xnor2_1 _3203_ (.Y(_2284_),
    .A(_2268_),
    .B(_2283_));
 sg13g2_xor2_1 _3204_ (.B(_2284_),
    .A(_2272_),
    .X(_2285_));
 sg13g2_nand2b_1 _3205_ (.Y(_2286_),
    .B(_2285_),
    .A_N(_2271_));
 sg13g2_xnor2_1 _3206_ (.Y(_2287_),
    .A(_2271_),
    .B(_2285_));
 sg13g2_nand2_1 _3207_ (.Y(_2288_),
    .A(_2262_),
    .B(_2287_));
 sg13g2_o21ai_1 _3208_ (.B1(_2226_),
    .Y(_2289_),
    .A1(_2217_),
    .A2(_2224_));
 sg13g2_and2_2 _3209_ (.A(net842),
    .B(net848),
    .X(_2290_));
 sg13g2_nand2_2 _3210_ (.Y(_2291_),
    .A(net843),
    .B(net849));
 sg13g2_xnor2_1 _3211_ (.Y(_2292_),
    .A(_2225_),
    .B(_2239_));
 sg13g2_nand2b_1 _3212_ (.Y(_2293_),
    .B(_2292_),
    .A_N(_2241_));
 sg13g2_xnor2_1 _3213_ (.Y(_2294_),
    .A(_2241_),
    .B(_2292_));
 sg13g2_nand2_1 _3214_ (.Y(_2295_),
    .A(_2289_),
    .B(_2294_));
 sg13g2_and2_2 _3215_ (.A(net863),
    .B(net869),
    .X(_2296_));
 sg13g2_nand2_2 _3216_ (.Y(_2297_),
    .A(net863),
    .B(net869));
 sg13g2_o21ai_1 _3217_ (.B1(net798),
    .Y(_2298_),
    .A1(net864),
    .A2(net869));
 sg13g2_nand2b_2 _3218_ (.Y(_2299_),
    .B(_2297_),
    .A_N(_2298_));
 sg13g2_xnor2_1 _3219_ (.Y(_2300_),
    .A(_2289_),
    .B(_2294_));
 sg13g2_o21ai_1 _3220_ (.B1(_2295_),
    .Y(_2301_),
    .A1(net723),
    .A2(_2300_));
 sg13g2_a21o_1 _3221_ (.A2(_2259_),
    .A1(_2251_),
    .B1(_2258_),
    .X(_2302_));
 sg13g2_o21ai_1 _3222_ (.B1(_2293_),
    .Y(_2303_),
    .A1(_1538_),
    .A2(_2291_));
 sg13g2_nor2_2 _3223_ (.A(_1373_),
    .B(_1406_),
    .Y(_2304_));
 sg13g2_nand2_2 _3224_ (.Y(_2305_),
    .A(net802),
    .B(net843));
 sg13g2_xor2_1 _3225_ (.B(_2276_),
    .A(_2274_),
    .X(_2306_));
 sg13g2_nand2_1 _3226_ (.Y(_2307_),
    .A(_2304_),
    .B(_2306_));
 sg13g2_xor2_1 _3227_ (.B(_2306_),
    .A(_2304_),
    .X(_2308_));
 sg13g2_nand2_1 _3228_ (.Y(_2309_),
    .A(_2303_),
    .B(_2308_));
 sg13g2_xnor2_1 _3229_ (.Y(_2310_),
    .A(_2303_),
    .B(_2308_));
 sg13g2_xor2_1 _3230_ (.B(_2310_),
    .A(net723),
    .X(_2311_));
 sg13g2_xnor2_1 _3231_ (.Y(_2312_),
    .A(_2302_),
    .B(_2311_));
 sg13g2_nor2b_1 _3232_ (.A(_2312_),
    .B_N(_2301_),
    .Y(_2313_));
 sg13g2_xor2_1 _3233_ (.B(_2312_),
    .A(_2301_),
    .X(_2314_));
 sg13g2_xnor2_1 _3234_ (.Y(_2315_),
    .A(_2262_),
    .B(_2287_));
 sg13g2_o21ai_1 _3235_ (.B1(_2288_),
    .Y(_2316_),
    .A1(_2314_),
    .A2(_2315_));
 sg13g2_o21ai_1 _3236_ (.B1(_2309_),
    .Y(_2317_),
    .A1(_2299_),
    .A2(_2310_));
 sg13g2_o21ai_1 _3237_ (.B1(_2269_),
    .Y(_2318_),
    .A1(_2263_),
    .A2(_2270_));
 sg13g2_o21ai_1 _3238_ (.B1(_2307_),
    .Y(_2319_),
    .A1(_2240_),
    .A2(_2305_));
 sg13g2_nand2_1 _3239_ (.Y(_2320_),
    .A(net799),
    .B(net849));
 sg13g2_xor2_1 _3240_ (.B(_2320_),
    .A(_2305_),
    .X(_2321_));
 sg13g2_nand2_1 _3241_ (.Y(_2322_),
    .A(_2304_),
    .B(_2321_));
 sg13g2_xor2_1 _3242_ (.B(_2321_),
    .A(_2304_),
    .X(_2323_));
 sg13g2_nand2_1 _3243_ (.Y(_2324_),
    .A(_2319_),
    .B(_2323_));
 sg13g2_xnor2_1 _3244_ (.Y(_2325_),
    .A(_2319_),
    .B(_2323_));
 sg13g2_xor2_1 _3245_ (.B(_2325_),
    .A(_2299_),
    .X(_2326_));
 sg13g2_xnor2_1 _3246_ (.Y(_2327_),
    .A(_2318_),
    .B(_2326_));
 sg13g2_nor2b_1 _3247_ (.A(_2327_),
    .B_N(_2317_),
    .Y(_2328_));
 sg13g2_xor2_1 _3248_ (.B(_2327_),
    .A(_2317_),
    .X(_2329_));
 sg13g2_o21ai_1 _3249_ (.B1(_2286_),
    .Y(_2330_),
    .A1(_2272_),
    .A2(_2284_));
 sg13g2_nand2_2 _3250_ (.Y(_2331_),
    .A(net810),
    .B(net825));
 sg13g2_nand2_1 _3251_ (.Y(_2332_),
    .A(net815),
    .B(net824));
 sg13g2_nor2_1 _3252_ (.A(_2265_),
    .B(_2331_),
    .Y(_2333_));
 sg13g2_a22oi_1 _3253_ (.Y(_2334_),
    .B1(net830),
    .B2(net810),
    .A2(net825),
    .A1(net814));
 sg13g2_nor2_2 _3254_ (.A(_2333_),
    .B(_2334_),
    .Y(_2335_));
 sg13g2_nand2_2 _3255_ (.Y(_2336_),
    .A(net805),
    .B(net837));
 sg13g2_inv_1 _3256_ (.Y(_2337_),
    .A(_2336_));
 sg13g2_xnor2_1 _3257_ (.Y(_2338_),
    .A(_2335_),
    .B(_2336_));
 sg13g2_a21oi_2 _3258_ (.B1(_2282_),
    .Y(_2339_),
    .A2(_2283_),
    .A1(_2268_));
 sg13g2_nand2_1 _3259_ (.Y(_2340_),
    .A(_2278_),
    .B(_2280_));
 sg13g2_nor2_1 _3260_ (.A(_1373_),
    .B(net849),
    .Y(_2341_));
 sg13g2_nor2b_1 _3261_ (.A(_2305_),
    .B_N(_2341_),
    .Y(_2342_));
 sg13g2_xnor2_1 _3262_ (.Y(_2343_),
    .A(_2305_),
    .B(_2341_));
 sg13g2_xnor2_1 _3263_ (.Y(_2344_),
    .A(_2336_),
    .B(_2343_));
 sg13g2_nand2_1 _3264_ (.Y(_2345_),
    .A(_2340_),
    .B(_2344_));
 sg13g2_xnor2_1 _3265_ (.Y(_2346_),
    .A(_2340_),
    .B(_2344_));
 sg13g2_xnor2_1 _3266_ (.Y(_2347_),
    .A(net818),
    .B(_2335_));
 sg13g2_xor2_1 _3267_ (.B(_2347_),
    .A(_2346_),
    .X(_2348_));
 sg13g2_nor2b_1 _3268_ (.A(_2339_),
    .B_N(_2348_),
    .Y(_2349_));
 sg13g2_xnor2_1 _3269_ (.Y(_2350_),
    .A(_2339_),
    .B(_2348_));
 sg13g2_xor2_1 _3270_ (.B(_2350_),
    .A(_2338_),
    .X(_2351_));
 sg13g2_nand2_1 _3271_ (.Y(_2352_),
    .A(_2330_),
    .B(_2351_));
 sg13g2_xnor2_1 _3272_ (.Y(_2353_),
    .A(_2330_),
    .B(_2351_));
 sg13g2_xor2_1 _3273_ (.B(_2353_),
    .A(_2329_),
    .X(_2354_));
 sg13g2_and2_1 _3274_ (.A(_2316_),
    .B(_2354_),
    .X(_2355_));
 sg13g2_a21o_1 _3275_ (.A2(_2311_),
    .A1(_2302_),
    .B1(_2313_),
    .X(_2356_));
 sg13g2_xor2_1 _3276_ (.B(_2354_),
    .A(_2316_),
    .X(_2357_));
 sg13g2_a21oi_1 _3277_ (.A1(_2356_),
    .A2(_2357_),
    .Y(_2358_),
    .B1(_2355_));
 sg13g2_a21o_1 _3278_ (.A2(_2326_),
    .A1(_2318_),
    .B1(_2328_),
    .X(_2359_));
 sg13g2_o21ai_1 _3279_ (.B1(_2352_),
    .Y(_2360_),
    .A1(_2329_),
    .A2(_2353_));
 sg13g2_o21ai_1 _3280_ (.B1(_2324_),
    .Y(_2361_),
    .A1(net723),
    .A2(_2325_));
 sg13g2_o21ai_1 _3281_ (.B1(_2267_),
    .Y(_2362_),
    .A1(_1560_),
    .A2(_2252_));
 sg13g2_nand2_2 _3282_ (.Y(_2363_),
    .A(_2290_),
    .B(_2304_));
 sg13g2_or2_1 _3283_ (.X(_2364_),
    .B(net849),
    .A(net843));
 sg13g2_nand2_1 _3284_ (.Y(_2365_),
    .A(_2291_),
    .B(_2364_));
 sg13g2_mux2_1 _3285_ (.A0(_2277_),
    .A1(_2304_),
    .S(_2365_),
    .X(_2366_));
 sg13g2_o21ai_1 _3286_ (.B1(_2322_),
    .Y(_2367_),
    .A1(_2186_),
    .A2(_2291_));
 sg13g2_o21ai_1 _3287_ (.B1(_2363_),
    .Y(_2368_),
    .A1(_2366_),
    .A2(_2367_));
 sg13g2_xnor2_1 _3288_ (.Y(_2369_),
    .A(net723),
    .B(_2368_));
 sg13g2_nand2b_1 _3289_ (.Y(_2370_),
    .B(_2362_),
    .A_N(_2369_));
 sg13g2_xor2_1 _3290_ (.B(_2369_),
    .A(_2362_),
    .X(_2371_));
 sg13g2_nand2b_1 _3291_ (.Y(_2372_),
    .B(_2361_),
    .A_N(_2371_));
 sg13g2_xnor2_1 _3292_ (.Y(_2373_),
    .A(_2361_),
    .B(_2371_));
 sg13g2_a21oi_1 _3293_ (.A1(_2338_),
    .A2(_2350_),
    .Y(_2374_),
    .B1(_2349_));
 sg13g2_a21oi_1 _3294_ (.A1(_2335_),
    .A2(_2337_),
    .Y(_2375_),
    .B1(_2333_));
 sg13g2_a21oi_1 _3295_ (.A1(net818),
    .A2(_2335_),
    .Y(_2376_),
    .B1(_2333_));
 sg13g2_nand2_2 _3296_ (.Y(_2377_),
    .A(net802),
    .B(net837));
 sg13g2_nand2_2 _3297_ (.Y(_2378_),
    .A(net805),
    .B(net830));
 sg13g2_inv_1 _3298_ (.Y(_2379_),
    .A(_2378_));
 sg13g2_xor2_1 _3299_ (.B(_2378_),
    .A(_2331_),
    .X(_2380_));
 sg13g2_nand2b_1 _3300_ (.Y(_2381_),
    .B(_2380_),
    .A_N(_2377_));
 sg13g2_xnor2_1 _3301_ (.Y(_2382_),
    .A(_2377_),
    .B(_2380_));
 sg13g2_inv_1 _3302_ (.Y(_2383_),
    .A(_2382_));
 sg13g2_xnor2_1 _3303_ (.Y(_2384_),
    .A(_2376_),
    .B(_2382_));
 sg13g2_nand2b_1 _3304_ (.Y(_2385_),
    .B(_2384_),
    .A_N(_2375_));
 sg13g2_xor2_1 _3305_ (.B(_2384_),
    .A(_2375_),
    .X(_2386_));
 sg13g2_o21ai_1 _3306_ (.B1(_2345_),
    .Y(_2387_),
    .A1(_2346_),
    .A2(_2347_));
 sg13g2_a21o_1 _3307_ (.A2(_2343_),
    .A1(_2337_),
    .B1(_2342_),
    .X(_2388_));
 sg13g2_nand2b_1 _3308_ (.Y(_2389_),
    .B(net798),
    .A_N(net843));
 sg13g2_nor2_1 _3309_ (.A(_2377_),
    .B(_2389_),
    .Y(_2390_));
 sg13g2_xor2_1 _3310_ (.B(_2389_),
    .A(_2377_),
    .X(_2391_));
 sg13g2_xnor2_1 _3311_ (.Y(_2392_),
    .A(_2378_),
    .B(_2391_));
 sg13g2_nand2_1 _3312_ (.Y(_2393_),
    .A(_2388_),
    .B(_2392_));
 sg13g2_nor2_1 _3313_ (.A(_2388_),
    .B(_2392_),
    .Y(_2394_));
 sg13g2_xor2_1 _3314_ (.B(_2392_),
    .A(_2388_),
    .X(_2395_));
 sg13g2_xnor2_1 _3315_ (.Y(_2396_),
    .A(_2331_),
    .B(_2395_));
 sg13g2_nand2_1 _3316_ (.Y(_2397_),
    .A(_2387_),
    .B(_2396_));
 sg13g2_nor2_1 _3317_ (.A(_2387_),
    .B(_2396_),
    .Y(_2398_));
 sg13g2_xor2_1 _3318_ (.B(_2396_),
    .A(_2387_),
    .X(_2399_));
 sg13g2_xnor2_1 _3319_ (.Y(_2400_),
    .A(_2386_),
    .B(_2399_));
 sg13g2_nor2b_1 _3320_ (.A(_2374_),
    .B_N(_2400_),
    .Y(_2401_));
 sg13g2_xnor2_1 _3321_ (.Y(_2402_),
    .A(_2374_),
    .B(_2400_));
 sg13g2_xor2_1 _3322_ (.B(_2402_),
    .A(_2373_),
    .X(_2403_));
 sg13g2_nand2_1 _3323_ (.Y(_2404_),
    .A(_2360_),
    .B(_2403_));
 sg13g2_xnor2_1 _3324_ (.Y(_2405_),
    .A(_2360_),
    .B(_2403_));
 sg13g2_nand2b_1 _3325_ (.Y(_2406_),
    .B(_2359_),
    .A_N(_2405_));
 sg13g2_xor2_1 _3326_ (.B(_2405_),
    .A(_2359_),
    .X(_2407_));
 sg13g2_nand2_2 _3327_ (.Y(_2408_),
    .A(net800),
    .B(_2296_));
 sg13g2_xor2_1 _3328_ (.B(_2407_),
    .A(_2358_),
    .X(_2409_));
 sg13g2_nand2b_1 _3329_ (.Y(_2410_),
    .B(_2409_),
    .A_N(_2408_));
 sg13g2_o21ai_1 _3330_ (.B1(_2410_),
    .Y(_2411_),
    .A1(_2358_),
    .A2(_2407_));
 sg13g2_and2_1 _3331_ (.A(_2370_),
    .B(_2372_),
    .X(_2412_));
 sg13g2_a21o_1 _3332_ (.A2(_2402_),
    .A1(_2373_),
    .B1(_2401_),
    .X(_2413_));
 sg13g2_a22oi_1 _3333_ (.Y(_2414_),
    .B1(_2364_),
    .B2(_2277_),
    .A2(_2304_),
    .A1(_2291_));
 sg13g2_xnor2_1 _3334_ (.Y(_2415_),
    .A(net723),
    .B(_2414_));
 sg13g2_o21ai_1 _3335_ (.B1(_2385_),
    .Y(_2416_),
    .A1(_2376_),
    .A2(_2383_));
 sg13g2_nand2b_1 _3336_ (.Y(_2417_),
    .B(_2416_),
    .A_N(_2415_));
 sg13g2_xor2_1 _3337_ (.B(_2416_),
    .A(_2415_),
    .X(_2418_));
 sg13g2_o21ai_1 _3338_ (.B1(_2363_),
    .Y(_2419_),
    .A1(net723),
    .A2(_2368_));
 sg13g2_inv_1 _3339_ (.Y(_2420_),
    .A(_2419_));
 sg13g2_xnor2_1 _3340_ (.Y(_2421_),
    .A(_2418_),
    .B(_2419_));
 sg13g2_o21ai_1 _3341_ (.B1(_2397_),
    .Y(_2422_),
    .A1(_2386_),
    .A2(_2398_));
 sg13g2_o21ai_1 _3342_ (.B1(_2381_),
    .Y(_2423_),
    .A1(_1538_),
    .A2(_2252_));
 sg13g2_nand2_1 _3343_ (.Y(_2424_),
    .A(net798),
    .B(net837));
 sg13g2_nand2_1 _3344_ (.Y(_2425_),
    .A(net805),
    .B(net826));
 sg13g2_nand2_2 _3345_ (.Y(_2426_),
    .A(net802),
    .B(net830));
 sg13g2_nand2_1 _3346_ (.Y(_2427_),
    .A(net802),
    .B(net826));
 sg13g2_xor2_1 _3347_ (.B(_2426_),
    .A(_2425_),
    .X(_2428_));
 sg13g2_nand2b_1 _3348_ (.Y(_2429_),
    .B(_2428_),
    .A_N(_2424_));
 sg13g2_xnor2_1 _3349_ (.Y(_2430_),
    .A(_2424_),
    .B(_2428_));
 sg13g2_and2_1 _3350_ (.A(_1549_),
    .B(_2430_),
    .X(_2431_));
 sg13g2_xnor2_1 _3351_ (.Y(_2432_),
    .A(_1560_),
    .B(_2430_));
 sg13g2_xor2_1 _3352_ (.B(_2432_),
    .A(_2423_),
    .X(_2433_));
 sg13g2_o21ai_1 _3353_ (.B1(_2393_),
    .Y(_2434_),
    .A1(_2331_),
    .A2(_2394_));
 sg13g2_a21oi_1 _3354_ (.A1(_2379_),
    .A2(_2391_),
    .Y(_2435_),
    .B1(_2390_));
 sg13g2_nand2b_1 _3355_ (.Y(_2436_),
    .B(net798),
    .A_N(net839));
 sg13g2_xor2_1 _3356_ (.B(_2436_),
    .A(_2426_),
    .X(_2437_));
 sg13g2_nand2b_1 _3357_ (.Y(_2438_),
    .B(_2437_),
    .A_N(_2425_));
 sg13g2_xnor2_1 _3358_ (.Y(_2439_),
    .A(_2425_),
    .B(_2437_));
 sg13g2_nor2b_1 _3359_ (.A(_2435_),
    .B_N(_2439_),
    .Y(_2440_));
 sg13g2_xnor2_1 _3360_ (.Y(_2441_),
    .A(_2435_),
    .B(_2439_));
 sg13g2_xnor2_1 _3361_ (.Y(_2442_),
    .A(_0026_),
    .B(_2441_));
 sg13g2_and2_1 _3362_ (.A(_2434_),
    .B(_2442_),
    .X(_2443_));
 sg13g2_xor2_1 _3363_ (.B(_2442_),
    .A(_2434_),
    .X(_2444_));
 sg13g2_xor2_1 _3364_ (.B(_2444_),
    .A(_2433_),
    .X(_2445_));
 sg13g2_and2_1 _3365_ (.A(_2422_),
    .B(_2445_),
    .X(_2446_));
 sg13g2_xor2_1 _3366_ (.B(_2445_),
    .A(_2422_),
    .X(_2447_));
 sg13g2_xor2_1 _3367_ (.B(_2447_),
    .A(_2421_),
    .X(_2448_));
 sg13g2_nand2_1 _3368_ (.Y(_2449_),
    .A(_2413_),
    .B(_2448_));
 sg13g2_xnor2_1 _3369_ (.Y(_2450_),
    .A(_2413_),
    .B(_2448_));
 sg13g2_xnor2_1 _3370_ (.Y(_2451_),
    .A(_2412_),
    .B(_2450_));
 sg13g2_a21oi_1 _3371_ (.A1(_2404_),
    .A2(_2406_),
    .Y(_2452_),
    .B1(_2451_));
 sg13g2_and3_1 _3372_ (.X(_2453_),
    .A(_2404_),
    .B(_2406_),
    .C(_2451_));
 sg13g2_nor2_1 _3373_ (.A(_2452_),
    .B(_2453_),
    .Y(_2454_));
 sg13g2_xnor2_1 _3374_ (.Y(_2455_),
    .A(_2408_),
    .B(_2454_));
 sg13g2_and2_1 _3375_ (.A(_2411_),
    .B(_2455_),
    .X(_2456_));
 sg13g2_or2_1 _3376_ (.X(_2457_),
    .B(_2455_),
    .A(_2411_));
 sg13g2_nand2b_1 _3377_ (.Y(_2458_),
    .B(_2457_),
    .A_N(_2456_));
 sg13g2_nor2_2 _3378_ (.A(_1560_),
    .B(_2297_),
    .Y(_2459_));
 sg13g2_nand2_1 _3379_ (.Y(_2460_),
    .A(_1549_),
    .B(_2296_));
 sg13g2_a22oi_1 _3380_ (.Y(_2461_),
    .B1(net870),
    .B2(\system_inst.neuron.v[9] ),
    .A2(net863),
    .A1(net821));
 sg13g2_nor2_2 _3381_ (.A(_2459_),
    .B(_2461_),
    .Y(_2462_));
 sg13g2_inv_1 _3382_ (.Y(_2463_),
    .A(_2462_));
 sg13g2_nand2_2 _3383_ (.Y(_2464_),
    .A(net828),
    .B(net856));
 sg13g2_nand2_2 _3384_ (.Y(_2465_),
    .A(net823),
    .B(net861));
 sg13g2_nand2_1 _3385_ (.Y(_2466_),
    .A(net834),
    .B(net847));
 sg13g2_xor2_1 _3386_ (.B(_2465_),
    .A(_2464_),
    .X(_2467_));
 sg13g2_nand2b_1 _3387_ (.Y(_2468_),
    .B(_2467_),
    .A_N(_2466_));
 sg13g2_o21ai_1 _3388_ (.B1(_2468_),
    .Y(_2469_),
    .A1(_2464_),
    .A2(_2465_));
 sg13g2_nand2_2 _3389_ (.Y(_2470_),
    .A(net834),
    .B(net841));
 sg13g2_and4_1 _3390_ (.A(net823),
    .B(net829),
    .C(net848),
    .D(net856),
    .X(_2471_));
 sg13g2_a22oi_1 _3391_ (.Y(_2472_),
    .B1(net856),
    .B2(net823),
    .A2(net848),
    .A1(net829));
 sg13g2_nor3_1 _3392_ (.A(_2470_),
    .B(_2471_),
    .C(_2472_),
    .Y(_2473_));
 sg13g2_o21ai_1 _3393_ (.B1(_2470_),
    .Y(_2474_),
    .A1(_2471_),
    .A2(_2472_));
 sg13g2_nor2b_2 _3394_ (.A(_2473_),
    .B_N(_2474_),
    .Y(_2475_));
 sg13g2_nand2_1 _3395_ (.Y(_2476_),
    .A(_2469_),
    .B(_2475_));
 sg13g2_xnor2_1 _3396_ (.Y(_2477_),
    .A(_2469_),
    .B(_2475_));
 sg13g2_nor2_1 _3397_ (.A(_2463_),
    .B(_2477_),
    .Y(_2478_));
 sg13g2_and2_2 _3398_ (.A(net820),
    .B(net856),
    .X(_2479_));
 sg13g2_nand2_2 _3399_ (.Y(_2480_),
    .A(net810),
    .B(net864));
 sg13g2_and4_2 _3400_ (.A(net809),
    .B(net816),
    .C(net863),
    .D(net870),
    .X(_2481_));
 sg13g2_a22oi_1 _3401_ (.Y(_2482_),
    .B1(net870),
    .B2(net809),
    .A2(net863),
    .A1(net816));
 sg13g2_nor2_2 _3402_ (.A(_2481_),
    .B(_2482_),
    .Y(_2483_));
 sg13g2_inv_1 _3403_ (.Y(_2484_),
    .A(_2483_));
 sg13g2_xnor2_1 _3404_ (.Y(_2485_),
    .A(_2479_),
    .B(_2483_));
 sg13g2_or2_2 _3405_ (.X(_2486_),
    .B(_2473_),
    .A(_2471_));
 sg13g2_nor2_1 _3406_ (.A(_2252_),
    .B(_2291_),
    .Y(_2487_));
 sg13g2_a22oi_1 _3407_ (.Y(_2488_),
    .B1(net848),
    .B2(net824),
    .A2(net842),
    .A1(net829));
 sg13g2_a21oi_2 _3408_ (.B1(_2488_),
    .Y(_2489_),
    .A2(_2290_),
    .A1(_2251_));
 sg13g2_xnor2_1 _3409_ (.Y(_2490_),
    .A(net836),
    .B(_2489_));
 sg13g2_nor2_1 _3410_ (.A(_2460_),
    .B(_2490_),
    .Y(_2491_));
 sg13g2_xnor2_1 _3411_ (.Y(_2492_),
    .A(_2459_),
    .B(_2490_));
 sg13g2_xnor2_1 _3412_ (.Y(_2493_),
    .A(_2486_),
    .B(_2492_));
 sg13g2_or2_1 _3413_ (.X(_2494_),
    .B(_2493_),
    .A(_2485_));
 sg13g2_xnor2_1 _3414_ (.Y(_2495_),
    .A(_2485_),
    .B(_2493_));
 sg13g2_or3_1 _3415_ (.A(_2463_),
    .B(_2477_),
    .C(_2495_),
    .X(_2496_));
 sg13g2_xor2_1 _3416_ (.B(_2495_),
    .A(_2478_),
    .X(_2497_));
 sg13g2_a21o_1 _3417_ (.A2(net848),
    .A1(net833),
    .B1(_0029_),
    .X(_2498_));
 sg13g2_nand3_1 _3418_ (.B(net848),
    .C(_0029_),
    .A(net833),
    .Y(_2499_));
 sg13g2_a21oi_2 _3419_ (.B1(_2464_),
    .Y(_2500_),
    .A2(_2499_),
    .A1(_2498_));
 sg13g2_a21oi_1 _3420_ (.A1(net836),
    .A2(_2290_),
    .Y(_2501_),
    .B1(_2500_));
 sg13g2_nor2b_1 _3421_ (.A(_2501_),
    .B_N(_2475_),
    .Y(_2502_));
 sg13g2_xnor2_1 _3422_ (.Y(_2503_),
    .A(_2475_),
    .B(_2501_));
 sg13g2_a21oi_1 _3423_ (.A1(_2462_),
    .A2(_2503_),
    .Y(_2504_),
    .B1(_2502_));
 sg13g2_xor2_1 _3424_ (.B(_2489_),
    .A(_2479_),
    .X(_2505_));
 sg13g2_nand2_1 _3425_ (.Y(_2506_),
    .A(_2486_),
    .B(_2505_));
 sg13g2_xnor2_1 _3426_ (.Y(_2507_),
    .A(_2486_),
    .B(_2505_));
 sg13g2_xnor2_1 _3427_ (.Y(_2508_),
    .A(_2484_),
    .B(_2507_));
 sg13g2_xor2_1 _3428_ (.B(_2508_),
    .A(_2476_),
    .X(_2509_));
 sg13g2_nand2b_1 _3429_ (.Y(_2510_),
    .B(_2509_),
    .A_N(_2504_));
 sg13g2_xor2_1 _3430_ (.B(_2509_),
    .A(_2504_),
    .X(_2511_));
 sg13g2_o21ai_1 _3431_ (.B1(_2496_),
    .Y(_2512_),
    .A1(_2497_),
    .A2(_2511_));
 sg13g2_o21ai_1 _3432_ (.B1(_2506_),
    .Y(_2513_),
    .A1(_2484_),
    .A2(_2507_));
 sg13g2_a21o_1 _3433_ (.A2(_2492_),
    .A1(_2486_),
    .B1(_2491_),
    .X(_2514_));
 sg13g2_nor2_1 _3434_ (.A(_1538_),
    .B(_2297_),
    .Y(_2515_));
 sg13g2_xor2_1 _3435_ (.B(_2480_),
    .A(_2215_),
    .X(_2516_));
 sg13g2_a21oi_1 _3436_ (.A1(_2479_),
    .A2(_2489_),
    .Y(_2517_),
    .B1(_2487_));
 sg13g2_nand2_2 _3437_ (.Y(_2518_),
    .A(net816),
    .B(net857));
 sg13g2_nand2_2 _3438_ (.Y(_2519_),
    .A(net820),
    .B(net848));
 sg13g2_nand2_2 _3439_ (.Y(_2520_),
    .A(net824),
    .B(net842));
 sg13g2_xor2_1 _3440_ (.B(_2520_),
    .A(_2519_),
    .X(_2521_));
 sg13g2_nand2b_1 _3441_ (.Y(_2522_),
    .B(_2521_),
    .A_N(_2518_));
 sg13g2_xnor2_1 _3442_ (.Y(_2523_),
    .A(_2518_),
    .B(_2521_));
 sg13g2_nor2b_1 _3443_ (.A(_2517_),
    .B_N(_2523_),
    .Y(_2524_));
 sg13g2_xnor2_1 _3444_ (.Y(_2525_),
    .A(_2517_),
    .B(_2523_));
 sg13g2_xor2_1 _3445_ (.B(_2525_),
    .A(_2516_),
    .X(_2526_));
 sg13g2_xnor2_1 _3446_ (.Y(_2527_),
    .A(_2514_),
    .B(_2526_));
 sg13g2_nor2b_1 _3447_ (.A(_2527_),
    .B_N(_2513_),
    .Y(_2528_));
 sg13g2_xor2_1 _3448_ (.B(_2527_),
    .A(_2513_),
    .X(_2529_));
 sg13g2_nand2_1 _3449_ (.Y(_2530_),
    .A(net810),
    .B(net856));
 sg13g2_xor2_1 _3450_ (.B(_2518_),
    .A(_2480_),
    .X(_2531_));
 sg13g2_nand2b_1 _3451_ (.Y(_2532_),
    .B(_2531_),
    .A_N(_2519_));
 sg13g2_xnor2_1 _3452_ (.Y(_2533_),
    .A(_2519_),
    .B(_2531_));
 sg13g2_nand2b_1 _3453_ (.Y(_2534_),
    .B(_2533_),
    .A_N(_2215_));
 sg13g2_xnor2_1 _3454_ (.Y(_2535_),
    .A(_2215_),
    .B(_2533_));
 sg13g2_a21oi_1 _3455_ (.A1(net836),
    .A2(_2489_),
    .Y(_2536_),
    .B1(_2487_));
 sg13g2_a21oi_1 _3456_ (.A1(_2479_),
    .A2(_2483_),
    .Y(_2537_),
    .B1(_2481_));
 sg13g2_xor2_1 _3457_ (.B(_2537_),
    .A(_2520_),
    .X(_2538_));
 sg13g2_nand2b_1 _3458_ (.Y(_2539_),
    .B(_2538_),
    .A_N(_2536_));
 sg13g2_xnor2_1 _3459_ (.Y(_2540_),
    .A(_2536_),
    .B(_2538_));
 sg13g2_nand2_1 _3460_ (.Y(_2541_),
    .A(_2535_),
    .B(_2540_));
 sg13g2_xnor2_1 _3461_ (.Y(_2542_),
    .A(_2535_),
    .B(_2540_));
 sg13g2_nor2_1 _3462_ (.A(_2494_),
    .B(_2542_),
    .Y(_2543_));
 sg13g2_xor2_1 _3463_ (.B(_2542_),
    .A(_2494_),
    .X(_2544_));
 sg13g2_nor2b_1 _3464_ (.A(_2529_),
    .B_N(_2544_),
    .Y(_2545_));
 sg13g2_xnor2_1 _3465_ (.Y(_2546_),
    .A(_2529_),
    .B(_2544_));
 sg13g2_o21ai_1 _3466_ (.B1(_2510_),
    .Y(_2547_),
    .A1(_2476_),
    .A2(_2508_));
 sg13g2_xnor2_1 _3467_ (.Y(_2548_),
    .A(_2512_),
    .B(_2546_));
 sg13g2_nor2b_1 _3468_ (.A(_2548_),
    .B_N(_2547_),
    .Y(_2549_));
 sg13g2_a21oi_2 _3469_ (.B1(_2549_),
    .Y(_2550_),
    .A2(_2546_),
    .A1(_2512_));
 sg13g2_a21o_1 _3470_ (.A2(_2526_),
    .A1(_2514_),
    .B1(_2528_),
    .X(_2551_));
 sg13g2_nor2_1 _3471_ (.A(_2543_),
    .B(_2545_),
    .Y(_2552_));
 sg13g2_a22oi_1 _3472_ (.Y(_2553_),
    .B1(net869),
    .B2(net802),
    .A2(net864),
    .A1(net805));
 sg13g2_nor2_2 _3473_ (.A(_2216_),
    .B(_2553_),
    .Y(_2554_));
 sg13g2_nand2_1 _3474_ (.Y(_2555_),
    .A(_1549_),
    .B(_2290_));
 sg13g2_a22oi_1 _3475_ (.Y(_2556_),
    .B1(net849),
    .B2(net814),
    .A2(net843),
    .A1(net818));
 sg13g2_a21oi_1 _3476_ (.A1(_1549_),
    .A2(_2290_),
    .Y(_2557_),
    .B1(_2556_));
 sg13g2_xnor2_1 _3477_ (.Y(_2558_),
    .A(_2530_),
    .B(_2557_));
 sg13g2_nand2_1 _3478_ (.Y(_2559_),
    .A(_2554_),
    .B(_2558_));
 sg13g2_xnor2_1 _3479_ (.Y(_2560_),
    .A(_2554_),
    .B(_2558_));
 sg13g2_nor2_1 _3480_ (.A(_2534_),
    .B(_2560_),
    .Y(_2561_));
 sg13g2_xor2_1 _3481_ (.B(_2560_),
    .A(_2534_),
    .X(_2562_));
 sg13g2_and2_2 _3482_ (.A(net827),
    .B(net833),
    .X(_2563_));
 sg13g2_nand2_2 _3483_ (.Y(_2564_),
    .A(net829),
    .B(net836));
 sg13g2_o21ai_1 _3484_ (.B1(_2532_),
    .Y(_2565_),
    .A1(_2480_),
    .A2(_2518_));
 sg13g2_nor2b_1 _3485_ (.A(_0027_),
    .B_N(_2565_),
    .Y(_2566_));
 sg13g2_xnor2_1 _3486_ (.Y(_2567_),
    .A(_0027_),
    .B(_2565_));
 sg13g2_xnor2_1 _3487_ (.Y(_2568_),
    .A(_2564_),
    .B(_2567_));
 sg13g2_xnor2_1 _3488_ (.Y(_2569_),
    .A(_2562_),
    .B(_2568_));
 sg13g2_nor2_1 _3489_ (.A(_2541_),
    .B(_2569_),
    .Y(_2570_));
 sg13g2_xor2_1 _3490_ (.B(_2569_),
    .A(_2541_),
    .X(_2571_));
 sg13g2_a21o_1 _3491_ (.A2(_2525_),
    .A1(_2516_),
    .B1(_2524_),
    .X(_2572_));
 sg13g2_o21ai_1 _3492_ (.B1(_2539_),
    .Y(_2573_),
    .A1(_2520_),
    .A2(_2537_));
 sg13g2_o21ai_1 _3493_ (.B1(_2522_),
    .Y(_2574_),
    .A1(_2519_),
    .A2(_2520_));
 sg13g2_and2_1 _3494_ (.A(_2558_),
    .B(_2574_),
    .X(_2575_));
 sg13g2_xor2_1 _3495_ (.B(_2574_),
    .A(_2558_),
    .X(_2576_));
 sg13g2_xnor2_1 _3496_ (.Y(_2577_),
    .A(_2554_),
    .B(_2576_));
 sg13g2_nand2b_1 _3497_ (.Y(_2578_),
    .B(_2573_),
    .A_N(_2577_));
 sg13g2_xor2_1 _3498_ (.B(_2577_),
    .A(_2573_),
    .X(_2579_));
 sg13g2_nand2b_1 _3499_ (.Y(_2580_),
    .B(_2572_),
    .A_N(_2579_));
 sg13g2_xnor2_1 _3500_ (.Y(_2581_),
    .A(_2572_),
    .B(_2579_));
 sg13g2_xnor2_1 _3501_ (.Y(_2582_),
    .A(_2571_),
    .B(_2581_));
 sg13g2_nor2_1 _3502_ (.A(_2552_),
    .B(_2582_),
    .Y(_2583_));
 sg13g2_xor2_1 _3503_ (.B(_2582_),
    .A(_2552_),
    .X(_2584_));
 sg13g2_xnor2_1 _3504_ (.Y(_2585_),
    .A(_2551_),
    .B(_2584_));
 sg13g2_nor2_1 _3505_ (.A(_2550_),
    .B(_2585_),
    .Y(_2586_));
 sg13g2_xor2_1 _3506_ (.B(_2585_),
    .A(_2550_),
    .X(_2587_));
 sg13g2_a21oi_1 _3507_ (.A1(_2515_),
    .A2(_2587_),
    .Y(_2588_),
    .B1(_2586_));
 sg13g2_a21oi_2 _3508_ (.B1(_2583_),
    .Y(_2589_),
    .A2(_2584_),
    .A1(_2551_));
 sg13g2_nand2_1 _3509_ (.Y(_2590_),
    .A(_2578_),
    .B(_2580_));
 sg13g2_a21oi_1 _3510_ (.A1(_2571_),
    .A2(_2581_),
    .Y(_2591_),
    .B1(_2570_));
 sg13g2_a21o_1 _3511_ (.A2(_2576_),
    .A1(_2554_),
    .B1(_2575_),
    .X(_2592_));
 sg13g2_a21oi_1 _3512_ (.A1(_2563_),
    .A2(_2567_),
    .Y(_2593_),
    .B1(_2566_));
 sg13g2_o21ai_1 _3513_ (.B1(_2555_),
    .Y(_2594_),
    .A1(_2530_),
    .A2(_2556_));
 sg13g2_xnor2_1 _3514_ (.Y(_2595_),
    .A(_2217_),
    .B(_2227_));
 sg13g2_nand2_1 _3515_ (.Y(_2596_),
    .A(_2594_),
    .B(_2595_));
 sg13g2_xnor2_1 _3516_ (.Y(_2597_),
    .A(_2594_),
    .B(_2595_));
 sg13g2_xnor2_1 _3517_ (.Y(_2598_),
    .A(_2220_),
    .B(_2597_));
 sg13g2_nor2_1 _3518_ (.A(_2593_),
    .B(_2598_),
    .Y(_2599_));
 sg13g2_xor2_1 _3519_ (.B(_2598_),
    .A(_2593_),
    .X(_2600_));
 sg13g2_xor2_1 _3520_ (.B(_2600_),
    .A(_2592_),
    .X(_2601_));
 sg13g2_a21oi_1 _3521_ (.A1(_2562_),
    .A2(_2568_),
    .Y(_2602_),
    .B1(_2561_));
 sg13g2_xnor2_1 _3522_ (.Y(_2603_),
    .A(_2223_),
    .B(_2230_));
 sg13g2_nor2_1 _3523_ (.A(_2559_),
    .B(_2603_),
    .Y(_2604_));
 sg13g2_xor2_1 _3524_ (.B(_2603_),
    .A(_2559_),
    .X(_2605_));
 sg13g2_nand2_1 _3525_ (.Y(_2606_),
    .A(net825),
    .B(net837));
 sg13g2_nand2b_1 _3526_ (.Y(_2607_),
    .B(_2594_),
    .A_N(_2228_));
 sg13g2_xnor2_1 _3527_ (.Y(_2608_),
    .A(_2228_),
    .B(_2594_));
 sg13g2_nand2b_1 _3528_ (.Y(_2609_),
    .B(_2608_),
    .A_N(_2606_));
 sg13g2_xnor2_1 _3529_ (.Y(_2610_),
    .A(_2606_),
    .B(_2608_));
 sg13g2_xnor2_1 _3530_ (.Y(_2611_),
    .A(_2605_),
    .B(_2610_));
 sg13g2_nor2_1 _3531_ (.A(_2602_),
    .B(_2611_),
    .Y(_2612_));
 sg13g2_xor2_1 _3532_ (.B(_2611_),
    .A(_2602_),
    .X(_2613_));
 sg13g2_xor2_1 _3533_ (.B(_2613_),
    .A(_2601_),
    .X(_2614_));
 sg13g2_nor2b_1 _3534_ (.A(_2591_),
    .B_N(_2614_),
    .Y(_2615_));
 sg13g2_xnor2_1 _3535_ (.Y(_2616_),
    .A(_2591_),
    .B(_2614_));
 sg13g2_xnor2_1 _3536_ (.Y(_2617_),
    .A(_2590_),
    .B(_2616_));
 sg13g2_nor2_1 _3537_ (.A(_2589_),
    .B(_2617_),
    .Y(_2618_));
 sg13g2_xor2_1 _3538_ (.B(_2617_),
    .A(_2589_),
    .X(_2619_));
 sg13g2_and2_1 _3539_ (.A(_2216_),
    .B(_2619_),
    .X(_2620_));
 sg13g2_xor2_1 _3540_ (.B(_2619_),
    .A(_2216_),
    .X(_2621_));
 sg13g2_nor2b_1 _3541_ (.A(_2588_),
    .B_N(_2621_),
    .Y(_2622_));
 sg13g2_xnor2_1 _3542_ (.Y(_2623_),
    .A(_2588_),
    .B(_2621_));
 sg13g2_xor2_1 _3543_ (.B(_2587_),
    .A(_2515_),
    .X(_2624_));
 sg13g2_nand2_2 _3544_ (.Y(_2625_),
    .A(net821),
    .B(net870));
 sg13g2_and4_2 _3545_ (.A(net823),
    .B(net827),
    .C(net862),
    .D(net867),
    .X(_2626_));
 sg13g2_nand2_2 _3546_ (.Y(_2627_),
    .A(_2251_),
    .B(_2296_));
 sg13g2_nand2_1 _3547_ (.Y(_2628_),
    .A(net833),
    .B(net854));
 sg13g2_a22oi_1 _3548_ (.Y(_2629_),
    .B1(net867),
    .B2(net823),
    .A2(net862),
    .A1(net828));
 sg13g2_or2_2 _3549_ (.X(_2630_),
    .B(_2629_),
    .A(_2626_));
 sg13g2_nor2_1 _3550_ (.A(_2628_),
    .B(_2630_),
    .Y(_2631_));
 sg13g2_xnor2_1 _3551_ (.Y(_2632_),
    .A(_2466_),
    .B(_2467_));
 sg13g2_o21ai_1 _3552_ (.B1(_2632_),
    .Y(_2633_),
    .A1(_2626_),
    .A2(_2631_));
 sg13g2_or3_1 _3553_ (.A(_2626_),
    .B(_2631_),
    .C(_2632_),
    .X(_2634_));
 sg13g2_and2_1 _3554_ (.A(_2633_),
    .B(_2634_),
    .X(_2635_));
 sg13g2_nand2b_1 _3555_ (.Y(_2636_),
    .B(_2635_),
    .A_N(_2625_));
 sg13g2_xnor2_1 _3556_ (.Y(_2637_),
    .A(_2463_),
    .B(_2477_));
 sg13g2_or2_1 _3557_ (.X(_2638_),
    .B(_2637_),
    .A(_2636_));
 sg13g2_xnor2_1 _3558_ (.Y(_2639_),
    .A(_2636_),
    .B(_2637_));
 sg13g2_and3_1 _3559_ (.X(_2640_),
    .A(_2464_),
    .B(_2498_),
    .C(_2499_));
 sg13g2_or3_1 _3560_ (.A(_2291_),
    .B(_2500_),
    .C(_2640_),
    .X(_2641_));
 sg13g2_o21ai_1 _3561_ (.B1(_2291_),
    .Y(_2642_),
    .A1(_2500_),
    .A2(_2640_));
 sg13g2_nand2_1 _3562_ (.Y(_2643_),
    .A(_2254_),
    .B(_2296_));
 sg13g2_xor2_1 _3563_ (.B(_2625_),
    .A(_2465_),
    .X(_2644_));
 sg13g2_nand3_1 _3564_ (.B(_2642_),
    .C(_2644_),
    .A(_2641_),
    .Y(_2645_));
 sg13g2_and2_1 _3565_ (.A(_2641_),
    .B(_2645_),
    .X(_2646_));
 sg13g2_xnor2_1 _3566_ (.Y(_2647_),
    .A(_2462_),
    .B(_2503_));
 sg13g2_xor2_1 _3567_ (.B(_2647_),
    .A(_2633_),
    .X(_2648_));
 sg13g2_nand2b_1 _3568_ (.Y(_2649_),
    .B(_2648_),
    .A_N(_2646_));
 sg13g2_xor2_1 _3569_ (.B(_2648_),
    .A(_2646_),
    .X(_2650_));
 sg13g2_o21ai_1 _3570_ (.B1(_2638_),
    .Y(_2651_),
    .A1(_2639_),
    .A2(_2650_));
 sg13g2_xor2_1 _3571_ (.B(_2511_),
    .A(_2497_),
    .X(_2652_));
 sg13g2_and2_1 _3572_ (.A(_2651_),
    .B(_2652_),
    .X(_2653_));
 sg13g2_o21ai_1 _3573_ (.B1(_2649_),
    .Y(_2654_),
    .A1(_2633_),
    .A2(_2647_));
 sg13g2_xor2_1 _3574_ (.B(_2652_),
    .A(_2651_),
    .X(_2655_));
 sg13g2_a21oi_2 _3575_ (.B1(_2653_),
    .Y(_2656_),
    .A2(_2655_),
    .A1(_2654_));
 sg13g2_xor2_1 _3576_ (.B(_2548_),
    .A(_2547_),
    .X(_2657_));
 sg13g2_xor2_1 _3577_ (.B(_2657_),
    .A(_2656_),
    .X(_2658_));
 sg13g2_nand2_1 _3578_ (.Y(_2659_),
    .A(_2481_),
    .B(_2658_));
 sg13g2_o21ai_1 _3579_ (.B1(_2659_),
    .Y(_2660_),
    .A1(_2656_),
    .A2(_2657_));
 sg13g2_and2_1 _3580_ (.A(_2624_),
    .B(_2660_),
    .X(_2661_));
 sg13g2_xnor2_1 _3581_ (.Y(_2662_),
    .A(_2624_),
    .B(_2660_));
 sg13g2_xnor2_1 _3582_ (.Y(_2663_),
    .A(_2625_),
    .B(_2635_));
 sg13g2_o21ai_1 _3583_ (.B1(net854),
    .Y(_2664_),
    .A1(net833),
    .A2(net841));
 sg13g2_nand2b_1 _3584_ (.Y(_2665_),
    .B(_2470_),
    .A_N(_2664_));
 sg13g2_nand3_1 _3585_ (.B(net841),
    .C(net854),
    .A(net833),
    .Y(_2666_));
 sg13g2_o21ai_1 _3586_ (.B1(_2666_),
    .Y(_2667_),
    .A1(_2630_),
    .A2(_2665_));
 sg13g2_inv_1 _3587_ (.Y(_2668_),
    .A(_2667_));
 sg13g2_nor2_2 _3588_ (.A(_2297_),
    .B(_2564_),
    .Y(_2669_));
 sg13g2_nand2_2 _3589_ (.Y(_2670_),
    .A(_2296_),
    .B(_2563_));
 sg13g2_xor2_1 _3590_ (.B(_2630_),
    .A(_2628_),
    .X(_2671_));
 sg13g2_and2_1 _3591_ (.A(_2669_),
    .B(_2671_),
    .X(_2672_));
 sg13g2_a21o_1 _3592_ (.A2(_2642_),
    .A1(_2641_),
    .B1(_2644_),
    .X(_2673_));
 sg13g2_and3_1 _3593_ (.X(_2674_),
    .A(_2645_),
    .B(_2672_),
    .C(_2673_));
 sg13g2_a21oi_1 _3594_ (.A1(_2645_),
    .A2(_2673_),
    .Y(_2675_),
    .B1(_2672_));
 sg13g2_o21ai_1 _3595_ (.B1(_2668_),
    .Y(_2676_),
    .A1(_2674_),
    .A2(_2675_));
 sg13g2_or3_1 _3596_ (.A(_2668_),
    .B(_2674_),
    .C(_2675_),
    .X(_2677_));
 sg13g2_and3_1 _3597_ (.X(_2678_),
    .A(_2663_),
    .B(_2676_),
    .C(_2677_));
 sg13g2_xor2_1 _3598_ (.B(_2650_),
    .A(_2639_),
    .X(_2679_));
 sg13g2_nand2_1 _3599_ (.Y(_2680_),
    .A(_2678_),
    .B(_2679_));
 sg13g2_nor2b_1 _3600_ (.A(_2674_),
    .B_N(_2677_),
    .Y(_2681_));
 sg13g2_xnor2_1 _3601_ (.Y(_2682_),
    .A(_2678_),
    .B(_2679_));
 sg13g2_o21ai_1 _3602_ (.B1(_2680_),
    .Y(_2683_),
    .A1(_2681_),
    .A2(_2682_));
 sg13g2_xnor2_1 _3603_ (.Y(_2684_),
    .A(_2654_),
    .B(_2655_));
 sg13g2_nand2b_1 _3604_ (.Y(_2685_),
    .B(_2683_),
    .A_N(_2684_));
 sg13g2_xor2_1 _3605_ (.B(_2684_),
    .A(_2683_),
    .X(_2686_));
 sg13g2_o21ai_1 _3606_ (.B1(_2685_),
    .Y(_2687_),
    .A1(_2460_),
    .A2(_2686_));
 sg13g2_inv_1 _3607_ (.Y(_2688_),
    .A(_2687_));
 sg13g2_xor2_1 _3608_ (.B(_2658_),
    .A(_2481_),
    .X(_2689_));
 sg13g2_inv_1 _3609_ (.Y(_2690_),
    .A(_2689_));
 sg13g2_xnor2_1 _3610_ (.Y(_2691_),
    .A(_2459_),
    .B(_2686_));
 sg13g2_xnor2_1 _3611_ (.Y(_2692_),
    .A(_2670_),
    .B(_2671_));
 sg13g2_xnor2_1 _3612_ (.Y(_2693_),
    .A(_2630_),
    .B(_2665_));
 sg13g2_a22oi_1 _3613_ (.Y(_2694_),
    .B1(net867),
    .B2(net828),
    .A2(net862),
    .A1(net833));
 sg13g2_nor2_2 _3614_ (.A(_2669_),
    .B(_2694_),
    .Y(_2695_));
 sg13g2_o21ai_1 _3615_ (.B1(net847),
    .Y(_2696_),
    .A1(net854),
    .A2(_2695_));
 sg13g2_or2_1 _3616_ (.X(_2697_),
    .B(_2696_),
    .A(_2693_));
 sg13g2_inv_1 _3617_ (.Y(_2698_),
    .A(_2697_));
 sg13g2_xor2_1 _3618_ (.B(_2696_),
    .A(_2693_),
    .X(_2699_));
 sg13g2_nand2_1 _3619_ (.Y(_2700_),
    .A(_2692_),
    .B(_2699_));
 sg13g2_a21oi_1 _3620_ (.A1(_2676_),
    .A2(_2677_),
    .Y(_2701_),
    .B1(_2663_));
 sg13g2_or3_1 _3621_ (.A(_2678_),
    .B(_2700_),
    .C(_2701_),
    .X(_2702_));
 sg13g2_o21ai_1 _3622_ (.B1(_2700_),
    .Y(_2703_),
    .A1(_2678_),
    .A2(_2701_));
 sg13g2_nand3_1 _3623_ (.B(_2702_),
    .C(_2703_),
    .A(_2698_),
    .Y(_2704_));
 sg13g2_and2_1 _3624_ (.A(_2702_),
    .B(_2704_),
    .X(_2705_));
 sg13g2_xor2_1 _3625_ (.B(_2682_),
    .A(_2681_),
    .X(_2706_));
 sg13g2_nand2b_1 _3626_ (.Y(_2707_),
    .B(_2706_),
    .A_N(_2705_));
 sg13g2_nor2b_1 _3627_ (.A(_2706_),
    .B_N(_2705_),
    .Y(_2708_));
 sg13g2_xnor2_1 _3628_ (.Y(_2709_),
    .A(_2705_),
    .B(_2706_));
 sg13g2_o21ai_1 _3629_ (.B1(_2707_),
    .Y(_2710_),
    .A1(_2643_),
    .A2(_2708_));
 sg13g2_nand2_1 _3630_ (.Y(_2711_),
    .A(_2691_),
    .B(_2710_));
 sg13g2_xor2_1 _3631_ (.B(_2710_),
    .A(_2691_),
    .X(_2712_));
 sg13g2_and2_1 _3632_ (.A(net841),
    .B(net861),
    .X(_2713_));
 sg13g2_a22oi_1 _3633_ (.Y(_2714_),
    .B1(net867),
    .B2(net841),
    .A2(net861),
    .A1(net847));
 sg13g2_and4_1 _3634_ (.A(net841),
    .B(net847),
    .C(net861),
    .D(net867),
    .X(_2715_));
 sg13g2_nand4_1 _3635_ (.B(net847),
    .C(net861),
    .A(net840),
    .Y(_2716_),
    .D(net867));
 sg13g2_a21oi_2 _3636_ (.B1(_2714_),
    .Y(_2717_),
    .A2(_2716_),
    .A1(_1406_));
 sg13g2_nand2_2 _3637_ (.Y(_2718_),
    .A(net833),
    .B(net867));
 sg13g2_or2_1 _3638_ (.X(_2719_),
    .B(_2470_),
    .A(_2297_));
 sg13g2_mux2_1 _3639_ (.A0(_2717_),
    .A1(_2713_),
    .S(_2718_),
    .X(_2720_));
 sg13g2_xnor2_1 _3640_ (.Y(_2721_),
    .A(_2275_),
    .B(_2695_));
 sg13g2_inv_1 _3641_ (.Y(_2722_),
    .A(_2721_));
 sg13g2_nand2_1 _3642_ (.Y(_2723_),
    .A(_2720_),
    .B(_2722_));
 sg13g2_xnor2_1 _3643_ (.Y(_2724_),
    .A(_2720_),
    .B(_2721_));
 sg13g2_nand2_1 _3644_ (.Y(_2725_),
    .A(_2695_),
    .B(_2724_));
 sg13g2_xnor2_1 _3645_ (.Y(_2726_),
    .A(_2692_),
    .B(_2699_));
 sg13g2_xor2_1 _3646_ (.B(_2726_),
    .A(_2725_),
    .X(_2727_));
 sg13g2_a21oi_2 _3647_ (.B1(_2726_),
    .Y(_2728_),
    .A2(_2725_),
    .A1(_2723_));
 sg13g2_a21o_1 _3648_ (.A2(_2703_),
    .A1(_2702_),
    .B1(_2698_),
    .X(_2729_));
 sg13g2_nand3_1 _3649_ (.B(_2728_),
    .C(_2729_),
    .A(_2704_),
    .Y(_2730_));
 sg13g2_a21oi_1 _3650_ (.A1(_2704_),
    .A2(_2729_),
    .Y(_2731_),
    .B1(_2728_));
 sg13g2_a21o_1 _3651_ (.A2(_2729_),
    .A1(_2704_),
    .B1(_2728_),
    .X(_2732_));
 sg13g2_and3_1 _3652_ (.X(_2733_),
    .A(_2626_),
    .B(_2730_),
    .C(_2732_));
 sg13g2_o21ai_1 _3653_ (.B1(_2730_),
    .Y(_2734_),
    .A1(_2627_),
    .A2(_2731_));
 sg13g2_xnor2_1 _3654_ (.Y(_2735_),
    .A(_2643_),
    .B(_2709_));
 sg13g2_nor2_1 _3655_ (.A(_2734_),
    .B(_2735_),
    .Y(_2736_));
 sg13g2_or2_1 _3656_ (.X(_2737_),
    .B(_2735_),
    .A(_2734_));
 sg13g2_xnor2_1 _3657_ (.Y(_2738_),
    .A(_2275_),
    .B(_2720_));
 sg13g2_xor2_1 _3658_ (.B(_2718_),
    .A(_2717_),
    .X(_2739_));
 sg13g2_nor3_1 _3659_ (.A(net855),
    .B(_2714_),
    .C(_2715_),
    .Y(_2740_));
 sg13g2_nor2_1 _3660_ (.A(_1395_),
    .B(_1417_),
    .Y(_2741_));
 sg13g2_nand3_1 _3661_ (.B(net861),
    .C(net867),
    .A(net847),
    .Y(_2742_));
 sg13g2_nand2_1 _3662_ (.Y(_2743_),
    .A(net855),
    .B(_2296_));
 sg13g2_and2_1 _3663_ (.A(net855),
    .B(_2742_),
    .X(_2744_));
 sg13g2_o21ai_1 _3664_ (.B1(_2744_),
    .Y(_2745_),
    .A1(net861),
    .A2(_2741_));
 sg13g2_o21ai_1 _3665_ (.B1(_2745_),
    .Y(_2746_),
    .A1(net854),
    .A2(_2741_));
 sg13g2_or2_1 _3666_ (.X(_2747_),
    .B(_2742_),
    .A(_1406_));
 sg13g2_nor2b_2 _3667_ (.A(_2740_),
    .B_N(_2747_),
    .Y(_2748_));
 sg13g2_nor2_1 _3668_ (.A(_2739_),
    .B(_2748_),
    .Y(_2749_));
 sg13g2_xnor2_1 _3669_ (.Y(_2750_),
    .A(_2739_),
    .B(_2748_));
 sg13g2_nor3_1 _3670_ (.A(_2718_),
    .B(_2738_),
    .C(_2750_),
    .Y(_2751_));
 sg13g2_o21ai_1 _3671_ (.B1(_2738_),
    .Y(_2752_),
    .A1(_2718_),
    .A2(_2750_));
 sg13g2_nor2b_1 _3672_ (.A(_2751_),
    .B_N(_2752_),
    .Y(_2753_));
 sg13g2_a21oi_1 _3673_ (.A1(_2749_),
    .A2(_2752_),
    .Y(_2754_),
    .B1(_2751_));
 sg13g2_xnor2_1 _3674_ (.Y(_2755_),
    .A(_2723_),
    .B(_2727_));
 sg13g2_nor2b_1 _3675_ (.A(_2754_),
    .B_N(_2755_),
    .Y(_2756_));
 sg13g2_xnor2_1 _3676_ (.Y(_2757_),
    .A(_2754_),
    .B(_2755_));
 sg13g2_a21oi_1 _3677_ (.A1(_2669_),
    .A2(_2757_),
    .Y(_2758_),
    .B1(_2756_));
 sg13g2_a21oi_1 _3678_ (.A1(_2730_),
    .A2(_2732_),
    .Y(_2759_),
    .B1(_2626_));
 sg13g2_nor3_1 _3679_ (.A(_2733_),
    .B(_2758_),
    .C(_2759_),
    .Y(_2760_));
 sg13g2_xnor2_1 _3680_ (.Y(_2761_),
    .A(_2717_),
    .B(_2748_));
 sg13g2_nor2b_1 _3681_ (.A(_2745_),
    .B_N(_2761_),
    .Y(_2762_));
 sg13g2_xor2_1 _3682_ (.B(_2753_),
    .A(_2749_),
    .X(_2763_));
 sg13g2_nand2_1 _3683_ (.Y(_2764_),
    .A(_2762_),
    .B(_2763_));
 sg13g2_xnor2_1 _3684_ (.Y(_2765_),
    .A(_2762_),
    .B(_2763_));
 sg13g2_o21ai_1 _3685_ (.B1(_2764_),
    .Y(_2766_),
    .A1(_2719_),
    .A2(_2765_));
 sg13g2_xnor2_1 _3686_ (.Y(_2767_),
    .A(_2670_),
    .B(_2757_));
 sg13g2_xnor2_1 _3687_ (.Y(_2768_),
    .A(_2766_),
    .B(_2767_));
 sg13g2_xnor2_1 _3688_ (.Y(_2769_),
    .A(_2745_),
    .B(_2761_));
 sg13g2_and2_1 _3689_ (.A(_2715_),
    .B(_2769_),
    .X(_2770_));
 sg13g2_xor2_1 _3690_ (.B(_2765_),
    .A(_2719_),
    .X(_2771_));
 sg13g2_and2_1 _3691_ (.A(_2770_),
    .B(_2771_),
    .X(_2772_));
 sg13g2_xnor2_1 _3692_ (.Y(_2773_),
    .A(_2715_),
    .B(_2769_));
 sg13g2_nand3_1 _3693_ (.B(_0032_),
    .C(_2296_),
    .A(net854),
    .Y(_2774_));
 sg13g2_nor3_1 _3694_ (.A(_2746_),
    .B(_2773_),
    .C(_2774_),
    .Y(_2775_));
 sg13g2_or2_1 _3695_ (.X(_2776_),
    .B(_2771_),
    .A(_2770_));
 sg13g2_o21ai_1 _3696_ (.B1(_2776_),
    .Y(_2777_),
    .A1(_2772_),
    .A2(_2775_));
 sg13g2_nand2b_1 _3697_ (.Y(_2778_),
    .B(net854),
    .A_N(_0032_));
 sg13g2_nor2_1 _3698_ (.A(_2291_),
    .B(_2778_),
    .Y(_2779_));
 sg13g2_a22oi_1 _3699_ (.Y(_2780_),
    .B1(_2779_),
    .B2(_2669_),
    .A2(_2767_),
    .A1(_2766_));
 sg13g2_o21ai_1 _3700_ (.B1(_2780_),
    .Y(_2781_),
    .A1(_2768_),
    .A2(_2777_));
 sg13g2_o21ai_1 _3701_ (.B1(_2758_),
    .Y(_2782_),
    .A1(_2733_),
    .A2(_2759_));
 sg13g2_nor2b_1 _3702_ (.A(_2760_),
    .B_N(_2782_),
    .Y(_2783_));
 sg13g2_a21oi_1 _3703_ (.A1(_2781_),
    .A2(_2782_),
    .Y(_2784_),
    .B1(_2760_));
 sg13g2_a221oi_1 _3704_ (.B2(_2782_),
    .C1(_2760_),
    .B1(_2781_),
    .A1(_2734_),
    .Y(_2785_),
    .A2(_2735_));
 sg13g2_nor2_1 _3705_ (.A(_2736_),
    .B(_2785_),
    .Y(_2786_));
 sg13g2_nand3b_1 _3706_ (.B(_2712_),
    .C(_2737_),
    .Y(_2787_),
    .A_N(_2785_));
 sg13g2_a22oi_1 _3707_ (.Y(_2788_),
    .B1(_2691_),
    .B2(_2710_),
    .A2(_2689_),
    .A1(_2687_));
 sg13g2_a22oi_1 _3708_ (.Y(_2789_),
    .B1(_2787_),
    .B2(_2788_),
    .A2(_2690_),
    .A1(_2688_));
 sg13g2_a221oi_1 _3709_ (.B2(_2788_),
    .C1(_2662_),
    .B1(_2787_),
    .A1(_2688_),
    .Y(_2790_),
    .A2(_2690_));
 sg13g2_nor2_1 _3710_ (.A(_2661_),
    .B(_2790_),
    .Y(_2791_));
 sg13g2_a21o_1 _3711_ (.A2(_2661_),
    .A1(_2623_),
    .B1(_2622_),
    .X(_2792_));
 sg13g2_a21oi_1 _3712_ (.A1(_2623_),
    .A2(_2790_),
    .Y(_2793_),
    .B1(_2792_));
 sg13g2_a21o_1 _3713_ (.A2(_2790_),
    .A1(_2623_),
    .B1(_2792_),
    .X(_2794_));
 sg13g2_a21oi_1 _3714_ (.A1(_2590_),
    .A2(_2616_),
    .Y(_2795_),
    .B1(_2615_));
 sg13g2_a21oi_1 _3715_ (.A1(_2592_),
    .A2(_2600_),
    .Y(_2796_),
    .B1(_2599_));
 sg13g2_a21oi_1 _3716_ (.A1(_2601_),
    .A2(_2613_),
    .Y(_2797_),
    .B1(_2612_));
 sg13g2_o21ai_1 _3717_ (.B1(_2596_),
    .Y(_2798_),
    .A1(_2220_),
    .A2(_2597_));
 sg13g2_nand2_1 _3718_ (.Y(_2799_),
    .A(_2607_),
    .B(_2609_));
 sg13g2_xor2_1 _3719_ (.B(_2300_),
    .A(net723),
    .X(_2800_));
 sg13g2_xnor2_1 _3720_ (.Y(_2801_),
    .A(_2799_),
    .B(_2800_));
 sg13g2_nor2b_1 _3721_ (.A(_2801_),
    .B_N(_2798_),
    .Y(_2802_));
 sg13g2_xor2_1 _3722_ (.B(_2801_),
    .A(_2798_),
    .X(_2803_));
 sg13g2_a21oi_1 _3723_ (.A1(_2605_),
    .A2(_2610_),
    .Y(_2804_),
    .B1(_2604_));
 sg13g2_xnor2_1 _3724_ (.Y(_2805_),
    .A(_2260_),
    .B(_2261_));
 sg13g2_xor2_1 _3725_ (.B(_2805_),
    .A(_2804_),
    .X(_2806_));
 sg13g2_nand2b_1 _3726_ (.Y(_2807_),
    .B(_2806_),
    .A_N(_2803_));
 sg13g2_xnor2_1 _3727_ (.Y(_2808_),
    .A(_2803_),
    .B(_2806_));
 sg13g2_nand2b_1 _3728_ (.Y(_2809_),
    .B(_2808_),
    .A_N(_2797_));
 sg13g2_xnor2_1 _3729_ (.Y(_2810_),
    .A(_2797_),
    .B(_2808_));
 sg13g2_nand2b_1 _3730_ (.Y(_2811_),
    .B(_2810_),
    .A_N(_2796_));
 sg13g2_xnor2_1 _3731_ (.Y(_2812_),
    .A(_2796_),
    .B(_2810_));
 sg13g2_nor2b_1 _3732_ (.A(_2795_),
    .B_N(_2812_),
    .Y(_2813_));
 sg13g2_o21ai_1 _3733_ (.B1(net798),
    .Y(_2814_),
    .A1(net869),
    .A2(_2214_));
 sg13g2_xnor2_1 _3734_ (.Y(_2815_),
    .A(_2795_),
    .B(_2812_));
 sg13g2_nor2b_1 _3735_ (.A(_2814_),
    .B_N(_2815_),
    .Y(_2816_));
 sg13g2_nand2_1 _3736_ (.Y(_2817_),
    .A(_2809_),
    .B(_2811_));
 sg13g2_a21o_1 _3737_ (.A2(_2800_),
    .A1(_2799_),
    .B1(_2802_),
    .X(_2818_));
 sg13g2_inv_1 _3738_ (.Y(_2819_),
    .A(_2818_));
 sg13g2_o21ai_1 _3739_ (.B1(_2807_),
    .Y(_2820_),
    .A1(_2804_),
    .A2(_2805_));
 sg13g2_xor2_1 _3740_ (.B(_2315_),
    .A(_2314_),
    .X(_2821_));
 sg13g2_nand2_1 _3741_ (.Y(_2822_),
    .A(_2820_),
    .B(_2821_));
 sg13g2_xnor2_1 _3742_ (.Y(_2823_),
    .A(_2820_),
    .B(_2821_));
 sg13g2_xnor2_1 _3743_ (.Y(_2824_),
    .A(_2819_),
    .B(_2823_));
 sg13g2_nand2b_1 _3744_ (.Y(_2825_),
    .B(_2817_),
    .A_N(_2824_));
 sg13g2_xor2_1 _3745_ (.B(_2824_),
    .A(_2817_),
    .X(_2826_));
 sg13g2_xor2_1 _3746_ (.B(_2826_),
    .A(_2408_),
    .X(_2827_));
 sg13g2_o21ai_1 _3747_ (.B1(_2827_),
    .Y(_2828_),
    .A1(_2813_),
    .A2(_2816_));
 sg13g2_xnor2_1 _3748_ (.Y(_2829_),
    .A(_2814_),
    .B(_2815_));
 sg13g2_o21ai_1 _3749_ (.B1(_2829_),
    .Y(_2830_),
    .A1(_2618_),
    .A2(_2620_));
 sg13g2_inv_1 _3750_ (.Y(_2831_),
    .A(_2830_));
 sg13g2_nand2_1 _3751_ (.Y(_2832_),
    .A(_2828_),
    .B(_2830_));
 sg13g2_nor3_1 _3752_ (.A(_2813_),
    .B(_2816_),
    .C(_2827_),
    .Y(_2833_));
 sg13g2_inv_1 _3753_ (.Y(_2834_),
    .A(_2833_));
 sg13g2_nor3_2 _3754_ (.A(_2618_),
    .B(_2620_),
    .C(_2829_),
    .Y(_2835_));
 sg13g2_o21ai_1 _3755_ (.B1(_2828_),
    .Y(_2836_),
    .A1(_2833_),
    .A2(_2835_));
 sg13g2_o21ai_1 _3756_ (.B1(_2836_),
    .Y(_2837_),
    .A1(_2794_),
    .A2(_2832_));
 sg13g2_o21ai_1 _3757_ (.B1(_2822_),
    .Y(_2838_),
    .A1(_2819_),
    .A2(_2823_));
 sg13g2_xnor2_1 _3758_ (.Y(_2839_),
    .A(_2356_),
    .B(_2357_));
 sg13g2_nand2b_1 _3759_ (.Y(_2840_),
    .B(_2838_),
    .A_N(_2839_));
 sg13g2_xnor2_1 _3760_ (.Y(_2841_),
    .A(_2838_),
    .B(_2839_));
 sg13g2_nand2b_1 _3761_ (.Y(_2842_),
    .B(_2841_),
    .A_N(_2408_));
 sg13g2_xnor2_1 _3762_ (.Y(_2843_),
    .A(_2408_),
    .B(_2841_));
 sg13g2_o21ai_1 _3763_ (.B1(_2825_),
    .Y(_2844_),
    .A1(_2408_),
    .A2(_2826_));
 sg13g2_nand2_1 _3764_ (.Y(_2845_),
    .A(_2843_),
    .B(_2844_));
 sg13g2_nor2_1 _3765_ (.A(_2843_),
    .B(_2844_),
    .Y(_2846_));
 sg13g2_xor2_1 _3766_ (.B(_2844_),
    .A(_2843_),
    .X(_2847_));
 sg13g2_xor2_1 _3767_ (.B(_2409_),
    .A(_2408_),
    .X(_2848_));
 sg13g2_nand3_1 _3768_ (.B(_2842_),
    .C(_2848_),
    .A(_2840_),
    .Y(_2849_));
 sg13g2_a21o_1 _3769_ (.A2(_2842_),
    .A1(_2840_),
    .B1(_2848_),
    .X(_2850_));
 sg13g2_and2_1 _3770_ (.A(_2849_),
    .B(_2850_),
    .X(_2851_));
 sg13g2_nand2_1 _3771_ (.Y(_2852_),
    .A(_2847_),
    .B(_2851_));
 sg13g2_nand2b_1 _3772_ (.Y(_2853_),
    .B(_2849_),
    .A_N(_2845_));
 sg13g2_and2_1 _3773_ (.A(_2850_),
    .B(_2853_),
    .X(_2854_));
 sg13g2_o21ai_1 _3774_ (.B1(_2854_),
    .Y(_2855_),
    .A1(_2837_),
    .A2(_2852_));
 sg13g2_a21oi_2 _3775_ (.B1(_2456_),
    .Y(_2856_),
    .A2(_2855_),
    .A1(_2457_));
 sg13g2_o21ai_1 _3776_ (.B1(_2449_),
    .Y(_2857_),
    .A1(_2412_),
    .A2(_2450_));
 sg13g2_a21oi_1 _3777_ (.A1(_2421_),
    .A2(_2447_),
    .Y(_2858_),
    .B1(_2446_));
 sg13g2_o21ai_1 _3778_ (.B1(_2417_),
    .Y(_2859_),
    .A1(_2418_),
    .A2(_2420_));
 sg13g2_a21oi_1 _3779_ (.A1(_2433_),
    .A2(_2444_),
    .Y(_2860_),
    .B1(_2443_));
 sg13g2_nor2_1 _3780_ (.A(_1373_),
    .B(_2563_),
    .Y(_2861_));
 sg13g2_o21ai_1 _3781_ (.B1(_2861_),
    .Y(_2862_),
    .A1(net830),
    .A2(net837));
 sg13g2_o21ai_1 _3782_ (.B1(_2438_),
    .Y(_2863_),
    .A1(_2426_),
    .A2(_2436_));
 sg13g2_xnor2_1 _3783_ (.Y(_2864_),
    .A(_2862_),
    .B(_2863_));
 sg13g2_a21oi_1 _3784_ (.A1(_2378_),
    .A2(_2429_),
    .Y(_2865_),
    .B1(_2427_));
 sg13g2_a21o_1 _3785_ (.A2(_2429_),
    .A1(_2427_),
    .B1(_2865_),
    .X(_2866_));
 sg13g2_nand2_2 _3786_ (.Y(_2867_),
    .A(net811),
    .B(net819));
 sg13g2_xnor2_1 _3787_ (.Y(_2868_),
    .A(_2427_),
    .B(_2867_));
 sg13g2_nor2_1 _3788_ (.A(_1373_),
    .B(net831),
    .Y(_2869_));
 sg13g2_xnor2_1 _3789_ (.Y(_2870_),
    .A(_2868_),
    .B(_2869_));
 sg13g2_nand3_1 _3790_ (.B(_2363_),
    .C(_2414_),
    .A(net723),
    .Y(_2871_));
 sg13g2_o21ai_1 _3791_ (.B1(_2871_),
    .Y(_2872_),
    .A1(_2363_),
    .A2(_2415_));
 sg13g2_xnor2_1 _3792_ (.Y(_2873_),
    .A(_2864_),
    .B(_2870_));
 sg13g2_xnor2_1 _3793_ (.Y(_2874_),
    .A(_2866_),
    .B(_2872_));
 sg13g2_xnor2_1 _3794_ (.Y(_2875_),
    .A(_2873_),
    .B(_2874_));
 sg13g2_a21oi_1 _3795_ (.A1(_1450_),
    .A2(_2441_),
    .Y(_2876_),
    .B1(_2440_));
 sg13g2_a21oi_1 _3796_ (.A1(_2423_),
    .A2(_2432_),
    .Y(_2877_),
    .B1(_2431_));
 sg13g2_xnor2_1 _3797_ (.Y(_2878_),
    .A(_2876_),
    .B(_2877_));
 sg13g2_xnor2_1 _3798_ (.Y(_2879_),
    .A(_2875_),
    .B(_2878_));
 sg13g2_xnor2_1 _3799_ (.Y(_2880_),
    .A(_2860_),
    .B(_2879_));
 sg13g2_xnor2_1 _3800_ (.Y(_2881_),
    .A(_2859_),
    .B(_2880_));
 sg13g2_xnor2_1 _3801_ (.Y(_2882_),
    .A(_2858_),
    .B(_2881_));
 sg13g2_xnor2_1 _3802_ (.Y(_2883_),
    .A(_2857_),
    .B(_2882_));
 sg13g2_mux2_1 _3803_ (.A0(_2453_),
    .A1(_2452_),
    .S(_2408_),
    .X(_2884_));
 sg13g2_xnor2_1 _3804_ (.Y(_2885_),
    .A(_2883_),
    .B(_2884_));
 sg13g2_xnor2_1 _3805_ (.Y(_2886_),
    .A(_2856_),
    .B(_2885_));
 sg13g2_nor2b_1 _3806_ (.A(_2886_),
    .B_N(\system_inst.neuron.u[13] ),
    .Y(_2887_));
 sg13g2_nor2b_1 _3807_ (.A(net742),
    .B_N(net681),
    .Y(_2888_));
 sg13g2_nand2b_1 _3808_ (.Y(_2889_),
    .B(net681),
    .A_N(net742));
 sg13g2_nor2_1 _3809_ (.A(net799),
    .B(_2888_),
    .Y(_2890_));
 sg13g2_nor2_1 _3810_ (.A(_2887_),
    .B(_2888_),
    .Y(_2891_));
 sg13g2_mux2_1 _3811_ (.A0(net681),
    .A1(_2891_),
    .S(_1373_),
    .X(_2892_));
 sg13g2_xnor2_1 _3812_ (.Y(_2893_),
    .A(_2175_),
    .B(_2212_));
 sg13g2_nand2_1 _3813_ (.Y(_2894_),
    .A(_2892_),
    .B(_2893_));
 sg13g2_and2_1 _3814_ (.A(_2213_),
    .B(_2894_),
    .X(_2895_));
 sg13g2_a21oi_1 _3815_ (.A1(_2196_),
    .A2(_2211_),
    .Y(_2896_),
    .B1(_2205_));
 sg13g2_inv_1 _3816_ (.Y(_2897_),
    .A(_2896_));
 sg13g2_xor2_1 _3817_ (.B(_2891_),
    .A(net9),
    .X(_2898_));
 sg13g2_xnor2_1 _3818_ (.Y(_2899_),
    .A(_2897_),
    .B(_2898_));
 sg13g2_nor2_1 _3819_ (.A(_2186_),
    .B(_2899_),
    .Y(_2900_));
 sg13g2_xor2_1 _3820_ (.B(_2899_),
    .A(_2186_),
    .X(_2901_));
 sg13g2_nor2b_1 _3821_ (.A(_2895_),
    .B_N(_2901_),
    .Y(_0108_));
 sg13g2_o21ai_1 _3822_ (.B1(_2889_),
    .Y(_0109_),
    .A1(net742),
    .A2(_1373_));
 sg13g2_xnor2_1 _3823_ (.Y(_0110_),
    .A(_2895_),
    .B(_2901_));
 sg13g2_a21oi_1 _3824_ (.A1(_0109_),
    .A2(_0110_),
    .Y(_0111_),
    .B1(_0108_));
 sg13g2_a21oi_1 _3825_ (.A1(_2897_),
    .A2(_2898_),
    .Y(_0112_),
    .B1(_2900_));
 sg13g2_o21ai_1 _3826_ (.B1(_2889_),
    .Y(_0113_),
    .A1(net9),
    .A2(_2887_));
 sg13g2_xnor2_1 _3827_ (.Y(_0114_),
    .A(net799),
    .B(_0113_));
 sg13g2_xor2_1 _3828_ (.B(_0114_),
    .A(_0112_),
    .X(_0115_));
 sg13g2_nand2b_1 _3829_ (.Y(_0116_),
    .B(_0115_),
    .A_N(_0111_));
 sg13g2_xnor2_1 _3830_ (.Y(_0117_),
    .A(_0111_),
    .B(_0115_));
 sg13g2_nand2_1 _3831_ (.Y(_0118_),
    .A(net815),
    .B(net6));
 sg13g2_xor2_1 _3832_ (.B(net7),
    .A(net811),
    .X(_0119_));
 sg13g2_nand2b_1 _3833_ (.Y(_0120_),
    .B(_0119_),
    .A_N(_0118_));
 sg13g2_nor2_1 _3834_ (.A(\system_inst.neuron.u[12] ),
    .B(_1384_),
    .Y(_0121_));
 sg13g2_xnor2_1 _3835_ (.Y(_0122_),
    .A(\system_inst.neuron.u[12] ),
    .B(net803));
 sg13g2_xnor2_1 _3836_ (.Y(_0123_),
    .A(_0118_),
    .B(_0119_));
 sg13g2_nand2_1 _3837_ (.Y(_0124_),
    .A(_0122_),
    .B(_0123_));
 sg13g2_and2_1 _3838_ (.A(_0120_),
    .B(_0124_),
    .X(_0125_));
 sg13g2_xor2_1 _3839_ (.B(_2155_),
    .A(_2145_),
    .X(_0126_));
 sg13g2_nand2b_1 _3840_ (.Y(_0127_),
    .B(_0126_),
    .A_N(_0125_));
 sg13g2_nand2_1 _3841_ (.Y(_0128_),
    .A(net681),
    .B(_0121_));
 sg13g2_xnor2_1 _3842_ (.Y(_0129_),
    .A(net681),
    .B(_0121_));
 sg13g2_xnor2_1 _3843_ (.Y(_0130_),
    .A(_0125_),
    .B(_0126_));
 sg13g2_nand2b_1 _3844_ (.Y(_0131_),
    .B(_0130_),
    .A_N(_0129_));
 sg13g2_and2_1 _3845_ (.A(_0127_),
    .B(_0131_),
    .X(_0132_));
 sg13g2_xnor2_1 _3846_ (.Y(_0133_),
    .A(_2892_),
    .B(_2893_));
 sg13g2_xor2_1 _3847_ (.B(_0133_),
    .A(_0132_),
    .X(_0134_));
 sg13g2_nand2b_1 _3848_ (.Y(_0135_),
    .B(_0134_),
    .A_N(_0128_));
 sg13g2_o21ai_1 _3849_ (.B1(_0135_),
    .Y(_0136_),
    .A1(_0132_),
    .A2(_0133_));
 sg13g2_xor2_1 _3850_ (.B(_0110_),
    .A(_0109_),
    .X(_0137_));
 sg13g2_nor2_1 _3851_ (.A(_0136_),
    .B(_0137_),
    .Y(_0138_));
 sg13g2_xor2_1 _3852_ (.B(_0134_),
    .A(_0128_),
    .X(_0139_));
 sg13g2_xor2_1 _3853_ (.B(net6),
    .A(net814),
    .X(_0140_));
 sg13g2_nand2_1 _3854_ (.Y(_0141_),
    .A(net5),
    .B(_0140_));
 sg13g2_nor2b_1 _3855_ (.A(\system_inst.neuron.u[11] ),
    .B_N(net806),
    .Y(_0142_));
 sg13g2_xor2_1 _3856_ (.B(net806),
    .A(\system_inst.neuron.u[11] ),
    .X(_0143_));
 sg13g2_xnor2_1 _3857_ (.Y(_0144_),
    .A(net5),
    .B(_0140_));
 sg13g2_o21ai_1 _3858_ (.B1(_0141_),
    .Y(_0145_),
    .A1(_0143_),
    .A2(_0144_));
 sg13g2_xor2_1 _3859_ (.B(_0123_),
    .A(_0122_),
    .X(_0146_));
 sg13g2_nand2_1 _3860_ (.Y(_0147_),
    .A(_0145_),
    .B(_0146_));
 sg13g2_o21ai_1 _3861_ (.B1(_2845_),
    .Y(_0148_),
    .A1(_2837_),
    .A2(_2846_));
 sg13g2_xor2_1 _3862_ (.B(_0148_),
    .A(_2851_),
    .X(_0149_));
 sg13g2_xnor2_1 _3863_ (.Y(_0150_),
    .A(_2458_),
    .B(_2855_));
 sg13g2_xor2_1 _3864_ (.B(_2855_),
    .A(_2458_),
    .X(_0151_));
 sg13g2_o21ai_1 _3865_ (.B1(net681),
    .Y(_0152_),
    .A1(_0149_),
    .A2(_0150_));
 sg13g2_inv_1 _3866_ (.Y(_0153_),
    .A(_0152_));
 sg13g2_xnor2_1 _3867_ (.Y(_0154_),
    .A(_2623_),
    .B(_2791_));
 sg13g2_nand2_1 _3868_ (.Y(_0155_),
    .A(_2828_),
    .B(_2834_));
 sg13g2_nor2_1 _3869_ (.A(_2831_),
    .B(_2835_),
    .Y(_0156_));
 sg13g2_o21ai_1 _3870_ (.B1(_2830_),
    .Y(_0157_),
    .A1(_2793_),
    .A2(_2835_));
 sg13g2_xor2_1 _3871_ (.B(_0157_),
    .A(_0155_),
    .X(_0158_));
 sg13g2_nand2b_1 _3872_ (.Y(_0159_),
    .B(_0154_),
    .A_N(_0158_));
 sg13g2_xnor2_1 _3873_ (.Y(_0160_),
    .A(_2837_),
    .B(_2847_));
 sg13g2_xnor2_1 _3874_ (.Y(_0161_),
    .A(_2793_),
    .B(_0156_));
 sg13g2_nand2_1 _3875_ (.Y(_0162_),
    .A(_0160_),
    .B(_0161_));
 sg13g2_inv_1 _3876_ (.Y(_0163_),
    .A(_0162_));
 sg13g2_xnor2_1 _3877_ (.Y(_0164_),
    .A(_0160_),
    .B(_0161_));
 sg13g2_nor2_1 _3878_ (.A(_0159_),
    .B(_0164_),
    .Y(_0165_));
 sg13g2_xor2_1 _3879_ (.B(_0164_),
    .A(_0159_),
    .X(_0166_));
 sg13g2_xnor2_1 _3880_ (.Y(_0167_),
    .A(_2662_),
    .B(_2789_));
 sg13g2_nand2_1 _3881_ (.Y(_0168_),
    .A(_0161_),
    .B(_0167_));
 sg13g2_inv_1 _3882_ (.Y(_0169_),
    .A(_0168_));
 sg13g2_xnor2_1 _3883_ (.Y(_0170_),
    .A(_0154_),
    .B(_0158_));
 sg13g2_or2_1 _3884_ (.X(_0171_),
    .B(_0170_),
    .A(_0169_));
 sg13g2_nand2_1 _3885_ (.Y(_0172_),
    .A(_0169_),
    .B(_0170_));
 sg13g2_xor2_1 _3886_ (.B(_2689_),
    .A(_2687_),
    .X(_0173_));
 sg13g2_a21oi_1 _3887_ (.A1(_2711_),
    .A2(_2787_),
    .Y(_0174_),
    .B1(_0173_));
 sg13g2_and3_1 _3888_ (.X(_0175_),
    .A(_2711_),
    .B(_2787_),
    .C(_0173_));
 sg13g2_nor2_1 _3889_ (.A(_0174_),
    .B(_0175_),
    .Y(_0176_));
 sg13g2_inv_1 _3890_ (.Y(_0177_),
    .A(_0176_));
 sg13g2_nand2_1 _3891_ (.Y(_0178_),
    .A(_0154_),
    .B(_0177_));
 sg13g2_xnor2_1 _3892_ (.Y(_0179_),
    .A(_0161_),
    .B(_0167_));
 sg13g2_or2_1 _3893_ (.X(_0180_),
    .B(_0179_),
    .A(_0178_));
 sg13g2_xor2_1 _3894_ (.B(_0179_),
    .A(_0178_),
    .X(_0181_));
 sg13g2_xnor2_1 _3895_ (.Y(_0182_),
    .A(_2712_),
    .B(_2786_));
 sg13g2_inv_1 _3896_ (.Y(_0183_),
    .A(_0182_));
 sg13g2_nand2_2 _3897_ (.Y(_0184_),
    .A(_0167_),
    .B(_0183_));
 sg13g2_inv_1 _3898_ (.Y(_0185_),
    .A(_0184_));
 sg13g2_xnor2_1 _3899_ (.Y(_0186_),
    .A(_0154_),
    .B(_0176_));
 sg13g2_xnor2_1 _3900_ (.Y(_0187_),
    .A(_0154_),
    .B(_0177_));
 sg13g2_nand2_1 _3901_ (.Y(_0188_),
    .A(_0184_),
    .B(_0187_));
 sg13g2_xor2_1 _3902_ (.B(_2735_),
    .A(_2734_),
    .X(_0189_));
 sg13g2_xnor2_1 _3903_ (.Y(_0190_),
    .A(_2784_),
    .B(_0189_));
 sg13g2_o21ai_1 _3904_ (.B1(_0190_),
    .Y(_0191_),
    .A1(_0174_),
    .A2(_0175_));
 sg13g2_xnor2_1 _3905_ (.Y(_0192_),
    .A(_0167_),
    .B(_0183_));
 sg13g2_nor2_1 _3906_ (.A(_0191_),
    .B(_0192_),
    .Y(_0193_));
 sg13g2_xor2_1 _3907_ (.B(_0192_),
    .A(_0191_),
    .X(_0194_));
 sg13g2_xnor2_1 _3908_ (.Y(_0195_),
    .A(_2781_),
    .B(_2783_));
 sg13g2_nor2_1 _3909_ (.A(_0182_),
    .B(_0195_),
    .Y(_0196_));
 sg13g2_or3_1 _3910_ (.A(_0174_),
    .B(_0175_),
    .C(_0190_),
    .X(_0197_));
 sg13g2_nand2_1 _3911_ (.Y(_0198_),
    .A(_0191_),
    .B(_0197_));
 sg13g2_nand3_1 _3912_ (.B(_0196_),
    .C(_0197_),
    .A(_0191_),
    .Y(_0199_));
 sg13g2_a21oi_1 _3913_ (.A1(_0191_),
    .A2(_0197_),
    .Y(_0200_),
    .B1(_0196_));
 sg13g2_xor2_1 _3914_ (.B(_0195_),
    .A(_0182_),
    .X(_0201_));
 sg13g2_nand2b_1 _3915_ (.Y(_0202_),
    .B(_2776_),
    .A_N(_2772_));
 sg13g2_nor2_1 _3916_ (.A(_2747_),
    .B(_2773_),
    .Y(_0203_));
 sg13g2_a21oi_1 _3917_ (.A1(_2776_),
    .A2(_0203_),
    .Y(_0204_),
    .B1(_2772_));
 sg13g2_xnor2_1 _3918_ (.Y(_0205_),
    .A(_2768_),
    .B(_0204_));
 sg13g2_inv_1 _3919_ (.Y(_0206_),
    .A(_0205_));
 sg13g2_nand2_1 _3920_ (.Y(_0207_),
    .A(_0190_),
    .B(_0206_));
 sg13g2_inv_1 _3921_ (.Y(_0208_),
    .A(_0207_));
 sg13g2_xnor2_1 _3922_ (.Y(_0209_),
    .A(_0190_),
    .B(_0205_));
 sg13g2_xor2_1 _3923_ (.B(_0203_),
    .A(_0202_),
    .X(_0210_));
 sg13g2_xnor2_1 _3924_ (.Y(_0211_),
    .A(_2747_),
    .B(_2773_));
 sg13g2_xnor2_1 _3925_ (.Y(_0212_),
    .A(_2743_),
    .B(_2746_));
 sg13g2_o21ai_1 _3926_ (.B1(_2778_),
    .Y(_0213_),
    .A1(net854),
    .A2(net861));
 sg13g2_nand2_1 _3927_ (.Y(_0214_),
    .A(_0195_),
    .B(_0210_));
 sg13g2_nor2_1 _3928_ (.A(_0205_),
    .B(_0211_),
    .Y(_0215_));
 sg13g2_nand2_1 _3929_ (.Y(_0216_),
    .A(_0205_),
    .B(_0211_));
 sg13g2_or3_1 _3930_ (.A(_1417_),
    .B(_0211_),
    .C(_0213_),
    .X(_0217_));
 sg13g2_xor2_1 _3931_ (.B(_2774_),
    .A(_2746_),
    .X(_0218_));
 sg13g2_nand2b_1 _3932_ (.Y(_0219_),
    .B(_0218_),
    .A_N(_0217_));
 sg13g2_a22oi_1 _3933_ (.Y(_0220_),
    .B1(_0219_),
    .B2(_0210_),
    .A2(_0217_),
    .A1(_0212_));
 sg13g2_o21ai_1 _3934_ (.B1(_0216_),
    .Y(_0221_),
    .A1(_0215_),
    .A2(_0220_));
 sg13g2_o21ai_1 _3935_ (.B1(_0221_),
    .Y(_0222_),
    .A1(_0195_),
    .A2(_0210_));
 sg13g2_nand2_1 _3936_ (.Y(_0223_),
    .A(_0214_),
    .B(_0222_));
 sg13g2_and3_1 _3937_ (.X(_0224_),
    .A(_0209_),
    .B(_0214_),
    .C(_0222_));
 sg13g2_nor2_1 _3938_ (.A(_0208_),
    .B(_0224_),
    .Y(_0225_));
 sg13g2_o21ai_1 _3939_ (.B1(_0201_),
    .Y(_0226_),
    .A1(_0208_),
    .A2(_0224_));
 sg13g2_xnor2_1 _3940_ (.Y(_0227_),
    .A(_0196_),
    .B(_0198_));
 sg13g2_a21oi_2 _3941_ (.B1(_0200_),
    .Y(_0228_),
    .A2(_0226_),
    .A1(_0199_));
 sg13g2_a21oi_1 _3942_ (.A1(_0194_),
    .A2(_0228_),
    .Y(_0229_),
    .B1(_0193_));
 sg13g2_a221oi_1 _3943_ (.B2(_0228_),
    .C1(_0193_),
    .B1(_0194_),
    .A1(_0185_),
    .Y(_0230_),
    .A2(_0186_));
 sg13g2_xnor2_1 _3944_ (.Y(_0231_),
    .A(_0184_),
    .B(_0186_));
 sg13g2_a21oi_1 _3945_ (.A1(_0184_),
    .A2(_0187_),
    .Y(_0232_),
    .B1(_0230_));
 sg13g2_nand3b_1 _3946_ (.B(_0181_),
    .C(_0188_),
    .Y(_0233_),
    .A_N(_0230_));
 sg13g2_nand2_1 _3947_ (.Y(_0234_),
    .A(_0180_),
    .B(_0233_));
 sg13g2_nand3_1 _3948_ (.B(_0180_),
    .C(_0233_),
    .A(_0172_),
    .Y(_0235_));
 sg13g2_and2_1 _3949_ (.A(_0171_),
    .B(_0172_),
    .X(_0236_));
 sg13g2_nand3_1 _3950_ (.B(_0171_),
    .C(_0235_),
    .A(_0166_),
    .Y(_0237_));
 sg13g2_nor2b_1 _3951_ (.A(_0158_),
    .B_N(_0149_),
    .Y(_0238_));
 sg13g2_xnor2_1 _3952_ (.Y(_0239_),
    .A(_0149_),
    .B(_0158_));
 sg13g2_a21oi_1 _3953_ (.A1(_0163_),
    .A2(_0239_),
    .Y(_0240_),
    .B1(_0165_));
 sg13g2_nor2_1 _3954_ (.A(_0163_),
    .B(_0239_),
    .Y(_0241_));
 sg13g2_a21o_1 _3955_ (.A2(_0240_),
    .A1(_0237_),
    .B1(_0241_),
    .X(_0242_));
 sg13g2_nand2_1 _3956_ (.Y(_0243_),
    .A(_0150_),
    .B(_0160_));
 sg13g2_nor2b_1 _3957_ (.A(_0149_),
    .B_N(net681),
    .Y(_0244_));
 sg13g2_xor2_1 _3958_ (.B(_0149_),
    .A(net681),
    .X(_0245_));
 sg13g2_nor2b_1 _3959_ (.A(_0243_),
    .B_N(_0245_),
    .Y(_0246_));
 sg13g2_nand2b_1 _3960_ (.Y(_0247_),
    .B(_0245_),
    .A_N(_0243_));
 sg13g2_xnor2_1 _3961_ (.Y(_0248_),
    .A(_0151_),
    .B(_0160_));
 sg13g2_and2_1 _3962_ (.A(_0238_),
    .B(_0248_),
    .X(_0249_));
 sg13g2_nand2b_1 _3963_ (.Y(_0250_),
    .B(_0243_),
    .A_N(_0245_));
 sg13g2_a21oi_1 _3964_ (.A1(_0249_),
    .A2(_0250_),
    .Y(_0251_),
    .B1(_0246_));
 sg13g2_o21ai_1 _3965_ (.B1(_0250_),
    .Y(_0252_),
    .A1(_0238_),
    .A2(_0248_));
 sg13g2_a22oi_1 _3966_ (.Y(_0253_),
    .B1(_0252_),
    .B2(_0247_),
    .A2(_0251_),
    .A1(_0242_));
 sg13g2_xnor2_1 _3967_ (.Y(_0254_),
    .A(_0151_),
    .B(_0244_));
 sg13g2_inv_1 _3968_ (.Y(_0255_),
    .A(_0254_));
 sg13g2_and2_1 _3969_ (.A(_0253_),
    .B(_0254_),
    .X(_0256_));
 sg13g2_nor2_1 _3970_ (.A(_0153_),
    .B(_0256_),
    .Y(_0257_));
 sg13g2_o21ai_1 _3971_ (.B1(_0142_),
    .Y(_0258_),
    .A1(_0153_),
    .A2(_0256_));
 sg13g2_xor2_1 _3972_ (.B(_0257_),
    .A(_0142_),
    .X(_0259_));
 sg13g2_xnor2_1 _3973_ (.Y(_0260_),
    .A(_0145_),
    .B(_0146_));
 sg13g2_o21ai_1 _3974_ (.B1(_0147_),
    .Y(_0261_),
    .A1(_0259_),
    .A2(_0260_));
 sg13g2_xnor2_1 _3975_ (.Y(_0262_),
    .A(_0129_),
    .B(_0130_));
 sg13g2_xnor2_1 _3976_ (.Y(_0263_),
    .A(_0261_),
    .B(_0262_));
 sg13g2_nor2_1 _3977_ (.A(_0258_),
    .B(_0263_),
    .Y(_0264_));
 sg13g2_a21oi_1 _3978_ (.A1(_0261_),
    .A2(_0262_),
    .Y(_0265_),
    .B1(_0264_));
 sg13g2_or2_1 _3979_ (.X(_0266_),
    .B(_0265_),
    .A(_0139_));
 sg13g2_nand2_1 _3980_ (.Y(_0267_),
    .A(_0136_),
    .B(_0137_));
 sg13g2_a21o_1 _3981_ (.A2(_0267_),
    .A1(_0266_),
    .B1(_0138_),
    .X(_0268_));
 sg13g2_nor2b_1 _3982_ (.A(_0138_),
    .B_N(_0267_),
    .Y(_0269_));
 sg13g2_xnor2_1 _3983_ (.Y(_0270_),
    .A(_0139_),
    .B(_0265_));
 sg13g2_inv_1 _3984_ (.Y(_0271_),
    .A(_0270_));
 sg13g2_nand2_1 _3985_ (.Y(_0272_),
    .A(_0269_),
    .B(_0271_));
 sg13g2_xor2_1 _3986_ (.B(net820),
    .A(net811),
    .X(_0273_));
 sg13g2_xnor2_1 _3987_ (.Y(_0274_),
    .A(net5),
    .B(net4));
 sg13g2_nand2_1 _3988_ (.Y(_0275_),
    .A(_0273_),
    .B(_0274_));
 sg13g2_o21ai_1 _3989_ (.B1(_0275_),
    .Y(_0276_),
    .A1(net5),
    .A2(_1439_));
 sg13g2_xor2_1 _3990_ (.B(_0144_),
    .A(_0143_),
    .X(_0277_));
 sg13g2_and2_1 _3991_ (.A(_0276_),
    .B(_0277_),
    .X(_0278_));
 sg13g2_xnor2_1 _3992_ (.Y(_0279_),
    .A(_0253_),
    .B(_0255_));
 sg13g2_nand2b_1 _3993_ (.Y(_0280_),
    .B(_0279_),
    .A_N(_2867_));
 sg13g2_inv_1 _3994_ (.Y(_0281_),
    .A(_0280_));
 sg13g2_xnor2_1 _3995_ (.Y(_0282_),
    .A(_2867_),
    .B(_0279_));
 sg13g2_xor2_1 _3996_ (.B(_0277_),
    .A(_0276_),
    .X(_0283_));
 sg13g2_a21oi_1 _3997_ (.A1(_0282_),
    .A2(_0283_),
    .Y(_0284_),
    .B1(_0278_));
 sg13g2_xnor2_1 _3998_ (.Y(_0285_),
    .A(_0259_),
    .B(_0260_));
 sg13g2_nor2_1 _3999_ (.A(_0284_),
    .B(_0285_),
    .Y(_0286_));
 sg13g2_xor2_1 _4000_ (.B(_0285_),
    .A(_0284_),
    .X(_0287_));
 sg13g2_a21oi_1 _4001_ (.A1(_0281_),
    .A2(_0287_),
    .Y(_0288_),
    .B1(_0286_));
 sg13g2_xor2_1 _4002_ (.B(_0263_),
    .A(_0258_),
    .X(_0289_));
 sg13g2_nor2b_1 _4003_ (.A(_0288_),
    .B_N(_0289_),
    .Y(_0290_));
 sg13g2_nand2b_1 _4004_ (.Y(_0291_),
    .B(_0288_),
    .A_N(_0289_));
 sg13g2_xnor2_1 _4005_ (.Y(_0292_),
    .A(_0280_),
    .B(_0287_));
 sg13g2_nand2_1 _4006_ (.Y(_0293_),
    .A(net831),
    .B(net3));
 sg13g2_nor2_1 _4007_ (.A(net4),
    .B(_0293_),
    .Y(_0294_));
 sg13g2_nor2b_1 _4008_ (.A(_1626_),
    .B_N(_2332_),
    .Y(_0295_));
 sg13g2_xnor2_1 _4009_ (.Y(_0296_),
    .A(_1439_),
    .B(_0293_));
 sg13g2_a21oi_1 _4010_ (.A1(_0295_),
    .A2(_0296_),
    .Y(_0297_),
    .B1(_0294_));
 sg13g2_xor2_1 _4011_ (.B(_0274_),
    .A(_0273_),
    .X(_0298_));
 sg13g2_inv_1 _4012_ (.Y(_0299_),
    .A(_0298_));
 sg13g2_xnor2_1 _4013_ (.Y(_0300_),
    .A(_0297_),
    .B(_0299_));
 sg13g2_inv_1 _4014_ (.Y(_0301_),
    .A(_0300_));
 sg13g2_nor2_1 _4015_ (.A(\system_inst.neuron.u[10] ),
    .B(_2332_),
    .Y(_0302_));
 sg13g2_xnor2_1 _4016_ (.Y(_0303_),
    .A(\system_inst.neuron.u[10] ),
    .B(_2332_));
 sg13g2_nand2_1 _4017_ (.Y(_0304_),
    .A(_0247_),
    .B(_0250_));
 sg13g2_xnor2_1 _4018_ (.Y(_0305_),
    .A(_0238_),
    .B(_0248_));
 sg13g2_nor2_1 _4019_ (.A(_0242_),
    .B(_0305_),
    .Y(_0306_));
 sg13g2_o21ai_1 _4020_ (.B1(_0304_),
    .Y(_0307_),
    .A1(_0249_),
    .A2(_0306_));
 sg13g2_or3_1 _4021_ (.A(_0249_),
    .B(_0304_),
    .C(_0306_),
    .X(_0308_));
 sg13g2_a21o_1 _4022_ (.A2(_0308_),
    .A1(_0307_),
    .B1(_0303_),
    .X(_0309_));
 sg13g2_nand3_1 _4023_ (.B(_0307_),
    .C(_0308_),
    .A(_0303_),
    .Y(_0310_));
 sg13g2_nand3_1 _4024_ (.B(_0309_),
    .C(_0310_),
    .A(_0301_),
    .Y(_0311_));
 sg13g2_o21ai_1 _4025_ (.B1(_0311_),
    .Y(_0312_),
    .A1(_0297_),
    .A2(_0299_));
 sg13g2_xnor2_1 _4026_ (.Y(_0313_),
    .A(_0282_),
    .B(_0283_));
 sg13g2_nor2b_1 _4027_ (.A(_0313_),
    .B_N(_0312_),
    .Y(_0314_));
 sg13g2_nor2b_1 _4028_ (.A(_0302_),
    .B_N(_0309_),
    .Y(_0315_));
 sg13g2_xor2_1 _4029_ (.B(_0313_),
    .A(_0312_),
    .X(_0316_));
 sg13g2_nor2_1 _4030_ (.A(_0315_),
    .B(_0316_),
    .Y(_0317_));
 sg13g2_o21ai_1 _4031_ (.B1(_0292_),
    .Y(_0318_),
    .A1(_0314_),
    .A2(_0317_));
 sg13g2_nand2b_1 _4032_ (.Y(_0319_),
    .B(_0318_),
    .A_N(_0290_));
 sg13g2_and2_1 _4033_ (.A(_0291_),
    .B(_0319_),
    .X(_0320_));
 sg13g2_nand2_1 _4034_ (.Y(_0321_),
    .A(net836),
    .B(net2));
 sg13g2_xor2_1 _4035_ (.B(net3),
    .A(net832),
    .X(_0322_));
 sg13g2_nor2b_1 _4036_ (.A(_0321_),
    .B_N(_0322_),
    .Y(_0323_));
 sg13g2_xnor2_1 _4037_ (.Y(_0324_),
    .A(_0321_),
    .B(_0322_));
 sg13g2_nand2b_1 _4038_ (.Y(_0325_),
    .B(net820),
    .A_N(\system_inst.neuron.u[8] ));
 sg13g2_xnor2_1 _4039_ (.Y(_0326_),
    .A(\system_inst.neuron.u[8] ),
    .B(net820));
 sg13g2_a21oi_1 _4040_ (.A1(_0324_),
    .A2(_0326_),
    .Y(_0327_),
    .B1(_0323_));
 sg13g2_xor2_1 _4041_ (.B(_0296_),
    .A(_0295_),
    .X(_0328_));
 sg13g2_nor2b_1 _4042_ (.A(_0327_),
    .B_N(_0328_),
    .Y(_0329_));
 sg13g2_xnor2_1 _4043_ (.Y(_0330_),
    .A(_0327_),
    .B(_0328_));
 sg13g2_xnor2_1 _4044_ (.Y(_0331_),
    .A(_0242_),
    .B(_0305_));
 sg13g2_xor2_1 _4045_ (.B(_0325_),
    .A(\system_inst.neuron.u[9] ),
    .X(_0332_));
 sg13g2_nand2b_1 _4046_ (.Y(_0333_),
    .B(_0332_),
    .A_N(_0331_));
 sg13g2_xnor2_1 _4047_ (.Y(_0334_),
    .A(_0331_),
    .B(_0332_));
 sg13g2_a21o_1 _4048_ (.A2(_0334_),
    .A1(_0330_),
    .B1(_0329_),
    .X(_0335_));
 sg13g2_a21o_1 _4049_ (.A2(_0310_),
    .A1(_0309_),
    .B1(_0301_),
    .X(_0336_));
 sg13g2_nand3_1 _4050_ (.B(_0335_),
    .C(_0336_),
    .A(_0311_),
    .Y(_0337_));
 sg13g2_o21ai_1 _4051_ (.B1(_0333_),
    .Y(_0338_),
    .A1(\system_inst.neuron.u[9] ),
    .A2(_0325_));
 sg13g2_a21o_1 _4052_ (.A2(_0336_),
    .A1(_0311_),
    .B1(_0335_),
    .X(_0339_));
 sg13g2_nand3_1 _4053_ (.B(_0338_),
    .C(_0339_),
    .A(_0337_),
    .Y(_0340_));
 sg13g2_and2_1 _4054_ (.A(_0337_),
    .B(_0340_),
    .X(_0341_));
 sg13g2_xnor2_1 _4055_ (.Y(_0342_),
    .A(_0315_),
    .B(_0316_));
 sg13g2_nand2_1 _4056_ (.Y(_0343_),
    .A(_0341_),
    .B(_0342_));
 sg13g2_a21o_1 _4057_ (.A2(_0339_),
    .A1(_0337_),
    .B1(_0338_),
    .X(_0344_));
 sg13g2_nand2_1 _4058_ (.Y(_0345_),
    .A(_0340_),
    .B(_0344_));
 sg13g2_nor2b_1 _4059_ (.A(\system_inst.neuron.u[7] ),
    .B_N(net824),
    .Y(_0346_));
 sg13g2_xor2_1 _4060_ (.B(net824),
    .A(\system_inst.neuron.u[7] ),
    .X(_0347_));
 sg13g2_xor2_1 _4061_ (.B(net2),
    .A(net836),
    .X(_0348_));
 sg13g2_nor2b_1 _4062_ (.A(_0347_),
    .B_N(_0348_),
    .Y(_0349_));
 sg13g2_inv_1 _4063_ (.Y(_0350_),
    .A(_0349_));
 sg13g2_xnor2_1 _4064_ (.Y(_0351_),
    .A(_0324_),
    .B(_0326_));
 sg13g2_nor2_1 _4065_ (.A(_0350_),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_xnor2_1 _4066_ (.Y(_0353_),
    .A(_0162_),
    .B(_0239_));
 sg13g2_nor2b_1 _4067_ (.A(_0165_),
    .B_N(_0237_),
    .Y(_0354_));
 sg13g2_xnor2_1 _4068_ (.Y(_0355_),
    .A(_0353_),
    .B(_0354_));
 sg13g2_nand2_1 _4069_ (.Y(_0356_),
    .A(_0346_),
    .B(_0355_));
 sg13g2_xor2_1 _4070_ (.B(_0355_),
    .A(_0346_),
    .X(_0357_));
 sg13g2_xnor2_1 _4071_ (.Y(_0358_),
    .A(_0349_),
    .B(_0351_));
 sg13g2_a21oi_1 _4072_ (.A1(_0357_),
    .A2(_0358_),
    .Y(_0359_),
    .B1(_0352_));
 sg13g2_xnor2_1 _4073_ (.Y(_0360_),
    .A(_0330_),
    .B(_0334_));
 sg13g2_or2_1 _4074_ (.X(_0361_),
    .B(_0360_),
    .A(_0359_));
 sg13g2_xnor2_1 _4075_ (.Y(_0362_),
    .A(_0359_),
    .B(_0360_));
 sg13g2_o21ai_1 _4076_ (.B1(_0361_),
    .Y(_0363_),
    .A1(_0356_),
    .A2(_0362_));
 sg13g2_inv_1 _4077_ (.Y(_0364_),
    .A(_0363_));
 sg13g2_nand3_1 _4078_ (.B(_0344_),
    .C(_0363_),
    .A(_0340_),
    .Y(_0365_));
 sg13g2_o21ai_1 _4079_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_0341_),
    .A2(_0342_));
 sg13g2_nor2b_1 _4080_ (.A(\system_inst.neuron.u[6] ),
    .B_N(net829),
    .Y(_0367_));
 sg13g2_xor2_1 _4081_ (.B(net829),
    .A(\system_inst.neuron.u[6] ),
    .X(_0368_));
 sg13g2_xnor2_1 _4082_ (.Y(_0369_),
    .A(_0234_),
    .B(_0236_));
 sg13g2_nor2_1 _4083_ (.A(_0368_),
    .B(_0369_),
    .Y(_0370_));
 sg13g2_xor2_1 _4084_ (.B(_0369_),
    .A(_0368_),
    .X(_0371_));
 sg13g2_nand2_1 _4085_ (.Y(_0372_),
    .A(net842),
    .B(_0371_));
 sg13g2_xnor2_1 _4086_ (.Y(_0373_),
    .A(_0347_),
    .B(_0348_));
 sg13g2_nand3_1 _4087_ (.B(_0371_),
    .C(_0373_),
    .A(net842),
    .Y(_0374_));
 sg13g2_nor2_1 _4088_ (.A(_0367_),
    .B(_0370_),
    .Y(_0375_));
 sg13g2_a21o_1 _4089_ (.A2(_0235_),
    .A1(_0171_),
    .B1(_0166_),
    .X(_0376_));
 sg13g2_and2_1 _4090_ (.A(_0237_),
    .B(_0376_),
    .X(_0377_));
 sg13g2_o21ai_1 _4091_ (.B1(_0377_),
    .Y(_0378_),
    .A1(_0367_),
    .A2(_0370_));
 sg13g2_xor2_1 _4092_ (.B(_0377_),
    .A(_0375_),
    .X(_0379_));
 sg13g2_a21oi_1 _4093_ (.A1(net845),
    .A2(_0371_),
    .Y(_0380_),
    .B1(_0373_));
 sg13g2_xnor2_1 _4094_ (.Y(_0381_),
    .A(_0372_),
    .B(_0373_));
 sg13g2_o21ai_1 _4095_ (.B1(_0374_),
    .Y(_0382_),
    .A1(_0379_),
    .A2(_0380_));
 sg13g2_xor2_1 _4096_ (.B(_0358_),
    .A(_0357_),
    .X(_0383_));
 sg13g2_nand2_1 _4097_ (.Y(_0384_),
    .A(_0382_),
    .B(_0383_));
 sg13g2_xnor2_1 _4098_ (.Y(_0385_),
    .A(_0382_),
    .B(_0383_));
 sg13g2_o21ai_1 _4099_ (.B1(_0384_),
    .Y(_0386_),
    .A1(_0378_),
    .A2(_0385_));
 sg13g2_xor2_1 _4100_ (.B(_0362_),
    .A(_0356_),
    .X(_0387_));
 sg13g2_nand2_1 _4101_ (.Y(_0388_),
    .A(_0386_),
    .B(_0387_));
 sg13g2_or2_1 _4102_ (.X(_0389_),
    .B(_0387_),
    .A(_0386_));
 sg13g2_xor2_1 _4103_ (.B(_0385_),
    .A(_0378_),
    .X(_0390_));
 sg13g2_xor2_1 _4104_ (.B(_0232_),
    .A(_0181_),
    .X(_0391_));
 sg13g2_nor2b_1 _4105_ (.A(\system_inst.neuron.u[5] ),
    .B_N(net836),
    .Y(_0392_));
 sg13g2_xnor2_1 _4106_ (.Y(_0393_),
    .A(\system_inst.neuron.u[5] ),
    .B(net836));
 sg13g2_xnor2_1 _4107_ (.Y(_0394_),
    .A(_0391_),
    .B(_0393_));
 sg13g2_or2_1 _4108_ (.X(_0395_),
    .B(_0394_),
    .A(_1395_));
 sg13g2_xnor2_1 _4109_ (.Y(_0396_),
    .A(net842),
    .B(_0371_));
 sg13g2_nor2_1 _4110_ (.A(_0395_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_a21oi_1 _4111_ (.A1(_0391_),
    .A2(_0393_),
    .Y(_0398_),
    .B1(_0392_));
 sg13g2_xnor2_1 _4112_ (.Y(_0399_),
    .A(_0395_),
    .B(_0396_));
 sg13g2_nor2_1 _4113_ (.A(_0398_),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_xnor2_1 _4114_ (.Y(_0401_),
    .A(_0379_),
    .B(_0381_));
 sg13g2_o21ai_1 _4115_ (.B1(_0401_),
    .Y(_0402_),
    .A1(_0397_),
    .A2(_0400_));
 sg13g2_xnor2_1 _4116_ (.Y(_0403_),
    .A(_1395_),
    .B(_0394_));
 sg13g2_nor2b_1 _4117_ (.A(\system_inst.neuron.u[4] ),
    .B_N(net842),
    .Y(_0404_));
 sg13g2_nand2b_1 _4118_ (.Y(_0405_),
    .B(\system_inst.neuron.u[4] ),
    .A_N(net842));
 sg13g2_nand2b_1 _4119_ (.Y(_0406_),
    .B(_0405_),
    .A_N(_0404_));
 sg13g2_xnor2_1 _4120_ (.Y(_0407_),
    .A(_0229_),
    .B(_0231_));
 sg13g2_xnor2_1 _4121_ (.Y(_0408_),
    .A(_0406_),
    .B(_0407_));
 sg13g2_nand2_1 _4122_ (.Y(_0409_),
    .A(net856),
    .B(_0408_));
 sg13g2_nor2_1 _4123_ (.A(_0403_),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_a21o_1 _4124_ (.A2(_0407_),
    .A1(_0405_),
    .B1(_0404_),
    .X(_0411_));
 sg13g2_xor2_1 _4125_ (.B(_0409_),
    .A(_0403_),
    .X(_0412_));
 sg13g2_a21oi_1 _4126_ (.A1(_0411_),
    .A2(_0412_),
    .Y(_0413_),
    .B1(_0410_));
 sg13g2_xnor2_1 _4127_ (.Y(_0414_),
    .A(_0398_),
    .B(_0399_));
 sg13g2_nor2_1 _4128_ (.A(_0413_),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_xnor2_1 _4129_ (.Y(_0416_),
    .A(_0411_),
    .B(_0412_));
 sg13g2_xor2_1 _4130_ (.B(net851),
    .A(\system_inst.neuron.u[3] ),
    .X(_0417_));
 sg13g2_xor2_1 _4131_ (.B(_0228_),
    .A(_0194_),
    .X(_0418_));
 sg13g2_nand2b_1 _4132_ (.Y(_0419_),
    .B(_0418_),
    .A_N(_0417_));
 sg13g2_xnor2_1 _4133_ (.Y(_0420_),
    .A(_0417_),
    .B(_0418_));
 sg13g2_nand2_1 _4134_ (.Y(_0421_),
    .A(net863),
    .B(_0420_));
 sg13g2_xnor2_1 _4135_ (.Y(_0422_),
    .A(net863),
    .B(_0420_));
 sg13g2_xnor2_1 _4136_ (.Y(_0423_),
    .A(\system_inst.neuron.u[2] ),
    .B(net858));
 sg13g2_xnor2_1 _4137_ (.Y(_0424_),
    .A(_0226_),
    .B(_0227_));
 sg13g2_nand2_1 _4138_ (.Y(_0425_),
    .A(_0423_),
    .B(_0424_));
 sg13g2_xnor2_1 _4139_ (.Y(_0426_),
    .A(_0423_),
    .B(_0424_));
 sg13g2_or2_1 _4140_ (.X(_0427_),
    .B(_0426_),
    .A(_1417_));
 sg13g2_nor2_1 _4141_ (.A(_0422_),
    .B(_0427_),
    .Y(_0428_));
 sg13g2_o21ai_1 _4142_ (.B1(_0425_),
    .Y(_0429_),
    .A1(\system_inst.neuron.u[2] ),
    .A2(_1406_));
 sg13g2_xor2_1 _4143_ (.B(_0427_),
    .A(_0422_),
    .X(_0430_));
 sg13g2_a21oi_1 _4144_ (.A1(_0429_),
    .A2(_0430_),
    .Y(_0431_),
    .B1(_0428_));
 sg13g2_nor2b_1 _4145_ (.A(\system_inst.neuron.u[1] ),
    .B_N(net862),
    .Y(_0432_));
 sg13g2_xnor2_1 _4146_ (.Y(_0433_),
    .A(_0201_),
    .B(_0225_));
 sg13g2_xnor2_1 _4147_ (.Y(_0434_),
    .A(\system_inst.neuron.u[1] ),
    .B(net862));
 sg13g2_a21oi_1 _4148_ (.A1(_0433_),
    .A2(_0434_),
    .Y(_0435_),
    .B1(_0432_));
 sg13g2_xnor2_1 _4149_ (.Y(_0436_),
    .A(_1417_),
    .B(_0426_));
 sg13g2_nor2_1 _4150_ (.A(_0435_),
    .B(_0436_),
    .Y(_0437_));
 sg13g2_xnor2_1 _4151_ (.Y(_0438_),
    .A(_0433_),
    .B(_0434_));
 sg13g2_xnor2_1 _4152_ (.Y(_0439_),
    .A(_0209_),
    .B(_0223_));
 sg13g2_nand3_1 _4153_ (.B(net868),
    .C(_0439_),
    .A(_1362_),
    .Y(_0440_));
 sg13g2_nor3_1 _4154_ (.A(_1362_),
    .B(net868),
    .C(_0439_),
    .Y(_0441_));
 sg13g2_a221oi_1 _4155_ (.B2(_0440_),
    .C1(_0441_),
    .B1(_0438_),
    .A1(_0435_),
    .Y(_0442_),
    .A2(_0436_));
 sg13g2_nor2_1 _4156_ (.A(_0437_),
    .B(_0442_),
    .Y(_0443_));
 sg13g2_xnor2_1 _4157_ (.Y(_0444_),
    .A(_0429_),
    .B(_0430_));
 sg13g2_nor2_1 _4158_ (.A(_0443_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_o21ai_1 _4159_ (.B1(_0431_),
    .Y(_0446_),
    .A1(_0443_),
    .A2(_0444_));
 sg13g2_o21ai_1 _4160_ (.B1(_0419_),
    .Y(_0447_),
    .A1(\system_inst.neuron.u[3] ),
    .A2(_1395_));
 sg13g2_xnor2_1 _4161_ (.Y(_0448_),
    .A(_0031_),
    .B(_0408_));
 sg13g2_nor2b_1 _4162_ (.A(_0421_),
    .B_N(_0448_),
    .Y(_0449_));
 sg13g2_xor2_1 _4163_ (.B(_0448_),
    .A(_0421_),
    .X(_0450_));
 sg13g2_nor2b_1 _4164_ (.A(_0450_),
    .B_N(_0447_),
    .Y(_0451_));
 sg13g2_xnor2_1 _4165_ (.Y(_0452_),
    .A(_0447_),
    .B(_0450_));
 sg13g2_a22oi_1 _4166_ (.Y(_0453_),
    .B1(_0446_),
    .B2(_0452_),
    .A2(_0445_),
    .A1(_0428_));
 sg13g2_nor2_1 _4167_ (.A(_0449_),
    .B(_0451_),
    .Y(_0454_));
 sg13g2_nor2_1 _4168_ (.A(_0416_),
    .B(_0453_),
    .Y(_0455_));
 sg13g2_a21oi_1 _4169_ (.A1(_0416_),
    .A2(_0453_),
    .Y(_0456_),
    .B1(_0454_));
 sg13g2_nor3_1 _4170_ (.A(_0415_),
    .B(_0455_),
    .C(_0456_),
    .Y(_0457_));
 sg13g2_nor3_1 _4171_ (.A(_0397_),
    .B(_0400_),
    .C(_0401_),
    .Y(_0458_));
 sg13g2_a21o_1 _4172_ (.A2(_0414_),
    .A1(_0413_),
    .B1(_0458_),
    .X(_0459_));
 sg13g2_o21ai_1 _4173_ (.B1(_0402_),
    .Y(_0460_),
    .A1(_0457_),
    .A2(_0459_));
 sg13g2_nand3_1 _4174_ (.B(_0390_),
    .C(_0460_),
    .A(_0389_),
    .Y(_0461_));
 sg13g2_a22oi_1 _4175_ (.Y(_0462_),
    .B1(_0388_),
    .B2(_0461_),
    .A2(_0364_),
    .A1(_0345_));
 sg13g2_o21ai_1 _4176_ (.B1(_0343_),
    .Y(_0463_),
    .A1(_0366_),
    .A2(_0462_));
 sg13g2_or3_1 _4177_ (.A(_0292_),
    .B(_0314_),
    .C(_0317_),
    .X(_0464_));
 sg13g2_nor2b_1 _4178_ (.A(_0290_),
    .B_N(_0291_),
    .Y(_0465_));
 sg13g2_and2_1 _4179_ (.A(_0318_),
    .B(_0464_),
    .X(_0466_));
 sg13g2_nand3b_1 _4180_ (.B(_0465_),
    .C(_0466_),
    .Y(_0467_),
    .A_N(_0463_));
 sg13g2_nor2b_2 _4181_ (.A(_0320_),
    .B_N(_0467_),
    .Y(_0468_));
 sg13g2_o21ai_1 _4182_ (.B1(_0268_),
    .Y(_0469_),
    .A1(_0272_),
    .A2(_0468_));
 sg13g2_o21ai_1 _4183_ (.B1(_0116_),
    .Y(_0470_),
    .A1(_0112_),
    .A2(_0114_));
 sg13g2_a21oi_1 _4184_ (.A1(_0117_),
    .A2(_0469_),
    .Y(_0471_),
    .B1(_0470_));
 sg13g2_xnor2_1 _4185_ (.Y(_0472_),
    .A(_0023_),
    .B(net9));
 sg13g2_o21ai_1 _4186_ (.B1(_2890_),
    .Y(_0473_),
    .A1(_2887_),
    .A2(_0472_));
 sg13g2_xnor2_1 _4187_ (.Y(_0474_),
    .A(_0471_),
    .B(_0473_));
 sg13g2_o21ai_1 _4188_ (.B1(_0266_),
    .Y(_0475_),
    .A1(_0270_),
    .A2(_0468_));
 sg13g2_xnor2_1 _4189_ (.Y(_0476_),
    .A(_0269_),
    .B(_0475_));
 sg13g2_xnor2_1 _4190_ (.Y(_0477_),
    .A(_0117_),
    .B(_0469_));
 sg13g2_xnor2_1 _4191_ (.Y(_0478_),
    .A(_0270_),
    .B(_0468_));
 sg13g2_nand2b_1 _4192_ (.Y(_0479_),
    .B(_0466_),
    .A_N(_0463_));
 sg13g2_nand2_1 _4193_ (.Y(_0480_),
    .A(_0318_),
    .B(_0479_));
 sg13g2_xnor2_1 _4194_ (.Y(_0481_),
    .A(_0465_),
    .B(_0480_));
 sg13g2_and4_1 _4195_ (.A(_0476_),
    .B(_0477_),
    .C(_0478_),
    .D(_0481_),
    .X(_0482_));
 sg13g2_nor2_1 _4196_ (.A(_0474_),
    .B(_0482_),
    .Y(_0483_));
 sg13g2_inv_1 _4197_ (.Y(_0484_),
    .A(net670));
 sg13g2_nand2_2 _4198_ (.Y(_0485_),
    .A(net727),
    .B(net669));
 sg13g2_xnor2_1 _4199_ (.Y(_0486_),
    .A(_1417_),
    .B(_0485_));
 sg13g2_nor2_1 _4200_ (.A(_2095_),
    .B(_0486_),
    .Y(_0036_));
 sg13g2_nand2_1 _4201_ (.Y(_0487_),
    .A(net182),
    .B(net669));
 sg13g2_and2_2 _4202_ (.A(net721),
    .B(net727),
    .X(_0488_));
 sg13g2_nand2_1 _4203_ (.Y(_0489_),
    .A(net722),
    .B(net727));
 sg13g2_xor2_1 _4204_ (.B(_0487_),
    .A(_0032_),
    .X(_0490_));
 sg13g2_a22oi_1 _4205_ (.Y(_0491_),
    .B1(_0488_),
    .B2(_0490_),
    .A2(net724),
    .A1(net864));
 sg13g2_nor2_1 _4206_ (.A(net873),
    .B(_0491_),
    .Y(_0037_));
 sg13g2_a21oi_1 _4207_ (.A1(_1428_),
    .A2(_0032_),
    .Y(_0492_),
    .B1(net863));
 sg13g2_nor2b_1 _4208_ (.A(_0485_),
    .B_N(_0492_),
    .Y(_0493_));
 sg13g2_xnor2_1 _4209_ (.Y(_0494_),
    .A(net857),
    .B(_0493_));
 sg13g2_nor2_1 _4210_ (.A(_2095_),
    .B(_0494_),
    .Y(_0038_));
 sg13g2_o21ai_1 _4211_ (.B1(_0031_),
    .Y(_0495_),
    .A1(net857),
    .A2(_0492_));
 sg13g2_nor2_1 _4212_ (.A(_0484_),
    .B(_0495_),
    .Y(_0496_));
 sg13g2_xnor2_1 _4213_ (.Y(_0497_),
    .A(net150),
    .B(_0496_));
 sg13g2_a22oi_1 _4214_ (.Y(_0498_),
    .B1(_0488_),
    .B2(_0497_),
    .A2(_2079_),
    .A1(net850));
 sg13g2_nor2_1 _4215_ (.A(net873),
    .B(_0498_),
    .Y(_0039_));
 sg13g2_a21oi_1 _4216_ (.A1(_0030_),
    .A2(_0495_),
    .Y(_0499_),
    .B1(net850));
 sg13g2_nor2b_1 _4217_ (.A(_0485_),
    .B_N(_0499_),
    .Y(_0500_));
 sg13g2_a21oi_1 _4218_ (.A1(net844),
    .A2(_0500_),
    .Y(_0501_),
    .B1(_2095_));
 sg13g2_o21ai_1 _4219_ (.B1(_0501_),
    .Y(_0502_),
    .A1(net844),
    .A2(_0500_));
 sg13g2_inv_1 _4220_ (.Y(_0040_),
    .A(_0502_));
 sg13g2_nand2_1 _4221_ (.Y(_0503_),
    .A(net838),
    .B(net724));
 sg13g2_o21ai_1 _4222_ (.B1(_0029_),
    .Y(_0504_),
    .A1(net844),
    .A2(_0499_));
 sg13g2_or2_1 _4223_ (.X(_0505_),
    .B(_0504_),
    .A(_0484_));
 sg13g2_a21oi_1 _4224_ (.A1(net165),
    .A2(_0505_),
    .Y(_0506_),
    .B1(_0489_));
 sg13g2_o21ai_1 _4225_ (.B1(_0506_),
    .Y(_0507_),
    .A1(net165),
    .A2(_0505_));
 sg13g2_a21oi_1 _4226_ (.A1(_0503_),
    .A2(_0507_),
    .Y(_0041_),
    .B1(net873));
 sg13g2_a21oi_1 _4227_ (.A1(net195),
    .A2(_0504_),
    .Y(_0508_),
    .B1(net838));
 sg13g2_nor2b_1 _4228_ (.A(_0485_),
    .B_N(_0508_),
    .Y(_0509_));
 sg13g2_o21ai_1 _4229_ (.B1(_2104_),
    .Y(_0510_),
    .A1(net831),
    .A2(_0509_));
 sg13g2_a21oi_1 _4230_ (.A1(net831),
    .A2(_0509_),
    .Y(_0042_),
    .B1(_0510_));
 sg13g2_o21ai_1 _4231_ (.B1(_0027_),
    .Y(_0511_),
    .A1(net830),
    .A2(_0508_));
 sg13g2_nor2_1 _4232_ (.A(_0484_),
    .B(_0511_),
    .Y(_0512_));
 sg13g2_a21oi_1 _4233_ (.A1(net825),
    .A2(_0512_),
    .Y(_0513_),
    .B1(net709));
 sg13g2_o21ai_1 _4234_ (.B1(_0513_),
    .Y(_0514_),
    .A1(net825),
    .A2(_0512_));
 sg13g2_a22oi_1 _4235_ (.Y(_0515_),
    .B1(_2087_),
    .B2(net112),
    .A2(net724),
    .A1(net825));
 sg13g2_a21oi_1 _4236_ (.A1(_0514_),
    .A2(_0515_),
    .Y(_0043_),
    .B1(net873));
 sg13g2_or2_1 _4237_ (.X(_0516_),
    .B(_0511_),
    .A(net825));
 sg13g2_nand2_1 _4238_ (.Y(_0517_),
    .A(net669),
    .B(_0516_));
 sg13g2_xnor2_1 _4239_ (.Y(_0518_),
    .A(net818),
    .B(net669));
 sg13g2_a21oi_1 _4240_ (.A1(_0517_),
    .A2(_0518_),
    .Y(_0519_),
    .B1(net709));
 sg13g2_o21ai_1 _4241_ (.B1(_0519_),
    .Y(_0520_),
    .A1(net818),
    .A2(_0517_));
 sg13g2_a22oi_1 _4242_ (.Y(_0521_),
    .B1(_2087_),
    .B2(net110),
    .A2(net724),
    .A1(net819));
 sg13g2_nand3_1 _4243_ (.B(_0520_),
    .C(_0521_),
    .A(net883),
    .Y(_0044_));
 sg13g2_xnor2_1 _4244_ (.Y(_0522_),
    .A(_0026_),
    .B(net669));
 sg13g2_o21ai_1 _4245_ (.B1(net669),
    .Y(_0523_),
    .A1(net819),
    .A2(_0516_));
 sg13g2_xnor2_1 _4246_ (.Y(_0524_),
    .A(_0522_),
    .B(_0523_));
 sg13g2_nand2_1 _4247_ (.Y(_0525_),
    .A(\system_inst.internal_param_c[2] ),
    .B(\system_inst.internal_param_c[1] ));
 sg13g2_xnor2_1 _4248_ (.Y(_0526_),
    .A(net131),
    .B(net130));
 sg13g2_o21ai_1 _4249_ (.B1(net883),
    .Y(_0527_),
    .A1(net815),
    .A2(net727));
 sg13g2_a221oi_1 _4250_ (.B2(_2087_),
    .C1(_0527_),
    .B1(_0526_),
    .A1(_0488_),
    .Y(_0045_),
    .A2(_0524_));
 sg13g2_nor2_1 _4251_ (.A(net819),
    .B(_0516_),
    .Y(_0528_));
 sg13g2_a21oi_2 _4252_ (.B1(_0026_),
    .Y(_0529_),
    .A2(_0528_),
    .A1(net669));
 sg13g2_xnor2_1 _4253_ (.Y(_0530_),
    .A(_0025_),
    .B(net670));
 sg13g2_inv_1 _4254_ (.Y(_0531_),
    .A(_0530_));
 sg13g2_a21oi_1 _4255_ (.A1(_0529_),
    .A2(_0531_),
    .Y(_0532_),
    .B1(net709));
 sg13g2_o21ai_1 _4256_ (.B1(_0532_),
    .Y(_0533_),
    .A1(_0529_),
    .A2(_0531_));
 sg13g2_nand2_1 _4257_ (.Y(_0534_),
    .A(net171),
    .B(_0525_));
 sg13g2_xnor2_1 _4258_ (.Y(_0535_),
    .A(net171),
    .B(_0525_));
 sg13g2_a22oi_1 _4259_ (.Y(_0536_),
    .B1(_2087_),
    .B2(net172),
    .A2(net724),
    .A1(net811));
 sg13g2_nand3_1 _4260_ (.B(_0533_),
    .C(_0536_),
    .A(net883),
    .Y(_0046_));
 sg13g2_a22oi_1 _4261_ (.Y(_0537_),
    .B1(_0529_),
    .B2(_0531_),
    .A2(_0484_),
    .A1(net812));
 sg13g2_xor2_1 _4262_ (.B(net670),
    .A(net808),
    .X(_0538_));
 sg13g2_xor2_1 _4263_ (.B(_0538_),
    .A(_0537_),
    .X(_0539_));
 sg13g2_nand2_1 _4264_ (.Y(_0540_),
    .A(net710),
    .B(_0539_));
 sg13g2_xnor2_1 _4265_ (.Y(_0541_),
    .A(net124),
    .B(_0534_));
 sg13g2_a22oi_1 _4266_ (.Y(_0542_),
    .B1(_2087_),
    .B2(_0541_),
    .A2(net724),
    .A1(net808));
 sg13g2_nand3_1 _4267_ (.B(_0540_),
    .C(_0542_),
    .A(net883),
    .Y(_0047_));
 sg13g2_nor2_1 _4268_ (.A(_0530_),
    .B(_0538_),
    .Y(_0543_));
 sg13g2_nor2_1 _4269_ (.A(_1648_),
    .B(net669),
    .Y(_0544_));
 sg13g2_a21o_1 _4270_ (.A2(_0543_),
    .A1(_0529_),
    .B1(_0544_),
    .X(_0545_));
 sg13g2_xor2_1 _4271_ (.B(net670),
    .A(_0024_),
    .X(_0546_));
 sg13g2_nand2_1 _4272_ (.Y(_0547_),
    .A(_0545_),
    .B(_0546_));
 sg13g2_a21oi_1 _4273_ (.A1(_0545_),
    .A2(_0546_),
    .Y(_0548_),
    .B1(net709));
 sg13g2_o21ai_1 _4274_ (.B1(_0548_),
    .Y(_0549_),
    .A1(_0545_),
    .A2(_0546_));
 sg13g2_nor2_1 _4275_ (.A(\system_inst.internal_param_c[4] ),
    .B(\system_inst.internal_param_c[3] ),
    .Y(_0550_));
 sg13g2_and2_1 _4276_ (.A(_0525_),
    .B(_0550_),
    .X(_0551_));
 sg13g2_nor2b_1 _4277_ (.A(net136),
    .B_N(_0551_),
    .Y(_0552_));
 sg13g2_inv_1 _4278_ (.Y(_0553_),
    .A(_0552_));
 sg13g2_xor2_1 _4279_ (.B(_0551_),
    .A(net136),
    .X(_0554_));
 sg13g2_a22oi_1 _4280_ (.Y(_0555_),
    .B1(_2087_),
    .B2(_0554_),
    .A2(net724),
    .A1(net803));
 sg13g2_nand3_1 _4281_ (.B(_0549_),
    .C(_0555_),
    .A(net883),
    .Y(_0048_));
 sg13g2_o21ai_1 _4282_ (.B1(_0547_),
    .Y(_0556_),
    .A1(_1384_),
    .A2(net670));
 sg13g2_xnor2_1 _4283_ (.Y(_0557_),
    .A(_0023_),
    .B(net670));
 sg13g2_xnor2_1 _4284_ (.Y(_0558_),
    .A(_0556_),
    .B(_0557_));
 sg13g2_nand2b_1 _4285_ (.Y(_0559_),
    .B(_0552_),
    .A_N(net126));
 sg13g2_a21oi_1 _4286_ (.A1(net126),
    .A2(_0553_),
    .Y(_0560_),
    .B1(net721));
 sg13g2_a221oi_1 _4287_ (.B2(_0560_),
    .C1(net724),
    .B1(_0559_),
    .A1(net721),
    .Y(_0561_),
    .A2(_0558_));
 sg13g2_o21ai_1 _4288_ (.B1(net883),
    .Y(_0562_),
    .A1(net799),
    .A2(net727));
 sg13g2_nor2_1 _4289_ (.A(_0561_),
    .B(_0562_),
    .Y(_0049_));
 sg13g2_nand3_1 _4290_ (.B(net760),
    .C(_2296_),
    .A(net758),
    .Y(_0563_));
 sg13g2_nand2_1 _4291_ (.Y(_0564_),
    .A(net754),
    .B(net866));
 sg13g2_and4_1 _4292_ (.A(net756),
    .B(net759),
    .C(net852),
    .D(net859),
    .X(_0565_));
 sg13g2_a22oi_1 _4293_ (.Y(_0566_),
    .B1(net859),
    .B2(net756),
    .A2(net852),
    .A1(net759));
 sg13g2_nor3_1 _4294_ (.A(_0564_),
    .B(_0565_),
    .C(_0566_),
    .Y(_0567_));
 sg13g2_o21ai_1 _4295_ (.B1(_0564_),
    .Y(_0568_),
    .A1(_0565_),
    .A2(_0566_));
 sg13g2_nor2b_1 _4296_ (.A(_0567_),
    .B_N(_0568_),
    .Y(_0569_));
 sg13g2_nand2b_1 _4297_ (.Y(_0570_),
    .B(_0569_),
    .A_N(_0563_));
 sg13g2_a22oi_1 _4298_ (.Y(_0571_),
    .B1(net852),
    .B2(net756),
    .A2(net846),
    .A1(net759));
 sg13g2_nand4_1 _4299_ (.B(net759),
    .C(net846),
    .A(net756),
    .Y(_0572_),
    .D(net852));
 sg13g2_nor2b_1 _4300_ (.A(_0571_),
    .B_N(_0572_),
    .Y(_0573_));
 sg13g2_and4_1 _4301_ (.A(net751),
    .B(net754),
    .C(net859),
    .D(net866),
    .X(_0574_));
 sg13g2_a22oi_1 _4302_ (.Y(_0575_),
    .B1(net866),
    .B2(net751),
    .A2(net859),
    .A1(net754));
 sg13g2_nor2_1 _4303_ (.A(_0574_),
    .B(_0575_),
    .Y(_0576_));
 sg13g2_nand2_1 _4304_ (.Y(_0577_),
    .A(_0573_),
    .B(_0576_));
 sg13g2_xnor2_1 _4305_ (.Y(_0578_),
    .A(_0573_),
    .B(_0576_));
 sg13g2_or2_1 _4306_ (.X(_0579_),
    .B(_0567_),
    .A(_0565_));
 sg13g2_nand2b_1 _4307_ (.Y(_0580_),
    .B(_0579_),
    .A_N(_0578_));
 sg13g2_xor2_1 _4308_ (.B(_0579_),
    .A(_0578_),
    .X(_0581_));
 sg13g2_xor2_1 _4309_ (.B(_0581_),
    .A(_0570_),
    .X(_0582_));
 sg13g2_and2_1 _4310_ (.A(net761),
    .B(_0582_),
    .X(_0583_));
 sg13g2_xnor2_1 _4311_ (.Y(_0584_),
    .A(_0563_),
    .B(_0569_));
 sg13g2_nand2_1 _4312_ (.Y(_0585_),
    .A(net764),
    .B(_0584_));
 sg13g2_nand2_1 _4313_ (.Y(_0586_),
    .A(net761),
    .B(_0584_));
 sg13g2_nand2_1 _4314_ (.Y(_0587_),
    .A(net764),
    .B(_0582_));
 sg13g2_or2_1 _4315_ (.X(_0588_),
    .B(_0587_),
    .A(_0586_));
 sg13g2_o21ai_1 _4316_ (.B1(_0580_),
    .Y(_0589_),
    .A1(_0570_),
    .A2(_0581_));
 sg13g2_nand2_1 _4317_ (.Y(_0590_),
    .A(net759),
    .B(net840));
 sg13g2_nand2_1 _4318_ (.Y(_0591_),
    .A(net756),
    .B(net846));
 sg13g2_nand3_1 _4319_ (.B(net846),
    .C(_0574_),
    .A(net756),
    .Y(_0592_));
 sg13g2_xnor2_1 _4320_ (.Y(_0593_),
    .A(_0574_),
    .B(_0591_));
 sg13g2_nand2b_1 _4321_ (.Y(_0594_),
    .B(_0593_),
    .A_N(_0590_));
 sg13g2_xnor2_1 _4322_ (.Y(_0595_),
    .A(_0590_),
    .B(_0593_));
 sg13g2_nand2_1 _4323_ (.Y(_0596_),
    .A(net754),
    .B(net853));
 sg13g2_and4_1 _4324_ (.A(net749),
    .B(net751),
    .C(net859),
    .D(net866),
    .X(_0597_));
 sg13g2_nand4_1 _4325_ (.B(net751),
    .C(net859),
    .A(net749),
    .Y(_0598_),
    .D(net866));
 sg13g2_a22oi_1 _4326_ (.Y(_0599_),
    .B1(net866),
    .B2(net749),
    .A2(net860),
    .A1(net751));
 sg13g2_nor3_1 _4327_ (.A(_0596_),
    .B(_0597_),
    .C(_0599_),
    .Y(_0600_));
 sg13g2_o21ai_1 _4328_ (.B1(_0596_),
    .Y(_0601_),
    .A1(_0597_),
    .A2(_0599_));
 sg13g2_nor2b_1 _4329_ (.A(_0600_),
    .B_N(_0601_),
    .Y(_0602_));
 sg13g2_nand2_1 _4330_ (.Y(_0603_),
    .A(_0595_),
    .B(_0602_));
 sg13g2_xnor2_1 _4331_ (.Y(_0604_),
    .A(_0595_),
    .B(_0602_));
 sg13g2_nor2_1 _4332_ (.A(_0577_),
    .B(_0604_),
    .Y(_0605_));
 sg13g2_xnor2_1 _4333_ (.Y(_0606_),
    .A(_0577_),
    .B(_0604_));
 sg13g2_nor2_1 _4334_ (.A(_0572_),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_xor2_1 _4335_ (.B(_0606_),
    .A(_0572_),
    .X(_0608_));
 sg13g2_nand2_1 _4336_ (.Y(_0609_),
    .A(_0589_),
    .B(_0608_));
 sg13g2_inv_1 _4337_ (.Y(_0610_),
    .A(_0609_));
 sg13g2_xor2_1 _4338_ (.B(_0608_),
    .A(_0589_),
    .X(_0611_));
 sg13g2_and2_1 _4339_ (.A(_1472_),
    .B(_0584_),
    .X(_0612_));
 sg13g2_xor2_1 _4340_ (.B(_0612_),
    .A(_0583_),
    .X(_0613_));
 sg13g2_and3_1 _4341_ (.X(_0614_),
    .A(net764),
    .B(net705),
    .C(_0613_));
 sg13g2_a21oi_1 _4342_ (.A1(net764),
    .A2(net705),
    .Y(_0615_),
    .B1(_0613_));
 sg13g2_nor2_1 _4343_ (.A(_0614_),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_nor3_1 _4344_ (.A(_0588_),
    .B(_0614_),
    .C(_0615_),
    .Y(_0617_));
 sg13g2_xnor2_1 _4345_ (.Y(_0618_),
    .A(_0588_),
    .B(_0616_));
 sg13g2_inv_1 _4346_ (.Y(_0619_),
    .A(_0618_));
 sg13g2_nor2_1 _4347_ (.A(_0605_),
    .B(_0607_),
    .Y(_0620_));
 sg13g2_and2_1 _4348_ (.A(_0592_),
    .B(_0594_),
    .X(_0621_));
 sg13g2_inv_1 _4349_ (.Y(_0622_),
    .A(_0621_));
 sg13g2_nand2_1 _4350_ (.Y(_0623_),
    .A(net747),
    .B(net866));
 sg13g2_nand2_1 _4351_ (.Y(_0624_),
    .A(net754),
    .B(net846));
 sg13g2_nand2_1 _4352_ (.Y(_0625_),
    .A(net749),
    .B(net852));
 sg13g2_and4_1 _4353_ (.A(net749),
    .B(net751),
    .C(net852),
    .D(net859),
    .X(_0626_));
 sg13g2_a22oi_1 _4354_ (.Y(_0627_),
    .B1(net859),
    .B2(net749),
    .A2(net852),
    .A1(net751));
 sg13g2_nor2_1 _4355_ (.A(_0626_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_nor3_1 _4356_ (.A(_0624_),
    .B(_0626_),
    .C(_0627_),
    .Y(_0629_));
 sg13g2_xnor2_1 _4357_ (.Y(_0630_),
    .A(_0624_),
    .B(_0628_));
 sg13g2_nand2b_1 _4358_ (.Y(_0631_),
    .B(_0630_),
    .A_N(_0623_));
 sg13g2_xnor2_1 _4359_ (.Y(_0632_),
    .A(_0623_),
    .B(_0630_));
 sg13g2_nand2_1 _4360_ (.Y(_0633_),
    .A(net759),
    .B(net835));
 sg13g2_o21ai_1 _4361_ (.B1(_0598_),
    .Y(_0634_),
    .A1(_0596_),
    .A2(_0599_));
 sg13g2_nand2_1 _4362_ (.Y(_0635_),
    .A(net756),
    .B(net840));
 sg13g2_nand2b_1 _4363_ (.Y(_0636_),
    .B(_0634_),
    .A_N(_0635_));
 sg13g2_xnor2_1 _4364_ (.Y(_0637_),
    .A(_0634_),
    .B(_0635_));
 sg13g2_nand2b_1 _4365_ (.Y(_0638_),
    .B(_0637_),
    .A_N(_0633_));
 sg13g2_xnor2_1 _4366_ (.Y(_0639_),
    .A(_0633_),
    .B(_0637_));
 sg13g2_nand2_1 _4367_ (.Y(_0640_),
    .A(_0632_),
    .B(_0639_));
 sg13g2_xnor2_1 _4368_ (.Y(_0641_),
    .A(_0632_),
    .B(_0639_));
 sg13g2_nor2_1 _4369_ (.A(_0603_),
    .B(_0641_),
    .Y(_0642_));
 sg13g2_xor2_1 _4370_ (.B(_0641_),
    .A(_0603_),
    .X(_0643_));
 sg13g2_xnor2_1 _4371_ (.Y(_0644_),
    .A(_0621_),
    .B(_0643_));
 sg13g2_nor2b_1 _4372_ (.A(_0620_),
    .B_N(_0644_),
    .Y(_0645_));
 sg13g2_xnor2_1 _4373_ (.Y(_0646_),
    .A(_0620_),
    .B(_0644_));
 sg13g2_a21o_1 _4374_ (.A2(_0646_),
    .A1(_0610_),
    .B1(_0645_),
    .X(_0647_));
 sg13g2_a21oi_2 _4375_ (.B1(_0642_),
    .Y(_0648_),
    .A2(_0643_),
    .A1(_0622_));
 sg13g2_nand2_2 _4376_ (.Y(_0649_),
    .A(_0636_),
    .B(_0638_));
 sg13g2_nand2_2 _4377_ (.Y(_0650_),
    .A(net745),
    .B(net860));
 sg13g2_nor2_1 _4378_ (.A(_0623_),
    .B(_0650_),
    .Y(_0651_));
 sg13g2_a22oi_1 _4379_ (.Y(_0652_),
    .B1(net866),
    .B2(net745),
    .A2(net860),
    .A1(net747));
 sg13g2_nor2_1 _4380_ (.A(_0651_),
    .B(_0652_),
    .Y(_0653_));
 sg13g2_nand2_1 _4381_ (.Y(_0654_),
    .A(net754),
    .B(net840));
 sg13g2_nand2_1 _4382_ (.Y(_0655_),
    .A(net752),
    .B(net846));
 sg13g2_or2_1 _4383_ (.X(_0656_),
    .B(_0655_),
    .A(_0625_));
 sg13g2_xor2_1 _4384_ (.B(_0655_),
    .A(_0625_),
    .X(_0657_));
 sg13g2_nand2b_1 _4385_ (.Y(_0658_),
    .B(_0657_),
    .A_N(_0654_));
 sg13g2_xnor2_1 _4386_ (.Y(_0659_),
    .A(_0654_),
    .B(_0657_));
 sg13g2_nand2_1 _4387_ (.Y(_0660_),
    .A(_0653_),
    .B(_0659_));
 sg13g2_xnor2_1 _4388_ (.Y(_0661_),
    .A(_0653_),
    .B(_0659_));
 sg13g2_nor2_1 _4389_ (.A(_0631_),
    .B(_0661_),
    .Y(_0662_));
 sg13g2_xor2_1 _4390_ (.B(_0661_),
    .A(_0631_),
    .X(_0663_));
 sg13g2_nand2_1 _4391_ (.Y(_0664_),
    .A(net759),
    .B(net827));
 sg13g2_or2_1 _4392_ (.X(_0665_),
    .B(_0629_),
    .A(_0626_));
 sg13g2_nand2_1 _4393_ (.Y(_0666_),
    .A(net756),
    .B(net835));
 sg13g2_nand2b_1 _4394_ (.Y(_0667_),
    .B(_0665_),
    .A_N(_0666_));
 sg13g2_xnor2_1 _4395_ (.Y(_0668_),
    .A(_0665_),
    .B(_0666_));
 sg13g2_nand2b_1 _4396_ (.Y(_0669_),
    .B(_0668_),
    .A_N(_0664_));
 sg13g2_xnor2_1 _4397_ (.Y(_0670_),
    .A(_0664_),
    .B(_0668_));
 sg13g2_xnor2_1 _4398_ (.Y(_0671_),
    .A(_0663_),
    .B(_0670_));
 sg13g2_nor2_1 _4399_ (.A(_0640_),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_xor2_1 _4400_ (.B(_0671_),
    .A(_0640_),
    .X(_0673_));
 sg13g2_xnor2_1 _4401_ (.Y(_0674_),
    .A(_0649_),
    .B(_0673_));
 sg13g2_nor2_1 _4402_ (.A(_0648_),
    .B(_0674_),
    .Y(_0675_));
 sg13g2_xor2_1 _4403_ (.B(_0674_),
    .A(_0648_),
    .X(_0676_));
 sg13g2_xnor2_1 _4404_ (.Y(_0677_),
    .A(_0647_),
    .B(_0676_));
 sg13g2_nor2_1 _4405_ (.A(\system_inst.neuron.u[1] ),
    .B(_0677_),
    .Y(_0678_));
 sg13g2_xnor2_1 _4406_ (.Y(_0679_),
    .A(_0609_),
    .B(_0646_));
 sg13g2_nand2b_2 _4407_ (.Y(_0680_),
    .B(\system_inst.neuron.u[0] ),
    .A_N(_0679_));
 sg13g2_xnor2_1 _4408_ (.Y(_0681_),
    .A(_1351_),
    .B(_0677_));
 sg13g2_a21oi_2 _4409_ (.B1(_0678_),
    .Y(_0682_),
    .A2(_0681_),
    .A1(_0680_));
 sg13g2_a21oi_1 _4410_ (.A1(_0647_),
    .A2(_0676_),
    .Y(_0683_),
    .B1(_0675_));
 sg13g2_a21oi_2 _4411_ (.B1(_0672_),
    .Y(_0684_),
    .A2(_0673_),
    .A1(_0649_));
 sg13g2_nand2_1 _4412_ (.Y(_0685_),
    .A(_0667_),
    .B(_0669_));
 sg13g2_a21oi_1 _4413_ (.A1(_0663_),
    .A2(_0670_),
    .Y(_0686_),
    .B1(_0662_));
 sg13g2_nand2_1 _4414_ (.Y(_0687_),
    .A(net747),
    .B(net852));
 sg13g2_nand2_1 _4415_ (.Y(_0688_),
    .A(net744),
    .B(net865));
 sg13g2_nand2_1 _4416_ (.Y(_0689_),
    .A(net744),
    .B(net868));
 sg13g2_xor2_1 _4417_ (.B(_0689_),
    .A(_0650_),
    .X(_0690_));
 sg13g2_nand2b_1 _4418_ (.Y(_0691_),
    .B(_0690_),
    .A_N(_0687_));
 sg13g2_xnor2_1 _4419_ (.Y(_0692_),
    .A(_0687_),
    .B(_0690_));
 sg13g2_and2_1 _4420_ (.A(_0651_),
    .B(_0692_),
    .X(_0693_));
 sg13g2_xor2_1 _4421_ (.B(_0692_),
    .A(_0651_),
    .X(_0694_));
 sg13g2_nand2_1 _4422_ (.Y(_0695_),
    .A(net754),
    .B(net835));
 sg13g2_nand2_2 _4423_ (.Y(_0696_),
    .A(net749),
    .B(net840));
 sg13g2_nor2_1 _4424_ (.A(_0655_),
    .B(_0696_),
    .Y(_0697_));
 sg13g2_or2_1 _4425_ (.X(_0698_),
    .B(_0696_),
    .A(_0655_));
 sg13g2_a22oi_1 _4426_ (.Y(_0699_),
    .B1(net846),
    .B2(net749),
    .A2(net840),
    .A1(net751));
 sg13g2_nor2_1 _4427_ (.A(_0697_),
    .B(_0699_),
    .Y(_0700_));
 sg13g2_xnor2_1 _4428_ (.Y(_0701_),
    .A(_0695_),
    .B(_0700_));
 sg13g2_xnor2_1 _4429_ (.Y(_0702_),
    .A(_0694_),
    .B(_0701_));
 sg13g2_nor2_1 _4430_ (.A(_0660_),
    .B(_0702_),
    .Y(_0703_));
 sg13g2_xor2_1 _4431_ (.B(_0702_),
    .A(_0660_),
    .X(_0704_));
 sg13g2_nand2_1 _4432_ (.Y(_0705_),
    .A(net759),
    .B(net822));
 sg13g2_and2_1 _4433_ (.A(_0656_),
    .B(_0658_),
    .X(_0706_));
 sg13g2_nand2_1 _4434_ (.Y(_0707_),
    .A(net757),
    .B(net827));
 sg13g2_xor2_1 _4435_ (.B(_0707_),
    .A(_0706_),
    .X(_0708_));
 sg13g2_nand2b_1 _4436_ (.Y(_0709_),
    .B(_0708_),
    .A_N(_0705_));
 sg13g2_xnor2_1 _4437_ (.Y(_0710_),
    .A(_0705_),
    .B(_0708_));
 sg13g2_xnor2_1 _4438_ (.Y(_0711_),
    .A(_0704_),
    .B(_0710_));
 sg13g2_nor2_1 _4439_ (.A(_0686_),
    .B(_0711_),
    .Y(_0712_));
 sg13g2_xor2_1 _4440_ (.B(_0711_),
    .A(_0686_),
    .X(_0713_));
 sg13g2_xnor2_1 _4441_ (.Y(_0714_),
    .A(_0685_),
    .B(_0713_));
 sg13g2_or2_1 _4442_ (.X(_0715_),
    .B(_0714_),
    .A(_0684_));
 sg13g2_and2_1 _4443_ (.A(_0684_),
    .B(_0714_),
    .X(_0716_));
 sg13g2_xor2_1 _4444_ (.B(_0714_),
    .A(_0684_),
    .X(_0717_));
 sg13g2_xnor2_1 _4445_ (.Y(_0718_),
    .A(_0683_),
    .B(_0717_));
 sg13g2_xnor2_1 _4446_ (.Y(_0719_),
    .A(_0022_),
    .B(_0718_));
 sg13g2_xor2_1 _4447_ (.B(_0719_),
    .A(_0682_),
    .X(_0720_));
 sg13g2_xnor2_1 _4448_ (.Y(_0721_),
    .A(_0682_),
    .B(_0719_));
 sg13g2_xor2_1 _4449_ (.B(_0681_),
    .A(_0680_),
    .X(_0722_));
 sg13g2_xnor2_1 _4450_ (.Y(_0723_),
    .A(_0680_),
    .B(_0681_));
 sg13g2_nor2_1 _4451_ (.A(net740),
    .B(_0723_),
    .Y(_0724_));
 sg13g2_nand2_1 _4452_ (.Y(_0725_),
    .A(net767),
    .B(net702));
 sg13g2_xnor2_1 _4453_ (.Y(_0726_),
    .A(_1362_),
    .B(_0679_));
 sg13g2_nand2_1 _4454_ (.Y(_0727_),
    .A(net770),
    .B(net703));
 sg13g2_nor2_1 _4455_ (.A(net734),
    .B(_0723_),
    .Y(_0728_));
 sg13g2_and2_1 _4456_ (.A(net767),
    .B(net703),
    .X(_0729_));
 sg13g2_nand2_1 _4457_ (.Y(_0730_),
    .A(net767),
    .B(net703));
 sg13g2_nand3_1 _4458_ (.B(net701),
    .C(_0729_),
    .A(net770),
    .Y(_0731_));
 sg13g2_o21ai_1 _4459_ (.B1(_0730_),
    .Y(_0732_),
    .A1(net734),
    .A2(_0723_));
 sg13g2_o21ai_1 _4460_ (.B1(_0729_),
    .Y(_0733_),
    .A1(net734),
    .A2(_0723_));
 sg13g2_nand3_1 _4461_ (.B(net701),
    .C(_0730_),
    .A(net770),
    .Y(_0734_));
 sg13g2_and4_1 _4462_ (.A(net776),
    .B(net699),
    .C(_0731_),
    .D(_0732_),
    .X(_0735_));
 sg13g2_nand4_1 _4463_ (.B(net699),
    .C(_0731_),
    .A(net776),
    .Y(_0736_),
    .D(_0732_));
 sg13g2_a22oi_1 _4464_ (.Y(_0737_),
    .B1(_0731_),
    .B2(_0732_),
    .A2(net699),
    .A1(net776));
 sg13g2_a22oi_1 _4465_ (.Y(_0738_),
    .B1(_0733_),
    .B2(_0734_),
    .A2(net699),
    .A1(net776));
 sg13g2_and4_1 _4466_ (.A(net776),
    .B(net699),
    .C(_0733_),
    .D(_0734_),
    .X(_0739_));
 sg13g2_nor3_2 _4467_ (.A(_0619_),
    .B(_0735_),
    .C(_0737_),
    .Y(_0740_));
 sg13g2_o21ai_1 _4468_ (.B1(_0618_),
    .Y(_0741_),
    .A1(_0738_),
    .A2(_0739_));
 sg13g2_nor2_1 _4469_ (.A(_0617_),
    .B(_0740_),
    .Y(_0742_));
 sg13g2_nand2b_1 _4470_ (.Y(_0743_),
    .B(_0741_),
    .A_N(_0617_));
 sg13g2_nand2b_1 _4471_ (.Y(_0744_),
    .B(_0718_),
    .A_N(\system_inst.neuron.u[2] ));
 sg13g2_o21ai_1 _4472_ (.B1(_0744_),
    .Y(_0745_),
    .A1(_0682_),
    .A2(_0719_));
 sg13g2_o21ai_1 _4473_ (.B1(_0715_),
    .Y(_0746_),
    .A1(_0683_),
    .A2(_0716_));
 sg13g2_a21oi_1 _4474_ (.A1(_0685_),
    .A2(_0713_),
    .Y(_0747_),
    .B1(_0712_));
 sg13g2_o21ai_1 _4475_ (.B1(_0709_),
    .Y(_0748_),
    .A1(_0706_),
    .A2(_0707_));
 sg13g2_a21oi_1 _4476_ (.A1(_0704_),
    .A2(_0710_),
    .Y(_0749_),
    .B1(_0703_));
 sg13g2_a21o_1 _4477_ (.A2(_0701_),
    .A1(_0694_),
    .B1(_0693_),
    .X(_0750_));
 sg13g2_o21ai_1 _4478_ (.B1(_0691_),
    .Y(_0751_),
    .A1(_0650_),
    .A2(_0689_));
 sg13g2_nand2_1 _4479_ (.Y(_0752_),
    .A(net747),
    .B(net847));
 sg13g2_nand2_2 _4480_ (.Y(_0753_),
    .A(net744),
    .B(net853));
 sg13g2_nand2_1 _4481_ (.Y(_0754_),
    .A(net745),
    .B(net853));
 sg13g2_xor2_1 _4482_ (.B(_0754_),
    .A(_0688_),
    .X(_0755_));
 sg13g2_nand2b_1 _4483_ (.Y(_0756_),
    .B(_0755_),
    .A_N(_0752_));
 sg13g2_xnor2_1 _4484_ (.Y(_0757_),
    .A(_0752_),
    .B(_0755_));
 sg13g2_xnor2_1 _4485_ (.Y(_0758_),
    .A(_0751_),
    .B(_0757_));
 sg13g2_nand2_1 _4486_ (.Y(_0759_),
    .A(net754),
    .B(net827));
 sg13g2_nand2_1 _4487_ (.Y(_0760_),
    .A(net750),
    .B(net835));
 sg13g2_nand2_1 _4488_ (.Y(_0761_),
    .A(net752),
    .B(net835));
 sg13g2_xor2_1 _4489_ (.B(_0761_),
    .A(_0696_),
    .X(_0762_));
 sg13g2_nand2b_1 _4490_ (.Y(_0763_),
    .B(_0762_),
    .A_N(_0759_));
 sg13g2_xnor2_1 _4491_ (.Y(_0764_),
    .A(_0759_),
    .B(_0762_));
 sg13g2_nor2b_1 _4492_ (.A(_0758_),
    .B_N(_0764_),
    .Y(_0765_));
 sg13g2_xnor2_1 _4493_ (.Y(_0766_),
    .A(_0758_),
    .B(_0764_));
 sg13g2_nand2_1 _4494_ (.Y(_0767_),
    .A(_0750_),
    .B(_0766_));
 sg13g2_xnor2_1 _4495_ (.Y(_0768_),
    .A(_0750_),
    .B(_0766_));
 sg13g2_nand2_1 _4496_ (.Y(_0769_),
    .A(net760),
    .B(net817));
 sg13g2_o21ai_1 _4497_ (.B1(_0698_),
    .Y(_0770_),
    .A1(_0695_),
    .A2(_0699_));
 sg13g2_nand2_1 _4498_ (.Y(_0771_),
    .A(net757),
    .B(net822));
 sg13g2_nand2b_1 _4499_ (.Y(_0772_),
    .B(_0770_),
    .A_N(_0771_));
 sg13g2_xnor2_1 _4500_ (.Y(_0773_),
    .A(_0770_),
    .B(_0771_));
 sg13g2_nand2b_1 _4501_ (.Y(_0774_),
    .B(_0773_),
    .A_N(_0769_));
 sg13g2_xnor2_1 _4502_ (.Y(_0775_),
    .A(_0769_),
    .B(_0773_));
 sg13g2_inv_1 _4503_ (.Y(_0776_),
    .A(_0775_));
 sg13g2_xnor2_1 _4504_ (.Y(_0777_),
    .A(_0768_),
    .B(_0775_));
 sg13g2_nor2b_1 _4505_ (.A(_0749_),
    .B_N(_0777_),
    .Y(_0778_));
 sg13g2_xnor2_1 _4506_ (.Y(_0779_),
    .A(_0749_),
    .B(_0777_));
 sg13g2_xnor2_1 _4507_ (.Y(_0780_),
    .A(_0748_),
    .B(_0779_));
 sg13g2_nor2_1 _4508_ (.A(_0747_),
    .B(_0780_),
    .Y(_0781_));
 sg13g2_xor2_1 _4509_ (.B(_0780_),
    .A(_0747_),
    .X(_0782_));
 sg13g2_xor2_1 _4510_ (.B(_0782_),
    .A(_0746_),
    .X(_0783_));
 sg13g2_and2_1 _4511_ (.A(_0021_),
    .B(_0783_),
    .X(_0784_));
 sg13g2_or2_1 _4512_ (.X(_0785_),
    .B(_0783_),
    .A(_0021_));
 sg13g2_xnor2_1 _4513_ (.Y(_0786_),
    .A(_0021_),
    .B(_0783_));
 sg13g2_xnor2_1 _4514_ (.Y(_0787_),
    .A(_0745_),
    .B(_0786_));
 sg13g2_xor2_1 _4515_ (.B(_0786_),
    .A(_0745_),
    .X(_0788_));
 sg13g2_nor2_2 _4516_ (.A(net740),
    .B(_0721_),
    .Y(_0789_));
 sg13g2_nand2_1 _4517_ (.Y(_0790_),
    .A(net767),
    .B(net700));
 sg13g2_nand2_1 _4518_ (.Y(_0791_),
    .A(net771),
    .B(net700));
 sg13g2_inv_1 _4519_ (.Y(_0792_),
    .A(_0791_));
 sg13g2_nor3_1 _4520_ (.A(net734),
    .B(_0721_),
    .C(_0725_),
    .Y(_0793_));
 sg13g2_nand3_1 _4521_ (.B(net699),
    .C(_0728_),
    .A(net767),
    .Y(_0794_));
 sg13g2_a21oi_1 _4522_ (.A1(net770),
    .A2(net700),
    .Y(_0795_),
    .B1(_0724_));
 sg13g2_o21ai_1 _4523_ (.B1(_0725_),
    .Y(_0796_),
    .A1(net734),
    .A2(_0721_));
 sg13g2_a21oi_1 _4524_ (.A1(net770),
    .A2(net700),
    .Y(_0797_),
    .B1(_0725_));
 sg13g2_nor3_1 _4525_ (.A(net734),
    .B(_0721_),
    .C(_0724_),
    .Y(_0798_));
 sg13g2_nor4_2 _4526_ (.A(net732),
    .B(net696),
    .C(_0793_),
    .Y(_0799_),
    .D(_0795_));
 sg13g2_a22oi_1 _4527_ (.Y(_0800_),
    .B1(_0794_),
    .B2(_0796_),
    .A2(net697),
    .A1(net777));
 sg13g2_nor4_1 _4528_ (.A(net732),
    .B(net696),
    .C(_0797_),
    .D(_0798_),
    .Y(_0801_));
 sg13g2_a221oi_1 _4529_ (.B2(_0728_),
    .C1(_0795_),
    .B1(_0789_),
    .A1(net776),
    .Y(_0802_),
    .A2(net697));
 sg13g2_a21oi_2 _4530_ (.B1(_0614_),
    .Y(_0803_),
    .A2(_0612_),
    .A1(_0583_));
 sg13g2_nand2_1 _4531_ (.Y(_0804_),
    .A(net764),
    .B(net703));
 sg13g2_and2_1 _4532_ (.A(_1472_),
    .B(_0611_),
    .X(_0805_));
 sg13g2_a22oi_1 _4533_ (.Y(_0806_),
    .B1(_0611_),
    .B2(net761),
    .A2(_0582_),
    .A1(_1472_));
 sg13g2_a21o_1 _4534_ (.A2(_0805_),
    .A1(_0583_),
    .B1(_0806_),
    .X(_0807_));
 sg13g2_nor2_1 _4535_ (.A(_0804_),
    .B(_0807_),
    .Y(_0808_));
 sg13g2_xor2_1 _4536_ (.B(_0807_),
    .A(_0804_),
    .X(_0809_));
 sg13g2_nor2b_1 _4537_ (.A(_0803_),
    .B_N(_0809_),
    .Y(_0810_));
 sg13g2_xnor2_1 _4538_ (.Y(_0811_),
    .A(_0803_),
    .B(_0809_));
 sg13g2_xor2_1 _4539_ (.B(_0809_),
    .A(_0803_),
    .X(_0812_));
 sg13g2_nor3_2 _4540_ (.A(_0799_),
    .B(_0800_),
    .C(_0812_),
    .Y(_0813_));
 sg13g2_o21ai_1 _4541_ (.B1(_0811_),
    .Y(_0814_),
    .A1(_0801_),
    .A2(_0802_));
 sg13g2_nor3_1 _4542_ (.A(_0801_),
    .B(_0802_),
    .C(_0811_),
    .Y(_0815_));
 sg13g2_o21ai_1 _4543_ (.B1(_0812_),
    .Y(_0816_),
    .A1(_0799_),
    .A2(_0800_));
 sg13g2_nor3_1 _4544_ (.A(_0742_),
    .B(_0813_),
    .C(_0815_),
    .Y(_0817_));
 sg13g2_a21oi_2 _4545_ (.B1(_0784_),
    .Y(_0818_),
    .A2(_0785_),
    .A1(_0745_));
 sg13g2_a21oi_1 _4546_ (.A1(_0746_),
    .A2(_0782_),
    .Y(_0819_),
    .B1(_0781_));
 sg13g2_a21oi_2 _4547_ (.B1(_0778_),
    .Y(_0820_),
    .A2(_0779_),
    .A1(_0748_));
 sg13g2_nand2_1 _4548_ (.Y(_0821_),
    .A(_0772_),
    .B(_0774_));
 sg13g2_inv_1 _4549_ (.Y(_0822_),
    .A(_0821_));
 sg13g2_o21ai_1 _4550_ (.B1(_0767_),
    .Y(_0823_),
    .A1(_0768_),
    .A2(_0776_));
 sg13g2_a21o_1 _4551_ (.A2(_0757_),
    .A1(_0751_),
    .B1(_0765_),
    .X(_0824_));
 sg13g2_o21ai_1 _4552_ (.B1(_0756_),
    .Y(_0825_),
    .A1(_0650_),
    .A2(_0753_));
 sg13g2_nand2_1 _4553_ (.Y(_0826_),
    .A(net747),
    .B(net840));
 sg13g2_nand2_1 _4554_ (.Y(_0827_),
    .A(net744),
    .B(net851));
 sg13g2_nand2_1 _4555_ (.Y(_0828_),
    .A(net745),
    .B(net846));
 sg13g2_xor2_1 _4556_ (.B(_0828_),
    .A(_0753_),
    .X(_0829_));
 sg13g2_nand2b_1 _4557_ (.Y(_0830_),
    .B(_0829_),
    .A_N(_0826_));
 sg13g2_xnor2_1 _4558_ (.Y(_0831_),
    .A(_0826_),
    .B(_0829_));
 sg13g2_xnor2_1 _4559_ (.Y(_0832_),
    .A(_0825_),
    .B(_0831_));
 sg13g2_nand2_1 _4560_ (.Y(_0833_),
    .A(net755),
    .B(net822));
 sg13g2_nand2_1 _4561_ (.Y(_0834_),
    .A(net750),
    .B(net827));
 sg13g2_nand2_1 _4562_ (.Y(_0835_),
    .A(net752),
    .B(net827));
 sg13g2_xor2_1 _4563_ (.B(_0835_),
    .A(_0760_),
    .X(_0836_));
 sg13g2_nand2b_1 _4564_ (.Y(_0837_),
    .B(_0836_),
    .A_N(_0833_));
 sg13g2_xnor2_1 _4565_ (.Y(_0838_),
    .A(_0833_),
    .B(_0836_));
 sg13g2_nor2b_1 _4566_ (.A(_0832_),
    .B_N(_0838_),
    .Y(_0839_));
 sg13g2_xnor2_1 _4567_ (.Y(_0840_),
    .A(_0832_),
    .B(_0838_));
 sg13g2_nand2_1 _4568_ (.Y(_0841_),
    .A(_0824_),
    .B(_0840_));
 sg13g2_xnor2_1 _4569_ (.Y(_0842_),
    .A(_0824_),
    .B(_0840_));
 sg13g2_nand2_1 _4570_ (.Y(_0843_),
    .A(net760),
    .B(net813));
 sg13g2_o21ai_1 _4571_ (.B1(_0763_),
    .Y(_0844_),
    .A1(_0696_),
    .A2(_0761_));
 sg13g2_nand2_1 _4572_ (.Y(_0845_),
    .A(net757),
    .B(net817));
 sg13g2_nand2b_1 _4573_ (.Y(_0846_),
    .B(_0844_),
    .A_N(_0845_));
 sg13g2_xnor2_1 _4574_ (.Y(_0847_),
    .A(_0844_),
    .B(_0845_));
 sg13g2_nand2b_1 _4575_ (.Y(_0848_),
    .B(_0847_),
    .A_N(_0843_));
 sg13g2_xnor2_1 _4576_ (.Y(_0849_),
    .A(_0843_),
    .B(_0847_));
 sg13g2_inv_1 _4577_ (.Y(_0850_),
    .A(_0849_));
 sg13g2_xnor2_1 _4578_ (.Y(_0851_),
    .A(_0842_),
    .B(_0849_));
 sg13g2_nand2_1 _4579_ (.Y(_0852_),
    .A(_0823_),
    .B(_0851_));
 sg13g2_xnor2_1 _4580_ (.Y(_0853_),
    .A(_0823_),
    .B(_0851_));
 sg13g2_xnor2_1 _4581_ (.Y(_0854_),
    .A(_0822_),
    .B(_0853_));
 sg13g2_or2_1 _4582_ (.X(_0855_),
    .B(_0854_),
    .A(_0820_));
 sg13g2_and2_1 _4583_ (.A(_0820_),
    .B(_0854_),
    .X(_0856_));
 sg13g2_xor2_1 _4584_ (.B(_0854_),
    .A(_0820_),
    .X(_0857_));
 sg13g2_xnor2_1 _4585_ (.Y(_0858_),
    .A(_0819_),
    .B(_0857_));
 sg13g2_xnor2_1 _4586_ (.Y(_0859_),
    .A(_0015_),
    .B(_0858_));
 sg13g2_nand2b_1 _4587_ (.Y(_0860_),
    .B(_0858_),
    .A_N(\system_inst.neuron.u[4] ));
 sg13g2_o21ai_1 _4588_ (.B1(_0860_),
    .Y(_0861_),
    .A1(_0818_),
    .A2(_0859_));
 sg13g2_o21ai_1 _4589_ (.B1(_0855_),
    .Y(_0862_),
    .A1(_0819_),
    .A2(_0856_));
 sg13g2_o21ai_1 _4590_ (.B1(_0852_),
    .Y(_0863_),
    .A1(_0822_),
    .A2(_0853_));
 sg13g2_nand2_1 _4591_ (.Y(_0864_),
    .A(_0846_),
    .B(_0848_));
 sg13g2_inv_1 _4592_ (.Y(_0865_),
    .A(_0864_));
 sg13g2_o21ai_1 _4593_ (.B1(_0841_),
    .Y(_0866_),
    .A1(_0842_),
    .A2(_0850_));
 sg13g2_a21o_1 _4594_ (.A2(_0831_),
    .A1(_0825_),
    .B1(_0839_),
    .X(_0867_));
 sg13g2_o21ai_1 _4595_ (.B1(_0830_),
    .Y(_0868_),
    .A1(_0753_),
    .A2(_0828_));
 sg13g2_nand2_1 _4596_ (.Y(_0869_),
    .A(net747),
    .B(net835));
 sg13g2_nand2_1 _4597_ (.Y(_0870_),
    .A(net744),
    .B(net841));
 sg13g2_nand2_1 _4598_ (.Y(_0871_),
    .A(net745),
    .B(net840));
 sg13g2_xor2_1 _4599_ (.B(_0871_),
    .A(_0827_),
    .X(_0872_));
 sg13g2_nand2b_1 _4600_ (.Y(_0873_),
    .B(_0872_),
    .A_N(_0869_));
 sg13g2_xnor2_1 _4601_ (.Y(_0874_),
    .A(_0869_),
    .B(_0872_));
 sg13g2_xnor2_1 _4602_ (.Y(_0875_),
    .A(_0868_),
    .B(_0874_));
 sg13g2_nand2_1 _4603_ (.Y(_0876_),
    .A(net755),
    .B(net817));
 sg13g2_nand2_2 _4604_ (.Y(_0877_),
    .A(\system_inst.internal_param_b[4] ),
    .B(net822));
 sg13g2_nand2_1 _4605_ (.Y(_0878_),
    .A(net752),
    .B(net822));
 sg13g2_xor2_1 _4606_ (.B(_0878_),
    .A(_0834_),
    .X(_0879_));
 sg13g2_nand2b_1 _4607_ (.Y(_0880_),
    .B(_0879_),
    .A_N(_0876_));
 sg13g2_xnor2_1 _4608_ (.Y(_0881_),
    .A(_0876_),
    .B(_0879_));
 sg13g2_nor2b_1 _4609_ (.A(_0875_),
    .B_N(_0881_),
    .Y(_0882_));
 sg13g2_xnor2_1 _4610_ (.Y(_0883_),
    .A(_0875_),
    .B(_0881_));
 sg13g2_nand2_1 _4611_ (.Y(_0884_),
    .A(_0867_),
    .B(_0883_));
 sg13g2_xnor2_1 _4612_ (.Y(_0885_),
    .A(_0867_),
    .B(_0883_));
 sg13g2_nand2_1 _4613_ (.Y(_0886_),
    .A(net760),
    .B(net812));
 sg13g2_o21ai_1 _4614_ (.B1(_0837_),
    .Y(_0887_),
    .A1(_0760_),
    .A2(_0835_));
 sg13g2_nand2_1 _4615_ (.Y(_0888_),
    .A(net757),
    .B(net813));
 sg13g2_nand2b_1 _4616_ (.Y(_0889_),
    .B(_0887_),
    .A_N(_0888_));
 sg13g2_xnor2_1 _4617_ (.Y(_0890_),
    .A(_0887_),
    .B(_0888_));
 sg13g2_nand2b_1 _4618_ (.Y(_0891_),
    .B(_0890_),
    .A_N(_0886_));
 sg13g2_xnor2_1 _4619_ (.Y(_0892_),
    .A(_0886_),
    .B(_0890_));
 sg13g2_inv_1 _4620_ (.Y(_0893_),
    .A(_0892_));
 sg13g2_xnor2_1 _4621_ (.Y(_0894_),
    .A(_0885_),
    .B(_0892_));
 sg13g2_nand2_1 _4622_ (.Y(_0895_),
    .A(_0866_),
    .B(_0894_));
 sg13g2_xnor2_1 _4623_ (.Y(_0896_),
    .A(_0866_),
    .B(_0894_));
 sg13g2_xnor2_1 _4624_ (.Y(_0897_),
    .A(_0865_),
    .B(_0896_));
 sg13g2_nor2b_1 _4625_ (.A(_0897_),
    .B_N(_0863_),
    .Y(_0898_));
 sg13g2_xor2_1 _4626_ (.B(_0897_),
    .A(_0863_),
    .X(_0899_));
 sg13g2_inv_1 _4627_ (.Y(_0900_),
    .A(_0899_));
 sg13g2_xnor2_1 _4628_ (.Y(_0901_),
    .A(_0862_),
    .B(_0899_));
 sg13g2_and2_1 _4629_ (.A(_0014_),
    .B(_0901_),
    .X(_0902_));
 sg13g2_or2_1 _4630_ (.X(_0903_),
    .B(_0901_),
    .A(_0014_));
 sg13g2_xnor2_1 _4631_ (.Y(_0904_),
    .A(_0014_),
    .B(_0901_));
 sg13g2_xnor2_1 _4632_ (.Y(_0905_),
    .A(_0861_),
    .B(_0904_));
 sg13g2_xor2_1 _4633_ (.B(_0904_),
    .A(_0861_),
    .X(_0906_));
 sg13g2_nand2_2 _4634_ (.Y(_0907_),
    .A(_0731_),
    .B(_0736_));
 sg13g2_xor2_1 _4635_ (.B(_0859_),
    .A(_0818_),
    .X(_0908_));
 sg13g2_xnor2_1 _4636_ (.Y(_0909_),
    .A(_0818_),
    .B(_0859_));
 sg13g2_nor2_1 _4637_ (.A(net728),
    .B(_0909_),
    .Y(_0910_));
 sg13g2_nand3_1 _4638_ (.B(_0907_),
    .C(net695),
    .A(net783),
    .Y(_0911_));
 sg13g2_a21o_1 _4639_ (.A2(net695),
    .A1(net783),
    .B1(_0907_),
    .X(_0912_));
 sg13g2_nand4_1 _4640_ (.B(_0731_),
    .C(_0736_),
    .A(net783),
    .Y(_0913_),
    .D(net695));
 sg13g2_o21ai_1 _4641_ (.B1(_0907_),
    .Y(_0914_),
    .A1(net728),
    .A2(_0909_));
 sg13g2_and4_1 _4642_ (.A(net790),
    .B(net693),
    .C(_0911_),
    .D(_0912_),
    .X(_0915_));
 sg13g2_a22oi_1 _4643_ (.Y(_0916_),
    .B1(_0911_),
    .B2(_0912_),
    .A2(net693),
    .A1(net789));
 sg13g2_and4_1 _4644_ (.A(net789),
    .B(net693),
    .C(_0913_),
    .D(_0914_),
    .X(_0917_));
 sg13g2_a22oi_1 _4645_ (.Y(_0918_),
    .B1(_0913_),
    .B2(_0914_),
    .A2(net693),
    .A1(net789));
 sg13g2_a21oi_1 _4646_ (.A1(_0814_),
    .A2(_0816_),
    .Y(_0919_),
    .B1(_0743_));
 sg13g2_a21oi_1 _4647_ (.A1(_0814_),
    .A2(_0816_),
    .Y(_0920_),
    .B1(_0742_));
 sg13g2_nor3_1 _4648_ (.A(_0743_),
    .B(_0813_),
    .C(_0815_),
    .Y(_0921_));
 sg13g2_or4_2 _4649_ (.A(_0817_),
    .B(_0915_),
    .C(_0916_),
    .D(_0919_),
    .X(_0922_));
 sg13g2_nor2b_1 _4650_ (.A(_0817_),
    .B_N(_0922_),
    .Y(_0923_));
 sg13g2_nand2b_1 _4651_ (.Y(_0924_),
    .B(_0922_),
    .A_N(_0817_));
 sg13g2_a21o_1 _4652_ (.A2(_0903_),
    .A1(_0861_),
    .B1(_0902_),
    .X(_0925_));
 sg13g2_a21o_1 _4653_ (.A2(_0900_),
    .A1(_0862_),
    .B1(_0898_),
    .X(_0926_));
 sg13g2_o21ai_1 _4654_ (.B1(_0895_),
    .Y(_0927_),
    .A1(_0865_),
    .A2(_0896_));
 sg13g2_nand2_1 _4655_ (.Y(_0928_),
    .A(_0889_),
    .B(_0891_));
 sg13g2_inv_1 _4656_ (.Y(_0929_),
    .A(_0928_));
 sg13g2_o21ai_1 _4657_ (.B1(_0884_),
    .Y(_0930_),
    .A1(_0885_),
    .A2(_0893_));
 sg13g2_a21o_1 _4658_ (.A2(_0874_),
    .A1(_0868_),
    .B1(_0882_),
    .X(_0931_));
 sg13g2_o21ai_1 _4659_ (.B1(_0873_),
    .Y(_0932_),
    .A1(_0827_),
    .A2(_0871_));
 sg13g2_nand2_1 _4660_ (.Y(_0933_),
    .A(net747),
    .B(net828));
 sg13g2_nand2_1 _4661_ (.Y(_0934_),
    .A(net743),
    .B(net834));
 sg13g2_nand2_1 _4662_ (.Y(_0935_),
    .A(net745),
    .B(net834));
 sg13g2_xor2_1 _4663_ (.B(_0935_),
    .A(_0870_),
    .X(_0936_));
 sg13g2_nand2b_1 _4664_ (.Y(_0937_),
    .B(_0936_),
    .A_N(_0933_));
 sg13g2_xnor2_1 _4665_ (.Y(_0938_),
    .A(_0933_),
    .B(_0936_));
 sg13g2_xnor2_1 _4666_ (.Y(_0939_),
    .A(_0932_),
    .B(_0938_));
 sg13g2_nand2_2 _4667_ (.Y(_0940_),
    .A(\system_inst.internal_param_b[2] ),
    .B(net813));
 sg13g2_nand2_1 _4668_ (.Y(_0941_),
    .A(net750),
    .B(net817));
 sg13g2_nand2_1 _4669_ (.Y(_0942_),
    .A(net752),
    .B(net817));
 sg13g2_xor2_1 _4670_ (.B(_0942_),
    .A(_0877_),
    .X(_0943_));
 sg13g2_nand2b_1 _4671_ (.Y(_0944_),
    .B(_0943_),
    .A_N(_0940_));
 sg13g2_xnor2_1 _4672_ (.Y(_0945_),
    .A(_0940_),
    .B(_0943_));
 sg13g2_nor2b_1 _4673_ (.A(_0939_),
    .B_N(_0945_),
    .Y(_0946_));
 sg13g2_xnor2_1 _4674_ (.Y(_0947_),
    .A(_0939_),
    .B(_0945_));
 sg13g2_nand2_1 _4675_ (.Y(_0948_),
    .A(_0931_),
    .B(_0947_));
 sg13g2_xnor2_1 _4676_ (.Y(_0949_),
    .A(_0931_),
    .B(_0947_));
 sg13g2_nand2_1 _4677_ (.Y(_0950_),
    .A(net760),
    .B(net807));
 sg13g2_o21ai_1 _4678_ (.B1(_0880_),
    .Y(_0951_),
    .A1(_0834_),
    .A2(_0878_));
 sg13g2_nand2_1 _4679_ (.Y(_0952_),
    .A(net757),
    .B(net812));
 sg13g2_nand2b_1 _4680_ (.Y(_0953_),
    .B(_0951_),
    .A_N(_0952_));
 sg13g2_xnor2_1 _4681_ (.Y(_0954_),
    .A(_0951_),
    .B(_0952_));
 sg13g2_nand2b_1 _4682_ (.Y(_0955_),
    .B(_0954_),
    .A_N(_0950_));
 sg13g2_xnor2_1 _4683_ (.Y(_0956_),
    .A(_0950_),
    .B(_0954_));
 sg13g2_inv_1 _4684_ (.Y(_0957_),
    .A(_0956_));
 sg13g2_xnor2_1 _4685_ (.Y(_0958_),
    .A(_0949_),
    .B(_0956_));
 sg13g2_nand2_1 _4686_ (.Y(_0959_),
    .A(_0930_),
    .B(_0958_));
 sg13g2_xnor2_1 _4687_ (.Y(_0960_),
    .A(_0930_),
    .B(_0958_));
 sg13g2_xnor2_1 _4688_ (.Y(_0961_),
    .A(_0929_),
    .B(_0960_));
 sg13g2_nor2b_1 _4689_ (.A(_0961_),
    .B_N(_0927_),
    .Y(_0962_));
 sg13g2_xor2_1 _4690_ (.B(_0961_),
    .A(_0927_),
    .X(_0963_));
 sg13g2_inv_1 _4691_ (.Y(_0964_),
    .A(_0963_));
 sg13g2_xnor2_1 _4692_ (.Y(_0965_),
    .A(_0926_),
    .B(_0964_));
 sg13g2_xnor2_1 _4693_ (.Y(_0966_),
    .A(_0013_),
    .B(_0965_));
 sg13g2_xor2_1 _4694_ (.B(_0966_),
    .A(_0925_),
    .X(_0967_));
 sg13g2_xnor2_1 _4695_ (.Y(_0968_),
    .A(_0925_),
    .B(_0966_));
 sg13g2_or2_1 _4696_ (.X(_0969_),
    .B(_0799_),
    .A(_0793_));
 sg13g2_nand3_1 _4697_ (.B(net693),
    .C(_0969_),
    .A(net784),
    .Y(_0970_));
 sg13g2_a21o_1 _4698_ (.A2(net693),
    .A1(net784),
    .B1(_0969_),
    .X(_0971_));
 sg13g2_or3_1 _4699_ (.A(net728),
    .B(_0906_),
    .C(_0969_),
    .X(_0972_));
 sg13g2_o21ai_1 _4700_ (.B1(_0969_),
    .Y(_0973_),
    .A1(net728),
    .A2(_0906_));
 sg13g2_and4_1 _4701_ (.A(net791),
    .B(net689),
    .C(_0970_),
    .D(_0971_),
    .X(_0974_));
 sg13g2_nand4_1 _4702_ (.B(net689),
    .C(_0970_),
    .A(net791),
    .Y(_0975_),
    .D(_0971_));
 sg13g2_a22oi_1 _4703_ (.Y(_0976_),
    .B1(_0970_),
    .B2(_0971_),
    .A2(net689),
    .A1(net791));
 sg13g2_and4_1 _4704_ (.A(net791),
    .B(net689),
    .C(_0972_),
    .D(_0973_),
    .X(_0977_));
 sg13g2_a22oi_1 _4705_ (.Y(_0978_),
    .B1(_0972_),
    .B2(_0973_),
    .A2(net689),
    .A1(net791));
 sg13g2_nor2_1 _4706_ (.A(_0810_),
    .B(_0813_),
    .Y(_0979_));
 sg13g2_nand2b_1 _4707_ (.Y(_0980_),
    .B(_0814_),
    .A_N(_0810_));
 sg13g2_nor2_2 _4708_ (.A(net740),
    .B(_0788_),
    .Y(_0981_));
 sg13g2_nand2_1 _4709_ (.Y(_0982_),
    .A(net768),
    .B(net698));
 sg13g2_nor3_1 _4710_ (.A(net740),
    .B(net696),
    .C(_0791_),
    .Y(_0983_));
 sg13g2_nand3_1 _4711_ (.B(net698),
    .C(_0789_),
    .A(net771),
    .Y(_0984_));
 sg13g2_a21oi_1 _4712_ (.A1(net771),
    .A2(net698),
    .Y(_0985_),
    .B1(_0789_));
 sg13g2_o21ai_1 _4713_ (.B1(_0790_),
    .Y(_0986_),
    .A1(net735),
    .A2(net696));
 sg13g2_a21oi_1 _4714_ (.A1(net771),
    .A2(net698),
    .Y(_0987_),
    .B1(_0790_));
 sg13g2_nor3_1 _4715_ (.A(net734),
    .B(net696),
    .C(_0789_),
    .Y(_0988_));
 sg13g2_nor4_2 _4716_ (.A(net732),
    .B(_0909_),
    .C(_0983_),
    .Y(_0989_),
    .D(_0985_));
 sg13g2_a22oi_1 _4717_ (.Y(_0990_),
    .B1(_0984_),
    .B2(_0986_),
    .A2(net694),
    .A1(net778));
 sg13g2_nor4_2 _4718_ (.A(net732),
    .B(_0909_),
    .C(_0987_),
    .Y(_0991_),
    .D(_0988_));
 sg13g2_a221oi_1 _4719_ (.B2(_0792_),
    .C1(_0985_),
    .B1(_0981_),
    .A1(net778),
    .Y(_0992_),
    .A2(net694));
 sg13g2_a21oi_1 _4720_ (.A1(_0583_),
    .A2(_0805_),
    .Y(_0993_),
    .B1(_0808_));
 sg13g2_nand2_1 _4721_ (.Y(_0994_),
    .A(net764),
    .B(net702));
 sg13g2_nand3_1 _4722_ (.B(net704),
    .C(_0805_),
    .A(net761),
    .Y(_0995_));
 sg13g2_a21o_1 _4723_ (.A2(net704),
    .A1(net761),
    .B1(_0805_),
    .X(_0996_));
 sg13g2_nand2_1 _4724_ (.Y(_0997_),
    .A(_0995_),
    .B(_0996_));
 sg13g2_xor2_1 _4725_ (.B(_0997_),
    .A(_0994_),
    .X(_0998_));
 sg13g2_nor2b_1 _4726_ (.A(_0993_),
    .B_N(_0998_),
    .Y(_0999_));
 sg13g2_xor2_1 _4727_ (.B(_0998_),
    .A(_0993_),
    .X(_1000_));
 sg13g2_inv_1 _4728_ (.Y(_1001_),
    .A(_1000_));
 sg13g2_nor3_2 _4729_ (.A(_0989_),
    .B(_0990_),
    .C(_1000_),
    .Y(_1002_));
 sg13g2_o21ai_1 _4730_ (.B1(_1001_),
    .Y(_1003_),
    .A1(_0991_),
    .A2(_0992_));
 sg13g2_nor3_2 _4731_ (.A(_0991_),
    .B(_0992_),
    .C(_1001_),
    .Y(_1004_));
 sg13g2_o21ai_1 _4732_ (.B1(_1000_),
    .Y(_1005_),
    .A1(_0989_),
    .A2(_0990_));
 sg13g2_nor3_2 _4733_ (.A(_0979_),
    .B(_1002_),
    .C(_1004_),
    .Y(_1006_));
 sg13g2_a21oi_1 _4734_ (.A1(_1003_),
    .A2(_1005_),
    .Y(_1007_),
    .B1(_0980_));
 sg13g2_a21oi_1 _4735_ (.A1(_1003_),
    .A2(_1005_),
    .Y(_1008_),
    .B1(_0979_));
 sg13g2_nor3_2 _4736_ (.A(_0980_),
    .B(_1002_),
    .C(_1004_),
    .Y(_1009_));
 sg13g2_nor4_2 _4737_ (.A(_0974_),
    .B(_0976_),
    .C(_1006_),
    .Y(_1010_),
    .D(_1007_));
 sg13g2_or4_1 _4738_ (.A(_0974_),
    .B(_0976_),
    .C(_1006_),
    .D(_1007_),
    .X(_1011_));
 sg13g2_nor4_2 _4739_ (.A(_0977_),
    .B(_0978_),
    .C(_1008_),
    .Y(_1012_),
    .D(_1009_));
 sg13g2_or4_1 _4740_ (.A(_0977_),
    .B(_0978_),
    .C(_1008_),
    .D(_1009_),
    .X(_1013_));
 sg13g2_nor3_1 _4741_ (.A(_0923_),
    .B(_1010_),
    .C(_1012_),
    .Y(_1014_));
 sg13g2_nand3_1 _4742_ (.B(_1011_),
    .C(_1013_),
    .A(_0924_),
    .Y(_1015_));
 sg13g2_a21oi_2 _4743_ (.B1(_0915_),
    .Y(_1016_),
    .A2(_0910_),
    .A1(_0907_));
 sg13g2_inv_1 _4744_ (.Y(_1017_),
    .A(_1016_));
 sg13g2_a21oi_1 _4745_ (.A1(_1011_),
    .A2(_1013_),
    .Y(_1018_),
    .B1(_0924_));
 sg13g2_o21ai_1 _4746_ (.B1(_0923_),
    .Y(_1019_),
    .A1(_1010_),
    .A2(_1012_));
 sg13g2_nor3_2 _4747_ (.A(_1014_),
    .B(_1016_),
    .C(_1018_),
    .Y(_1020_));
 sg13g2_nor2_1 _4748_ (.A(_1014_),
    .B(_1020_),
    .Y(_1021_));
 sg13g2_o21ai_1 _4749_ (.B1(_1015_),
    .Y(_1022_),
    .A1(_1016_),
    .A2(_1018_));
 sg13g2_nand2_1 _4750_ (.Y(_1023_),
    .A(_0970_),
    .B(_0975_));
 sg13g2_nor2_1 _4751_ (.A(_1006_),
    .B(_1010_),
    .Y(_1024_));
 sg13g2_nor2_1 _4752_ (.A(_0999_),
    .B(_1002_),
    .Y(_1025_));
 sg13g2_nand2b_1 _4753_ (.Y(_1026_),
    .B(_1003_),
    .A_N(_0999_));
 sg13g2_o21ai_1 _4754_ (.B1(_0995_),
    .Y(_1027_),
    .A1(_0994_),
    .A2(_0997_));
 sg13g2_nand2_1 _4755_ (.Y(_1028_),
    .A(net765),
    .B(net700));
 sg13g2_nand2_1 _4756_ (.Y(_1029_),
    .A(net762),
    .B(net702));
 sg13g2_nand2_1 _4757_ (.Y(_1030_),
    .A(\system_inst.internal_param_a[7] ),
    .B(net704));
 sg13g2_xor2_1 _4758_ (.B(_1030_),
    .A(_1029_),
    .X(_1031_));
 sg13g2_nand2b_1 _4759_ (.Y(_1032_),
    .B(_1031_),
    .A_N(_1028_));
 sg13g2_xnor2_1 _4760_ (.Y(_1033_),
    .A(_1028_),
    .B(_1031_));
 sg13g2_xor2_1 _4761_ (.B(_1033_),
    .A(_1027_),
    .X(_1034_));
 sg13g2_xnor2_1 _4762_ (.Y(_1035_),
    .A(_1027_),
    .B(_1033_));
 sg13g2_nor2_1 _4763_ (.A(net740),
    .B(_0909_),
    .Y(_1036_));
 sg13g2_nand2_1 _4764_ (.Y(_1037_),
    .A(net768),
    .B(net694));
 sg13g2_nand2_1 _4765_ (.Y(_1038_),
    .A(net772),
    .B(net694));
 sg13g2_inv_1 _4766_ (.Y(_1039_),
    .A(_1038_));
 sg13g2_nand3_1 _4767_ (.B(net694),
    .C(_0981_),
    .A(net772),
    .Y(_1040_));
 sg13g2_o21ai_1 _4768_ (.B1(_0982_),
    .Y(_1041_),
    .A1(net735),
    .A2(_0909_));
 sg13g2_o21ai_1 _4769_ (.B1(_0981_),
    .Y(_1042_),
    .A1(net735),
    .A2(_0909_));
 sg13g2_nand3_1 _4770_ (.B(net694),
    .C(_0982_),
    .A(net772),
    .Y(_1043_));
 sg13g2_and4_1 _4771_ (.A(net779),
    .B(net692),
    .C(_1040_),
    .D(_1041_),
    .X(_1044_));
 sg13g2_a22oi_1 _4772_ (.Y(_1045_),
    .B1(_1040_),
    .B2(_1041_),
    .A2(net692),
    .A1(net779));
 sg13g2_and4_1 _4773_ (.A(net779),
    .B(net692),
    .C(_1042_),
    .D(_1043_),
    .X(_1046_));
 sg13g2_a22oi_1 _4774_ (.Y(_1047_),
    .B1(_1042_),
    .B2(_1043_),
    .A2(net692),
    .A1(net779));
 sg13g2_nor3_2 _4775_ (.A(_1035_),
    .B(_1044_),
    .C(_1045_),
    .Y(_1048_));
 sg13g2_o21ai_1 _4776_ (.B1(_1034_),
    .Y(_1049_),
    .A1(_1046_),
    .A2(_1047_));
 sg13g2_nor3_1 _4777_ (.A(_1034_),
    .B(_1046_),
    .C(_1047_),
    .Y(_1050_));
 sg13g2_o21ai_1 _4778_ (.B1(_1035_),
    .Y(_1051_),
    .A1(_1044_),
    .A2(_1045_));
 sg13g2_nor3_1 _4779_ (.A(_1025_),
    .B(_1048_),
    .C(_1050_),
    .Y(_1052_));
 sg13g2_a21oi_1 _4780_ (.A1(_1049_),
    .A2(_1051_),
    .Y(_1053_),
    .B1(_1026_));
 sg13g2_a21oi_1 _4781_ (.A1(_1049_),
    .A2(_1051_),
    .Y(_1054_),
    .B1(_1025_));
 sg13g2_nor3_1 _4782_ (.A(_1026_),
    .B(_1048_),
    .C(_1050_),
    .Y(_1055_));
 sg13g2_nor2_1 _4783_ (.A(\system_inst.neuron.u[6] ),
    .B(_0965_),
    .Y(_1056_));
 sg13g2_a21oi_2 _4784_ (.B1(_1056_),
    .Y(_1057_),
    .A2(_0966_),
    .A1(_0925_));
 sg13g2_a21oi_1 _4785_ (.A1(_0926_),
    .A2(_0964_),
    .Y(_1058_),
    .B1(_0962_));
 sg13g2_o21ai_1 _4786_ (.B1(_0959_),
    .Y(_1059_),
    .A1(_0929_),
    .A2(_0960_));
 sg13g2_nand2_1 _4787_ (.Y(_1060_),
    .A(_0953_),
    .B(_0955_));
 sg13g2_inv_1 _4788_ (.Y(_1061_),
    .A(_1060_));
 sg13g2_o21ai_1 _4789_ (.B1(_0948_),
    .Y(_1062_),
    .A1(_0949_),
    .A2(_0957_));
 sg13g2_a21o_1 _4790_ (.A2(_0938_),
    .A1(_0932_),
    .B1(_0946_),
    .X(_1063_));
 sg13g2_o21ai_1 _4791_ (.B1(_0937_),
    .Y(_1064_),
    .A1(_0870_),
    .A2(_0935_));
 sg13g2_nand2_1 _4792_ (.Y(_1065_),
    .A(net748),
    .B(net822));
 sg13g2_nand2_1 _4793_ (.Y(_1066_),
    .A(net743),
    .B(net827));
 sg13g2_nand2_1 _4794_ (.Y(_1067_),
    .A(net746),
    .B(net828));
 sg13g2_xor2_1 _4795_ (.B(_1067_),
    .A(_0934_),
    .X(_1068_));
 sg13g2_nand2b_1 _4796_ (.Y(_1069_),
    .B(_1068_),
    .A_N(_1065_));
 sg13g2_xnor2_1 _4797_ (.Y(_1070_),
    .A(_1065_),
    .B(_1068_));
 sg13g2_xnor2_1 _4798_ (.Y(_1071_),
    .A(_1064_),
    .B(_1070_));
 sg13g2_nand2_1 _4799_ (.Y(_1072_),
    .A(net755),
    .B(net809));
 sg13g2_nand2_2 _4800_ (.Y(_1073_),
    .A(net753),
    .B(net813));
 sg13g2_xor2_1 _4801_ (.B(_1073_),
    .A(_0941_),
    .X(_1074_));
 sg13g2_nand2b_1 _4802_ (.Y(_1075_),
    .B(_1074_),
    .A_N(_1072_));
 sg13g2_xnor2_1 _4803_ (.Y(_1076_),
    .A(_1072_),
    .B(_1074_));
 sg13g2_nor2b_1 _4804_ (.A(_1071_),
    .B_N(_1076_),
    .Y(_1077_));
 sg13g2_xnor2_1 _4805_ (.Y(_1078_),
    .A(_1071_),
    .B(_1076_));
 sg13g2_nand2_1 _4806_ (.Y(_1079_),
    .A(_1063_),
    .B(_1078_));
 sg13g2_xnor2_1 _4807_ (.Y(_1080_),
    .A(_1063_),
    .B(_1078_));
 sg13g2_nand2_1 _4808_ (.Y(_1081_),
    .A(net760),
    .B(net804));
 sg13g2_o21ai_1 _4809_ (.B1(_0944_),
    .Y(_1082_),
    .A1(_0877_),
    .A2(_0942_));
 sg13g2_nand2_1 _4810_ (.Y(_1083_),
    .A(net757),
    .B(net807));
 sg13g2_nand2b_1 _4811_ (.Y(_1084_),
    .B(_1082_),
    .A_N(_1083_));
 sg13g2_xnor2_1 _4812_ (.Y(_1085_),
    .A(_1082_),
    .B(_1083_));
 sg13g2_nand2b_1 _4813_ (.Y(_1086_),
    .B(_1085_),
    .A_N(_1081_));
 sg13g2_xnor2_1 _4814_ (.Y(_1087_),
    .A(_1081_),
    .B(_1085_));
 sg13g2_inv_1 _4815_ (.Y(_1088_),
    .A(_1087_));
 sg13g2_xnor2_1 _4816_ (.Y(_1089_),
    .A(_1080_),
    .B(_1087_));
 sg13g2_nand2_1 _4817_ (.Y(_1090_),
    .A(_1062_),
    .B(_1089_));
 sg13g2_xnor2_1 _4818_ (.Y(_1091_),
    .A(_1062_),
    .B(_1089_));
 sg13g2_xnor2_1 _4819_ (.Y(_1092_),
    .A(_1061_),
    .B(_1091_));
 sg13g2_nand2b_1 _4820_ (.Y(_1093_),
    .B(_1059_),
    .A_N(_1092_));
 sg13g2_xor2_1 _4821_ (.B(_1092_),
    .A(_1059_),
    .X(_1094_));
 sg13g2_xor2_1 _4822_ (.B(_1094_),
    .A(_1058_),
    .X(_1095_));
 sg13g2_nand2_1 _4823_ (.Y(_1096_),
    .A(_0012_),
    .B(_1095_));
 sg13g2_xnor2_1 _4824_ (.Y(_1097_),
    .A(_0012_),
    .B(_1095_));
 sg13g2_xor2_1 _4825_ (.B(_1097_),
    .A(_1057_),
    .X(_1098_));
 sg13g2_xnor2_1 _4826_ (.Y(_1099_),
    .A(_1057_),
    .B(_1097_));
 sg13g2_or2_2 _4827_ (.X(_1100_),
    .B(_0989_),
    .A(_0983_));
 sg13g2_and3_1 _4828_ (.X(_1101_),
    .A(net788),
    .B(net689),
    .C(_1100_));
 sg13g2_nand3_1 _4829_ (.B(net689),
    .C(_1100_),
    .A(net785),
    .Y(_1102_));
 sg13g2_a21o_1 _4830_ (.A2(net689),
    .A1(net785),
    .B1(_1100_),
    .X(_1103_));
 sg13g2_or3_1 _4831_ (.A(net729),
    .B(net688),
    .C(_1100_),
    .X(_1104_));
 sg13g2_o21ai_1 _4832_ (.B1(_1100_),
    .Y(_1105_),
    .A1(net729),
    .A2(net688));
 sg13g2_and4_1 _4833_ (.A(net793),
    .B(net686),
    .C(_1102_),
    .D(_1103_),
    .X(_1106_));
 sg13g2_a22oi_1 _4834_ (.Y(_1107_),
    .B1(_1102_),
    .B2(_1103_),
    .A2(net686),
    .A1(net793));
 sg13g2_and4_1 _4835_ (.A(net793),
    .B(net686),
    .C(_1104_),
    .D(_1105_),
    .X(_1108_));
 sg13g2_a22oi_1 _4836_ (.Y(_1109_),
    .B1(_1104_),
    .B2(_1105_),
    .A2(net686),
    .A1(net793));
 sg13g2_nor4_2 _4837_ (.A(_1052_),
    .B(_1053_),
    .C(_1106_),
    .Y(_1110_),
    .D(_1107_));
 sg13g2_nor4_1 _4838_ (.A(_1054_),
    .B(_1055_),
    .C(_1108_),
    .D(_1109_),
    .Y(_1111_));
 sg13g2_or3_1 _4839_ (.A(_1024_),
    .B(_1110_),
    .C(_1111_),
    .X(_1112_));
 sg13g2_o21ai_1 _4840_ (.B1(_1024_),
    .Y(_1113_),
    .A1(_1110_),
    .A2(_1111_));
 sg13g2_nand3_1 _4841_ (.B(_1112_),
    .C(_1113_),
    .A(_1023_),
    .Y(_1114_));
 sg13g2_a21o_1 _4842_ (.A2(_1113_),
    .A1(_1112_),
    .B1(_1023_),
    .X(_1115_));
 sg13g2_nand3_1 _4843_ (.B(_1114_),
    .C(_1115_),
    .A(_1022_),
    .Y(_1116_));
 sg13g2_a21oi_1 _4844_ (.A1(_1114_),
    .A2(_1115_),
    .Y(_1117_),
    .B1(_1022_));
 sg13g2_a21oi_1 _4845_ (.A1(_1114_),
    .A2(_1115_),
    .Y(_1118_),
    .B1(_1021_));
 sg13g2_nand3_1 _4846_ (.B(_1114_),
    .C(_1115_),
    .A(_1021_),
    .Y(_1119_));
 sg13g2_nor2b_1 _4847_ (.A(_1118_),
    .B_N(_1119_),
    .Y(_1120_));
 sg13g2_nand2_2 _4848_ (.Y(_1121_),
    .A(net767),
    .B(net705));
 sg13g2_xor2_1 _4849_ (.B(_1121_),
    .A(_0727_),
    .X(_1122_));
 sg13g2_a21o_1 _4850_ (.A2(net701),
    .A1(net776),
    .B1(_1122_),
    .X(_1123_));
 sg13g2_nand3_1 _4851_ (.B(net701),
    .C(_1122_),
    .A(net776),
    .Y(_1124_));
 sg13g2_xor2_1 _4852_ (.B(_0587_),
    .A(_0586_),
    .X(_1125_));
 sg13g2_and3_1 _4853_ (.X(_1126_),
    .A(_1123_),
    .B(_1124_),
    .C(_1125_));
 sg13g2_inv_1 _4854_ (.Y(_1127_),
    .A(_1126_));
 sg13g2_nor3_1 _4855_ (.A(_0618_),
    .B(_0738_),
    .C(_0739_),
    .Y(_1128_));
 sg13g2_o21ai_1 _4856_ (.B1(_0619_),
    .Y(_1129_),
    .A1(_0735_),
    .A2(_0737_));
 sg13g2_nor3_1 _4857_ (.A(_0740_),
    .B(_1127_),
    .C(_1128_),
    .Y(_1130_));
 sg13g2_o21ai_1 _4858_ (.B1(_1124_),
    .Y(_1131_),
    .A1(_0727_),
    .A2(_1121_));
 sg13g2_nand3_1 _4859_ (.B(net697),
    .C(_1131_),
    .A(net783),
    .Y(_1132_));
 sg13g2_a21o_1 _4860_ (.A2(net697),
    .A1(net783),
    .B1(_1131_),
    .X(_1133_));
 sg13g2_or3_1 _4861_ (.A(net728),
    .B(net696),
    .C(_1131_),
    .X(_1134_));
 sg13g2_o21ai_1 _4862_ (.B1(_1131_),
    .Y(_1135_),
    .A1(net728),
    .A2(net696));
 sg13g2_and4_1 _4863_ (.A(net789),
    .B(net695),
    .C(_1132_),
    .D(_1133_),
    .X(_1136_));
 sg13g2_nand4_1 _4864_ (.B(net695),
    .C(_1132_),
    .A(net789),
    .Y(_1137_),
    .D(_1133_));
 sg13g2_a22oi_1 _4865_ (.Y(_1138_),
    .B1(_1132_),
    .B2(_1133_),
    .A2(net695),
    .A1(net789));
 sg13g2_and4_1 _4866_ (.A(net789),
    .B(net695),
    .C(_1134_),
    .D(_1135_),
    .X(_1139_));
 sg13g2_a22oi_1 _4867_ (.Y(_1140_),
    .B1(_1134_),
    .B2(_1135_),
    .A2(net695),
    .A1(net789));
 sg13g2_a21oi_1 _4868_ (.A1(_0741_),
    .A2(_1129_),
    .Y(_1141_),
    .B1(_1126_));
 sg13g2_a21oi_1 _4869_ (.A1(_0741_),
    .A2(_1129_),
    .Y(_1142_),
    .B1(_1127_));
 sg13g2_nor3_1 _4870_ (.A(_0740_),
    .B(_1126_),
    .C(_1128_),
    .Y(_1143_));
 sg13g2_or4_1 _4871_ (.A(_1130_),
    .B(_1136_),
    .C(_1138_),
    .D(_1141_),
    .X(_1144_));
 sg13g2_nand2b_1 _4872_ (.Y(_1145_),
    .B(_1144_),
    .A_N(_1130_));
 sg13g2_or4_1 _4873_ (.A(_0917_),
    .B(_0918_),
    .C(_0920_),
    .D(_0921_),
    .X(_1146_));
 sg13g2_nand3_1 _4874_ (.B(_1145_),
    .C(_1146_),
    .A(_0922_),
    .Y(_1147_));
 sg13g2_nand2_1 _4875_ (.Y(_1148_),
    .A(_1132_),
    .B(_1137_));
 sg13g2_a21o_1 _4876_ (.A2(_1146_),
    .A1(_0922_),
    .B1(_1145_),
    .X(_1149_));
 sg13g2_nand3_1 _4877_ (.B(_1148_),
    .C(_1149_),
    .A(_1147_),
    .Y(_1150_));
 sg13g2_and2_1 _4878_ (.A(_1147_),
    .B(_1150_),
    .X(_1151_));
 sg13g2_a21oi_1 _4879_ (.A1(_1015_),
    .A2(_1019_),
    .Y(_1152_),
    .B1(_1017_));
 sg13g2_o21ai_1 _4880_ (.B1(_1151_),
    .Y(_1153_),
    .A1(_1020_),
    .A2(_1152_));
 sg13g2_nor3_1 _4881_ (.A(_1020_),
    .B(_1151_),
    .C(_1152_),
    .Y(_1154_));
 sg13g2_a21o_1 _4882_ (.A2(_1149_),
    .A1(_1147_),
    .B1(_1148_),
    .X(_1155_));
 sg13g2_a21oi_1 _4883_ (.A1(_1123_),
    .A2(_1124_),
    .Y(_1156_),
    .B1(_1125_));
 sg13g2_or2_1 _4884_ (.X(_1157_),
    .B(_1156_),
    .A(_1126_));
 sg13g2_nand2_2 _4885_ (.Y(_1158_),
    .A(net770),
    .B(_0582_));
 sg13g2_nor2_1 _4886_ (.A(_1121_),
    .B(_1158_),
    .Y(_1159_));
 sg13g2_a22oi_1 _4887_ (.Y(_1160_),
    .B1(net705),
    .B2(net770),
    .A2(_0582_),
    .A1(net767));
 sg13g2_nor2_1 _4888_ (.A(_1159_),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_nand3_1 _4889_ (.B(net703),
    .C(_1161_),
    .A(net777),
    .Y(_1162_));
 sg13g2_a21o_1 _4890_ (.A2(net703),
    .A1(net778),
    .B1(_1161_),
    .X(_1163_));
 sg13g2_and2_1 _4891_ (.A(_1162_),
    .B(_1163_),
    .X(_1165_));
 sg13g2_nor2b_1 _4892_ (.A(_0585_),
    .B_N(_1165_),
    .Y(_1166_));
 sg13g2_nor2b_1 _4893_ (.A(_1157_),
    .B_N(_1166_),
    .Y(_1167_));
 sg13g2_xnor2_1 _4894_ (.Y(_1168_),
    .A(_1157_),
    .B(_1166_));
 sg13g2_nand2_1 _4895_ (.Y(_1169_),
    .A(net790),
    .B(net697));
 sg13g2_o21ai_1 _4896_ (.B1(_1162_),
    .Y(_1170_),
    .A1(_1121_),
    .A2(_1158_));
 sg13g2_nor2_1 _4897_ (.A(net728),
    .B(_0721_),
    .Y(_1171_));
 sg13g2_nand2_1 _4898_ (.Y(_1172_),
    .A(_1170_),
    .B(_1171_));
 sg13g2_xnor2_1 _4899_ (.Y(_1173_),
    .A(_1170_),
    .B(_1171_));
 sg13g2_xor2_1 _4900_ (.B(_1173_),
    .A(_1169_),
    .X(_1174_));
 sg13g2_a21o_1 _4901_ (.A2(_1174_),
    .A1(_1168_),
    .B1(_1167_),
    .X(_1176_));
 sg13g2_or4_1 _4902_ (.A(_1139_),
    .B(_1140_),
    .C(_1142_),
    .D(_1143_),
    .X(_1177_));
 sg13g2_nand3_1 _4903_ (.B(_1176_),
    .C(_1177_),
    .A(_1144_),
    .Y(_1178_));
 sg13g2_o21ai_1 _4904_ (.B1(_1172_),
    .Y(_1179_),
    .A1(_1169_),
    .A2(_1173_));
 sg13g2_inv_1 _4905_ (.Y(_1180_),
    .A(_1179_));
 sg13g2_a21oi_1 _4906_ (.A1(_1144_),
    .A2(_1177_),
    .Y(_1181_),
    .B1(_1176_));
 sg13g2_a21o_1 _4907_ (.A2(_1177_),
    .A1(_1144_),
    .B1(_1176_),
    .X(_1182_));
 sg13g2_and3_1 _4908_ (.X(_1183_),
    .A(_1178_),
    .B(_1179_),
    .C(_1182_));
 sg13g2_o21ai_1 _4909_ (.B1(_1178_),
    .Y(_1184_),
    .A1(_1180_),
    .A2(_1181_));
 sg13g2_nand3_1 _4910_ (.B(_1155_),
    .C(_1184_),
    .A(_1150_),
    .Y(_1185_));
 sg13g2_a21oi_1 _4911_ (.A1(_1150_),
    .A2(_1155_),
    .Y(_1187_),
    .B1(_1184_));
 sg13g2_a21oi_1 _4912_ (.A1(_1178_),
    .A2(_1182_),
    .Y(_1188_),
    .B1(_1179_));
 sg13g2_nand2_1 _4913_ (.Y(_1189_),
    .A(net790),
    .B(net699));
 sg13g2_nand2_1 _4914_ (.Y(_1190_),
    .A(net767),
    .B(_0584_));
 sg13g2_nand2_1 _4915_ (.Y(_1191_),
    .A(net777),
    .B(net705));
 sg13g2_xor2_1 _4916_ (.B(_1190_),
    .A(_1158_),
    .X(_1192_));
 sg13g2_nand3_1 _4917_ (.B(net705),
    .C(_1192_),
    .A(net777),
    .Y(_1193_));
 sg13g2_o21ai_1 _4918_ (.B1(_1193_),
    .Y(_1194_),
    .A1(_1158_),
    .A2(_1190_));
 sg13g2_nand3_1 _4919_ (.B(net701),
    .C(_1194_),
    .A(net784),
    .Y(_1195_));
 sg13g2_a21o_1 _4920_ (.A2(net701),
    .A1(net783),
    .B1(_1194_),
    .X(_1196_));
 sg13g2_nand2_1 _4921_ (.Y(_1198_),
    .A(_1195_),
    .B(_1196_));
 sg13g2_xor2_1 _4922_ (.B(_1198_),
    .A(_1189_),
    .X(_1199_));
 sg13g2_xnor2_1 _4923_ (.Y(_1200_),
    .A(_0585_),
    .B(_1165_));
 sg13g2_nand2_1 _4924_ (.Y(_1201_),
    .A(_1199_),
    .B(_1200_));
 sg13g2_xnor2_1 _4925_ (.Y(_1202_),
    .A(_1168_),
    .B(_1174_));
 sg13g2_nor2_1 _4926_ (.A(_1201_),
    .B(_1202_),
    .Y(_1203_));
 sg13g2_o21ai_1 _4927_ (.B1(_1195_),
    .Y(_1204_),
    .A1(_1189_),
    .A2(_1198_));
 sg13g2_inv_1 _4928_ (.Y(_1205_),
    .A(_1204_));
 sg13g2_nand2_1 _4929_ (.Y(_1206_),
    .A(_1201_),
    .B(_1202_));
 sg13g2_xnor2_1 _4930_ (.Y(_1207_),
    .A(_1201_),
    .B(_1202_));
 sg13g2_a21oi_1 _4931_ (.A1(_1204_),
    .A2(_1206_),
    .Y(_1209_),
    .B1(_1203_));
 sg13g2_o21ai_1 _4932_ (.B1(_1209_),
    .Y(_1210_),
    .A1(_1183_),
    .A2(_1188_));
 sg13g2_nor3_1 _4933_ (.A(_1183_),
    .B(_1188_),
    .C(_1209_),
    .Y(_1211_));
 sg13g2_xor2_1 _4934_ (.B(_1200_),
    .A(_1199_),
    .X(_1212_));
 sg13g2_nand2_1 _4935_ (.Y(_1213_),
    .A(net777),
    .B(_0584_));
 sg13g2_nor2_1 _4936_ (.A(_1158_),
    .B(_1213_),
    .Y(_1214_));
 sg13g2_nand2_1 _4937_ (.Y(_1215_),
    .A(net784),
    .B(net703));
 sg13g2_nand3_1 _4938_ (.B(net703),
    .C(_1214_),
    .A(net783),
    .Y(_1216_));
 sg13g2_xnor2_1 _4939_ (.Y(_1217_),
    .A(_1214_),
    .B(_1215_));
 sg13g2_nand3_1 _4940_ (.B(net701),
    .C(_1217_),
    .A(net790),
    .Y(_1218_));
 sg13g2_a21o_1 _4941_ (.A2(net701),
    .A1(net790),
    .B1(_1217_),
    .X(_1220_));
 sg13g2_nand2_1 _4942_ (.Y(_1221_),
    .A(_1218_),
    .B(_1220_));
 sg13g2_xor2_1 _4943_ (.B(_1192_),
    .A(_1191_),
    .X(_1222_));
 sg13g2_nor2_1 _4944_ (.A(_1221_),
    .B(_1222_),
    .Y(_1223_));
 sg13g2_nand2_1 _4945_ (.Y(_1224_),
    .A(_1212_),
    .B(_1223_));
 sg13g2_and2_1 _4946_ (.A(_1216_),
    .B(_1218_),
    .X(_1225_));
 sg13g2_nand2_1 _4947_ (.Y(_1226_),
    .A(net784),
    .B(_0582_));
 sg13g2_nand2_1 _4948_ (.Y(_1227_),
    .A(net791),
    .B(net705));
 sg13g2_a21oi_1 _4949_ (.A1(_1226_),
    .A2(_1227_),
    .Y(_1228_),
    .B1(_1213_));
 sg13g2_nor2_1 _4950_ (.A(_1226_),
    .B(_1227_),
    .Y(_1229_));
 sg13g2_or2_1 _4951_ (.X(_1231_),
    .B(net705),
    .A(net777));
 sg13g2_nand4_1 _4952_ (.B(net790),
    .C(_0582_),
    .A(net783),
    .Y(_1232_),
    .D(_0584_));
 sg13g2_a21oi_1 _4953_ (.A1(_1191_),
    .A2(_1231_),
    .Y(_1233_),
    .B1(_1232_));
 sg13g2_nor3_1 _4954_ (.A(_1228_),
    .B(_1229_),
    .C(_1233_),
    .Y(_1234_));
 sg13g2_nand2_1 _4955_ (.Y(_1235_),
    .A(_1229_),
    .B(_1233_));
 sg13g2_nand2_1 _4956_ (.Y(_1236_),
    .A(net784),
    .B(_0611_));
 sg13g2_nand2_1 _4957_ (.Y(_1237_),
    .A(net791),
    .B(net704));
 sg13g2_nor2_1 _4958_ (.A(_1215_),
    .B(_1227_),
    .Y(_1238_));
 sg13g2_xor2_1 _4959_ (.B(_1237_),
    .A(_1236_),
    .X(_1239_));
 sg13g2_a22oi_1 _4960_ (.Y(_1240_),
    .B1(_0584_),
    .B2(net770),
    .A2(_0582_),
    .A1(net777));
 sg13g2_nor2_1 _4961_ (.A(_1214_),
    .B(_1240_),
    .Y(_1242_));
 sg13g2_xnor2_1 _4962_ (.Y(_1243_),
    .A(_1239_),
    .B(_1242_));
 sg13g2_a21o_1 _4963_ (.A2(_1243_),
    .A1(_1235_),
    .B1(_1234_),
    .X(_1244_));
 sg13g2_a21oi_1 _4964_ (.A1(_1239_),
    .A2(_1242_),
    .Y(_1245_),
    .B1(_1238_));
 sg13g2_nand2_1 _4965_ (.Y(_1246_),
    .A(_1244_),
    .B(_1245_));
 sg13g2_xor2_1 _4966_ (.B(_1222_),
    .A(_1221_),
    .X(_1247_));
 sg13g2_nor2_1 _4967_ (.A(_1244_),
    .B(_1245_),
    .Y(_1248_));
 sg13g2_o21ai_1 _4968_ (.B1(_1246_),
    .Y(_1249_),
    .A1(_1247_),
    .A2(_1248_));
 sg13g2_or2_1 _4969_ (.X(_1250_),
    .B(_1249_),
    .A(_1225_));
 sg13g2_or2_1 _4970_ (.X(_1251_),
    .B(_1250_),
    .A(_1224_));
 sg13g2_and2_1 _4971_ (.A(_1205_),
    .B(_1207_),
    .X(_1253_));
 sg13g2_and2_1 _4972_ (.A(_1225_),
    .B(_1249_),
    .X(_1254_));
 sg13g2_nor2_1 _4973_ (.A(_1212_),
    .B(_1223_),
    .Y(_1255_));
 sg13g2_a22oi_1 _4974_ (.Y(_1256_),
    .B1(_1255_),
    .B2(_1250_),
    .A2(_1254_),
    .A1(_1224_));
 sg13g2_o21ai_1 _4975_ (.B1(_1256_),
    .Y(_1257_),
    .A1(_1205_),
    .A2(_1207_));
 sg13g2_o21ai_1 _4976_ (.B1(_1251_),
    .Y(_1258_),
    .A1(_1253_),
    .A2(_1257_));
 sg13g2_a21oi_1 _4977_ (.A1(_1210_),
    .A2(_1258_),
    .Y(_1259_),
    .B1(_1211_));
 sg13g2_o21ai_1 _4978_ (.B1(_1185_),
    .Y(_1260_),
    .A1(_1187_),
    .A2(_1259_));
 sg13g2_a21oi_2 _4979_ (.B1(_1154_),
    .Y(_1261_),
    .A2(_1260_),
    .A1(_1153_));
 sg13g2_xnor2_1 _4980_ (.Y(_1262_),
    .A(_1120_),
    .B(_1261_));
 sg13g2_nand2_1 _4981_ (.Y(_1264_),
    .A(_1472_),
    .B(net691));
 sg13g2_nor2_2 _4982_ (.A(_0019_),
    .B(_0906_),
    .Y(_1265_));
 sg13g2_nand2_1 _4983_ (.Y(_1266_),
    .A(net763),
    .B(net691));
 sg13g2_inv_1 _4984_ (.Y(_1267_),
    .A(_1266_));
 sg13g2_nand2_1 _4985_ (.Y(_1268_),
    .A(net766),
    .B(net687));
 sg13g2_xor2_1 _4986_ (.B(_1266_),
    .A(_1265_),
    .X(_1269_));
 sg13g2_nor2_1 _4987_ (.A(_1268_),
    .B(_1269_),
    .Y(_1270_));
 sg13g2_a21oi_2 _4988_ (.B1(_1270_),
    .Y(_1271_),
    .A2(_1267_),
    .A1(_1265_));
 sg13g2_o21ai_1 _4989_ (.B1(_1096_),
    .Y(_1272_),
    .A1(_1057_),
    .A2(_1097_));
 sg13g2_o21ai_1 _4990_ (.B1(_1093_),
    .Y(_1273_),
    .A1(_1058_),
    .A2(_1094_));
 sg13g2_o21ai_1 _4991_ (.B1(_1090_),
    .Y(_1275_),
    .A1(_1061_),
    .A2(_1091_));
 sg13g2_nand2_1 _4992_ (.Y(_1276_),
    .A(_1084_),
    .B(_1086_));
 sg13g2_inv_1 _4993_ (.Y(_1277_),
    .A(_1276_));
 sg13g2_o21ai_1 _4994_ (.B1(_1079_),
    .Y(_1278_),
    .A1(_1080_),
    .A2(_1088_));
 sg13g2_nand2_1 _4995_ (.Y(_1279_),
    .A(net760),
    .B(net800));
 sg13g2_o21ai_1 _4996_ (.B1(_1075_),
    .Y(_1280_),
    .A1(_0941_),
    .A2(_1073_));
 sg13g2_nand2_1 _4997_ (.Y(_1281_),
    .A(net758),
    .B(net804));
 sg13g2_nand2b_1 _4998_ (.Y(_1282_),
    .B(_1280_),
    .A_N(_1281_));
 sg13g2_xnor2_1 _4999_ (.Y(_1283_),
    .A(_1280_),
    .B(_1281_));
 sg13g2_nand2b_1 _5000_ (.Y(_1284_),
    .B(_1283_),
    .A_N(_1279_));
 sg13g2_xnor2_1 _5001_ (.Y(_1286_),
    .A(_1279_),
    .B(_1283_));
 sg13g2_inv_1 _5002_ (.Y(_1287_),
    .A(_1286_));
 sg13g2_a21o_1 _5003_ (.A2(_1070_),
    .A1(_1064_),
    .B1(_1077_),
    .X(_1288_));
 sg13g2_nand2_1 _5004_ (.Y(_1289_),
    .A(net755),
    .B(net807));
 sg13g2_nand2_2 _5005_ (.Y(_1290_),
    .A(\system_inst.internal_param_b[4] ),
    .B(net809));
 sg13g2_nor2_1 _5006_ (.A(_1073_),
    .B(_1290_),
    .Y(_1291_));
 sg13g2_or2_1 _5007_ (.X(_1292_),
    .B(_1290_),
    .A(_1073_));
 sg13g2_a22oi_1 _5008_ (.Y(_1293_),
    .B1(net813),
    .B2(net750),
    .A2(net809),
    .A1(net753));
 sg13g2_nor2_1 _5009_ (.A(_1291_),
    .B(_1293_),
    .Y(_1294_));
 sg13g2_xnor2_1 _5010_ (.Y(_1295_),
    .A(_1289_),
    .B(_1294_));
 sg13g2_inv_1 _5011_ (.Y(_1297_),
    .A(_1295_));
 sg13g2_o21ai_1 _5012_ (.B1(_1069_),
    .Y(_1298_),
    .A1(_0934_),
    .A2(_1067_));
 sg13g2_nand2_1 _5013_ (.Y(_1299_),
    .A(net747),
    .B(net817));
 sg13g2_nand2_1 _5014_ (.Y(_1300_),
    .A(net744),
    .B(net822));
 sg13g2_nand2_1 _5015_ (.Y(_1301_),
    .A(net745),
    .B(net822));
 sg13g2_xor2_1 _5016_ (.B(_1301_),
    .A(_1066_),
    .X(_1302_));
 sg13g2_nand2b_1 _5017_ (.Y(_1303_),
    .B(_1302_),
    .A_N(_1299_));
 sg13g2_xnor2_1 _5018_ (.Y(_1304_),
    .A(_1299_),
    .B(_1302_));
 sg13g2_nand2_1 _5019_ (.Y(_1305_),
    .A(_1298_),
    .B(_1304_));
 sg13g2_xnor2_1 _5020_ (.Y(_1306_),
    .A(_1298_),
    .B(_1304_));
 sg13g2_xnor2_1 _5021_ (.Y(_1308_),
    .A(_1295_),
    .B(_1306_));
 sg13g2_nand2_1 _5022_ (.Y(_1309_),
    .A(_1288_),
    .B(_1308_));
 sg13g2_xnor2_1 _5023_ (.Y(_1310_),
    .A(_1288_),
    .B(_1308_));
 sg13g2_xnor2_1 _5024_ (.Y(_1311_),
    .A(_1287_),
    .B(_1310_));
 sg13g2_nand2b_1 _5025_ (.Y(_1312_),
    .B(_1278_),
    .A_N(_1311_));
 sg13g2_xor2_1 _5026_ (.B(_1311_),
    .A(_1278_),
    .X(_1313_));
 sg13g2_xnor2_1 _5027_ (.Y(_1314_),
    .A(_1277_),
    .B(_1313_));
 sg13g2_nor2b_1 _5028_ (.A(_1314_),
    .B_N(_1275_),
    .Y(_1315_));
 sg13g2_xor2_1 _5029_ (.B(_1314_),
    .A(_1275_),
    .X(_1316_));
 sg13g2_inv_1 _5030_ (.Y(_1317_),
    .A(_1316_));
 sg13g2_xnor2_1 _5031_ (.Y(_1319_),
    .A(_1273_),
    .B(_1317_));
 sg13g2_xnor2_1 _5032_ (.Y(_1320_),
    .A(_0011_),
    .B(_1319_));
 sg13g2_xor2_1 _5033_ (.B(_1320_),
    .A(_1272_),
    .X(_1321_));
 sg13g2_xnor2_1 _5034_ (.Y(_1322_),
    .A(_1272_),
    .B(_1320_));
 sg13g2_nand2_1 _5035_ (.Y(_1323_),
    .A(net766),
    .B(_1321_));
 sg13g2_nor2_1 _5036_ (.A(_0019_),
    .B(_1099_),
    .Y(_1324_));
 sg13g2_nand2_1 _5037_ (.Y(_1325_),
    .A(net763),
    .B(net687));
 sg13g2_xnor2_1 _5038_ (.Y(_1326_),
    .A(_1264_),
    .B(_1325_));
 sg13g2_nor2_1 _5039_ (.A(_1323_),
    .B(_1326_),
    .Y(_1327_));
 sg13g2_xor2_1 _5040_ (.B(_1326_),
    .A(_1323_),
    .X(_1328_));
 sg13g2_nor2b_1 _5041_ (.A(_1271_),
    .B_N(_1328_),
    .Y(_1330_));
 sg13g2_a21oi_2 _5042_ (.B1(_1315_),
    .Y(_1331_),
    .A2(_1317_),
    .A1(_1273_));
 sg13g2_o21ai_1 _5043_ (.B1(_1312_),
    .Y(_1332_),
    .A1(_1277_),
    .A2(_1313_));
 sg13g2_nand2_1 _5044_ (.Y(_1333_),
    .A(_1282_),
    .B(_1284_));
 sg13g2_inv_1 _5045_ (.Y(_1334_),
    .A(_1333_));
 sg13g2_o21ai_1 _5046_ (.B1(_1309_),
    .Y(_1335_),
    .A1(_1287_),
    .A2(_1310_));
 sg13g2_o21ai_1 _5047_ (.B1(_1292_),
    .Y(_1336_),
    .A1(_1289_),
    .A2(_1293_));
 sg13g2_nand2_1 _5048_ (.Y(_1337_),
    .A(net758),
    .B(net800));
 sg13g2_nand2b_1 _5049_ (.Y(_1338_),
    .B(_1336_),
    .A_N(_1337_));
 sg13g2_xnor2_1 _5050_ (.Y(_1339_),
    .A(_1336_),
    .B(_1337_));
 sg13g2_inv_1 _5051_ (.Y(_1341_),
    .A(_1339_));
 sg13g2_o21ai_1 _5052_ (.B1(_1305_),
    .Y(_1342_),
    .A1(_1297_),
    .A2(_1306_));
 sg13g2_o21ai_1 _5053_ (.B1(_1303_),
    .Y(_1343_),
    .A1(_1066_),
    .A2(_1301_));
 sg13g2_nand2_1 _5054_ (.Y(_1344_),
    .A(net748),
    .B(net813));
 sg13g2_nand2_1 _5055_ (.Y(_1345_),
    .A(net743),
    .B(net817));
 sg13g2_nand2_1 _5056_ (.Y(_1346_),
    .A(net746),
    .B(net817));
 sg13g2_xor2_1 _5057_ (.B(_1346_),
    .A(_1300_),
    .X(_1347_));
 sg13g2_nand2b_1 _5058_ (.Y(_1348_),
    .B(_1347_),
    .A_N(_1344_));
 sg13g2_xnor2_1 _5059_ (.Y(_1349_),
    .A(_1344_),
    .B(_1347_));
 sg13g2_xnor2_1 _5060_ (.Y(_1350_),
    .A(_1343_),
    .B(_1349_));
 sg13g2_nand2_1 _5061_ (.Y(_1352_),
    .A(net755),
    .B(net804));
 sg13g2_nand2_1 _5062_ (.Y(_1353_),
    .A(net750),
    .B(net807));
 sg13g2_nand2_1 _5063_ (.Y(_1354_),
    .A(net753),
    .B(net807));
 sg13g2_xor2_1 _5064_ (.B(_1354_),
    .A(_1290_),
    .X(_1355_));
 sg13g2_nand2b_1 _5065_ (.Y(_1356_),
    .B(_1355_),
    .A_N(_1352_));
 sg13g2_xnor2_1 _5066_ (.Y(_1357_),
    .A(_1352_),
    .B(_1355_));
 sg13g2_nor2b_1 _5067_ (.A(_1350_),
    .B_N(_1357_),
    .Y(_1358_));
 sg13g2_xnor2_1 _5068_ (.Y(_1359_),
    .A(_1350_),
    .B(_1357_));
 sg13g2_nand2_1 _5069_ (.Y(_1360_),
    .A(_1342_),
    .B(_1359_));
 sg13g2_xnor2_1 _5070_ (.Y(_1361_),
    .A(_1342_),
    .B(_1359_));
 sg13g2_xnor2_1 _5071_ (.Y(_1363_),
    .A(_1339_),
    .B(_1361_));
 sg13g2_nand2_1 _5072_ (.Y(_1364_),
    .A(_1335_),
    .B(_1363_));
 sg13g2_xnor2_1 _5073_ (.Y(_1365_),
    .A(_1335_),
    .B(_1363_));
 sg13g2_xnor2_1 _5074_ (.Y(_1366_),
    .A(_1334_),
    .B(_1365_));
 sg13g2_nand2b_1 _5075_ (.Y(_1367_),
    .B(_1332_),
    .A_N(_1366_));
 sg13g2_xor2_1 _5076_ (.B(_1366_),
    .A(_1332_),
    .X(_1368_));
 sg13g2_xor2_1 _5077_ (.B(_1368_),
    .A(_1331_),
    .X(_1369_));
 sg13g2_nand2_1 _5078_ (.Y(_1370_),
    .A(_0010_),
    .B(_1369_));
 sg13g2_nor2_1 _5079_ (.A(\system_inst.neuron.u[8] ),
    .B(_1319_),
    .Y(_1371_));
 sg13g2_a21oi_2 _5080_ (.B1(_1371_),
    .Y(_1372_),
    .A2(_1320_),
    .A1(_1272_));
 sg13g2_xnor2_1 _5081_ (.Y(_1374_),
    .A(_0010_),
    .B(_1369_));
 sg13g2_o21ai_1 _5082_ (.B1(_1370_),
    .Y(_1375_),
    .A1(_1372_),
    .A2(_1374_));
 sg13g2_o21ai_1 _5083_ (.B1(_1367_),
    .Y(_1376_),
    .A1(_1331_),
    .A2(_1368_));
 sg13g2_o21ai_1 _5084_ (.B1(_1364_),
    .Y(_1377_),
    .A1(_1334_),
    .A2(_1365_));
 sg13g2_o21ai_1 _5085_ (.B1(_1360_),
    .Y(_1378_),
    .A1(_1341_),
    .A2(_1361_));
 sg13g2_o21ai_1 _5086_ (.B1(_1356_),
    .Y(_1379_),
    .A1(_1290_),
    .A2(_1354_));
 sg13g2_inv_1 _5087_ (.Y(_1380_),
    .A(_1379_));
 sg13g2_a21o_1 _5088_ (.A2(_1349_),
    .A1(_1343_),
    .B1(_1358_),
    .X(_1381_));
 sg13g2_o21ai_1 _5089_ (.B1(_1348_),
    .Y(_1382_),
    .A1(_1300_),
    .A2(_1346_));
 sg13g2_nand2_1 _5090_ (.Y(_1383_),
    .A(net748),
    .B(net809));
 sg13g2_nand2_1 _5091_ (.Y(_1385_),
    .A(net743),
    .B(net813));
 sg13g2_nand2_1 _5092_ (.Y(_1386_),
    .A(net746),
    .B(net813));
 sg13g2_xor2_1 _5093_ (.B(_1386_),
    .A(_1345_),
    .X(_1387_));
 sg13g2_nand2b_1 _5094_ (.Y(_1388_),
    .B(_1387_),
    .A_N(_1383_));
 sg13g2_xnor2_1 _5095_ (.Y(_1389_),
    .A(_1383_),
    .B(_1387_));
 sg13g2_xnor2_1 _5096_ (.Y(_1390_),
    .A(_1382_),
    .B(_1389_));
 sg13g2_nand2_1 _5097_ (.Y(_1391_),
    .A(net755),
    .B(net800));
 sg13g2_nand2_1 _5098_ (.Y(_1392_),
    .A(net753),
    .B(net804));
 sg13g2_xor2_1 _5099_ (.B(_1392_),
    .A(_1353_),
    .X(_1393_));
 sg13g2_nand2b_1 _5100_ (.Y(_1394_),
    .B(_1393_),
    .A_N(_1391_));
 sg13g2_xnor2_1 _5101_ (.Y(_1396_),
    .A(_1391_),
    .B(_1393_));
 sg13g2_nor2b_1 _5102_ (.A(_1390_),
    .B_N(_1396_),
    .Y(_1397_));
 sg13g2_xnor2_1 _5103_ (.Y(_1398_),
    .A(_1390_),
    .B(_1396_));
 sg13g2_nand2_1 _5104_ (.Y(_1399_),
    .A(_1381_),
    .B(_1398_));
 sg13g2_xnor2_1 _5105_ (.Y(_1400_),
    .A(_1381_),
    .B(_1398_));
 sg13g2_xnor2_1 _5106_ (.Y(_1401_),
    .A(_1380_),
    .B(_1400_));
 sg13g2_nand2b_1 _5107_ (.Y(_1402_),
    .B(_1378_),
    .A_N(_1401_));
 sg13g2_xor2_1 _5108_ (.B(_1401_),
    .A(_1378_),
    .X(_1403_));
 sg13g2_xor2_1 _5109_ (.B(_1403_),
    .A(_1338_),
    .X(_1404_));
 sg13g2_and2_1 _5110_ (.A(_1377_),
    .B(_1404_),
    .X(_1405_));
 sg13g2_xnor2_1 _5111_ (.Y(_1407_),
    .A(_1377_),
    .B(_1404_));
 sg13g2_inv_1 _5112_ (.Y(_1408_),
    .A(_1407_));
 sg13g2_xnor2_1 _5113_ (.Y(_1409_),
    .A(_1376_),
    .B(_1408_));
 sg13g2_xnor2_1 _5114_ (.Y(_1410_),
    .A(_0009_),
    .B(_1409_));
 sg13g2_nor2_1 _5115_ (.A(\system_inst.neuron.u[10] ),
    .B(_1409_),
    .Y(_1411_));
 sg13g2_a21oi_2 _5116_ (.B1(_1411_),
    .Y(_1412_),
    .A2(_1410_),
    .A1(_1375_));
 sg13g2_o21ai_1 _5117_ (.B1(_1399_),
    .Y(_1413_),
    .A1(_1380_),
    .A2(_1400_));
 sg13g2_o21ai_1 _5118_ (.B1(_1394_),
    .Y(_1414_),
    .A1(_1353_),
    .A2(_1392_));
 sg13g2_a21o_1 _5119_ (.A2(_1389_),
    .A1(_1382_),
    .B1(_1397_),
    .X(_1415_));
 sg13g2_a22oi_1 _5120_ (.Y(_1416_),
    .B1(net804),
    .B2(net750),
    .A2(net800),
    .A1(net753));
 sg13g2_nand2_1 _5121_ (.Y(_1418_),
    .A(net750),
    .B(net800));
 sg13g2_or2_1 _5122_ (.X(_1419_),
    .B(_1418_),
    .A(_1392_));
 sg13g2_nand2b_1 _5123_ (.Y(_1420_),
    .B(_1419_),
    .A_N(_1416_));
 sg13g2_o21ai_1 _5124_ (.B1(_1388_),
    .Y(_1421_),
    .A1(_1345_),
    .A2(_1386_));
 sg13g2_nand2_1 _5125_ (.Y(_1422_),
    .A(net748),
    .B(net807));
 sg13g2_nand2_1 _5126_ (.Y(_1423_),
    .A(net746),
    .B(net809));
 sg13g2_or2_1 _5127_ (.X(_1424_),
    .B(_1423_),
    .A(_1385_));
 sg13g2_xnor2_1 _5128_ (.Y(_1425_),
    .A(_1385_),
    .B(_1423_));
 sg13g2_xor2_1 _5129_ (.B(_1425_),
    .A(_1422_),
    .X(_1426_));
 sg13g2_nand2_1 _5130_ (.Y(_1427_),
    .A(_1421_),
    .B(_1426_));
 sg13g2_xnor2_1 _5131_ (.Y(_1429_),
    .A(_1421_),
    .B(_1426_));
 sg13g2_xnor2_1 _5132_ (.Y(_1430_),
    .A(_1420_),
    .B(_1429_));
 sg13g2_nor2b_1 _5133_ (.A(_1430_),
    .B_N(_1415_),
    .Y(_1431_));
 sg13g2_xor2_1 _5134_ (.B(_1430_),
    .A(_1415_),
    .X(_1432_));
 sg13g2_nor2b_1 _5135_ (.A(_1432_),
    .B_N(_1414_),
    .Y(_1433_));
 sg13g2_xnor2_1 _5136_ (.Y(_1434_),
    .A(_1414_),
    .B(_1432_));
 sg13g2_nand2_1 _5137_ (.Y(_1435_),
    .A(_1413_),
    .B(_1434_));
 sg13g2_xnor2_1 _5138_ (.Y(_1436_),
    .A(_1413_),
    .B(_1434_));
 sg13g2_o21ai_1 _5139_ (.B1(_1402_),
    .Y(_1437_),
    .A1(_1338_),
    .A2(_1403_));
 sg13g2_nand2b_1 _5140_ (.Y(_1438_),
    .B(_1437_),
    .A_N(_1436_));
 sg13g2_xor2_1 _5141_ (.B(_1437_),
    .A(_1436_),
    .X(_1440_));
 sg13g2_a21oi_1 _5142_ (.A1(_1376_),
    .A2(_1408_),
    .Y(_1441_),
    .B1(_1405_));
 sg13g2_xor2_1 _5143_ (.B(_1441_),
    .A(_1440_),
    .X(_1442_));
 sg13g2_nand2_1 _5144_ (.Y(_1443_),
    .A(_0008_),
    .B(_1442_));
 sg13g2_xnor2_1 _5145_ (.Y(_1444_),
    .A(_0008_),
    .B(_1442_));
 sg13g2_xor2_1 _5146_ (.B(_1444_),
    .A(_1412_),
    .X(_1445_));
 sg13g2_xnor2_1 _5147_ (.Y(_1446_),
    .A(_1412_),
    .B(_1444_));
 sg13g2_xor2_1 _5148_ (.B(_1374_),
    .A(_1372_),
    .X(_1447_));
 sg13g2_xnor2_1 _5149_ (.Y(_1448_),
    .A(_1372_),
    .B(_1374_));
 sg13g2_xor2_1 _5150_ (.B(_1410_),
    .A(_1375_),
    .X(_1449_));
 sg13g2_xnor2_1 _5151_ (.Y(_1451_),
    .A(_1375_),
    .B(_1410_));
 sg13g2_nor2_1 _5152_ (.A(net741),
    .B(_1451_),
    .Y(_1452_));
 sg13g2_nand2_2 _5153_ (.Y(_1453_),
    .A(net769),
    .B(net677));
 sg13g2_nor2_1 _5154_ (.A(net741),
    .B(net678),
    .Y(_1454_));
 sg13g2_nor3_1 _5155_ (.A(net738),
    .B(net678),
    .C(_1453_),
    .Y(_1455_));
 sg13g2_nand3_1 _5156_ (.B(net677),
    .C(_1454_),
    .A(net775),
    .Y(_1456_));
 sg13g2_a21o_1 _5157_ (.A2(net677),
    .A1(net774),
    .B1(_1454_),
    .X(_1457_));
 sg13g2_and4_1 _5158_ (.A(net781),
    .B(net675),
    .C(_1456_),
    .D(_1457_),
    .X(_1458_));
 sg13g2_a22oi_1 _5159_ (.Y(_1459_),
    .B1(_1456_),
    .B2(_1457_),
    .A2(net675),
    .A1(net781));
 sg13g2_nor2_1 _5160_ (.A(_1458_),
    .B(_1459_),
    .Y(_1460_));
 sg13g2_xnor2_1 _5161_ (.Y(_1462_),
    .A(_1271_),
    .B(_1328_));
 sg13g2_a21oi_1 _5162_ (.A1(_1460_),
    .A2(_1462_),
    .Y(_1463_),
    .B1(_1330_));
 sg13g2_a21o_1 _5163_ (.A2(_1462_),
    .A1(_1460_),
    .B1(_1330_),
    .X(_1464_));
 sg13g2_o21ai_1 _5164_ (.B1(_1443_),
    .Y(_1465_),
    .A1(_1412_),
    .A2(_1444_));
 sg13g2_o21ai_1 _5165_ (.B1(_1427_),
    .Y(_1466_),
    .A1(_1420_),
    .A2(_1429_));
 sg13g2_o21ai_1 _5166_ (.B1(_1424_),
    .Y(_1467_),
    .A1(_1422_),
    .A2(_1425_));
 sg13g2_nand2_1 _5167_ (.Y(_1468_),
    .A(net748),
    .B(net804));
 sg13g2_nand2_1 _5168_ (.Y(_1469_),
    .A(net743),
    .B(net807));
 sg13g2_nor2_1 _5169_ (.A(_1423_),
    .B(_1469_),
    .Y(_1470_));
 sg13g2_a22oi_1 _5170_ (.Y(_1471_),
    .B1(net809),
    .B2(net743),
    .A2(net807),
    .A1(net746));
 sg13g2_nor2_1 _5171_ (.A(_1470_),
    .B(_1471_),
    .Y(_1473_));
 sg13g2_nor3_1 _5172_ (.A(_1468_),
    .B(_1470_),
    .C(_1471_),
    .Y(_1474_));
 sg13g2_xnor2_1 _5173_ (.Y(_1475_),
    .A(_1468_),
    .B(_1473_));
 sg13g2_xnor2_1 _5174_ (.Y(_1476_),
    .A(_1467_),
    .B(_1475_));
 sg13g2_nor2_1 _5175_ (.A(_1418_),
    .B(_1476_),
    .Y(_1477_));
 sg13g2_xor2_1 _5176_ (.B(_1476_),
    .A(_1418_),
    .X(_1478_));
 sg13g2_nand2_1 _5177_ (.Y(_1479_),
    .A(_1466_),
    .B(_1478_));
 sg13g2_xnor2_1 _5178_ (.Y(_1480_),
    .A(_1466_),
    .B(_1478_));
 sg13g2_xor2_1 _5179_ (.B(_1480_),
    .A(_1419_),
    .X(_1481_));
 sg13g2_o21ai_1 _5180_ (.B1(_1481_),
    .Y(_1482_),
    .A1(_1431_),
    .A2(_1433_));
 sg13g2_or3_1 _5181_ (.A(_1431_),
    .B(_1433_),
    .C(_1481_),
    .X(_1484_));
 sg13g2_nand2_1 _5182_ (.Y(_1485_),
    .A(_1482_),
    .B(_1484_));
 sg13g2_nor2_1 _5183_ (.A(_1435_),
    .B(_1485_),
    .Y(_1486_));
 sg13g2_xor2_1 _5184_ (.B(_1485_),
    .A(_1435_),
    .X(_1487_));
 sg13g2_o21ai_1 _5185_ (.B1(_1438_),
    .Y(_1488_),
    .A1(_1440_),
    .A2(_1441_));
 sg13g2_xor2_1 _5186_ (.B(_1488_),
    .A(_1487_),
    .X(_1489_));
 sg13g2_xnor2_1 _5187_ (.Y(_1490_),
    .A(_1483_),
    .B(_1489_));
 sg13g2_xor2_1 _5188_ (.B(_1490_),
    .A(_1465_),
    .X(_1491_));
 sg13g2_xnor2_1 _5189_ (.Y(_1492_),
    .A(_1465_),
    .B(_1490_));
 sg13g2_nor3_1 _5190_ (.A(net738),
    .B(_1446_),
    .C(_1453_),
    .Y(_1493_));
 sg13g2_nand3_1 _5191_ (.B(net675),
    .C(_1452_),
    .A(net774),
    .Y(_1495_));
 sg13g2_o21ai_1 _5192_ (.B1(_1453_),
    .Y(_1496_),
    .A1(net738),
    .A2(_1446_));
 sg13g2_nand3_1 _5193_ (.B(net675),
    .C(_1453_),
    .A(net774),
    .Y(_1497_));
 sg13g2_o21ai_1 _5194_ (.B1(_1452_),
    .Y(_1498_),
    .A1(net738),
    .A2(_1446_));
 sg13g2_and4_1 _5195_ (.A(net782),
    .B(_1491_),
    .C(_1495_),
    .D(_1496_),
    .X(_1499_));
 sg13g2_a22oi_1 _5196_ (.Y(_1500_),
    .B1(_1495_),
    .B2(_1496_),
    .A2(net673),
    .A1(net782));
 sg13g2_and4_1 _5197_ (.A(net782),
    .B(net673),
    .C(_1497_),
    .D(_1498_),
    .X(_1501_));
 sg13g2_a22oi_1 _5198_ (.Y(_1502_),
    .B1(_1497_),
    .B2(_1498_),
    .A2(net673),
    .A1(net782));
 sg13g2_a21oi_2 _5199_ (.B1(_1327_),
    .Y(_1503_),
    .A2(_1324_),
    .A1(_1267_));
 sg13g2_inv_1 _5200_ (.Y(_1504_),
    .A(_1503_));
 sg13g2_nand2_1 _5201_ (.Y(_1506_),
    .A(net766),
    .B(net680));
 sg13g2_nor2_1 _5202_ (.A(_0019_),
    .B(_1322_),
    .Y(_1507_));
 sg13g2_nor3_1 _5203_ (.A(_0019_),
    .B(_1322_),
    .C(_1325_),
    .Y(_1508_));
 sg13g2_a21oi_1 _5204_ (.A1(net763),
    .A2(net684),
    .Y(_1509_),
    .B1(_1324_));
 sg13g2_or2_1 _5205_ (.X(_1510_),
    .B(_1509_),
    .A(_1508_));
 sg13g2_nor2_1 _5206_ (.A(_1506_),
    .B(_1510_),
    .Y(_1511_));
 sg13g2_xor2_1 _5207_ (.B(_1510_),
    .A(_1506_),
    .X(_1512_));
 sg13g2_xor2_1 _5208_ (.B(_1512_),
    .A(_1503_),
    .X(_1513_));
 sg13g2_inv_1 _5209_ (.Y(_1514_),
    .A(_1513_));
 sg13g2_nor3_2 _5210_ (.A(_1499_),
    .B(_1500_),
    .C(_1513_),
    .Y(_1515_));
 sg13g2_o21ai_1 _5211_ (.B1(_1514_),
    .Y(_1517_),
    .A1(_1501_),
    .A2(_1502_));
 sg13g2_nor3_1 _5212_ (.A(_1501_),
    .B(_1502_),
    .C(_1514_),
    .Y(_1518_));
 sg13g2_o21ai_1 _5213_ (.B1(_1513_),
    .Y(_1519_),
    .A1(_1499_),
    .A2(_1500_));
 sg13g2_nor3_1 _5214_ (.A(_1463_),
    .B(_1515_),
    .C(_1518_),
    .Y(_1520_));
 sg13g2_a21oi_1 _5215_ (.A1(_1487_),
    .A2(_1488_),
    .Y(_1521_),
    .B1(_1486_));
 sg13g2_o21ai_1 _5216_ (.B1(_1479_),
    .Y(_1522_),
    .A1(_1419_),
    .A2(_1480_));
 sg13g2_nand2_1 _5217_ (.Y(_1523_),
    .A(net748),
    .B(net800));
 sg13g2_nand2_1 _5218_ (.Y(_1524_),
    .A(net743),
    .B(net804));
 sg13g2_nand2_1 _5219_ (.Y(_1525_),
    .A(net746),
    .B(net804));
 sg13g2_xor2_1 _5220_ (.B(_1525_),
    .A(_1469_),
    .X(_1526_));
 sg13g2_nand2b_1 _5221_ (.Y(_1528_),
    .B(_1526_),
    .A_N(_1523_));
 sg13g2_xnor2_1 _5222_ (.Y(_1529_),
    .A(_1523_),
    .B(_1526_));
 sg13g2_nor3_1 _5223_ (.A(_1470_),
    .B(_1474_),
    .C(_1529_),
    .Y(_1530_));
 sg13g2_o21ai_1 _5224_ (.B1(_1529_),
    .Y(_1531_),
    .A1(_1470_),
    .A2(_1474_));
 sg13g2_nor2b_1 _5225_ (.A(_1530_),
    .B_N(_1531_),
    .Y(_1532_));
 sg13g2_a21oi_1 _5226_ (.A1(_1467_),
    .A2(_1475_),
    .Y(_1533_),
    .B1(_1477_));
 sg13g2_xnor2_1 _5227_ (.Y(_1534_),
    .A(_1532_),
    .B(_1533_));
 sg13g2_nand2_1 _5228_ (.Y(_1535_),
    .A(_1522_),
    .B(_1534_));
 sg13g2_xnor2_1 _5229_ (.Y(_1536_),
    .A(_1522_),
    .B(_1534_));
 sg13g2_or2_1 _5230_ (.X(_1537_),
    .B(_1536_),
    .A(_1482_));
 sg13g2_xor2_1 _5231_ (.B(_1536_),
    .A(_1482_),
    .X(_1539_));
 sg13g2_inv_1 _5232_ (.Y(_1540_),
    .A(_1539_));
 sg13g2_xnor2_1 _5233_ (.Y(_1541_),
    .A(_1521_),
    .B(_1539_));
 sg13g2_nand2_1 _5234_ (.Y(_1542_),
    .A(_0034_),
    .B(_1541_));
 sg13g2_a22oi_1 _5235_ (.Y(_1543_),
    .B1(_1490_),
    .B2(_1465_),
    .A2(_1489_),
    .A1(_1164_));
 sg13g2_xnor2_1 _5236_ (.Y(_1544_),
    .A(_0034_),
    .B(_1541_));
 sg13g2_o21ai_1 _5237_ (.B1(_1542_),
    .Y(_1545_),
    .A1(_1543_),
    .A2(_1544_));
 sg13g2_o21ai_1 _5238_ (.B1(_1537_),
    .Y(_1546_),
    .A1(_1521_),
    .A2(_1540_));
 sg13g2_a21oi_1 _5239_ (.A1(_1531_),
    .A2(_1533_),
    .Y(_1547_),
    .B1(_1530_));
 sg13g2_o21ai_1 _5240_ (.B1(_1528_),
    .Y(_1548_),
    .A1(_1469_),
    .A2(_1525_));
 sg13g2_nand2_1 _5241_ (.Y(_1550_),
    .A(net746),
    .B(net800));
 sg13g2_xnor2_1 _5242_ (.Y(_1551_),
    .A(_1524_),
    .B(_1550_));
 sg13g2_xnor2_1 _5243_ (.Y(_1552_),
    .A(_1548_),
    .B(_1551_));
 sg13g2_xnor2_1 _5244_ (.Y(_1553_),
    .A(_1547_),
    .B(_1552_));
 sg13g2_xnor2_1 _5245_ (.Y(_1554_),
    .A(_1535_),
    .B(_1553_));
 sg13g2_xor2_1 _5246_ (.B(_1554_),
    .A(_1546_),
    .X(_1555_));
 sg13g2_nor2_1 _5247_ (.A(net742),
    .B(_1555_),
    .Y(_1556_));
 sg13g2_xor2_1 _5248_ (.B(_1555_),
    .A(net742),
    .X(_1557_));
 sg13g2_nand2_1 _5249_ (.Y(_1558_),
    .A(_1545_),
    .B(_1557_));
 sg13g2_xor2_1 _5250_ (.B(_1557_),
    .A(_1545_),
    .X(_1559_));
 sg13g2_nor2_1 _5251_ (.A(_1455_),
    .B(_1458_),
    .Y(_1561_));
 sg13g2_or2_1 _5252_ (.X(_1562_),
    .B(_1458_),
    .A(_1455_));
 sg13g2_xor2_1 _5253_ (.B(_1544_),
    .A(_1543_),
    .X(_1563_));
 sg13g2_nand3_1 _5254_ (.B(_1562_),
    .C(_1563_),
    .A(net786),
    .Y(_1564_));
 sg13g2_a21o_1 _5255_ (.A2(_1563_),
    .A1(net786),
    .B1(_1562_),
    .X(_1565_));
 sg13g2_nand3_1 _5256_ (.B(_1561_),
    .C(_1563_),
    .A(net786),
    .Y(_1566_));
 sg13g2_a21o_1 _5257_ (.A2(_1563_),
    .A1(net786),
    .B1(_1561_),
    .X(_1567_));
 sg13g2_and4_1 _5258_ (.A(net795),
    .B(_1559_),
    .C(_1564_),
    .D(_1565_),
    .X(_1568_));
 sg13g2_nand4_1 _5259_ (.B(_1559_),
    .C(_1564_),
    .A(net795),
    .Y(_1569_),
    .D(_1565_));
 sg13g2_a22oi_1 _5260_ (.Y(_1570_),
    .B1(_1564_),
    .B2(_1565_),
    .A2(_1559_),
    .A1(net795));
 sg13g2_and4_1 _5261_ (.A(net795),
    .B(_1559_),
    .C(_1566_),
    .D(_1567_),
    .X(_1572_));
 sg13g2_a22oi_1 _5262_ (.Y(_1573_),
    .B1(_1566_),
    .B2(_1567_),
    .A2(_1559_),
    .A1(net795));
 sg13g2_a21oi_1 _5263_ (.A1(_1517_),
    .A2(_1519_),
    .Y(_1574_),
    .B1(_1464_));
 sg13g2_a21oi_1 _5264_ (.A1(_1517_),
    .A2(_1519_),
    .Y(_1575_),
    .B1(_1463_));
 sg13g2_nor3_1 _5265_ (.A(_1464_),
    .B(_1515_),
    .C(_1518_),
    .Y(_1576_));
 sg13g2_or4_1 _5266_ (.A(_1520_),
    .B(_1568_),
    .C(_1570_),
    .D(_1574_),
    .X(_1577_));
 sg13g2_nand2b_1 _5267_ (.Y(_1578_),
    .B(_1577_),
    .A_N(_1520_));
 sg13g2_xnor2_1 _5268_ (.Y(_1579_),
    .A(_1494_),
    .B(_1556_));
 sg13g2_mux2_1 _5269_ (.A0(_1494_),
    .A1(_1579_),
    .S(_1558_),
    .X(_1580_));
 sg13g2_nand2_1 _5270_ (.Y(_1581_),
    .A(net796),
    .B(_1580_));
 sg13g2_or2_1 _5271_ (.X(_1583_),
    .B(_1499_),
    .A(_1493_));
 sg13g2_and3_1 _5272_ (.X(_1584_),
    .A(net787),
    .B(_1559_),
    .C(_1583_));
 sg13g2_inv_1 _5273_ (.Y(_1585_),
    .A(_1584_));
 sg13g2_a21oi_1 _5274_ (.A1(net788),
    .A2(_1559_),
    .Y(_1586_),
    .B1(_1583_));
 sg13g2_or2_1 _5275_ (.X(_1587_),
    .B(_1586_),
    .A(_1584_));
 sg13g2_xor2_1 _5276_ (.B(_1587_),
    .A(_1581_),
    .X(_1588_));
 sg13g2_a21oi_2 _5277_ (.B1(_1515_),
    .Y(_1589_),
    .A2(_1512_),
    .A1(_1504_));
 sg13g2_nand2_1 _5278_ (.Y(_1590_),
    .A(net782),
    .B(_1563_));
 sg13g2_nor2_1 _5279_ (.A(_0020_),
    .B(_1492_),
    .Y(_1591_));
 sg13g2_nor2_1 _5280_ (.A(_0020_),
    .B(_1446_),
    .Y(_1592_));
 sg13g2_nor2_1 _5281_ (.A(net739),
    .B(_1492_),
    .Y(_1594_));
 sg13g2_xnor2_1 _5282_ (.Y(_1595_),
    .A(_1592_),
    .B(_1594_));
 sg13g2_nor2_1 _5283_ (.A(_1590_),
    .B(_1595_),
    .Y(_1596_));
 sg13g2_xor2_1 _5284_ (.B(_1595_),
    .A(_1590_),
    .X(_1597_));
 sg13g2_nor2_2 _5285_ (.A(_1508_),
    .B(_1511_),
    .Y(_1598_));
 sg13g2_nand2_1 _5286_ (.Y(_1599_),
    .A(net766),
    .B(net677));
 sg13g2_nand2_1 _5287_ (.Y(_1600_),
    .A(_1472_),
    .B(net680));
 sg13g2_nand3_1 _5288_ (.B(net680),
    .C(_1507_),
    .A(net763),
    .Y(_1601_));
 sg13g2_a21o_1 _5289_ (.A2(net680),
    .A1(net763),
    .B1(_1507_),
    .X(_1602_));
 sg13g2_nand2_1 _5290_ (.Y(_1603_),
    .A(_1601_),
    .B(_1602_));
 sg13g2_xor2_1 _5291_ (.B(_1603_),
    .A(_1599_),
    .X(_1605_));
 sg13g2_nor2b_1 _5292_ (.A(_1598_),
    .B_N(_1605_),
    .Y(_1606_));
 sg13g2_xor2_1 _5293_ (.B(_1605_),
    .A(_1598_),
    .X(_1607_));
 sg13g2_inv_1 _5294_ (.Y(_1608_),
    .A(_1607_));
 sg13g2_xnor2_1 _5295_ (.Y(_1609_),
    .A(_1597_),
    .B(_1608_));
 sg13g2_nor2_1 _5296_ (.A(_1589_),
    .B(_1609_),
    .Y(_1610_));
 sg13g2_xor2_1 _5297_ (.B(_1609_),
    .A(_1589_),
    .X(_1611_));
 sg13g2_xnor2_1 _5298_ (.Y(_1612_),
    .A(_1588_),
    .B(_1611_));
 sg13g2_nor2b_1 _5299_ (.A(_1612_),
    .B_N(_1578_),
    .Y(_1613_));
 sg13g2_nand2_1 _5300_ (.Y(_1614_),
    .A(_1564_),
    .B(_1569_));
 sg13g2_xnor2_1 _5301_ (.Y(_1616_),
    .A(_1578_),
    .B(_1612_));
 sg13g2_a21oi_2 _5302_ (.B1(_1613_),
    .Y(_1617_),
    .A2(_1616_),
    .A1(_1614_));
 sg13g2_nand2_1 _5303_ (.Y(_1618_),
    .A(net766),
    .B(net674));
 sg13g2_nand2_1 _5304_ (.Y(_1619_),
    .A(net774),
    .B(_1563_));
 sg13g2_o21ai_1 _5305_ (.B1(_1601_),
    .Y(_1620_),
    .A1(_1599_),
    .A2(_1603_));
 sg13g2_nand2_1 _5306_ (.Y(_1621_),
    .A(net763),
    .B(net677));
 sg13g2_xnor2_1 _5307_ (.Y(_1622_),
    .A(_1600_),
    .B(_1621_));
 sg13g2_xnor2_1 _5308_ (.Y(_1623_),
    .A(_1620_),
    .B(_1622_));
 sg13g2_xnor2_1 _5309_ (.Y(_1624_),
    .A(_1591_),
    .B(_1623_));
 sg13g2_xnor2_1 _5310_ (.Y(_1625_),
    .A(_1619_),
    .B(_1624_));
 sg13g2_xnor2_1 _5311_ (.Y(_1627_),
    .A(_1618_),
    .B(_1625_));
 sg13g2_nand2_1 _5312_ (.Y(_1628_),
    .A(_1545_),
    .B(_1555_));
 sg13g2_nand3_1 _5313_ (.B(_1579_),
    .C(_1628_),
    .A(net796),
    .Y(_1629_));
 sg13g2_nand2_1 _5314_ (.Y(_1630_),
    .A(net781),
    .B(_1559_));
 sg13g2_a21oi_1 _5315_ (.A1(_1597_),
    .A2(_1608_),
    .Y(_1631_),
    .B1(_1606_));
 sg13g2_o21ai_1 _5316_ (.B1(_1585_),
    .Y(_1632_),
    .A1(_1581_),
    .A2(_1587_));
 sg13g2_nand2_1 _5317_ (.Y(_1633_),
    .A(net786),
    .B(_1580_));
 sg13g2_xnor2_1 _5318_ (.Y(_1634_),
    .A(_1627_),
    .B(_1630_));
 sg13g2_xnor2_1 _5319_ (.Y(_1635_),
    .A(_1632_),
    .B(_1634_));
 sg13g2_xor2_1 _5320_ (.B(_1631_),
    .A(_1629_),
    .X(_1636_));
 sg13g2_xnor2_1 _5321_ (.Y(_1638_),
    .A(_1633_),
    .B(_1636_));
 sg13g2_xnor2_1 _5322_ (.Y(_1639_),
    .A(_1635_),
    .B(_1638_));
 sg13g2_a21oi_1 _5323_ (.A1(_1592_),
    .A2(_1594_),
    .Y(_1640_),
    .B1(_1596_));
 sg13g2_a21oi_1 _5324_ (.A1(_1588_),
    .A2(_1611_),
    .Y(_1641_),
    .B1(_1610_));
 sg13g2_xor2_1 _5325_ (.B(_1641_),
    .A(_1640_),
    .X(_1642_));
 sg13g2_xnor2_1 _5326_ (.Y(_1643_),
    .A(_1639_),
    .B(_1642_));
 sg13g2_xnor2_1 _5327_ (.Y(_1644_),
    .A(_1617_),
    .B(_1643_));
 sg13g2_xor2_1 _5328_ (.B(_1643_),
    .A(_1617_),
    .X(_1645_));
 sg13g2_and2_2 _5329_ (.A(net762),
    .B(_0908_),
    .X(_1646_));
 sg13g2_nand2_1 _5330_ (.Y(_1647_),
    .A(net765),
    .B(net691));
 sg13g2_a22oi_1 _5331_ (.Y(_1649_),
    .B1(net694),
    .B2(_1472_),
    .A2(net692),
    .A1(net762));
 sg13g2_a21oi_1 _5332_ (.A1(_1265_),
    .A2(_1646_),
    .Y(_1650_),
    .B1(_1649_));
 sg13g2_nor2b_1 _5333_ (.A(_1647_),
    .B_N(_1650_),
    .Y(_1651_));
 sg13g2_a21oi_2 _5334_ (.B1(_1651_),
    .Y(_1652_),
    .A2(_1646_),
    .A1(_1265_));
 sg13g2_xor2_1 _5335_ (.B(_1269_),
    .A(_1268_),
    .X(_1653_));
 sg13g2_nor2b_1 _5336_ (.A(_1652_),
    .B_N(_1653_),
    .Y(_1654_));
 sg13g2_nor2_1 _5337_ (.A(net738),
    .B(_1322_),
    .Y(_1655_));
 sg13g2_nor2_1 _5338_ (.A(net741),
    .B(net682),
    .Y(_1656_));
 sg13g2_nand2_1 _5339_ (.Y(_1657_),
    .A(net769),
    .B(net684));
 sg13g2_nor3_1 _5340_ (.A(net738),
    .B(_1448_),
    .C(_1657_),
    .Y(_1658_));
 sg13g2_nand3_1 _5341_ (.B(net680),
    .C(_1655_),
    .A(net769),
    .Y(_1660_));
 sg13g2_a21oi_1 _5342_ (.A1(net774),
    .A2(net680),
    .Y(_1661_),
    .B1(_1656_));
 sg13g2_o21ai_1 _5343_ (.B1(_1657_),
    .Y(_1662_),
    .A1(net738),
    .A2(net678));
 sg13g2_a21oi_1 _5344_ (.A1(net774),
    .A2(net680),
    .Y(_1663_),
    .B1(_1657_));
 sg13g2_nor3_1 _5345_ (.A(net738),
    .B(net678),
    .C(_1656_),
    .Y(_1664_));
 sg13g2_nor4_2 _5346_ (.A(net733),
    .B(_1451_),
    .C(_1658_),
    .Y(_1665_),
    .D(_1661_));
 sg13g2_a22oi_1 _5347_ (.Y(_1666_),
    .B1(_1660_),
    .B2(_1662_),
    .A2(net677),
    .A1(net781));
 sg13g2_nor4_1 _5348_ (.A(net733),
    .B(_1451_),
    .C(_1663_),
    .D(_1664_),
    .Y(_1667_));
 sg13g2_a221oi_1 _5349_ (.B2(_1655_),
    .C1(_1661_),
    .B1(_1454_),
    .A1(net781),
    .Y(_1668_),
    .A2(net676));
 sg13g2_xnor2_1 _5350_ (.Y(_1669_),
    .A(_1652_),
    .B(_1653_));
 sg13g2_xor2_1 _5351_ (.B(_1653_),
    .A(_1652_),
    .X(_1671_));
 sg13g2_nor3_2 _5352_ (.A(_1665_),
    .B(_1666_),
    .C(_1671_),
    .Y(_1672_));
 sg13g2_o21ai_1 _5353_ (.B1(_1669_),
    .Y(_1673_),
    .A1(_1667_),
    .A2(_1668_));
 sg13g2_nor2_1 _5354_ (.A(_1654_),
    .B(_1672_),
    .Y(_1674_));
 sg13g2_xnor2_1 _5355_ (.Y(_1675_),
    .A(_1460_),
    .B(_1462_));
 sg13g2_nor2_1 _5356_ (.A(_1674_),
    .B(_1675_),
    .Y(_1676_));
 sg13g2_or2_1 _5357_ (.X(_1677_),
    .B(_1665_),
    .A(_1658_));
 sg13g2_nor2_1 _5358_ (.A(net730),
    .B(_1492_),
    .Y(_1678_));
 sg13g2_nand3_1 _5359_ (.B(_1491_),
    .C(_1677_),
    .A(net786),
    .Y(_1679_));
 sg13g2_a21o_1 _5360_ (.A2(net673),
    .A1(net786),
    .B1(_1677_),
    .X(_1680_));
 sg13g2_and4_1 _5361_ (.A(net795),
    .B(_1563_),
    .C(_1679_),
    .D(_1680_),
    .X(_1682_));
 sg13g2_a22oi_1 _5362_ (.Y(_1683_),
    .B1(_1679_),
    .B2(_1680_),
    .A2(_1563_),
    .A1(net795));
 sg13g2_nor2_1 _5363_ (.A(_1682_),
    .B(_1683_),
    .Y(_1684_));
 sg13g2_xor2_1 _5364_ (.B(_1675_),
    .A(_1674_),
    .X(_1685_));
 sg13g2_a21oi_1 _5365_ (.A1(_1684_),
    .A2(_1685_),
    .Y(_1686_),
    .B1(_1676_));
 sg13g2_a21o_1 _5366_ (.A2(_1685_),
    .A1(_1684_),
    .B1(_1676_),
    .X(_1687_));
 sg13g2_or4_1 _5367_ (.A(_1572_),
    .B(_1573_),
    .C(_1575_),
    .D(_1576_),
    .X(_1688_));
 sg13g2_nand3_1 _5368_ (.B(_1687_),
    .C(_1688_),
    .A(_1577_),
    .Y(_1689_));
 sg13g2_a21oi_1 _5369_ (.A1(_1677_),
    .A2(_1678_),
    .Y(_1690_),
    .B1(_1682_));
 sg13g2_a21oi_1 _5370_ (.A1(_1577_),
    .A2(_1688_),
    .Y(_1691_),
    .B1(_1686_));
 sg13g2_nand3_1 _5371_ (.B(_1686_),
    .C(_1688_),
    .A(_1577_),
    .Y(_1693_));
 sg13g2_nor2b_1 _5372_ (.A(_1691_),
    .B_N(_1693_),
    .Y(_1694_));
 sg13g2_o21ai_1 _5373_ (.B1(_1689_),
    .Y(_1695_),
    .A1(_1690_),
    .A2(_1694_));
 sg13g2_xnor2_1 _5374_ (.Y(_1696_),
    .A(_1614_),
    .B(_1616_));
 sg13g2_nand2b_1 _5375_ (.Y(_1697_),
    .B(_1695_),
    .A_N(_1696_));
 sg13g2_and2_1 _5376_ (.A(_1644_),
    .B(_1697_),
    .X(_1698_));
 sg13g2_nand2b_1 _5377_ (.Y(_1699_),
    .B(_1696_),
    .A_N(_1695_));
 sg13g2_nor2_2 _5378_ (.A(_0019_),
    .B(net696),
    .Y(_1700_));
 sg13g2_nand2_1 _5379_ (.Y(_1701_),
    .A(net765),
    .B(_0905_));
 sg13g2_xor2_1 _5380_ (.B(_1700_),
    .A(_1646_),
    .X(_1702_));
 sg13g2_nor2b_1 _5381_ (.A(_1701_),
    .B_N(_1702_),
    .Y(_1704_));
 sg13g2_a21oi_2 _5382_ (.B1(_1704_),
    .Y(_1705_),
    .A2(_1700_),
    .A1(_1646_));
 sg13g2_xnor2_1 _5383_ (.Y(_1706_),
    .A(_1647_),
    .B(_1650_));
 sg13g2_nor2b_1 _5384_ (.A(_1705_),
    .B_N(_1706_),
    .Y(_1707_));
 sg13g2_nor2_1 _5385_ (.A(net737),
    .B(net685),
    .Y(_1708_));
 sg13g2_nor2_1 _5386_ (.A(net741),
    .B(_1099_),
    .Y(_1709_));
 sg13g2_nand2_1 _5387_ (.Y(_1710_),
    .A(net768),
    .B(net687));
 sg13g2_nor3_1 _5388_ (.A(net736),
    .B(net682),
    .C(_1710_),
    .Y(_1711_));
 sg13g2_nand3_1 _5389_ (.B(net684),
    .C(_1708_),
    .A(net768),
    .Y(_1712_));
 sg13g2_a21oi_1 _5390_ (.A1(net774),
    .A2(net684),
    .Y(_1713_),
    .B1(_1709_));
 sg13g2_o21ai_1 _5391_ (.B1(_1710_),
    .Y(_1714_),
    .A1(net736),
    .A2(net682));
 sg13g2_a21oi_1 _5392_ (.A1(net774),
    .A2(net684),
    .Y(_1715_),
    .B1(_1710_));
 sg13g2_nor3_1 _5393_ (.A(net737),
    .B(net682),
    .C(_1709_),
    .Y(_1716_));
 sg13g2_nor4_2 _5394_ (.A(net733),
    .B(net678),
    .C(_1711_),
    .Y(_1717_),
    .D(_1713_));
 sg13g2_a22oi_1 _5395_ (.Y(_1718_),
    .B1(_1712_),
    .B2(_1714_),
    .A2(net679),
    .A1(net781));
 sg13g2_nor4_1 _5396_ (.A(net733),
    .B(net678),
    .C(_1715_),
    .D(_1716_),
    .Y(_1719_));
 sg13g2_a221oi_1 _5397_ (.B2(_1708_),
    .C1(_1713_),
    .B1(_1656_),
    .A1(net781),
    .Y(_1720_),
    .A2(net679));
 sg13g2_xnor2_1 _5398_ (.Y(_1721_),
    .A(_1705_),
    .B(_1706_));
 sg13g2_xor2_1 _5399_ (.B(_1706_),
    .A(_1705_),
    .X(_1722_));
 sg13g2_nor3_1 _5400_ (.A(_1717_),
    .B(_1718_),
    .C(_1722_),
    .Y(_1723_));
 sg13g2_o21ai_1 _5401_ (.B1(_1721_),
    .Y(_1724_),
    .A1(_1719_),
    .A2(_1720_));
 sg13g2_nor2_1 _5402_ (.A(_1707_),
    .B(_1723_),
    .Y(_1725_));
 sg13g2_nand2b_1 _5403_ (.Y(_1726_),
    .B(_1724_),
    .A_N(_1707_));
 sg13g2_nor3_1 _5404_ (.A(_1667_),
    .B(_1668_),
    .C(_1669_),
    .Y(_1727_));
 sg13g2_o21ai_1 _5405_ (.B1(_1671_),
    .Y(_1728_),
    .A1(_1665_),
    .A2(_1666_));
 sg13g2_nor3_1 _5406_ (.A(_1672_),
    .B(_1725_),
    .C(_1727_),
    .Y(_1729_));
 sg13g2_or2_2 _5407_ (.X(_1730_),
    .B(_1717_),
    .A(_1711_));
 sg13g2_nor2_1 _5408_ (.A(net730),
    .B(_1446_),
    .Y(_1731_));
 sg13g2_nand3_1 _5409_ (.B(net674),
    .C(_1730_),
    .A(net787),
    .Y(_1732_));
 sg13g2_a21o_1 _5410_ (.A2(net674),
    .A1(net787),
    .B1(_1730_),
    .X(_1733_));
 sg13g2_or3_1 _5411_ (.A(net730),
    .B(_1446_),
    .C(_1730_),
    .X(_1734_));
 sg13g2_o21ai_1 _5412_ (.B1(_1730_),
    .Y(_1735_),
    .A1(net730),
    .A2(_1446_));
 sg13g2_and4_1 _5413_ (.A(net796),
    .B(net673),
    .C(_1732_),
    .D(_1733_),
    .X(_1736_));
 sg13g2_a22oi_1 _5414_ (.Y(_1737_),
    .B1(_1732_),
    .B2(_1733_),
    .A2(net673),
    .A1(net796));
 sg13g2_and4_1 _5415_ (.A(net796),
    .B(net673),
    .C(_1734_),
    .D(_1735_),
    .X(_1738_));
 sg13g2_a22oi_1 _5416_ (.Y(_1739_),
    .B1(_1734_),
    .B2(_1735_),
    .A2(net673),
    .A1(net794));
 sg13g2_a21oi_1 _5417_ (.A1(_1673_),
    .A2(_1728_),
    .Y(_1740_),
    .B1(_1726_));
 sg13g2_a21oi_1 _5418_ (.A1(_1673_),
    .A2(_1728_),
    .Y(_1741_),
    .B1(_1725_));
 sg13g2_nor3_1 _5419_ (.A(_1672_),
    .B(_1726_),
    .C(_1727_),
    .Y(_1742_));
 sg13g2_nor4_2 _5420_ (.A(_1729_),
    .B(_1736_),
    .C(_1737_),
    .Y(_1743_),
    .D(_1740_));
 sg13g2_or2_1 _5421_ (.X(_1744_),
    .B(_1743_),
    .A(_1729_));
 sg13g2_xor2_1 _5422_ (.B(_1685_),
    .A(_1684_),
    .X(_1745_));
 sg13g2_nand2_1 _5423_ (.Y(_1746_),
    .A(_1744_),
    .B(_1745_));
 sg13g2_a21oi_1 _5424_ (.A1(_1730_),
    .A2(_1731_),
    .Y(_1747_),
    .B1(_1736_));
 sg13g2_xnor2_1 _5425_ (.Y(_1748_),
    .A(_1744_),
    .B(_1745_));
 sg13g2_o21ai_1 _5426_ (.B1(_1746_),
    .Y(_1749_),
    .A1(_1747_),
    .A2(_1748_));
 sg13g2_xor2_1 _5427_ (.B(_1694_),
    .A(_1690_),
    .X(_1750_));
 sg13g2_nand2_1 _5428_ (.Y(_1751_),
    .A(_1749_),
    .B(_1750_));
 sg13g2_nor2_1 _5429_ (.A(_0019_),
    .B(_0721_),
    .Y(_1752_));
 sg13g2_nand3_1 _5430_ (.B(net698),
    .C(_1752_),
    .A(net761),
    .Y(_1753_));
 sg13g2_nand2_1 _5431_ (.Y(_1754_),
    .A(net764),
    .B(net694));
 sg13g2_a21o_1 _5432_ (.A2(net697),
    .A1(net761),
    .B1(_1752_),
    .X(_1755_));
 sg13g2_and2_1 _5433_ (.A(_1753_),
    .B(_1755_),
    .X(_1756_));
 sg13g2_nand2b_1 _5434_ (.Y(_1757_),
    .B(_1756_),
    .A_N(_1754_));
 sg13g2_and2_2 _5435_ (.A(_1753_),
    .B(_1757_),
    .X(_1758_));
 sg13g2_xnor2_1 _5436_ (.Y(_1759_),
    .A(_1701_),
    .B(_1702_));
 sg13g2_nor2b_1 _5437_ (.A(_1758_),
    .B_N(_1759_),
    .Y(_1760_));
 sg13g2_nor2_1 _5438_ (.A(net736),
    .B(net688),
    .Y(_1761_));
 sg13g2_nor2_1 _5439_ (.A(net740),
    .B(net688),
    .Y(_1762_));
 sg13g2_nand2_1 _5440_ (.Y(_1763_),
    .A(net769),
    .B(net691));
 sg13g2_nor3_1 _5441_ (.A(net736),
    .B(net685),
    .C(_1763_),
    .Y(_1764_));
 sg13g2_nand3_1 _5442_ (.B(net687),
    .C(_1761_),
    .A(net768),
    .Y(_1765_));
 sg13g2_a21oi_1 _5443_ (.A1(net773),
    .A2(net687),
    .Y(_1766_),
    .B1(_1762_));
 sg13g2_o21ai_1 _5444_ (.B1(_1763_),
    .Y(_1767_),
    .A1(net736),
    .A2(net685));
 sg13g2_a21oi_1 _5445_ (.A1(net773),
    .A2(net687),
    .Y(_1768_),
    .B1(_1763_));
 sg13g2_nor3_1 _5446_ (.A(net736),
    .B(net685),
    .C(_1762_),
    .Y(_1769_));
 sg13g2_nor4_2 _5447_ (.A(net733),
    .B(net682),
    .C(_1764_),
    .Y(_1770_),
    .D(_1766_));
 sg13g2_a22oi_1 _5448_ (.Y(_1771_),
    .B1(_1765_),
    .B2(_1767_),
    .A2(net684),
    .A1(net780));
 sg13g2_nor4_2 _5449_ (.A(net733),
    .B(net682),
    .C(_1768_),
    .Y(_1772_),
    .D(_1769_));
 sg13g2_a221oi_1 _5450_ (.B2(_1761_),
    .C1(_1766_),
    .B1(_1709_),
    .A1(net780),
    .Y(_1773_),
    .A2(net684));
 sg13g2_xnor2_1 _5451_ (.Y(_1774_),
    .A(_1758_),
    .B(_1759_));
 sg13g2_xor2_1 _5452_ (.B(_1759_),
    .A(_1758_),
    .X(_1775_));
 sg13g2_nor3_2 _5453_ (.A(_1770_),
    .B(_1771_),
    .C(_1775_),
    .Y(_1776_));
 sg13g2_o21ai_1 _5454_ (.B1(_1774_),
    .Y(_1777_),
    .A1(_1772_),
    .A2(_1773_));
 sg13g2_nor2_1 _5455_ (.A(_1760_),
    .B(_1776_),
    .Y(_1778_));
 sg13g2_nand2b_1 _5456_ (.Y(_1779_),
    .B(_1777_),
    .A_N(_1760_));
 sg13g2_nor3_1 _5457_ (.A(_1719_),
    .B(_1720_),
    .C(_1721_),
    .Y(_1780_));
 sg13g2_o21ai_1 _5458_ (.B1(_1722_),
    .Y(_1781_),
    .A1(_1717_),
    .A2(_1718_));
 sg13g2_nor3_1 _5459_ (.A(_1723_),
    .B(_1778_),
    .C(_1780_),
    .Y(_1782_));
 sg13g2_or2_1 _5460_ (.X(_1783_),
    .B(_1770_),
    .A(_1764_));
 sg13g2_nand3_1 _5461_ (.B(net676),
    .C(_1783_),
    .A(net787),
    .Y(_1784_));
 sg13g2_a21o_1 _5462_ (.A2(net676),
    .A1(net787),
    .B1(_1783_),
    .X(_1785_));
 sg13g2_or3_1 _5463_ (.A(net730),
    .B(_1451_),
    .C(_1783_),
    .X(_1786_));
 sg13g2_o21ai_1 _5464_ (.B1(_1783_),
    .Y(_1787_),
    .A1(net730),
    .A2(_1451_));
 sg13g2_and4_1 _5465_ (.A(net794),
    .B(net674),
    .C(_1784_),
    .D(_1785_),
    .X(_1788_));
 sg13g2_nand4_1 _5466_ (.B(net674),
    .C(_1784_),
    .A(net794),
    .Y(_1789_),
    .D(_1785_));
 sg13g2_a22oi_1 _5467_ (.Y(_1790_),
    .B1(_1784_),
    .B2(_1785_),
    .A2(net674),
    .A1(net794));
 sg13g2_and4_1 _5468_ (.A(net794),
    .B(net674),
    .C(_1786_),
    .D(_1787_),
    .X(_1791_));
 sg13g2_a22oi_1 _5469_ (.Y(_1792_),
    .B1(_1786_),
    .B2(_1787_),
    .A2(net674),
    .A1(net794));
 sg13g2_a21oi_1 _5470_ (.A1(_1724_),
    .A2(_1781_),
    .Y(_1793_),
    .B1(_1779_));
 sg13g2_a21oi_1 _5471_ (.A1(_1724_),
    .A2(_1781_),
    .Y(_1795_),
    .B1(_1778_));
 sg13g2_nor3_1 _5472_ (.A(_1723_),
    .B(_1779_),
    .C(_1780_),
    .Y(_1796_));
 sg13g2_or4_1 _5473_ (.A(_1782_),
    .B(_1788_),
    .C(_1790_),
    .D(_1793_),
    .X(_1797_));
 sg13g2_nor2b_1 _5474_ (.A(_1782_),
    .B_N(_1797_),
    .Y(_1798_));
 sg13g2_nor4_2 _5475_ (.A(_1738_),
    .B(_1739_),
    .C(_1741_),
    .Y(_1799_),
    .D(_1742_));
 sg13g2_nor3_1 _5476_ (.A(_1743_),
    .B(_1798_),
    .C(_1799_),
    .Y(_1800_));
 sg13g2_or3_1 _5477_ (.A(_1743_),
    .B(_1798_),
    .C(_1799_),
    .X(_1801_));
 sg13g2_nand2_1 _5478_ (.Y(_1802_),
    .A(_1784_),
    .B(_1789_));
 sg13g2_o21ai_1 _5479_ (.B1(_1798_),
    .Y(_1803_),
    .A1(_1743_),
    .A2(_1799_));
 sg13g2_and3_1 _5480_ (.X(_1804_),
    .A(_1801_),
    .B(_1802_),
    .C(_1803_));
 sg13g2_nor2_1 _5481_ (.A(_1800_),
    .B(_1804_),
    .Y(_1806_));
 sg13g2_xnor2_1 _5482_ (.Y(_1807_),
    .A(_1747_),
    .B(_1748_));
 sg13g2_nor2_1 _5483_ (.A(_1806_),
    .B(_1807_),
    .Y(_1808_));
 sg13g2_nor3_1 _5484_ (.A(_0019_),
    .B(_0721_),
    .C(_1029_),
    .Y(_1809_));
 sg13g2_and2_1 _5485_ (.A(net765),
    .B(net697),
    .X(_1810_));
 sg13g2_nand2_1 _5486_ (.Y(_1811_),
    .A(net764),
    .B(net697));
 sg13g2_a22oi_1 _5487_ (.Y(_1812_),
    .B1(net702),
    .B2(_1472_),
    .A2(net699),
    .A1(net761));
 sg13g2_nor2_1 _5488_ (.A(_1809_),
    .B(_1812_),
    .Y(_1813_));
 sg13g2_a21oi_2 _5489_ (.B1(_1809_),
    .Y(_1814_),
    .A2(_1813_),
    .A1(_1810_));
 sg13g2_xnor2_1 _5490_ (.Y(_1815_),
    .A(_1754_),
    .B(_1756_));
 sg13g2_nor2b_1 _5491_ (.A(_1814_),
    .B_N(_1815_),
    .Y(_1817_));
 sg13g2_nand2_1 _5492_ (.Y(_1818_),
    .A(net773),
    .B(net692));
 sg13g2_inv_1 _5493_ (.Y(_1819_),
    .A(_1818_));
 sg13g2_nor2_2 _5494_ (.A(net740),
    .B(_0906_),
    .Y(_1820_));
 sg13g2_nand2_1 _5495_ (.Y(_1821_),
    .A(net768),
    .B(_0905_));
 sg13g2_nor3_1 _5496_ (.A(net740),
    .B(net688),
    .C(_1818_),
    .Y(_1822_));
 sg13g2_nand3_1 _5497_ (.B(net690),
    .C(_1820_),
    .A(net772),
    .Y(_1823_));
 sg13g2_a21oi_1 _5498_ (.A1(net772),
    .A2(net690),
    .Y(_1824_),
    .B1(_1820_));
 sg13g2_o21ai_1 _5499_ (.B1(_1821_),
    .Y(_1825_),
    .A1(net736),
    .A2(net688));
 sg13g2_a21oi_1 _5500_ (.A1(net772),
    .A2(net690),
    .Y(_1826_),
    .B1(_1821_));
 sg13g2_nor3_1 _5501_ (.A(net736),
    .B(net688),
    .C(_1820_),
    .Y(_1828_));
 sg13g2_nor4_2 _5502_ (.A(net732),
    .B(net685),
    .C(_1822_),
    .Y(_1829_),
    .D(_1824_));
 sg13g2_a22oi_1 _5503_ (.Y(_1830_),
    .B1(_1823_),
    .B2(_1825_),
    .A2(net686),
    .A1(net779));
 sg13g2_nor4_2 _5504_ (.A(net732),
    .B(net685),
    .C(_1826_),
    .Y(_1831_),
    .D(_1828_));
 sg13g2_a221oi_1 _5505_ (.B2(_1819_),
    .C1(_1824_),
    .B1(_1762_),
    .A1(net779),
    .Y(_1832_),
    .A2(net686));
 sg13g2_xnor2_1 _5506_ (.Y(_1833_),
    .A(_1814_),
    .B(_1815_));
 sg13g2_xor2_1 _5507_ (.B(_1815_),
    .A(_1814_),
    .X(_1834_));
 sg13g2_nor3_2 _5508_ (.A(_1829_),
    .B(_1830_),
    .C(_1834_),
    .Y(_1835_));
 sg13g2_o21ai_1 _5509_ (.B1(_1833_),
    .Y(_1836_),
    .A1(_1831_),
    .A2(_1832_));
 sg13g2_nor2_1 _5510_ (.A(_1817_),
    .B(_1835_),
    .Y(_1837_));
 sg13g2_nand2b_1 _5511_ (.Y(_1838_),
    .B(_1836_),
    .A_N(_1817_));
 sg13g2_nor3_1 _5512_ (.A(_1772_),
    .B(_1773_),
    .C(_1774_),
    .Y(_1839_));
 sg13g2_o21ai_1 _5513_ (.B1(_1775_),
    .Y(_1840_),
    .A1(_1770_),
    .A2(_1771_));
 sg13g2_nor3_1 _5514_ (.A(_1776_),
    .B(_1837_),
    .C(_1839_),
    .Y(_1841_));
 sg13g2_or2_1 _5515_ (.X(_1842_),
    .B(_1829_),
    .A(_1822_));
 sg13g2_nand3_1 _5516_ (.B(net679),
    .C(_1842_),
    .A(net787),
    .Y(_1843_));
 sg13g2_a21o_1 _5517_ (.A2(net679),
    .A1(net787),
    .B1(_1842_),
    .X(_1844_));
 sg13g2_or3_1 _5518_ (.A(net730),
    .B(net678),
    .C(_1842_),
    .X(_1845_));
 sg13g2_o21ai_1 _5519_ (.B1(_1842_),
    .Y(_1846_),
    .A1(net730),
    .A2(net678));
 sg13g2_and4_1 _5520_ (.A(net794),
    .B(net676),
    .C(_1843_),
    .D(_1844_),
    .X(_1847_));
 sg13g2_nand4_1 _5521_ (.B(net676),
    .C(_1843_),
    .A(net794),
    .Y(_1849_),
    .D(_1844_));
 sg13g2_a22oi_1 _5522_ (.Y(_1850_),
    .B1(_1843_),
    .B2(_1844_),
    .A2(net676),
    .A1(net792));
 sg13g2_and4_1 _5523_ (.A(net792),
    .B(net676),
    .C(_1845_),
    .D(_1846_),
    .X(_1851_));
 sg13g2_a22oi_1 _5524_ (.Y(_1852_),
    .B1(_1845_),
    .B2(_1846_),
    .A2(net676),
    .A1(net792));
 sg13g2_a21oi_1 _5525_ (.A1(_1777_),
    .A2(_1840_),
    .Y(_1853_),
    .B1(_1838_));
 sg13g2_a21oi_1 _5526_ (.A1(_1777_),
    .A2(_1840_),
    .Y(_1854_),
    .B1(_1837_));
 sg13g2_nor3_1 _5527_ (.A(_1776_),
    .B(_1838_),
    .C(_1839_),
    .Y(_1855_));
 sg13g2_nor4_1 _5528_ (.A(_1841_),
    .B(_1847_),
    .C(_1850_),
    .D(_1853_),
    .Y(_1856_));
 sg13g2_or4_1 _5529_ (.A(_1841_),
    .B(_1847_),
    .C(_1850_),
    .D(_1853_),
    .X(_1857_));
 sg13g2_nand2b_1 _5530_ (.Y(_1858_),
    .B(_1857_),
    .A_N(_1841_));
 sg13g2_or4_1 _5531_ (.A(_1791_),
    .B(_1792_),
    .C(_1795_),
    .D(_1796_),
    .X(_1860_));
 sg13g2_nand3_1 _5532_ (.B(_1858_),
    .C(_1860_),
    .A(_1797_),
    .Y(_1861_));
 sg13g2_nand2_1 _5533_ (.Y(_1862_),
    .A(_1843_),
    .B(_1849_));
 sg13g2_a21o_1 _5534_ (.A2(_1860_),
    .A1(_1797_),
    .B1(_1858_),
    .X(_1863_));
 sg13g2_nand3_1 _5535_ (.B(_1862_),
    .C(_1863_),
    .A(_1861_),
    .Y(_1864_));
 sg13g2_and2_1 _5536_ (.A(_1861_),
    .B(_1864_),
    .X(_1865_));
 sg13g2_a21oi_1 _5537_ (.A1(_1801_),
    .A2(_1803_),
    .Y(_1866_),
    .B1(_1802_));
 sg13g2_nor3_1 _5538_ (.A(_1804_),
    .B(_1865_),
    .C(_1866_),
    .Y(_1867_));
 sg13g2_o21ai_1 _5539_ (.B1(_1032_),
    .Y(_1868_),
    .A1(_1029_),
    .A2(_1030_));
 sg13g2_xnor2_1 _5540_ (.Y(_1869_),
    .A(_1811_),
    .B(_1813_));
 sg13g2_nor3_1 _5541_ (.A(net741),
    .B(_0906_),
    .C(_1038_),
    .Y(_1871_));
 sg13g2_nand3_1 _5542_ (.B(net693),
    .C(_1036_),
    .A(net772),
    .Y(_1872_));
 sg13g2_a21oi_1 _5543_ (.A1(net772),
    .A2(net692),
    .Y(_1873_),
    .B1(_1036_));
 sg13g2_o21ai_1 _5544_ (.B1(_1037_),
    .Y(_1874_),
    .A1(net734),
    .A2(_0906_));
 sg13g2_a21oi_1 _5545_ (.A1(net773),
    .A2(net692),
    .Y(_1875_),
    .B1(_1037_));
 sg13g2_nor3_1 _5546_ (.A(net735),
    .B(_0906_),
    .C(_1036_),
    .Y(_1876_));
 sg13g2_nor4_2 _5547_ (.A(net732),
    .B(_0968_),
    .C(_1871_),
    .Y(_1877_),
    .D(_1873_));
 sg13g2_a22oi_1 _5548_ (.Y(_1878_),
    .B1(_1872_),
    .B2(_1874_),
    .A2(net690),
    .A1(net779));
 sg13g2_nor4_2 _5549_ (.A(net732),
    .B(net688),
    .C(_1875_),
    .Y(_1879_),
    .D(_1876_));
 sg13g2_a221oi_1 _5550_ (.B2(_1820_),
    .C1(_1873_),
    .B1(_1039_),
    .A1(net779),
    .Y(_1880_),
    .A2(net690));
 sg13g2_xnor2_1 _5551_ (.Y(_1882_),
    .A(_1868_),
    .B(_1869_));
 sg13g2_inv_1 _5552_ (.Y(_1883_),
    .A(_1882_));
 sg13g2_nor3_2 _5553_ (.A(_1877_),
    .B(_1878_),
    .C(_1882_),
    .Y(_1884_));
 sg13g2_o21ai_1 _5554_ (.B1(_1883_),
    .Y(_1885_),
    .A1(_1879_),
    .A2(_1880_));
 sg13g2_a21oi_1 _5555_ (.A1(_1868_),
    .A2(_1869_),
    .Y(_1886_),
    .B1(_1884_));
 sg13g2_a21o_1 _5556_ (.A2(_1869_),
    .A1(_1868_),
    .B1(_1884_),
    .X(_1887_));
 sg13g2_nor3_1 _5557_ (.A(_1831_),
    .B(_1832_),
    .C(_1833_),
    .Y(_1888_));
 sg13g2_o21ai_1 _5558_ (.B1(_1834_),
    .Y(_1889_),
    .A1(_1829_),
    .A2(_1830_));
 sg13g2_nor3_1 _5559_ (.A(_1835_),
    .B(_1886_),
    .C(_1888_),
    .Y(_1890_));
 sg13g2_or2_1 _5560_ (.X(_1891_),
    .B(_1877_),
    .A(_1871_));
 sg13g2_and3_1 _5561_ (.X(_1893_),
    .A(net785),
    .B(net683),
    .C(_1891_));
 sg13g2_nand3_1 _5562_ (.B(net683),
    .C(_1891_),
    .A(net785),
    .Y(_1894_));
 sg13g2_a21o_1 _5563_ (.A2(net683),
    .A1(net785),
    .B1(_1891_),
    .X(_1895_));
 sg13g2_or3_1 _5564_ (.A(net728),
    .B(net682),
    .C(_1891_),
    .X(_1896_));
 sg13g2_o21ai_1 _5565_ (.B1(_1891_),
    .Y(_1897_),
    .A1(net729),
    .A2(net682));
 sg13g2_and4_1 _5566_ (.A(net792),
    .B(net679),
    .C(_1894_),
    .D(_1895_),
    .X(_1898_));
 sg13g2_a22oi_1 _5567_ (.Y(_1899_),
    .B1(_1894_),
    .B2(_1895_),
    .A2(net679),
    .A1(net792));
 sg13g2_and4_1 _5568_ (.A(net793),
    .B(net679),
    .C(_1896_),
    .D(_1897_),
    .X(_1900_));
 sg13g2_a22oi_1 _5569_ (.Y(_1901_),
    .B1(_1896_),
    .B2(_1897_),
    .A2(net679),
    .A1(net797));
 sg13g2_a21oi_1 _5570_ (.A1(_1836_),
    .A2(_1889_),
    .Y(_1902_),
    .B1(_1887_));
 sg13g2_a21oi_1 _5571_ (.A1(_1836_),
    .A2(_1889_),
    .Y(_1904_),
    .B1(_1886_));
 sg13g2_nor3_1 _5572_ (.A(_1835_),
    .B(_1887_),
    .C(_1888_),
    .Y(_1905_));
 sg13g2_or4_1 _5573_ (.A(_1890_),
    .B(_1898_),
    .C(_1899_),
    .D(_1902_),
    .X(_1906_));
 sg13g2_nor2b_1 _5574_ (.A(_1890_),
    .B_N(_1906_),
    .Y(_1907_));
 sg13g2_nand2b_1 _5575_ (.Y(_1908_),
    .B(_1906_),
    .A_N(_1890_));
 sg13g2_nor4_1 _5576_ (.A(_1851_),
    .B(_1852_),
    .C(_1854_),
    .D(_1855_),
    .Y(_1909_));
 sg13g2_or4_1 _5577_ (.A(_1851_),
    .B(_1852_),
    .C(_1854_),
    .D(_1855_),
    .X(_1910_));
 sg13g2_nor3_1 _5578_ (.A(_1856_),
    .B(_1907_),
    .C(_1909_),
    .Y(_1911_));
 sg13g2_nand3_1 _5579_ (.B(_1908_),
    .C(_1910_),
    .A(_1857_),
    .Y(_1912_));
 sg13g2_nor2_1 _5580_ (.A(_1893_),
    .B(_1898_),
    .Y(_1913_));
 sg13g2_or2_1 _5581_ (.X(_1915_),
    .B(_1898_),
    .A(_1893_));
 sg13g2_a21oi_1 _5582_ (.A1(_1857_),
    .A2(_1910_),
    .Y(_1916_),
    .B1(_1908_));
 sg13g2_o21ai_1 _5583_ (.B1(_1907_),
    .Y(_1917_),
    .A1(_1856_),
    .A2(_1909_));
 sg13g2_nor3_1 _5584_ (.A(_1911_),
    .B(_1913_),
    .C(_1916_),
    .Y(_1918_));
 sg13g2_nor2_1 _5585_ (.A(_1911_),
    .B(_1918_),
    .Y(_1919_));
 sg13g2_o21ai_1 _5586_ (.B1(_1912_),
    .Y(_1920_),
    .A1(_1913_),
    .A2(_1916_));
 sg13g2_a21o_1 _5587_ (.A2(_1863_),
    .A1(_1861_),
    .B1(_1862_),
    .X(_1921_));
 sg13g2_nand3_1 _5588_ (.B(_1920_),
    .C(_1921_),
    .A(_1864_),
    .Y(_1922_));
 sg13g2_a21oi_1 _5589_ (.A1(_1027_),
    .A2(_1033_),
    .Y(_1923_),
    .B1(_1048_));
 sg13g2_a21o_1 _5590_ (.A2(_1033_),
    .A1(_1027_),
    .B1(_1048_),
    .X(_1924_));
 sg13g2_nor3_1 _5591_ (.A(_1879_),
    .B(_1880_),
    .C(_1883_),
    .Y(_1925_));
 sg13g2_o21ai_1 _5592_ (.B1(_1882_),
    .Y(_1926_),
    .A1(_1877_),
    .A2(_1878_));
 sg13g2_nor3_1 _5593_ (.A(_1884_),
    .B(_1923_),
    .C(_1925_),
    .Y(_1927_));
 sg13g2_a21o_1 _5594_ (.A2(_1039_),
    .A1(_0981_),
    .B1(_1044_),
    .X(_1928_));
 sg13g2_nand3_1 _5595_ (.B(net686),
    .C(_1928_),
    .A(net785),
    .Y(_1929_));
 sg13g2_a21o_1 _5596_ (.A2(net686),
    .A1(net785),
    .B1(_1928_),
    .X(_1930_));
 sg13g2_or3_1 _5597_ (.A(net729),
    .B(net685),
    .C(_1928_),
    .X(_1931_));
 sg13g2_o21ai_1 _5598_ (.B1(_1928_),
    .Y(_1932_),
    .A1(net729),
    .A2(net685));
 sg13g2_and4_1 _5599_ (.A(net792),
    .B(net683),
    .C(_1929_),
    .D(_1930_),
    .X(_1933_));
 sg13g2_nand4_1 _5600_ (.B(net683),
    .C(_1929_),
    .A(net792),
    .Y(_1934_),
    .D(_1930_));
 sg13g2_a22oi_1 _5601_ (.Y(_1935_),
    .B1(_1929_),
    .B2(_1930_),
    .A2(net683),
    .A1(net792));
 sg13g2_and4_1 _5602_ (.A(net793),
    .B(net683),
    .C(_1931_),
    .D(_1932_),
    .X(_1936_));
 sg13g2_a22oi_1 _5603_ (.Y(_1937_),
    .B1(_1931_),
    .B2(_1932_),
    .A2(net683),
    .A1(net793));
 sg13g2_a21oi_1 _5604_ (.A1(_1885_),
    .A2(_1926_),
    .Y(_1938_),
    .B1(_1924_));
 sg13g2_a21oi_1 _5605_ (.A1(_1885_),
    .A2(_1926_),
    .Y(_1939_),
    .B1(_1923_));
 sg13g2_nor3_1 _5606_ (.A(_1884_),
    .B(_1924_),
    .C(_1925_),
    .Y(_1940_));
 sg13g2_or4_1 _5607_ (.A(_1927_),
    .B(_1933_),
    .C(_1935_),
    .D(_1938_),
    .X(_1941_));
 sg13g2_nand2b_1 _5608_ (.Y(_1942_),
    .B(_1941_),
    .A_N(_1927_));
 sg13g2_or4_1 _5609_ (.A(_1900_),
    .B(_1901_),
    .C(_1904_),
    .D(_1905_),
    .X(_1943_));
 sg13g2_nand3_1 _5610_ (.B(_1942_),
    .C(_1943_),
    .A(_1906_),
    .Y(_1944_));
 sg13g2_nand2_1 _5611_ (.Y(_1946_),
    .A(_1929_),
    .B(_1934_));
 sg13g2_a21o_1 _5612_ (.A2(_1943_),
    .A1(_1906_),
    .B1(_1942_),
    .X(_1947_));
 sg13g2_nand3_1 _5613_ (.B(_1946_),
    .C(_1947_),
    .A(_1944_),
    .Y(_1948_));
 sg13g2_and2_1 _5614_ (.A(_1944_),
    .B(_1948_),
    .X(_1949_));
 sg13g2_a21oi_1 _5615_ (.A1(_1912_),
    .A2(_1917_),
    .Y(_1950_),
    .B1(_1915_));
 sg13g2_nor3_1 _5616_ (.A(_1918_),
    .B(_1949_),
    .C(_1950_),
    .Y(_1951_));
 sg13g2_or2_1 _5617_ (.X(_1952_),
    .B(_1110_),
    .A(_1052_));
 sg13g2_or4_1 _5618_ (.A(_1936_),
    .B(_1937_),
    .C(_1939_),
    .D(_1940_),
    .X(_1953_));
 sg13g2_nand3_1 _5619_ (.B(_1952_),
    .C(_1953_),
    .A(_1941_),
    .Y(_1954_));
 sg13g2_nor2_1 _5620_ (.A(_1101_),
    .B(_1106_),
    .Y(_1955_));
 sg13g2_or2_1 _5621_ (.X(_1957_),
    .B(_1106_),
    .A(_1101_));
 sg13g2_a21oi_1 _5622_ (.A1(_1941_),
    .A2(_1953_),
    .Y(_1958_),
    .B1(_1952_));
 sg13g2_a21o_1 _5623_ (.A2(_1953_),
    .A1(_1941_),
    .B1(_1952_),
    .X(_1959_));
 sg13g2_and3_1 _5624_ (.X(_1960_),
    .A(_1954_),
    .B(_1957_),
    .C(_1959_));
 sg13g2_o21ai_1 _5625_ (.B1(_1954_),
    .Y(_1961_),
    .A1(_1955_),
    .A2(_1958_));
 sg13g2_a21o_1 _5626_ (.A2(_1947_),
    .A1(_1944_),
    .B1(_1946_),
    .X(_1962_));
 sg13g2_and2_1 _5627_ (.A(_1948_),
    .B(_1962_),
    .X(_1963_));
 sg13g2_nand3_1 _5628_ (.B(_1961_),
    .C(_1962_),
    .A(_1948_),
    .Y(_1964_));
 sg13g2_and2_1 _5629_ (.A(_1112_),
    .B(_1114_),
    .X(_1965_));
 sg13g2_a21oi_1 _5630_ (.A1(_1954_),
    .A2(_1959_),
    .Y(_1966_),
    .B1(_1957_));
 sg13g2_nor3_1 _5631_ (.A(_1960_),
    .B(_1965_),
    .C(_1966_),
    .Y(_1968_));
 sg13g2_o21ai_1 _5632_ (.B1(_1116_),
    .Y(_1969_),
    .A1(_1117_),
    .A2(_1261_));
 sg13g2_o21ai_1 _5633_ (.B1(_1965_),
    .Y(_1970_),
    .A1(_1960_),
    .A2(_1966_));
 sg13g2_nor2b_1 _5634_ (.A(_1968_),
    .B_N(_1970_),
    .Y(_1971_));
 sg13g2_a21oi_2 _5635_ (.B1(_1968_),
    .Y(_1972_),
    .A2(_1970_),
    .A1(_1969_));
 sg13g2_a21oi_1 _5636_ (.A1(_1948_),
    .A2(_1962_),
    .Y(_1973_),
    .B1(_1961_));
 sg13g2_xnor2_1 _5637_ (.Y(_1974_),
    .A(_1961_),
    .B(_1963_));
 sg13g2_o21ai_1 _5638_ (.B1(_1964_),
    .Y(_1975_),
    .A1(_1972_),
    .A2(_1973_));
 sg13g2_o21ai_1 _5639_ (.B1(_1949_),
    .Y(_1976_),
    .A1(_1918_),
    .A2(_1950_));
 sg13g2_nand2b_1 _5640_ (.Y(_1977_),
    .B(_1976_),
    .A_N(_1951_));
 sg13g2_a21oi_1 _5641_ (.A1(_1975_),
    .A2(_1976_),
    .Y(_1978_),
    .B1(_1951_));
 sg13g2_a21oi_1 _5642_ (.A1(_1864_),
    .A2(_1921_),
    .Y(_1979_),
    .B1(_1920_));
 sg13g2_a21oi_1 _5643_ (.A1(_1864_),
    .A2(_1921_),
    .Y(_1980_),
    .B1(_1919_));
 sg13g2_nand3_1 _5644_ (.B(_1919_),
    .C(_1921_),
    .A(_1864_),
    .Y(_1981_));
 sg13g2_nand2b_1 _5645_ (.Y(_1982_),
    .B(_1981_),
    .A_N(_1980_));
 sg13g2_o21ai_1 _5646_ (.B1(_1922_),
    .Y(_1983_),
    .A1(_1978_),
    .A2(_1979_));
 sg13g2_o21ai_1 _5647_ (.B1(_1865_),
    .Y(_1984_),
    .A1(_1804_),
    .A2(_1866_));
 sg13g2_nor2b_1 _5648_ (.A(_1867_),
    .B_N(_1984_),
    .Y(_1985_));
 sg13g2_a21oi_1 _5649_ (.A1(_1983_),
    .A2(_1984_),
    .Y(_1986_),
    .B1(_1867_));
 sg13g2_inv_1 _5650_ (.Y(_1987_),
    .A(_1986_));
 sg13g2_xor2_1 _5651_ (.B(_1807_),
    .A(_1806_),
    .X(_1989_));
 sg13g2_a21oi_2 _5652_ (.B1(_1808_),
    .Y(_1990_),
    .A2(_1989_),
    .A1(_1987_));
 sg13g2_xnor2_1 _5653_ (.Y(_1991_),
    .A(_1749_),
    .B(_1750_));
 sg13g2_o21ai_1 _5654_ (.B1(_1751_),
    .Y(_1992_),
    .A1(_1990_),
    .A2(_1991_));
 sg13g2_o21ai_1 _5655_ (.B1(_1699_),
    .Y(_1993_),
    .A1(_1645_),
    .A2(_1992_));
 sg13g2_a21oi_1 _5656_ (.A1(_1644_),
    .A2(_1697_),
    .Y(_1994_),
    .B1(_1992_));
 sg13g2_mux2_1 _5657_ (.A0(_1698_),
    .A1(_1994_),
    .S(_1993_),
    .X(_1995_));
 sg13g2_a21oi_1 _5658_ (.A1(_1262_),
    .A2(net671),
    .Y(_1996_),
    .B1(net709));
 sg13g2_a21oi_1 _5659_ (.A1(_1262_),
    .A2(net671),
    .Y(_1997_),
    .B1(_1362_));
 sg13g2_xnor2_1 _5660_ (.Y(_1998_),
    .A(net156),
    .B(_1996_));
 sg13g2_nor2_1 _5661_ (.A(net875),
    .B(_1998_),
    .Y(_0051_));
 sg13g2_xnor2_1 _5662_ (.Y(_2000_),
    .A(_1969_),
    .B(_1971_));
 sg13g2_a21oi_1 _5663_ (.A1(net671),
    .A2(_2000_),
    .Y(_2001_),
    .B1(_1351_));
 sg13g2_nand3_1 _5664_ (.B(net671),
    .C(_2000_),
    .A(_1351_),
    .Y(_2002_));
 sg13g2_nor2b_1 _5665_ (.A(_2001_),
    .B_N(_2002_),
    .Y(_2003_));
 sg13g2_xnor2_1 _5666_ (.Y(_2004_),
    .A(_1997_),
    .B(_2003_));
 sg13g2_o21ai_1 _5667_ (.B1(net878),
    .Y(_2005_),
    .A1(net179),
    .A2(net710));
 sg13g2_a21oi_1 _5668_ (.A1(net710),
    .A2(_2004_),
    .Y(_0052_),
    .B1(_2005_));
 sg13g2_a21o_1 _5669_ (.A2(_2002_),
    .A1(_1997_),
    .B1(_2001_),
    .X(_2006_));
 sg13g2_xnor2_1 _5670_ (.Y(_2007_),
    .A(_1972_),
    .B(_1974_));
 sg13g2_and2_1 _5671_ (.A(net671),
    .B(_2007_),
    .X(_2009_));
 sg13g2_xnor2_1 _5672_ (.Y(_2010_),
    .A(\system_inst.neuron.u[2] ),
    .B(_2009_));
 sg13g2_xnor2_1 _5673_ (.Y(_2011_),
    .A(_2006_),
    .B(_2010_));
 sg13g2_o21ai_1 _5674_ (.B1(net878),
    .Y(_2012_),
    .A1(net180),
    .A2(net710));
 sg13g2_a21oi_1 _5675_ (.A1(net710),
    .A2(_2011_),
    .Y(_0053_),
    .B1(_2012_));
 sg13g2_xnor2_1 _5676_ (.Y(_2013_),
    .A(_1975_),
    .B(_1977_));
 sg13g2_nand2b_1 _5677_ (.Y(_2014_),
    .B(net671),
    .A_N(_2013_));
 sg13g2_nand2_1 _5678_ (.Y(_2015_),
    .A(\system_inst.neuron.u[3] ),
    .B(_2014_));
 sg13g2_xor2_1 _5679_ (.B(_2014_),
    .A(\system_inst.neuron.u[3] ),
    .X(_2016_));
 sg13g2_inv_1 _5680_ (.Y(_2017_),
    .A(_2016_));
 sg13g2_nor2_1 _5681_ (.A(_0022_),
    .B(_2009_),
    .Y(_2018_));
 sg13g2_a21oi_1 _5682_ (.A1(_2006_),
    .A2(_2010_),
    .Y(_2019_),
    .B1(_2018_));
 sg13g2_xnor2_1 _5683_ (.Y(_2020_),
    .A(_2017_),
    .B(_2019_));
 sg13g2_o21ai_1 _5684_ (.B1(net878),
    .Y(_2021_),
    .A1(net175),
    .A2(net710));
 sg13g2_a21oi_1 _5685_ (.A1(net710),
    .A2(_2020_),
    .Y(_0054_),
    .B1(_2021_));
 sg13g2_o21ai_1 _5686_ (.B1(_1794_),
    .Y(_2022_),
    .A1(\system_inst.loader.state[4] ),
    .A2(\system_inst.loader.state[0] ));
 sg13g2_nor3_1 _5687_ (.A(\system_inst.loader.state[1] ),
    .B(_1859_),
    .C(_1892_),
    .Y(_2023_));
 sg13g2_o21ai_1 _5688_ (.B1(_2022_),
    .Y(_2024_),
    .A1(net719),
    .A2(_2023_));
 sg13g2_nand2_1 _5689_ (.Y(_2025_),
    .A(_1892_),
    .B(net719));
 sg13g2_a21oi_1 _5690_ (.A1(net146),
    .A2(_2024_),
    .Y(_2026_),
    .B1(net871));
 sg13g2_nand2_1 _5691_ (.Y(_0055_),
    .A(_2025_),
    .B(_2026_));
 sg13g2_nor3_1 _5692_ (.A(\system_inst.loader.shift_reg[2] ),
    .B(\system_inst.loader.shift_reg[1] ),
    .C(net192),
    .Y(_2028_));
 sg13g2_nor4_1 _5693_ (.A(\system_inst.loader.shift_reg[6] ),
    .B(\system_inst.loader.shift_reg[5] ),
    .C(\system_inst.loader.shift_reg[4] ),
    .D(\system_inst.loader.shift_reg[3] ),
    .Y(_2029_));
 sg13g2_a21oi_2 _5694_ (.B1(net12),
    .Y(_2030_),
    .A2(_2029_),
    .A1(net193));
 sg13g2_o21ai_1 _5695_ (.B1(net880),
    .Y(_2031_),
    .A1(net795),
    .A2(net712));
 sg13g2_a21oi_1 _5696_ (.A1(net712),
    .A2(net194),
    .Y(_0056_),
    .B1(_2031_));
 sg13g2_a21oi_1 _5697_ (.A1(net128),
    .A2(net712),
    .Y(_2032_),
    .B1(net874));
 sg13g2_o21ai_1 _5698_ (.B1(_2032_),
    .Y(_0057_),
    .A1(net731),
    .A2(net711));
 sg13g2_o21ai_1 _5699_ (.B1(net879),
    .Y(_2033_),
    .A1(net781),
    .A2(net711));
 sg13g2_a21oi_1 _5700_ (.A1(_1241_),
    .A2(net711),
    .Y(_0058_),
    .B1(_2033_));
 sg13g2_a21oi_1 _5701_ (.A1(net137),
    .A2(net711),
    .Y(_2035_),
    .B1(net874));
 sg13g2_o21ai_1 _5702_ (.B1(_2035_),
    .Y(_0059_),
    .A1(net739),
    .A2(net712));
 sg13g2_a21oi_1 _5703_ (.A1(net149),
    .A2(net713),
    .Y(_2036_),
    .B1(net875));
 sg13g2_o21ai_1 _5704_ (.B1(_2036_),
    .Y(_0060_),
    .A1(net741),
    .A2(net713));
 sg13g2_o21ai_1 _5705_ (.B1(net879),
    .Y(_2037_),
    .A1(net766),
    .A2(net711));
 sg13g2_a21oi_1 _5706_ (.A1(_1219_),
    .A2(net711),
    .Y(_0061_),
    .B1(_2037_));
 sg13g2_o21ai_1 _5707_ (.B1(net879),
    .Y(_2038_),
    .A1(net763),
    .A2(net711));
 sg13g2_a21oi_1 _5708_ (.A1(_1208_),
    .A2(net711),
    .Y(_0062_),
    .B1(_2038_));
 sg13g2_o21ai_1 _5709_ (.B1(net878),
    .Y(_2039_),
    .A1(\system_inst.internal_param_a[7] ),
    .A2(net713));
 sg13g2_a21oi_1 _5710_ (.A1(_1197_),
    .A2(net713),
    .Y(_0063_),
    .B1(_2039_));
 sg13g2_o21ai_1 _5711_ (.B1(net876),
    .Y(_2041_),
    .A1(net163),
    .A2(net714));
 sg13g2_a21oi_1 _5712_ (.A1(net714),
    .A2(_2030_),
    .Y(_0064_),
    .B1(_2041_));
 sg13g2_a21oi_1 _5713_ (.A1(net758),
    .A2(_2034_),
    .Y(_2042_),
    .B1(net875));
 sg13g2_o21ai_1 _5714_ (.B1(_2042_),
    .Y(_0065_),
    .A1(_1252_),
    .A2(_2034_));
 sg13g2_o21ai_1 _5715_ (.B1(net876),
    .Y(_2043_),
    .A1(net755),
    .A2(net715));
 sg13g2_a21oi_1 _5716_ (.A1(_1241_),
    .A2(net714),
    .Y(_0066_),
    .B1(_2043_));
 sg13g2_a21oi_1 _5717_ (.A1(net753),
    .A2(_2034_),
    .Y(_2044_),
    .B1(net875));
 sg13g2_o21ai_1 _5718_ (.B1(_2044_),
    .Y(_0067_),
    .A1(_1230_),
    .A2(_2034_));
 sg13g2_a21oi_1 _5719_ (.A1(net149),
    .A2(net714),
    .Y(_2045_),
    .B1(net875));
 sg13g2_o21ai_1 _5720_ (.B1(_2045_),
    .Y(_0068_),
    .A1(_1296_),
    .A2(net714));
 sg13g2_o21ai_1 _5721_ (.B1(net877),
    .Y(_2046_),
    .A1(net748),
    .A2(net714));
 sg13g2_a21oi_1 _5722_ (.A1(_1219_),
    .A2(net715),
    .Y(_0069_),
    .B1(_2046_));
 sg13g2_o21ai_1 _5723_ (.B1(net876),
    .Y(_2047_),
    .A1(net745),
    .A2(net715));
 sg13g2_a21oi_1 _5724_ (.A1(_1208_),
    .A2(net715),
    .Y(_0070_),
    .B1(_2047_));
 sg13g2_o21ai_1 _5725_ (.B1(net876),
    .Y(_2048_),
    .A1(net743),
    .A2(net714));
 sg13g2_a21oi_1 _5726_ (.A1(_1197_),
    .A2(net714),
    .Y(_0071_),
    .B1(_2048_));
 sg13g2_a21oi_1 _5727_ (.A1(net12),
    .A2(_1988_),
    .Y(_2049_),
    .B1(net871));
 sg13g2_o21ai_1 _5728_ (.B1(_2049_),
    .Y(_0072_),
    .A1(_1285_),
    .A2(_1988_));
 sg13g2_a21oi_1 _5729_ (.A1(net130),
    .A2(net716),
    .Y(_2050_),
    .B1(net872));
 sg13g2_o21ai_1 _5730_ (.B1(_2050_),
    .Y(_0073_),
    .A1(_1252_),
    .A2(net716));
 sg13g2_a21oi_1 _5731_ (.A1(net131),
    .A2(net716),
    .Y(_2052_),
    .B1(net872));
 sg13g2_o21ai_1 _5732_ (.B1(_2052_),
    .Y(_0074_),
    .A1(_1241_),
    .A2(net716));
 sg13g2_a21oi_1 _5733_ (.A1(net117),
    .A2(net716),
    .Y(_2053_),
    .B1(net872));
 sg13g2_o21ai_1 _5734_ (.B1(_2053_),
    .Y(_0075_),
    .A1(_1230_),
    .A2(net716));
 sg13g2_a21oi_1 _5735_ (.A1(\system_inst.loader.shift_reg[3] ),
    .A2(_1988_),
    .Y(_2054_),
    .B1(net872));
 sg13g2_o21ai_1 _5736_ (.B1(_2054_),
    .Y(_0076_),
    .A1(_1274_),
    .A2(_1988_));
 sg13g2_a21oi_1 _5737_ (.A1(net136),
    .A2(_1999_),
    .Y(_2055_),
    .B1(net872));
 sg13g2_o21ai_1 _5738_ (.B1(_2055_),
    .Y(_0077_),
    .A1(_1219_),
    .A2(net716));
 sg13g2_o21ai_1 _5739_ (.B1(net882),
    .Y(_2056_),
    .A1(net126),
    .A2(_1988_));
 sg13g2_a21oi_1 _5740_ (.A1(_1208_),
    .A2(_1988_),
    .Y(_0078_),
    .B1(_2056_));
 sg13g2_o21ai_1 _5741_ (.B1(net876),
    .Y(_2058_),
    .A1(net151),
    .A2(net717));
 sg13g2_a21oi_1 _5742_ (.A1(net717),
    .A2(_2030_),
    .Y(_0079_),
    .B1(_2058_));
 sg13g2_o21ai_1 _5743_ (.B1(net876),
    .Y(_2059_),
    .A1(net155),
    .A2(net717));
 sg13g2_a21oi_1 _5744_ (.A1(_1252_),
    .A2(net717),
    .Y(_0080_),
    .B1(_2059_));
 sg13g2_o21ai_1 _5745_ (.B1(net877),
    .Y(_2060_),
    .A1(net145),
    .A2(net717));
 sg13g2_a21oi_1 _5746_ (.A1(_1241_),
    .A2(net717),
    .Y(_0081_),
    .B1(_2060_));
 sg13g2_o21ai_1 _5747_ (.B1(net876),
    .Y(_2061_),
    .A1(net148),
    .A2(net717));
 sg13g2_a21oi_1 _5748_ (.A1(_1230_),
    .A2(net717),
    .Y(_0082_),
    .B1(_2061_));
 sg13g2_a21oi_1 _5749_ (.A1(\system_inst.loader.shift_reg[3] ),
    .A2(net718),
    .Y(_2062_),
    .B1(net874));
 sg13g2_o21ai_1 _5750_ (.B1(_2062_),
    .Y(_0083_),
    .A1(_1263_),
    .A2(net718));
 sg13g2_o21ai_1 _5751_ (.B1(net881),
    .Y(_2063_),
    .A1(net161),
    .A2(net718));
 sg13g2_a21oi_1 _5752_ (.A1(_1219_),
    .A2(net718),
    .Y(_0084_),
    .B1(_2063_));
 sg13g2_o21ai_1 _5753_ (.B1(net880),
    .Y(_2064_),
    .A1(net144),
    .A2(net719));
 sg13g2_a21oi_1 _5754_ (.A1(_1208_),
    .A2(net719),
    .Y(_0085_),
    .B1(_2064_));
 sg13g2_o21ai_1 _5755_ (.B1(net880),
    .Y(_2065_),
    .A1(net140),
    .A2(net719));
 sg13g2_a21oi_1 _5756_ (.A1(_1197_),
    .A2(_1956_),
    .Y(_0086_),
    .B1(_2065_));
 sg13g2_nor3_1 _5757_ (.A(\system_inst.loader.state[2] ),
    .B(\system_inst.loader.state[3] ),
    .C(_1527_),
    .Y(_2066_));
 sg13g2_a21oi_1 _5758_ (.A1(_1505_),
    .A2(_2066_),
    .Y(_2067_),
    .B1(net11));
 sg13g2_and3_1 _5759_ (.X(_2068_),
    .A(_0035_),
    .B(_1892_),
    .C(_2066_));
 sg13g2_nand2_1 _5760_ (.Y(_2069_),
    .A(net1),
    .B(_2022_));
 sg13g2_nor3_1 _5761_ (.A(_2067_),
    .B(_2068_),
    .C(_2069_),
    .Y(_2071_));
 sg13g2_o21ai_1 _5762_ (.B1(_1892_),
    .Y(_2072_),
    .A1(_0016_),
    .A2(_1848_));
 sg13g2_nand2_2 _5763_ (.Y(_2073_),
    .A(_1505_),
    .B(_2072_));
 sg13g2_nand2_1 _5764_ (.Y(_2074_),
    .A(net12),
    .B(_2073_));
 sg13g2_o21ai_1 _5765_ (.B1(net882),
    .Y(_2075_),
    .A1(net128),
    .A2(net706));
 sg13g2_a21oi_1 _5766_ (.A1(net706),
    .A2(_2074_),
    .Y(_0087_),
    .B1(_2075_));
 sg13g2_nand2_1 _5767_ (.Y(_2076_),
    .A(net128),
    .B(_2073_));
 sg13g2_o21ai_1 _5768_ (.B1(net879),
    .Y(_2077_),
    .A1(\system_inst.loader.shift_reg[1] ),
    .A2(net706));
 sg13g2_a21oi_1 _5769_ (.A1(net706),
    .A2(_2076_),
    .Y(_0088_),
    .B1(_2077_));
 sg13g2_nand2_1 _5770_ (.Y(_2078_),
    .A(net139),
    .B(_2073_));
 sg13g2_o21ai_1 _5771_ (.B1(net879),
    .Y(_2080_),
    .A1(net137),
    .A2(net706));
 sg13g2_a21oi_1 _5772_ (.A1(net706),
    .A2(_2078_),
    .Y(_0089_),
    .B1(_2080_));
 sg13g2_nand2_1 _5773_ (.Y(_2081_),
    .A(net137),
    .B(_2073_));
 sg13g2_o21ai_1 _5774_ (.B1(net880),
    .Y(_2082_),
    .A1(\system_inst.loader.shift_reg[3] ),
    .A2(net706));
 sg13g2_a21oi_1 _5775_ (.A1(net707),
    .A2(_2081_),
    .Y(_0090_),
    .B1(_2082_));
 sg13g2_nand2_1 _5776_ (.Y(_2083_),
    .A(net149),
    .B(_2073_));
 sg13g2_o21ai_1 _5777_ (.B1(net882),
    .Y(_2084_),
    .A1(net121),
    .A2(net707));
 sg13g2_a21oi_1 _5778_ (.A1(net706),
    .A2(_2083_),
    .Y(_0091_),
    .B1(_2084_));
 sg13g2_nand2_1 _5779_ (.Y(_2085_),
    .A(net121),
    .B(_2073_));
 sg13g2_o21ai_1 _5780_ (.B1(net882),
    .Y(_2086_),
    .A1(net119),
    .A2(net707));
 sg13g2_a21oi_1 _5781_ (.A1(net707),
    .A2(_2085_),
    .Y(_0092_),
    .B1(_2086_));
 sg13g2_nand2_1 _5782_ (.Y(_2088_),
    .A(net119),
    .B(_2073_));
 sg13g2_o21ai_1 _5783_ (.B1(net879),
    .Y(_2089_),
    .A1(\system_inst.loader.shift_reg[6] ),
    .A2(net707));
 sg13g2_a21oi_1 _5784_ (.A1(net707),
    .A2(_2088_),
    .Y(_0093_),
    .B1(_2089_));
 sg13g2_a21oi_1 _5785_ (.A1(_2024_),
    .A2(net708),
    .Y(_2090_),
    .B1(net111));
 sg13g2_a21oi_1 _5786_ (.A1(net111),
    .A2(net708),
    .Y(_2091_),
    .B1(net871));
 sg13g2_nor2b_1 _5787_ (.A(_2090_),
    .B_N(_2091_),
    .Y(_0094_));
 sg13g2_a21oi_1 _5788_ (.A1(\system_inst.loader.bit_count[0] ),
    .A2(net708),
    .Y(_2092_),
    .B1(net105));
 sg13g2_o21ai_1 _5789_ (.B1(_1848_),
    .Y(_2093_),
    .A1(\system_inst.loader.state[1] ),
    .A2(_1892_));
 sg13g2_a21oi_1 _5790_ (.A1(net708),
    .A2(_2093_),
    .Y(_2094_),
    .B1(net871));
 sg13g2_nor2b_1 _5791_ (.A(net106),
    .B_N(_2094_),
    .Y(_0095_));
 sg13g2_xor2_1 _5792_ (.B(_1848_),
    .A(_0016_),
    .X(_2096_));
 sg13g2_o21ai_1 _5793_ (.B1(_2096_),
    .Y(_2097_),
    .A1(\system_inst.loader.state[1] ),
    .A2(_1892_));
 sg13g2_o21ai_1 _5794_ (.B1(net882),
    .Y(_2098_),
    .A1(net113),
    .A2(net708));
 sg13g2_a21oi_1 _5795_ (.A1(net708),
    .A2(_2097_),
    .Y(_0096_),
    .B1(_2098_));
 sg13g2_o21ai_1 _5796_ (.B1(_2015_),
    .Y(_2099_),
    .A1(_2017_),
    .A2(_2019_));
 sg13g2_xnor2_1 _5797_ (.Y(_2100_),
    .A(_1978_),
    .B(_1982_));
 sg13g2_nand2b_1 _5798_ (.Y(_2101_),
    .B(net671),
    .A_N(_2100_));
 sg13g2_inv_1 _5799_ (.Y(_2102_),
    .A(_2101_));
 sg13g2_xor2_1 _5800_ (.B(_2101_),
    .A(\system_inst.neuron.u[4] ),
    .X(_2103_));
 sg13g2_nand2_1 _5801_ (.Y(_2105_),
    .A(_2099_),
    .B(_2103_));
 sg13g2_o21ai_1 _5802_ (.B1(net720),
    .Y(_2106_),
    .A1(_2099_),
    .A2(_2103_));
 sg13g2_nand2b_1 _5803_ (.Y(_2107_),
    .B(_2105_),
    .A_N(_2106_));
 sg13g2_nand2_1 _5804_ (.Y(_2108_),
    .A(\system_inst.neuron.u[4] ),
    .B(net151));
 sg13g2_xor2_1 _5805_ (.B(net151),
    .A(\system_inst.neuron.u[4] ),
    .X(_2109_));
 sg13g2_o21ai_1 _5806_ (.B1(net709),
    .Y(_2110_),
    .A1(net725),
    .A2(_2109_));
 sg13g2_o21ai_1 _5807_ (.B1(net878),
    .Y(_2111_),
    .A1(net190),
    .A2(net726));
 sg13g2_a21oi_1 _5808_ (.A1(_2107_),
    .A2(_2110_),
    .Y(_0097_),
    .B1(_2111_));
 sg13g2_o21ai_1 _5809_ (.B1(_2105_),
    .Y(_2112_),
    .A1(_0015_),
    .A2(_2102_));
 sg13g2_xnor2_1 _5810_ (.Y(_2113_),
    .A(_1983_),
    .B(_1985_));
 sg13g2_a21oi_1 _5811_ (.A1(net672),
    .A2(_2113_),
    .Y(_2115_),
    .B1(_1186_));
 sg13g2_and3_1 _5812_ (.X(_2116_),
    .A(_1186_),
    .B(net672),
    .C(_2113_));
 sg13g2_nor2_1 _5813_ (.A(_2115_),
    .B(_2116_),
    .Y(_2117_));
 sg13g2_xnor2_1 _5814_ (.Y(_2118_),
    .A(_2112_),
    .B(_2117_));
 sg13g2_xnor2_1 _5815_ (.Y(_2119_),
    .A(\system_inst.neuron.u[5] ),
    .B(\system_inst.internal_param_d[1] ));
 sg13g2_nor2_1 _5816_ (.A(_2108_),
    .B(_2119_),
    .Y(_2120_));
 sg13g2_xnor2_1 _5817_ (.Y(_2121_),
    .A(_2108_),
    .B(_2119_));
 sg13g2_o21ai_1 _5818_ (.B1(net876),
    .Y(_2122_),
    .A1(net186),
    .A2(net726));
 sg13g2_a221oi_1 _5819_ (.B2(_2087_),
    .C1(_2122_),
    .B1(_2121_),
    .A1(net710),
    .Y(_0098_),
    .A2(_2118_));
 sg13g2_xnor2_1 _5820_ (.Y(_2123_),
    .A(\system_inst.neuron.u[6] ),
    .B(\system_inst.internal_param_d[2] ));
 sg13g2_a21oi_1 _5821_ (.A1(\system_inst.neuron.u[5] ),
    .A2(\system_inst.internal_param_d[1] ),
    .Y(_2125_),
    .B1(_2120_));
 sg13g2_nor2_1 _5822_ (.A(_2123_),
    .B(_2125_),
    .Y(_2126_));
 sg13g2_a21o_1 _5823_ (.A2(_2125_),
    .A1(_2123_),
    .B1(net720),
    .X(_2127_));
 sg13g2_o21ai_1 _5824_ (.B1(net726),
    .Y(_2128_),
    .A1(_2126_),
    .A2(_2127_));
 sg13g2_a221oi_1 _5825_ (.B2(_2099_),
    .C1(_2115_),
    .B1(_2103_),
    .A1(_1461_),
    .Y(_2129_),
    .A2(_2101_));
 sg13g2_xnor2_1 _5826_ (.Y(_2130_),
    .A(_1987_),
    .B(_1989_));
 sg13g2_nand2_1 _5827_ (.Y(_2131_),
    .A(net672),
    .B(_2130_));
 sg13g2_xnor2_1 _5828_ (.Y(_2132_),
    .A(\system_inst.neuron.u[6] ),
    .B(_2131_));
 sg13g2_nor3_2 _5829_ (.A(_2116_),
    .B(_2129_),
    .C(_2132_),
    .Y(_2133_));
 sg13g2_o21ai_1 _5830_ (.B1(_2132_),
    .Y(_2134_),
    .A1(_2116_),
    .A2(_2129_));
 sg13g2_nand2_1 _5831_ (.Y(_2136_),
    .A(net720),
    .B(_2134_));
 sg13g2_nor2_1 _5832_ (.A(_2133_),
    .B(_2136_),
    .Y(_2137_));
 sg13g2_o21ai_1 _5833_ (.B1(net877),
    .Y(_2138_),
    .A1(_2128_),
    .A2(_2137_));
 sg13g2_a21oi_1 _5834_ (.A1(_1175_),
    .A2(net725),
    .Y(_0099_),
    .B1(_2138_));
 sg13g2_a21oi_1 _5835_ (.A1(net672),
    .A2(_2130_),
    .Y(_2139_),
    .B1(_0013_));
 sg13g2_xnor2_1 _5836_ (.Y(_2140_),
    .A(_1990_),
    .B(_1991_));
 sg13g2_nand2_1 _5837_ (.Y(_2141_),
    .A(net671),
    .B(_2140_));
 sg13g2_nand2_1 _5838_ (.Y(_2142_),
    .A(\system_inst.neuron.u[7] ),
    .B(_2141_));
 sg13g2_xor2_1 _5839_ (.B(_2141_),
    .A(\system_inst.neuron.u[7] ),
    .X(_2143_));
 sg13g2_or3_1 _5840_ (.A(_2133_),
    .B(_2139_),
    .C(_2143_),
    .X(_2144_));
 sg13g2_o21ai_1 _5841_ (.B1(_2143_),
    .Y(_2146_),
    .A1(_2133_),
    .A2(_2139_));
 sg13g2_nand3_1 _5842_ (.B(_2144_),
    .C(_2146_),
    .A(net720),
    .Y(_2147_));
 sg13g2_xnor2_1 _5843_ (.Y(_2148_),
    .A(\system_inst.neuron.u[7] ),
    .B(\system_inst.internal_param_d[3] ));
 sg13g2_a21oi_1 _5844_ (.A1(\system_inst.neuron.u[6] ),
    .A2(\system_inst.internal_param_d[2] ),
    .Y(_2149_),
    .B1(_2126_));
 sg13g2_nor2_1 _5845_ (.A(_2148_),
    .B(_2149_),
    .Y(_2150_));
 sg13g2_xor2_1 _5846_ (.B(_2149_),
    .A(_2148_),
    .X(_2151_));
 sg13g2_o21ai_1 _5847_ (.B1(net709),
    .Y(_2152_),
    .A1(net725),
    .A2(_2151_));
 sg13g2_o21ai_1 _5848_ (.B1(net877),
    .Y(_2153_),
    .A1(net188),
    .A2(net726));
 sg13g2_a21oi_1 _5849_ (.A1(_2147_),
    .A2(_2152_),
    .Y(_0100_),
    .B1(_2153_));
 sg13g2_a21oi_1 _5850_ (.A1(_2142_),
    .A2(_2146_),
    .Y(_2154_),
    .B1(_0011_));
 sg13g2_nand3_1 _5851_ (.B(_2142_),
    .C(_2146_),
    .A(_0011_),
    .Y(_2156_));
 sg13g2_nor2b_1 _5852_ (.A(_2154_),
    .B_N(_2156_),
    .Y(_2157_));
 sg13g2_xnor2_1 _5853_ (.Y(_2158_),
    .A(\system_inst.neuron.u[8] ),
    .B(\system_inst.internal_param_d[4] ));
 sg13g2_a21oi_1 _5854_ (.A1(\system_inst.neuron.u[7] ),
    .A2(\system_inst.internal_param_d[3] ),
    .Y(_2159_),
    .B1(_2150_));
 sg13g2_nor2_1 _5855_ (.A(_2158_),
    .B(_2159_),
    .Y(_2160_));
 sg13g2_nand2_1 _5856_ (.Y(_2161_),
    .A(_2158_),
    .B(_2159_));
 sg13g2_nor2_1 _5857_ (.A(net722),
    .B(_2160_),
    .Y(_2162_));
 sg13g2_a221oi_1 _5858_ (.B2(_2162_),
    .C1(net725),
    .B1(_2161_),
    .A1(net722),
    .Y(_2163_),
    .A2(_2157_));
 sg13g2_o21ai_1 _5859_ (.B1(net877),
    .Y(_2164_),
    .A1(net185),
    .A2(net727));
 sg13g2_nor2_1 _5860_ (.A(_2163_),
    .B(_2164_),
    .Y(_0101_));
 sg13g2_xnor2_1 _5861_ (.Y(_2166_),
    .A(net177),
    .B(_2154_));
 sg13g2_nor2_1 _5862_ (.A(net709),
    .B(_2166_),
    .Y(_2167_));
 sg13g2_a21oi_2 _5863_ (.B1(_2160_),
    .Y(_2168_),
    .A2(net122),
    .A1(\system_inst.neuron.u[8] ));
 sg13g2_nand2_1 _5864_ (.Y(_2169_),
    .A(\system_inst.neuron.u[9] ),
    .B(\system_inst.internal_param_d[5] ));
 sg13g2_nor2_1 _5865_ (.A(\system_inst.neuron.u[9] ),
    .B(\system_inst.internal_param_d[5] ),
    .Y(_2170_));
 sg13g2_xor2_1 _5866_ (.B(net161),
    .A(\system_inst.neuron.u[9] ),
    .X(_2171_));
 sg13g2_o21ai_1 _5867_ (.B1(_2087_),
    .Y(_2172_),
    .A1(_2168_),
    .A2(_2171_));
 sg13g2_a21oi_1 _5868_ (.A1(_2168_),
    .A2(_2171_),
    .Y(_2173_),
    .B1(_2172_));
 sg13g2_o21ai_1 _5869_ (.B1(net881),
    .Y(_2174_),
    .A1(\system_inst.neuron.u[9] ),
    .A2(net726));
 sg13g2_nor3_1 _5870_ (.A(_2167_),
    .B(_2173_),
    .C(_2174_),
    .Y(_0102_));
 sg13g2_nand2_1 _5871_ (.Y(_2176_),
    .A(\system_inst.neuron.u[9] ),
    .B(\system_inst.neuron.u[8] ));
 sg13g2_a21oi_2 _5872_ (.B1(_2176_),
    .Y(_2177_),
    .A2(_2146_),
    .A1(_2142_));
 sg13g2_nor2b_1 _5873_ (.A(_0009_),
    .B_N(_2177_),
    .Y(_2178_));
 sg13g2_xnor2_1 _5874_ (.Y(_2179_),
    .A(_0009_),
    .B(_2177_));
 sg13g2_xor2_1 _5875_ (.B(\system_inst.internal_param_d[6] ),
    .A(\system_inst.neuron.u[10] ),
    .X(_2180_));
 sg13g2_o21ai_1 _5876_ (.B1(_2169_),
    .Y(_2181_),
    .A1(_2168_),
    .A2(_2170_));
 sg13g2_and2_1 _5877_ (.A(_2180_),
    .B(_2181_),
    .X(_2182_));
 sg13g2_or2_1 _5878_ (.X(_2183_),
    .B(_2181_),
    .A(_2180_));
 sg13g2_nor2_1 _5879_ (.A(net721),
    .B(_2182_),
    .Y(_2184_));
 sg13g2_a221oi_1 _5880_ (.B2(_2184_),
    .C1(net725),
    .B1(_2183_),
    .A1(net721),
    .Y(_2185_),
    .A2(_2179_));
 sg13g2_o21ai_1 _5881_ (.B1(net881),
    .Y(_2187_),
    .A1(net189),
    .A2(net727));
 sg13g2_nor2_1 _5882_ (.A(_2185_),
    .B(_2187_),
    .Y(_0103_));
 sg13g2_xnor2_1 _5883_ (.Y(_2188_),
    .A(_0008_),
    .B(_2178_));
 sg13g2_xor2_1 _5884_ (.B(\system_inst.internal_param_d[7] ),
    .A(\system_inst.neuron.u[11] ),
    .X(_2189_));
 sg13g2_a21o_1 _5885_ (.A2(\system_inst.internal_param_d[6] ),
    .A1(\system_inst.neuron.u[10] ),
    .B1(_2182_),
    .X(_2190_));
 sg13g2_and2_1 _5886_ (.A(_2189_),
    .B(_2190_),
    .X(_2191_));
 sg13g2_nor2_1 _5887_ (.A(_2189_),
    .B(_2190_),
    .Y(_2192_));
 sg13g2_nor3_1 _5888_ (.A(net721),
    .B(_2191_),
    .C(_2192_),
    .Y(_2193_));
 sg13g2_a21oi_1 _5889_ (.A1(net721),
    .A2(_2188_),
    .Y(_2194_),
    .B1(_2193_));
 sg13g2_o21ai_1 _5890_ (.B1(net879),
    .Y(_2195_),
    .A1(net183),
    .A2(_2070_));
 sg13g2_a21oi_1 _5891_ (.A1(_2070_),
    .A2(_2194_),
    .Y(_0104_),
    .B1(_2195_));
 sg13g2_nand3_1 _5892_ (.B(\system_inst.neuron.u[10] ),
    .C(_2177_),
    .A(\system_inst.neuron.u[11] ),
    .Y(_2197_));
 sg13g2_a21o_1 _5893_ (.A2(\system_inst.internal_param_d[7] ),
    .A1(\system_inst.neuron.u[11] ),
    .B1(_2191_),
    .X(_2198_));
 sg13g2_nor2_1 _5894_ (.A(net720),
    .B(_2198_),
    .Y(_2199_));
 sg13g2_a21oi_1 _5895_ (.A1(net720),
    .A2(_2197_),
    .Y(_2200_),
    .B1(_2199_));
 sg13g2_xnor2_1 _5896_ (.Y(_2201_),
    .A(_1483_),
    .B(_2200_));
 sg13g2_o21ai_1 _5897_ (.B1(net877),
    .Y(_2202_),
    .A1(\system_inst.neuron.u[12] ),
    .A2(net726));
 sg13g2_a21oi_1 _5898_ (.A1(net726),
    .A2(_2201_),
    .Y(_0105_),
    .B1(_2202_));
 sg13g2_nand4_1 _5899_ (.B(\system_inst.neuron.u[10] ),
    .C(_1483_),
    .A(\system_inst.neuron.u[11] ),
    .Y(_2203_),
    .D(_2177_));
 sg13g2_xnor2_1 _5900_ (.Y(_2204_),
    .A(_1494_),
    .B(_2203_));
 sg13g2_a21oi_1 _5901_ (.A1(\system_inst.neuron.u[12] ),
    .A2(_2198_),
    .Y(_2206_),
    .B1(net742));
 sg13g2_nand3_1 _5902_ (.B(net191),
    .C(_2198_),
    .A(net742),
    .Y(_2207_));
 sg13g2_nor2_1 _5903_ (.A(net722),
    .B(_2206_),
    .Y(_2208_));
 sg13g2_a221oi_1 _5904_ (.B2(_2208_),
    .C1(net725),
    .B1(_2207_),
    .A1(net720),
    .Y(_2209_),
    .A2(_2204_));
 sg13g2_o21ai_1 _5905_ (.B1(net879),
    .Y(_2210_),
    .A1(net742),
    .A2(net726));
 sg13g2_nor2_1 _5906_ (.A(_2209_),
    .B(_2210_),
    .Y(_0106_));
 sg13g2_nor3_1 _5907_ (.A(net873),
    .B(net721),
    .C(_2079_),
    .Y(_0107_));
 sg13g2_dfrbp_1 _5908_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net93),
    .D(_0036_),
    .Q_N(_0033_),
    .Q(\system_inst.neuron.membrane_scaled[1] ));
 sg13g2_dfrbp_1 _5909_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net72),
    .D(_0037_),
    .Q_N(_0032_),
    .Q(\system_inst.neuron.membrane_scaled[2] ));
 sg13g2_dfrbp_1 _5910_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net70),
    .D(_0038_),
    .Q_N(_0031_),
    .Q(\system_inst.neuron.membrane_scaled[3] ));
 sg13g2_dfrbp_1 _5911_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net68),
    .D(_0039_),
    .Q_N(_0030_),
    .Q(\system_inst.neuron.membrane_scaled[4] ));
 sg13g2_dfrbp_1 _5912_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net66),
    .D(_0040_),
    .Q_N(_0029_),
    .Q(\system_inst.neuron.membrane_scaled[5] ));
 sg13g2_dfrbp_1 _5913_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net64),
    .D(_0041_),
    .Q_N(_0028_),
    .Q(\system_inst.neuron.membrane_scaled[6] ));
 sg13g2_dfrbp_1 _5914_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net62),
    .D(_0042_),
    .Q_N(_0027_),
    .Q(\system_inst.neuron.membrane_scaled[7] ));
 sg13g2_dfrbp_1 _5915_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net60),
    .D(_0043_),
    .Q_N(_2945_),
    .Q(\system_inst.neuron.membrane_scaled[8] ));
 sg13g2_dfrbp_1 _5916_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net58),
    .D(_0044_),
    .Q_N(_2944_),
    .Q(\system_inst.neuron.v[8] ));
 sg13g2_dfrbp_1 _5917_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net56),
    .D(_0045_),
    .Q_N(_0026_),
    .Q(\system_inst.neuron.v[9] ));
 sg13g2_dfrbp_1 _5918_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net54),
    .D(_0046_),
    .Q_N(_0025_),
    .Q(\system_inst.neuron.v[10] ));
 sg13g2_dfrbp_1 _5919_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net52),
    .D(_0047_),
    .Q_N(_2943_),
    .Q(\system_inst.neuron.v[11] ));
 sg13g2_dfrbp_1 _5920_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net50),
    .D(_0048_),
    .Q_N(_0024_),
    .Q(\system_inst.neuron.v[12] ));
 sg13g2_dfrbp_1 _5921_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net48),
    .D(_0049_),
    .Q_N(_0023_),
    .Q(\system_inst.neuron.v[13] ));
 sg13g2_dfrbp_1 _5922_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net46),
    .D(_0050_),
    .Q_N(_2942_),
    .Q(\system_inst.loader.load_enable_prev ));
 sg13g2_dfrbp_1 _5923_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net45),
    .D(_0051_),
    .Q_N(_2941_),
    .Q(\system_inst.neuron.u[0] ));
 sg13g2_dfrbp_1 _5924_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net43),
    .D(_0052_),
    .Q_N(_2940_),
    .Q(\system_inst.neuron.u[1] ));
 sg13g2_dfrbp_1 _5925_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net41),
    .D(_0053_),
    .Q_N(_0022_),
    .Q(\system_inst.neuron.u[2] ));
 sg13g2_dfrbp_1 _5926_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net39),
    .D(net176),
    .Q_N(_0021_),
    .Q(\system_inst.neuron.u[3] ));
 sg13g2_dfrbp_1 _5927_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net37),
    .D(net147),
    .Q_N(_2939_),
    .Q(params_ready_internal));
 sg13g2_dfrbp_1 _5928_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net35),
    .D(_0056_),
    .Q_N(_2938_),
    .Q(\system_inst.internal_param_a[0] ));
 sg13g2_dfrbp_1 _5929_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net33),
    .D(_0057_),
    .Q_N(_2937_),
    .Q(\system_inst.internal_param_a[1] ));
 sg13g2_dfrbp_1 _5930_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net31),
    .D(_0058_),
    .Q_N(_2936_),
    .Q(\system_inst.internal_param_a[2] ));
 sg13g2_dfrbp_1 _5931_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net29),
    .D(_0059_),
    .Q_N(_2935_),
    .Q(\system_inst.internal_param_a[3] ));
 sg13g2_dfrbp_1 _5932_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net27),
    .D(_0060_),
    .Q_N(_0020_),
    .Q(\system_inst.internal_param_a[4] ));
 sg13g2_dfrbp_1 _5933_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net25),
    .D(_0061_),
    .Q_N(_2934_),
    .Q(\system_inst.internal_param_a[5] ));
 sg13g2_dfrbp_1 _5934_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net23),
    .D(_0062_),
    .Q_N(_2933_),
    .Q(\system_inst.internal_param_a[6] ));
 sg13g2_dfrbp_1 _5935_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net99),
    .D(net143),
    .Q_N(_0019_),
    .Q(\system_inst.internal_param_a[7] ));
 sg13g2_dfrbp_1 _5936_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net91),
    .D(net164),
    .Q_N(_2932_),
    .Q(\system_inst.internal_param_b[0] ));
 sg13g2_dfrbp_1 _5937_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net89),
    .D(net154),
    .Q_N(_2931_),
    .Q(\system_inst.internal_param_b[1] ));
 sg13g2_dfrbp_1 _5938_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net87),
    .D(_0066_),
    .Q_N(_2930_),
    .Q(\system_inst.internal_param_b[2] ));
 sg13g2_dfrbp_1 _5939_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net85),
    .D(_0067_),
    .Q_N(_2929_),
    .Q(\system_inst.internal_param_b[3] ));
 sg13g2_dfrbp_1 _5940_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net83),
    .D(_0068_),
    .Q_N(_2928_),
    .Q(\system_inst.internal_param_b[4] ));
 sg13g2_dfrbp_1 _5941_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net81),
    .D(_0069_),
    .Q_N(_2927_),
    .Q(\system_inst.internal_param_b[5] ));
 sg13g2_dfrbp_1 _5942_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net79),
    .D(_0070_),
    .Q_N(_2926_),
    .Q(\system_inst.internal_param_b[6] ));
 sg13g2_dfrbp_1 _5943_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net77),
    .D(_0071_),
    .Q_N(_2925_),
    .Q(\system_inst.internal_param_b[7] ));
 sg13g2_dfrbp_1 _5944_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net75),
    .D(_0072_),
    .Q_N(_2924_),
    .Q(\system_inst.internal_param_c[0] ));
 sg13g2_dfrbp_1 _5945_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net73),
    .D(_0073_),
    .Q_N(_0018_),
    .Q(\system_inst.internal_param_c[1] ));
 sg13g2_dfrbp_1 _5946_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net69),
    .D(net132),
    .Q_N(_2923_),
    .Q(\system_inst.internal_param_c[2] ));
 sg13g2_dfrbp_1 _5947_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net65),
    .D(net118),
    .Q_N(_0017_),
    .Q(\system_inst.internal_param_c[3] ));
 sg13g2_dfrbp_1 _5948_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net61),
    .D(net125),
    .Q_N(_2922_),
    .Q(\system_inst.internal_param_c[4] ));
 sg13g2_dfrbp_1 _5949_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net57),
    .D(_0077_),
    .Q_N(_2921_),
    .Q(\system_inst.internal_param_c[5] ));
 sg13g2_dfrbp_1 _5950_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net53),
    .D(_0078_),
    .Q_N(_2920_),
    .Q(\system_inst.internal_param_c[6] ));
 sg13g2_dfrbp_1 _5951_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net49),
    .D(net152),
    .Q_N(_2919_),
    .Q(\system_inst.internal_param_d[0] ));
 sg13g2_dfrbp_1 _5952_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net44),
    .D(_0080_),
    .Q_N(_2918_),
    .Q(\system_inst.internal_param_d[1] ));
 sg13g2_dfrbp_1 _5953_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net40),
    .D(_0081_),
    .Q_N(_2917_),
    .Q(\system_inst.internal_param_d[2] ));
 sg13g2_dfrbp_1 _5954_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net36),
    .D(_0082_),
    .Q_N(_2916_),
    .Q(\system_inst.internal_param_d[3] ));
 sg13g2_dfrbp_1 _5955_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net32),
    .D(net123),
    .Q_N(_2915_),
    .Q(\system_inst.internal_param_d[4] ));
 sg13g2_dfrbp_1 _5956_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net28),
    .D(_0084_),
    .Q_N(_2914_),
    .Q(\system_inst.internal_param_d[5] ));
 sg13g2_dfrbp_1 _5957_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net24),
    .D(_0085_),
    .Q_N(_2913_),
    .Q(\system_inst.internal_param_d[6] ));
 sg13g2_dfrbp_1 _5958_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net92),
    .D(net141),
    .Q_N(_2912_),
    .Q(\system_inst.internal_param_d[7] ));
 sg13g2_dfrbp_1 _5959_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net88),
    .D(_0087_),
    .Q_N(_2911_),
    .Q(\system_inst.loader.shift_reg[0] ));
 sg13g2_dfrbp_1 _5960_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net84),
    .D(net129),
    .Q_N(_2910_),
    .Q(\system_inst.loader.shift_reg[1] ));
 sg13g2_dfrbp_1 _5961_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net80),
    .D(_0089_),
    .Q_N(_2909_),
    .Q(\system_inst.loader.shift_reg[2] ));
 sg13g2_dfrbp_1 _5962_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net76),
    .D(net138),
    .Q_N(_2908_),
    .Q(\system_inst.loader.shift_reg[3] ));
 sg13g2_dfrbp_1 _5963_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net71),
    .D(_0091_),
    .Q_N(_2907_),
    .Q(\system_inst.loader.shift_reg[4] ));
 sg13g2_dfrbp_1 _5964_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net63),
    .D(_0092_),
    .Q_N(_2906_),
    .Q(\system_inst.loader.shift_reg[5] ));
 sg13g2_dfrbp_1 _5965_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net55),
    .D(net120),
    .Q_N(_2905_),
    .Q(\system_inst.loader.shift_reg[6] ));
 sg13g2_dfrbp_1 _5966_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net47),
    .D(_0094_),
    .Q_N(_2904_),
    .Q(\system_inst.loader.bit_count[0] ));
 sg13g2_dfrbp_1 _5967_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net38),
    .D(net107),
    .Q_N(_2903_),
    .Q(\system_inst.loader.bit_count[1] ));
 sg13g2_dfrbp_1 _5968_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net30),
    .D(net114),
    .Q_N(_0016_),
    .Q(\system_inst.loader.bit_count[2] ));
 sg13g2_dfrbp_1 _5969_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net22),
    .D(_0097_),
    .Q_N(_0015_),
    .Q(\system_inst.neuron.u[4] ));
 sg13g2_dfrbp_1 _5970_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net86),
    .D(net187),
    .Q_N(_0014_),
    .Q(\system_inst.neuron.u[5] ));
 sg13g2_dfrbp_1 _5971_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net78),
    .D(_0099_),
    .Q_N(_0013_),
    .Q(\system_inst.neuron.u[6] ));
 sg13g2_dfrbp_1 _5972_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net67),
    .D(_0100_),
    .Q_N(_0012_),
    .Q(\system_inst.neuron.u[7] ));
 sg13g2_dfrbp_1 _5973_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net51),
    .D(_0101_),
    .Q_N(_0011_),
    .Q(\system_inst.neuron.u[8] ));
 sg13g2_dfrbp_1 _5974_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net34),
    .D(net178),
    .Q_N(_0010_),
    .Q(\system_inst.neuron.u[9] ));
 sg13g2_dfrbp_1 _5975_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net90),
    .D(_0103_),
    .Q_N(_0009_),
    .Q(\system_inst.neuron.u[10] ));
 sg13g2_dfrbp_1 _5976_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net74),
    .D(net184),
    .Q_N(_0008_),
    .Q(\system_inst.neuron.u[11] ));
 sg13g2_dfrbp_1 _5977_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net42),
    .D(net158),
    .Q_N(_0007_),
    .Q(\system_inst.neuron.u[12] ));
 sg13g2_dfrbp_1 _5978_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net94),
    .D(_0106_),
    .Q_N(_0034_),
    .Q(\system_inst.neuron.u[13] ));
 sg13g2_dfrbp_1 _5979_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net95),
    .D(_0000_),
    .Q_N(_2946_),
    .Q(\system_inst.loader.state[0] ));
 sg13g2_dfrbp_1 _5980_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net96),
    .D(_0001_),
    .Q_N(_0035_),
    .Q(\system_inst.loader.state[1] ));
 sg13g2_dfrbp_1 _5981_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net97),
    .D(_0002_),
    .Q_N(_2947_),
    .Q(\system_inst.loader.state[2] ));
 sg13g2_dfrbp_1 _5982_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net98),
    .D(_0003_),
    .Q_N(_2948_),
    .Q(\system_inst.loader.state[3] ));
 sg13g2_dfrbp_1 _5983_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net59),
    .D(_0004_),
    .Q_N(_2949_),
    .Q(\system_inst.loader.state[4] ));
 sg13g2_dfrbp_1 _5984_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net82),
    .D(net109),
    .Q_N(_0006_),
    .Q(\system_inst.loader.state[5] ));
 sg13g2_dfrbp_1 _5985_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net26),
    .D(_0107_),
    .Q_N(_2902_),
    .Q(spike_out_internal));
 sg13g2_tiehi _5934__23 (.L_HI(net23));
 sg13g2_tiehi _5957__24 (.L_HI(net24));
 sg13g2_tiehi _5933__25 (.L_HI(net25));
 sg13g2_tiehi _5985__26 (.L_HI(net26));
 sg13g2_tiehi _5932__27 (.L_HI(net27));
 sg13g2_tiehi _5956__28 (.L_HI(net28));
 sg13g2_tiehi _5931__29 (.L_HI(net29));
 sg13g2_tiehi _5968__30 (.L_HI(net30));
 sg13g2_tiehi _5930__31 (.L_HI(net31));
 sg13g2_tiehi _5955__32 (.L_HI(net32));
 sg13g2_tiehi _5929__33 (.L_HI(net33));
 sg13g2_tiehi _5974__34 (.L_HI(net34));
 sg13g2_tiehi _5928__35 (.L_HI(net35));
 sg13g2_tiehi _5954__36 (.L_HI(net36));
 sg13g2_tiehi _5927__37 (.L_HI(net37));
 sg13g2_tiehi _5967__38 (.L_HI(net38));
 sg13g2_tiehi _5926__39 (.L_HI(net39));
 sg13g2_tiehi _5953__40 (.L_HI(net40));
 sg13g2_tiehi _5925__41 (.L_HI(net41));
 sg13g2_tiehi _5977__42 (.L_HI(net42));
 sg13g2_tiehi _5924__43 (.L_HI(net43));
 sg13g2_tiehi _5952__44 (.L_HI(net44));
 sg13g2_tiehi _5923__45 (.L_HI(net45));
 sg13g2_tiehi _5922__46 (.L_HI(net46));
 sg13g2_tiehi _5966__47 (.L_HI(net47));
 sg13g2_tiehi _5921__48 (.L_HI(net48));
 sg13g2_tiehi _5951__49 (.L_HI(net49));
 sg13g2_tiehi _5920__50 (.L_HI(net50));
 sg13g2_tiehi _5973__51 (.L_HI(net51));
 sg13g2_tiehi _5919__52 (.L_HI(net52));
 sg13g2_tiehi _5950__53 (.L_HI(net53));
 sg13g2_tiehi _5918__54 (.L_HI(net54));
 sg13g2_tiehi _5965__55 (.L_HI(net55));
 sg13g2_tiehi _5917__56 (.L_HI(net56));
 sg13g2_tiehi _5949__57 (.L_HI(net57));
 sg13g2_tiehi _5916__58 (.L_HI(net58));
 sg13g2_tiehi _5983__59 (.L_HI(net59));
 sg13g2_tiehi _5915__60 (.L_HI(net60));
 sg13g2_tiehi _5948__61 (.L_HI(net61));
 sg13g2_tiehi _5914__62 (.L_HI(net62));
 sg13g2_tiehi _5964__63 (.L_HI(net63));
 sg13g2_tiehi _5913__64 (.L_HI(net64));
 sg13g2_tiehi _5947__65 (.L_HI(net65));
 sg13g2_tiehi _5912__66 (.L_HI(net66));
 sg13g2_tiehi _5972__67 (.L_HI(net67));
 sg13g2_tiehi _5911__68 (.L_HI(net68));
 sg13g2_tiehi _5946__69 (.L_HI(net69));
 sg13g2_tiehi _5910__70 (.L_HI(net70));
 sg13g2_tiehi _5963__71 (.L_HI(net71));
 sg13g2_tiehi _5909__72 (.L_HI(net72));
 sg13g2_tiehi _5945__73 (.L_HI(net73));
 sg13g2_tiehi _5976__74 (.L_HI(net74));
 sg13g2_tiehi _5944__75 (.L_HI(net75));
 sg13g2_tiehi _5962__76 (.L_HI(net76));
 sg13g2_tiehi _5943__77 (.L_HI(net77));
 sg13g2_tiehi _5971__78 (.L_HI(net78));
 sg13g2_tiehi _5942__79 (.L_HI(net79));
 sg13g2_tiehi _5961__80 (.L_HI(net80));
 sg13g2_tiehi _5941__81 (.L_HI(net81));
 sg13g2_tiehi _5984__82 (.L_HI(net82));
 sg13g2_tiehi _5940__83 (.L_HI(net83));
 sg13g2_tiehi _5960__84 (.L_HI(net84));
 sg13g2_tiehi _5939__85 (.L_HI(net85));
 sg13g2_tiehi _5970__86 (.L_HI(net86));
 sg13g2_tiehi _5938__87 (.L_HI(net87));
 sg13g2_tiehi _5959__88 (.L_HI(net88));
 sg13g2_tiehi _5937__89 (.L_HI(net89));
 sg13g2_tiehi _5975__90 (.L_HI(net90));
 sg13g2_tiehi _5936__91 (.L_HI(net91));
 sg13g2_tiehi _5958__92 (.L_HI(net92));
 sg13g2_tiehi _5908__93 (.L_HI(net93));
 sg13g2_tiehi _5978__94 (.L_HI(net94));
 sg13g2_tiehi _5979__95 (.L_HI(net95));
 sg13g2_tiehi _5980__96 (.L_HI(net96));
 sg13g2_tiehi _5981__97 (.L_HI(net97));
 sg13g2_tiehi _5982__98 (.L_HI(net98));
 sg13g2_tiehi _5935__99 (.L_HI(net99));
 sg13g2_tiehi tt_um_iz_neuron_100 (.L_HI(net100));
 sg13g2_tiehi tt_um_iz_neuron_101 (.L_HI(net101));
 sg13g2_tiehi tt_um_iz_neuron_102 (.L_HI(net102));
 sg13g2_tiehi tt_um_iz_neuron_103 (.L_HI(net103));
 sg13g2_tiehi tt_um_iz_neuron_104 (.L_HI(net104));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_iz_neuron_14 (.L_LO(net14));
 sg13g2_tielo tt_um_iz_neuron_15 (.L_LO(net15));
 sg13g2_tielo tt_um_iz_neuron_16 (.L_LO(net16));
 sg13g2_tielo tt_um_iz_neuron_17 (.L_LO(net17));
 sg13g2_tielo tt_um_iz_neuron_18 (.L_LO(net18));
 sg13g2_tielo tt_um_iz_neuron_19 (.L_LO(net19));
 sg13g2_tielo tt_um_iz_neuron_20 (.L_LO(net20));
 sg13g2_tielo tt_um_iz_neuron_21 (.L_LO(net21));
 sg13g2_tiehi _5969__22 (.L_HI(net22));
 sg13g2_buf_1 _6078_ (.A(spike_out_internal),
    .X(uio_out[0]));
 sg13g2_buf_1 _6079_ (.A(params_ready_internal),
    .X(uio_out[1]));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(_0483_));
 sg13g2_buf_2 fanout670 (.A(_0483_),
    .X(net670));
 sg13g2_buf_4 fanout671 (.X(net671),
    .A(_1995_));
 sg13g2_buf_1 fanout672 (.A(_1995_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_1491_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_1445_),
    .X(net674));
 sg13g2_buf_1 fanout675 (.A(_1445_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_1449_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_1449_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_1448_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(_1447_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_1447_),
    .X(net680));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(_2886_));
 sg13g2_buf_2 fanout682 (.A(_1322_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(net684),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_1321_),
    .X(net684));
 sg13g2_buf_4 fanout685 (.X(net685),
    .A(_1099_));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_1098_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_0968_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(net691),
    .X(net689));
 sg13g2_buf_1 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_0967_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_0905_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_0908_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(_0908_),
    .X(net695));
 sg13g2_buf_4 fanout696 (.X(net696),
    .A(_0788_));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(_0787_));
 sg13g2_buf_2 fanout698 (.A(_0787_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_0720_),
    .X(net699));
 sg13g2_buf_1 fanout700 (.A(_0720_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_0722_),
    .X(net701));
 sg13g2_buf_1 fanout702 (.A(_0722_),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_0726_),
    .X(net703));
 sg13g2_buf_1 fanout704 (.A(_0726_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_0611_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(net708),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_2071_),
    .X(net708));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(_0489_));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(_0488_));
 sg13g2_buf_2 fanout711 (.A(net713),
    .X(net711));
 sg13g2_buf_1 fanout712 (.A(net713),
    .X(net712));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(_2051_));
 sg13g2_buf_2 fanout714 (.A(_2027_),
    .X(net714));
 sg13g2_buf_1 fanout715 (.A(_2027_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_1999_),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(net719),
    .X(net717));
 sg13g2_buf_1 fanout718 (.A(net719),
    .X(net718));
 sg13g2_buf_4 fanout719 (.X(net719),
    .A(_1956_));
 sg13g2_buf_2 fanout720 (.A(net722),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(net722),
    .X(net721));
 sg13g2_buf_4 fanout722 (.X(net722),
    .A(_1582_));
 sg13g2_buf_4 fanout723 (.X(net723),
    .A(_2299_));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(net725));
 sg13g2_buf_4 fanout725 (.X(net725),
    .A(_2079_));
 sg13g2_buf_2 fanout726 (.A(net727),
    .X(net726));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(_2070_));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(net731));
 sg13g2_buf_2 fanout729 (.A(net731),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(net731),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_1340_),
    .X(net731));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(_1329_));
 sg13g2_buf_2 fanout733 (.A(_1329_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(net737),
    .X(net734));
 sg13g2_buf_1 fanout735 (.A(net737),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(net737),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(net739),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(net739),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_1318_),
    .X(net739));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(net741));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(_1307_));
 sg13g2_buf_2 fanout742 (.A(\system_inst.neuron.u[13] ),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(net744),
    .X(net743));
 sg13g2_buf_4 fanout744 (.X(net744),
    .A(\system_inst.internal_param_b[7] ));
 sg13g2_buf_4 fanout745 (.X(net745),
    .A(net170));
 sg13g2_buf_2 fanout746 (.A(\system_inst.internal_param_b[6] ),
    .X(net746));
 sg13g2_buf_4 fanout747 (.X(net747),
    .A(\system_inst.internal_param_b[5] ));
 sg13g2_buf_2 fanout748 (.A(net173),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(net750),
    .X(net749));
 sg13g2_buf_4 fanout750 (.X(net750),
    .A(\system_inst.internal_param_b[4] ));
 sg13g2_buf_2 fanout751 (.A(net752),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(net753),
    .X(net752));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(net162));
 sg13g2_buf_2 fanout754 (.A(net755),
    .X(net754));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(net168));
 sg13g2_buf_2 fanout756 (.A(net757),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(net758),
    .X(net757));
 sg13g2_buf_4 fanout758 (.X(net758),
    .A(net153));
 sg13g2_buf_2 fanout759 (.A(net760),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(\system_inst.internal_param_b[0] ),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(net762),
    .X(net761));
 sg13g2_buf_1 fanout762 (.A(net763),
    .X(net762));
 sg13g2_buf_4 fanout763 (.X(net763),
    .A(net167));
 sg13g2_buf_2 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(net766),
    .X(net765));
 sg13g2_buf_4 fanout766 (.X(net766),
    .A(net169));
 sg13g2_buf_2 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_4 fanout768 (.X(net768),
    .A(\system_inst.internal_param_a[4] ));
 sg13g2_buf_2 fanout769 (.A(\system_inst.internal_param_a[4] ),
    .X(net769));
 sg13g2_buf_4 fanout770 (.X(net770),
    .A(net775));
 sg13g2_buf_1 fanout771 (.A(net775),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(net773),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(net775),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_4 fanout775 (.X(net775),
    .A(\system_inst.internal_param_a[3] ));
 sg13g2_buf_2 fanout776 (.A(net777),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(net780),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(net780),
    .X(net779));
 sg13g2_buf_1 fanout780 (.A(\system_inst.internal_param_a[2] ),
    .X(net780));
 sg13g2_buf_4 fanout781 (.X(net781),
    .A(\system_inst.internal_param_a[2] ));
 sg13g2_buf_1 fanout782 (.A(\system_inst.internal_param_a[2] ),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(net784),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(net785),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(net788),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(net788),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(\system_inst.internal_param_a[1] ),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(net790),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(net791),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(net797),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(net793),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(net797),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(net796),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(net796),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(net797),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(\system_inst.internal_param_a[0] ));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(net799));
 sg13g2_buf_4 fanout799 (.X(net799),
    .A(net801));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(\system_inst.neuron.v[13] ));
 sg13g2_buf_2 fanout801 (.A(\system_inst.neuron.v[13] ),
    .X(net801));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(net803));
 sg13g2_buf_4 fanout803 (.X(net803),
    .A(net174));
 sg13g2_buf_4 fanout804 (.X(net804),
    .A(\system_inst.neuron.v[12] ));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(net806));
 sg13g2_buf_4 fanout806 (.X(net806),
    .A(net808));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(\system_inst.neuron.v[11] ));
 sg13g2_buf_2 fanout808 (.A(\system_inst.neuron.v[11] ),
    .X(net808));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(net812));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(net811));
 sg13g2_buf_4 fanout811 (.X(net811),
    .A(net812));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(\system_inst.neuron.v[10] ));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(\system_inst.neuron.v[9] ));
 sg13g2_buf_4 fanout814 (.X(net814),
    .A(net816));
 sg13g2_buf_2 fanout815 (.A(net816),
    .X(net815));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(\system_inst.neuron.v[9] ));
 sg13g2_buf_2 fanout817 (.A(net821),
    .X(net817));
 sg13g2_buf_4 fanout818 (.X(net818),
    .A(net821));
 sg13g2_buf_2 fanout819 (.A(net821),
    .X(net819));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(net821));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(\system_inst.neuron.v[8] ));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(\system_inst.neuron.membrane_scaled[8] ));
 sg13g2_buf_2 fanout823 (.A(\system_inst.neuron.membrane_scaled[8] ),
    .X(net823));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(net826));
 sg13g2_buf_4 fanout825 (.X(net825),
    .A(net826));
 sg13g2_buf_2 fanout826 (.A(\system_inst.neuron.membrane_scaled[8] ),
    .X(net826));
 sg13g2_buf_4 fanout827 (.X(net827),
    .A(\system_inst.neuron.membrane_scaled[7] ));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(\system_inst.neuron.membrane_scaled[7] ));
 sg13g2_buf_4 fanout829 (.X(net829),
    .A(net832));
 sg13g2_buf_4 fanout830 (.X(net830),
    .A(net832));
 sg13g2_buf_2 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(\system_inst.neuron.membrane_scaled[7] ),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(net834),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(net835),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(net839),
    .X(net835));
 sg13g2_buf_4 fanout836 (.X(net836),
    .A(net839));
 sg13g2_buf_4 fanout837 (.X(net837),
    .A(net838));
 sg13g2_buf_2 fanout838 (.A(net839),
    .X(net838));
 sg13g2_buf_4 fanout839 (.X(net839),
    .A(\system_inst.neuron.membrane_scaled[6] ));
 sg13g2_buf_4 fanout840 (.X(net840),
    .A(net845));
 sg13g2_buf_4 fanout841 (.X(net841),
    .A(net845));
 sg13g2_buf_2 fanout842 (.A(net845),
    .X(net842));
 sg13g2_buf_4 fanout843 (.X(net843),
    .A(net844));
 sg13g2_buf_2 fanout844 (.A(net845),
    .X(net844));
 sg13g2_buf_4 fanout845 (.X(net845),
    .A(\system_inst.neuron.membrane_scaled[5] ));
 sg13g2_buf_2 fanout846 (.A(net847),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(net851),
    .X(net847));
 sg13g2_buf_4 fanout848 (.X(net848),
    .A(net851));
 sg13g2_buf_2 fanout849 (.A(net850),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net851),
    .X(net850));
 sg13g2_buf_4 fanout851 (.X(net851),
    .A(\system_inst.neuron.membrane_scaled[4] ));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net858),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(net855),
    .X(net854));
 sg13g2_buf_1 fanout855 (.A(net858),
    .X(net855));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(net858));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(net858));
 sg13g2_buf_4 fanout858 (.X(net858),
    .A(\system_inst.neuron.membrane_scaled[3] ));
 sg13g2_buf_2 fanout859 (.A(net860),
    .X(net859));
 sg13g2_buf_1 fanout860 (.A(net865),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(net862),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(net865),
    .X(net862));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(net865));
 sg13g2_buf_2 fanout864 (.A(net865),
    .X(net864));
 sg13g2_buf_4 fanout865 (.X(net865),
    .A(\system_inst.neuron.membrane_scaled[2] ));
 sg13g2_buf_2 fanout866 (.A(net868),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(net868),
    .X(net867));
 sg13g2_buf_4 fanout868 (.X(net868),
    .A(\system_inst.neuron.membrane_scaled[1] ));
 sg13g2_buf_2 fanout869 (.A(net870),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(\system_inst.neuron.membrane_scaled[1] ),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(net872),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(net873),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(net874),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(net875),
    .X(net874));
 sg13g2_buf_4 fanout875 (.X(net875),
    .A(_1516_));
 sg13g2_buf_2 fanout876 (.A(net877),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(net878),
    .X(net877));
 sg13g2_buf_4 fanout878 (.X(net878),
    .A(net884));
 sg13g2_buf_2 fanout879 (.A(net881),
    .X(net879));
 sg13g2_buf_1 fanout880 (.A(net881),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(net884),
    .X(net881));
 sg13g2_buf_4 fanout882 (.X(net882),
    .A(net883));
 sg13g2_buf_4 fanout883 (.X(net883),
    .A(net884));
 sg13g2_buf_2 fanout884 (.A(rst_n),
    .X(net884));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_4 input2 (.X(net2),
    .A(ui_in[0]));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[1]));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_4 input5 (.X(net5),
    .A(ui_in[3]));
 sg13g2_buf_2 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[2]),
    .X(net12));
 sg13g2_tielo tt_um_iz_neuron_13 (.L_LO(net13));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\system_inst.loader.bit_count[1] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold2 (.A(_2092_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0095_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold4 (.A(\system_inst.loader.state[5] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0005_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0018_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold7 (.A(\system_inst.loader.bit_count[0] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold8 (.A(\system_inst.internal_param_c[0] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold9 (.A(\system_inst.loader.bit_count[2] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0096_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold11 (.A(\system_inst.loader.state[3] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold12 (.A(_1914_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold13 (.A(\system_inst.internal_param_c[3] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0075_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold15 (.A(\system_inst.loader.shift_reg[5] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0093_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold17 (.A(\system_inst.loader.shift_reg[4] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold18 (.A(\system_inst.internal_param_d[4] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0083_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold20 (.A(\system_inst.internal_param_c[4] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0076_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold22 (.A(\system_inst.internal_param_c[6] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold23 (.A(\system_inst.loader.state[1] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold24 (.A(\system_inst.loader.shift_reg[0] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0088_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold26 (.A(\system_inst.internal_param_c[1] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold27 (.A(\system_inst.internal_param_c[2] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0074_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold29 (.A(\system_inst.loader.state[4] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold30 (.A(_1967_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold31 (.A(\system_inst.loader.state[2] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold32 (.A(\system_inst.internal_param_c[5] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold33 (.A(\system_inst.loader.shift_reg[2] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0090_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold35 (.A(\system_inst.loader.shift_reg[1] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold36 (.A(\system_inst.internal_param_d[7] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0086_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold38 (.A(\system_inst.loader.shift_reg[6] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0063_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold40 (.A(\system_inst.internal_param_d[6] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold41 (.A(\system_inst.internal_param_d[2] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold42 (.A(params_ready_internal),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0055_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold44 (.A(\system_inst.internal_param_d[3] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold45 (.A(\system_inst.loader.shift_reg[3] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0030_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold47 (.A(\system_inst.internal_param_d[0] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0079_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold49 (.A(\system_inst.internal_param_b[1] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0065_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold51 (.A(\system_inst.internal_param_d[1] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold52 (.A(\system_inst.neuron.u[0] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0007_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0105_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0016_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold56 (.A(\system_inst.internal_param_b[4] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold57 (.A(\system_inst.internal_param_d[5] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold58 (.A(\system_inst.internal_param_b[3] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold59 (.A(\system_inst.internal_param_b[0] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0064_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0028_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold62 (.A(\system_inst.loader.state[0] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold63 (.A(\system_inst.internal_param_a[6] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold64 (.A(\system_inst.internal_param_b[2] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold65 (.A(\system_inst.internal_param_a[5] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold66 (.A(\system_inst.internal_param_b[6] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0017_),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0535_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold69 (.A(\system_inst.internal_param_b[5] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold70 (.A(\system_inst.neuron.v[12] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold71 (.A(\system_inst.neuron.u[3] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0054_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0010_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0102_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold75 (.A(\system_inst.neuron.u[1] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold76 (.A(\system_inst.neuron.u[2] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold77 (.A(\system_inst.neuron.u[6] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0033_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold79 (.A(\system_inst.neuron.u[11] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0104_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold81 (.A(\system_inst.neuron.u[8] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold82 (.A(\system_inst.neuron.u[5] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0098_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold84 (.A(\system_inst.neuron.u[7] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold85 (.A(\system_inst.neuron.u[10] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold86 (.A(\system_inst.neuron.u[4] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold87 (.A(\system_inst.neuron.u[12] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold88 (.A(\system_inst.loader.shift_reg[0] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold89 (.A(_2028_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold90 (.A(_2030_),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0028_),
    .X(net195));
 sg13g2_antennanp ANTENNA_1 (.A(_0055_));
 sg13g2_antennanp ANTENNA_2 (.A(_0055_));
 sg13g2_antennanp ANTENNA_3 (.A(_0055_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_fill_2 FILLER_0_336 ();
 sg13g2_fill_1 FILLER_0_338 ();
 sg13g2_decap_4 FILLER_0_345 ();
 sg13g2_fill_2 FILLER_0_349 ();
 sg13g2_decap_4 FILLER_0_374 ();
 sg13g2_decap_4 FILLER_0_396 ();
 sg13g2_fill_2 FILLER_0_400 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_4 FILLER_1_322 ();
 sg13g2_fill_2 FILLER_1_326 ();
 sg13g2_decap_4 FILLER_1_333 ();
 sg13g2_fill_1 FILLER_1_358 ();
 sg13g2_fill_1 FILLER_1_366 ();
 sg13g2_fill_1 FILLER_1_379 ();
 sg13g2_fill_1 FILLER_1_388 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_fill_1 FILLER_2_322 ();
 sg13g2_fill_2 FILLER_2_333 ();
 sg13g2_fill_1 FILLER_2_335 ();
 sg13g2_decap_4 FILLER_2_346 ();
 sg13g2_fill_1 FILLER_2_350 ();
 sg13g2_decap_4 FILLER_2_359 ();
 sg13g2_fill_1 FILLER_2_363 ();
 sg13g2_fill_1 FILLER_2_386 ();
 sg13g2_fill_2 FILLER_2_395 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_4 FILLER_3_259 ();
 sg13g2_fill_1 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_269 ();
 sg13g2_decap_8 FILLER_3_276 ();
 sg13g2_decap_8 FILLER_3_283 ();
 sg13g2_decap_8 FILLER_3_290 ();
 sg13g2_decap_8 FILLER_3_297 ();
 sg13g2_decap_8 FILLER_3_304 ();
 sg13g2_decap_8 FILLER_3_311 ();
 sg13g2_decap_8 FILLER_3_318 ();
 sg13g2_decap_4 FILLER_3_325 ();
 sg13g2_fill_1 FILLER_3_334 ();
 sg13g2_fill_1 FILLER_3_349 ();
 sg13g2_fill_1 FILLER_3_363 ();
 sg13g2_fill_1 FILLER_3_384 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_4 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_286 ();
 sg13g2_decap_8 FILLER_4_293 ();
 sg13g2_decap_8 FILLER_4_300 ();
 sg13g2_decap_8 FILLER_4_307 ();
 sg13g2_decap_8 FILLER_4_314 ();
 sg13g2_fill_1 FILLER_4_321 ();
 sg13g2_fill_2 FILLER_4_358 ();
 sg13g2_fill_2 FILLER_4_372 ();
 sg13g2_fill_1 FILLER_4_374 ();
 sg13g2_fill_2 FILLER_4_385 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_fill_2 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_174 ();
 sg13g2_decap_8 FILLER_5_181 ();
 sg13g2_decap_8 FILLER_5_188 ();
 sg13g2_decap_8 FILLER_5_195 ();
 sg13g2_decap_8 FILLER_5_202 ();
 sg13g2_decap_8 FILLER_5_209 ();
 sg13g2_decap_8 FILLER_5_216 ();
 sg13g2_decap_8 FILLER_5_223 ();
 sg13g2_decap_4 FILLER_5_230 ();
 sg13g2_fill_2 FILLER_5_238 ();
 sg13g2_fill_1 FILLER_5_250 ();
 sg13g2_fill_2 FILLER_5_259 ();
 sg13g2_fill_1 FILLER_5_261 ();
 sg13g2_fill_1 FILLER_5_275 ();
 sg13g2_fill_1 FILLER_5_284 ();
 sg13g2_fill_1 FILLER_5_293 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_fill_1 FILLER_5_330 ();
 sg13g2_fill_2 FILLER_5_336 ();
 sg13g2_fill_2 FILLER_5_348 ();
 sg13g2_fill_1 FILLER_5_359 ();
 sg13g2_fill_2 FILLER_5_369 ();
 sg13g2_fill_1 FILLER_5_371 ();
 sg13g2_fill_1 FILLER_5_384 ();
 sg13g2_fill_2 FILLER_5_398 ();
 sg13g2_fill_1 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_4 FILLER_6_154 ();
 sg13g2_fill_1 FILLER_6_158 ();
 sg13g2_decap_8 FILLER_6_183 ();
 sg13g2_decap_8 FILLER_6_190 ();
 sg13g2_decap_8 FILLER_6_197 ();
 sg13g2_decap_8 FILLER_6_204 ();
 sg13g2_decap_8 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_218 ();
 sg13g2_fill_2 FILLER_6_225 ();
 sg13g2_fill_1 FILLER_6_227 ();
 sg13g2_fill_1 FILLER_6_259 ();
 sg13g2_fill_2 FILLER_6_268 ();
 sg13g2_fill_1 FILLER_6_270 ();
 sg13g2_fill_1 FILLER_6_283 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_fill_1 FILLER_6_315 ();
 sg13g2_decap_4 FILLER_6_334 ();
 sg13g2_fill_1 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_4 FILLER_7_140 ();
 sg13g2_decap_4 FILLER_7_147 ();
 sg13g2_fill_1 FILLER_7_179 ();
 sg13g2_decap_8 FILLER_7_192 ();
 sg13g2_decap_8 FILLER_7_199 ();
 sg13g2_decap_8 FILLER_7_206 ();
 sg13g2_decap_8 FILLER_7_213 ();
 sg13g2_decap_8 FILLER_7_220 ();
 sg13g2_decap_4 FILLER_7_227 ();
 sg13g2_fill_2 FILLER_7_231 ();
 sg13g2_decap_4 FILLER_7_238 ();
 sg13g2_fill_1 FILLER_7_242 ();
 sg13g2_fill_2 FILLER_7_267 ();
 sg13g2_fill_1 FILLER_7_269 ();
 sg13g2_fill_2 FILLER_7_293 ();
 sg13g2_fill_2 FILLER_7_302 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_fill_2 FILLER_7_315 ();
 sg13g2_fill_1 FILLER_7_317 ();
 sg13g2_fill_1 FILLER_7_323 ();
 sg13g2_decap_4 FILLER_7_328 ();
 sg13g2_fill_2 FILLER_7_339 ();
 sg13g2_fill_1 FILLER_7_341 ();
 sg13g2_fill_2 FILLER_7_354 ();
 sg13g2_fill_2 FILLER_7_379 ();
 sg13g2_fill_1 FILLER_7_381 ();
 sg13g2_fill_1 FILLER_7_401 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_fill_1 FILLER_8_133 ();
 sg13g2_decap_4 FILLER_8_164 ();
 sg13g2_decap_8 FILLER_8_204 ();
 sg13g2_decap_8 FILLER_8_211 ();
 sg13g2_decap_8 FILLER_8_218 ();
 sg13g2_decap_4 FILLER_8_225 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_fill_1 FILLER_8_249 ();
 sg13g2_fill_2 FILLER_8_263 ();
 sg13g2_fill_1 FILLER_8_321 ();
 sg13g2_fill_2 FILLER_8_338 ();
 sg13g2_fill_1 FILLER_8_356 ();
 sg13g2_fill_2 FILLER_8_388 ();
 sg13g2_fill_1 FILLER_8_390 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_fill_2 FILLER_9_158 ();
 sg13g2_fill_1 FILLER_9_160 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_191 ();
 sg13g2_decap_8 FILLER_9_198 ();
 sg13g2_decap_8 FILLER_9_205 ();
 sg13g2_decap_8 FILLER_9_212 ();
 sg13g2_decap_8 FILLER_9_219 ();
 sg13g2_fill_1 FILLER_9_226 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_fill_2 FILLER_9_245 ();
 sg13g2_decap_4 FILLER_9_289 ();
 sg13g2_decap_4 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_fill_2 FILLER_9_327 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_fill_2 FILLER_9_341 ();
 sg13g2_fill_1 FILLER_9_343 ();
 sg13g2_fill_1 FILLER_9_349 ();
 sg13g2_fill_2 FILLER_9_366 ();
 sg13g2_fill_1 FILLER_9_368 ();
 sg13g2_fill_2 FILLER_9_377 ();
 sg13g2_fill_1 FILLER_9_379 ();
 sg13g2_fill_2 FILLER_9_390 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_fill_2 FILLER_10_189 ();
 sg13g2_fill_1 FILLER_10_191 ();
 sg13g2_decap_4 FILLER_10_202 ();
 sg13g2_fill_2 FILLER_10_206 ();
 sg13g2_fill_2 FILLER_10_213 ();
 sg13g2_fill_1 FILLER_10_215 ();
 sg13g2_fill_1 FILLER_10_227 ();
 sg13g2_fill_2 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_fill_2 FILLER_10_263 ();
 sg13g2_decap_4 FILLER_10_274 ();
 sg13g2_fill_1 FILLER_10_278 ();
 sg13g2_decap_4 FILLER_10_309 ();
 sg13g2_fill_1 FILLER_10_313 ();
 sg13g2_fill_2 FILLER_10_328 ();
 sg13g2_fill_1 FILLER_10_353 ();
 sg13g2_fill_2 FILLER_10_359 ();
 sg13g2_fill_1 FILLER_10_380 ();
 sg13g2_fill_2 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_4 FILLER_11_150 ();
 sg13g2_fill_1 FILLER_11_154 ();
 sg13g2_fill_2 FILLER_11_165 ();
 sg13g2_fill_1 FILLER_11_167 ();
 sg13g2_decap_8 FILLER_11_183 ();
 sg13g2_fill_1 FILLER_11_190 ();
 sg13g2_fill_2 FILLER_11_206 ();
 sg13g2_fill_2 FILLER_11_212 ();
 sg13g2_fill_1 FILLER_11_214 ();
 sg13g2_fill_2 FILLER_11_224 ();
 sg13g2_fill_1 FILLER_11_230 ();
 sg13g2_fill_1 FILLER_11_261 ();
 sg13g2_fill_2 FILLER_11_270 ();
 sg13g2_fill_2 FILLER_11_286 ();
 sg13g2_fill_1 FILLER_11_321 ();
 sg13g2_fill_1 FILLER_11_337 ();
 sg13g2_fill_2 FILLER_11_398 ();
 sg13g2_fill_1 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_fill_2 FILLER_12_119 ();
 sg13g2_decap_4 FILLER_12_125 ();
 sg13g2_fill_1 FILLER_12_161 ();
 sg13g2_fill_2 FILLER_12_167 ();
 sg13g2_fill_1 FILLER_12_169 ();
 sg13g2_fill_2 FILLER_12_180 ();
 sg13g2_fill_1 FILLER_12_182 ();
 sg13g2_fill_1 FILLER_12_188 ();
 sg13g2_decap_4 FILLER_12_194 ();
 sg13g2_fill_1 FILLER_12_198 ();
 sg13g2_fill_2 FILLER_12_212 ();
 sg13g2_fill_1 FILLER_12_214 ();
 sg13g2_fill_1 FILLER_12_260 ();
 sg13g2_decap_4 FILLER_12_273 ();
 sg13g2_fill_2 FILLER_12_281 ();
 sg13g2_fill_1 FILLER_12_291 ();
 sg13g2_decap_4 FILLER_12_302 ();
 sg13g2_fill_2 FILLER_12_321 ();
 sg13g2_decap_4 FILLER_12_331 ();
 sg13g2_fill_1 FILLER_12_350 ();
 sg13g2_fill_2 FILLER_12_360 ();
 sg13g2_decap_4 FILLER_12_367 ();
 sg13g2_fill_1 FILLER_12_383 ();
 sg13g2_fill_1 FILLER_12_394 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_4 FILLER_13_112 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_decap_4 FILLER_13_147 ();
 sg13g2_fill_2 FILLER_13_186 ();
 sg13g2_decap_4 FILLER_13_201 ();
 sg13g2_fill_1 FILLER_13_205 ();
 sg13g2_fill_1 FILLER_13_220 ();
 sg13g2_fill_1 FILLER_13_226 ();
 sg13g2_fill_1 FILLER_13_251 ();
 sg13g2_fill_1 FILLER_13_264 ();
 sg13g2_fill_1 FILLER_13_323 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_377 ();
 sg13g2_fill_2 FILLER_13_383 ();
 sg13g2_fill_1 FILLER_13_385 ();
 sg13g2_fill_2 FILLER_13_392 ();
 sg13g2_fill_1 FILLER_13_394 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_4 FILLER_14_119 ();
 sg13g2_fill_1 FILLER_14_123 ();
 sg13g2_fill_2 FILLER_14_162 ();
 sg13g2_fill_1 FILLER_14_164 ();
 sg13g2_fill_2 FILLER_14_188 ();
 sg13g2_fill_1 FILLER_14_190 ();
 sg13g2_fill_2 FILLER_14_212 ();
 sg13g2_fill_2 FILLER_14_219 ();
 sg13g2_fill_1 FILLER_14_221 ();
 sg13g2_fill_2 FILLER_14_227 ();
 sg13g2_fill_1 FILLER_14_229 ();
 sg13g2_fill_1 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_300 ();
 sg13g2_fill_2 FILLER_14_307 ();
 sg13g2_fill_2 FILLER_14_319 ();
 sg13g2_fill_1 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_fill_1 FILLER_14_336 ();
 sg13g2_fill_1 FILLER_14_347 ();
 sg13g2_fill_1 FILLER_14_358 ();
 sg13g2_fill_2 FILLER_14_364 ();
 sg13g2_fill_1 FILLER_14_370 ();
 sg13g2_fill_1 FILLER_14_391 ();
 sg13g2_fill_2 FILLER_14_396 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_4 FILLER_15_117 ();
 sg13g2_fill_1 FILLER_15_129 ();
 sg13g2_decap_4 FILLER_15_145 ();
 sg13g2_fill_1 FILLER_15_169 ();
 sg13g2_fill_2 FILLER_15_177 ();
 sg13g2_fill_1 FILLER_15_199 ();
 sg13g2_fill_2 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_240 ();
 sg13g2_decap_4 FILLER_15_246 ();
 sg13g2_fill_1 FILLER_15_250 ();
 sg13g2_fill_1 FILLER_15_270 ();
 sg13g2_decap_4 FILLER_15_280 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_fill_1 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_4 FILLER_16_98 ();
 sg13g2_fill_2 FILLER_16_102 ();
 sg13g2_fill_2 FILLER_16_145 ();
 sg13g2_fill_1 FILLER_16_147 ();
 sg13g2_fill_2 FILLER_16_164 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_decap_8 FILLER_16_185 ();
 sg13g2_fill_1 FILLER_16_192 ();
 sg13g2_fill_2 FILLER_16_220 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_fill_2 FILLER_16_320 ();
 sg13g2_decap_4 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_332 ();
 sg13g2_decap_4 FILLER_16_350 ();
 sg13g2_fill_2 FILLER_16_368 ();
 sg13g2_fill_2 FILLER_16_393 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_4 FILLER_17_98 ();
 sg13g2_fill_1 FILLER_17_102 ();
 sg13g2_decap_8 FILLER_17_111 ();
 sg13g2_fill_2 FILLER_17_118 ();
 sg13g2_fill_1 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_136 ();
 sg13g2_fill_2 FILLER_17_143 ();
 sg13g2_fill_1 FILLER_17_173 ();
 sg13g2_fill_1 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_188 ();
 sg13g2_fill_2 FILLER_17_195 ();
 sg13g2_fill_2 FILLER_17_205 ();
 sg13g2_fill_1 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_229 ();
 sg13g2_decap_4 FILLER_17_244 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_fill_2 FILLER_17_258 ();
 sg13g2_fill_1 FILLER_17_260 ();
 sg13g2_fill_2 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_decap_8 FILLER_17_274 ();
 sg13g2_fill_1 FILLER_17_281 ();
 sg13g2_fill_2 FILLER_17_304 ();
 sg13g2_fill_2 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_373 ();
 sg13g2_fill_2 FILLER_17_390 ();
 sg13g2_fill_2 FILLER_17_397 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_4 FILLER_18_91 ();
 sg13g2_fill_2 FILLER_18_121 ();
 sg13g2_fill_2 FILLER_18_144 ();
 sg13g2_decap_4 FILLER_18_151 ();
 sg13g2_fill_1 FILLER_18_168 ();
 sg13g2_fill_2 FILLER_18_177 ();
 sg13g2_fill_2 FILLER_18_194 ();
 sg13g2_fill_2 FILLER_18_206 ();
 sg13g2_fill_1 FILLER_18_208 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_fill_1 FILLER_18_228 ();
 sg13g2_decap_4 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_253 ();
 sg13g2_fill_1 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_292 ();
 sg13g2_fill_2 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_381 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_4 FILLER_19_98 ();
 sg13g2_fill_2 FILLER_19_102 ();
 sg13g2_fill_2 FILLER_19_109 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_191 ();
 sg13g2_fill_1 FILLER_19_193 ();
 sg13g2_fill_1 FILLER_19_206 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_4 FILLER_19_297 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_308 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_fill_1 FILLER_19_342 ();
 sg13g2_fill_2 FILLER_19_366 ();
 sg13g2_fill_1 FILLER_19_368 ();
 sg13g2_decap_4 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_fill_2 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_107 ();
 sg13g2_fill_2 FILLER_20_113 ();
 sg13g2_fill_1 FILLER_20_115 ();
 sg13g2_fill_1 FILLER_20_126 ();
 sg13g2_fill_2 FILLER_20_135 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_149 ();
 sg13g2_fill_1 FILLER_20_156 ();
 sg13g2_decap_4 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_177 ();
 sg13g2_decap_4 FILLER_20_184 ();
 sg13g2_fill_2 FILLER_20_192 ();
 sg13g2_fill_2 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_224 ();
 sg13g2_fill_1 FILLER_20_239 ();
 sg13g2_fill_2 FILLER_20_253 ();
 sg13g2_fill_2 FILLER_20_267 ();
 sg13g2_fill_1 FILLER_20_281 ();
 sg13g2_decap_4 FILLER_20_292 ();
 sg13g2_fill_2 FILLER_20_334 ();
 sg13g2_fill_2 FILLER_20_382 ();
 sg13g2_fill_1 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_4 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_95 ();
 sg13g2_fill_2 FILLER_21_117 ();
 sg13g2_fill_2 FILLER_21_126 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_fill_2 FILLER_21_166 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_210 ();
 sg13g2_fill_2 FILLER_21_220 ();
 sg13g2_fill_2 FILLER_21_234 ();
 sg13g2_fill_1 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_245 ();
 sg13g2_decap_4 FILLER_21_328 ();
 sg13g2_fill_2 FILLER_21_340 ();
 sg13g2_decap_4 FILLER_21_360 ();
 sg13g2_fill_2 FILLER_21_373 ();
 sg13g2_fill_1 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_4 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_134 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_143 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_179 ();
 sg13g2_fill_2 FILLER_22_189 ();
 sg13g2_fill_1 FILLER_22_191 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_fill_2 FILLER_22_224 ();
 sg13g2_fill_1 FILLER_22_226 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_fill_2 FILLER_22_258 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_decap_4 FILLER_22_279 ();
 sg13g2_decap_4 FILLER_22_288 ();
 sg13g2_fill_1 FILLER_22_292 ();
 sg13g2_decap_4 FILLER_22_298 ();
 sg13g2_decap_4 FILLER_22_307 ();
 sg13g2_fill_1 FILLER_22_311 ();
 sg13g2_decap_4 FILLER_22_324 ();
 sg13g2_decap_4 FILLER_22_348 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_fill_2 FILLER_22_375 ();
 sg13g2_decap_4 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_4 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_95 ();
 sg13g2_fill_2 FILLER_23_144 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_225 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_decap_8 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_fill_1 FILLER_23_262 ();
 sg13g2_fill_1 FILLER_23_300 ();
 sg13g2_fill_2 FILLER_23_317 ();
 sg13g2_fill_2 FILLER_23_335 ();
 sg13g2_fill_1 FILLER_23_337 ();
 sg13g2_fill_2 FILLER_23_359 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_382 ();
 sg13g2_fill_1 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_109 ();
 sg13g2_fill_1 FILLER_24_111 ();
 sg13g2_fill_2 FILLER_24_117 ();
 sg13g2_fill_1 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_128 ();
 sg13g2_fill_1 FILLER_24_130 ();
 sg13g2_fill_2 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_fill_2 FILLER_24_144 ();
 sg13g2_fill_1 FILLER_24_146 ();
 sg13g2_fill_1 FILLER_24_167 ();
 sg13g2_decap_4 FILLER_24_176 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_decap_4 FILLER_24_186 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_2 FILLER_24_195 ();
 sg13g2_fill_1 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_236 ();
 sg13g2_fill_1 FILLER_24_245 ();
 sg13g2_fill_2 FILLER_24_263 ();
 sg13g2_decap_4 FILLER_24_274 ();
 sg13g2_fill_2 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_311 ();
 sg13g2_decap_4 FILLER_24_329 ();
 sg13g2_decap_4 FILLER_24_338 ();
 sg13g2_fill_2 FILLER_24_347 ();
 sg13g2_decap_4 FILLER_24_359 ();
 sg13g2_fill_1 FILLER_24_363 ();
 sg13g2_fill_1 FILLER_24_369 ();
 sg13g2_fill_1 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_4 FILLER_25_91 ();
 sg13g2_fill_2 FILLER_25_127 ();
 sg13g2_decap_4 FILLER_25_169 ();
 sg13g2_fill_1 FILLER_25_173 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_200 ();
 sg13g2_decap_8 FILLER_25_206 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_fill_2 FILLER_25_252 ();
 sg13g2_decap_4 FILLER_25_290 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_decap_4 FILLER_25_303 ();
 sg13g2_fill_2 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_fill_1 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_91 ();
 sg13g2_fill_2 FILLER_26_101 ();
 sg13g2_decap_8 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_118 ();
 sg13g2_fill_1 FILLER_26_125 ();
 sg13g2_decap_4 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_fill_1 FILLER_26_209 ();
 sg13g2_decap_4 FILLER_26_215 ();
 sg13g2_fill_2 FILLER_26_226 ();
 sg13g2_fill_2 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_272 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_fill_1 FILLER_26_294 ();
 sg13g2_fill_2 FILLER_26_307 ();
 sg13g2_fill_1 FILLER_26_309 ();
 sg13g2_decap_4 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_367 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_4 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_fill_1 FILLER_27_124 ();
 sg13g2_fill_2 FILLER_27_136 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_decap_4 FILLER_27_173 ();
 sg13g2_decap_4 FILLER_27_186 ();
 sg13g2_fill_2 FILLER_27_190 ();
 sg13g2_fill_1 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_fill_2 FILLER_27_282 ();
 sg13g2_fill_2 FILLER_27_292 ();
 sg13g2_fill_1 FILLER_27_298 ();
 sg13g2_decap_4 FILLER_27_307 ();
 sg13g2_fill_1 FILLER_27_316 ();
 sg13g2_fill_2 FILLER_27_361 ();
 sg13g2_fill_1 FILLER_27_368 ();
 sg13g2_decap_4 FILLER_27_382 ();
 sg13g2_fill_2 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_fill_2 FILLER_28_104 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_1 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_213 ();
 sg13g2_fill_2 FILLER_28_220 ();
 sg13g2_decap_8 FILLER_28_227 ();
 sg13g2_fill_2 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_fill_1 FILLER_28_242 ();
 sg13g2_fill_1 FILLER_28_273 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_fill_2 FILLER_28_287 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_fill_2 FILLER_28_342 ();
 sg13g2_fill_1 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_111 ();
 sg13g2_fill_1 FILLER_29_113 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_126 ();
 sg13g2_decap_4 FILLER_29_144 ();
 sg13g2_fill_2 FILLER_29_148 ();
 sg13g2_decap_8 FILLER_29_156 ();
 sg13g2_decap_4 FILLER_29_166 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_decap_4 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_223 ();
 sg13g2_decap_4 FILLER_29_228 ();
 sg13g2_fill_1 FILLER_29_281 ();
 sg13g2_decap_8 FILLER_29_298 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_313 ();
 sg13g2_fill_2 FILLER_29_334 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_fill_1 FILLER_29_367 ();
 sg13g2_fill_2 FILLER_29_373 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_125 ();
 sg13g2_fill_2 FILLER_30_148 ();
 sg13g2_fill_2 FILLER_30_172 ();
 sg13g2_fill_1 FILLER_30_174 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_4 FILLER_30_196 ();
 sg13g2_fill_1 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_234 ();
 sg13g2_decap_4 FILLER_30_248 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_267 ();
 sg13g2_fill_1 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_313 ();
 sg13g2_fill_2 FILLER_30_362 ();
 sg13g2_decap_4 FILLER_30_380 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_4 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_130 ();
 sg13g2_fill_1 FILLER_31_135 ();
 sg13g2_decap_4 FILLER_31_141 ();
 sg13g2_fill_2 FILLER_31_155 ();
 sg13g2_fill_2 FILLER_31_180 ();
 sg13g2_fill_1 FILLER_31_182 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_206 ();
 sg13g2_fill_1 FILLER_31_208 ();
 sg13g2_fill_2 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_decap_4 FILLER_31_240 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_fill_2 FILLER_31_273 ();
 sg13g2_decap_4 FILLER_31_315 ();
 sg13g2_fill_2 FILLER_31_327 ();
 sg13g2_fill_1 FILLER_31_329 ();
 sg13g2_decap_4 FILLER_31_338 ();
 sg13g2_fill_2 FILLER_31_353 ();
 sg13g2_fill_2 FILLER_31_368 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_4 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_88 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_fill_2 FILLER_32_161 ();
 sg13g2_fill_2 FILLER_32_171 ();
 sg13g2_decap_4 FILLER_32_178 ();
 sg13g2_fill_2 FILLER_32_182 ();
 sg13g2_fill_2 FILLER_32_216 ();
 sg13g2_fill_2 FILLER_32_248 ();
 sg13g2_decap_4 FILLER_32_255 ();
 sg13g2_fill_2 FILLER_32_259 ();
 sg13g2_fill_2 FILLER_32_293 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_fill_2 FILLER_32_318 ();
 sg13g2_fill_1 FILLER_32_320 ();
 sg13g2_decap_4 FILLER_32_328 ();
 sg13g2_fill_1 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_353 ();
 sg13g2_fill_1 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_88 ();
 sg13g2_decap_4 FILLER_33_102 ();
 sg13g2_decap_4 FILLER_33_113 ();
 sg13g2_fill_2 FILLER_33_117 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_208 ();
 sg13g2_fill_2 FILLER_33_220 ();
 sg13g2_fill_1 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_246 ();
 sg13g2_decap_4 FILLER_33_302 ();
 sg13g2_decap_4 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_decap_4 FILLER_33_360 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_4 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_88 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_118 ();
 sg13g2_fill_2 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_127 ();
 sg13g2_fill_2 FILLER_34_132 ();
 sg13g2_fill_2 FILLER_34_144 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_4 FILLER_34_182 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_fill_1 FILLER_34_234 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_273 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_fill_1 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_363 ();
 sg13g2_decap_4 FILLER_34_404 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_4 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_121 ();
 sg13g2_fill_1 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_137 ();
 sg13g2_fill_1 FILLER_35_139 ();
 sg13g2_fill_2 FILLER_35_172 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_fill_1 FILLER_35_206 ();
 sg13g2_fill_2 FILLER_35_211 ();
 sg13g2_fill_2 FILLER_35_222 ();
 sg13g2_fill_1 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_242 ();
 sg13g2_fill_2 FILLER_35_257 ();
 sg13g2_fill_1 FILLER_35_259 ();
 sg13g2_decap_4 FILLER_35_324 ();
 sg13g2_decap_4 FILLER_35_335 ();
 sg13g2_decap_4 FILLER_35_356 ();
 sg13g2_fill_2 FILLER_35_389 ();
 sg13g2_fill_1 FILLER_35_391 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_4 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_88 ();
 sg13g2_fill_2 FILLER_36_102 ();
 sg13g2_decap_4 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_fill_2 FILLER_36_128 ();
 sg13g2_fill_2 FILLER_36_136 ();
 sg13g2_fill_2 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_168 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_188 ();
 sg13g2_fill_1 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_229 ();
 sg13g2_fill_2 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_244 ();
 sg13g2_fill_2 FILLER_36_252 ();
 sg13g2_fill_2 FILLER_36_262 ();
 sg13g2_decap_4 FILLER_36_273 ();
 sg13g2_fill_1 FILLER_36_277 ();
 sg13g2_fill_2 FILLER_36_291 ();
 sg13g2_fill_1 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_decap_8 FILLER_36_328 ();
 sg13g2_fill_1 FILLER_36_361 ();
 sg13g2_fill_1 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_fill_1 FILLER_37_84 ();
 sg13g2_fill_2 FILLER_37_101 ();
 sg13g2_fill_1 FILLER_37_103 ();
 sg13g2_fill_2 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_138 ();
 sg13g2_decap_4 FILLER_37_154 ();
 sg13g2_fill_2 FILLER_37_158 ();
 sg13g2_fill_2 FILLER_37_165 ();
 sg13g2_fill_1 FILLER_37_167 ();
 sg13g2_decap_4 FILLER_37_185 ();
 sg13g2_fill_1 FILLER_37_189 ();
 sg13g2_fill_2 FILLER_37_203 ();
 sg13g2_fill_1 FILLER_37_205 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_fill_2 FILLER_37_245 ();
 sg13g2_fill_1 FILLER_37_247 ();
 sg13g2_fill_2 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_258 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_fill_2 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_304 ();
 sg13g2_fill_1 FILLER_37_310 ();
 sg13g2_fill_1 FILLER_37_323 ();
 sg13g2_decap_4 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_350 ();
 sg13g2_fill_1 FILLER_37_361 ();
 sg13g2_fill_2 FILLER_37_367 ();
 sg13g2_fill_1 FILLER_37_369 ();
 sg13g2_fill_2 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_88 ();
 sg13g2_decap_8 FILLER_38_94 ();
 sg13g2_decap_4 FILLER_38_113 ();
 sg13g2_fill_1 FILLER_38_117 ();
 sg13g2_fill_2 FILLER_38_128 ();
 sg13g2_fill_2 FILLER_38_147 ();
 sg13g2_fill_2 FILLER_38_185 ();
 sg13g2_fill_2 FILLER_38_207 ();
 sg13g2_decap_4 FILLER_38_217 ();
 sg13g2_decap_4 FILLER_38_225 ();
 sg13g2_fill_2 FILLER_38_303 ();
 sg13g2_decap_4 FILLER_38_356 ();
 sg13g2_fill_2 FILLER_38_378 ();
 sg13g2_fill_2 FILLER_38_396 ();
 sg13g2_fill_1 FILLER_38_398 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_4 FILLER_39_77 ();
 sg13g2_fill_1 FILLER_39_110 ();
 sg13g2_fill_2 FILLER_39_126 ();
 sg13g2_fill_1 FILLER_39_141 ();
 sg13g2_fill_1 FILLER_39_150 ();
 sg13g2_fill_2 FILLER_39_178 ();
 sg13g2_decap_4 FILLER_39_185 ();
 sg13g2_fill_1 FILLER_39_189 ();
 sg13g2_fill_1 FILLER_39_218 ();
 sg13g2_decap_8 FILLER_39_227 ();
 sg13g2_fill_2 FILLER_39_264 ();
 sg13g2_fill_2 FILLER_39_284 ();
 sg13g2_fill_1 FILLER_39_286 ();
 sg13g2_fill_2 FILLER_39_369 ();
 sg13g2_fill_2 FILLER_39_391 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_4 FILLER_40_117 ();
 sg13g2_decap_4 FILLER_40_147 ();
 sg13g2_fill_2 FILLER_40_184 ();
 sg13g2_fill_1 FILLER_40_186 ();
 sg13g2_fill_2 FILLER_40_197 ();
 sg13g2_fill_1 FILLER_40_199 ();
 sg13g2_fill_1 FILLER_40_209 ();
 sg13g2_fill_2 FILLER_40_230 ();
 sg13g2_fill_2 FILLER_40_244 ();
 sg13g2_fill_2 FILLER_40_275 ();
 sg13g2_fill_1 FILLER_40_346 ();
 sg13g2_decap_4 FILLER_40_366 ();
 sg13g2_decap_4 FILLER_40_380 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_fill_2 FILLER_41_104 ();
 sg13g2_fill_1 FILLER_41_106 ();
 sg13g2_fill_1 FILLER_41_111 ();
 sg13g2_fill_2 FILLER_41_117 ();
 sg13g2_fill_1 FILLER_41_124 ();
 sg13g2_fill_2 FILLER_41_129 ();
 sg13g2_fill_2 FILLER_41_137 ();
 sg13g2_fill_2 FILLER_41_174 ();
 sg13g2_fill_1 FILLER_41_176 ();
 sg13g2_fill_2 FILLER_41_181 ();
 sg13g2_fill_1 FILLER_41_183 ();
 sg13g2_fill_1 FILLER_41_227 ();
 sg13g2_decap_8 FILLER_41_257 ();
 sg13g2_fill_2 FILLER_41_264 ();
 sg13g2_fill_1 FILLER_41_266 ();
 sg13g2_fill_1 FILLER_41_280 ();
 sg13g2_decap_4 FILLER_41_286 ();
 sg13g2_fill_1 FILLER_41_290 ();
 sg13g2_fill_2 FILLER_41_299 ();
 sg13g2_decap_8 FILLER_41_306 ();
 sg13g2_decap_4 FILLER_41_313 ();
 sg13g2_decap_8 FILLER_41_341 ();
 sg13g2_decap_4 FILLER_41_354 ();
 sg13g2_fill_1 FILLER_41_369 ();
 sg13g2_decap_4 FILLER_41_379 ();
 sg13g2_fill_1 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_fill_2 FILLER_42_77 ();
 sg13g2_fill_1 FILLER_42_86 ();
 sg13g2_fill_2 FILLER_42_134 ();
 sg13g2_fill_1 FILLER_42_148 ();
 sg13g2_fill_1 FILLER_42_157 ();
 sg13g2_fill_2 FILLER_42_178 ();
 sg13g2_fill_2 FILLER_42_185 ();
 sg13g2_decap_4 FILLER_42_196 ();
 sg13g2_fill_1 FILLER_42_217 ();
 sg13g2_fill_2 FILLER_42_234 ();
 sg13g2_fill_1 FILLER_42_241 ();
 sg13g2_fill_1 FILLER_42_247 ();
 sg13g2_fill_2 FILLER_42_258 ();
 sg13g2_fill_1 FILLER_42_260 ();
 sg13g2_fill_2 FILLER_42_265 ();
 sg13g2_fill_1 FILLER_42_280 ();
 sg13g2_decap_8 FILLER_42_321 ();
 sg13g2_decap_4 FILLER_42_342 ();
 sg13g2_fill_2 FILLER_42_398 ();
 sg13g2_fill_1 FILLER_42_400 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_4 FILLER_43_70 ();
 sg13g2_fill_1 FILLER_43_74 ();
 sg13g2_decap_8 FILLER_43_104 ();
 sg13g2_decap_8 FILLER_43_111 ();
 sg13g2_fill_2 FILLER_43_118 ();
 sg13g2_fill_2 FILLER_43_137 ();
 sg13g2_fill_2 FILLER_43_147 ();
 sg13g2_fill_1 FILLER_43_149 ();
 sg13g2_fill_2 FILLER_43_158 ();
 sg13g2_fill_1 FILLER_43_178 ();
 sg13g2_fill_2 FILLER_43_187 ();
 sg13g2_fill_1 FILLER_43_189 ();
 sg13g2_decap_4 FILLER_43_203 ();
 sg13g2_fill_1 FILLER_43_207 ();
 sg13g2_fill_2 FILLER_43_216 ();
 sg13g2_fill_2 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_288 ();
 sg13g2_decap_8 FILLER_43_295 ();
 sg13g2_decap_4 FILLER_43_302 ();
 sg13g2_fill_2 FILLER_43_306 ();
 sg13g2_fill_1 FILLER_43_326 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_fill_2 FILLER_43_365 ();
 sg13g2_fill_1 FILLER_43_377 ();
 sg13g2_fill_2 FILLER_43_392 ();
 sg13g2_fill_1 FILLER_43_394 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_fill_2 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_88 ();
 sg13g2_fill_1 FILLER_44_95 ();
 sg13g2_fill_1 FILLER_44_112 ();
 sg13g2_fill_1 FILLER_44_121 ();
 sg13g2_decap_4 FILLER_44_136 ();
 sg13g2_fill_1 FILLER_44_140 ();
 sg13g2_decap_4 FILLER_44_146 ();
 sg13g2_fill_2 FILLER_44_150 ();
 sg13g2_decap_4 FILLER_44_191 ();
 sg13g2_fill_2 FILLER_44_216 ();
 sg13g2_fill_1 FILLER_44_218 ();
 sg13g2_fill_2 FILLER_44_225 ();
 sg13g2_fill_1 FILLER_44_227 ();
 sg13g2_fill_2 FILLER_44_237 ();
 sg13g2_decap_8 FILLER_44_244 ();
 sg13g2_fill_2 FILLER_44_251 ();
 sg13g2_fill_1 FILLER_44_264 ();
 sg13g2_decap_4 FILLER_44_304 ();
 sg13g2_fill_1 FILLER_44_308 ();
 sg13g2_fill_1 FILLER_44_345 ();
 sg13g2_fill_2 FILLER_44_355 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_fill_1 FILLER_45_77 ();
 sg13g2_decap_4 FILLER_45_86 ();
 sg13g2_fill_2 FILLER_45_98 ();
 sg13g2_decap_4 FILLER_45_105 ();
 sg13g2_fill_1 FILLER_45_114 ();
 sg13g2_decap_4 FILLER_45_120 ();
 sg13g2_fill_1 FILLER_45_124 ();
 sg13g2_fill_2 FILLER_45_143 ();
 sg13g2_decap_8 FILLER_45_153 ();
 sg13g2_fill_2 FILLER_45_160 ();
 sg13g2_fill_2 FILLER_45_166 ();
 sg13g2_fill_2 FILLER_45_173 ();
 sg13g2_fill_2 FILLER_45_199 ();
 sg13g2_fill_2 FILLER_45_214 ();
 sg13g2_fill_2 FILLER_45_224 ();
 sg13g2_fill_2 FILLER_45_244 ();
 sg13g2_fill_2 FILLER_45_254 ();
 sg13g2_fill_1 FILLER_45_256 ();
 sg13g2_decap_8 FILLER_45_277 ();
 sg13g2_fill_1 FILLER_45_338 ();
 sg13g2_fill_2 FILLER_45_347 ();
 sg13g2_fill_2 FILLER_45_376 ();
 sg13g2_fill_1 FILLER_45_378 ();
 sg13g2_fill_1 FILLER_45_389 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_fill_2 FILLER_46_82 ();
 sg13g2_fill_1 FILLER_46_84 ();
 sg13g2_fill_2 FILLER_46_113 ();
 sg13g2_fill_1 FILLER_46_115 ();
 sg13g2_decap_8 FILLER_46_134 ();
 sg13g2_decap_4 FILLER_46_141 ();
 sg13g2_fill_1 FILLER_46_145 ();
 sg13g2_fill_1 FILLER_46_152 ();
 sg13g2_decap_4 FILLER_46_161 ();
 sg13g2_fill_1 FILLER_46_177 ();
 sg13g2_fill_2 FILLER_46_190 ();
 sg13g2_fill_1 FILLER_46_192 ();
 sg13g2_decap_4 FILLER_46_200 ();
 sg13g2_decap_4 FILLER_46_214 ();
 sg13g2_fill_2 FILLER_46_231 ();
 sg13g2_fill_1 FILLER_46_233 ();
 sg13g2_fill_1 FILLER_46_260 ();
 sg13g2_fill_1 FILLER_46_311 ();
 sg13g2_fill_1 FILLER_46_359 ();
 sg13g2_fill_1 FILLER_46_369 ();
 sg13g2_fill_1 FILLER_46_393 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_fill_2 FILLER_47_83 ();
 sg13g2_fill_2 FILLER_47_95 ();
 sg13g2_fill_1 FILLER_47_97 ();
 sg13g2_decap_8 FILLER_47_104 ();
 sg13g2_fill_1 FILLER_47_116 ();
 sg13g2_fill_2 FILLER_47_165 ();
 sg13g2_fill_1 FILLER_47_167 ();
 sg13g2_decap_4 FILLER_47_178 ();
 sg13g2_fill_1 FILLER_47_182 ();
 sg13g2_fill_2 FILLER_47_200 ();
 sg13g2_fill_1 FILLER_47_202 ();
 sg13g2_fill_2 FILLER_47_220 ();
 sg13g2_fill_1 FILLER_47_222 ();
 sg13g2_fill_1 FILLER_47_255 ();
 sg13g2_decap_4 FILLER_47_266 ();
 sg13g2_fill_1 FILLER_47_270 ();
 sg13g2_fill_2 FILLER_47_323 ();
 sg13g2_fill_2 FILLER_47_367 ();
 sg13g2_fill_1 FILLER_47_385 ();
 sg13g2_fill_2 FILLER_47_406 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_fill_2 FILLER_48_63 ();
 sg13g2_decap_4 FILLER_48_98 ();
 sg13g2_fill_2 FILLER_48_115 ();
 sg13g2_fill_1 FILLER_48_117 ();
 sg13g2_fill_2 FILLER_48_123 ();
 sg13g2_fill_1 FILLER_48_125 ();
 sg13g2_fill_2 FILLER_48_149 ();
 sg13g2_fill_1 FILLER_48_151 ();
 sg13g2_fill_2 FILLER_48_189 ();
 sg13g2_fill_2 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_206 ();
 sg13g2_fill_2 FILLER_48_213 ();
 sg13g2_fill_1 FILLER_48_215 ();
 sg13g2_decap_4 FILLER_48_228 ();
 sg13g2_fill_1 FILLER_48_232 ();
 sg13g2_fill_2 FILLER_48_281 ();
 sg13g2_fill_1 FILLER_48_308 ();
 sg13g2_fill_2 FILLER_48_359 ();
 sg13g2_fill_1 FILLER_48_361 ();
 sg13g2_fill_2 FILLER_48_379 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_fill_2 FILLER_49_70 ();
 sg13g2_fill_2 FILLER_49_81 ();
 sg13g2_fill_2 FILLER_49_132 ();
 sg13g2_fill_1 FILLER_49_139 ();
 sg13g2_fill_2 FILLER_49_156 ();
 sg13g2_decap_4 FILLER_49_176 ();
 sg13g2_fill_1 FILLER_49_188 ();
 sg13g2_fill_1 FILLER_49_200 ();
 sg13g2_fill_2 FILLER_49_212 ();
 sg13g2_fill_2 FILLER_49_227 ();
 sg13g2_fill_2 FILLER_49_241 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_4 FILLER_49_262 ();
 sg13g2_fill_2 FILLER_49_266 ();
 sg13g2_fill_1 FILLER_49_272 ();
 sg13g2_fill_2 FILLER_49_283 ();
 sg13g2_fill_2 FILLER_49_331 ();
 sg13g2_fill_2 FILLER_49_357 ();
 sg13g2_fill_2 FILLER_49_369 ();
 sg13g2_fill_1 FILLER_49_371 ();
 sg13g2_fill_1 FILLER_49_399 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_fill_1 FILLER_50_70 ();
 sg13g2_fill_2 FILLER_50_79 ();
 sg13g2_decap_8 FILLER_50_89 ();
 sg13g2_fill_2 FILLER_50_99 ();
 sg13g2_fill_1 FILLER_50_101 ();
 sg13g2_fill_2 FILLER_50_120 ();
 sg13g2_fill_1 FILLER_50_122 ();
 sg13g2_fill_1 FILLER_50_130 ();
 sg13g2_fill_2 FILLER_50_136 ();
 sg13g2_fill_1 FILLER_50_138 ();
 sg13g2_fill_2 FILLER_50_144 ();
 sg13g2_fill_1 FILLER_50_155 ();
 sg13g2_fill_2 FILLER_50_166 ();
 sg13g2_fill_2 FILLER_50_184 ();
 sg13g2_fill_1 FILLER_50_212 ();
 sg13g2_fill_2 FILLER_50_217 ();
 sg13g2_fill_1 FILLER_50_236 ();
 sg13g2_fill_1 FILLER_50_360 ();
 sg13g2_fill_2 FILLER_50_386 ();
 sg13g2_fill_1 FILLER_50_396 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_4 FILLER_51_63 ();
 sg13g2_fill_2 FILLER_51_67 ();
 sg13g2_fill_1 FILLER_51_107 ();
 sg13g2_fill_2 FILLER_51_119 ();
 sg13g2_fill_1 FILLER_51_121 ();
 sg13g2_fill_2 FILLER_51_130 ();
 sg13g2_fill_1 FILLER_51_137 ();
 sg13g2_fill_2 FILLER_51_154 ();
 sg13g2_fill_1 FILLER_51_176 ();
 sg13g2_fill_1 FILLER_51_181 ();
 sg13g2_fill_2 FILLER_51_201 ();
 sg13g2_decap_8 FILLER_51_215 ();
 sg13g2_fill_2 FILLER_51_222 ();
 sg13g2_fill_2 FILLER_51_265 ();
 sg13g2_fill_1 FILLER_51_267 ();
 sg13g2_fill_1 FILLER_51_286 ();
 sg13g2_fill_2 FILLER_51_304 ();
 sg13g2_fill_2 FILLER_51_348 ();
 sg13g2_fill_1 FILLER_51_350 ();
 sg13g2_fill_2 FILLER_51_358 ();
 sg13g2_fill_2 FILLER_51_372 ();
 sg13g2_fill_1 FILLER_51_374 ();
 sg13g2_fill_2 FILLER_51_384 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_fill_2 FILLER_52_63 ();
 sg13g2_fill_1 FILLER_52_65 ();
 sg13g2_decap_4 FILLER_52_79 ();
 sg13g2_fill_2 FILLER_52_106 ();
 sg13g2_fill_1 FILLER_52_108 ();
 sg13g2_fill_2 FILLER_52_130 ();
 sg13g2_fill_1 FILLER_52_132 ();
 sg13g2_decap_4 FILLER_52_152 ();
 sg13g2_fill_1 FILLER_52_156 ();
 sg13g2_fill_1 FILLER_52_162 ();
 sg13g2_fill_2 FILLER_52_176 ();
 sg13g2_fill_2 FILLER_52_191 ();
 sg13g2_fill_1 FILLER_52_246 ();
 sg13g2_fill_2 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_394 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_fill_2 FILLER_53_63 ();
 sg13g2_fill_1 FILLER_53_65 ();
 sg13g2_fill_2 FILLER_53_87 ();
 sg13g2_decap_4 FILLER_53_94 ();
 sg13g2_decap_4 FILLER_53_103 ();
 sg13g2_fill_1 FILLER_53_107 ();
 sg13g2_fill_2 FILLER_53_121 ();
 sg13g2_fill_1 FILLER_53_123 ();
 sg13g2_decap_4 FILLER_53_129 ();
 sg13g2_fill_1 FILLER_53_133 ();
 sg13g2_fill_2 FILLER_53_147 ();
 sg13g2_fill_2 FILLER_53_181 ();
 sg13g2_fill_1 FILLER_53_204 ();
 sg13g2_fill_2 FILLER_53_214 ();
 sg13g2_decap_8 FILLER_53_220 ();
 sg13g2_fill_1 FILLER_53_227 ();
 sg13g2_fill_1 FILLER_53_232 ();
 sg13g2_fill_1 FILLER_53_242 ();
 sg13g2_fill_2 FILLER_53_248 ();
 sg13g2_fill_2 FILLER_53_272 ();
 sg13g2_fill_2 FILLER_53_344 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_4 FILLER_54_63 ();
 sg13g2_fill_2 FILLER_54_67 ();
 sg13g2_fill_1 FILLER_54_77 ();
 sg13g2_fill_2 FILLER_54_87 ();
 sg13g2_fill_1 FILLER_54_89 ();
 sg13g2_fill_2 FILLER_54_263 ();
 sg13g2_fill_1 FILLER_54_278 ();
 sg13g2_fill_2 FILLER_54_289 ();
 sg13g2_fill_2 FILLER_54_295 ();
 sg13g2_fill_2 FILLER_54_304 ();
 sg13g2_fill_1 FILLER_54_311 ();
 sg13g2_fill_2 FILLER_54_321 ();
 sg13g2_fill_2 FILLER_54_393 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_fill_1 FILLER_55_104 ();
 sg13g2_fill_2 FILLER_55_110 ();
 sg13g2_fill_1 FILLER_55_151 ();
 sg13g2_fill_1 FILLER_55_165 ();
 sg13g2_fill_1 FILLER_55_171 ();
 sg13g2_fill_2 FILLER_55_177 ();
 sg13g2_fill_2 FILLER_55_208 ();
 sg13g2_fill_1 FILLER_55_210 ();
 sg13g2_fill_2 FILLER_55_224 ();
 sg13g2_fill_2 FILLER_55_234 ();
 sg13g2_fill_1 FILLER_55_236 ();
 sg13g2_fill_2 FILLER_55_245 ();
 sg13g2_fill_1 FILLER_55_269 ();
 sg13g2_fill_2 FILLER_55_278 ();
 sg13g2_fill_1 FILLER_55_280 ();
 sg13g2_fill_1 FILLER_55_320 ();
 sg13g2_fill_1 FILLER_55_338 ();
 sg13g2_fill_2 FILLER_55_364 ();
 sg13g2_fill_1 FILLER_55_376 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_4 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_79 ();
 sg13g2_fill_1 FILLER_56_110 ();
 sg13g2_fill_1 FILLER_56_124 ();
 sg13g2_fill_2 FILLER_56_130 ();
 sg13g2_decap_4 FILLER_56_152 ();
 sg13g2_fill_1 FILLER_56_183 ();
 sg13g2_fill_2 FILLER_56_194 ();
 sg13g2_fill_2 FILLER_56_203 ();
 sg13g2_fill_2 FILLER_56_218 ();
 sg13g2_fill_1 FILLER_56_285 ();
 sg13g2_fill_2 FILLER_56_291 ();
 sg13g2_fill_2 FILLER_56_302 ();
 sg13g2_fill_1 FILLER_56_340 ();
 sg13g2_fill_1 FILLER_56_346 ();
 sg13g2_fill_2 FILLER_56_389 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_4 FILLER_57_70 ();
 sg13g2_fill_2 FILLER_57_74 ();
 sg13g2_fill_2 FILLER_57_80 ();
 sg13g2_fill_1 FILLER_57_82 ();
 sg13g2_fill_2 FILLER_57_98 ();
 sg13g2_fill_1 FILLER_57_100 ();
 sg13g2_fill_1 FILLER_57_121 ();
 sg13g2_fill_1 FILLER_57_145 ();
 sg13g2_decap_8 FILLER_57_158 ();
 sg13g2_decap_4 FILLER_57_165 ();
 sg13g2_fill_1 FILLER_57_169 ();
 sg13g2_fill_2 FILLER_57_177 ();
 sg13g2_fill_1 FILLER_57_179 ();
 sg13g2_fill_1 FILLER_57_209 ();
 sg13g2_fill_2 FILLER_57_252 ();
 sg13g2_fill_1 FILLER_57_341 ();
 sg13g2_fill_2 FILLER_57_350 ();
 sg13g2_fill_1 FILLER_57_369 ();
 sg13g2_fill_1 FILLER_57_381 ();
 sg13g2_fill_1 FILLER_57_387 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_fill_2 FILLER_58_134 ();
 sg13g2_fill_2 FILLER_58_143 ();
 sg13g2_decap_8 FILLER_58_153 ();
 sg13g2_fill_2 FILLER_58_197 ();
 sg13g2_fill_1 FILLER_58_204 ();
 sg13g2_fill_2 FILLER_58_215 ();
 sg13g2_fill_1 FILLER_58_230 ();
 sg13g2_fill_1 FILLER_58_248 ();
 sg13g2_fill_1 FILLER_58_273 ();
 sg13g2_fill_2 FILLER_58_300 ();
 sg13g2_fill_2 FILLER_58_310 ();
 sg13g2_fill_2 FILLER_58_336 ();
 sg13g2_fill_1 FILLER_58_343 ();
 sg13g2_fill_2 FILLER_58_361 ();
 sg13g2_fill_1 FILLER_58_363 ();
 sg13g2_fill_1 FILLER_58_372 ();
 sg13g2_fill_2 FILLER_58_390 ();
 sg13g2_fill_1 FILLER_58_400 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_4 FILLER_59_70 ();
 sg13g2_fill_2 FILLER_59_74 ();
 sg13g2_fill_2 FILLER_59_98 ();
 sg13g2_fill_1 FILLER_59_100 ();
 sg13g2_fill_2 FILLER_59_109 ();
 sg13g2_fill_1 FILLER_59_111 ();
 sg13g2_fill_1 FILLER_59_136 ();
 sg13g2_decap_8 FILLER_59_142 ();
 sg13g2_fill_1 FILLER_59_149 ();
 sg13g2_decap_8 FILLER_59_176 ();
 sg13g2_decap_4 FILLER_59_183 ();
 sg13g2_fill_1 FILLER_59_187 ();
 sg13g2_fill_2 FILLER_59_203 ();
 sg13g2_fill_1 FILLER_59_205 ();
 sg13g2_fill_1 FILLER_59_221 ();
 sg13g2_fill_1 FILLER_59_291 ();
 sg13g2_fill_2 FILLER_59_372 ();
 sg13g2_fill_1 FILLER_59_374 ();
 sg13g2_fill_1 FILLER_59_381 ();
 sg13g2_fill_2 FILLER_59_400 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_4 FILLER_60_70 ();
 sg13g2_fill_1 FILLER_60_74 ();
 sg13g2_fill_2 FILLER_60_88 ();
 sg13g2_fill_1 FILLER_60_90 ();
 sg13g2_fill_1 FILLER_60_102 ();
 sg13g2_fill_2 FILLER_60_108 ();
 sg13g2_fill_2 FILLER_60_130 ();
 sg13g2_decap_4 FILLER_60_145 ();
 sg13g2_fill_2 FILLER_60_159 ();
 sg13g2_fill_1 FILLER_60_181 ();
 sg13g2_fill_2 FILLER_60_209 ();
 sg13g2_fill_2 FILLER_60_224 ();
 sg13g2_fill_1 FILLER_60_226 ();
 sg13g2_fill_1 FILLER_60_273 ();
 sg13g2_fill_1 FILLER_60_288 ();
 sg13g2_fill_1 FILLER_60_367 ();
 sg13g2_fill_1 FILLER_60_376 ();
 sg13g2_fill_1 FILLER_60_392 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_fill_2 FILLER_61_77 ();
 sg13g2_fill_1 FILLER_61_79 ();
 sg13g2_decap_4 FILLER_61_85 ();
 sg13g2_fill_1 FILLER_61_89 ();
 sg13g2_fill_2 FILLER_61_98 ();
 sg13g2_fill_1 FILLER_61_100 ();
 sg13g2_fill_2 FILLER_61_124 ();
 sg13g2_fill_1 FILLER_61_141 ();
 sg13g2_fill_2 FILLER_61_170 ();
 sg13g2_fill_2 FILLER_61_177 ();
 sg13g2_fill_1 FILLER_61_179 ();
 sg13g2_fill_1 FILLER_61_217 ();
 sg13g2_fill_2 FILLER_61_239 ();
 sg13g2_fill_1 FILLER_61_241 ();
 sg13g2_fill_2 FILLER_61_276 ();
 sg13g2_fill_2 FILLER_61_309 ();
 sg13g2_fill_1 FILLER_61_340 ();
 sg13g2_fill_1 FILLER_61_356 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_fill_1 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_97 ();
 sg13g2_fill_1 FILLER_62_104 ();
 sg13g2_fill_2 FILLER_62_133 ();
 sg13g2_fill_1 FILLER_62_143 ();
 sg13g2_fill_2 FILLER_62_160 ();
 sg13g2_fill_1 FILLER_62_162 ();
 sg13g2_fill_2 FILLER_62_173 ();
 sg13g2_fill_1 FILLER_62_183 ();
 sg13g2_fill_1 FILLER_62_208 ();
 sg13g2_fill_1 FILLER_62_226 ();
 sg13g2_fill_2 FILLER_62_257 ();
 sg13g2_fill_1 FILLER_62_259 ();
 sg13g2_fill_2 FILLER_62_265 ();
 sg13g2_fill_1 FILLER_62_267 ();
 sg13g2_fill_1 FILLER_62_282 ();
 sg13g2_fill_2 FILLER_62_302 ();
 sg13g2_fill_2 FILLER_62_309 ();
 sg13g2_fill_1 FILLER_62_319 ();
 sg13g2_fill_2 FILLER_62_368 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_fill_2 FILLER_63_70 ();
 sg13g2_fill_1 FILLER_63_72 ();
 sg13g2_decap_4 FILLER_63_110 ();
 sg13g2_fill_2 FILLER_63_145 ();
 sg13g2_fill_1 FILLER_63_147 ();
 sg13g2_fill_2 FILLER_63_200 ();
 sg13g2_fill_1 FILLER_63_202 ();
 sg13g2_fill_2 FILLER_63_208 ();
 sg13g2_fill_1 FILLER_63_210 ();
 sg13g2_fill_1 FILLER_63_221 ();
 sg13g2_fill_2 FILLER_63_235 ();
 sg13g2_fill_2 FILLER_63_244 ();
 sg13g2_fill_2 FILLER_63_294 ();
 sg13g2_fill_1 FILLER_63_296 ();
 sg13g2_fill_2 FILLER_63_317 ();
 sg13g2_fill_1 FILLER_63_319 ();
 sg13g2_fill_1 FILLER_63_338 ();
 sg13g2_fill_2 FILLER_63_354 ();
 sg13g2_fill_1 FILLER_63_373 ();
 sg13g2_fill_2 FILLER_63_379 ();
 sg13g2_fill_2 FILLER_63_389 ();
 sg13g2_fill_1 FILLER_63_391 ();
 sg13g2_fill_1 FILLER_63_400 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_fill_2 FILLER_64_77 ();
 sg13g2_fill_1 FILLER_64_79 ();
 sg13g2_decap_4 FILLER_64_88 ();
 sg13g2_fill_1 FILLER_64_92 ();
 sg13g2_fill_2 FILLER_64_101 ();
 sg13g2_fill_1 FILLER_64_103 ();
 sg13g2_fill_1 FILLER_64_122 ();
 sg13g2_fill_1 FILLER_64_138 ();
 sg13g2_fill_2 FILLER_64_182 ();
 sg13g2_fill_1 FILLER_64_184 ();
 sg13g2_fill_2 FILLER_64_218 ();
 sg13g2_fill_1 FILLER_64_240 ();
 sg13g2_fill_2 FILLER_64_246 ();
 sg13g2_fill_2 FILLER_64_262 ();
 sg13g2_fill_1 FILLER_64_264 ();
 sg13g2_fill_2 FILLER_64_274 ();
 sg13g2_fill_1 FILLER_64_296 ();
 sg13g2_fill_2 FILLER_64_307 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_fill_1 FILLER_65_77 ();
 sg13g2_decap_4 FILLER_65_86 ();
 sg13g2_fill_1 FILLER_65_103 ();
 sg13g2_fill_2 FILLER_65_110 ();
 sg13g2_fill_1 FILLER_65_112 ();
 sg13g2_fill_1 FILLER_65_150 ();
 sg13g2_fill_2 FILLER_65_203 ();
 sg13g2_fill_1 FILLER_65_205 ();
 sg13g2_fill_2 FILLER_65_232 ();
 sg13g2_fill_2 FILLER_65_242 ();
 sg13g2_fill_1 FILLER_65_286 ();
 sg13g2_fill_2 FILLER_65_302 ();
 sg13g2_fill_1 FILLER_65_330 ();
 sg13g2_fill_1 FILLER_65_344 ();
 sg13g2_fill_1 FILLER_65_353 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_4 FILLER_66_70 ();
 sg13g2_fill_1 FILLER_66_74 ();
 sg13g2_fill_1 FILLER_66_93 ();
 sg13g2_fill_1 FILLER_66_100 ();
 sg13g2_fill_1 FILLER_66_107 ();
 sg13g2_fill_2 FILLER_66_119 ();
 sg13g2_fill_1 FILLER_66_121 ();
 sg13g2_fill_1 FILLER_66_153 ();
 sg13g2_fill_2 FILLER_66_159 ();
 sg13g2_fill_1 FILLER_66_161 ();
 sg13g2_fill_1 FILLER_66_171 ();
 sg13g2_fill_2 FILLER_66_177 ();
 sg13g2_fill_2 FILLER_66_199 ();
 sg13g2_fill_2 FILLER_66_206 ();
 sg13g2_fill_2 FILLER_66_213 ();
 sg13g2_fill_1 FILLER_66_215 ();
 sg13g2_fill_1 FILLER_66_269 ();
 sg13g2_fill_2 FILLER_66_292 ();
 sg13g2_fill_1 FILLER_66_294 ();
 sg13g2_fill_1 FILLER_66_355 ();
 sg13g2_fill_1 FILLER_66_364 ();
 sg13g2_fill_1 FILLER_66_392 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_fill_2 FILLER_67_77 ();
 sg13g2_fill_1 FILLER_67_79 ();
 sg13g2_fill_1 FILLER_67_108 ();
 sg13g2_fill_2 FILLER_67_129 ();
 sg13g2_fill_2 FILLER_67_141 ();
 sg13g2_fill_2 FILLER_67_161 ();
 sg13g2_fill_1 FILLER_67_163 ();
 sg13g2_fill_2 FILLER_67_302 ();
 sg13g2_fill_1 FILLER_67_304 ();
 sg13g2_fill_1 FILLER_67_339 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_fill_2 FILLER_68_99 ();
 sg13g2_fill_1 FILLER_68_130 ();
 sg13g2_fill_2 FILLER_68_139 ();
 sg13g2_fill_1 FILLER_68_141 ();
 sg13g2_fill_2 FILLER_68_151 ();
 sg13g2_fill_2 FILLER_68_158 ();
 sg13g2_fill_1 FILLER_68_160 ();
 sg13g2_fill_1 FILLER_68_166 ();
 sg13g2_fill_2 FILLER_68_176 ();
 sg13g2_fill_1 FILLER_68_178 ();
 sg13g2_fill_2 FILLER_68_197 ();
 sg13g2_fill_2 FILLER_68_216 ();
 sg13g2_fill_2 FILLER_68_223 ();
 sg13g2_fill_1 FILLER_68_225 ();
 sg13g2_fill_1 FILLER_68_254 ();
 sg13g2_fill_1 FILLER_68_269 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_4 FILLER_69_77 ();
 sg13g2_fill_1 FILLER_69_81 ();
 sg13g2_fill_1 FILLER_69_86 ();
 sg13g2_fill_2 FILLER_69_121 ();
 sg13g2_fill_2 FILLER_69_152 ();
 sg13g2_fill_2 FILLER_69_162 ();
 sg13g2_fill_1 FILLER_69_164 ();
 sg13g2_fill_1 FILLER_69_180 ();
 sg13g2_fill_2 FILLER_69_233 ();
 sg13g2_fill_1 FILLER_69_274 ();
 sg13g2_fill_1 FILLER_69_284 ();
 sg13g2_fill_2 FILLER_69_329 ();
 sg13g2_fill_2 FILLER_69_389 ();
 sg13g2_fill_1 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_4 FILLER_70_70 ();
 sg13g2_fill_1 FILLER_70_74 ();
 sg13g2_fill_1 FILLER_70_100 ();
 sg13g2_fill_1 FILLER_70_105 ();
 sg13g2_fill_1 FILLER_70_119 ();
 sg13g2_fill_2 FILLER_70_149 ();
 sg13g2_fill_1 FILLER_70_160 ();
 sg13g2_fill_2 FILLER_70_179 ();
 sg13g2_fill_1 FILLER_70_181 ();
 sg13g2_fill_1 FILLER_70_187 ();
 sg13g2_fill_2 FILLER_70_204 ();
 sg13g2_fill_2 FILLER_70_284 ();
 sg13g2_fill_2 FILLER_70_315 ();
 sg13g2_fill_1 FILLER_70_317 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_fill_2 FILLER_71_77 ();
 sg13g2_fill_2 FILLER_71_108 ();
 sg13g2_fill_1 FILLER_71_120 ();
 sg13g2_fill_2 FILLER_71_153 ();
 sg13g2_fill_1 FILLER_71_169 ();
 sg13g2_fill_2 FILLER_71_187 ();
 sg13g2_fill_1 FILLER_71_189 ();
 sg13g2_fill_1 FILLER_71_216 ();
 sg13g2_fill_2 FILLER_71_241 ();
 sg13g2_fill_2 FILLER_71_300 ();
 sg13g2_fill_1 FILLER_71_302 ();
 sg13g2_fill_1 FILLER_71_317 ();
 sg13g2_fill_2 FILLER_71_347 ();
 sg13g2_fill_2 FILLER_71_380 ();
 sg13g2_fill_1 FILLER_71_391 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_4 FILLER_72_70 ();
 sg13g2_fill_2 FILLER_72_74 ();
 sg13g2_fill_1 FILLER_72_91 ();
 sg13g2_fill_2 FILLER_72_144 ();
 sg13g2_fill_1 FILLER_72_154 ();
 sg13g2_fill_2 FILLER_72_178 ();
 sg13g2_fill_2 FILLER_72_253 ();
 sg13g2_fill_1 FILLER_72_314 ();
 sg13g2_fill_2 FILLER_72_367 ();
 sg13g2_fill_2 FILLER_72_380 ();
 sg13g2_fill_1 FILLER_72_382 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_4 FILLER_73_70 ();
 sg13g2_fill_1 FILLER_73_130 ();
 sg13g2_fill_1 FILLER_73_139 ();
 sg13g2_fill_2 FILLER_73_148 ();
 sg13g2_fill_1 FILLER_73_150 ();
 sg13g2_fill_2 FILLER_73_174 ();
 sg13g2_fill_2 FILLER_73_205 ();
 sg13g2_fill_1 FILLER_73_224 ();
 sg13g2_fill_2 FILLER_73_234 ();
 sg13g2_fill_1 FILLER_73_236 ();
 sg13g2_fill_1 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_fill_2 FILLER_74_63 ();
 sg13g2_fill_1 FILLER_74_65 ();
 sg13g2_fill_1 FILLER_74_100 ();
 sg13g2_fill_2 FILLER_74_157 ();
 sg13g2_fill_2 FILLER_74_181 ();
 sg13g2_fill_1 FILLER_74_183 ();
 sg13g2_fill_2 FILLER_74_234 ();
 sg13g2_fill_2 FILLER_74_253 ();
 sg13g2_fill_1 FILLER_74_255 ();
 sg13g2_fill_1 FILLER_74_313 ();
 sg13g2_fill_2 FILLER_74_380 ();
 sg13g2_fill_1 FILLER_74_382 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_fill_2 FILLER_75_70 ();
 sg13g2_fill_1 FILLER_75_72 ();
 sg13g2_fill_1 FILLER_75_105 ();
 sg13g2_fill_1 FILLER_75_122 ();
 sg13g2_fill_2 FILLER_75_152 ();
 sg13g2_fill_1 FILLER_75_154 ();
 sg13g2_fill_1 FILLER_75_189 ();
 sg13g2_fill_1 FILLER_75_205 ();
 sg13g2_fill_1 FILLER_75_268 ();
 sg13g2_fill_1 FILLER_75_346 ();
 sg13g2_fill_2 FILLER_75_356 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_fill_2 FILLER_76_108 ();
 sg13g2_fill_2 FILLER_76_149 ();
 sg13g2_fill_2 FILLER_76_268 ();
 sg13g2_fill_1 FILLER_76_270 ();
 sg13g2_fill_2 FILLER_76_322 ();
 sg13g2_fill_2 FILLER_76_333 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_fill_2 FILLER_77_77 ();
 sg13g2_fill_1 FILLER_77_123 ();
 sg13g2_fill_1 FILLER_77_132 ();
 sg13g2_fill_2 FILLER_77_172 ();
 sg13g2_fill_1 FILLER_77_174 ();
 sg13g2_fill_2 FILLER_77_181 ();
 sg13g2_fill_1 FILLER_77_183 ();
 sg13g2_fill_1 FILLER_77_218 ();
 sg13g2_fill_1 FILLER_77_266 ();
 sg13g2_fill_1 FILLER_77_305 ();
 sg13g2_fill_1 FILLER_77_346 ();
 sg13g2_fill_1 FILLER_77_355 ();
 sg13g2_fill_1 FILLER_77_369 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_fill_2 FILLER_78_77 ();
 sg13g2_fill_2 FILLER_78_264 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_4 FILLER_79_70 ();
 sg13g2_fill_2 FILLER_79_159 ();
 sg13g2_fill_2 FILLER_79_181 ();
 sg13g2_fill_2 FILLER_79_254 ();
 sg13g2_fill_1 FILLER_79_261 ();
 sg13g2_fill_2 FILLER_79_326 ();
 sg13g2_fill_2 FILLER_79_347 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_fill_1 FILLER_80_76 ();
 sg13g2_fill_2 FILLER_80_118 ();
 sg13g2_fill_1 FILLER_80_378 ();
 sg13g2_fill_2 FILLER_80_406 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net100;
 assign uio_oe[1] = net101;
 assign uio_oe[2] = net102;
 assign uio_oe[3] = net103;
 assign uio_oe[4] = net104;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
 assign uio_out[2] = net16;
 assign uio_out[3] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
endmodule
