module tt_um_pwm_block (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \MemCell.counter[0] ;
 wire \MemCell.counter[1] ;
 wire \MemCell.counter_value[0] ;
 wire \MemCell.counter_value[10] ;
 wire \MemCell.counter_value[11] ;
 wire \MemCell.counter_value[12] ;
 wire \MemCell.counter_value[13] ;
 wire \MemCell.counter_value[14] ;
 wire \MemCell.counter_value[15] ;
 wire \MemCell.counter_value[16] ;
 wire \MemCell.counter_value[17] ;
 wire \MemCell.counter_value[18] ;
 wire \MemCell.counter_value[19] ;
 wire \MemCell.counter_value[1] ;
 wire \MemCell.counter_value[20] ;
 wire \MemCell.counter_value[21] ;
 wire \MemCell.counter_value[22] ;
 wire \MemCell.counter_value[23] ;
 wire \MemCell.counter_value[24] ;
 wire \MemCell.counter_value[25] ;
 wire \MemCell.counter_value[26] ;
 wire \MemCell.counter_value[27] ;
 wire \MemCell.counter_value[28] ;
 wire \MemCell.counter_value[29] ;
 wire \MemCell.counter_value[2] ;
 wire \MemCell.counter_value[30] ;
 wire \MemCell.counter_value[31] ;
 wire \MemCell.counter_value[3] ;
 wire \MemCell.counter_value[4] ;
 wire \MemCell.counter_value[5] ;
 wire \MemCell.counter_value[6] ;
 wire \MemCell.counter_value[7] ;
 wire \MemCell.counter_value[8] ;
 wire \MemCell.counter_value[9] ;
 wire \MemCell.curr_state[0] ;
 wire \MemCell.curr_state[1] ;
 wire \MemCell.curr_state[2] ;
 wire \MemCell.dc1_reg[0][0] ;
 wire \MemCell.dc1_reg[0][1] ;
 wire \MemCell.dc1_reg[0][2] ;
 wire \MemCell.dc1_reg[0][3] ;
 wire \MemCell.dc1_reg[0][4] ;
 wire \MemCell.dc1_reg[0][5] ;
 wire \MemCell.dc1_reg[0][6] ;
 wire \MemCell.dc1_reg[0][7] ;
 wire \MemCell.dc1_reg[1][0] ;
 wire \MemCell.dc1_reg[1][1] ;
 wire \MemCell.dc1_reg[1][2] ;
 wire \MemCell.dc1_reg[1][3] ;
 wire \MemCell.dc1_reg[1][4] ;
 wire \MemCell.dc1_reg[1][5] ;
 wire \MemCell.dc1_reg[1][6] ;
 wire \MemCell.dc1_reg[1][7] ;
 wire \MemCell.dc1_reg[2][0] ;
 wire \MemCell.dc1_reg[2][1] ;
 wire \MemCell.dc1_reg[2][2] ;
 wire \MemCell.dc1_reg[2][3] ;
 wire \MemCell.dc1_reg[2][4] ;
 wire \MemCell.dc1_reg[2][5] ;
 wire \MemCell.dc1_reg[2][6] ;
 wire \MemCell.dc1_reg[2][7] ;
 wire \MemCell.dc1_reg[3][0] ;
 wire \MemCell.dc1_reg[3][1] ;
 wire \MemCell.dc1_reg[3][2] ;
 wire \MemCell.dc1_reg[3][3] ;
 wire \MemCell.dc1_reg[3][4] ;
 wire \MemCell.dc1_reg[3][5] ;
 wire \MemCell.dc1_reg[3][6] ;
 wire \MemCell.dc1_reg[3][7] ;
 wire \MemCell.dc2_reg[0][0] ;
 wire \MemCell.dc2_reg[0][1] ;
 wire \MemCell.dc2_reg[0][2] ;
 wire \MemCell.dc2_reg[0][3] ;
 wire \MemCell.dc2_reg[0][4] ;
 wire \MemCell.dc2_reg[0][5] ;
 wire \MemCell.dc2_reg[0][6] ;
 wire \MemCell.dc2_reg[0][7] ;
 wire \MemCell.dc2_reg[1][0] ;
 wire \MemCell.dc2_reg[1][1] ;
 wire \MemCell.dc2_reg[1][2] ;
 wire \MemCell.dc2_reg[1][3] ;
 wire \MemCell.dc2_reg[1][4] ;
 wire \MemCell.dc2_reg[1][5] ;
 wire \MemCell.dc2_reg[1][6] ;
 wire \MemCell.dc2_reg[1][7] ;
 wire \MemCell.dc2_reg[2][0] ;
 wire \MemCell.dc2_reg[2][1] ;
 wire \MemCell.dc2_reg[2][2] ;
 wire \MemCell.dc2_reg[2][3] ;
 wire \MemCell.dc2_reg[2][4] ;
 wire \MemCell.dc2_reg[2][5] ;
 wire \MemCell.dc2_reg[2][6] ;
 wire \MemCell.dc2_reg[2][7] ;
 wire \MemCell.dc2_reg[3][0] ;
 wire \MemCell.dc2_reg[3][1] ;
 wire \MemCell.dc2_reg[3][2] ;
 wire \MemCell.dc2_reg[3][3] ;
 wire \MemCell.dc2_reg[3][4] ;
 wire \MemCell.dc2_reg[3][5] ;
 wire \MemCell.dc2_reg[3][6] ;
 wire \MemCell.dc2_reg[3][7] ;
 wire \MemCell.dc3_reg[0][0] ;
 wire \MemCell.dc3_reg[0][1] ;
 wire \MemCell.dc3_reg[0][2] ;
 wire \MemCell.dc3_reg[0][3] ;
 wire \MemCell.dc3_reg[0][4] ;
 wire \MemCell.dc3_reg[0][5] ;
 wire \MemCell.dc3_reg[0][6] ;
 wire \MemCell.dc3_reg[0][7] ;
 wire \MemCell.dc3_reg[1][0] ;
 wire \MemCell.dc3_reg[1][1] ;
 wire \MemCell.dc3_reg[1][2] ;
 wire \MemCell.dc3_reg[1][3] ;
 wire \MemCell.dc3_reg[1][4] ;
 wire \MemCell.dc3_reg[1][5] ;
 wire \MemCell.dc3_reg[1][6] ;
 wire \MemCell.dc3_reg[1][7] ;
 wire \MemCell.dc3_reg[2][0] ;
 wire \MemCell.dc3_reg[2][1] ;
 wire \MemCell.dc3_reg[2][2] ;
 wire \MemCell.dc3_reg[2][3] ;
 wire \MemCell.dc3_reg[2][4] ;
 wire \MemCell.dc3_reg[2][5] ;
 wire \MemCell.dc3_reg[2][6] ;
 wire \MemCell.dc3_reg[2][7] ;
 wire \MemCell.dc3_reg[3][0] ;
 wire \MemCell.dc3_reg[3][1] ;
 wire \MemCell.dc3_reg[3][2] ;
 wire \MemCell.dc3_reg[3][3] ;
 wire \MemCell.dc3_reg[3][4] ;
 wire \MemCell.dc3_reg[3][5] ;
 wire \MemCell.dc3_reg[3][6] ;
 wire \MemCell.dc3_reg[3][7] ;
 wire \MemCell.enable_pwm ;
 wire \MemCell.next_state[0] ;
 wire \MemCell.next_state[1] ;
 wire \MemCell.next_state[2] ;
 wire \MemCell.o_RX_Byte[0] ;
 wire \MemCell.o_RX_Byte[1] ;
 wire \MemCell.o_RX_Byte[2] ;
 wire \MemCell.o_RX_Byte[3] ;
 wire \MemCell.o_RX_Byte[4] ;
 wire \MemCell.o_RX_Byte[5] ;
 wire \MemCell.o_RX_Byte[6] ;
 wire \MemCell.o_RX_Byte[7] ;
 wire \MemCell.o_RX_DV ;
 wire \MemCell.prescale_reg[0][0] ;
 wire \MemCell.prescale_reg[0][1] ;
 wire \MemCell.prescale_reg[0][2] ;
 wire \MemCell.prescale_reg[0][3] ;
 wire \MemCell.prescale_reg[0][4] ;
 wire \MemCell.prescale_reg[0][5] ;
 wire \MemCell.prescale_reg[0][6] ;
 wire \MemCell.prescale_reg[0][7] ;
 wire \MemCell.prescale_reg[1][0] ;
 wire \MemCell.prescale_reg[1][1] ;
 wire \MemCell.prescale_reg[1][2] ;
 wire \MemCell.prescale_reg[1][3] ;
 wire \MemCell.prescale_reg[1][4] ;
 wire \MemCell.prescale_reg[1][5] ;
 wire \MemCell.prescale_reg[1][6] ;
 wire \MemCell.prescale_reg[1][7] ;
 wire \MemCell.prescale_reg[2][0] ;
 wire \MemCell.prescale_reg[2][1] ;
 wire \MemCell.prescale_reg[2][2] ;
 wire \MemCell.prescale_reg[2][3] ;
 wire \MemCell.prescale_reg[2][4] ;
 wire \MemCell.prescale_reg[2][5] ;
 wire \MemCell.prescale_reg[2][6] ;
 wire \MemCell.prescale_reg[2][7] ;
 wire \MemCell.prescale_reg[3][0] ;
 wire \MemCell.prescale_reg[3][1] ;
 wire \MemCell.prescale_reg[3][2] ;
 wire \MemCell.prescale_reg[3][3] ;
 wire \MemCell.prescale_reg[3][4] ;
 wire \MemCell.prescale_reg[3][5] ;
 wire \MemCell.prescale_reg[3][6] ;
 wire \MemCell.prescale_reg[3][7] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire \pwm_module.counter0[0] ;
 wire \pwm_module.counter0[10] ;
 wire \pwm_module.counter0[11] ;
 wire \pwm_module.counter0[12] ;
 wire \pwm_module.counter0[13] ;
 wire \pwm_module.counter0[14] ;
 wire \pwm_module.counter0[15] ;
 wire \pwm_module.counter0[16] ;
 wire \pwm_module.counter0[17] ;
 wire \pwm_module.counter0[18] ;
 wire \pwm_module.counter0[19] ;
 wire \pwm_module.counter0[1] ;
 wire \pwm_module.counter0[20] ;
 wire \pwm_module.counter0[21] ;
 wire \pwm_module.counter0[22] ;
 wire \pwm_module.counter0[23] ;
 wire \pwm_module.counter0[24] ;
 wire \pwm_module.counter0[25] ;
 wire \pwm_module.counter0[26] ;
 wire \pwm_module.counter0[27] ;
 wire \pwm_module.counter0[28] ;
 wire \pwm_module.counter0[29] ;
 wire \pwm_module.counter0[2] ;
 wire \pwm_module.counter0[30] ;
 wire \pwm_module.counter0[31] ;
 wire \pwm_module.counter0[3] ;
 wire \pwm_module.counter0[4] ;
 wire \pwm_module.counter0[5] ;
 wire \pwm_module.counter0[6] ;
 wire \pwm_module.counter0[7] ;
 wire \pwm_module.counter0[8] ;
 wire \pwm_module.counter0[9] ;
 wire \pwm_module.counter1[0] ;
 wire \pwm_module.counter1[10] ;
 wire \pwm_module.counter1[11] ;
 wire \pwm_module.counter1[12] ;
 wire \pwm_module.counter1[13] ;
 wire \pwm_module.counter1[14] ;
 wire \pwm_module.counter1[15] ;
 wire \pwm_module.counter1[16] ;
 wire \pwm_module.counter1[17] ;
 wire \pwm_module.counter1[18] ;
 wire \pwm_module.counter1[19] ;
 wire \pwm_module.counter1[1] ;
 wire \pwm_module.counter1[20] ;
 wire \pwm_module.counter1[21] ;
 wire \pwm_module.counter1[22] ;
 wire \pwm_module.counter1[23] ;
 wire \pwm_module.counter1[24] ;
 wire \pwm_module.counter1[25] ;
 wire \pwm_module.counter1[26] ;
 wire \pwm_module.counter1[27] ;
 wire \pwm_module.counter1[28] ;
 wire \pwm_module.counter1[29] ;
 wire \pwm_module.counter1[2] ;
 wire \pwm_module.counter1[30] ;
 wire \pwm_module.counter1[31] ;
 wire \pwm_module.counter1[3] ;
 wire \pwm_module.counter1[4] ;
 wire \pwm_module.counter1[5] ;
 wire \pwm_module.counter1[6] ;
 wire \pwm_module.counter1[7] ;
 wire \pwm_module.counter1[8] ;
 wire \pwm_module.counter1[9] ;
 wire \pwm_module.counter2[0] ;
 wire \pwm_module.counter2[10] ;
 wire \pwm_module.counter2[11] ;
 wire \pwm_module.counter2[12] ;
 wire \pwm_module.counter2[13] ;
 wire \pwm_module.counter2[14] ;
 wire \pwm_module.counter2[15] ;
 wire \pwm_module.counter2[16] ;
 wire \pwm_module.counter2[17] ;
 wire \pwm_module.counter2[18] ;
 wire \pwm_module.counter2[19] ;
 wire \pwm_module.counter2[1] ;
 wire \pwm_module.counter2[20] ;
 wire \pwm_module.counter2[21] ;
 wire \pwm_module.counter2[22] ;
 wire \pwm_module.counter2[23] ;
 wire \pwm_module.counter2[24] ;
 wire \pwm_module.counter2[25] ;
 wire \pwm_module.counter2[26] ;
 wire \pwm_module.counter2[27] ;
 wire \pwm_module.counter2[28] ;
 wire \pwm_module.counter2[29] ;
 wire \pwm_module.counter2[2] ;
 wire \pwm_module.counter2[30] ;
 wire \pwm_module.counter2[31] ;
 wire \pwm_module.counter2[3] ;
 wire \pwm_module.counter2[4] ;
 wire \pwm_module.counter2[5] ;
 wire \pwm_module.counter2[6] ;
 wire \pwm_module.counter2[7] ;
 wire \pwm_module.counter2[8] ;
 wire \pwm_module.counter2[9] ;
 wire \pwm_module.prescaler0[0] ;
 wire \pwm_module.prescaler0[10] ;
 wire \pwm_module.prescaler0[11] ;
 wire \pwm_module.prescaler0[12] ;
 wire \pwm_module.prescaler0[13] ;
 wire \pwm_module.prescaler0[14] ;
 wire \pwm_module.prescaler0[15] ;
 wire \pwm_module.prescaler0[16] ;
 wire \pwm_module.prescaler0[17] ;
 wire \pwm_module.prescaler0[18] ;
 wire \pwm_module.prescaler0[19] ;
 wire \pwm_module.prescaler0[1] ;
 wire \pwm_module.prescaler0[20] ;
 wire \pwm_module.prescaler0[21] ;
 wire \pwm_module.prescaler0[22] ;
 wire \pwm_module.prescaler0[23] ;
 wire \pwm_module.prescaler0[24] ;
 wire \pwm_module.prescaler0[25] ;
 wire \pwm_module.prescaler0[26] ;
 wire \pwm_module.prescaler0[27] ;
 wire \pwm_module.prescaler0[28] ;
 wire \pwm_module.prescaler0[29] ;
 wire \pwm_module.prescaler0[2] ;
 wire \pwm_module.prescaler0[30] ;
 wire \pwm_module.prescaler0[31] ;
 wire \pwm_module.prescaler0[3] ;
 wire \pwm_module.prescaler0[4] ;
 wire \pwm_module.prescaler0[5] ;
 wire \pwm_module.prescaler0[6] ;
 wire \pwm_module.prescaler0[7] ;
 wire \pwm_module.prescaler0[8] ;
 wire \pwm_module.prescaler0[9] ;
 wire \pwm_module.prescaler1[0] ;
 wire \pwm_module.prescaler1[10] ;
 wire \pwm_module.prescaler1[11] ;
 wire \pwm_module.prescaler1[12] ;
 wire \pwm_module.prescaler1[13] ;
 wire \pwm_module.prescaler1[14] ;
 wire \pwm_module.prescaler1[15] ;
 wire \pwm_module.prescaler1[16] ;
 wire \pwm_module.prescaler1[17] ;
 wire \pwm_module.prescaler1[18] ;
 wire \pwm_module.prescaler1[19] ;
 wire \pwm_module.prescaler1[1] ;
 wire \pwm_module.prescaler1[20] ;
 wire \pwm_module.prescaler1[21] ;
 wire \pwm_module.prescaler1[22] ;
 wire \pwm_module.prescaler1[23] ;
 wire \pwm_module.prescaler1[24] ;
 wire \pwm_module.prescaler1[25] ;
 wire \pwm_module.prescaler1[26] ;
 wire \pwm_module.prescaler1[27] ;
 wire \pwm_module.prescaler1[28] ;
 wire \pwm_module.prescaler1[29] ;
 wire \pwm_module.prescaler1[2] ;
 wire \pwm_module.prescaler1[30] ;
 wire \pwm_module.prescaler1[31] ;
 wire \pwm_module.prescaler1[3] ;
 wire \pwm_module.prescaler1[4] ;
 wire \pwm_module.prescaler1[5] ;
 wire \pwm_module.prescaler1[6] ;
 wire \pwm_module.prescaler1[7] ;
 wire \pwm_module.prescaler1[8] ;
 wire \pwm_module.prescaler1[9] ;
 wire \pwm_module.prescaler2[0] ;
 wire \pwm_module.prescaler2[10] ;
 wire \pwm_module.prescaler2[11] ;
 wire \pwm_module.prescaler2[12] ;
 wire \pwm_module.prescaler2[13] ;
 wire \pwm_module.prescaler2[14] ;
 wire \pwm_module.prescaler2[15] ;
 wire \pwm_module.prescaler2[16] ;
 wire \pwm_module.prescaler2[17] ;
 wire \pwm_module.prescaler2[18] ;
 wire \pwm_module.prescaler2[19] ;
 wire \pwm_module.prescaler2[1] ;
 wire \pwm_module.prescaler2[20] ;
 wire \pwm_module.prescaler2[21] ;
 wire \pwm_module.prescaler2[22] ;
 wire \pwm_module.prescaler2[23] ;
 wire \pwm_module.prescaler2[24] ;
 wire \pwm_module.prescaler2[25] ;
 wire \pwm_module.prescaler2[26] ;
 wire \pwm_module.prescaler2[27] ;
 wire \pwm_module.prescaler2[28] ;
 wire \pwm_module.prescaler2[29] ;
 wire \pwm_module.prescaler2[2] ;
 wire \pwm_module.prescaler2[30] ;
 wire \pwm_module.prescaler2[31] ;
 wire \pwm_module.prescaler2[3] ;
 wire \pwm_module.prescaler2[4] ;
 wire \pwm_module.prescaler2[5] ;
 wire \pwm_module.prescaler2[6] ;
 wire \pwm_module.prescaler2[7] ;
 wire \pwm_module.prescaler2[8] ;
 wire \pwm_module.prescaler2[9] ;
 wire reg_ui0;
 wire reg_ui1;
 wire \spi_module.r2_RX_Done ;
 wire \spi_module.r3_RX_Done ;
 wire \spi_module.r_RX_Bit_Count[0] ;
 wire \spi_module.r_RX_Bit_Count[1] ;
 wire \spi_module.r_RX_Bit_Count[2] ;
 wire \spi_module.r_RX_Byte[0] ;
 wire \spi_module.r_RX_Byte[1] ;
 wire \spi_module.r_RX_Byte[2] ;
 wire \spi_module.r_RX_Byte[3] ;
 wire \spi_module.r_RX_Byte[4] ;
 wire \spi_module.r_RX_Byte[5] ;
 wire \spi_module.r_RX_Byte[6] ;
 wire \spi_module.r_RX_Byte[7] ;
 wire \spi_module.r_RX_Done ;
 wire \spi_module.r_Temp_RX_Byte[0] ;
 wire \spi_module.r_Temp_RX_Byte[1] ;
 wire \spi_module.r_Temp_RX_Byte[2] ;
 wire \spi_module.r_Temp_RX_Byte[3] ;
 wire \spi_module.r_Temp_RX_Byte[4] ;
 wire \spi_module.r_Temp_RX_Byte[5] ;
 wire \spi_module.r_Temp_RX_Byte[6] ;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net7;
 wire clknet_leaf_0_clk;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;

 sg13g2_inv_1 _2689_ (.Y(_2313_),
    .A(net391));
 sg13g2_inv_1 _2690_ (.Y(_2314_),
    .A(\pwm_module.prescaler1[22] ));
 sg13g2_inv_1 _2691_ (.Y(_2315_),
    .A(net464));
 sg13g2_inv_1 _2692_ (.Y(_2316_),
    .A(net442));
 sg13g2_inv_1 _2693_ (.Y(_2317_),
    .A(net505));
 sg13g2_inv_1 _2694_ (.Y(_2318_),
    .A(\pwm_module.counter2[2] ));
 sg13g2_inv_1 _2695_ (.Y(_2319_),
    .A(\pwm_module.counter2[5] ));
 sg13g2_inv_1 _2696_ (.Y(_2320_),
    .A(\pwm_module.counter2[4] ));
 sg13g2_inv_1 _2697_ (.Y(_2321_),
    .A(\pwm_module.counter2[14] ));
 sg13g2_inv_1 _2698_ (.Y(_2322_),
    .A(\pwm_module.counter2[13] ));
 sg13g2_inv_1 _2699_ (.Y(_2323_),
    .A(net89));
 sg13g2_inv_1 _2700_ (.Y(_2324_),
    .A(_0131_));
 sg13g2_inv_1 _2701_ (.Y(_2325_),
    .A(net528));
 sg13g2_inv_1 _2702_ (.Y(_2326_),
    .A(_0127_));
 sg13g2_inv_1 _2703_ (.Y(_2327_),
    .A(net481));
 sg13g2_inv_1 _2704_ (.Y(_2328_),
    .A(_0128_));
 sg13g2_inv_1 _2705_ (.Y(_2329_),
    .A(_0129_));
 sg13g2_inv_1 _2706_ (.Y(_2330_),
    .A(net522));
 sg13g2_inv_1 _2707_ (.Y(_2331_),
    .A(_0126_));
 sg13g2_inv_1 _2708_ (.Y(_2332_),
    .A(net184));
 sg13g2_inv_1 _2709_ (.Y(_2333_),
    .A(_0189_));
 sg13g2_inv_1 _2710_ (.Y(_2334_),
    .A(\pwm_module.prescaler2[10] ));
 sg13g2_inv_1 _2711_ (.Y(_2335_),
    .A(_0190_));
 sg13g2_inv_1 _2712_ (.Y(_2336_),
    .A(_0194_));
 sg13g2_inv_1 _2713_ (.Y(_2337_),
    .A(_0197_));
 sg13g2_inv_1 _2714_ (.Y(_2338_),
    .A(\pwm_module.prescaler2[22] ));
 sg13g2_inv_1 _2715_ (.Y(_2339_),
    .A(net410));
 sg13g2_inv_1 _2716_ (.Y(_2340_),
    .A(net512));
 sg13g2_inv_1 _2717_ (.Y(_2341_),
    .A(net572));
 sg13g2_inv_1 _2718_ (.Y(_2342_),
    .A(net244));
 sg13g2_inv_1 _2719_ (.Y(_2343_),
    .A(net575));
 sg13g2_inv_1 _2720_ (.Y(_2344_),
    .A(\MemCell.o_RX_Byte[1] ));
 sg13g2_inv_1 _2721_ (.Y(_2345_),
    .A(\MemCell.o_RX_Byte[2] ));
 sg13g2_inv_1 _2722_ (.Y(_2346_),
    .A(\MemCell.o_RX_DV ));
 sg13g2_inv_2 _2723_ (.Y(_2347_),
    .A(net3));
 sg13g2_inv_1 _2724_ (.Y(_2348_),
    .A(net483));
 sg13g2_inv_1 _2725_ (.Y(_2349_),
    .A(net552));
 sg13g2_inv_1 _2726_ (.Y(_2350_),
    .A(net564));
 sg13g2_inv_1 _2727_ (.Y(_2351_),
    .A(\pwm_module.counter0[22] ));
 sg13g2_inv_2 _2728_ (.Y(_2352_),
    .A(net525));
 sg13g2_inv_1 _2729_ (.Y(_2353_),
    .A(net554));
 sg13g2_inv_1 _2730_ (.Y(_2354_),
    .A(\pwm_module.counter0[12] ));
 sg13g2_inv_1 _2731_ (.Y(_2355_),
    .A(_0164_));
 sg13g2_inv_1 _2732_ (.Y(_2356_),
    .A(net774));
 sg13g2_inv_1 _2733_ (.Y(_2357_),
    .A(net308));
 sg13g2_inv_1 _2734_ (.Y(_2358_),
    .A(net390));
 sg13g2_inv_1 _2735_ (.Y(_2359_),
    .A(_0105_));
 sg13g2_inv_1 _2736_ (.Y(_2360_),
    .A(\pwm_module.counter1[22] ));
 sg13g2_inv_1 _2737_ (.Y(_2361_),
    .A(_0107_));
 sg13g2_inv_1 _2738_ (.Y(_2362_),
    .A(\pwm_module.counter1[21] ));
 sg13g2_inv_1 _2739_ (.Y(_2363_),
    .A(_0112_));
 sg13g2_inv_1 _2740_ (.Y(_2364_),
    .A(net549));
 sg13g2_inv_1 _2741_ (.Y(_2365_),
    .A(\pwm_module.counter1[6] ));
 sg13g2_inv_1 _2742_ (.Y(_2366_),
    .A(net477));
 sg13g2_inv_2 _2743_ (.Y(_2367_),
    .A(net441));
 sg13g2_inv_1 _2744_ (.Y(_2368_),
    .A(net551));
 sg13g2_inv_1 _2745_ (.Y(_2369_),
    .A(_0122_));
 sg13g2_inv_1 _2746_ (.Y(_2370_),
    .A(net770));
 sg13g2_inv_1 _2747_ (.Y(_2371_),
    .A(\MemCell.dc3_reg[2][2] ));
 sg13g2_inv_1 _2748_ (.Y(_2372_),
    .A(net337));
 sg13g2_inv_1 _2749_ (.Y(_2373_),
    .A(\MemCell.enable_pwm ));
 sg13g2_inv_1 _2750_ (.Y(_2374_),
    .A(\pwm_module.prescaler1[6] ));
 sg13g2_inv_1 _2751_ (.Y(_2375_),
    .A(\pwm_module.prescaler1[14] ));
 sg13g2_inv_1 _2752_ (.Y(_2376_),
    .A(_0172_));
 sg13g2_inv_1 _2753_ (.Y(_2377_),
    .A(net379));
 sg13g2_inv_1 _2754_ (.Y(_2378_),
    .A(net270));
 sg13g2_inv_1 _2755_ (.Y(_2379_),
    .A(\pwm_module.prescaler0[6] ));
 sg13g2_inv_1 _2756_ (.Y(_2380_),
    .A(net405));
 sg13g2_inv_1 _2757_ (.Y(_2381_),
    .A(_0206_));
 sg13g2_inv_1 _2758_ (.Y(_2382_),
    .A(\pwm_module.prescaler0[11] ));
 sg13g2_inv_1 _2759_ (.Y(_2383_),
    .A(_0207_));
 sg13g2_inv_1 _2760_ (.Y(_2384_),
    .A(\pwm_module.prescaler0[10] ));
 sg13g2_inv_1 _2761_ (.Y(_2385_),
    .A(net526));
 sg13g2_inv_1 _2762_ (.Y(_2386_),
    .A(\pwm_module.prescaler0[22] ));
 sg13g2_inv_1 _2763_ (.Y(_2387_),
    .A(\pwm_module.prescaler0[16] ));
 sg13g2_inv_1 _2764_ (.Y(_0219_),
    .A(net763));
 sg13g2_inv_1 _2765_ (.Y(_2388_),
    .A(net50));
 sg13g2_inv_1 _2766_ (.Y(_2389_),
    .A(net247));
 sg13g2_inv_1 _2767_ (.Y(_2390_),
    .A(net152));
 sg13g2_inv_1 _2768_ (.Y(_2391_),
    .A(net58));
 sg13g2_inv_1 _2769_ (.Y(_2397_),
    .A(_0166_));
 sg13g2_nand2b_1 _2770_ (.Y(_2392_),
    .B(\spi_module.r_RX_Bit_Count[1] ),
    .A_N(\spi_module.r_RX_Bit_Count[0] ));
 sg13g2_nand3_1 _2771_ (.B(\spi_module.r_RX_Bit_Count[0] ),
    .C(\spi_module.r_RX_Bit_Count[2] ),
    .A(\spi_module.r_RX_Bit_Count[1] ),
    .Y(_2393_));
 sg13g2_o21ai_1 _2772_ (.B1(\spi_module.r_RX_Done ),
    .Y(_2394_),
    .A1(\spi_module.r_RX_Bit_Count[2] ),
    .A2(_2392_));
 sg13g2_nand2_1 _2773_ (.Y(_0278_),
    .A(_2393_),
    .B(_2394_));
 sg13g2_nor2_2 _2774_ (.A(net4),
    .B(\MemCell.enable_pwm ),
    .Y(_2395_));
 sg13g2_or2_2 _2775_ (.X(_2396_),
    .B(\MemCell.enable_pwm ),
    .A(net4));
 sg13g2_nand2b_2 _2776_ (.Y(_0506_),
    .B(\MemCell.prescale_reg[3][6] ),
    .A_N(net786));
 sg13g2_xnor2_1 _2777_ (.Y(_0507_),
    .A(\pwm_module.prescaler1[30] ),
    .B(_0506_));
 sg13g2_nor2b_2 _2778_ (.A(net786),
    .B_N(\MemCell.prescale_reg[3][5] ),
    .Y(_0508_));
 sg13g2_nor2_1 _2779_ (.A(_0184_),
    .B(_0508_),
    .Y(_0509_));
 sg13g2_nor2b_1 _2780_ (.A(net786),
    .B_N(\MemCell.prescale_reg[3][7] ),
    .Y(_0510_));
 sg13g2_nor2_1 _2781_ (.A(_0185_),
    .B(net719),
    .Y(_0511_));
 sg13g2_nor3_1 _2782_ (.A(_0507_),
    .B(_0509_),
    .C(_0511_),
    .Y(_0512_));
 sg13g2_nor2b_2 _2783_ (.A(net786),
    .B_N(\MemCell.prescale_reg[3][4] ),
    .Y(_0513_));
 sg13g2_nand2b_2 _2784_ (.Y(_0514_),
    .B(\MemCell.prescale_reg[3][4] ),
    .A_N(net786));
 sg13g2_a22oi_1 _2785_ (.Y(_0515_),
    .B1(_0513_),
    .B2(_2316_),
    .A2(_0508_),
    .A1(_0184_));
 sg13g2_inv_1 _2786_ (.Y(_0516_),
    .A(_0515_));
 sg13g2_nor2b_1 _2787_ (.A(net785),
    .B_N(\MemCell.prescale_reg[3][0] ),
    .Y(_0517_));
 sg13g2_nand2b_2 _2788_ (.Y(_0518_),
    .B(\MemCell.prescale_reg[3][0] ),
    .A_N(net785));
 sg13g2_nor2b_2 _2789_ (.A(net785),
    .B_N(\MemCell.prescale_reg[3][1] ),
    .Y(_0519_));
 sg13g2_nand2b_2 _2790_ (.Y(_0520_),
    .B(\MemCell.prescale_reg[3][1] ),
    .A_N(net785));
 sg13g2_nand3b_1 _2791_ (.B(\MemCell.prescale_reg[3][1] ),
    .C(_0182_),
    .Y(_0521_),
    .A_N(net786));
 sg13g2_o21ai_1 _2792_ (.B1(_0521_),
    .Y(_0522_),
    .A1(\pwm_module.prescaler1[24] ),
    .A2(_0518_));
 sg13g2_nor2b_2 _2793_ (.A(net785),
    .B_N(\MemCell.prescale_reg[3][2] ),
    .Y(_0523_));
 sg13g2_nand2b_1 _2794_ (.Y(_0524_),
    .B(\MemCell.prescale_reg[3][2] ),
    .A_N(net785));
 sg13g2_nor2_1 _2795_ (.A(\pwm_module.prescaler1[26] ),
    .B(_0524_),
    .Y(_0525_));
 sg13g2_xnor2_1 _2796_ (.Y(_0526_),
    .A(\pwm_module.prescaler1[26] ),
    .B(_0523_));
 sg13g2_nor2b_2 _2797_ (.A(net785),
    .B_N(\MemCell.prescale_reg[3][3] ),
    .Y(_0527_));
 sg13g2_nand2b_2 _2798_ (.Y(_0528_),
    .B(\MemCell.prescale_reg[3][3] ),
    .A_N(net785));
 sg13g2_nand2b_1 _2799_ (.Y(_0529_),
    .B(_0528_),
    .A_N(_0183_));
 sg13g2_nand2_1 _2800_ (.Y(_0530_),
    .A(_2315_),
    .B(_0520_));
 sg13g2_nand4_1 _2801_ (.B(_0526_),
    .C(_0529_),
    .A(_0522_),
    .Y(_0531_),
    .D(_0530_));
 sg13g2_and2_1 _2802_ (.A(_0183_),
    .B(_0527_),
    .X(_0532_));
 sg13g2_nand2_1 _2803_ (.Y(_0533_),
    .A(_0183_),
    .B(_0527_));
 sg13g2_a21oi_1 _2804_ (.A1(_0525_),
    .A2(_0529_),
    .Y(_0534_),
    .B1(_0532_));
 sg13g2_a22oi_1 _2805_ (.Y(_0535_),
    .B1(_0531_),
    .B2(_0534_),
    .A2(_0514_),
    .A1(\pwm_module.prescaler1[28] ));
 sg13g2_o21ai_1 _2806_ (.B1(_0512_),
    .Y(_0536_),
    .A1(_0516_),
    .A2(_0535_));
 sg13g2_a22oi_1 _2807_ (.Y(_0537_),
    .B1(_0520_),
    .B2(_2315_),
    .A2(net719),
    .A1(_0185_));
 sg13g2_and4_1 _2808_ (.A(_0526_),
    .B(_0529_),
    .C(_0533_),
    .D(_0537_),
    .X(_0538_));
 sg13g2_a221oi_1 _2809_ (.B2(\pwm_module.prescaler1[24] ),
    .C1(_0522_),
    .B1(_0518_),
    .A1(\pwm_module.prescaler1[28] ),
    .Y(_0539_),
    .A2(_0514_));
 sg13g2_nand4_1 _2810_ (.B(_0515_),
    .C(_0538_),
    .A(_0512_),
    .Y(_0540_),
    .D(_0539_));
 sg13g2_nor2b_1 _2811_ (.A(net784),
    .B_N(\MemCell.prescale_reg[2][6] ),
    .Y(_0541_));
 sg13g2_nand2b_2 _2812_ (.Y(_0542_),
    .B(\MemCell.prescale_reg[2][6] ),
    .A_N(net783));
 sg13g2_nor2b_2 _2813_ (.A(net784),
    .B_N(\MemCell.prescale_reg[2][7] ),
    .Y(_0543_));
 sg13g2_a22oi_1 _2814_ (.Y(_0544_),
    .B1(_0543_),
    .B2(_0181_),
    .A2(_0541_),
    .A1(_2314_));
 sg13g2_or2_1 _2815_ (.X(_0545_),
    .B(_0543_),
    .A(_0181_));
 sg13g2_nor2b_1 _2816_ (.A(net783),
    .B_N(\MemCell.prescale_reg[2][5] ),
    .Y(_0546_));
 sg13g2_nand2b_2 _2817_ (.Y(_0547_),
    .B(\MemCell.prescale_reg[2][5] ),
    .A_N(net784));
 sg13g2_a22oi_1 _2818_ (.Y(_0548_),
    .B1(_0547_),
    .B2(_2313_),
    .A2(_0542_),
    .A1(\pwm_module.prescaler1[22] ));
 sg13g2_and3_1 _2819_ (.X(_0549_),
    .A(_0544_),
    .B(_0545_),
    .C(_0548_));
 sg13g2_nor2b_2 _2820_ (.A(net783),
    .B_N(\MemCell.prescale_reg[2][4] ),
    .Y(_0550_));
 sg13g2_a22oi_1 _2821_ (.Y(_0551_),
    .B1(_0550_),
    .B2(_0179_),
    .A2(_0546_),
    .A1(_0180_));
 sg13g2_inv_1 _2822_ (.Y(_0552_),
    .A(_0551_));
 sg13g2_nor2_1 _2823_ (.A(_0179_),
    .B(_0550_),
    .Y(_0553_));
 sg13g2_nand4_1 _2824_ (.B(_0545_),
    .C(_0548_),
    .A(_0544_),
    .Y(_0554_),
    .D(_0551_));
 sg13g2_or2_1 _2825_ (.X(_0555_),
    .B(_0554_),
    .A(_0553_));
 sg13g2_nor2b_2 _2826_ (.A(net783),
    .B_N(\MemCell.prescale_reg[2][3] ),
    .Y(_0556_));
 sg13g2_nand2b_1 _2827_ (.Y(_0557_),
    .B(\MemCell.prescale_reg[2][3] ),
    .A_N(net783));
 sg13g2_nand3b_1 _2828_ (.B(\MemCell.prescale_reg[2][3] ),
    .C(_0178_),
    .Y(_0558_),
    .A_N(net784));
 sg13g2_nand2b_2 _2829_ (.Y(_0559_),
    .B(\MemCell.prescale_reg[2][2] ),
    .A_N(net783));
 sg13g2_o21ai_1 _2830_ (.B1(_0558_),
    .Y(_0560_),
    .A1(\pwm_module.prescaler1[18] ),
    .A2(_0559_));
 sg13g2_nor2b_1 _2831_ (.A(net784),
    .B_N(\MemCell.prescale_reg[2][1] ),
    .Y(_0561_));
 sg13g2_nand2b_2 _2832_ (.Y(_0562_),
    .B(\MemCell.prescale_reg[2][1] ),
    .A_N(net784));
 sg13g2_a22oi_1 _2833_ (.Y(_0563_),
    .B1(_0562_),
    .B2(_2377_),
    .A2(_0559_),
    .A1(\pwm_module.prescaler1[18] ));
 sg13g2_nand2b_1 _2834_ (.Y(_0564_),
    .B(_0557_),
    .A_N(_0178_));
 sg13g2_nand2b_2 _2835_ (.Y(_0565_),
    .B(\MemCell.prescale_reg[2][0] ),
    .A_N(net783));
 sg13g2_nor2_1 _2836_ (.A(\pwm_module.prescaler1[16] ),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_nor2_1 _2837_ (.A(_2377_),
    .B(_0562_),
    .Y(_0567_));
 sg13g2_nor3_1 _2838_ (.A(_0560_),
    .B(_0566_),
    .C(_0567_),
    .Y(_0568_));
 sg13g2_o21ai_1 _2839_ (.B1(_0564_),
    .Y(_0569_),
    .A1(_0560_),
    .A2(_0563_));
 sg13g2_or4_1 _2840_ (.A(_0553_),
    .B(_0554_),
    .C(_0568_),
    .D(_0569_),
    .X(_0570_));
 sg13g2_nor2b_1 _2841_ (.A(_0544_),
    .B_N(_0545_),
    .Y(_0571_));
 sg13g2_a21oi_1 _2842_ (.A1(_0549_),
    .A2(_0552_),
    .Y(_0572_),
    .B1(_0571_));
 sg13g2_a21o_1 _2843_ (.A2(_0572_),
    .A1(_0570_),
    .B1(_0540_),
    .X(_0573_));
 sg13g2_nor3_1 _2844_ (.A(\pwm_module.prescaler1[30] ),
    .B(_0506_),
    .C(_0511_),
    .Y(_0574_));
 sg13g2_a21oi_1 _2845_ (.A1(_0185_),
    .A2(net719),
    .Y(_0575_),
    .B1(_0574_));
 sg13g2_and3_1 _2846_ (.X(_0576_),
    .A(_0536_),
    .B(_0573_),
    .C(_0575_));
 sg13g2_nor2b_1 _2847_ (.A(net780),
    .B_N(\MemCell.prescale_reg[0][6] ),
    .Y(_0577_));
 sg13g2_nand2b_2 _2848_ (.Y(_0578_),
    .B(\MemCell.prescale_reg[0][6] ),
    .A_N(net779));
 sg13g2_nor2b_2 _2849_ (.A(net780),
    .B_N(\MemCell.prescale_reg[0][7] ),
    .Y(_0579_));
 sg13g2_a22oi_1 _2850_ (.Y(_0580_),
    .B1(_0579_),
    .B2(_0171_),
    .A2(_0577_),
    .A1(_2374_));
 sg13g2_inv_1 _2851_ (.Y(_0581_),
    .A(_0580_));
 sg13g2_or2_1 _2852_ (.X(_0582_),
    .B(_0579_),
    .A(_0171_));
 sg13g2_nand2_1 _2853_ (.Y(_0583_),
    .A(\pwm_module.prescaler1[6] ),
    .B(_0578_));
 sg13g2_and3_1 _2854_ (.X(_0584_),
    .A(_0580_),
    .B(_0582_),
    .C(_0583_));
 sg13g2_nand2b_2 _2855_ (.Y(_0585_),
    .B(\MemCell.prescale_reg[0][4] ),
    .A_N(net780));
 sg13g2_or2_1 _2856_ (.X(_0586_),
    .B(_0585_),
    .A(\pwm_module.prescaler1[4] ));
 sg13g2_nor2b_2 _2857_ (.A(net780),
    .B_N(\MemCell.prescale_reg[0][5] ),
    .Y(_0587_));
 sg13g2_nand2b_1 _2858_ (.Y(_0588_),
    .B(\MemCell.prescale_reg[0][5] ),
    .A_N(net779));
 sg13g2_nor2_1 _2859_ (.A(_0170_),
    .B(_0587_),
    .Y(_0589_));
 sg13g2_nand2b_1 _2860_ (.Y(_0590_),
    .B(_0588_),
    .A_N(_0170_));
 sg13g2_nand2_1 _2861_ (.Y(_0591_),
    .A(_0170_),
    .B(_0587_));
 sg13g2_a22oi_1 _2862_ (.Y(_0592_),
    .B1(_0587_),
    .B2(_0170_),
    .A2(_0585_),
    .A1(\pwm_module.prescaler1[4] ));
 sg13g2_nand4_1 _2863_ (.B(_0586_),
    .C(_0590_),
    .A(_0584_),
    .Y(_0593_),
    .D(_0592_));
 sg13g2_nand2b_2 _2864_ (.Y(_0594_),
    .B(\MemCell.prescale_reg[0][2] ),
    .A_N(net779));
 sg13g2_nor2b_2 _2865_ (.A(net779),
    .B_N(\MemCell.prescale_reg[0][3] ),
    .Y(_0595_));
 sg13g2_nand3b_1 _2866_ (.B(\MemCell.prescale_reg[0][3] ),
    .C(_0169_),
    .Y(_0596_),
    .A_N(net779));
 sg13g2_o21ai_1 _2867_ (.B1(_0596_),
    .Y(_0597_),
    .A1(\pwm_module.prescaler1[2] ),
    .A2(_0594_));
 sg13g2_nor2_1 _2868_ (.A(_0169_),
    .B(_0595_),
    .Y(_0598_));
 sg13g2_or2_1 _2869_ (.X(_0599_),
    .B(_0595_),
    .A(_0169_));
 sg13g2_and2_1 _2870_ (.A(\pwm_module.prescaler1[2] ),
    .B(_0594_),
    .X(_0600_));
 sg13g2_nor3_1 _2871_ (.A(_0597_),
    .B(_0598_),
    .C(_0600_),
    .Y(_0601_));
 sg13g2_nor2_2 _2872_ (.A(net779),
    .B(\MemCell.prescale_reg[0][0] ),
    .Y(_0602_));
 sg13g2_nand2b_2 _2873_ (.Y(_0603_),
    .B(\MemCell.prescale_reg[0][1] ),
    .A_N(net779));
 sg13g2_a22oi_1 _2874_ (.Y(_0604_),
    .B1(_0603_),
    .B2(\pwm_module.prescaler1[1] ),
    .A2(_0602_),
    .A1(\pwm_module.prescaler1[0] ));
 sg13g2_nor2_1 _2875_ (.A(\pwm_module.prescaler1[1] ),
    .B(_0603_),
    .Y(_0605_));
 sg13g2_or2_1 _2876_ (.X(_0606_),
    .B(_0605_),
    .A(_0604_));
 sg13g2_a22oi_1 _2877_ (.Y(_0607_),
    .B1(_0601_),
    .B2(_0606_),
    .A2(_0599_),
    .A1(_0597_));
 sg13g2_o21ai_1 _2878_ (.B1(_0591_),
    .Y(_0608_),
    .A1(_0586_),
    .A2(_0589_));
 sg13g2_a22oi_1 _2879_ (.Y(_0609_),
    .B1(_0584_),
    .B2(_0608_),
    .A2(_0582_),
    .A1(_0581_));
 sg13g2_o21ai_1 _2880_ (.B1(_0609_),
    .Y(_0610_),
    .A1(_0593_),
    .A2(_0607_));
 sg13g2_nor2b_1 _2881_ (.A(net782),
    .B_N(\MemCell.prescale_reg[1][6] ),
    .Y(_0611_));
 sg13g2_nand2b_2 _2882_ (.Y(_0612_),
    .B(\MemCell.prescale_reg[1][6] ),
    .A_N(net782));
 sg13g2_nor2b_2 _2883_ (.A(net782),
    .B_N(\MemCell.prescale_reg[1][7] ),
    .Y(_0613_));
 sg13g2_a22oi_1 _2884_ (.Y(_0614_),
    .B1(_0613_),
    .B2(_0176_),
    .A2(_0611_),
    .A1(_2375_));
 sg13g2_or2_1 _2885_ (.X(_0615_),
    .B(_0613_),
    .A(_0176_));
 sg13g2_nand2_1 _2886_ (.Y(_0616_),
    .A(\pwm_module.prescaler1[14] ),
    .B(_0612_));
 sg13g2_nor2b_2 _2887_ (.A(net787),
    .B_N(\MemCell.prescale_reg[1][5] ),
    .Y(_0617_));
 sg13g2_nor2_1 _2888_ (.A(_0175_),
    .B(_0617_),
    .Y(_0618_));
 sg13g2_nand3_1 _2889_ (.B(_0615_),
    .C(_0616_),
    .A(_0614_),
    .Y(_0619_));
 sg13g2_nor2b_2 _2890_ (.A(net782),
    .B_N(\MemCell.prescale_reg[1][4] ),
    .Y(_0620_));
 sg13g2_a22oi_1 _2891_ (.Y(_0621_),
    .B1(_0620_),
    .B2(_0174_),
    .A2(_0617_),
    .A1(_0175_));
 sg13g2_or2_1 _2892_ (.X(_0622_),
    .B(_0620_),
    .A(_0174_));
 sg13g2_nand3b_1 _2893_ (.B(_0621_),
    .C(_0622_),
    .Y(_0623_),
    .A_N(_0618_));
 sg13g2_nor2_1 _2894_ (.A(_0619_),
    .B(_0623_),
    .Y(_0624_));
 sg13g2_nand2b_2 _2895_ (.Y(_0625_),
    .B(\MemCell.prescale_reg[1][1] ),
    .A_N(net781));
 sg13g2_nor2b_2 _2896_ (.A(net781),
    .B_N(\MemCell.prescale_reg[1][2] ),
    .Y(_0626_));
 sg13g2_nand2b_1 _2897_ (.Y(_0627_),
    .B(\MemCell.prescale_reg[1][2] ),
    .A_N(net781));
 sg13g2_a22oi_1 _2898_ (.Y(_0628_),
    .B1(_0627_),
    .B2(\pwm_module.prescaler1[10] ),
    .A2(_0625_),
    .A1(_2376_));
 sg13g2_nor2b_2 _2899_ (.A(net781),
    .B_N(\MemCell.prescale_reg[1][3] ),
    .Y(_0629_));
 sg13g2_nand2b_1 _2900_ (.Y(_0630_),
    .B(\MemCell.prescale_reg[1][3] ),
    .A_N(net781));
 sg13g2_nor2_1 _2901_ (.A(_0173_),
    .B(_0629_),
    .Y(_0631_));
 sg13g2_nand2b_2 _2902_ (.Y(_0632_),
    .B(\MemCell.prescale_reg[1][0] ),
    .A_N(net781));
 sg13g2_a21oi_1 _2903_ (.A1(\pwm_module.prescaler1[8] ),
    .A2(_0632_),
    .Y(_0633_),
    .B1(_0631_));
 sg13g2_nand3b_1 _2904_ (.B(\MemCell.prescale_reg[1][3] ),
    .C(_0173_),
    .Y(_0634_),
    .A_N(net781));
 sg13g2_o21ai_1 _2905_ (.B1(_0634_),
    .Y(_0635_),
    .A1(\pwm_module.prescaler1[10] ),
    .A2(_0627_));
 sg13g2_nand3b_1 _2906_ (.B(\MemCell.prescale_reg[1][1] ),
    .C(_0172_),
    .Y(_0636_),
    .A_N(net780));
 sg13g2_o21ai_1 _2907_ (.B1(_0636_),
    .Y(_0637_),
    .A1(\pwm_module.prescaler1[8] ),
    .A2(_0632_));
 sg13g2_nor2_1 _2908_ (.A(_0635_),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_and4_2 _2909_ (.A(_0624_),
    .B(_0628_),
    .C(_0633_),
    .D(_0638_),
    .X(_0639_));
 sg13g2_a21oi_1 _2910_ (.A1(_0628_),
    .A2(_0637_),
    .Y(_0640_),
    .B1(_0635_));
 sg13g2_nor4_1 _2911_ (.A(_0619_),
    .B(_0623_),
    .C(_0631_),
    .D(_0640_),
    .Y(_0641_));
 sg13g2_nor2b_1 _2912_ (.A(_0614_),
    .B_N(_0615_),
    .Y(_0642_));
 sg13g2_nor3_1 _2913_ (.A(_0618_),
    .B(_0619_),
    .C(_0621_),
    .Y(_0643_));
 sg13g2_or3_1 _2914_ (.A(_0641_),
    .B(_0642_),
    .C(_0643_),
    .X(_0644_));
 sg13g2_a21oi_2 _2915_ (.B1(_0644_),
    .Y(_0645_),
    .A2(_0639_),
    .A1(_0610_));
 sg13g2_nand2_1 _2916_ (.Y(_0646_),
    .A(\pwm_module.prescaler1[16] ),
    .B(_0565_));
 sg13g2_nand4_1 _2917_ (.B(_0564_),
    .C(_0568_),
    .A(_0563_),
    .Y(_0647_),
    .D(_0646_));
 sg13g2_nor3_1 _2918_ (.A(_0540_),
    .B(_0555_),
    .C(_0647_),
    .Y(_0648_));
 sg13g2_or3_1 _2919_ (.A(_0540_),
    .B(_0555_),
    .C(_0647_),
    .X(_0649_));
 sg13g2_o21ai_1 _2920_ (.B1(_0576_),
    .Y(_0650_),
    .A1(_0645_),
    .A2(_0649_));
 sg13g2_nor2_1 _2921_ (.A(\pwm_module.prescaler1[0] ),
    .B(_0602_),
    .Y(_0651_));
 sg13g2_nor2_1 _2922_ (.A(_0605_),
    .B(_0651_),
    .Y(_0652_));
 sg13g2_nor2b_1 _2923_ (.A(_0593_),
    .B_N(_0601_),
    .Y(_0653_));
 sg13g2_and4_2 _2924_ (.A(_0604_),
    .B(_0639_),
    .C(_0652_),
    .D(_0653_),
    .X(_0654_));
 sg13g2_a21oi_2 _2925_ (.B1(_2395_),
    .Y(_0655_),
    .A2(_0654_),
    .A1(_0648_));
 sg13g2_nand2_1 _2926_ (.Y(_0656_),
    .A(net696),
    .B(net693));
 sg13g2_and3_1 _2927_ (.X(_0657_),
    .A(net579),
    .B(\pwm_module.prescaler1[1] ),
    .C(net226));
 sg13g2_nand4_1 _2928_ (.B(\pwm_module.prescaler1[1] ),
    .C(\pwm_module.prescaler1[3] ),
    .A(\pwm_module.prescaler1[0] ),
    .Y(_0658_),
    .D(\pwm_module.prescaler1[2] ));
 sg13g2_nand2_2 _2929_ (.Y(_0659_),
    .A(\pwm_module.prescaler1[5] ),
    .B(\pwm_module.prescaler1[4] ));
 sg13g2_nor2_1 _2930_ (.A(_0658_),
    .B(_0659_),
    .Y(_0660_));
 sg13g2_nand2_1 _2931_ (.Y(_0661_),
    .A(\pwm_module.prescaler1[7] ),
    .B(net449));
 sg13g2_nor3_1 _2932_ (.A(_0658_),
    .B(_0659_),
    .C(_0661_),
    .Y(_0662_));
 sg13g2_nand2_1 _2933_ (.Y(_0663_),
    .A(\pwm_module.prescaler1[9] ),
    .B(\pwm_module.prescaler1[8] ));
 sg13g2_nor4_2 _2934_ (.A(_0658_),
    .B(_0659_),
    .C(_0661_),
    .Y(_0664_),
    .D(_0663_));
 sg13g2_and2_1 _2935_ (.A(\pwm_module.prescaler1[11] ),
    .B(\pwm_module.prescaler1[10] ),
    .X(_0665_));
 sg13g2_nand2_1 _2936_ (.Y(_0666_),
    .A(_0664_),
    .B(_0665_));
 sg13g2_and2_1 _2937_ (.A(\pwm_module.prescaler1[13] ),
    .B(\pwm_module.prescaler1[12] ),
    .X(_0667_));
 sg13g2_nor2b_1 _2938_ (.A(_0666_),
    .B_N(_0667_),
    .Y(_0668_));
 sg13g2_and2_1 _2939_ (.A(\pwm_module.prescaler1[15] ),
    .B(\pwm_module.prescaler1[14] ),
    .X(_0669_));
 sg13g2_and2_1 _2940_ (.A(_0668_),
    .B(_0669_),
    .X(_0670_));
 sg13g2_nand4_1 _2941_ (.B(_0665_),
    .C(_0667_),
    .A(_0664_),
    .Y(_0671_),
    .D(_0669_));
 sg13g2_and2_1 _2942_ (.A(net469),
    .B(_0670_),
    .X(_0672_));
 sg13g2_and3_1 _2943_ (.X(_0673_),
    .A(\pwm_module.prescaler1[17] ),
    .B(\pwm_module.prescaler1[16] ),
    .C(_0670_));
 sg13g2_nand2_1 _2944_ (.Y(_0674_),
    .A(\pwm_module.prescaler1[18] ),
    .B(_0673_));
 sg13g2_xnor2_1 _2945_ (.Y(_0675_),
    .A(net465),
    .B(_0673_));
 sg13g2_nor2_1 _2946_ (.A(net675),
    .B(net466),
    .Y(_0041_));
 sg13g2_xnor2_1 _2947_ (.Y(_0676_),
    .A(net122),
    .B(_0674_));
 sg13g2_nor2_1 _2948_ (.A(net675),
    .B(net123),
    .Y(_0042_));
 sg13g2_nand4_1 _2949_ (.B(\pwm_module.prescaler1[19] ),
    .C(\pwm_module.prescaler1[17] ),
    .A(\pwm_module.prescaler1[18] ),
    .Y(_0677_),
    .D(\pwm_module.prescaler1[16] ));
 sg13g2_nor3_1 _2950_ (.A(net407),
    .B(_0671_),
    .C(_0677_),
    .Y(_0678_));
 sg13g2_o21ai_1 _2951_ (.B1(net407),
    .Y(_0679_),
    .A1(_0671_),
    .A2(_0677_));
 sg13g2_inv_1 _2952_ (.Y(_0680_),
    .A(net408));
 sg13g2_nor3_1 _2953_ (.A(net675),
    .B(_0678_),
    .C(_0680_),
    .Y(_0044_));
 sg13g2_xnor2_1 _2954_ (.Y(_0681_),
    .A(_2313_),
    .B(_0678_));
 sg13g2_nor2_1 _2955_ (.A(net675),
    .B(net392),
    .Y(_0045_));
 sg13g2_nand2_1 _2956_ (.Y(_0682_),
    .A(\pwm_module.prescaler1[21] ),
    .B(\pwm_module.prescaler1[20] ));
 sg13g2_nor3_1 _2957_ (.A(_0671_),
    .B(_0677_),
    .C(_0682_),
    .Y(_0683_));
 sg13g2_nand2_1 _2958_ (.Y(_0684_),
    .A(\pwm_module.prescaler1[22] ),
    .B(_0683_));
 sg13g2_xnor2_1 _2959_ (.Y(_0685_),
    .A(net451),
    .B(_0683_));
 sg13g2_nor2_1 _2960_ (.A(net675),
    .B(net452),
    .Y(_0046_));
 sg13g2_xnor2_1 _2961_ (.Y(_0686_),
    .A(net192),
    .B(_0684_));
 sg13g2_nor2_1 _2962_ (.A(net675),
    .B(net193),
    .Y(_0047_));
 sg13g2_nand2_1 _2963_ (.Y(_0687_),
    .A(net451),
    .B(\pwm_module.prescaler1[23] ));
 sg13g2_nor4_2 _2964_ (.A(_0671_),
    .B(_0677_),
    .C(_0682_),
    .Y(_0688_),
    .D(_0687_));
 sg13g2_and2_1 _2965_ (.A(net453),
    .B(_0688_),
    .X(_0689_));
 sg13g2_nor2_1 _2966_ (.A(net453),
    .B(_0688_),
    .Y(_0690_));
 sg13g2_nor3_1 _2967_ (.A(net679),
    .B(_0689_),
    .C(net454),
    .Y(_0048_));
 sg13g2_xnor2_1 _2968_ (.Y(_0691_),
    .A(_2315_),
    .B(_0689_));
 sg13g2_nor2_1 _2969_ (.A(net678),
    .B(_0691_),
    .Y(_0049_));
 sg13g2_nand2_1 _2970_ (.Y(_0692_),
    .A(\pwm_module.prescaler1[25] ),
    .B(_0689_));
 sg13g2_nand3_1 _2971_ (.B(\pwm_module.prescaler1[25] ),
    .C(_0688_),
    .A(net453),
    .Y(_0693_));
 sg13g2_nand3_1 _2972_ (.B(\pwm_module.prescaler1[26] ),
    .C(_0689_),
    .A(\pwm_module.prescaler1[25] ),
    .Y(_0694_));
 sg13g2_xor2_1 _2973_ (.B(_0693_),
    .A(net529),
    .X(_0695_));
 sg13g2_nor2_1 _2974_ (.A(net678),
    .B(net530),
    .Y(_0050_));
 sg13g2_xnor2_1 _2975_ (.Y(_0696_),
    .A(net388),
    .B(_0694_));
 sg13g2_nor2_1 _2976_ (.A(net678),
    .B(net389),
    .Y(_0051_));
 sg13g2_nand2_1 _2977_ (.Y(_0697_),
    .A(\pwm_module.prescaler1[26] ),
    .B(\pwm_module.prescaler1[27] ));
 sg13g2_nor2_1 _2978_ (.A(_0693_),
    .B(_0697_),
    .Y(_0698_));
 sg13g2_nor2_1 _2979_ (.A(net442),
    .B(_0698_),
    .Y(_0699_));
 sg13g2_nor3_2 _2980_ (.A(_2316_),
    .B(_0692_),
    .C(_0697_),
    .Y(_0700_));
 sg13g2_nor3_1 _2981_ (.A(net678),
    .B(net443),
    .C(_0700_),
    .Y(_0052_));
 sg13g2_nor2b_1 _2982_ (.A(_0700_),
    .B_N(net100),
    .Y(_0701_));
 sg13g2_nor2b_1 _2983_ (.A(net100),
    .B_N(_0700_),
    .Y(_0702_));
 sg13g2_nor3_1 _2984_ (.A(net678),
    .B(_0701_),
    .C(_0702_),
    .Y(_0053_));
 sg13g2_a21oi_1 _2985_ (.A1(net80),
    .A2(_0700_),
    .Y(_0703_),
    .B1(\pwm_module.prescaler1[30] ));
 sg13g2_nand3_1 _2986_ (.B(\pwm_module.prescaler1[30] ),
    .C(_0700_),
    .A(net80),
    .Y(_0704_));
 sg13g2_inv_1 _2987_ (.Y(_0705_),
    .A(_0704_));
 sg13g2_nor3_1 _2988_ (.A(net678),
    .B(net81),
    .C(_0705_),
    .Y(_0055_));
 sg13g2_a21oi_1 _2989_ (.A1(net393),
    .A2(_0704_),
    .Y(_0706_),
    .B1(net678));
 sg13g2_nor2_1 _2990_ (.A(net393),
    .B(_0704_),
    .Y(_0707_));
 sg13g2_nor2b_1 _2991_ (.A(net394),
    .B_N(_0706_),
    .Y(_0056_));
 sg13g2_nand3b_1 _2992_ (.B(\MemCell.prescale_reg[1][7] ),
    .C(_0193_),
    .Y(_0708_),
    .A_N(net782));
 sg13g2_o21ai_1 _2993_ (.B1(_0708_),
    .Y(_0709_),
    .A1(\pwm_module.prescaler2[14] ),
    .A2(_0612_));
 sg13g2_nand2_1 _2994_ (.Y(_0710_),
    .A(\pwm_module.prescaler2[14] ),
    .B(_0612_));
 sg13g2_or2_1 _2995_ (.X(_0711_),
    .B(_0613_),
    .A(_0193_));
 sg13g2_nand3b_1 _2996_ (.B(_0710_),
    .C(_0711_),
    .Y(_0712_),
    .A_N(_0709_));
 sg13g2_nand3b_1 _2997_ (.B(\MemCell.prescale_reg[1][5] ),
    .C(_0192_),
    .Y(_0713_),
    .A_N(net782));
 sg13g2_nand3b_1 _2998_ (.B(\MemCell.prescale_reg[1][4] ),
    .C(_0191_),
    .Y(_0714_),
    .A_N(net782));
 sg13g2_nand2_1 _2999_ (.Y(_0715_),
    .A(_0713_),
    .B(_0714_));
 sg13g2_nor2_1 _3000_ (.A(_0192_),
    .B(_0617_),
    .Y(_0716_));
 sg13g2_or2_1 _3001_ (.X(_0717_),
    .B(_0617_),
    .A(_0192_));
 sg13g2_or2_1 _3002_ (.X(_0718_),
    .B(_0620_),
    .A(_0191_));
 sg13g2_o21ai_1 _3003_ (.B1(_0718_),
    .Y(_0719_),
    .A1(_0190_),
    .A2(_0629_));
 sg13g2_nor4_1 _3004_ (.A(_0712_),
    .B(_0715_),
    .C(_0716_),
    .D(_0719_),
    .Y(_0720_));
 sg13g2_nor2_1 _3005_ (.A(_2334_),
    .B(_0626_),
    .Y(_0721_));
 sg13g2_nor2_1 _3006_ (.A(\pwm_module.prescaler2[8] ),
    .B(_0632_),
    .Y(_0722_));
 sg13g2_nand2_1 _3007_ (.Y(_0723_),
    .A(_2333_),
    .B(_0625_));
 sg13g2_a22oi_1 _3008_ (.Y(_0724_),
    .B1(_0629_),
    .B2(_0190_),
    .A2(_0626_),
    .A1(_2334_));
 sg13g2_nor2_1 _3009_ (.A(_2333_),
    .B(_0625_),
    .Y(_0725_));
 sg13g2_xor2_1 _3010_ (.B(_0632_),
    .A(\pwm_module.prescaler2[8] ),
    .X(_0726_));
 sg13g2_nand4_1 _3011_ (.B(_0714_),
    .C(_0717_),
    .A(_0713_),
    .Y(_0727_),
    .D(_0718_));
 sg13g2_a22oi_1 _3012_ (.Y(_0728_),
    .B1(_0630_),
    .B2(_2335_),
    .A2(_0627_),
    .A1(\pwm_module.prescaler2[10] ));
 sg13g2_xnor2_1 _3013_ (.Y(_0729_),
    .A(_0189_),
    .B(_0625_));
 sg13g2_nand4_1 _3014_ (.B(_0726_),
    .C(_0728_),
    .A(_0724_),
    .Y(_0730_),
    .D(_0729_));
 sg13g2_nor3_2 _3015_ (.A(_0712_),
    .B(_0727_),
    .C(_0730_),
    .Y(_0731_));
 sg13g2_nand2_1 _3016_ (.Y(_0732_),
    .A(_0187_),
    .B(_0587_));
 sg13g2_o21ai_1 _3017_ (.B1(_0732_),
    .Y(_0733_),
    .A1(\pwm_module.prescaler2[4] ),
    .A2(_0585_));
 sg13g2_nor2_1 _3018_ (.A(_0188_),
    .B(_0579_),
    .Y(_0734_));
 sg13g2_nand3b_1 _3019_ (.B(\MemCell.prescale_reg[0][7] ),
    .C(_0188_),
    .Y(_0735_),
    .A_N(net780));
 sg13g2_o21ai_1 _3020_ (.B1(_0735_),
    .Y(_0736_),
    .A1(\pwm_module.prescaler2[6] ),
    .A2(_0578_));
 sg13g2_and2_1 _3021_ (.A(\pwm_module.prescaler2[6] ),
    .B(_0578_),
    .X(_0737_));
 sg13g2_nor2_1 _3022_ (.A(_0187_),
    .B(_0587_),
    .Y(_0738_));
 sg13g2_nor4_2 _3023_ (.A(_0734_),
    .B(_0736_),
    .C(_0737_),
    .Y(_0739_),
    .D(_0738_));
 sg13g2_a21oi_1 _3024_ (.A1(\pwm_module.prescaler2[4] ),
    .A2(_0585_),
    .Y(_0740_),
    .B1(_0733_));
 sg13g2_nand3_1 _3025_ (.B(_0739_),
    .C(_0740_),
    .A(_0731_),
    .Y(_0741_));
 sg13g2_nand3b_1 _3026_ (.B(\MemCell.prescale_reg[0][3] ),
    .C(_0186_),
    .Y(_0742_),
    .A_N(net779));
 sg13g2_o21ai_1 _3027_ (.B1(_0742_),
    .Y(_0743_),
    .A1(\pwm_module.prescaler2[2] ),
    .A2(_0594_));
 sg13g2_or2_1 _3028_ (.X(_0744_),
    .B(_0595_),
    .A(_0186_));
 sg13g2_nand2_1 _3029_ (.Y(_0745_),
    .A(\pwm_module.prescaler2[2] ),
    .B(_0594_));
 sg13g2_nand3b_1 _3030_ (.B(_0744_),
    .C(_0745_),
    .Y(_0746_),
    .A_N(_0743_));
 sg13g2_nor2_1 _3031_ (.A(\pwm_module.prescaler2[1] ),
    .B(_0603_),
    .Y(_0747_));
 sg13g2_nand2_1 _3032_ (.Y(_0748_),
    .A(\pwm_module.prescaler2[0] ),
    .B(_0602_));
 sg13g2_xor2_1 _3033_ (.B(_0603_),
    .A(\pwm_module.prescaler2[1] ),
    .X(_0749_));
 sg13g2_nand2_1 _3034_ (.Y(_0750_),
    .A(_0748_),
    .B(_0749_));
 sg13g2_a21oi_1 _3035_ (.A1(_0748_),
    .A2(_0749_),
    .Y(_0751_),
    .B1(_0747_));
 sg13g2_nand2_1 _3036_ (.Y(_0752_),
    .A(_0743_),
    .B(_0744_));
 sg13g2_o21ai_1 _3037_ (.B1(_0752_),
    .Y(_0753_),
    .A1(_0746_),
    .A2(_0751_));
 sg13g2_nand4_1 _3038_ (.B(_0739_),
    .C(_0740_),
    .A(_0731_),
    .Y(_0754_),
    .D(_0753_));
 sg13g2_nor2b_1 _3039_ (.A(_0734_),
    .B_N(_0736_),
    .Y(_0755_));
 sg13g2_a21o_1 _3040_ (.A2(_0739_),
    .A1(_0733_),
    .B1(_0755_),
    .X(_0756_));
 sg13g2_nand2_1 _3041_ (.Y(_0757_),
    .A(_0709_),
    .B(_0711_));
 sg13g2_nand2_1 _3042_ (.Y(_0758_),
    .A(_0715_),
    .B(_0717_));
 sg13g2_o21ai_1 _3043_ (.B1(_0757_),
    .Y(_0759_),
    .A1(_0712_),
    .A2(_0758_));
 sg13g2_a21oi_1 _3044_ (.A1(_0722_),
    .A2(_0723_),
    .Y(_0760_),
    .B1(_0725_));
 sg13g2_o21ai_1 _3045_ (.B1(_0724_),
    .Y(_0761_),
    .A1(_0721_),
    .A2(_0760_));
 sg13g2_a221oi_1 _3046_ (.B2(_0720_),
    .C1(_0759_),
    .B1(_0761_),
    .A1(_0731_),
    .Y(_0762_),
    .A2(_0756_));
 sg13g2_or2_1 _3047_ (.X(_0763_),
    .B(net719),
    .A(_0123_));
 sg13g2_nor2_1 _3048_ (.A(\pwm_module.prescaler2[30] ),
    .B(_0506_),
    .Y(_0764_));
 sg13g2_nand2_1 _3049_ (.Y(_0765_),
    .A(_0123_),
    .B(net719));
 sg13g2_or2_1 _3050_ (.X(_0766_),
    .B(_0508_),
    .A(_0201_));
 sg13g2_xor2_1 _3051_ (.B(_0506_),
    .A(\pwm_module.prescaler2[30] ),
    .X(_0767_));
 sg13g2_nand4_1 _3052_ (.B(_0765_),
    .C(_0766_),
    .A(_0763_),
    .Y(_0768_),
    .D(_0767_));
 sg13g2_a22oi_1 _3053_ (.Y(_0769_),
    .B1(_0513_),
    .B2(_2343_),
    .A2(_0508_),
    .A1(_0201_));
 sg13g2_o21ai_1 _3054_ (.B1(_0769_),
    .Y(_0770_),
    .A1(_2343_),
    .A2(_0513_));
 sg13g2_nor2_1 _3055_ (.A(_0768_),
    .B(_0770_),
    .Y(_0771_));
 sg13g2_a22oi_1 _3056_ (.Y(_0772_),
    .B1(_0524_),
    .B2(\pwm_module.prescaler2[26] ),
    .A2(_0520_),
    .A1(_2340_));
 sg13g2_a22oi_1 _3057_ (.Y(_0773_),
    .B1(_0528_),
    .B2(_2342_),
    .A2(_0518_),
    .A1(\pwm_module.prescaler2[24] ));
 sg13g2_a22oi_1 _3058_ (.Y(_0774_),
    .B1(_0527_),
    .B2(_0200_),
    .A2(_0523_),
    .A1(_2341_));
 sg13g2_a22oi_1 _3059_ (.Y(_0775_),
    .B1(_0519_),
    .B2(_0199_),
    .A2(_0517_),
    .A1(_2339_));
 sg13g2_nand4_1 _3060_ (.B(_0773_),
    .C(_0774_),
    .A(_0772_),
    .Y(_0776_),
    .D(_0775_));
 sg13g2_nor3_2 _3061_ (.A(_0768_),
    .B(_0770_),
    .C(_0776_),
    .Y(_0777_));
 sg13g2_a22oi_1 _3062_ (.Y(_0778_),
    .B1(_0543_),
    .B2(_0198_),
    .A2(_0541_),
    .A1(_2338_));
 sg13g2_or2_1 _3063_ (.X(_0779_),
    .B(_0543_),
    .A(_0198_));
 sg13g2_a22oi_1 _3064_ (.Y(_0780_),
    .B1(_0547_),
    .B2(_2337_),
    .A2(_0542_),
    .A1(\pwm_module.prescaler2[22] ));
 sg13g2_and3_1 _3065_ (.X(_0781_),
    .A(_0778_),
    .B(_0779_),
    .C(_0780_));
 sg13g2_nand3b_1 _3066_ (.B(\MemCell.prescale_reg[2][4] ),
    .C(_0196_),
    .Y(_0782_),
    .A_N(net783));
 sg13g2_o21ai_1 _3067_ (.B1(_0782_),
    .Y(_0783_),
    .A1(_2337_),
    .A2(_0547_));
 sg13g2_nor2_1 _3068_ (.A(_0196_),
    .B(_0550_),
    .Y(_0784_));
 sg13g2_nor2_1 _3069_ (.A(_0783_),
    .B(_0784_),
    .Y(_0785_));
 sg13g2_nand2_1 _3070_ (.Y(_0786_),
    .A(_0781_),
    .B(_0785_));
 sg13g2_nand2_1 _3071_ (.Y(_0787_),
    .A(_0195_),
    .B(_0556_));
 sg13g2_xnor2_1 _3072_ (.Y(_0788_),
    .A(_0195_),
    .B(_0557_));
 sg13g2_nor2_1 _3073_ (.A(\pwm_module.prescaler2[18] ),
    .B(_0559_),
    .Y(_0789_));
 sg13g2_xor2_1 _3074_ (.B(_0559_),
    .A(\pwm_module.prescaler2[18] ),
    .X(_0790_));
 sg13g2_and2_1 _3075_ (.A(_0788_),
    .B(_0790_),
    .X(_0791_));
 sg13g2_nand3b_1 _3076_ (.B(\MemCell.prescale_reg[2][1] ),
    .C(_0194_),
    .Y(_0792_),
    .A_N(net784));
 sg13g2_o21ai_1 _3077_ (.B1(_0792_),
    .Y(_0793_),
    .A1(\pwm_module.prescaler2[16] ),
    .A2(_0565_));
 sg13g2_nand2_1 _3078_ (.Y(_0794_),
    .A(_2336_),
    .B(_0562_));
 sg13g2_a22oi_1 _3079_ (.Y(_0795_),
    .B1(_0565_),
    .B2(\pwm_module.prescaler2[16] ),
    .A2(_0562_),
    .A1(_2336_));
 sg13g2_nor2b_1 _3080_ (.A(_0793_),
    .B_N(_0795_),
    .Y(_0796_));
 sg13g2_and4_2 _3081_ (.A(_0781_),
    .B(_0785_),
    .C(_0791_),
    .D(_0796_),
    .X(_0797_));
 sg13g2_nand2_1 _3082_ (.Y(_0798_),
    .A(_0777_),
    .B(_0797_));
 sg13g2_a21o_1 _3083_ (.A2(_0762_),
    .A1(_0754_),
    .B1(_0798_),
    .X(_0799_));
 sg13g2_nand4_1 _3084_ (.B(_0790_),
    .C(_0793_),
    .A(_0788_),
    .Y(_0800_),
    .D(_0794_));
 sg13g2_o21ai_1 _3085_ (.B1(_0789_),
    .Y(_0801_),
    .A1(_0195_),
    .A2(_0556_));
 sg13g2_and3_1 _3086_ (.X(_0802_),
    .A(_0787_),
    .B(_0800_),
    .C(_0801_));
 sg13g2_nor2b_1 _3087_ (.A(_0778_),
    .B_N(_0779_),
    .Y(_0803_));
 sg13g2_a21oi_1 _3088_ (.A1(_0781_),
    .A2(_0783_),
    .Y(_0804_),
    .B1(_0803_));
 sg13g2_o21ai_1 _3089_ (.B1(_0804_),
    .Y(_0805_),
    .A1(_0786_),
    .A2(_0802_));
 sg13g2_nand2b_1 _3090_ (.Y(_0806_),
    .B(_0772_),
    .A_N(_0775_));
 sg13g2_a22oi_1 _3091_ (.Y(_0807_),
    .B1(_0774_),
    .B2(_0806_),
    .A2(_0528_),
    .A1(_2342_));
 sg13g2_or2_1 _3092_ (.X(_0808_),
    .B(_0769_),
    .A(_0768_));
 sg13g2_o21ai_1 _3093_ (.B1(_0764_),
    .Y(_0809_),
    .A1(_0123_),
    .A2(net719));
 sg13g2_nand3_1 _3094_ (.B(_0808_),
    .C(_0809_),
    .A(_0765_),
    .Y(_0810_));
 sg13g2_a221oi_1 _3095_ (.B2(_0771_),
    .C1(_0810_),
    .B1(_0807_),
    .A1(_0777_),
    .Y(_0811_),
    .A2(_0805_));
 sg13g2_nor2_1 _3096_ (.A(\pwm_module.prescaler2[0] ),
    .B(_0602_),
    .Y(_0812_));
 sg13g2_nor3_2 _3097_ (.A(_0746_),
    .B(_0750_),
    .C(_0812_),
    .Y(_0813_));
 sg13g2_nand3_1 _3098_ (.B(_0797_),
    .C(_0813_),
    .A(_0777_),
    .Y(_0814_));
 sg13g2_o21ai_1 _3099_ (.B1(_2396_),
    .Y(_0815_),
    .A1(_0741_),
    .A2(_0814_));
 sg13g2_a21oi_1 _3100_ (.A1(_0799_),
    .A2(_0811_),
    .Y(_0816_),
    .B1(_0815_));
 sg13g2_nor2b_1 _3101_ (.A(net283),
    .B_N(net682),
    .Y(_0064_));
 sg13g2_xor2_1 _3102_ (.B(net561),
    .A(net283),
    .X(_0817_));
 sg13g2_and2_1 _3103_ (.A(net682),
    .B(_0817_),
    .X(_0075_));
 sg13g2_and3_1 _3104_ (.X(_0818_),
    .A(\pwm_module.prescaler2[0] ),
    .B(\pwm_module.prescaler2[1] ),
    .C(\pwm_module.prescaler2[2] ));
 sg13g2_a21oi_1 _3105_ (.A1(net283),
    .A2(\pwm_module.prescaler2[1] ),
    .Y(_0819_),
    .B1(net547));
 sg13g2_nor2_1 _3106_ (.A(_0818_),
    .B(net548),
    .Y(_0820_));
 sg13g2_and2_1 _3107_ (.A(net682),
    .B(_0820_),
    .X(_0086_));
 sg13g2_xnor2_1 _3108_ (.Y(_0821_),
    .A(net427),
    .B(_0818_));
 sg13g2_and2_1 _3109_ (.A(net682),
    .B(net428),
    .X(_0089_));
 sg13g2_and4_2 _3110_ (.A(\pwm_module.prescaler2[0] ),
    .B(\pwm_module.prescaler2[1] ),
    .C(\pwm_module.prescaler2[2] ),
    .D(\pwm_module.prescaler2[3] ),
    .X(_0822_));
 sg13g2_nor2_1 _3111_ (.A(net412),
    .B(_0822_),
    .Y(_0823_));
 sg13g2_and2_1 _3112_ (.A(\pwm_module.prescaler2[4] ),
    .B(_0822_),
    .X(_0824_));
 sg13g2_nand2b_1 _3113_ (.Y(_0825_),
    .B(net682),
    .A_N(_0824_));
 sg13g2_nor2_1 _3114_ (.A(net413),
    .B(_0825_),
    .Y(_0090_));
 sg13g2_xnor2_1 _3115_ (.Y(_0826_),
    .A(net402),
    .B(_0824_));
 sg13g2_and2_1 _3116_ (.A(net682),
    .B(_0826_),
    .X(_0091_));
 sg13g2_a21oi_1 _3117_ (.A1(\pwm_module.prescaler2[5] ),
    .A2(_0824_),
    .Y(_0827_),
    .B1(net242));
 sg13g2_and3_1 _3118_ (.X(_0828_),
    .A(\pwm_module.prescaler2[5] ),
    .B(\pwm_module.prescaler2[6] ),
    .C(_0824_));
 sg13g2_nand2b_1 _3119_ (.Y(_0829_),
    .B(net682),
    .A_N(_0828_));
 sg13g2_nor2_1 _3120_ (.A(net243),
    .B(_0829_),
    .Y(_0092_));
 sg13g2_xnor2_1 _3121_ (.Y(_0830_),
    .A(net404),
    .B(_0828_));
 sg13g2_and2_1 _3122_ (.A(net682),
    .B(_0830_),
    .X(_0093_));
 sg13g2_and2_1 _3123_ (.A(\pwm_module.prescaler2[6] ),
    .B(\pwm_module.prescaler2[7] ),
    .X(_0831_));
 sg13g2_nand4_1 _3124_ (.B(\pwm_module.prescaler2[5] ),
    .C(_0822_),
    .A(\pwm_module.prescaler2[4] ),
    .Y(_0832_),
    .D(_0831_));
 sg13g2_nand3_1 _3125_ (.B(\pwm_module.prescaler2[8] ),
    .C(_0828_),
    .A(\pwm_module.prescaler2[7] ),
    .Y(_0833_));
 sg13g2_xnor2_1 _3126_ (.Y(_0834_),
    .A(net569),
    .B(_0832_));
 sg13g2_and2_1 _3127_ (.A(net683),
    .B(_0834_),
    .X(_0094_));
 sg13g2_xor2_1 _3128_ (.B(_0833_),
    .A(net431),
    .X(_0835_));
 sg13g2_and2_1 _3129_ (.A(net683),
    .B(net432),
    .X(_0095_));
 sg13g2_nand2_2 _3130_ (.Y(_0836_),
    .A(\pwm_module.prescaler2[8] ),
    .B(net543));
 sg13g2_nor3_2 _3131_ (.A(_2334_),
    .B(_0832_),
    .C(_0836_),
    .Y(_0837_));
 sg13g2_o21ai_1 _3132_ (.B1(_2334_),
    .Y(_0838_),
    .A1(_0832_),
    .A2(_0836_));
 sg13g2_nand2_1 _3133_ (.Y(_0839_),
    .A(net683),
    .B(net544));
 sg13g2_nor2_1 _3134_ (.A(_0837_),
    .B(_0839_),
    .Y(_0065_));
 sg13g2_xnor2_1 _3135_ (.Y(_0840_),
    .A(net492),
    .B(_0837_));
 sg13g2_and2_1 _3136_ (.A(net683),
    .B(net493),
    .X(_0066_));
 sg13g2_nand2_1 _3137_ (.Y(_0841_),
    .A(\pwm_module.prescaler2[11] ),
    .B(_0837_));
 sg13g2_nand2_1 _3138_ (.Y(_0842_),
    .A(\pwm_module.prescaler2[10] ),
    .B(\pwm_module.prescaler2[11] ));
 sg13g2_nor2_1 _3139_ (.A(net36),
    .B(_0841_),
    .Y(_0843_));
 sg13g2_nand2b_1 _3140_ (.Y(_0844_),
    .B(net683),
    .A_N(_0843_));
 sg13g2_a21oi_1 _3141_ (.A1(net36),
    .A2(_0841_),
    .Y(_0067_),
    .B1(_0844_));
 sg13g2_xnor2_1 _3142_ (.Y(_0845_),
    .A(net474),
    .B(_0843_));
 sg13g2_and2_1 _3143_ (.A(net683),
    .B(net475),
    .X(_0068_));
 sg13g2_nand2_1 _3144_ (.Y(_0846_),
    .A(\pwm_module.prescaler2[13] ),
    .B(\pwm_module.prescaler2[12] ));
 sg13g2_nor2_1 _3145_ (.A(_0841_),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_nor4_2 _3146_ (.A(_0832_),
    .B(_0836_),
    .C(_0842_),
    .Y(_0848_),
    .D(_0846_));
 sg13g2_or2_1 _3147_ (.X(_0849_),
    .B(_0848_),
    .A(net567));
 sg13g2_nand2_1 _3148_ (.Y(_0850_),
    .A(net567),
    .B(_0847_));
 sg13g2_and3_1 _3149_ (.X(_0069_),
    .A(net683),
    .B(net568),
    .C(_0850_));
 sg13g2_o21ai_1 _3150_ (.B1(net683),
    .Y(_0851_),
    .A1(net40),
    .A2(_0850_));
 sg13g2_a21oi_1 _3151_ (.A1(net40),
    .A2(_0850_),
    .Y(_0070_),
    .B1(_0851_));
 sg13g2_nand4_1 _3152_ (.B(net540),
    .C(\pwm_module.prescaler2[16] ),
    .A(net578),
    .Y(_0852_),
    .D(_0847_));
 sg13g2_nand3_1 _3153_ (.B(net540),
    .C(_0848_),
    .A(\pwm_module.prescaler2[14] ),
    .Y(_0853_));
 sg13g2_nand2b_1 _3154_ (.Y(_0854_),
    .B(net541),
    .A_N(\pwm_module.prescaler2[16] ));
 sg13g2_and3_1 _3155_ (.X(_0071_),
    .A(net690),
    .B(_0852_),
    .C(net542));
 sg13g2_o21ai_1 _3156_ (.B1(net690),
    .Y(_0855_),
    .A1(net42),
    .A2(_0852_));
 sg13g2_a21oi_1 _3157_ (.A1(net42),
    .A2(_0852_),
    .Y(_0072_),
    .B1(_0855_));
 sg13g2_nand2_1 _3158_ (.Y(_0856_),
    .A(\pwm_module.prescaler2[16] ),
    .B(\pwm_module.prescaler2[17] ));
 sg13g2_nor2_1 _3159_ (.A(_0853_),
    .B(_0856_),
    .Y(_0857_));
 sg13g2_or2_1 _3160_ (.X(_0858_),
    .B(_0857_),
    .A(net570));
 sg13g2_nand2_1 _3161_ (.Y(_0859_),
    .A(net570),
    .B(_0857_));
 sg13g2_and3_1 _3162_ (.X(_0073_),
    .A(net690),
    .B(net571),
    .C(_0859_));
 sg13g2_xor2_1 _3163_ (.B(_0859_),
    .A(net513),
    .X(_0860_));
 sg13g2_and2_1 _3164_ (.A(net690),
    .B(net514),
    .X(_0074_));
 sg13g2_and4_1 _3165_ (.A(\pwm_module.prescaler2[16] ),
    .B(\pwm_module.prescaler2[17] ),
    .C(\pwm_module.prescaler2[18] ),
    .D(\pwm_module.prescaler2[19] ),
    .X(_0861_));
 sg13g2_nand4_1 _3166_ (.B(\pwm_module.prescaler2[15] ),
    .C(_0848_),
    .A(\pwm_module.prescaler2[14] ),
    .Y(_0862_),
    .D(_0861_));
 sg13g2_nor2_1 _3167_ (.A(_0196_),
    .B(_0862_),
    .Y(_0863_));
 sg13g2_xor2_1 _3168_ (.B(_0862_),
    .A(net497),
    .X(_0864_));
 sg13g2_and2_1 _3169_ (.A(net690),
    .B(net498),
    .X(_0076_));
 sg13g2_xnor2_1 _3170_ (.Y(_0865_),
    .A(net384),
    .B(_0863_));
 sg13g2_and2_1 _3171_ (.A(net690),
    .B(net385),
    .X(_0077_));
 sg13g2_nand2_1 _3172_ (.Y(_0866_),
    .A(net508),
    .B(\pwm_module.prescaler2[20] ));
 sg13g2_nor2_1 _3173_ (.A(_0862_),
    .B(_0866_),
    .Y(_0867_));
 sg13g2_o21ai_1 _3174_ (.B1(_2338_),
    .Y(_0868_),
    .A1(_0862_),
    .A2(net509));
 sg13g2_nand2_1 _3175_ (.Y(_0869_),
    .A(\pwm_module.prescaler2[22] ),
    .B(_0867_));
 sg13g2_and3_1 _3176_ (.X(_0078_),
    .A(net690),
    .B(net510),
    .C(_0869_));
 sg13g2_o21ai_1 _3177_ (.B1(net689),
    .Y(_0870_),
    .A1(net54),
    .A2(_0869_));
 sg13g2_a21oi_1 _3178_ (.A1(net54),
    .A2(_0869_),
    .Y(_0079_),
    .B1(_0870_));
 sg13g2_nand3_1 _3179_ (.B(\pwm_module.prescaler2[23] ),
    .C(_0867_),
    .A(\pwm_module.prescaler2[22] ),
    .Y(_0871_));
 sg13g2_or2_1 _3180_ (.X(_0872_),
    .B(_0871_),
    .A(_2339_));
 sg13g2_nand2_1 _3181_ (.Y(_0873_),
    .A(net689),
    .B(_0872_));
 sg13g2_a21oi_1 _3182_ (.A1(_2339_),
    .A2(_0871_),
    .Y(_0080_),
    .B1(_0873_));
 sg13g2_xnor2_1 _3183_ (.Y(_0874_),
    .A(_2340_),
    .B(_0872_));
 sg13g2_and2_1 _3184_ (.A(net689),
    .B(_0874_),
    .X(_0081_));
 sg13g2_nand2_1 _3185_ (.Y(_0875_),
    .A(\pwm_module.prescaler2[24] ),
    .B(\pwm_module.prescaler2[25] ));
 sg13g2_nor2_1 _3186_ (.A(_0871_),
    .B(_0875_),
    .Y(_0876_));
 sg13g2_nor3_1 _3187_ (.A(_2341_),
    .B(_0871_),
    .C(_0875_),
    .Y(_0877_));
 sg13g2_xnor2_1 _3188_ (.Y(_0878_),
    .A(_2341_),
    .B(_0876_));
 sg13g2_and2_1 _3189_ (.A(net689),
    .B(_0878_),
    .X(_0082_));
 sg13g2_o21ai_1 _3190_ (.B1(net689),
    .Y(_0879_),
    .A1(_2342_),
    .A2(_0877_));
 sg13g2_a21oi_1 _3191_ (.A1(_2342_),
    .A2(_0877_),
    .Y(_0083_),
    .B1(_0879_));
 sg13g2_nand2_1 _3192_ (.Y(_0880_),
    .A(\pwm_module.prescaler2[26] ),
    .B(\pwm_module.prescaler2[27] ));
 sg13g2_nor3_2 _3193_ (.A(_0871_),
    .B(_0875_),
    .C(_0880_),
    .Y(_0881_));
 sg13g2_nand2_1 _3194_ (.Y(_0882_),
    .A(\pwm_module.prescaler2[28] ),
    .B(_0881_));
 sg13g2_xnor2_1 _3195_ (.Y(_0883_),
    .A(_2343_),
    .B(_0881_));
 sg13g2_and2_1 _3196_ (.A(net690),
    .B(net576),
    .X(_0084_));
 sg13g2_o21ai_1 _3197_ (.B1(net689),
    .Y(_0884_),
    .A1(net56),
    .A2(_0882_));
 sg13g2_a21oi_1 _3198_ (.A1(net56),
    .A2(_0882_),
    .Y(_0085_),
    .B1(_0884_));
 sg13g2_nand3_1 _3199_ (.B(net515),
    .C(_0881_),
    .A(\pwm_module.prescaler2[28] ),
    .Y(_0885_));
 sg13g2_nand2b_1 _3200_ (.Y(_0886_),
    .B(net516),
    .A_N(\pwm_module.prescaler2[30] ));
 sg13g2_nand4_1 _3201_ (.B(net515),
    .C(\pwm_module.prescaler2[30] ),
    .A(\pwm_module.prescaler2[28] ),
    .Y(_0887_),
    .D(_0881_));
 sg13g2_and3_1 _3202_ (.X(_0087_),
    .A(net689),
    .B(net517),
    .C(_0887_));
 sg13g2_xor2_1 _3203_ (.B(_0887_),
    .A(net503),
    .X(_0888_));
 sg13g2_and2_1 _3204_ (.A(net689),
    .B(net504),
    .X(_0088_));
 sg13g2_nand2_1 _3205_ (.Y(_0889_),
    .A(net415),
    .B(net559));
 sg13g2_xor2_1 _3206_ (.B(_0889_),
    .A(net753),
    .X(_0890_));
 sg13g2_nand2_1 _3207_ (.Y(_0891_),
    .A(\MemCell.curr_state[0] ),
    .B(_0144_));
 sg13g2_nand2_1 _3208_ (.Y(_0892_),
    .A(\MemCell.curr_state[0] ),
    .B(\MemCell.curr_state[1] ));
 sg13g2_nor2_2 _3209_ (.A(\MemCell.curr_state[2] ),
    .B(_0892_),
    .Y(_0893_));
 sg13g2_nor2b_1 _3210_ (.A(\MemCell.curr_state[1] ),
    .B_N(\MemCell.curr_state[2] ),
    .Y(_0894_));
 sg13g2_and2_1 _3211_ (.A(\MemCell.curr_state[0] ),
    .B(_0894_),
    .X(_0895_));
 sg13g2_nor2_1 _3212_ (.A(_0893_),
    .B(_0895_),
    .Y(_0896_));
 sg13g2_o21ai_1 _3213_ (.B1(_0896_),
    .Y(_0897_),
    .A1(\MemCell.curr_state[1] ),
    .A2(_0891_));
 sg13g2_nor2_1 _3214_ (.A(\MemCell.curr_state[0] ),
    .B(\MemCell.curr_state[1] ),
    .Y(_0898_));
 sg13g2_nor3_2 _3215_ (.A(\MemCell.curr_state[0] ),
    .B(\MemCell.curr_state[1] ),
    .C(net558),
    .Y(_0899_));
 sg13g2_nor2b_1 _3216_ (.A(\MemCell.curr_state[0] ),
    .B_N(\MemCell.curr_state[1] ),
    .Y(_0900_));
 sg13g2_nand2_1 _3217_ (.Y(_0901_),
    .A(net420),
    .B(_0900_));
 sg13g2_nand2_1 _3218_ (.Y(_0902_),
    .A(_0144_),
    .B(_0900_));
 sg13g2_nor2_1 _3219_ (.A(_0144_),
    .B(_0892_),
    .Y(_0903_));
 sg13g2_nor3_1 _3220_ (.A(_0897_),
    .B(_0899_),
    .C(_0903_),
    .Y(_0904_));
 sg13g2_and3_1 _3221_ (.X(_0905_),
    .A(_0901_),
    .B(_0902_),
    .C(_0904_));
 sg13g2_nor2_1 _3222_ (.A(net749),
    .B(net740),
    .Y(_0906_));
 sg13g2_nor4_1 _3223_ (.A(net744),
    .B(net732),
    .C(net736),
    .D(_2346_),
    .Y(_0907_));
 sg13g2_nand3_1 _3224_ (.B(_0906_),
    .C(_0907_),
    .A(_0905_),
    .Y(_0908_));
 sg13g2_and2_1 _3225_ (.A(net729),
    .B(\MemCell.counter[1] ),
    .X(_0909_));
 sg13g2_nand2_2 _3226_ (.Y(_0910_),
    .A(net729),
    .B(\MemCell.counter[1] ));
 sg13g2_a21oi_2 _3227_ (.B1(_0905_),
    .Y(_0911_),
    .A2(_0909_),
    .A1(\MemCell.o_RX_DV ));
 sg13g2_nand2_1 _3228_ (.Y(_0912_),
    .A(_0897_),
    .B(_0911_));
 sg13g2_o21ai_1 _3229_ (.B1(_0912_),
    .Y(\MemCell.next_state[0] ),
    .A1(_0890_),
    .A2(_0908_));
 sg13g2_nor2b_1 _3230_ (.A(_0893_),
    .B_N(_0902_),
    .Y(_0913_));
 sg13g2_nand2b_1 _3231_ (.Y(_0914_),
    .B(_0911_),
    .A_N(_0913_));
 sg13g2_o21ai_1 _3232_ (.B1(_0914_),
    .Y(\MemCell.next_state[1] ),
    .A1(net726),
    .A2(_0908_));
 sg13g2_o21ai_1 _3233_ (.B1(_0911_),
    .Y(_0915_),
    .A1(_0895_),
    .A2(_0899_));
 sg13g2_o21ai_1 _3234_ (.B1(_0915_),
    .Y(\MemCell.next_state[2] ),
    .A1(net722),
    .A2(_0908_));
 sg13g2_nand2b_1 _3235_ (.Y(_0916_),
    .B(\MemCell.dc1_reg[1][6] ),
    .A_N(net776));
 sg13g2_nor2b_1 _3236_ (.A(net776),
    .B_N(\MemCell.dc1_reg[1][7] ),
    .Y(_0917_));
 sg13g2_nor2_1 _3237_ (.A(_0153_),
    .B(_0917_),
    .Y(_0918_));
 sg13g2_xnor2_1 _3238_ (.Y(_0919_),
    .A(\pwm_module.counter0[14] ),
    .B(_0916_));
 sg13g2_nor2_1 _3239_ (.A(_0918_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_nor2b_1 _3240_ (.A(net776),
    .B_N(\MemCell.dc1_reg[1][5] ),
    .Y(_0921_));
 sg13g2_nand3_1 _3241_ (.B(_0920_),
    .C(_0921_),
    .A(_0154_),
    .Y(_0922_));
 sg13g2_nand2_1 _3242_ (.Y(_0923_),
    .A(_0153_),
    .B(_0917_));
 sg13g2_or3_1 _3243_ (.A(\pwm_module.counter0[14] ),
    .B(_0916_),
    .C(_0918_),
    .X(_0924_));
 sg13g2_xor2_1 _3244_ (.B(_0921_),
    .A(\pwm_module.counter0[13] ),
    .X(_0925_));
 sg13g2_nand2b_1 _3245_ (.Y(_0926_),
    .B(\MemCell.dc1_reg[1][4] ),
    .A_N(net776));
 sg13g2_a21oi_1 _3246_ (.A1(\pwm_module.counter0[12] ),
    .A2(_0926_),
    .Y(_0927_),
    .B1(_0925_));
 sg13g2_nand2_1 _3247_ (.Y(_0928_),
    .A(_0920_),
    .B(_0927_));
 sg13g2_nor2b_1 _3248_ (.A(net775),
    .B_N(\MemCell.dc1_reg[1][2] ),
    .Y(_0929_));
 sg13g2_xnor2_1 _3249_ (.Y(_0930_),
    .A(\pwm_module.counter0[10] ),
    .B(_0929_));
 sg13g2_nand3b_1 _3250_ (.B(\MemCell.dc1_reg[1][3] ),
    .C(_0156_),
    .Y(_0931_),
    .A_N(net775));
 sg13g2_a21o_1 _3251_ (.A2(\MemCell.dc1_reg[1][3] ),
    .A1(_2347_),
    .B1(_0156_),
    .X(_0932_));
 sg13g2_nand3_1 _3252_ (.B(_0931_),
    .C(_0932_),
    .A(_0930_),
    .Y(_0933_));
 sg13g2_nor2_1 _3253_ (.A(net775),
    .B(\MemCell.dc1_reg[1][1] ),
    .Y(_0934_));
 sg13g2_nor2_1 _3254_ (.A(\pwm_module.counter0[9] ),
    .B(_0934_),
    .Y(_0935_));
 sg13g2_xnor2_1 _3255_ (.Y(_0936_),
    .A(_0158_),
    .B(_0934_));
 sg13g2_nand2b_1 _3256_ (.Y(_0937_),
    .B(\MemCell.dc1_reg[1][0] ),
    .A_N(net776));
 sg13g2_nor2_1 _3257_ (.A(\pwm_module.counter0[8] ),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_a21oi_1 _3258_ (.A1(_0936_),
    .A2(_0938_),
    .Y(_0939_),
    .B1(_0935_));
 sg13g2_and2_1 _3259_ (.A(_0157_),
    .B(_0929_),
    .X(_0940_));
 sg13g2_nor2_1 _3260_ (.A(\pwm_module.counter0[12] ),
    .B(_0926_),
    .Y(_0941_));
 sg13g2_o21ai_1 _3261_ (.B1(_0931_),
    .Y(_0942_),
    .A1(\pwm_module.counter0[12] ),
    .A2(_0926_));
 sg13g2_a21oi_1 _3262_ (.A1(_0932_),
    .A2(_0940_),
    .Y(_0943_),
    .B1(_0942_));
 sg13g2_o21ai_1 _3263_ (.B1(_0943_),
    .Y(_0944_),
    .A1(_0933_),
    .A2(_0939_));
 sg13g2_nor2_1 _3264_ (.A(net777),
    .B(\MemCell.dc1_reg[0][6] ),
    .Y(_0945_));
 sg13g2_xor2_1 _3265_ (.B(_0945_),
    .A(_0160_),
    .X(_0946_));
 sg13g2_nor2_1 _3266_ (.A(net777),
    .B(\MemCell.dc1_reg[0][5] ),
    .Y(_0947_));
 sg13g2_nor2_1 _3267_ (.A(\pwm_module.counter0[5] ),
    .B(_0947_),
    .Y(_0948_));
 sg13g2_nor3_1 _3268_ (.A(net777),
    .B(\MemCell.dc1_reg[0][4] ),
    .C(_0162_),
    .Y(_0949_));
 sg13g2_xor2_1 _3269_ (.B(_0947_),
    .A(_0161_),
    .X(_0950_));
 sg13g2_nor2_1 _3270_ (.A(_0949_),
    .B(_0950_),
    .Y(_0951_));
 sg13g2_o21ai_1 _3271_ (.B1(_0162_),
    .Y(_0952_),
    .A1(net777),
    .A2(\MemCell.dc1_reg[0][4] ));
 sg13g2_nor2b_2 _3272_ (.A(net775),
    .B_N(\MemCell.dc1_reg[0][3] ),
    .Y(_0953_));
 sg13g2_nor2_1 _3273_ (.A(_0163_),
    .B(_0953_),
    .Y(_0954_));
 sg13g2_nand2b_1 _3274_ (.Y(_0955_),
    .B(\MemCell.dc1_reg[0][2] ),
    .A_N(net775));
 sg13g2_nor2_1 _3275_ (.A(\pwm_module.counter0[2] ),
    .B(_0955_),
    .Y(_0956_));
 sg13g2_a21oi_1 _3276_ (.A1(_0163_),
    .A2(_0953_),
    .Y(_0957_),
    .B1(_0956_));
 sg13g2_nand2b_1 _3277_ (.Y(_0958_),
    .B(\MemCell.dc1_reg[0][1] ),
    .A_N(net775));
 sg13g2_a22oi_1 _3278_ (.Y(_0959_),
    .B1(_0958_),
    .B2(_2355_),
    .A2(_0955_),
    .A1(\pwm_module.counter0[2] ));
 sg13g2_nand3b_1 _3279_ (.B(\MemCell.dc1_reg[0][1] ),
    .C(_0164_),
    .Y(_0960_),
    .A_N(net775));
 sg13g2_nor2_1 _3280_ (.A(net775),
    .B(\MemCell.dc1_reg[0][0] ),
    .Y(_0961_));
 sg13g2_nand3_1 _3281_ (.B(_0960_),
    .C(_0961_),
    .A(net754),
    .Y(_0962_));
 sg13g2_a221oi_1 _3282_ (.B2(_0962_),
    .C1(_0956_),
    .B1(_0959_),
    .A1(_0163_),
    .Y(_0963_),
    .A2(_0953_));
 sg13g2_o21ai_1 _3283_ (.B1(_0952_),
    .Y(_0964_),
    .A1(_0954_),
    .A2(_0963_));
 sg13g2_a21oi_1 _3284_ (.A1(_0951_),
    .A2(_0964_),
    .Y(_0965_),
    .B1(_0948_));
 sg13g2_nor2b_1 _3285_ (.A(net777),
    .B_N(\MemCell.dc1_reg[0][7] ),
    .Y(_0966_));
 sg13g2_nand2_1 _3286_ (.Y(_0967_),
    .A(_0159_),
    .B(_0966_));
 sg13g2_o21ai_1 _3287_ (.B1(_0967_),
    .Y(_0968_),
    .A1(\pwm_module.counter0[6] ),
    .A2(_0945_));
 sg13g2_inv_1 _3288_ (.Y(_0969_),
    .A(_0968_));
 sg13g2_o21ai_1 _3289_ (.B1(_0969_),
    .Y(_0970_),
    .A1(_0946_),
    .A2(_0965_));
 sg13g2_nor2_1 _3290_ (.A(_0938_),
    .B(_0941_),
    .Y(_0971_));
 sg13g2_o21ai_1 _3291_ (.B1(_0923_),
    .Y(_0972_),
    .A1(_0159_),
    .A2(_0966_));
 sg13g2_a21oi_1 _3292_ (.A1(\pwm_module.counter0[8] ),
    .A2(_0937_),
    .Y(_0973_),
    .B1(_0972_));
 sg13g2_nand3_1 _3293_ (.B(_0971_),
    .C(_0973_),
    .A(_0936_),
    .Y(_0974_));
 sg13g2_nor3_1 _3294_ (.A(_0928_),
    .B(_0933_),
    .C(_0974_),
    .Y(_0975_));
 sg13g2_nand2b_1 _3295_ (.Y(_0976_),
    .B(_0944_),
    .A_N(_0928_));
 sg13g2_nand4_1 _3296_ (.B(_0923_),
    .C(_0924_),
    .A(_0922_),
    .Y(_0977_),
    .D(_0976_));
 sg13g2_a21oi_1 _3297_ (.A1(_0970_),
    .A2(_0975_),
    .Y(_0978_),
    .B1(_0977_));
 sg13g2_nand2_1 _3298_ (.Y(_0979_),
    .A(net762),
    .B(\MemCell.dc1_reg[3][2] ));
 sg13g2_nand2_1 _3299_ (.Y(_0980_),
    .A(\pwm_module.counter0[26] ),
    .B(_0979_));
 sg13g2_nor2b_1 _3300_ (.A(net778),
    .B_N(\MemCell.dc1_reg[3][3] ),
    .Y(_0981_));
 sg13g2_o21ai_1 _3301_ (.B1(_0980_),
    .Y(_0982_),
    .A1(_0146_),
    .A2(_0981_));
 sg13g2_nand3_1 _3302_ (.B(net762),
    .C(_0167_),
    .A(\MemCell.dc1_reg[3][7] ),
    .Y(_0983_));
 sg13g2_nand2_1 _3303_ (.Y(_0984_),
    .A(net761),
    .B(\MemCell.dc1_reg[3][4] ));
 sg13g2_nand2_1 _3304_ (.Y(_0985_),
    .A(\pwm_module.counter0[28] ),
    .B(_0984_));
 sg13g2_nand2_1 _3305_ (.Y(_0986_),
    .A(_0983_),
    .B(_0985_));
 sg13g2_nand2_1 _3306_ (.Y(_0987_),
    .A(net761),
    .B(\MemCell.dc1_reg[3][6] ));
 sg13g2_nor2b_1 _3307_ (.A(net778),
    .B_N(\MemCell.dc1_reg[3][5] ),
    .Y(_0988_));
 sg13g2_nand2_1 _3308_ (.Y(_0989_),
    .A(_0145_),
    .B(_0988_));
 sg13g2_o21ai_1 _3309_ (.B1(_0989_),
    .Y(_0990_),
    .A1(\pwm_module.counter0[30] ),
    .A2(_0987_));
 sg13g2_a21oi_1 _3310_ (.A1(\MemCell.dc1_reg[3][7] ),
    .A2(net762),
    .Y(_0991_),
    .B1(_0167_));
 sg13g2_a21o_1 _3311_ (.A2(_0987_),
    .A1(\pwm_module.counter0[30] ),
    .B1(_0991_),
    .X(_0992_));
 sg13g2_nor4_1 _3312_ (.A(_0982_),
    .B(_0986_),
    .C(_0990_),
    .D(_0992_),
    .Y(_0993_));
 sg13g2_nand2_1 _3313_ (.Y(_0994_),
    .A(net762),
    .B(\MemCell.dc1_reg[3][0] ));
 sg13g2_nor2_1 _3314_ (.A(\pwm_module.counter0[24] ),
    .B(_0994_),
    .Y(_0995_));
 sg13g2_nand2_1 _3315_ (.Y(_0996_),
    .A(\pwm_module.counter0[24] ),
    .B(_0994_));
 sg13g2_nor2b_1 _3316_ (.A(net778),
    .B_N(\MemCell.dc1_reg[3][1] ),
    .Y(_0997_));
 sg13g2_nor2_1 _3317_ (.A(_0147_),
    .B(_0997_),
    .Y(_0998_));
 sg13g2_o21ai_1 _3318_ (.B1(_0996_),
    .Y(_0999_),
    .A1(_0145_),
    .A2(_0988_));
 sg13g2_nor3_1 _3319_ (.A(_0995_),
    .B(_0998_),
    .C(_0999_),
    .Y(_1000_));
 sg13g2_nor2_1 _3320_ (.A(\pwm_module.counter0[28] ),
    .B(_0984_),
    .Y(_1001_));
 sg13g2_a21oi_1 _3321_ (.A1(_0146_),
    .A2(_0981_),
    .Y(_1002_),
    .B1(_1001_));
 sg13g2_nor2_1 _3322_ (.A(\pwm_module.counter0[26] ),
    .B(_0979_),
    .Y(_1003_));
 sg13g2_a21oi_1 _3323_ (.A1(_0147_),
    .A2(_0997_),
    .Y(_1004_),
    .B1(_1003_));
 sg13g2_and2_1 _3324_ (.A(_1002_),
    .B(_1004_),
    .X(_1005_));
 sg13g2_nand3_1 _3325_ (.B(_1000_),
    .C(_1005_),
    .A(_0993_),
    .Y(_1006_));
 sg13g2_nor2b_1 _3326_ (.A(net778),
    .B_N(\MemCell.dc1_reg[2][3] ),
    .Y(_1007_));
 sg13g2_nor2_1 _3327_ (.A(_0151_),
    .B(_1007_),
    .Y(_1008_));
 sg13g2_nand3_1 _3328_ (.B(\MemCell.dc1_reg[2][7] ),
    .C(_0148_),
    .A(net761),
    .Y(_1009_));
 sg13g2_nand2b_1 _3329_ (.Y(_1010_),
    .B(_1009_),
    .A_N(_1008_));
 sg13g2_nand2_2 _3330_ (.Y(_1011_),
    .A(net761),
    .B(\MemCell.dc1_reg[2][6] ));
 sg13g2_nor2_1 _3331_ (.A(\pwm_module.counter0[22] ),
    .B(_1011_),
    .Y(_1012_));
 sg13g2_a21oi_1 _3332_ (.A1(net761),
    .A2(\MemCell.dc1_reg[2][7] ),
    .Y(_1013_),
    .B1(_0148_));
 sg13g2_nand2_1 _3333_ (.Y(_1014_),
    .A(net761),
    .B(\MemCell.dc1_reg[2][4] ));
 sg13g2_nor2_1 _3334_ (.A(\pwm_module.counter0[20] ),
    .B(_1014_),
    .Y(_1015_));
 sg13g2_nor2b_1 _3335_ (.A(net778),
    .B_N(\MemCell.dc1_reg[2][0] ),
    .Y(_1016_));
 sg13g2_nor2_1 _3336_ (.A(_2352_),
    .B(_1016_),
    .Y(_1017_));
 sg13g2_or4_1 _3337_ (.A(_1012_),
    .B(_1013_),
    .C(_1015_),
    .D(_1017_),
    .X(_1018_));
 sg13g2_nand2b_1 _3338_ (.Y(_1019_),
    .B(\MemCell.dc1_reg[2][2] ),
    .A_N(net778));
 sg13g2_nor2_1 _3339_ (.A(\pwm_module.counter0[18] ),
    .B(_1019_),
    .Y(_1020_));
 sg13g2_a21o_1 _3340_ (.A2(_1007_),
    .A1(_0151_),
    .B1(_1020_),
    .X(_1021_));
 sg13g2_nor2b_1 _3341_ (.A(net778),
    .B_N(\MemCell.dc1_reg[2][1] ),
    .Y(_1022_));
 sg13g2_a221oi_1 _3342_ (.B2(_0152_),
    .C1(_1021_),
    .B1(_1022_),
    .A1(_2352_),
    .Y(_1023_),
    .A2(_1016_));
 sg13g2_nand2_1 _3343_ (.Y(_1024_),
    .A(net761),
    .B(\MemCell.dc1_reg[2][5] ));
 sg13g2_xnor2_1 _3344_ (.Y(_1025_),
    .A(\pwm_module.counter0[21] ),
    .B(_1024_));
 sg13g2_a21oi_1 _3345_ (.A1(\pwm_module.counter0[20] ),
    .A2(_1014_),
    .Y(_1026_),
    .B1(_1025_));
 sg13g2_nand2_1 _3346_ (.Y(_1027_),
    .A(\pwm_module.counter0[18] ),
    .B(_1019_));
 sg13g2_nor2_1 _3347_ (.A(_0152_),
    .B(_1022_),
    .Y(_1028_));
 sg13g2_or2_1 _3348_ (.X(_1029_),
    .B(_1022_),
    .A(_0152_));
 sg13g2_a21oi_1 _3349_ (.A1(\pwm_module.counter0[22] ),
    .A2(_1011_),
    .Y(_1030_),
    .B1(_1028_));
 sg13g2_nand4_1 _3350_ (.B(_1026_),
    .C(_1027_),
    .A(_1023_),
    .Y(_1031_),
    .D(_1030_));
 sg13g2_nor4_2 _3351_ (.A(_1006_),
    .B(_1010_),
    .C(_1018_),
    .Y(_1032_),
    .D(_1031_));
 sg13g2_nand2b_1 _3352_ (.Y(_1033_),
    .B(_1032_),
    .A_N(_0978_));
 sg13g2_nand2b_1 _3353_ (.Y(_1034_),
    .B(_0995_),
    .A_N(_0998_));
 sg13g2_o21ai_1 _3354_ (.B1(_0985_),
    .Y(_1035_),
    .A1(_0145_),
    .A2(_0988_));
 sg13g2_a221oi_1 _3355_ (.B2(_1034_),
    .C1(_1035_),
    .B1(_1005_),
    .A1(_0982_),
    .Y(_1036_),
    .A2(_1002_));
 sg13g2_nor2_1 _3356_ (.A(_0990_),
    .B(_1036_),
    .Y(_1037_));
 sg13g2_or2_1 _3357_ (.X(_1038_),
    .B(_1037_),
    .A(_0992_));
 sg13g2_a21oi_1 _3358_ (.A1(_1027_),
    .A2(_1029_),
    .Y(_1039_),
    .B1(_1021_));
 sg13g2_nor3_1 _3359_ (.A(_1008_),
    .B(_1023_),
    .C(_1039_),
    .Y(_1040_));
 sg13g2_o21ai_1 _3360_ (.B1(_1026_),
    .Y(_1041_),
    .A1(_1015_),
    .A2(_1040_));
 sg13g2_nand3_1 _3361_ (.B(\MemCell.dc1_reg[2][5] ),
    .C(_0149_),
    .A(net761),
    .Y(_1042_));
 sg13g2_a22oi_1 _3362_ (.Y(_1043_),
    .B1(_1041_),
    .B2(_1042_),
    .A2(_1011_),
    .A1(\pwm_module.counter0[22] ));
 sg13g2_o21ai_1 _3363_ (.B1(_1009_),
    .Y(_1044_),
    .A1(\pwm_module.counter0[22] ),
    .A2(_1011_));
 sg13g2_nor2_1 _3364_ (.A(_1006_),
    .B(_1013_),
    .Y(_1045_));
 sg13g2_o21ai_1 _3365_ (.B1(_1045_),
    .Y(_1046_),
    .A1(_1043_),
    .A2(_1044_));
 sg13g2_nand4_1 _3366_ (.B(_1033_),
    .C(_1038_),
    .A(_0983_),
    .Y(_1047_),
    .D(_1046_));
 sg13g2_o21ai_1 _3367_ (.B1(_0952_),
    .Y(_1048_),
    .A1(_0163_),
    .A2(_0953_));
 sg13g2_nor2_1 _3368_ (.A(_0946_),
    .B(_1048_),
    .Y(_1049_));
 sg13g2_xnor2_1 _3369_ (.Y(_1050_),
    .A(_0165_),
    .B(_0961_));
 sg13g2_and4_1 _3370_ (.A(_0951_),
    .B(_0960_),
    .C(_0967_),
    .D(_1050_),
    .X(_1051_));
 sg13g2_and4_1 _3371_ (.A(_0957_),
    .B(_0959_),
    .C(_1049_),
    .D(_1051_),
    .X(_1052_));
 sg13g2_nand3_1 _3372_ (.B(_1032_),
    .C(_1052_),
    .A(_0975_),
    .Y(_1053_));
 sg13g2_and3_2 _3373_ (.X(_0096_),
    .A(_2396_),
    .B(_1047_),
    .C(_1053_));
 sg13g2_nand2_1 _3374_ (.Y(_1054_),
    .A(net757),
    .B(\MemCell.dc2_reg[3][6] ));
 sg13g2_nor2_1 _3375_ (.A(\pwm_module.counter1[30] ),
    .B(_1054_),
    .Y(_1055_));
 sg13g2_nor2b_1 _3376_ (.A(net774),
    .B_N(\MemCell.dc2_reg[3][7] ),
    .Y(_1056_));
 sg13g2_a21oi_1 _3377_ (.A1(_0202_),
    .A2(_1056_),
    .Y(_1057_),
    .B1(_1055_));
 sg13g2_nor2_1 _3378_ (.A(_0202_),
    .B(_1056_),
    .Y(_1058_));
 sg13g2_or2_1 _3379_ (.X(_1059_),
    .B(_1058_),
    .A(_1057_));
 sg13g2_nor2b_1 _3380_ (.A(net774),
    .B_N(\MemCell.dc2_reg[3][5] ),
    .Y(_1060_));
 sg13g2_a21oi_1 _3381_ (.A1(\pwm_module.counter1[30] ),
    .A2(_1054_),
    .Y(_1061_),
    .B1(_1058_));
 sg13g2_o21ai_1 _3382_ (.B1(_1061_),
    .Y(_1062_),
    .A1(_0103_),
    .A2(_1060_));
 sg13g2_and2_1 _3383_ (.A(_0103_),
    .B(_1060_),
    .X(_1063_));
 sg13g2_nand2_1 _3384_ (.Y(_1064_),
    .A(net757),
    .B(\MemCell.dc2_reg[3][4] ));
 sg13g2_nand2_1 _3385_ (.Y(_1065_),
    .A(\pwm_module.counter1[28] ),
    .B(_1064_));
 sg13g2_nand3_1 _3386_ (.B(\MemCell.dc2_reg[3][3] ),
    .C(_0104_),
    .A(net757),
    .Y(_1066_));
 sg13g2_o21ai_1 _3387_ (.B1(_1066_),
    .Y(_1067_),
    .A1(\pwm_module.counter1[28] ),
    .A2(_1064_));
 sg13g2_nand2_1 _3388_ (.Y(_1068_),
    .A(net757),
    .B(\MemCell.dc2_reg[3][2] ));
 sg13g2_a21oi_1 _3389_ (.A1(net757),
    .A2(\MemCell.dc2_reg[3][3] ),
    .Y(_1069_),
    .B1(_0104_));
 sg13g2_a21oi_1 _3390_ (.A1(\pwm_module.counter1[26] ),
    .A2(_1068_),
    .Y(_1070_),
    .B1(_1069_));
 sg13g2_nand3_1 _3391_ (.B(\MemCell.dc2_reg[3][1] ),
    .C(_0105_),
    .A(net757),
    .Y(_1071_));
 sg13g2_o21ai_1 _3392_ (.B1(_1071_),
    .Y(_1072_),
    .A1(\pwm_module.counter1[26] ),
    .A2(_1068_));
 sg13g2_a21o_1 _3393_ (.A2(\MemCell.dc2_reg[3][1] ),
    .A1(net757),
    .B1(_0105_),
    .X(_1073_));
 sg13g2_nand2_1 _3394_ (.Y(_1074_),
    .A(net757),
    .B(\MemCell.dc2_reg[3][0] ));
 sg13g2_nor2_1 _3395_ (.A(\pwm_module.counter1[24] ),
    .B(_1074_),
    .Y(_1075_));
 sg13g2_a21o_1 _3396_ (.A2(_1075_),
    .A1(_1073_),
    .B1(_1072_),
    .X(_1076_));
 sg13g2_a21o_1 _3397_ (.A2(_1076_),
    .A1(_1070_),
    .B1(_1067_),
    .X(_1077_));
 sg13g2_a21oi_1 _3398_ (.A1(_1065_),
    .A2(_1077_),
    .Y(_1078_),
    .B1(_1063_));
 sg13g2_o21ai_1 _3399_ (.B1(_1059_),
    .Y(_1079_),
    .A1(_1062_),
    .A2(_1078_));
 sg13g2_nand2_1 _3400_ (.Y(_1080_),
    .A(_1057_),
    .B(_1070_));
 sg13g2_nand2_1 _3401_ (.Y(_1081_),
    .A(\pwm_module.counter1[24] ),
    .B(_1074_));
 sg13g2_nor3_1 _3402_ (.A(_1063_),
    .B(_1072_),
    .C(_1075_),
    .Y(_1082_));
 sg13g2_nand4_1 _3403_ (.B(_1073_),
    .C(_1081_),
    .A(_1065_),
    .Y(_1083_),
    .D(_1082_));
 sg13g2_nor4_2 _3404_ (.A(_1062_),
    .B(_1067_),
    .C(_1080_),
    .Y(_1084_),
    .D(_1083_));
 sg13g2_nand3_1 _3405_ (.B(\MemCell.dc2_reg[2][7] ),
    .C(_0106_),
    .A(net759),
    .Y(_1085_));
 sg13g2_nand2_1 _3406_ (.Y(_1086_),
    .A(net759),
    .B(\MemCell.dc2_reg[2][6] ));
 sg13g2_a21oi_1 _3407_ (.A1(net758),
    .A2(\MemCell.dc2_reg[2][6] ),
    .Y(_1087_),
    .B1(_2360_));
 sg13g2_a21oi_1 _3408_ (.A1(net759),
    .A2(\MemCell.dc2_reg[2][7] ),
    .Y(_1088_),
    .B1(_0106_));
 sg13g2_nor2_1 _3409_ (.A(_1087_),
    .B(_1088_),
    .Y(_1089_));
 sg13g2_nor2b_2 _3410_ (.A(net774),
    .B_N(\MemCell.dc2_reg[2][5] ),
    .Y(_1090_));
 sg13g2_nand2_1 _3411_ (.Y(_1091_),
    .A(net759),
    .B(\MemCell.dc2_reg[2][4] ));
 sg13g2_a22oi_1 _3412_ (.Y(_1092_),
    .B1(_1091_),
    .B2(\pwm_module.counter1[20] ),
    .A2(_1090_),
    .A1(_2362_));
 sg13g2_o21ai_1 _3413_ (.B1(_1092_),
    .Y(_1093_),
    .A1(_2362_),
    .A2(_1090_));
 sg13g2_nand2b_1 _3414_ (.Y(_1094_),
    .B(\MemCell.dc2_reg[2][0] ),
    .A_N(net774));
 sg13g2_nand3b_1 _3415_ (.B(\MemCell.dc2_reg[2][1] ),
    .C(_0110_),
    .Y(_1095_),
    .A_N(net774));
 sg13g2_o21ai_1 _3416_ (.B1(_1095_),
    .Y(_1096_),
    .A1(\pwm_module.counter1[16] ),
    .A2(_1094_));
 sg13g2_nand2b_1 _3417_ (.Y(_1097_),
    .B(\MemCell.dc2_reg[2][2] ),
    .A_N(net774));
 sg13g2_a21oi_1 _3418_ (.A1(net758),
    .A2(\MemCell.dc2_reg[2][3] ),
    .Y(_1098_),
    .B1(_0109_));
 sg13g2_a21oi_1 _3419_ (.A1(\pwm_module.counter1[18] ),
    .A2(_1097_),
    .Y(_1099_),
    .B1(_1098_));
 sg13g2_a21o_1 _3420_ (.A2(\MemCell.dc2_reg[2][1] ),
    .A1(net758),
    .B1(_0110_),
    .X(_1100_));
 sg13g2_nand2_1 _3421_ (.Y(_1101_),
    .A(_1099_),
    .B(_1100_));
 sg13g2_nand3_1 _3422_ (.B(\MemCell.dc2_reg[2][3] ),
    .C(_0109_),
    .A(net758),
    .Y(_1102_));
 sg13g2_o21ai_1 _3423_ (.B1(_1102_),
    .Y(_1103_),
    .A1(\pwm_module.counter1[20] ),
    .A2(_1091_));
 sg13g2_nor2_1 _3424_ (.A(\pwm_module.counter1[18] ),
    .B(_1097_),
    .Y(_1104_));
 sg13g2_a21o_1 _3425_ (.A2(_1100_),
    .A1(_1096_),
    .B1(_1104_),
    .X(_1105_));
 sg13g2_a21oi_1 _3426_ (.A1(_1099_),
    .A2(_1105_),
    .Y(_1106_),
    .B1(_1103_));
 sg13g2_nor2_1 _3427_ (.A(\pwm_module.counter1[22] ),
    .B(_1086_),
    .Y(_1107_));
 sg13g2_nand2_1 _3428_ (.Y(_1108_),
    .A(_0107_),
    .B(_1090_));
 sg13g2_o21ai_1 _3429_ (.B1(_1108_),
    .Y(_1109_),
    .A1(_1093_),
    .A2(_1106_));
 sg13g2_o21ai_1 _3430_ (.B1(_1089_),
    .Y(_1110_),
    .A1(_1107_),
    .A2(_1109_));
 sg13g2_nand2_1 _3431_ (.Y(_1111_),
    .A(_1085_),
    .B(_1110_));
 sg13g2_nor2b_1 _3432_ (.A(net772),
    .B_N(\MemCell.dc2_reg[0][7] ),
    .Y(_1112_));
 sg13g2_nand2_1 _3433_ (.Y(_1113_),
    .A(_0117_),
    .B(_1112_));
 sg13g2_or2_1 _3434_ (.X(_1114_),
    .B(\MemCell.dc2_reg[0][6] ),
    .A(net772));
 sg13g2_a22oi_1 _3435_ (.Y(_1115_),
    .B1(_1114_),
    .B2(_2365_),
    .A2(_1112_),
    .A1(_0117_));
 sg13g2_xnor2_1 _3436_ (.Y(_1116_),
    .A(_0118_),
    .B(_1114_));
 sg13g2_nor2_1 _3437_ (.A(net772),
    .B(\MemCell.dc2_reg[0][5] ),
    .Y(_1117_));
 sg13g2_nor2_1 _3438_ (.A(\pwm_module.counter1[5] ),
    .B(_1117_),
    .Y(_1118_));
 sg13g2_xnor2_1 _3439_ (.Y(_1119_),
    .A(_0119_),
    .B(_1117_));
 sg13g2_o21ai_1 _3440_ (.B1(_0120_),
    .Y(_1120_),
    .A1(net772),
    .A2(\MemCell.dc2_reg[0][4] ));
 sg13g2_nor2b_1 _3441_ (.A(net772),
    .B_N(\MemCell.dc2_reg[0][3] ),
    .Y(_1121_));
 sg13g2_nand2_1 _3442_ (.Y(_1122_),
    .A(_0121_),
    .B(_1121_));
 sg13g2_nand2b_1 _3443_ (.Y(_1123_),
    .B(\MemCell.dc2_reg[0][2] ),
    .A_N(net773));
 sg13g2_o21ai_1 _3444_ (.B1(_1122_),
    .Y(_1124_),
    .A1(\pwm_module.counter1[2] ),
    .A2(_1123_));
 sg13g2_nand2_1 _3445_ (.Y(_1125_),
    .A(\pwm_module.counter1[2] ),
    .B(_1123_));
 sg13g2_nand2b_1 _3446_ (.Y(_1126_),
    .B(\MemCell.dc2_reg[0][1] ),
    .A_N(net772));
 sg13g2_nor2_1 _3447_ (.A(_2369_),
    .B(_1126_),
    .Y(_1127_));
 sg13g2_nor2_1 _3448_ (.A(net772),
    .B(\MemCell.dc2_reg[0][0] ),
    .Y(_1128_));
 sg13g2_a22oi_1 _3449_ (.Y(_1129_),
    .B1(_1128_),
    .B2(\pwm_module.counter1[0] ),
    .A2(_1126_),
    .A1(_2369_));
 sg13g2_o21ai_1 _3450_ (.B1(_1125_),
    .Y(_1130_),
    .A1(_1127_),
    .A2(_1129_));
 sg13g2_nor2b_1 _3451_ (.A(_1124_),
    .B_N(_1130_),
    .Y(_1131_));
 sg13g2_or3_1 _3452_ (.A(net772),
    .B(\MemCell.dc2_reg[0][4] ),
    .C(_0120_),
    .X(_1132_));
 sg13g2_o21ai_1 _3453_ (.B1(_1132_),
    .Y(_1133_),
    .A1(_0121_),
    .A2(_1121_));
 sg13g2_o21ai_1 _3454_ (.B1(_1120_),
    .Y(_1134_),
    .A1(_1131_),
    .A2(_1133_));
 sg13g2_a21oi_1 _3455_ (.A1(_1119_),
    .A2(_1134_),
    .Y(_1135_),
    .B1(_1118_));
 sg13g2_o21ai_1 _3456_ (.B1(_1115_),
    .Y(_1136_),
    .A1(_1116_),
    .A2(_1135_));
 sg13g2_nor2_1 _3457_ (.A(_0117_),
    .B(_1112_),
    .Y(_1137_));
 sg13g2_nor2b_1 _3458_ (.A(net773),
    .B_N(\MemCell.dc2_reg[1][7] ),
    .Y(_1138_));
 sg13g2_nor2_1 _3459_ (.A(_0111_),
    .B(_1138_),
    .Y(_1139_));
 sg13g2_inv_1 _3460_ (.Y(_1140_),
    .A(_1139_));
 sg13g2_nand2_1 _3461_ (.Y(_1141_),
    .A(net760),
    .B(\MemCell.dc2_reg[1][6] ));
 sg13g2_a21oi_1 _3462_ (.A1(\pwm_module.counter1[14] ),
    .A2(_1141_),
    .Y(_1142_),
    .B1(_1139_));
 sg13g2_nor2_1 _3463_ (.A(net773),
    .B(\MemCell.dc2_reg[1][1] ),
    .Y(_1143_));
 sg13g2_xnor2_1 _3464_ (.Y(_1144_),
    .A(_0116_),
    .B(_1143_));
 sg13g2_nor2_1 _3465_ (.A(\pwm_module.counter1[14] ),
    .B(_1141_),
    .Y(_1145_));
 sg13g2_a21oi_1 _3466_ (.A1(_0111_),
    .A2(_1138_),
    .Y(_1146_),
    .B1(_1145_));
 sg13g2_inv_1 _3467_ (.Y(_1147_),
    .A(_1146_));
 sg13g2_nand3_1 _3468_ (.B(_1144_),
    .C(_1146_),
    .A(_1142_),
    .Y(_1148_));
 sg13g2_nand2_1 _3469_ (.Y(_1149_),
    .A(net760),
    .B(\MemCell.dc2_reg[1][5] ));
 sg13g2_nand2_1 _3470_ (.Y(_1150_),
    .A(net759),
    .B(\MemCell.dc2_reg[1][4] ));
 sg13g2_xnor2_1 _3471_ (.Y(_1151_),
    .A(\pwm_module.counter1[13] ),
    .B(_1149_));
 sg13g2_a21o_1 _3472_ (.A2(_1150_),
    .A1(\pwm_module.counter1[12] ),
    .B1(_1151_),
    .X(_1152_));
 sg13g2_nor2b_1 _3473_ (.A(net773),
    .B_N(\MemCell.dc2_reg[1][3] ),
    .Y(_1153_));
 sg13g2_nor2_1 _3474_ (.A(_0114_),
    .B(_1153_),
    .Y(_1154_));
 sg13g2_and3_1 _3475_ (.X(_1155_),
    .A(net759),
    .B(\MemCell.dc2_reg[1][0] ),
    .C(_2364_));
 sg13g2_a21oi_1 _3476_ (.A1(net759),
    .A2(\MemCell.dc2_reg[1][0] ),
    .Y(_1156_),
    .B1(_2364_));
 sg13g2_nor3_1 _3477_ (.A(_1154_),
    .B(_1155_),
    .C(_1156_),
    .Y(_1157_));
 sg13g2_nor2_1 _3478_ (.A(\pwm_module.counter1[12] ),
    .B(_1150_),
    .Y(_1158_));
 sg13g2_a21oi_1 _3479_ (.A1(_0114_),
    .A2(_1153_),
    .Y(_1159_),
    .B1(_1158_));
 sg13g2_nor2b_1 _3480_ (.A(net773),
    .B_N(\MemCell.dc2_reg[1][2] ),
    .Y(_1160_));
 sg13g2_xor2_1 _3481_ (.B(_1160_),
    .A(\pwm_module.counter1[10] ),
    .X(_1161_));
 sg13g2_nand3b_1 _3482_ (.B(_1159_),
    .C(_1157_),
    .Y(_1162_),
    .A_N(_1161_));
 sg13g2_nor3_1 _3483_ (.A(_1148_),
    .B(_1152_),
    .C(_1162_),
    .Y(_1163_));
 sg13g2_nor2b_1 _3484_ (.A(_1137_),
    .B_N(_1163_),
    .Y(_1164_));
 sg13g2_nor2_1 _3485_ (.A(\pwm_module.counter1[9] ),
    .B(_1143_),
    .Y(_1165_));
 sg13g2_a21oi_1 _3486_ (.A1(_1144_),
    .A2(_1155_),
    .Y(_1166_),
    .B1(_1165_));
 sg13g2_nand2_1 _3487_ (.Y(_1167_),
    .A(_0115_),
    .B(_1160_));
 sg13g2_o21ai_1 _3488_ (.B1(_1167_),
    .Y(_1168_),
    .A1(_1161_),
    .A2(_1166_));
 sg13g2_nand2b_1 _3489_ (.Y(_1169_),
    .B(_1168_),
    .A_N(_1154_));
 sg13g2_a21o_1 _3490_ (.A2(_1169_),
    .A1(_1159_),
    .B1(_1152_),
    .X(_1170_));
 sg13g2_nand3_1 _3491_ (.B(\MemCell.dc2_reg[1][5] ),
    .C(_0112_),
    .A(net759),
    .Y(_1171_));
 sg13g2_nand2b_1 _3492_ (.Y(_1172_),
    .B(_1142_),
    .A_N(_1145_));
 sg13g2_a21oi_1 _3493_ (.A1(_1170_),
    .A2(_1171_),
    .Y(_1173_),
    .B1(_1172_));
 sg13g2_nor2_1 _3494_ (.A(_1116_),
    .B(_1137_),
    .Y(_1174_));
 sg13g2_nor2b_1 _3495_ (.A(_1133_),
    .B_N(_1120_),
    .Y(_1175_));
 sg13g2_nand4_1 _3496_ (.B(_1119_),
    .C(_1174_),
    .A(_1113_),
    .Y(_1176_),
    .D(_1175_));
 sg13g2_a221oi_1 _3497_ (.B2(_1136_),
    .C1(_1173_),
    .B1(_1164_),
    .A1(_1140_),
    .Y(_1177_),
    .A2(_1147_));
 sg13g2_or4_1 _3498_ (.A(_1087_),
    .B(_1088_),
    .C(_1096_),
    .D(_1103_),
    .X(_1178_));
 sg13g2_o21ai_1 _3499_ (.B1(_1085_),
    .Y(_1179_),
    .A1(\pwm_module.counter1[18] ),
    .A2(_1097_));
 sg13g2_a21oi_1 _3500_ (.A1(\pwm_module.counter1[16] ),
    .A2(_1094_),
    .Y(_1180_),
    .B1(_1107_));
 sg13g2_nand2b_1 _3501_ (.Y(_1181_),
    .B(_1180_),
    .A_N(_1179_));
 sg13g2_nor4_2 _3502_ (.A(_1093_),
    .B(_1101_),
    .C(_1178_),
    .Y(_1182_),
    .D(_1181_));
 sg13g2_a21oi_1 _3503_ (.A1(_1084_),
    .A2(_1111_),
    .Y(_1183_),
    .B1(_1079_));
 sg13g2_nand2_1 _3504_ (.Y(_1184_),
    .A(_1084_),
    .B(_1182_));
 sg13g2_o21ai_1 _3505_ (.B1(_1183_),
    .Y(_1185_),
    .A1(_1177_),
    .A2(_1184_));
 sg13g2_o21ai_1 _3506_ (.B1(_1125_),
    .Y(_1186_),
    .A1(\pwm_module.counter1[0] ),
    .A2(_1128_));
 sg13g2_nand2b_1 _3507_ (.Y(_1187_),
    .B(_1129_),
    .A_N(_1127_));
 sg13g2_nor4_2 _3508_ (.A(_1124_),
    .B(_1176_),
    .C(_1186_),
    .Y(_1188_),
    .D(_1187_));
 sg13g2_nand4_1 _3509_ (.B(_1163_),
    .C(_1182_),
    .A(_1084_),
    .Y(_1189_),
    .D(_1188_));
 sg13g2_and3_1 _3510_ (.X(_0097_),
    .A(_2396_),
    .B(_1185_),
    .C(_1189_));
 sg13g2_a21oi_1 _3511_ (.A1(\MemCell.dc3_reg[3][7] ),
    .A2(net755),
    .Y(_1190_),
    .B1(_0168_));
 sg13g2_nand2_1 _3512_ (.Y(_1191_),
    .A(net755),
    .B(\MemCell.dc3_reg[3][6] ));
 sg13g2_a21oi_1 _3513_ (.A1(\pwm_module.counter2[30] ),
    .A2(_1191_),
    .Y(_1192_),
    .B1(_1190_));
 sg13g2_nor2b_1 _3514_ (.A(net768),
    .B_N(\MemCell.dc3_reg[3][5] ),
    .Y(_1193_));
 sg13g2_nand2_1 _3515_ (.Y(_1194_),
    .A(_0124_),
    .B(_1193_));
 sg13g2_o21ai_1 _3516_ (.B1(_1194_),
    .Y(_1195_),
    .A1(\pwm_module.counter2[30] ),
    .A2(_1191_));
 sg13g2_nand2b_1 _3517_ (.Y(_1196_),
    .B(\MemCell.dc3_reg[3][4] ),
    .A_N(net768));
 sg13g2_nor2_1 _3518_ (.A(_0124_),
    .B(_1193_),
    .Y(_1197_));
 sg13g2_a21oi_1 _3519_ (.A1(\pwm_module.counter2[28] ),
    .A2(_1196_),
    .Y(_1198_),
    .B1(_1197_));
 sg13g2_nor2_1 _3520_ (.A(\pwm_module.counter2[28] ),
    .B(_1196_),
    .Y(_1199_));
 sg13g2_nor2b_1 _3521_ (.A(net768),
    .B_N(\MemCell.dc3_reg[3][3] ),
    .Y(_1200_));
 sg13g2_a21oi_1 _3522_ (.A1(_0125_),
    .A2(_1200_),
    .Y(_1201_),
    .B1(_1199_));
 sg13g2_nor2_1 _3523_ (.A(_0125_),
    .B(_1200_),
    .Y(_1202_));
 sg13g2_nand2_1 _3524_ (.Y(_1203_),
    .A(net755),
    .B(\MemCell.dc3_reg[3][2] ));
 sg13g2_nor2_1 _3525_ (.A(\pwm_module.counter2[26] ),
    .B(_1203_),
    .Y(_1204_));
 sg13g2_nor2b_1 _3526_ (.A(net768),
    .B_N(\MemCell.dc3_reg[3][1] ),
    .Y(_1205_));
 sg13g2_nor2_1 _3527_ (.A(_0126_),
    .B(_1205_),
    .Y(_1206_));
 sg13g2_a21oi_1 _3528_ (.A1(\pwm_module.counter2[26] ),
    .A2(_1203_),
    .Y(_1207_),
    .B1(_1206_));
 sg13g2_nand2b_1 _3529_ (.Y(_1208_),
    .B(\MemCell.dc3_reg[3][0] ),
    .A_N(net768));
 sg13g2_nor2_1 _3530_ (.A(\pwm_module.counter2[24] ),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_a21oi_1 _3531_ (.A1(_0126_),
    .A2(_1205_),
    .Y(_1210_),
    .B1(_1209_));
 sg13g2_a21o_1 _3532_ (.A2(_1205_),
    .A1(_0126_),
    .B1(_1209_),
    .X(_1211_));
 sg13g2_a21oi_1 _3533_ (.A1(_1207_),
    .A2(_1211_),
    .Y(_1212_),
    .B1(_1204_));
 sg13g2_o21ai_1 _3534_ (.B1(_1201_),
    .Y(_1213_),
    .A1(_1202_),
    .A2(_1212_));
 sg13g2_a21oi_1 _3535_ (.A1(_1198_),
    .A2(_1213_),
    .Y(_1214_),
    .B1(_1195_));
 sg13g2_nand2b_1 _3536_ (.Y(_1215_),
    .B(_1192_),
    .A_N(_1214_));
 sg13g2_nand3_1 _3537_ (.B(\MemCell.dc3_reg[3][7] ),
    .C(net755),
    .A(_0168_),
    .Y(_1216_));
 sg13g2_nor2b_1 _3538_ (.A(net768),
    .B_N(\MemCell.dc3_reg[2][5] ),
    .Y(_1217_));
 sg13g2_xnor2_1 _3539_ (.Y(_1218_),
    .A(\pwm_module.counter2[21] ),
    .B(_1217_));
 sg13g2_nand2_1 _3540_ (.Y(_1219_),
    .A(net755),
    .B(\MemCell.dc3_reg[2][4] ));
 sg13g2_nand2_1 _3541_ (.Y(_1220_),
    .A(\pwm_module.counter2[20] ),
    .B(_1219_));
 sg13g2_nand2_1 _3542_ (.Y(_1221_),
    .A(net755),
    .B(\MemCell.dc3_reg[2][6] ));
 sg13g2_nand2_1 _3543_ (.Y(_1222_),
    .A(\pwm_module.counter2[22] ),
    .B(_1221_));
 sg13g2_nand3_1 _3544_ (.B(_1220_),
    .C(_1222_),
    .A(_1218_),
    .Y(_1223_));
 sg13g2_nand2b_1 _3545_ (.Y(_1224_),
    .B(\MemCell.dc3_reg[2][0] ),
    .A_N(net768));
 sg13g2_nor2_1 _3546_ (.A(\pwm_module.counter2[16] ),
    .B(_1224_),
    .Y(_1225_));
 sg13g2_nor2b_1 _3547_ (.A(net769),
    .B_N(\MemCell.dc3_reg[2][1] ),
    .Y(_1226_));
 sg13g2_a21oi_1 _3548_ (.A1(_0131_),
    .A2(_1226_),
    .Y(_1227_),
    .B1(_1225_));
 sg13g2_o21ai_1 _3549_ (.B1(\pwm_module.counter2[18] ),
    .Y(_1228_),
    .A1(net769),
    .A2(_2371_));
 sg13g2_nor3_1 _3550_ (.A(\pwm_module.counter2[18] ),
    .B(net769),
    .C(_2371_),
    .Y(_1229_));
 sg13g2_nor2b_1 _3551_ (.A(net769),
    .B_N(\MemCell.dc3_reg[2][3] ),
    .Y(_1230_));
 sg13g2_nor2_1 _3552_ (.A(_0131_),
    .B(_1226_),
    .Y(_1231_));
 sg13g2_o21ai_1 _3553_ (.B1(_1228_),
    .Y(_1232_),
    .A1(_0130_),
    .A2(_1230_));
 sg13g2_nor4_1 _3554_ (.A(_1227_),
    .B(_1229_),
    .C(_1231_),
    .D(_1232_),
    .Y(_1233_));
 sg13g2_nor2_1 _3555_ (.A(\pwm_module.counter2[20] ),
    .B(_1219_),
    .Y(_1234_));
 sg13g2_nand2_1 _3556_ (.Y(_1235_),
    .A(_0130_),
    .B(_1230_));
 sg13g2_nor2b_1 _3557_ (.A(_1234_),
    .B_N(_1235_),
    .Y(_1236_));
 sg13g2_o21ai_1 _3558_ (.B1(_1229_),
    .Y(_1237_),
    .A1(_0130_),
    .A2(_1230_));
 sg13g2_nand2_1 _3559_ (.Y(_1238_),
    .A(_1235_),
    .B(_1237_));
 sg13g2_nor3_1 _3560_ (.A(_1233_),
    .B(_1234_),
    .C(_1238_),
    .Y(_1239_));
 sg13g2_nor2b_1 _3561_ (.A(net768),
    .B_N(\MemCell.dc3_reg[2][7] ),
    .Y(_1240_));
 sg13g2_nor2_1 _3562_ (.A(\pwm_module.counter2[22] ),
    .B(_1221_),
    .Y(_1241_));
 sg13g2_a21oi_1 _3563_ (.A1(_0127_),
    .A2(_1240_),
    .Y(_1242_),
    .B1(_1241_));
 sg13g2_nand3_1 _3564_ (.B(_1217_),
    .C(_1222_),
    .A(_0128_),
    .Y(_1243_));
 sg13g2_and2_1 _3565_ (.A(_1242_),
    .B(_1243_),
    .X(_1244_));
 sg13g2_o21ai_1 _3566_ (.B1(_1244_),
    .Y(_1245_),
    .A1(_1223_),
    .A2(_1239_));
 sg13g2_or2_1 _3567_ (.X(_1246_),
    .B(_1240_),
    .A(_0127_));
 sg13g2_nand2_1 _3568_ (.Y(_1247_),
    .A(\pwm_module.counter2[24] ),
    .B(_1208_));
 sg13g2_and4_1 _3569_ (.A(_1198_),
    .B(_1201_),
    .C(_1207_),
    .D(_1210_),
    .X(_1248_));
 sg13g2_nand4_1 _3570_ (.B(_1216_),
    .C(_1247_),
    .A(_1192_),
    .Y(_1249_),
    .D(_1248_));
 sg13g2_nor4_2 _3571_ (.A(_1195_),
    .B(_1202_),
    .C(_1204_),
    .Y(_1250_),
    .D(_1249_));
 sg13g2_nand3_1 _3572_ (.B(_1246_),
    .C(_1250_),
    .A(_1245_),
    .Y(_1251_));
 sg13g2_nand3_1 _3573_ (.B(_1216_),
    .C(_1251_),
    .A(_1215_),
    .Y(_1252_));
 sg13g2_nand3_1 _3574_ (.B(net756),
    .C(\MemCell.dc3_reg[0][7] ),
    .A(_0138_),
    .Y(_1253_));
 sg13g2_nor2_1 _3575_ (.A(net771),
    .B(\MemCell.dc3_reg[0][6] ),
    .Y(_1254_));
 sg13g2_o21ai_1 _3576_ (.B1(_1253_),
    .Y(_1255_),
    .A1(\pwm_module.counter2[6] ),
    .A2(_1254_));
 sg13g2_xnor2_1 _3577_ (.Y(_1256_),
    .A(_0139_),
    .B(_1254_));
 sg13g2_nor2_1 _3578_ (.A(net770),
    .B(\MemCell.dc3_reg[0][5] ),
    .Y(_1257_));
 sg13g2_or2_1 _3579_ (.X(_1258_),
    .B(_1257_),
    .A(\pwm_module.counter2[5] ));
 sg13g2_xor2_1 _3580_ (.B(_1257_),
    .A(_0140_),
    .X(_1259_));
 sg13g2_o21ai_1 _3581_ (.B1(_0141_),
    .Y(_1260_),
    .A1(net770),
    .A2(\MemCell.dc3_reg[0][4] ));
 sg13g2_inv_1 _3582_ (.Y(_1261_),
    .A(_1260_));
 sg13g2_nor2b_1 _3583_ (.A(net770),
    .B_N(\MemCell.dc3_reg[0][3] ),
    .Y(_1262_));
 sg13g2_nor2_1 _3584_ (.A(_0142_),
    .B(_1262_),
    .Y(_1263_));
 sg13g2_nor3_1 _3585_ (.A(net770),
    .B(\MemCell.dc3_reg[0][4] ),
    .C(_0141_),
    .Y(_1264_));
 sg13g2_nor2b_1 _3586_ (.A(net770),
    .B_N(\MemCell.dc3_reg[0][2] ),
    .Y(_1265_));
 sg13g2_nand2_1 _3587_ (.Y(_1266_),
    .A(net756),
    .B(\MemCell.dc3_reg[0][2] ));
 sg13g2_a22oi_1 _3588_ (.Y(_1267_),
    .B1(_1265_),
    .B2(_2318_),
    .A2(_1262_),
    .A1(_0142_));
 sg13g2_nor2_1 _3589_ (.A(_2318_),
    .B(_1265_),
    .Y(_1268_));
 sg13g2_nor2b_1 _3590_ (.A(net770),
    .B_N(\MemCell.dc3_reg[0][1] ),
    .Y(_1269_));
 sg13g2_nor2_1 _3591_ (.A(net770),
    .B(\MemCell.dc3_reg[0][0] ),
    .Y(_1270_));
 sg13g2_nand2_1 _3592_ (.Y(_1271_),
    .A(\pwm_module.counter2[0] ),
    .B(_1270_));
 sg13g2_o21ai_1 _3593_ (.B1(_1271_),
    .Y(_1272_),
    .A1(_0143_),
    .A2(_1269_));
 sg13g2_nand2_1 _3594_ (.Y(_1273_),
    .A(_0143_),
    .B(_1269_));
 sg13g2_a21o_1 _3595_ (.A2(\MemCell.dc3_reg[0][7] ),
    .A1(net756),
    .B1(_0138_),
    .X(_1274_));
 sg13g2_nor2b_1 _3596_ (.A(net771),
    .B_N(\MemCell.dc3_reg[1][2] ),
    .Y(_1275_));
 sg13g2_xnor2_1 _3597_ (.Y(_1276_),
    .A(\pwm_module.counter2[10] ),
    .B(_1275_));
 sg13g2_nor2_1 _3598_ (.A(net771),
    .B(\MemCell.dc3_reg[1][1] ),
    .Y(_1277_));
 sg13g2_xnor2_1 _3599_ (.Y(_1278_),
    .A(_0137_),
    .B(_1277_));
 sg13g2_nand2_1 _3600_ (.Y(_1279_),
    .A(net755),
    .B(\MemCell.dc3_reg[1][4] ));
 sg13g2_or2_1 _3601_ (.X(_1280_),
    .B(_1279_),
    .A(\pwm_module.counter2[12] ));
 sg13g2_nor2b_1 _3602_ (.A(net771),
    .B_N(\MemCell.dc3_reg[1][7] ),
    .Y(_1281_));
 sg13g2_nand2_1 _3603_ (.Y(_1282_),
    .A(_0132_),
    .B(_1281_));
 sg13g2_nand2_1 _3604_ (.Y(_1283_),
    .A(net755),
    .B(\MemCell.dc3_reg[1][6] ));
 sg13g2_nand2_1 _3605_ (.Y(_1284_),
    .A(\pwm_module.counter2[14] ),
    .B(_1283_));
 sg13g2_nor2_1 _3606_ (.A(\pwm_module.counter2[14] ),
    .B(_1283_),
    .Y(_1285_));
 sg13g2_o21ai_1 _3607_ (.B1(_1284_),
    .Y(_1286_),
    .A1(_0132_),
    .A2(_1281_));
 sg13g2_nor2_1 _3608_ (.A(_1285_),
    .B(_1286_),
    .Y(_1287_));
 sg13g2_nor2b_1 _3609_ (.A(net771),
    .B_N(\MemCell.dc3_reg[1][5] ),
    .Y(_1288_));
 sg13g2_a22oi_1 _3610_ (.Y(_1289_),
    .B1(_1288_),
    .B2(_2322_),
    .A2(_1279_),
    .A1(\pwm_module.counter2[12] ));
 sg13g2_o21ai_1 _3611_ (.B1(_1289_),
    .Y(_1290_),
    .A1(_2322_),
    .A2(_1288_));
 sg13g2_nand3_1 _3612_ (.B(net756),
    .C(\MemCell.dc3_reg[1][3] ),
    .A(_0135_),
    .Y(_1291_));
 sg13g2_nor3_1 _3613_ (.A(\pwm_module.counter2[8] ),
    .B(net771),
    .C(_2372_),
    .Y(_1292_));
 sg13g2_a21oi_1 _3614_ (.A1(net756),
    .A2(\MemCell.dc3_reg[1][3] ),
    .Y(_1293_),
    .B1(_0135_));
 sg13g2_o21ai_1 _3615_ (.B1(\pwm_module.counter2[8] ),
    .Y(_1294_),
    .A1(net771),
    .A2(_2372_));
 sg13g2_and2_1 _3616_ (.A(_0133_),
    .B(_1288_),
    .X(_1295_));
 sg13g2_and2_1 _3617_ (.A(_1280_),
    .B(_1291_),
    .X(_1296_));
 sg13g2_nor2_1 _3618_ (.A(\pwm_module.counter2[9] ),
    .B(_1277_),
    .Y(_1297_));
 sg13g2_a21o_1 _3619_ (.A2(_1292_),
    .A1(_1278_),
    .B1(_1297_),
    .X(_1298_));
 sg13g2_a22oi_1 _3620_ (.Y(_1299_),
    .B1(_1276_),
    .B2(_1298_),
    .A2(_1275_),
    .A1(_0136_));
 sg13g2_or2_1 _3621_ (.X(_1300_),
    .B(_1299_),
    .A(_1293_));
 sg13g2_nand3b_1 _3622_ (.B(_1276_),
    .C(_1291_),
    .Y(_1301_),
    .A_N(_1293_));
 sg13g2_a21oi_1 _3623_ (.A1(_1296_),
    .A2(_1300_),
    .Y(_1302_),
    .B1(_1290_));
 sg13g2_o21ai_1 _3624_ (.B1(_1287_),
    .Y(_1303_),
    .A1(_1295_),
    .A2(_1302_));
 sg13g2_o21ai_1 _3625_ (.B1(_1285_),
    .Y(_1304_),
    .A1(_0132_),
    .A2(_1281_));
 sg13g2_nor2_1 _3626_ (.A(_1290_),
    .B(_1301_),
    .Y(_1305_));
 sg13g2_nor2b_1 _3627_ (.A(_1292_),
    .B_N(_1294_),
    .Y(_1306_));
 sg13g2_and4_1 _3628_ (.A(_1278_),
    .B(_1280_),
    .C(_1282_),
    .D(_1306_),
    .X(_1307_));
 sg13g2_nand2_1 _3629_ (.Y(_1308_),
    .A(_1255_),
    .B(_1274_));
 sg13g2_nand3_1 _3630_ (.B(_1256_),
    .C(_1274_),
    .A(_1253_),
    .Y(_1309_));
 sg13g2_nor4_2 _3631_ (.A(_1259_),
    .B(_1261_),
    .C(_1264_),
    .Y(_1310_),
    .D(_1309_));
 sg13g2_nand2b_1 _3632_ (.Y(_1311_),
    .B(_1267_),
    .A_N(_1263_));
 sg13g2_a221oi_1 _3633_ (.B2(_1273_),
    .C1(_1311_),
    .B1(_1272_),
    .A1(\pwm_module.counter2[2] ),
    .Y(_1312_),
    .A2(_1266_));
 sg13g2_nor2_1 _3634_ (.A(_1263_),
    .B(_1267_),
    .Y(_1313_));
 sg13g2_o21ai_1 _3635_ (.B1(_1310_),
    .Y(_1314_),
    .A1(_1312_),
    .A2(_1313_));
 sg13g2_o21ai_1 _3636_ (.B1(_1258_),
    .Y(_1315_),
    .A1(_1259_),
    .A2(_1260_));
 sg13g2_nand2b_1 _3637_ (.Y(_1316_),
    .B(_1315_),
    .A_N(_1309_));
 sg13g2_nand3_1 _3638_ (.B(_1314_),
    .C(_1316_),
    .A(_1308_),
    .Y(_1317_));
 sg13g2_nand4_1 _3639_ (.B(_1305_),
    .C(_1307_),
    .A(_1287_),
    .Y(_1318_),
    .D(_1317_));
 sg13g2_nand4_1 _3640_ (.B(_1303_),
    .C(_1304_),
    .A(_1282_),
    .Y(_1319_),
    .D(_1318_));
 sg13g2_nand2_1 _3641_ (.Y(_1320_),
    .A(\pwm_module.counter2[16] ),
    .B(_1224_));
 sg13g2_and2_1 _3642_ (.A(_1246_),
    .B(_1320_),
    .X(_1321_));
 sg13g2_and4_1 _3643_ (.A(_1227_),
    .B(_1236_),
    .C(_1242_),
    .D(_1321_),
    .X(_1322_));
 sg13g2_nor4_1 _3644_ (.A(_1223_),
    .B(_1229_),
    .C(_1231_),
    .D(_1232_),
    .Y(_1323_));
 sg13g2_and3_1 _3645_ (.X(_1324_),
    .A(_1250_),
    .B(_1322_),
    .C(_1323_));
 sg13g2_a21oi_1 _3646_ (.A1(_1319_),
    .A2(_1324_),
    .Y(_1325_),
    .B1(_1252_));
 sg13g2_or2_1 _3647_ (.X(_1326_),
    .B(_1270_),
    .A(\pwm_module.counter2[0] ));
 sg13g2_nor3_1 _3648_ (.A(_1268_),
    .B(_1272_),
    .C(_1311_),
    .Y(_1327_));
 sg13g2_nand4_1 _3649_ (.B(_1310_),
    .C(_1326_),
    .A(_1273_),
    .Y(_1328_),
    .D(_1327_));
 sg13g2_nand4_1 _3650_ (.B(_1305_),
    .C(_1307_),
    .A(_1287_),
    .Y(_1329_),
    .D(_1324_));
 sg13g2_nor2_1 _3651_ (.A(_1328_),
    .B(_1329_),
    .Y(_1330_));
 sg13g2_nor3_2 _3652_ (.A(_2395_),
    .B(_1325_),
    .C(_1330_),
    .Y(_0098_));
 sg13g2_xor2_1 _3653_ (.B(\spi_module.r_RX_Bit_Count[0] ),
    .A(\spi_module.r_RX_Bit_Count[1] ),
    .X(_0100_));
 sg13g2_a21o_1 _3654_ (.A2(\spi_module.r_RX_Bit_Count[0] ),
    .A1(\spi_module.r_RX_Bit_Count[1] ),
    .B1(\spi_module.r_RX_Bit_Count[2] ),
    .X(_1331_));
 sg13g2_and2_1 _3655_ (.A(_2393_),
    .B(_1331_),
    .X(_0101_));
 sg13g2_nor4_1 _3656_ (.A(\MemCell.counter_value[21] ),
    .B(\MemCell.counter_value[20] ),
    .C(\MemCell.counter_value[23] ),
    .D(\MemCell.counter_value[22] ),
    .Y(_1332_));
 sg13g2_nor4_1 _3657_ (.A(\MemCell.counter_value[17] ),
    .B(\MemCell.counter_value[16] ),
    .C(\MemCell.counter_value[19] ),
    .D(\MemCell.counter_value[18] ),
    .Y(_1333_));
 sg13g2_nor4_2 _3658_ (.A(\MemCell.counter_value[25] ),
    .B(\MemCell.counter_value[24] ),
    .C(\MemCell.counter_value[27] ),
    .Y(_1334_),
    .D(\MemCell.counter_value[26] ));
 sg13g2_nor4_1 _3659_ (.A(\MemCell.counter_value[29] ),
    .B(\MemCell.counter_value[28] ),
    .C(\MemCell.counter_value[31] ),
    .D(\MemCell.counter_value[30] ),
    .Y(_1335_));
 sg13g2_and3_1 _3660_ (.X(_1336_),
    .A(_1332_),
    .B(_1333_),
    .C(_1335_));
 sg13g2_nor4_1 _3661_ (.A(\MemCell.counter_value[5] ),
    .B(\MemCell.counter_value[4] ),
    .C(\MemCell.counter_value[7] ),
    .D(\MemCell.counter_value[6] ),
    .Y(_1337_));
 sg13g2_nor4_1 _3662_ (.A(\MemCell.counter_value[1] ),
    .B(\MemCell.counter_value[0] ),
    .C(\MemCell.counter_value[3] ),
    .D(\MemCell.counter_value[2] ),
    .Y(_1338_));
 sg13g2_nor4_1 _3663_ (.A(\MemCell.counter_value[9] ),
    .B(\MemCell.counter_value[8] ),
    .C(\MemCell.counter_value[11] ),
    .D(\MemCell.counter_value[10] ),
    .Y(_1339_));
 sg13g2_nor4_1 _3664_ (.A(\MemCell.counter_value[13] ),
    .B(\MemCell.counter_value[12] ),
    .C(\MemCell.counter_value[15] ),
    .D(\MemCell.counter_value[14] ),
    .Y(_1340_));
 sg13g2_and3_2 _3665_ (.X(_1341_),
    .A(_1337_),
    .B(_1338_),
    .C(_1340_));
 sg13g2_nand4_1 _3666_ (.B(_1336_),
    .C(_1339_),
    .A(_1334_),
    .Y(uo_out[3]),
    .D(_1341_));
 sg13g2_nor4_1 _3667_ (.A(\MemCell.prescale_reg[3][3] ),
    .B(\MemCell.prescale_reg[3][2] ),
    .C(\MemCell.prescale_reg[3][1] ),
    .D(\MemCell.prescale_reg[3][0] ),
    .Y(_1342_));
 sg13g2_nor4_1 _3668_ (.A(\MemCell.prescale_reg[3][7] ),
    .B(\MemCell.prescale_reg[3][6] ),
    .C(\MemCell.prescale_reg[3][5] ),
    .D(\MemCell.prescale_reg[3][4] ),
    .Y(_1343_));
 sg13g2_and2_1 _3669_ (.A(_1342_),
    .B(_1343_),
    .X(_1344_));
 sg13g2_nor4_1 _3670_ (.A(\MemCell.prescale_reg[2][7] ),
    .B(\MemCell.prescale_reg[2][6] ),
    .C(\MemCell.prescale_reg[2][5] ),
    .D(\MemCell.prescale_reg[2][4] ),
    .Y(_1345_));
 sg13g2_nor4_1 _3671_ (.A(\MemCell.prescale_reg[2][3] ),
    .B(\MemCell.prescale_reg[2][2] ),
    .C(\MemCell.prescale_reg[2][1] ),
    .D(\MemCell.prescale_reg[2][0] ),
    .Y(_1346_));
 sg13g2_nor4_1 _3672_ (.A(\MemCell.prescale_reg[0][7] ),
    .B(\MemCell.prescale_reg[0][6] ),
    .C(\MemCell.prescale_reg[0][5] ),
    .D(\MemCell.prescale_reg[0][4] ),
    .Y(_1347_));
 sg13g2_nor4_2 _3673_ (.A(\MemCell.prescale_reg[0][0] ),
    .B(\MemCell.prescale_reg[0][1] ),
    .C(\MemCell.prescale_reg[0][3] ),
    .Y(_1348_),
    .D(\MemCell.prescale_reg[0][2] ));
 sg13g2_or2_1 _3674_ (.X(_1349_),
    .B(\MemCell.prescale_reg[1][6] ),
    .A(\MemCell.prescale_reg[1][7] ));
 sg13g2_nor4_1 _3675_ (.A(\MemCell.prescale_reg[1][3] ),
    .B(\MemCell.prescale_reg[1][2] ),
    .C(\MemCell.prescale_reg[1][1] ),
    .D(\MemCell.prescale_reg[1][0] ),
    .Y(_1350_));
 sg13g2_nand3_1 _3676_ (.B(_1348_),
    .C(_1350_),
    .A(_1347_),
    .Y(_1351_));
 sg13g2_nor4_2 _3677_ (.A(\MemCell.prescale_reg[1][5] ),
    .B(\MemCell.prescale_reg[1][4] ),
    .C(_1349_),
    .Y(_1352_),
    .D(_1351_));
 sg13g2_nand4_1 _3678_ (.B(_1345_),
    .C(_1346_),
    .A(_1344_),
    .Y(uo_out[4]),
    .D(_1352_));
 sg13g2_nor4_1 _3679_ (.A(\MemCell.dc1_reg[1][3] ),
    .B(\MemCell.dc1_reg[1][2] ),
    .C(\MemCell.dc1_reg[1][1] ),
    .D(\MemCell.dc1_reg[1][0] ),
    .Y(_1353_));
 sg13g2_nor4_1 _3680_ (.A(\MemCell.dc1_reg[1][7] ),
    .B(\MemCell.dc1_reg[1][6] ),
    .C(\MemCell.dc1_reg[1][5] ),
    .D(\MemCell.dc1_reg[1][4] ),
    .Y(_1354_));
 sg13g2_nor4_1 _3681_ (.A(\MemCell.dc1_reg[0][7] ),
    .B(\MemCell.dc1_reg[0][6] ),
    .C(\MemCell.dc1_reg[0][5] ),
    .D(\MemCell.dc1_reg[0][4] ),
    .Y(_1355_));
 sg13g2_nor4_1 _3682_ (.A(\MemCell.dc1_reg[0][3] ),
    .B(\MemCell.dc1_reg[0][2] ),
    .C(\MemCell.dc1_reg[0][1] ),
    .D(\MemCell.dc1_reg[0][0] ),
    .Y(_1356_));
 sg13g2_and3_1 _3683_ (.X(_1357_),
    .A(_1353_),
    .B(_1354_),
    .C(_1356_));
 sg13g2_nor4_1 _3684_ (.A(\MemCell.dc1_reg[3][3] ),
    .B(\MemCell.dc1_reg[3][2] ),
    .C(\MemCell.dc1_reg[3][1] ),
    .D(\MemCell.dc1_reg[3][0] ),
    .Y(_1358_));
 sg13g2_nor4_1 _3685_ (.A(\MemCell.dc1_reg[3][7] ),
    .B(\MemCell.dc1_reg[3][6] ),
    .C(\MemCell.dc1_reg[3][5] ),
    .D(\MemCell.dc1_reg[3][4] ),
    .Y(_1359_));
 sg13g2_nor4_1 _3686_ (.A(\MemCell.dc1_reg[2][7] ),
    .B(\MemCell.dc1_reg[2][6] ),
    .C(\MemCell.dc1_reg[2][5] ),
    .D(\MemCell.dc1_reg[2][4] ),
    .Y(_1360_));
 sg13g2_nor4_1 _3687_ (.A(\MemCell.dc1_reg[2][3] ),
    .B(\MemCell.dc1_reg[2][2] ),
    .C(\MemCell.dc1_reg[2][1] ),
    .D(\MemCell.dc1_reg[2][0] ),
    .Y(_1361_));
 sg13g2_and3_1 _3688_ (.X(_1362_),
    .A(_1358_),
    .B(_1359_),
    .C(_1361_));
 sg13g2_nand4_1 _3689_ (.B(_1357_),
    .C(_1360_),
    .A(_1355_),
    .Y(uo_out[5]),
    .D(_1362_));
 sg13g2_nor4_1 _3690_ (.A(\MemCell.dc2_reg[1][3] ),
    .B(\MemCell.dc2_reg[1][2] ),
    .C(\MemCell.dc2_reg[1][1] ),
    .D(\MemCell.dc2_reg[1][0] ),
    .Y(_1363_));
 sg13g2_nor4_1 _3691_ (.A(\MemCell.dc2_reg[1][7] ),
    .B(\MemCell.dc2_reg[1][6] ),
    .C(\MemCell.dc2_reg[1][5] ),
    .D(\MemCell.dc2_reg[1][4] ),
    .Y(_1364_));
 sg13g2_nor4_2 _3692_ (.A(\MemCell.dc2_reg[0][7] ),
    .B(\MemCell.dc2_reg[0][6] ),
    .C(\MemCell.dc2_reg[0][5] ),
    .Y(_1365_),
    .D(\MemCell.dc2_reg[0][4] ));
 sg13g2_nor4_2 _3693_ (.A(\MemCell.dc2_reg[0][3] ),
    .B(\MemCell.dc2_reg[0][2] ),
    .C(\MemCell.dc2_reg[0][1] ),
    .Y(_1366_),
    .D(\MemCell.dc2_reg[0][0] ));
 sg13g2_and3_1 _3694_ (.X(_1367_),
    .A(_1363_),
    .B(_1364_),
    .C(_1366_));
 sg13g2_nor4_2 _3695_ (.A(\MemCell.dc2_reg[3][3] ),
    .B(\MemCell.dc2_reg[3][2] ),
    .C(\MemCell.dc2_reg[3][1] ),
    .Y(_1368_),
    .D(\MemCell.dc2_reg[3][0] ));
 sg13g2_nor4_1 _3696_ (.A(\MemCell.dc2_reg[3][7] ),
    .B(\MemCell.dc2_reg[3][6] ),
    .C(\MemCell.dc2_reg[3][5] ),
    .D(\MemCell.dc2_reg[3][4] ),
    .Y(_1369_));
 sg13g2_nor4_1 _3697_ (.A(\MemCell.dc2_reg[2][7] ),
    .B(\MemCell.dc2_reg[2][6] ),
    .C(\MemCell.dc2_reg[2][5] ),
    .D(\MemCell.dc2_reg[2][4] ),
    .Y(_1370_));
 sg13g2_nor4_1 _3698_ (.A(\MemCell.dc2_reg[2][3] ),
    .B(\MemCell.dc2_reg[2][2] ),
    .C(\MemCell.dc2_reg[2][1] ),
    .D(\MemCell.dc2_reg[2][0] ),
    .Y(_1371_));
 sg13g2_and3_1 _3699_ (.X(_1372_),
    .A(_1368_),
    .B(_1369_),
    .C(_1371_));
 sg13g2_nand4_1 _3700_ (.B(_1367_),
    .C(_1370_),
    .A(_1365_),
    .Y(uo_out[6]),
    .D(_1372_));
 sg13g2_nor4_1 _3701_ (.A(\MemCell.dc3_reg[1][3] ),
    .B(\MemCell.dc3_reg[1][2] ),
    .C(\MemCell.dc3_reg[1][1] ),
    .D(\MemCell.dc3_reg[1][0] ),
    .Y(_1373_));
 sg13g2_nor4_1 _3702_ (.A(\MemCell.dc3_reg[1][7] ),
    .B(\MemCell.dc3_reg[1][6] ),
    .C(\MemCell.dc3_reg[1][5] ),
    .D(\MemCell.dc3_reg[1][4] ),
    .Y(_1374_));
 sg13g2_nor4_2 _3703_ (.A(\MemCell.dc3_reg[0][7] ),
    .B(\MemCell.dc3_reg[0][6] ),
    .C(\MemCell.dc3_reg[0][5] ),
    .Y(_1375_),
    .D(\MemCell.dc3_reg[0][4] ));
 sg13g2_nor4_2 _3704_ (.A(\MemCell.dc3_reg[0][3] ),
    .B(\MemCell.dc3_reg[0][2] ),
    .C(\MemCell.dc3_reg[0][1] ),
    .Y(_1376_),
    .D(\MemCell.dc3_reg[0][0] ));
 sg13g2_and3_1 _3705_ (.X(_1377_),
    .A(_1373_),
    .B(_1374_),
    .C(_1376_));
 sg13g2_nor4_1 _3706_ (.A(\MemCell.dc3_reg[3][3] ),
    .B(\MemCell.dc3_reg[3][2] ),
    .C(\MemCell.dc3_reg[3][1] ),
    .D(\MemCell.dc3_reg[3][0] ),
    .Y(_1378_));
 sg13g2_nor4_1 _3707_ (.A(\MemCell.dc3_reg[3][7] ),
    .B(\MemCell.dc3_reg[3][6] ),
    .C(\MemCell.dc3_reg[3][5] ),
    .D(\MemCell.dc3_reg[3][4] ),
    .Y(_1379_));
 sg13g2_nor4_1 _3708_ (.A(\MemCell.dc3_reg[2][7] ),
    .B(\MemCell.dc3_reg[2][6] ),
    .C(\MemCell.dc3_reg[2][5] ),
    .D(\MemCell.dc3_reg[2][4] ),
    .Y(_1380_));
 sg13g2_nor4_1 _3709_ (.A(\MemCell.dc3_reg[2][3] ),
    .B(\MemCell.dc3_reg[2][2] ),
    .C(\MemCell.dc3_reg[2][1] ),
    .D(\MemCell.dc3_reg[2][0] ),
    .Y(_1381_));
 sg13g2_and3_1 _3710_ (.X(_1382_),
    .A(_1378_),
    .B(_1379_),
    .C(_1381_));
 sg13g2_nand4_1 _3711_ (.B(_1377_),
    .C(_1380_),
    .A(_1375_),
    .Y(uo_out[7]),
    .D(_1382_));
 sg13g2_nor2b_2 _3712_ (.A(net375),
    .B_N(net35),
    .Y(_0099_));
 sg13g2_nand2_1 _3713_ (.Y(_1383_),
    .A(_0214_),
    .B(_0543_));
 sg13g2_a22oi_1 _3714_ (.Y(_1384_),
    .B1(_0543_),
    .B2(_0214_),
    .A2(_0541_),
    .A1(_2386_));
 sg13g2_o21ai_1 _3715_ (.B1(_1383_),
    .Y(_1385_),
    .A1(\pwm_module.prescaler0[22] ),
    .A2(_0542_));
 sg13g2_nand2_1 _3716_ (.Y(_1386_),
    .A(\pwm_module.prescaler0[22] ),
    .B(_0542_));
 sg13g2_nand2b_1 _3717_ (.Y(_1387_),
    .B(_0547_),
    .A_N(_0213_));
 sg13g2_a22oi_1 _3718_ (.Y(_1388_),
    .B1(_0550_),
    .B2(_0212_),
    .A2(_0546_),
    .A1(_0213_));
 sg13g2_and2_1 _3719_ (.A(_0211_),
    .B(_0556_),
    .X(_1389_));
 sg13g2_nor2_1 _3720_ (.A(_0211_),
    .B(_0556_),
    .Y(_1390_));
 sg13g2_nand2b_1 _3721_ (.Y(_1391_),
    .B(_0557_),
    .A_N(_0211_));
 sg13g2_and2_1 _3722_ (.A(\pwm_module.prescaler0[18] ),
    .B(_0559_),
    .X(_1392_));
 sg13g2_nor2_1 _3723_ (.A(\pwm_module.prescaler0[18] ),
    .B(_0559_),
    .Y(_1393_));
 sg13g2_or4_1 _3724_ (.A(_1389_),
    .B(_1390_),
    .C(_1392_),
    .D(_1393_),
    .X(_1394_));
 sg13g2_and2_1 _3725_ (.A(_0210_),
    .B(_0561_),
    .X(_1395_));
 sg13g2_nand2b_1 _3726_ (.Y(_1396_),
    .B(_0562_),
    .A_N(_0210_));
 sg13g2_nor2_1 _3727_ (.A(\pwm_module.prescaler0[16] ),
    .B(_0565_),
    .Y(_1397_));
 sg13g2_a21oi_1 _3728_ (.A1(_1396_),
    .A2(_1397_),
    .Y(_1398_),
    .B1(_1395_));
 sg13g2_a21oi_1 _3729_ (.A1(_1391_),
    .A2(_1393_),
    .Y(_1399_),
    .B1(_1389_));
 sg13g2_o21ai_1 _3730_ (.B1(_1399_),
    .Y(_1400_),
    .A1(_1394_),
    .A2(_1398_));
 sg13g2_or2_1 _3731_ (.X(_1401_),
    .B(_0543_),
    .A(_0214_));
 sg13g2_nor2_1 _3732_ (.A(_0218_),
    .B(_0508_),
    .Y(_1402_));
 sg13g2_a21oi_1 _3733_ (.A1(\pwm_module.prescaler0[28] ),
    .A2(_0514_),
    .Y(_1403_),
    .B1(_1402_));
 sg13g2_inv_1 _3734_ (.Y(_1404_),
    .A(_1403_));
 sg13g2_nand2_1 _3735_ (.Y(_1405_),
    .A(_0215_),
    .B(_0519_));
 sg13g2_a22oi_1 _3736_ (.Y(_1406_),
    .B1(_0527_),
    .B2(_0217_),
    .A2(_0519_),
    .A1(_0215_));
 sg13g2_nand2_1 _3737_ (.Y(_1407_),
    .A(_0218_),
    .B(_0508_));
 sg13g2_nand2_1 _3738_ (.Y(_1408_),
    .A(\pwm_module.prescaler0[24] ),
    .B(_0518_));
 sg13g2_nand4_1 _3739_ (.B(_1406_),
    .C(_1407_),
    .A(_1403_),
    .Y(_1409_),
    .D(_1408_));
 sg13g2_a22oi_1 _3740_ (.Y(_1410_),
    .B1(_0528_),
    .B2(_2385_),
    .A2(_0523_),
    .A1(_0216_));
 sg13g2_o21ai_1 _3741_ (.B1(_1410_),
    .Y(_1411_),
    .A1(_0216_),
    .A2(_0523_));
 sg13g2_nor2_1 _3742_ (.A(\pwm_module.prescaler0[30] ),
    .B(_0506_),
    .Y(_1412_));
 sg13g2_xor2_1 _3743_ (.B(_0506_),
    .A(\pwm_module.prescaler0[30] ),
    .X(_1413_));
 sg13g2_o21ai_1 _3744_ (.B1(_1413_),
    .Y(_1414_),
    .A1(_0102_),
    .A2(_0510_));
 sg13g2_inv_1 _3745_ (.Y(_1415_),
    .A(_1414_));
 sg13g2_nor2_1 _3746_ (.A(\pwm_module.prescaler0[28] ),
    .B(_0514_),
    .Y(_1416_));
 sg13g2_a21oi_1 _3747_ (.A1(_0102_),
    .A2(_0510_),
    .Y(_1417_),
    .B1(_1416_));
 sg13g2_nand2b_1 _3748_ (.Y(_1418_),
    .B(_0520_),
    .A_N(_0215_));
 sg13g2_nor2_1 _3749_ (.A(\pwm_module.prescaler0[24] ),
    .B(_0518_),
    .Y(_1419_));
 sg13g2_nand3b_1 _3750_ (.B(_1417_),
    .C(_1418_),
    .Y(_1420_),
    .A_N(_1419_));
 sg13g2_nor4_2 _3751_ (.A(_1409_),
    .B(_1411_),
    .C(_1414_),
    .Y(_1421_),
    .D(_1420_));
 sg13g2_nand2_1 _3752_ (.Y(_1422_),
    .A(_1418_),
    .B(_1419_));
 sg13g2_a21oi_1 _3753_ (.A1(_1405_),
    .A2(_1422_),
    .Y(_1423_),
    .B1(_1411_));
 sg13g2_a22oi_1 _3754_ (.Y(_1424_),
    .B1(_0527_),
    .B2(_0217_),
    .A2(_0523_),
    .A1(_0216_));
 sg13g2_a21oi_1 _3755_ (.A1(_2385_),
    .A2(_0528_),
    .Y(_1425_),
    .B1(_1424_));
 sg13g2_nor3_1 _3756_ (.A(_1416_),
    .B(_1423_),
    .C(_1425_),
    .Y(_1426_));
 sg13g2_o21ai_1 _3757_ (.B1(_1407_),
    .Y(_1427_),
    .A1(_1404_),
    .A2(_1426_));
 sg13g2_o21ai_1 _3758_ (.B1(_1412_),
    .Y(_1428_),
    .A1(_0102_),
    .A2(net719));
 sg13g2_nand4_1 _3759_ (.B(_1386_),
    .C(_1387_),
    .A(_1384_),
    .Y(_1429_),
    .D(_1401_));
 sg13g2_nor2_1 _3760_ (.A(_1388_),
    .B(_1429_),
    .Y(_1430_));
 sg13g2_o21ai_1 _3761_ (.B1(_1388_),
    .Y(_1431_),
    .A1(_0212_),
    .A2(_0550_));
 sg13g2_nor2_1 _3762_ (.A(_1429_),
    .B(_1431_),
    .Y(_1432_));
 sg13g2_a221oi_1 _3763_ (.B2(_1400_),
    .C1(_1430_),
    .B1(_1432_),
    .A1(_1385_),
    .Y(_1433_),
    .A2(_1401_));
 sg13g2_nand4_1 _3764_ (.B(_1407_),
    .C(_1417_),
    .A(_1403_),
    .Y(_1434_),
    .D(_1418_));
 sg13g2_nand3b_1 _3765_ (.B(_1406_),
    .C(_1408_),
    .Y(_1435_),
    .A_N(_1419_));
 sg13g2_or4_1 _3766_ (.A(_1411_),
    .B(_1414_),
    .C(_1434_),
    .D(_1435_),
    .X(_1436_));
 sg13g2_o21ai_1 _3767_ (.B1(_1428_),
    .Y(_1437_),
    .A1(_1433_),
    .A2(_1436_));
 sg13g2_a221oi_1 _3768_ (.B2(_1427_),
    .C1(_1437_),
    .B1(_1415_),
    .A1(_0102_),
    .Y(_1438_),
    .A2(net719));
 sg13g2_or2_1 _3769_ (.X(_1439_),
    .B(_0613_),
    .A(_0209_));
 sg13g2_o21ai_1 _3770_ (.B1(_1439_),
    .Y(_1440_),
    .A1(_0208_),
    .A2(_0617_));
 sg13g2_a21o_1 _3771_ (.A2(_0612_),
    .A1(\pwm_module.prescaler0[14] ),
    .B1(_1440_),
    .X(_1441_));
 sg13g2_nand2_1 _3772_ (.Y(_1442_),
    .A(_0208_),
    .B(_0617_));
 sg13g2_nand2b_1 _3773_ (.Y(_1443_),
    .B(_0620_),
    .A_N(\pwm_module.prescaler0[12] ));
 sg13g2_and2_1 _3774_ (.A(_1442_),
    .B(_1443_),
    .X(_1444_));
 sg13g2_nand2_1 _3775_ (.Y(_1445_),
    .A(_1442_),
    .B(_1443_));
 sg13g2_nand2b_1 _3776_ (.Y(_1446_),
    .B(\pwm_module.prescaler0[12] ),
    .A_N(_0620_));
 sg13g2_nand2_1 _3777_ (.Y(_1447_),
    .A(_0207_),
    .B(_0629_));
 sg13g2_a22oi_1 _3778_ (.Y(_1448_),
    .B1(_0629_),
    .B2(_0207_),
    .A2(_0626_),
    .A1(_2384_));
 sg13g2_a22oi_1 _3779_ (.Y(_1449_),
    .B1(_0630_),
    .B2(_2383_),
    .A2(_0625_),
    .A1(_2381_));
 sg13g2_xnor2_1 _3780_ (.Y(_1450_),
    .A(\pwm_module.prescaler0[10] ),
    .B(_0626_));
 sg13g2_nand3_1 _3781_ (.B(_1449_),
    .C(_1450_),
    .A(_1447_),
    .Y(_1451_));
 sg13g2_nand3b_1 _3782_ (.B(\MemCell.prescale_reg[1][1] ),
    .C(_0206_),
    .Y(_1452_),
    .A_N(net781));
 sg13g2_o21ai_1 _3783_ (.B1(_1452_),
    .Y(_1453_),
    .A1(\pwm_module.prescaler0[8] ),
    .A2(_0632_));
 sg13g2_and4_1 _3784_ (.A(_1447_),
    .B(_1449_),
    .C(_1450_),
    .D(_1453_),
    .X(_1454_));
 sg13g2_a21oi_1 _3785_ (.A1(_2383_),
    .A2(_0630_),
    .Y(_1455_),
    .B1(_1448_));
 sg13g2_o21ai_1 _3786_ (.B1(_1446_),
    .Y(_1456_),
    .A1(_1454_),
    .A2(_1455_));
 sg13g2_a21oi_1 _3787_ (.A1(_1444_),
    .A2(_1456_),
    .Y(_1457_),
    .B1(_1441_));
 sg13g2_nand2_1 _3788_ (.Y(_1458_),
    .A(_0209_),
    .B(_0613_));
 sg13g2_o21ai_1 _3789_ (.B1(_1458_),
    .Y(_1459_),
    .A1(\pwm_module.prescaler0[14] ),
    .A2(_0612_));
 sg13g2_nand2_1 _3790_ (.Y(_1460_),
    .A(\pwm_module.prescaler0[8] ),
    .B(_0632_));
 sg13g2_nand2_1 _3791_ (.Y(_1461_),
    .A(_1446_),
    .B(_1460_));
 sg13g2_or4_1 _3792_ (.A(_1445_),
    .B(_1453_),
    .C(_1459_),
    .D(_1461_),
    .X(_1462_));
 sg13g2_nor3_2 _3793_ (.A(_1441_),
    .B(_1451_),
    .C(_1462_),
    .Y(_1463_));
 sg13g2_a22oi_1 _3794_ (.Y(_1464_),
    .B1(_0579_),
    .B2(_0205_),
    .A2(_0577_),
    .A1(_2379_));
 sg13g2_or2_1 _3795_ (.X(_1465_),
    .B(_0585_),
    .A(\pwm_module.prescaler0[4] ));
 sg13g2_nand2_1 _3796_ (.Y(_1466_),
    .A(_0204_),
    .B(_0587_));
 sg13g2_and3_1 _3797_ (.X(_1467_),
    .A(_1464_),
    .B(_1465_),
    .C(_1466_));
 sg13g2_a22oi_1 _3798_ (.Y(_1468_),
    .B1(_0588_),
    .B2(_2378_),
    .A2(_0578_),
    .A1(\pwm_module.prescaler0[6] ));
 sg13g2_or2_1 _3799_ (.X(_1469_),
    .B(_0595_),
    .A(_0203_));
 sg13g2_nor2_1 _3800_ (.A(_0205_),
    .B(_0579_),
    .Y(_1470_));
 sg13g2_a21oi_1 _3801_ (.A1(\pwm_module.prescaler0[4] ),
    .A2(_0585_),
    .Y(_1471_),
    .B1(_1470_));
 sg13g2_nand4_1 _3802_ (.B(_1468_),
    .C(_1469_),
    .A(_1467_),
    .Y(_1472_),
    .D(_1471_));
 sg13g2_nand2_1 _3803_ (.Y(_1473_),
    .A(_0203_),
    .B(_0595_));
 sg13g2_o21ai_1 _3804_ (.B1(_1473_),
    .Y(_1474_),
    .A1(\pwm_module.prescaler0[2] ),
    .A2(_0594_));
 sg13g2_nand2_1 _3805_ (.Y(_1475_),
    .A(\pwm_module.prescaler0[2] ),
    .B(_0594_));
 sg13g2_a22oi_1 _3806_ (.Y(_1476_),
    .B1(_0603_),
    .B2(\pwm_module.prescaler0[1] ),
    .A2(_0602_),
    .A1(\pwm_module.prescaler0[0] ));
 sg13g2_nor2_1 _3807_ (.A(\pwm_module.prescaler0[1] ),
    .B(_0603_),
    .Y(_1477_));
 sg13g2_o21ai_1 _3808_ (.B1(_1475_),
    .Y(_1478_),
    .A1(_1476_),
    .A2(_1477_));
 sg13g2_nor2b_1 _3809_ (.A(_1474_),
    .B_N(_1478_),
    .Y(_1479_));
 sg13g2_and2_1 _3810_ (.A(_1468_),
    .B(_1471_),
    .X(_1480_));
 sg13g2_nand2_1 _3811_ (.Y(_1481_),
    .A(_1469_),
    .B(_1475_));
 sg13g2_nor2b_1 _3812_ (.A(_1468_),
    .B_N(_1464_),
    .Y(_1482_));
 sg13g2_or3_1 _3813_ (.A(_1467_),
    .B(_1470_),
    .C(_1482_),
    .X(_1483_));
 sg13g2_o21ai_1 _3814_ (.B1(_1483_),
    .Y(_1484_),
    .A1(_1472_),
    .A2(_1479_));
 sg13g2_a221oi_1 _3815_ (.B2(_1484_),
    .C1(_1457_),
    .B1(_1463_),
    .A1(_1439_),
    .Y(_1485_),
    .A2(_1459_));
 sg13g2_xnor2_1 _3816_ (.Y(_1486_),
    .A(_2387_),
    .B(_0565_));
 sg13g2_nand3b_1 _3817_ (.B(_1396_),
    .C(_1486_),
    .Y(_1487_),
    .A_N(_1395_));
 sg13g2_nor4_1 _3818_ (.A(_1394_),
    .B(_1429_),
    .C(_1431_),
    .D(_1487_),
    .Y(_1488_));
 sg13g2_nand2_1 _3819_ (.Y(_1489_),
    .A(_1421_),
    .B(_1488_));
 sg13g2_or2_1 _3820_ (.X(_1490_),
    .B(_1489_),
    .A(_1485_));
 sg13g2_nor2_1 _3821_ (.A(\pwm_module.prescaler0[0] ),
    .B(_0602_),
    .Y(_1491_));
 sg13g2_nand2b_1 _3822_ (.Y(_1492_),
    .B(_1476_),
    .A_N(_1477_));
 sg13g2_nor4_2 _3823_ (.A(_1474_),
    .B(_1481_),
    .C(_1491_),
    .Y(_1493_),
    .D(_1492_));
 sg13g2_nand4_1 _3824_ (.B(_1467_),
    .C(_1480_),
    .A(_1463_),
    .Y(_1494_),
    .D(_1493_));
 sg13g2_o21ai_1 _3825_ (.B1(_2396_),
    .Y(_1495_),
    .A1(_1489_),
    .A2(_1494_));
 sg13g2_a21oi_1 _3826_ (.A1(_1438_),
    .A2(_1490_),
    .Y(_1496_),
    .B1(_1495_));
 sg13g2_a21o_1 _3827_ (.A2(_1490_),
    .A1(_1438_),
    .B1(_1495_),
    .X(_1497_));
 sg13g2_nor2_1 _3828_ (.A(net238),
    .B(net661),
    .Y(_0000_));
 sg13g2_xnor2_1 _3829_ (.Y(_1498_),
    .A(net238),
    .B(net430));
 sg13g2_nor2_1 _3830_ (.A(net661),
    .B(_1498_),
    .Y(_0011_));
 sg13g2_and3_2 _3831_ (.X(_1499_),
    .A(net581),
    .B(\pwm_module.prescaler0[1] ),
    .C(net222));
 sg13g2_a21oi_1 _3832_ (.A1(\pwm_module.prescaler0[0] ),
    .A2(\pwm_module.prescaler0[1] ),
    .Y(_1500_),
    .B1(net222));
 sg13g2_nor3_1 _3833_ (.A(net660),
    .B(_1499_),
    .C(net223),
    .Y(_0022_));
 sg13g2_xor2_1 _3834_ (.B(_1499_),
    .A(net250),
    .X(_1501_));
 sg13g2_nor2_1 _3835_ (.A(net660),
    .B(net251),
    .Y(_0025_));
 sg13g2_and3_1 _3836_ (.X(_1502_),
    .A(\pwm_module.prescaler0[3] ),
    .B(\pwm_module.prescaler0[4] ),
    .C(_1499_));
 sg13g2_a21oi_1 _3837_ (.A1(\pwm_module.prescaler0[3] ),
    .A2(_1499_),
    .Y(_1503_),
    .B1(net317));
 sg13g2_nor3_1 _3838_ (.A(net660),
    .B(_1502_),
    .C(net318),
    .Y(_0026_));
 sg13g2_xnor2_1 _3839_ (.Y(_1504_),
    .A(_2378_),
    .B(_1502_));
 sg13g2_nor2_1 _3840_ (.A(net660),
    .B(net271),
    .Y(_0027_));
 sg13g2_and2_1 _3841_ (.A(\pwm_module.prescaler0[5] ),
    .B(\pwm_module.prescaler0[4] ),
    .X(_1505_));
 sg13g2_a21oi_1 _3842_ (.A1(net274),
    .A2(_1502_),
    .Y(_1506_),
    .B1(\pwm_module.prescaler0[6] ));
 sg13g2_and3_1 _3843_ (.X(_1507_),
    .A(net274),
    .B(\pwm_module.prescaler0[6] ),
    .C(_1502_));
 sg13g2_nor3_1 _3844_ (.A(net661),
    .B(net275),
    .C(_1507_),
    .Y(_0028_));
 sg13g2_xor2_1 _3845_ (.B(_1507_),
    .A(net257),
    .X(_1508_));
 sg13g2_nor2_1 _3846_ (.A(net660),
    .B(net258),
    .Y(_0029_));
 sg13g2_and2_1 _3847_ (.A(\pwm_module.prescaler0[7] ),
    .B(\pwm_module.prescaler0[6] ),
    .X(_1509_));
 sg13g2_and4_2 _3848_ (.A(\pwm_module.prescaler0[3] ),
    .B(_1499_),
    .C(_1505_),
    .D(_1509_),
    .X(_1510_));
 sg13g2_nand2_1 _3849_ (.Y(_1511_),
    .A(net523),
    .B(_1510_));
 sg13g2_o21ai_1 _3850_ (.B1(net668),
    .Y(_1512_),
    .A1(net523),
    .A2(_1510_));
 sg13g2_nor2b_1 _3851_ (.A(net524),
    .B_N(_1511_),
    .Y(_0030_));
 sg13g2_xnor2_1 _3852_ (.Y(_1513_),
    .A(net312),
    .B(_1511_));
 sg13g2_nor2_1 _3853_ (.A(net661),
    .B(net313),
    .Y(_0031_));
 sg13g2_nand3_1 _3854_ (.B(\pwm_module.prescaler0[8] ),
    .C(_1510_),
    .A(net459),
    .Y(_1514_));
 sg13g2_or2_1 _3855_ (.X(_1515_),
    .B(_1514_),
    .A(_2384_));
 sg13g2_nand2_1 _3856_ (.Y(_1516_),
    .A(net668),
    .B(_1515_));
 sg13g2_a21oi_1 _3857_ (.A1(_2384_),
    .A2(net460),
    .Y(_0001_),
    .B1(_1516_));
 sg13g2_xnor2_1 _3858_ (.Y(_1517_),
    .A(net333),
    .B(_1515_));
 sg13g2_nor2_1 _3859_ (.A(net661),
    .B(_1517_),
    .Y(_0002_));
 sg13g2_nor3_2 _3860_ (.A(_2382_),
    .B(_2384_),
    .C(_1514_),
    .Y(_1518_));
 sg13g2_nand2_1 _3861_ (.Y(_1519_),
    .A(net489),
    .B(_1518_));
 sg13g2_and4_1 _3862_ (.A(\pwm_module.prescaler0[9] ),
    .B(\pwm_module.prescaler0[8] ),
    .C(\pwm_module.prescaler0[11] ),
    .D(\pwm_module.prescaler0[10] ),
    .X(_1520_));
 sg13g2_o21ai_1 _3863_ (.B1(net668),
    .Y(_1521_),
    .A1(net489),
    .A2(_1518_));
 sg13g2_nor2b_1 _3864_ (.A(net490),
    .B_N(_1519_),
    .Y(_0003_));
 sg13g2_xnor2_1 _3865_ (.Y(_1522_),
    .A(net129),
    .B(_1519_));
 sg13g2_nor2_1 _3866_ (.A(net661),
    .B(net130),
    .Y(_0004_));
 sg13g2_nand3_1 _3867_ (.B(\pwm_module.prescaler0[12] ),
    .C(_1518_),
    .A(\pwm_module.prescaler0[13] ),
    .Y(_1523_));
 sg13g2_nand4_1 _3868_ (.B(\pwm_module.prescaler0[12] ),
    .C(_1510_),
    .A(\pwm_module.prescaler0[13] ),
    .Y(_1524_),
    .D(_1520_));
 sg13g2_or2_1 _3869_ (.X(_1525_),
    .B(_1523_),
    .A(_2380_));
 sg13g2_nand2_1 _3870_ (.Y(_1526_),
    .A(net668),
    .B(_1525_));
 sg13g2_a21oi_1 _3871_ (.A1(_2380_),
    .A2(_1524_),
    .Y(_0005_),
    .B1(_1526_));
 sg13g2_xnor2_1 _3872_ (.Y(_1527_),
    .A(net263),
    .B(_1525_));
 sg13g2_nor2_1 _3873_ (.A(net661),
    .B(_1527_),
    .Y(_0006_));
 sg13g2_nand2_2 _3874_ (.Y(_1528_),
    .A(\pwm_module.prescaler0[15] ),
    .B(\pwm_module.prescaler0[14] ));
 sg13g2_nor3_2 _3875_ (.A(_2387_),
    .B(_1523_),
    .C(_1528_),
    .Y(_1529_));
 sg13g2_nor2_1 _3876_ (.A(_1524_),
    .B(_1528_),
    .Y(_1530_));
 sg13g2_nor2_1 _3877_ (.A(net376),
    .B(_1530_),
    .Y(_1531_));
 sg13g2_nor3_1 _3878_ (.A(net663),
    .B(_1529_),
    .C(net377),
    .Y(_0007_));
 sg13g2_xor2_1 _3879_ (.B(_1529_),
    .A(net204),
    .X(_1532_));
 sg13g2_nor2_1 _3880_ (.A(net663),
    .B(net205),
    .Y(_0008_));
 sg13g2_a21oi_1 _3881_ (.A1(net328),
    .A2(_1529_),
    .Y(_1533_),
    .B1(\pwm_module.prescaler0[18] ));
 sg13g2_nand3_1 _3882_ (.B(net328),
    .C(_1529_),
    .A(\pwm_module.prescaler0[18] ),
    .Y(_1534_));
 sg13g2_nand2_1 _3883_ (.Y(_1535_),
    .A(_1496_),
    .B(_1534_));
 sg13g2_nor2_1 _3884_ (.A(net329),
    .B(_1535_),
    .Y(_0009_));
 sg13g2_xnor2_1 _3885_ (.Y(_1536_),
    .A(net324),
    .B(_1534_));
 sg13g2_nor2_1 _3886_ (.A(net663),
    .B(net325),
    .Y(_0010_));
 sg13g2_nand4_1 _3887_ (.B(\pwm_module.prescaler0[18] ),
    .C(\pwm_module.prescaler0[17] ),
    .A(\pwm_module.prescaler0[19] ),
    .Y(_1537_),
    .D(\pwm_module.prescaler0[16] ));
 sg13g2_or3_1 _3888_ (.A(_1524_),
    .B(_1528_),
    .C(_1537_),
    .X(_1538_));
 sg13g2_and2_1 _3889_ (.A(net353),
    .B(_1538_),
    .X(_1539_));
 sg13g2_nor2_1 _3890_ (.A(net353),
    .B(_1538_),
    .Y(_1540_));
 sg13g2_nor3_1 _3891_ (.A(net663),
    .B(net354),
    .C(_1540_),
    .Y(_0012_));
 sg13g2_xor2_1 _3892_ (.B(_1540_),
    .A(net187),
    .X(_1541_));
 sg13g2_nor2_1 _3893_ (.A(net663),
    .B(net188),
    .Y(_0013_));
 sg13g2_nand2_1 _3894_ (.Y(_1542_),
    .A(\pwm_module.prescaler0[20] ),
    .B(\pwm_module.prescaler0[21] ));
 sg13g2_nor4_2 _3895_ (.A(_1524_),
    .B(_1528_),
    .C(_1537_),
    .Y(_1543_),
    .D(_1542_));
 sg13g2_or2_1 _3896_ (.X(_1544_),
    .B(_1543_),
    .A(net565));
 sg13g2_nand2_1 _3897_ (.Y(_1545_),
    .A(net565),
    .B(_1543_));
 sg13g2_and3_1 _3898_ (.X(_0014_),
    .A(net669),
    .B(net566),
    .C(_1545_));
 sg13g2_xnor2_1 _3899_ (.Y(_1546_),
    .A(net305),
    .B(_1545_));
 sg13g2_nor2_1 _3900_ (.A(net663),
    .B(net306),
    .Y(_0015_));
 sg13g2_and3_1 _3901_ (.X(_1547_),
    .A(\pwm_module.prescaler0[23] ),
    .B(\pwm_module.prescaler0[22] ),
    .C(_1543_));
 sg13g2_or2_1 _3902_ (.X(_1548_),
    .B(_1547_),
    .A(net562));
 sg13g2_nand2_1 _3903_ (.Y(_1549_),
    .A(net562),
    .B(_1547_));
 sg13g2_and3_1 _3904_ (.X(_0016_),
    .A(net669),
    .B(net563),
    .C(_1549_));
 sg13g2_xnor2_1 _3905_ (.Y(_1550_),
    .A(net292),
    .B(_1549_));
 sg13g2_nor2_1 _3906_ (.A(net664),
    .B(net293),
    .Y(_0017_));
 sg13g2_nand3_1 _3907_ (.B(\pwm_module.prescaler0[24] ),
    .C(_1547_),
    .A(\pwm_module.prescaler0[25] ),
    .Y(_1551_));
 sg13g2_and2_1 _3908_ (.A(net486),
    .B(_1551_),
    .X(_1552_));
 sg13g2_nor2_1 _3909_ (.A(net486),
    .B(_1551_),
    .Y(_1553_));
 sg13g2_nor3_1 _3910_ (.A(net664),
    .B(_1552_),
    .C(net487),
    .Y(_0018_));
 sg13g2_xnor2_1 _3911_ (.Y(_1554_),
    .A(_2385_),
    .B(net487));
 sg13g2_nor2_1 _3912_ (.A(net663),
    .B(_1554_),
    .Y(_0019_));
 sg13g2_nand2_1 _3913_ (.Y(_1555_),
    .A(\pwm_module.prescaler0[26] ),
    .B(\pwm_module.prescaler0[27] ));
 sg13g2_nor2_2 _3914_ (.A(_1551_),
    .B(_1555_),
    .Y(_1556_));
 sg13g2_nor2_1 _3915_ (.A(net417),
    .B(_1556_),
    .Y(_1557_));
 sg13g2_and2_1 _3916_ (.A(net417),
    .B(_1556_),
    .X(_1558_));
 sg13g2_nor3_1 _3917_ (.A(net663),
    .B(net418),
    .C(_1558_),
    .Y(_0020_));
 sg13g2_xnor2_1 _3918_ (.Y(_1559_),
    .A(net416),
    .B(_1558_));
 sg13g2_and2_1 _3919_ (.A(net669),
    .B(_1559_),
    .X(_0021_));
 sg13g2_and2_1 _3920_ (.A(\pwm_module.prescaler0[28] ),
    .B(\pwm_module.prescaler0[29] ),
    .X(_1560_));
 sg13g2_a21oi_1 _3921_ (.A1(_1556_),
    .A2(_1560_),
    .Y(_1561_),
    .B1(net381));
 sg13g2_and3_1 _3922_ (.X(_1562_),
    .A(net381),
    .B(_1556_),
    .C(_1560_));
 sg13g2_nor3_1 _3923_ (.A(net664),
    .B(net382),
    .C(_1562_),
    .Y(_0023_));
 sg13g2_xnor2_1 _3924_ (.Y(_1563_),
    .A(net532),
    .B(_1562_));
 sg13g2_and2_1 _3925_ (.A(net669),
    .B(_1563_),
    .X(_0024_));
 sg13g2_nor2_1 _3926_ (.A(net357),
    .B(net670),
    .Y(_0032_));
 sg13g2_xnor2_1 _3927_ (.Y(_1564_),
    .A(net357),
    .B(net476));
 sg13g2_nor2_1 _3928_ (.A(net670),
    .B(_1564_),
    .Y(_0043_));
 sg13g2_a21oi_1 _3929_ (.A1(\pwm_module.prescaler1[0] ),
    .A2(\pwm_module.prescaler1[1] ),
    .Y(_1565_),
    .B1(net226));
 sg13g2_nor3_1 _3930_ (.A(net670),
    .B(_0657_),
    .C(net227),
    .Y(_0054_));
 sg13g2_xor2_1 _3931_ (.B(_0657_),
    .A(net423),
    .X(_1566_));
 sg13g2_nor2_1 _3932_ (.A(net670),
    .B(net424),
    .Y(_0057_));
 sg13g2_nand3_1 _3933_ (.B(\pwm_module.prescaler1[4] ),
    .C(_0657_),
    .A(\pwm_module.prescaler1[3] ),
    .Y(_1567_));
 sg13g2_xor2_1 _3934_ (.B(_0658_),
    .A(net501),
    .X(_1568_));
 sg13g2_nor2_1 _3935_ (.A(net670),
    .B(net502),
    .Y(_0058_));
 sg13g2_xnor2_1 _3936_ (.Y(_1569_),
    .A(net447),
    .B(_1567_));
 sg13g2_nor2_1 _3937_ (.A(net670),
    .B(net448),
    .Y(_0059_));
 sg13g2_nand2_1 _3938_ (.Y(_1570_),
    .A(\pwm_module.prescaler1[6] ),
    .B(_0660_));
 sg13g2_xnor2_1 _3939_ (.Y(_1571_),
    .A(net449),
    .B(_0660_));
 sg13g2_nor2_1 _3940_ (.A(net670),
    .B(net450),
    .Y(_0060_));
 sg13g2_xnor2_1 _3941_ (.Y(_1572_),
    .A(net111),
    .B(_1570_));
 sg13g2_nor2_1 _3942_ (.A(net670),
    .B(net112),
    .Y(_0061_));
 sg13g2_nand2_1 _3943_ (.Y(_1573_),
    .A(\pwm_module.prescaler1[8] ),
    .B(_0662_));
 sg13g2_xnor2_1 _3944_ (.Y(_1574_),
    .A(net472),
    .B(_0662_));
 sg13g2_nor2_1 _3945_ (.A(net673),
    .B(net473),
    .Y(_0062_));
 sg13g2_xnor2_1 _3946_ (.Y(_1575_),
    .A(net179),
    .B(_1573_));
 sg13g2_nor2_1 _3947_ (.A(net673),
    .B(net180),
    .Y(_0063_));
 sg13g2_nand2_1 _3948_ (.Y(_1576_),
    .A(\pwm_module.prescaler1[10] ),
    .B(_0664_));
 sg13g2_xnor2_1 _3949_ (.Y(_1577_),
    .A(net439),
    .B(_0664_));
 sg13g2_nor2_1 _3950_ (.A(net672),
    .B(net440),
    .Y(_0033_));
 sg13g2_xnor2_1 _3951_ (.Y(_1578_),
    .A(net267),
    .B(_1576_));
 sg13g2_nor2_1 _3952_ (.A(net672),
    .B(net268),
    .Y(_0034_));
 sg13g2_nor2_1 _3953_ (.A(_0174_),
    .B(_0666_),
    .Y(_1579_));
 sg13g2_xnor2_1 _3954_ (.Y(_1580_),
    .A(net338),
    .B(_0666_));
 sg13g2_nor2_1 _3955_ (.A(net672),
    .B(net339),
    .Y(_0035_));
 sg13g2_xor2_1 _3956_ (.B(_1579_),
    .A(net190),
    .X(_1581_));
 sg13g2_nor2_1 _3957_ (.A(net672),
    .B(net191),
    .Y(_0036_));
 sg13g2_nand2_1 _3958_ (.Y(_1582_),
    .A(\pwm_module.prescaler1[14] ),
    .B(_0668_));
 sg13g2_xnor2_1 _3959_ (.Y(_1583_),
    .A(net457),
    .B(_0668_));
 sg13g2_nor2_1 _3960_ (.A(net672),
    .B(net458),
    .Y(_0037_));
 sg13g2_xnor2_1 _3961_ (.Y(_1584_),
    .A(net142),
    .B(_1582_));
 sg13g2_nor2_1 _3962_ (.A(net672),
    .B(net143),
    .Y(_0038_));
 sg13g2_nor2_1 _3963_ (.A(net469),
    .B(_0670_),
    .Y(_1585_));
 sg13g2_nor3_1 _3964_ (.A(net675),
    .B(_0672_),
    .C(_1585_),
    .Y(_0039_));
 sg13g2_xnor2_1 _3965_ (.Y(_1586_),
    .A(_2377_),
    .B(_0672_));
 sg13g2_nor2_1 _3966_ (.A(net675),
    .B(net380),
    .Y(_0040_));
 sg13g2_nor2b_2 _3967_ (.A(net790),
    .B_N(\MemCell.counter_value[29] ),
    .Y(_1587_));
 sg13g2_xnor2_1 _3968_ (.Y(_1588_),
    .A(\pwm_module.counter0[29] ),
    .B(_1587_));
 sg13g2_nor2b_2 _3969_ (.A(net791),
    .B_N(\MemCell.counter_value[30] ),
    .Y(_1589_));
 sg13g2_nand2b_2 _3970_ (.Y(_1590_),
    .B(\MemCell.counter_value[30] ),
    .A_N(net791));
 sg13g2_nor2b_2 _3971_ (.A(net790),
    .B_N(\MemCell.counter_value[31] ),
    .Y(_1591_));
 sg13g2_nor2_1 _3972_ (.A(_0167_),
    .B(_1591_),
    .Y(_1592_));
 sg13g2_nor2b_2 _3973_ (.A(net790),
    .B_N(\MemCell.counter_value[26] ),
    .Y(_1593_));
 sg13g2_nand2b_2 _3974_ (.Y(_1594_),
    .B(\MemCell.counter_value[26] ),
    .A_N(net790));
 sg13g2_nor2b_2 _3975_ (.A(net790),
    .B_N(\MemCell.counter_value[27] ),
    .Y(_1595_));
 sg13g2_nand2_1 _3976_ (.Y(_1596_),
    .A(_0146_),
    .B(_1595_));
 sg13g2_o21ai_1 _3977_ (.B1(_1596_),
    .Y(_1597_),
    .A1(\pwm_module.counter0[26] ),
    .A2(_1594_));
 sg13g2_nor2b_2 _3978_ (.A(net790),
    .B_N(\MemCell.counter_value[25] ),
    .Y(_1598_));
 sg13g2_nand2b_1 _3979_ (.Y(_1599_),
    .B(\MemCell.counter_value[25] ),
    .A_N(net791));
 sg13g2_xnor2_1 _3980_ (.Y(_1600_),
    .A(\pwm_module.counter0[25] ),
    .B(_1598_));
 sg13g2_nand2b_2 _3981_ (.Y(_1601_),
    .B(\MemCell.counter_value[28] ),
    .A_N(net790));
 sg13g2_nand2b_2 _3982_ (.Y(_1602_),
    .B(\MemCell.counter_value[24] ),
    .A_N(net790));
 sg13g2_nor2_1 _3983_ (.A(\pwm_module.counter0[28] ),
    .B(_1601_),
    .Y(_1603_));
 sg13g2_or2_1 _3984_ (.X(_1604_),
    .B(_1595_),
    .A(_0146_));
 sg13g2_nor2_1 _3985_ (.A(\pwm_module.counter0[24] ),
    .B(_1602_),
    .Y(_1605_));
 sg13g2_xnor2_1 _3986_ (.Y(_1606_),
    .A(\pwm_module.counter0[30] ),
    .B(_1589_));
 sg13g2_xor2_1 _3987_ (.B(_1591_),
    .A(_0167_),
    .X(_1607_));
 sg13g2_nand2_1 _3988_ (.Y(_1608_),
    .A(_1606_),
    .B(_1607_));
 sg13g2_xor2_1 _3989_ (.B(_1601_),
    .A(\pwm_module.counter0[28] ),
    .X(_1609_));
 sg13g2_and4_1 _3990_ (.A(_1588_),
    .B(_1606_),
    .C(_1607_),
    .D(_1609_),
    .X(_1610_));
 sg13g2_nand4_1 _3991_ (.B(_1606_),
    .C(_1607_),
    .A(_1588_),
    .Y(_1611_),
    .D(_1609_));
 sg13g2_o21ai_1 _3992_ (.B1(_1604_),
    .Y(_1612_),
    .A1(_2349_),
    .A2(_1593_));
 sg13g2_xnor2_1 _3993_ (.Y(_1613_),
    .A(_2350_),
    .B(_1602_));
 sg13g2_nand2_1 _3994_ (.Y(_1614_),
    .A(_1600_),
    .B(_1613_));
 sg13g2_or4_1 _3995_ (.A(_1597_),
    .B(_1611_),
    .C(_1612_),
    .D(_1614_),
    .X(_1615_));
 sg13g2_nor2b_2 _3996_ (.A(net792),
    .B_N(\MemCell.counter_value[21] ),
    .Y(_1616_));
 sg13g2_nand2b_1 _3997_ (.Y(_1617_),
    .B(\MemCell.counter_value[21] ),
    .A_N(net793));
 sg13g2_xnor2_1 _3998_ (.Y(_1618_),
    .A(\pwm_module.counter0[21] ),
    .B(_1616_));
 sg13g2_nand2b_2 _3999_ (.Y(_1619_),
    .B(\MemCell.counter_value[16] ),
    .A_N(net788));
 sg13g2_nor2_1 _4000_ (.A(\pwm_module.counter0[16] ),
    .B(_1619_),
    .Y(_1620_));
 sg13g2_xnor2_1 _4001_ (.Y(_1621_),
    .A(_2352_),
    .B(_1619_));
 sg13g2_nor2b_2 _4002_ (.A(net792),
    .B_N(\MemCell.counter_value[23] ),
    .Y(_1622_));
 sg13g2_nand2b_1 _4003_ (.Y(_1623_),
    .B(\MemCell.counter_value[23] ),
    .A_N(net792));
 sg13g2_nor2b_2 _4004_ (.A(net792),
    .B_N(\MemCell.counter_value[22] ),
    .Y(_1624_));
 sg13g2_nand2b_1 _4005_ (.Y(_1625_),
    .B(\MemCell.counter_value[22] ),
    .A_N(net793));
 sg13g2_a22oi_1 _4006_ (.Y(_1626_),
    .B1(_1624_),
    .B2(_2351_),
    .A2(_1622_),
    .A1(_0148_));
 sg13g2_nor2b_2 _4007_ (.A(net789),
    .B_N(\MemCell.counter_value[17] ),
    .Y(_1627_));
 sg13g2_nand2b_1 _4008_ (.Y(_1628_),
    .B(\MemCell.counter_value[17] ),
    .A_N(net792));
 sg13g2_xnor2_1 _4009_ (.Y(_1629_),
    .A(\pwm_module.counter0[17] ),
    .B(_1627_));
 sg13g2_nor2_1 _4010_ (.A(_0148_),
    .B(_1622_),
    .Y(_1630_));
 sg13g2_nor2b_1 _4011_ (.A(net792),
    .B_N(\MemCell.counter_value[20] ),
    .Y(_1631_));
 sg13g2_nand2b_2 _4012_ (.Y(_1632_),
    .B(\MemCell.counter_value[20] ),
    .A_N(net792));
 sg13g2_nor2_1 _4013_ (.A(\pwm_module.counter0[20] ),
    .B(_1632_),
    .Y(_1633_));
 sg13g2_nor2_1 _4014_ (.A(_1630_),
    .B(_1633_),
    .Y(_1634_));
 sg13g2_nor2_1 _4015_ (.A(_2351_),
    .B(_1624_),
    .Y(_1635_));
 sg13g2_a21oi_1 _4016_ (.A1(\pwm_module.counter0[20] ),
    .A2(_1632_),
    .Y(_1636_),
    .B1(_1635_));
 sg13g2_nor2b_2 _4017_ (.A(net788),
    .B_N(\MemCell.counter_value[19] ),
    .Y(_1637_));
 sg13g2_nor2_1 _4018_ (.A(_0151_),
    .B(_1637_),
    .Y(_1638_));
 sg13g2_or2_1 _4019_ (.X(_1639_),
    .B(_1637_),
    .A(_0151_));
 sg13g2_and2_1 _4020_ (.A(_0151_),
    .B(_1637_),
    .X(_1640_));
 sg13g2_nand2b_2 _4021_ (.Y(_1641_),
    .B(\MemCell.counter_value[18] ),
    .A_N(net788));
 sg13g2_and2_1 _4022_ (.A(\pwm_module.counter0[18] ),
    .B(_1641_),
    .X(_1642_));
 sg13g2_nor2_1 _4023_ (.A(\pwm_module.counter0[18] ),
    .B(_1641_),
    .Y(_1643_));
 sg13g2_or4_1 _4024_ (.A(_1638_),
    .B(_1640_),
    .C(_1642_),
    .D(_1643_),
    .X(_1644_));
 sg13g2_nand4_1 _4025_ (.B(_1626_),
    .C(_1634_),
    .A(_1618_),
    .Y(_1645_),
    .D(_1636_));
 sg13g2_nand2_1 _4026_ (.Y(_1646_),
    .A(_1621_),
    .B(_1629_));
 sg13g2_nor4_2 _4027_ (.A(_1615_),
    .B(_1644_),
    .C(_1645_),
    .Y(_1647_),
    .D(_1646_));
 sg13g2_nor2b_2 _4028_ (.A(net788),
    .B_N(\MemCell.counter_value[15] ),
    .Y(_1648_));
 sg13g2_or2_1 _4029_ (.X(_1649_),
    .B(_1648_),
    .A(_0153_));
 sg13g2_nor2b_1 _4030_ (.A(net795),
    .B_N(\MemCell.counter_value[14] ),
    .Y(_1650_));
 sg13g2_nand2b_2 _4031_ (.Y(_1651_),
    .B(\MemCell.counter_value[14] ),
    .A_N(net795));
 sg13g2_nand3b_1 _4032_ (.B(\MemCell.counter_value[15] ),
    .C(_0153_),
    .Y(_1652_),
    .A_N(net788));
 sg13g2_o21ai_1 _4033_ (.B1(_1652_),
    .Y(_1653_),
    .A1(\pwm_module.counter0[14] ),
    .A2(_1651_));
 sg13g2_nand2_1 _4034_ (.Y(_1654_),
    .A(\pwm_module.counter0[14] ),
    .B(_1651_));
 sg13g2_nor2b_2 _4035_ (.A(net795),
    .B_N(\MemCell.counter_value[13] ),
    .Y(_1655_));
 sg13g2_nand2b_1 _4036_ (.Y(_1656_),
    .B(\MemCell.counter_value[13] ),
    .A_N(net795));
 sg13g2_xnor2_1 _4037_ (.Y(_1657_),
    .A(\pwm_module.counter0[13] ),
    .B(_1655_));
 sg13g2_nor2b_2 _4038_ (.A(net795),
    .B_N(\MemCell.counter_value[12] ),
    .Y(_1658_));
 sg13g2_o21ai_1 _4039_ (.B1(_1657_),
    .Y(_1659_),
    .A1(_2354_),
    .A2(_1658_));
 sg13g2_nor2_2 _4040_ (.A(\MemCell.counter_value[10] ),
    .B(net789),
    .Y(_1660_));
 sg13g2_xnor2_1 _4041_ (.Y(_1661_),
    .A(_0157_),
    .B(_1660_));
 sg13g2_nor2b_2 _4042_ (.A(net788),
    .B_N(\MemCell.counter_value[11] ),
    .Y(_1662_));
 sg13g2_nand3b_1 _4043_ (.B(\MemCell.counter_value[11] ),
    .C(_0156_),
    .Y(_1663_),
    .A_N(net788));
 sg13g2_or2_1 _4044_ (.X(_1664_),
    .B(_1662_),
    .A(_0156_));
 sg13g2_nand3_1 _4045_ (.B(_1663_),
    .C(_1664_),
    .A(_1661_),
    .Y(_1665_));
 sg13g2_nor2b_2 _4046_ (.A(net789),
    .B_N(\MemCell.counter_value[9] ),
    .Y(_1666_));
 sg13g2_xnor2_1 _4047_ (.Y(_1667_),
    .A(\pwm_module.counter0[9] ),
    .B(_1666_));
 sg13g2_nand2b_2 _4048_ (.Y(_1668_),
    .B(\MemCell.counter_value[8] ),
    .A_N(net788));
 sg13g2_nor2_1 _4049_ (.A(\pwm_module.counter0[8] ),
    .B(_1668_),
    .Y(_1669_));
 sg13g2_a22oi_1 _4050_ (.Y(_1670_),
    .B1(_1667_),
    .B2(_1669_),
    .A2(_1666_),
    .A1(_0158_));
 sg13g2_and2_1 _4051_ (.A(_2354_),
    .B(_1658_),
    .X(_1671_));
 sg13g2_o21ai_1 _4052_ (.B1(_1663_),
    .Y(_1672_),
    .A1(\pwm_module.counter0[10] ),
    .A2(_1660_));
 sg13g2_o21ai_1 _4053_ (.B1(_1672_),
    .Y(_1673_),
    .A1(_0156_),
    .A2(_1662_));
 sg13g2_nand3b_1 _4054_ (.B(_1654_),
    .C(_1649_),
    .Y(_1674_),
    .A_N(_1653_));
 sg13g2_a22oi_1 _4055_ (.Y(_1675_),
    .B1(_1657_),
    .B2(_1671_),
    .A2(_1655_),
    .A1(_0154_));
 sg13g2_nor2_1 _4056_ (.A(_1674_),
    .B(_1675_),
    .Y(_1676_));
 sg13g2_nor3_1 _4057_ (.A(_1659_),
    .B(_1671_),
    .C(_1674_),
    .Y(_1677_));
 sg13g2_o21ai_1 _4058_ (.B1(_1673_),
    .Y(_1678_),
    .A1(_1665_),
    .A2(_1670_));
 sg13g2_a221oi_1 _4059_ (.B2(_1678_),
    .C1(_1676_),
    .B1(_1677_),
    .A1(_1649_),
    .Y(_1679_),
    .A2(_1653_));
 sg13g2_nor2_2 _4060_ (.A(\MemCell.counter_value[7] ),
    .B(net794),
    .Y(_1680_));
 sg13g2_or2_1 _4061_ (.X(_1681_),
    .B(_1680_),
    .A(\pwm_module.counter0[7] ));
 sg13g2_nor2_2 _4062_ (.A(\MemCell.counter_value[6] ),
    .B(net794),
    .Y(_1682_));
 sg13g2_or2_1 _4063_ (.X(_1683_),
    .B(net795),
    .A(\MemCell.counter_value[6] ));
 sg13g2_o21ai_1 _4064_ (.B1(_1681_),
    .Y(_1684_),
    .A1(\pwm_module.counter0[6] ),
    .A2(_1682_));
 sg13g2_xnor2_1 _4065_ (.Y(_1685_),
    .A(_0160_),
    .B(_1682_));
 sg13g2_nor2_2 _4066_ (.A(\MemCell.counter_value[5] ),
    .B(net794),
    .Y(_1686_));
 sg13g2_or2_2 _4067_ (.X(_1687_),
    .B(net794),
    .A(\MemCell.counter_value[5] ));
 sg13g2_nand2b_1 _4068_ (.Y(_1688_),
    .B(_1687_),
    .A_N(\pwm_module.counter0[5] ));
 sg13g2_xnor2_1 _4069_ (.Y(_1689_),
    .A(_0161_),
    .B(_1686_));
 sg13g2_nor2b_2 _4070_ (.A(net794),
    .B_N(\MemCell.counter_value[4] ),
    .Y(_1690_));
 sg13g2_nor2b_2 _4071_ (.A(net794),
    .B_N(\MemCell.counter_value[3] ),
    .Y(_1691_));
 sg13g2_nand2_1 _4072_ (.Y(_1692_),
    .A(_0163_),
    .B(_1691_));
 sg13g2_nand2b_2 _4073_ (.Y(_1693_),
    .B(\MemCell.counter_value[2] ),
    .A_N(net794));
 sg13g2_o21ai_1 _4074_ (.B1(_1692_),
    .Y(_1694_),
    .A1(\pwm_module.counter0[2] ),
    .A2(_1693_));
 sg13g2_nor2_2 _4075_ (.A(\MemCell.counter_value[1] ),
    .B(net794),
    .Y(_1695_));
 sg13g2_a22oi_1 _4076_ (.Y(_1696_),
    .B1(_1695_),
    .B2(\pwm_module.counter0[1] ),
    .A2(_1693_),
    .A1(\pwm_module.counter0[2] ));
 sg13g2_or2_1 _4077_ (.X(_1697_),
    .B(_1695_),
    .A(\pwm_module.counter0[1] ));
 sg13g2_nand2b_2 _4078_ (.Y(_1698_),
    .B(\MemCell.counter_value[0] ),
    .A_N(net795));
 sg13g2_nand3_1 _4079_ (.B(_1697_),
    .C(_1698_),
    .A(net754),
    .Y(_1699_));
 sg13g2_a21o_1 _4080_ (.A2(_1699_),
    .A1(_1696_),
    .B1(_1694_),
    .X(_1700_));
 sg13g2_nand2_1 _4081_ (.Y(_1701_),
    .A(\pwm_module.counter0[8] ),
    .B(_1668_));
 sg13g2_nor2_1 _4082_ (.A(_1665_),
    .B(_1669_),
    .Y(_1702_));
 sg13g2_and4_1 _4083_ (.A(_1667_),
    .B(_1677_),
    .C(_1701_),
    .D(_1702_),
    .X(_1703_));
 sg13g2_nand4_1 _4084_ (.B(_1677_),
    .C(_1701_),
    .A(_1667_),
    .Y(_1704_),
    .D(_1702_));
 sg13g2_nand2_1 _4085_ (.Y(_1705_),
    .A(\pwm_module.counter0[7] ),
    .B(_1680_));
 sg13g2_nand3_1 _4086_ (.B(_1685_),
    .C(_1705_),
    .A(_1681_),
    .Y(_1706_));
 sg13g2_nand3_1 _4087_ (.B(_1689_),
    .C(_1690_),
    .A(_0162_),
    .Y(_1707_));
 sg13g2_a21oi_1 _4088_ (.A1(_1688_),
    .A2(_1707_),
    .Y(_1708_),
    .B1(_1706_));
 sg13g2_xnor2_1 _4089_ (.Y(_1709_),
    .A(_0162_),
    .B(_1690_));
 sg13g2_o21ai_1 _4090_ (.B1(_1689_),
    .Y(_1710_),
    .A1(_0163_),
    .A2(_1691_));
 sg13g2_nor3_1 _4091_ (.A(_1706_),
    .B(_1709_),
    .C(_1710_),
    .Y(_1711_));
 sg13g2_a221oi_1 _4092_ (.B2(_1700_),
    .C1(_1708_),
    .B1(_1711_),
    .A1(_1684_),
    .Y(_1712_),
    .A2(_1705_));
 sg13g2_o21ai_1 _4093_ (.B1(_1679_),
    .Y(_1713_),
    .A1(_1704_),
    .A2(_1712_));
 sg13g2_a22oi_1 _4094_ (.Y(_1714_),
    .B1(_1600_),
    .B2(_1605_),
    .A2(_1598_),
    .A1(_0147_));
 sg13g2_nor3_1 _4095_ (.A(_1597_),
    .B(_1612_),
    .C(_1714_),
    .Y(_1715_));
 sg13g2_a21o_1 _4096_ (.A2(_1604_),
    .A1(_1597_),
    .B1(_1715_),
    .X(_1716_));
 sg13g2_a22oi_1 _4097_ (.Y(_1717_),
    .B1(_1588_),
    .B2(_1603_),
    .A2(_1587_),
    .A1(_0145_));
 sg13g2_nor3_1 _4098_ (.A(\pwm_module.counter0[30] ),
    .B(_1590_),
    .C(_1592_),
    .Y(_1718_));
 sg13g2_a21oi_1 _4099_ (.A1(_0167_),
    .A2(_1591_),
    .Y(_1719_),
    .B1(_1718_));
 sg13g2_o21ai_1 _4100_ (.B1(_1719_),
    .Y(_1720_),
    .A1(_1608_),
    .A2(_1717_));
 sg13g2_a21oi_1 _4101_ (.A1(_1610_),
    .A2(_1716_),
    .Y(_1721_),
    .B1(_1720_));
 sg13g2_a22oi_1 _4102_ (.Y(_1722_),
    .B1(_1629_),
    .B2(_1620_),
    .A2(_1627_),
    .A1(_0152_));
 sg13g2_a22oi_1 _4103_ (.Y(_1723_),
    .B1(_1618_),
    .B2(_1633_),
    .A2(_1616_),
    .A1(_0149_));
 sg13g2_o21ai_1 _4104_ (.B1(_1626_),
    .Y(_1724_),
    .A1(_1635_),
    .A2(_1723_));
 sg13g2_nand2b_1 _4105_ (.Y(_1725_),
    .B(_1724_),
    .A_N(_1630_));
 sg13g2_a21oi_1 _4106_ (.A1(_1639_),
    .A2(_1643_),
    .Y(_1726_),
    .B1(_1640_));
 sg13g2_o21ai_1 _4107_ (.B1(_1726_),
    .Y(_1727_),
    .A1(_1644_),
    .A2(_1722_));
 sg13g2_nand2b_1 _4108_ (.Y(_1728_),
    .B(_1727_),
    .A_N(_1645_));
 sg13g2_a21oi_1 _4109_ (.A1(_1725_),
    .A2(_1728_),
    .Y(_1729_),
    .B1(_1615_));
 sg13g2_a21oi_1 _4110_ (.A1(_1647_),
    .A2(_1713_),
    .Y(_1730_),
    .B1(_1729_));
 sg13g2_xnor2_1 _4111_ (.Y(_1731_),
    .A(_0165_),
    .B(_1698_));
 sg13g2_and3_1 _4112_ (.X(_1732_),
    .A(_1696_),
    .B(_1697_),
    .C(_1731_));
 sg13g2_nor2b_1 _4113_ (.A(_1694_),
    .B_N(_1732_),
    .Y(_1733_));
 sg13g2_nand4_1 _4114_ (.B(_1703_),
    .C(_1711_),
    .A(_1647_),
    .Y(_1734_),
    .D(_1733_));
 sg13g2_nand2_1 _4115_ (.Y(_1735_),
    .A(_2396_),
    .B(_1734_));
 sg13g2_a21oi_2 _4116_ (.B1(_1735_),
    .Y(_1736_),
    .A2(_1730_),
    .A1(_1721_));
 sg13g2_nand2_1 _4117_ (.Y(_1737_),
    .A(net659),
    .B(_1736_));
 sg13g2_nand2_1 _4118_ (.Y(_1738_),
    .A(net79),
    .B(net665));
 sg13g2_o21ai_1 _4119_ (.B1(_1738_),
    .Y(_0223_),
    .A1(net754),
    .A2(net653));
 sg13g2_nor2_2 _4120_ (.A(net667),
    .B(_1736_),
    .Y(_1739_));
 sg13g2_and3_1 _4121_ (.X(_1740_),
    .A(net485),
    .B(net754),
    .C(net658));
 sg13g2_a21oi_1 _4122_ (.A1(net754),
    .A2(net658),
    .Y(_1741_),
    .B1(net485));
 sg13g2_nor3_1 _4123_ (.A(_1739_),
    .B(_1740_),
    .C(_1741_),
    .Y(_0224_));
 sg13g2_nand2_1 _4124_ (.Y(_1742_),
    .A(net527),
    .B(net665));
 sg13g2_nand3_1 _4125_ (.B(\pwm_module.counter0[1] ),
    .C(net754),
    .A(\pwm_module.counter0[2] ),
    .Y(_1743_));
 sg13g2_a21o_1 _4126_ (.A2(net754),
    .A1(net485),
    .B1(\pwm_module.counter0[2] ),
    .X(_1744_));
 sg13g2_nand2_1 _4127_ (.Y(_1745_),
    .A(_1743_),
    .B(_1744_));
 sg13g2_o21ai_1 _4128_ (.B1(_1742_),
    .Y(_0225_),
    .A1(net653),
    .A2(_1745_));
 sg13g2_nand2_1 _4129_ (.Y(_1746_),
    .A(net60),
    .B(net665));
 sg13g2_xnor2_1 _4130_ (.Y(_1747_),
    .A(_0163_),
    .B(_1743_));
 sg13g2_o21ai_1 _4131_ (.B1(_1746_),
    .Y(_0226_),
    .A1(net653),
    .A2(_1747_));
 sg13g2_and4_2 _4132_ (.A(\pwm_module.counter0[2] ),
    .B(\pwm_module.counter0[1] ),
    .C(net754),
    .D(net60),
    .X(_1748_));
 sg13g2_and3_1 _4133_ (.X(_1749_),
    .A(net102),
    .B(net658),
    .C(_1748_));
 sg13g2_a21oi_1 _4134_ (.A1(net658),
    .A2(_1748_),
    .Y(_1750_),
    .B1(net102));
 sg13g2_nand2_1 _4135_ (.Y(_1751_),
    .A(net102),
    .B(_1748_));
 sg13g2_nor3_1 _4136_ (.A(_1739_),
    .B(_1749_),
    .C(_1750_),
    .Y(_0227_));
 sg13g2_nand2_1 _4137_ (.Y(_1752_),
    .A(net252),
    .B(net665));
 sg13g2_xnor2_1 _4138_ (.Y(_1753_),
    .A(_0161_),
    .B(_1751_));
 sg13g2_o21ai_1 _4139_ (.B1(_1752_),
    .Y(_0228_),
    .A1(net654),
    .A2(_1753_));
 sg13g2_nand2_1 _4140_ (.Y(_1754_),
    .A(net290),
    .B(net665));
 sg13g2_nand3_1 _4141_ (.B(\pwm_module.counter0[4] ),
    .C(_1748_),
    .A(\pwm_module.counter0[5] ),
    .Y(_1755_));
 sg13g2_nor2_1 _4142_ (.A(_0160_),
    .B(_1755_),
    .Y(_1756_));
 sg13g2_xnor2_1 _4143_ (.Y(_1757_),
    .A(_0160_),
    .B(_1755_));
 sg13g2_o21ai_1 _4144_ (.B1(_1754_),
    .Y(_0229_),
    .A1(net654),
    .A2(_1757_));
 sg13g2_nand2_1 _4145_ (.Y(_1758_),
    .A(net265),
    .B(net665));
 sg13g2_xor2_1 _4146_ (.B(_1756_),
    .A(_0159_),
    .X(_1759_));
 sg13g2_o21ai_1 _4147_ (.B1(_1758_),
    .Y(_0230_),
    .A1(net653),
    .A2(_1759_));
 sg13g2_nand2_1 _4148_ (.Y(_1760_),
    .A(\pwm_module.counter0[6] ),
    .B(\pwm_module.counter0[7] ));
 sg13g2_nor2_1 _4149_ (.A(_1755_),
    .B(_1760_),
    .Y(_1761_));
 sg13g2_and3_1 _4150_ (.X(_1762_),
    .A(net494),
    .B(net659),
    .C(_1761_));
 sg13g2_a21oi_1 _4151_ (.A1(net659),
    .A2(_1761_),
    .Y(_1763_),
    .B1(net494));
 sg13g2_and2_1 _4152_ (.A(\pwm_module.counter0[8] ),
    .B(_1761_),
    .X(_1764_));
 sg13g2_nor3_1 _4153_ (.A(_1739_),
    .B(_1762_),
    .C(_1763_),
    .Y(_0231_));
 sg13g2_nand2_1 _4154_ (.Y(_1765_),
    .A(net367),
    .B(net665));
 sg13g2_xor2_1 _4155_ (.B(_1764_),
    .A(_0158_),
    .X(_1766_));
 sg13g2_o21ai_1 _4156_ (.B1(_1765_),
    .Y(_0232_),
    .A1(net654),
    .A2(_1766_));
 sg13g2_nand2_1 _4157_ (.Y(_1767_),
    .A(net455),
    .B(net666));
 sg13g2_nand2_1 _4158_ (.Y(_1768_),
    .A(\pwm_module.counter0[9] ),
    .B(\pwm_module.counter0[8] ));
 sg13g2_or3_1 _4159_ (.A(_1755_),
    .B(_1760_),
    .C(_1768_),
    .X(_1769_));
 sg13g2_nor2_1 _4160_ (.A(_0157_),
    .B(_1769_),
    .Y(_1770_));
 sg13g2_xnor2_1 _4161_ (.Y(_1771_),
    .A(_0157_),
    .B(_1769_));
 sg13g2_o21ai_1 _4162_ (.B1(_1767_),
    .Y(_0233_),
    .A1(net653),
    .A2(_1771_));
 sg13g2_nand2_1 _4163_ (.Y(_1772_),
    .A(net97),
    .B(net666));
 sg13g2_xor2_1 _4164_ (.B(_1770_),
    .A(_0156_),
    .X(_1773_));
 sg13g2_o21ai_1 _4165_ (.B1(_1772_),
    .Y(_0234_),
    .A1(net653),
    .A2(_1773_));
 sg13g2_nand2_1 _4166_ (.Y(_1774_),
    .A(\pwm_module.counter0[12] ),
    .B(net666));
 sg13g2_nand2_1 _4167_ (.Y(_1775_),
    .A(\pwm_module.counter0[10] ),
    .B(net97));
 sg13g2_nand4_1 _4168_ (.B(\pwm_module.counter0[9] ),
    .C(net97),
    .A(\pwm_module.counter0[10] ),
    .Y(_1776_),
    .D(_1764_));
 sg13g2_nor2_1 _4169_ (.A(net198),
    .B(_1776_),
    .Y(_1777_));
 sg13g2_xnor2_1 _4170_ (.Y(_1778_),
    .A(net198),
    .B(_1776_));
 sg13g2_o21ai_1 _4171_ (.B1(_1774_),
    .Y(_0235_),
    .A1(net653),
    .A2(_1778_));
 sg13g2_nand2_1 _4172_ (.Y(_1779_),
    .A(net434),
    .B(net666));
 sg13g2_xor2_1 _4173_ (.B(_1777_),
    .A(_0154_),
    .X(_1780_));
 sg13g2_o21ai_1 _4174_ (.B1(_1779_),
    .Y(_0236_),
    .A1(net653),
    .A2(_1780_));
 sg13g2_nand2_1 _4175_ (.Y(_1781_),
    .A(net434),
    .B(\pwm_module.counter0[12] ));
 sg13g2_or3_1 _4176_ (.A(net666),
    .B(_1776_),
    .C(_1781_),
    .X(_1782_));
 sg13g2_nor4_2 _4177_ (.A(_2353_),
    .B(_1769_),
    .C(_1775_),
    .Y(_1783_),
    .D(_1781_));
 sg13g2_a221oi_1 _4178_ (.B2(net658),
    .C1(_1739_),
    .B1(_1783_),
    .A1(_2353_),
    .Y(_0237_),
    .A2(_1782_));
 sg13g2_nand2_1 _4179_ (.Y(_1784_),
    .A(net70),
    .B(net665));
 sg13g2_xor2_1 _4180_ (.B(_1783_),
    .A(_0153_),
    .X(_1785_));
 sg13g2_o21ai_1 _4181_ (.B1(_1784_),
    .Y(_0238_),
    .A1(net654),
    .A2(_1785_));
 sg13g2_nand2_2 _4182_ (.Y(_1786_),
    .A(net70),
    .B(_1783_));
 sg13g2_nand2b_1 _4183_ (.Y(_1787_),
    .B(net658),
    .A_N(_1786_));
 sg13g2_nor2_1 _4184_ (.A(_2352_),
    .B(_1786_),
    .Y(_1788_));
 sg13g2_a221oi_1 _4185_ (.B2(net658),
    .C1(_1739_),
    .B1(_1788_),
    .A1(_2352_),
    .Y(_0239_),
    .A2(_1787_));
 sg13g2_nand2_1 _4186_ (.Y(_1789_),
    .A(net247),
    .B(net668));
 sg13g2_xor2_1 _4187_ (.B(_1788_),
    .A(_0152_),
    .X(_1790_));
 sg13g2_o21ai_1 _4188_ (.B1(_1789_),
    .Y(_0240_),
    .A1(net655),
    .A2(_1790_));
 sg13g2_nor3_1 _4189_ (.A(_2352_),
    .B(_2389_),
    .C(_1786_),
    .Y(_1791_));
 sg13g2_a21oi_1 _4190_ (.A1(net658),
    .A2(_1791_),
    .Y(_1792_),
    .B1(net479));
 sg13g2_nand2_1 _4191_ (.Y(_1793_),
    .A(\pwm_module.counter0[18] ),
    .B(_1791_));
 sg13g2_nor2_1 _4192_ (.A(net668),
    .B(_1793_),
    .Y(_1794_));
 sg13g2_nor3_1 _4193_ (.A(_1739_),
    .B(net480),
    .C(_1794_),
    .Y(_0241_));
 sg13g2_nand2_1 _4194_ (.Y(_1795_),
    .A(net52),
    .B(net667));
 sg13g2_xnor2_1 _4195_ (.Y(_1796_),
    .A(_0151_),
    .B(_1793_));
 sg13g2_o21ai_1 _4196_ (.B1(_1795_),
    .Y(_0242_),
    .A1(net655),
    .A2(_1796_));
 sg13g2_nand2_1 _4197_ (.Y(_1797_),
    .A(\pwm_module.counter0[20] ),
    .B(net667));
 sg13g2_nand4_1 _4198_ (.B(net525),
    .C(net52),
    .A(\pwm_module.counter0[18] ),
    .Y(_1798_),
    .D(\pwm_module.counter0[17] ));
 sg13g2_nor2_1 _4199_ (.A(_1786_),
    .B(_1798_),
    .Y(_1799_));
 sg13g2_or2_2 _4200_ (.X(_1800_),
    .B(_1798_),
    .A(_1786_));
 sg13g2_nor2_1 _4201_ (.A(net236),
    .B(_1800_),
    .Y(_1801_));
 sg13g2_xnor2_1 _4202_ (.Y(_1802_),
    .A(net236),
    .B(_1800_));
 sg13g2_o21ai_1 _4203_ (.B1(_1797_),
    .Y(_0243_),
    .A1(net655),
    .A2(_1802_));
 sg13g2_nand2_1 _4204_ (.Y(_1803_),
    .A(net425),
    .B(net667));
 sg13g2_xor2_1 _4205_ (.B(_1801_),
    .A(_0149_),
    .X(_1804_));
 sg13g2_o21ai_1 _4206_ (.B1(_1803_),
    .Y(_0244_),
    .A1(net655),
    .A2(_1804_));
 sg13g2_nand4_1 _4207_ (.B(net534),
    .C(net659),
    .A(net425),
    .Y(_1805_),
    .D(_1799_));
 sg13g2_nand3_1 _4208_ (.B(\pwm_module.counter0[21] ),
    .C(\pwm_module.counter0[20] ),
    .A(\pwm_module.counter0[22] ),
    .Y(_1806_));
 sg13g2_nor2_1 _4209_ (.A(_1800_),
    .B(_1806_),
    .Y(_1807_));
 sg13g2_a221oi_1 _4210_ (.B2(net662),
    .C1(_1739_),
    .B1(_1807_),
    .A1(_2351_),
    .Y(_0245_),
    .A2(net535));
 sg13g2_nand2_1 _4211_ (.Y(_1808_),
    .A(net50),
    .B(net667));
 sg13g2_xor2_1 _4212_ (.B(_1807_),
    .A(_0148_),
    .X(_1809_));
 sg13g2_o21ai_1 _4213_ (.B1(_1808_),
    .Y(_0246_),
    .A1(net655),
    .A2(_1809_));
 sg13g2_or3_1 _4214_ (.A(_2388_),
    .B(_1798_),
    .C(_1806_),
    .X(_1810_));
 sg13g2_nor2_1 _4215_ (.A(_1786_),
    .B(_1810_),
    .Y(_1811_));
 sg13g2_nand2_1 _4216_ (.Y(_1812_),
    .A(net662),
    .B(_1811_));
 sg13g2_nor4_2 _4217_ (.A(_2350_),
    .B(_2388_),
    .C(_1800_),
    .Y(_1813_),
    .D(_1806_));
 sg13g2_a221oi_1 _4218_ (.B2(net659),
    .C1(_1739_),
    .B1(_1813_),
    .A1(_2350_),
    .Y(_0247_),
    .A2(_1812_));
 sg13g2_nand2_1 _4219_ (.Y(_1814_),
    .A(net400),
    .B(net667));
 sg13g2_xor2_1 _4220_ (.B(_1813_),
    .A(_0147_),
    .X(_1815_));
 sg13g2_o21ai_1 _4221_ (.B1(_1814_),
    .Y(_0248_),
    .A1(_1737_),
    .A2(_1815_));
 sg13g2_nand3_1 _4222_ (.B(net400),
    .C(_1811_),
    .A(\pwm_module.counter0[24] ),
    .Y(_1816_));
 sg13g2_nand2b_1 _4223_ (.Y(_1817_),
    .B(net659),
    .A_N(_1816_));
 sg13g2_o21ai_1 _4224_ (.B1(_1736_),
    .Y(_1818_),
    .A1(_2349_),
    .A2(_1816_));
 sg13g2_a22oi_1 _4225_ (.Y(_0249_),
    .B1(_1818_),
    .B2(net659),
    .A2(_1817_),
    .A1(_2349_));
 sg13g2_nand2_1 _4226_ (.Y(_1819_),
    .A(net72),
    .B(net669));
 sg13g2_nand3_1 _4227_ (.B(\pwm_module.counter0[25] ),
    .C(_1813_),
    .A(\pwm_module.counter0[26] ),
    .Y(_1820_));
 sg13g2_xnor2_1 _4228_ (.Y(_1821_),
    .A(_0146_),
    .B(_1820_));
 sg13g2_o21ai_1 _4229_ (.B1(_1819_),
    .Y(_0250_),
    .A1(net655),
    .A2(_1821_));
 sg13g2_nand4_1 _4230_ (.B(\pwm_module.counter0[24] ),
    .C(net72),
    .A(\pwm_module.counter0[26] ),
    .Y(_1822_),
    .D(\pwm_module.counter0[25] ));
 sg13g2_nor3_2 _4231_ (.A(_1786_),
    .B(_1810_),
    .C(_1822_),
    .Y(_1823_));
 sg13g2_a21oi_1 _4232_ (.A1(net660),
    .A2(_1823_),
    .Y(_1824_),
    .B1(net537));
 sg13g2_nand2_1 _4233_ (.Y(_1825_),
    .A(\pwm_module.counter0[28] ),
    .B(_1823_));
 sg13g2_a21oi_1 _4234_ (.A1(_1736_),
    .A2(_1825_),
    .Y(_1826_),
    .B1(net668));
 sg13g2_nor2_1 _4235_ (.A(net538),
    .B(_1826_),
    .Y(_0251_));
 sg13g2_nand2_1 _4236_ (.Y(_1827_),
    .A(net326),
    .B(net669));
 sg13g2_xnor2_1 _4237_ (.Y(_1828_),
    .A(_0145_),
    .B(_1825_));
 sg13g2_o21ai_1 _4238_ (.B1(_1827_),
    .Y(_0252_),
    .A1(net655),
    .A2(_1828_));
 sg13g2_nand4_1 _4239_ (.B(net326),
    .C(net660),
    .A(\pwm_module.counter0[28] ),
    .Y(_1829_),
    .D(_1823_));
 sg13g2_nand4_1 _4240_ (.B(\pwm_module.counter0[28] ),
    .C(net326),
    .A(\pwm_module.counter0[30] ),
    .Y(_1830_),
    .D(_1823_));
 sg13g2_nand2_1 _4241_ (.Y(_1831_),
    .A(_1736_),
    .B(_1830_));
 sg13g2_a22oi_1 _4242_ (.Y(_0253_),
    .B1(_1831_),
    .B2(net660),
    .A2(_1829_),
    .A1(_2348_));
 sg13g2_nand2_1 _4243_ (.Y(_1832_),
    .A(net44),
    .B(net669));
 sg13g2_xnor2_1 _4244_ (.Y(_1833_),
    .A(_0167_),
    .B(_1830_));
 sg13g2_o21ai_1 _4245_ (.B1(_1832_),
    .Y(_0254_),
    .A1(net655),
    .A2(_1833_));
 sg13g2_mux2_1 _4246_ (.A0(net752),
    .A1(\spi_module.r_RX_Byte[0] ),
    .S(_0099_),
    .X(_0255_));
 sg13g2_nand2_1 _4247_ (.Y(_1834_),
    .A(\spi_module.r_RX_Byte[1] ),
    .B(_0099_));
 sg13g2_o21ai_1 _4248_ (.B1(_1834_),
    .Y(_0256_),
    .A1(net726),
    .A2(net718));
 sg13g2_nand2_1 _4249_ (.Y(_1835_),
    .A(\spi_module.r_RX_Byte[2] ),
    .B(_0099_));
 sg13g2_o21ai_1 _4250_ (.B1(_1835_),
    .Y(_0257_),
    .A1(net722),
    .A2(net718));
 sg13g2_mux2_1 _4251_ (.A0(net748),
    .A1(\spi_module.r_RX_Byte[3] ),
    .S(net718),
    .X(_0258_));
 sg13g2_mux2_1 _4252_ (.A0(net744),
    .A1(\spi_module.r_RX_Byte[4] ),
    .S(net718),
    .X(_0259_));
 sg13g2_mux2_1 _4253_ (.A0(net739),
    .A1(\spi_module.r_RX_Byte[5] ),
    .S(net718),
    .X(_0260_));
 sg13g2_mux2_1 _4254_ (.A0(net736),
    .A1(\spi_module.r_RX_Byte[6] ),
    .S(net718),
    .X(_0261_));
 sg13g2_mux2_1 _4255_ (.A0(net731),
    .A1(\spi_module.r_RX_Byte[7] ),
    .S(net718),
    .X(_0262_));
 sg13g2_mux2_1 _4256_ (.A0(net5),
    .A1(\spi_module.r_Temp_RX_Byte[0] ),
    .S(net764),
    .X(_0263_));
 sg13g2_mux2_1 _4257_ (.A0(\spi_module.r_Temp_RX_Byte[0] ),
    .A1(\spi_module.r_Temp_RX_Byte[1] ),
    .S(net764),
    .X(_0264_));
 sg13g2_mux2_1 _4258_ (.A0(\spi_module.r_Temp_RX_Byte[1] ),
    .A1(\spi_module.r_Temp_RX_Byte[2] ),
    .S(net764),
    .X(_0265_));
 sg13g2_mux2_1 _4259_ (.A0(\spi_module.r_Temp_RX_Byte[2] ),
    .A1(\spi_module.r_Temp_RX_Byte[3] ),
    .S(net763),
    .X(_0266_));
 sg13g2_mux2_1 _4260_ (.A0(\spi_module.r_Temp_RX_Byte[3] ),
    .A1(\spi_module.r_Temp_RX_Byte[4] ),
    .S(net763),
    .X(_0267_));
 sg13g2_mux2_1 _4261_ (.A0(\spi_module.r_Temp_RX_Byte[4] ),
    .A1(\spi_module.r_Temp_RX_Byte[5] ),
    .S(net763),
    .X(_0268_));
 sg13g2_mux2_1 _4262_ (.A0(\spi_module.r_Temp_RX_Byte[5] ),
    .A1(\spi_module.r_Temp_RX_Byte[6] ),
    .S(net763),
    .X(_0269_));
 sg13g2_nor2_2 _4263_ (.A(net764),
    .B(_2393_),
    .Y(_1836_));
 sg13g2_mux2_1 _4264_ (.A0(\spi_module.r_RX_Byte[0] ),
    .A1(net5),
    .S(_1836_),
    .X(_0270_));
 sg13g2_mux2_1 _4265_ (.A0(\spi_module.r_RX_Byte[1] ),
    .A1(\spi_module.r_Temp_RX_Byte[0] ),
    .S(_1836_),
    .X(_0271_));
 sg13g2_mux2_1 _4266_ (.A0(\spi_module.r_RX_Byte[2] ),
    .A1(\spi_module.r_Temp_RX_Byte[1] ),
    .S(_1836_),
    .X(_0272_));
 sg13g2_mux2_1 _4267_ (.A0(\spi_module.r_RX_Byte[3] ),
    .A1(\spi_module.r_Temp_RX_Byte[2] ),
    .S(_1836_),
    .X(_0273_));
 sg13g2_mux2_1 _4268_ (.A0(\spi_module.r_RX_Byte[4] ),
    .A1(\spi_module.r_Temp_RX_Byte[3] ),
    .S(_1836_),
    .X(_0274_));
 sg13g2_mux2_1 _4269_ (.A0(\spi_module.r_RX_Byte[5] ),
    .A1(\spi_module.r_Temp_RX_Byte[4] ),
    .S(_1836_),
    .X(_0275_));
 sg13g2_mux2_1 _4270_ (.A0(\spi_module.r_RX_Byte[6] ),
    .A1(\spi_module.r_Temp_RX_Byte[5] ),
    .S(_1836_),
    .X(_0276_));
 sg13g2_mux2_1 _4271_ (.A0(\spi_module.r_RX_Byte[7] ),
    .A1(\spi_module.r_Temp_RX_Byte[6] ),
    .S(_1836_),
    .X(_0277_));
 sg13g2_nor2_1 _4272_ (.A(\MemCell.curr_state[2] ),
    .B(_0898_),
    .Y(_1837_));
 sg13g2_nor2_1 _4273_ (.A(_0894_),
    .B(_1837_),
    .Y(_1838_));
 sg13g2_o21ai_1 _4274_ (.B1(\MemCell.o_RX_DV ),
    .Y(_1839_),
    .A1(_0894_),
    .A2(_1837_));
 sg13g2_nand3b_1 _4275_ (.B(_0899_),
    .C(\MemCell.o_RX_DV ),
    .Y(_1840_),
    .A_N(_1838_));
 sg13g2_nor2_2 _4276_ (.A(_0910_),
    .B(_1840_),
    .Y(_1841_));
 sg13g2_mux2_1 _4277_ (.A0(net215),
    .A1(net750),
    .S(net709),
    .X(_0279_));
 sg13g2_nor2_1 _4278_ (.A(net372),
    .B(net709),
    .Y(_1842_));
 sg13g2_a21oi_1 _4279_ (.A1(net724),
    .A2(net709),
    .Y(_0280_),
    .B1(_1842_));
 sg13g2_nor2_1 _4280_ (.A(net158),
    .B(_1841_),
    .Y(_1843_));
 sg13g2_a21oi_1 _4281_ (.A1(net720),
    .A2(_1841_),
    .Y(_0281_),
    .B1(_1843_));
 sg13g2_mux2_1 _4282_ (.A0(net361),
    .A1(net747),
    .S(net709),
    .X(_0282_));
 sg13g2_mux2_1 _4283_ (.A0(net146),
    .A1(net742),
    .S(net709),
    .X(_0283_));
 sg13g2_mux2_1 _4284_ (.A0(net131),
    .A1(net740),
    .S(net709),
    .X(_0284_));
 sg13g2_mux2_1 _4285_ (.A0(net175),
    .A1(net735),
    .S(net709),
    .X(_0285_));
 sg13g2_mux2_1 _4286_ (.A0(net154),
    .A1(net732),
    .S(net709),
    .X(_0286_));
 sg13g2_nand2b_2 _4287_ (.Y(_1844_),
    .B(\MemCell.counter[1] ),
    .A_N(net729));
 sg13g2_nand2_2 _4288_ (.Y(_1845_),
    .A(\MemCell.o_RX_DV ),
    .B(_0895_));
 sg13g2_nor2_2 _4289_ (.A(_1844_),
    .B(_1845_),
    .Y(_1846_));
 sg13g2_mux2_1 _4290_ (.A0(net133),
    .A1(net751),
    .S(net717),
    .X(_0287_));
 sg13g2_nor2_1 _4291_ (.A(net104),
    .B(net717),
    .Y(_1847_));
 sg13g2_a21oi_1 _4292_ (.A1(net725),
    .A2(net717),
    .Y(_0288_),
    .B1(_1847_));
 sg13g2_nor2_1 _4293_ (.A(net211),
    .B(net717),
    .Y(_1848_));
 sg13g2_a21oi_1 _4294_ (.A1(net721),
    .A2(net717),
    .Y(_0289_),
    .B1(_1848_));
 sg13g2_mux2_1 _4295_ (.A0(net189),
    .A1(net746),
    .S(net717),
    .X(_0290_));
 sg13g2_mux2_1 _4296_ (.A0(net116),
    .A1(net745),
    .S(_1846_),
    .X(_0291_));
 sg13g2_mux2_1 _4297_ (.A0(net137),
    .A1(net738),
    .S(_1846_),
    .X(_0292_));
 sg13g2_mux2_1 _4298_ (.A0(net164),
    .A1(net734),
    .S(net717),
    .X(_0293_));
 sg13g2_mux2_1 _4299_ (.A0(net136),
    .A1(net730),
    .S(net717),
    .X(_0294_));
 sg13g2_nor2_1 _4300_ (.A(_1840_),
    .B(_1844_),
    .Y(_1849_));
 sg13g2_mux2_1 _4301_ (.A0(net196),
    .A1(net752),
    .S(net708),
    .X(_0295_));
 sg13g2_nor2_1 _4302_ (.A(net322),
    .B(net708),
    .Y(_1850_));
 sg13g2_a21oi_1 _4303_ (.A1(net726),
    .A2(net708),
    .Y(_0296_),
    .B1(_1850_));
 sg13g2_nor2_1 _4304_ (.A(net155),
    .B(net708),
    .Y(_1851_));
 sg13g2_a21oi_1 _4305_ (.A1(net722),
    .A2(net708),
    .Y(_0297_),
    .B1(_1851_));
 sg13g2_mux2_1 _4306_ (.A0(net294),
    .A1(net748),
    .S(net708),
    .X(_0298_));
 sg13g2_mux2_1 _4307_ (.A0(net174),
    .A1(net743),
    .S(net708),
    .X(_0299_));
 sg13g2_mux2_1 _4308_ (.A0(net171),
    .A1(net739),
    .S(net708),
    .X(_0300_));
 sg13g2_mux2_1 _4309_ (.A0(net363),
    .A1(net735),
    .S(_1849_),
    .X(_0301_));
 sg13g2_mux2_1 _4310_ (.A0(net311),
    .A1(net732),
    .S(_1849_),
    .X(_0302_));
 sg13g2_nand2b_2 _4311_ (.Y(_1852_),
    .B(net729),
    .A_N(\MemCell.counter[1] ));
 sg13g2_nor2_2 _4312_ (.A(_1840_),
    .B(_1852_),
    .Y(_1853_));
 sg13g2_mux2_1 _4313_ (.A0(net287),
    .A1(net752),
    .S(_1853_),
    .X(_0303_));
 sg13g2_nor2_1 _4314_ (.A(net332),
    .B(net707),
    .Y(_1854_));
 sg13g2_a21oi_1 _4315_ (.A1(net726),
    .A2(net707),
    .Y(_0304_),
    .B1(_1854_));
 sg13g2_nor2_1 _4316_ (.A(net228),
    .B(net707),
    .Y(_1855_));
 sg13g2_a21oi_1 _4317_ (.A1(net722),
    .A2(net707),
    .Y(_0305_),
    .B1(_1855_));
 sg13g2_mux2_1 _4318_ (.A0(net119),
    .A1(net748),
    .S(net707),
    .X(_0306_));
 sg13g2_mux2_1 _4319_ (.A0(net203),
    .A1(net743),
    .S(_1853_),
    .X(_0307_));
 sg13g2_mux2_1 _4320_ (.A0(net262),
    .A1(net739),
    .S(net707),
    .X(_0308_));
 sg13g2_mux2_1 _4321_ (.A0(net177),
    .A1(net735),
    .S(net707),
    .X(_0309_));
 sg13g2_mux2_1 _4322_ (.A0(net170),
    .A1(net731),
    .S(net707),
    .X(_0310_));
 sg13g2_nor2_2 _4323_ (.A(net729),
    .B(\MemCell.counter[1] ),
    .Y(_1856_));
 sg13g2_nand2b_1 _4324_ (.Y(_1857_),
    .B(_1856_),
    .A_N(_1840_));
 sg13g2_mux2_1 _4325_ (.A0(net752),
    .A1(net362),
    .S(net706),
    .X(_0311_));
 sg13g2_nand2_1 _4326_ (.Y(_1858_),
    .A(net149),
    .B(_1857_));
 sg13g2_o21ai_1 _4327_ (.B1(_1858_),
    .Y(_0312_),
    .A1(net726),
    .A2(net706));
 sg13g2_nand2_1 _4328_ (.Y(_1859_),
    .A(net207),
    .B(_1857_));
 sg13g2_o21ai_1 _4329_ (.B1(_1859_),
    .Y(_0313_),
    .A1(net722),
    .A2(net706));
 sg13g2_mux2_1 _4330_ (.A0(net749),
    .A1(net355),
    .S(net706),
    .X(_0314_));
 sg13g2_mux2_1 _4331_ (.A0(net743),
    .A1(net419),
    .S(net706),
    .X(_0315_));
 sg13g2_mux2_1 _4332_ (.A0(net739),
    .A1(net364),
    .S(net706),
    .X(_0316_));
 sg13g2_mux2_1 _4333_ (.A0(net735),
    .A1(net330),
    .S(net706),
    .X(_0317_));
 sg13g2_mux2_1 _4334_ (.A0(net731),
    .A1(net374),
    .S(net706),
    .X(_0318_));
 sg13g2_nand2_2 _4335_ (.Y(_1860_),
    .A(\MemCell.o_RX_DV ),
    .B(_0893_));
 sg13g2_nor2_2 _4336_ (.A(_0910_),
    .B(_1860_),
    .Y(_1861_));
 sg13g2_mux2_1 _4337_ (.A0(net200),
    .A1(net750),
    .S(net716),
    .X(_0319_));
 sg13g2_nor2_1 _4338_ (.A(net105),
    .B(net716),
    .Y(_1862_));
 sg13g2_a21oi_1 _4339_ (.A1(net724),
    .A2(net716),
    .Y(_0320_),
    .B1(_1862_));
 sg13g2_nor2_1 _4340_ (.A(net256),
    .B(net716),
    .Y(_1863_));
 sg13g2_a21oi_1 _4341_ (.A1(net720),
    .A2(net716),
    .Y(_0321_),
    .B1(_1863_));
 sg13g2_mux2_1 _4342_ (.A0(net126),
    .A1(net747),
    .S(net716),
    .X(_0322_));
 sg13g2_mux2_1 _4343_ (.A0(net214),
    .A1(net742),
    .S(net716),
    .X(_0323_));
 sg13g2_mux2_1 _4344_ (.A0(net161),
    .A1(net738),
    .S(_1861_),
    .X(_0324_));
 sg13g2_mux2_1 _4345_ (.A0(net221),
    .A1(net734),
    .S(_1861_),
    .X(_0325_));
 sg13g2_mux2_1 _4346_ (.A0(net398),
    .A1(net730),
    .S(net716),
    .X(_0326_));
 sg13g2_nor2_2 _4347_ (.A(_1844_),
    .B(_1860_),
    .Y(_1864_));
 sg13g2_mux2_1 _4348_ (.A0(net151),
    .A1(net750),
    .S(net715),
    .X(_0327_));
 sg13g2_nor2_1 _4349_ (.A(net307),
    .B(net715),
    .Y(_1865_));
 sg13g2_a21oi_1 _4350_ (.A1(net724),
    .A2(net715),
    .Y(_0328_),
    .B1(_1865_));
 sg13g2_nor2_1 _4351_ (.A(net157),
    .B(net715),
    .Y(_1866_));
 sg13g2_a21oi_1 _4352_ (.A1(net720),
    .A2(net715),
    .Y(_0329_),
    .B1(_1866_));
 sg13g2_mux2_1 _4353_ (.A0(net115),
    .A1(net746),
    .S(net715),
    .X(_0330_));
 sg13g2_mux2_1 _4354_ (.A0(net225),
    .A1(net742),
    .S(_1864_),
    .X(_0331_));
 sg13g2_mux2_1 _4355_ (.A0(net346),
    .A1(net741),
    .S(net715),
    .X(_0332_));
 sg13g2_mux2_1 _4356_ (.A0(net232),
    .A1(net734),
    .S(_1864_),
    .X(_0333_));
 sg13g2_mux2_1 _4357_ (.A0(net278),
    .A1(net733),
    .S(net715),
    .X(_0334_));
 sg13g2_nor2_2 _4358_ (.A(_1852_),
    .B(_1860_),
    .Y(_1867_));
 sg13g2_mux2_1 _4359_ (.A0(net141),
    .A1(net750),
    .S(_1867_),
    .X(_0335_));
 sg13g2_nor2_1 _4360_ (.A(net370),
    .B(net714),
    .Y(_1868_));
 sg13g2_a21oi_1 _4361_ (.A1(net724),
    .A2(net714),
    .Y(_0336_),
    .B1(_1868_));
 sg13g2_nor2_1 _4362_ (.A(net114),
    .B(net714),
    .Y(_1869_));
 sg13g2_a21oi_1 _4363_ (.A1(net720),
    .A2(net714),
    .Y(_0337_),
    .B1(_1869_));
 sg13g2_mux2_1 _4364_ (.A0(net299),
    .A1(net746),
    .S(_1867_),
    .X(_0338_));
 sg13g2_mux2_1 _4365_ (.A0(net145),
    .A1(net742),
    .S(net714),
    .X(_0339_));
 sg13g2_mux2_1 _4366_ (.A0(net186),
    .A1(net738),
    .S(net714),
    .X(_0340_));
 sg13g2_mux2_1 _4367_ (.A0(net220),
    .A1(net734),
    .S(net714),
    .X(_0341_));
 sg13g2_mux2_1 _4368_ (.A0(net285),
    .A1(net730),
    .S(net714),
    .X(_0342_));
 sg13g2_nor3_2 _4369_ (.A(net729),
    .B(\MemCell.counter[1] ),
    .C(_1860_),
    .Y(_1870_));
 sg13g2_mux2_1 _4370_ (.A0(net139),
    .A1(net750),
    .S(net713),
    .X(_0343_));
 sg13g2_nor2_1 _4371_ (.A(net350),
    .B(net713),
    .Y(_1871_));
 sg13g2_a21oi_1 _4372_ (.A1(net724),
    .A2(net713),
    .Y(_0344_),
    .B1(_1871_));
 sg13g2_nor2_1 _4373_ (.A(net134),
    .B(net713),
    .Y(_1872_));
 sg13g2_a21oi_1 _4374_ (.A1(net720),
    .A2(net713),
    .Y(_0345_),
    .B1(_1872_));
 sg13g2_mux2_1 _4375_ (.A0(net239),
    .A1(net746),
    .S(net713),
    .X(_0346_));
 sg13g2_mux2_1 _4376_ (.A0(net358),
    .A1(net742),
    .S(_1870_),
    .X(_0347_));
 sg13g2_mux2_1 _4377_ (.A0(net169),
    .A1(net738),
    .S(_1870_),
    .X(_0348_));
 sg13g2_mux2_1 _4378_ (.A0(net241),
    .A1(net734),
    .S(net713),
    .X(_0349_));
 sg13g2_mux2_1 _4379_ (.A0(net259),
    .A1(net730),
    .S(net713),
    .X(_0350_));
 sg13g2_nor2_2 _4380_ (.A(_0902_),
    .B(_1839_),
    .Y(_1873_));
 sg13g2_nand2_2 _4381_ (.Y(_1874_),
    .A(_0909_),
    .B(_1873_));
 sg13g2_mux2_1 _4382_ (.A0(net752),
    .A1(net387),
    .S(net705),
    .X(_0351_));
 sg13g2_nand2_1 _4383_ (.Y(_1875_),
    .A(net310),
    .B(net705));
 sg13g2_o21ai_1 _4384_ (.B1(_1875_),
    .Y(_0352_),
    .A1(net726),
    .A2(net705));
 sg13g2_nand2_1 _4385_ (.Y(_1876_),
    .A(net224),
    .B(net705));
 sg13g2_o21ai_1 _4386_ (.B1(_1876_),
    .Y(_0353_),
    .A1(net722),
    .A2(net705));
 sg13g2_mux2_1 _4387_ (.A0(net748),
    .A1(net365),
    .S(net705),
    .X(_0354_));
 sg13g2_mux2_1 _4388_ (.A0(net743),
    .A1(net383),
    .S(net705),
    .X(_0355_));
 sg13g2_mux2_1 _4389_ (.A0(net740),
    .A1(net302),
    .S(_1874_),
    .X(_0356_));
 sg13g2_mux2_1 _4390_ (.A0(net735),
    .A1(net281),
    .S(_1874_),
    .X(_0357_));
 sg13g2_mux2_1 _4391_ (.A0(net731),
    .A1(net273),
    .S(net705),
    .X(_0358_));
 sg13g2_nand2b_2 _4392_ (.Y(_1877_),
    .B(_1873_),
    .A_N(_1844_));
 sg13g2_mux2_1 _4393_ (.A0(net752),
    .A1(net314),
    .S(net704),
    .X(_0359_));
 sg13g2_nand2_1 _4394_ (.Y(_1878_),
    .A(net321),
    .B(net704));
 sg13g2_o21ai_1 _4395_ (.B1(_1878_),
    .Y(_0360_),
    .A1(net726),
    .A2(net704));
 sg13g2_nand2_1 _4396_ (.Y(_1879_),
    .A(net74),
    .B(net704));
 sg13g2_o21ai_1 _4397_ (.B1(_1879_),
    .Y(_0361_),
    .A1(net722),
    .A2(net704));
 sg13g2_mux2_1 _4398_ (.A0(net748),
    .A1(net462),
    .S(net704),
    .X(_0362_));
 sg13g2_mux2_1 _4399_ (.A0(net743),
    .A1(net340),
    .S(_1877_),
    .X(_0363_));
 sg13g2_mux2_1 _4400_ (.A0(net740),
    .A1(net371),
    .S(_1877_),
    .X(_0364_));
 sg13g2_mux2_1 _4401_ (.A0(net736),
    .A1(net436),
    .S(net704),
    .X(_0365_));
 sg13g2_mux2_1 _4402_ (.A0(net731),
    .A1(net320),
    .S(net704),
    .X(_0366_));
 sg13g2_nor2_2 _4403_ (.A(_1845_),
    .B(_1852_),
    .Y(_1880_));
 sg13g2_nand2_1 _4404_ (.Y(_1881_),
    .A(net752),
    .B(net712));
 sg13g2_o21ai_1 _4405_ (.B1(_1881_),
    .Y(_0367_),
    .A1(_2372_),
    .A2(net712));
 sg13g2_nor2_1 _4406_ (.A(net99),
    .B(net712),
    .Y(_1882_));
 sg13g2_a21oi_1 _4407_ (.A1(net726),
    .A2(net712),
    .Y(_0368_),
    .B1(_1882_));
 sg13g2_nor2_1 _4408_ (.A(net150),
    .B(net712),
    .Y(_1883_));
 sg13g2_a21oi_1 _4409_ (.A1(net722),
    .A2(net712),
    .Y(_0369_),
    .B1(_1883_));
 sg13g2_mux2_1 _4410_ (.A0(net284),
    .A1(net748),
    .S(net712),
    .X(_0370_));
 sg13g2_mux2_1 _4411_ (.A0(net144),
    .A1(net743),
    .S(_1880_),
    .X(_0371_));
 sg13g2_mux2_1 _4412_ (.A0(net135),
    .A1(net739),
    .S(net712),
    .X(_0372_));
 sg13g2_mux2_1 _4413_ (.A0(net197),
    .A1(net735),
    .S(_1880_),
    .X(_0373_));
 sg13g2_mux2_1 _4414_ (.A0(net166),
    .A1(net731),
    .S(_1880_),
    .X(_0374_));
 sg13g2_nand2b_2 _4415_ (.Y(_1884_),
    .B(_1873_),
    .A_N(_1852_));
 sg13g2_mux2_1 _4416_ (.A0(net751),
    .A1(net335),
    .S(net703),
    .X(_0375_));
 sg13g2_nand2_1 _4417_ (.Y(_1885_),
    .A(net366),
    .B(net703));
 sg13g2_o21ai_1 _4418_ (.B1(_1885_),
    .Y(_0376_),
    .A1(net725),
    .A2(net703));
 sg13g2_nand2_1 _4419_ (.Y(_1886_),
    .A(net103),
    .B(net703));
 sg13g2_o21ai_1 _4420_ (.B1(_1886_),
    .Y(_0377_),
    .A1(net721),
    .A2(net703));
 sg13g2_mux2_1 _4421_ (.A0(net747),
    .A1(net471),
    .S(net703),
    .X(_0378_));
 sg13g2_mux2_1 _4422_ (.A0(net745),
    .A1(net437),
    .S(_1884_),
    .X(_0379_));
 sg13g2_mux2_1 _4423_ (.A0(net738),
    .A1(net433),
    .S(_1884_),
    .X(_0380_));
 sg13g2_mux2_1 _4424_ (.A0(net737),
    .A1(net395),
    .S(net703),
    .X(_0381_));
 sg13g2_mux2_1 _4425_ (.A0(net733),
    .A1(net348),
    .S(net703),
    .X(_0382_));
 sg13g2_nand2_2 _4426_ (.Y(_1887_),
    .A(_1856_),
    .B(_1873_));
 sg13g2_mux2_1 _4427_ (.A0(net750),
    .A1(net429),
    .S(net702),
    .X(_0383_));
 sg13g2_nand2_1 _4428_ (.Y(_1888_),
    .A(net108),
    .B(net702));
 sg13g2_o21ai_1 _4429_ (.B1(_1888_),
    .Y(_0384_),
    .A1(net724),
    .A2(net702));
 sg13g2_nand2_1 _4430_ (.Y(_1889_),
    .A(net183),
    .B(net702));
 sg13g2_o21ai_1 _4431_ (.B1(_1889_),
    .Y(_0385_),
    .A1(net720),
    .A2(net702));
 sg13g2_mux2_1 _4432_ (.A0(net747),
    .A1(net463),
    .S(net702),
    .X(_0386_));
 sg13g2_mux2_1 _4433_ (.A0(net742),
    .A1(net323),
    .S(_1887_),
    .X(_0387_));
 sg13g2_mux2_1 _4434_ (.A0(net738),
    .A1(net373),
    .S(_1887_),
    .X(_0388_));
 sg13g2_mux2_1 _4435_ (.A0(net734),
    .A1(net403),
    .S(net702),
    .X(_0389_));
 sg13g2_mux2_1 _4436_ (.A0(net730),
    .A1(net386),
    .S(net702),
    .X(_0390_));
 sg13g2_or3_2 _4437_ (.A(\MemCell.curr_state[1] ),
    .B(_0891_),
    .C(_1839_),
    .X(_1890_));
 sg13g2_nor2_2 _4438_ (.A(_0910_),
    .B(_1890_),
    .Y(_1891_));
 sg13g2_mux2_1 _4439_ (.A0(net282),
    .A1(net750),
    .S(net701),
    .X(_0391_));
 sg13g2_nor2_1 _4440_ (.A(net343),
    .B(net701),
    .Y(_1892_));
 sg13g2_a21oi_1 _4441_ (.A1(net724),
    .A2(net701),
    .Y(_0392_),
    .B1(_1892_));
 sg13g2_nor2_1 _4442_ (.A(net351),
    .B(net701),
    .Y(_1893_));
 sg13g2_a21oi_1 _4443_ (.A1(net721),
    .A2(net701),
    .Y(_0393_),
    .B1(_1893_));
 sg13g2_mux2_1 _4444_ (.A0(net249),
    .A1(net746),
    .S(net701),
    .X(_0394_));
 sg13g2_mux2_1 _4445_ (.A0(net156),
    .A1(net742),
    .S(_1891_),
    .X(_0395_));
 sg13g2_mux2_1 _4446_ (.A0(net208),
    .A1(net738),
    .S(_1891_),
    .X(_0396_));
 sg13g2_mux2_1 _4447_ (.A0(net298),
    .A1(net734),
    .S(net701),
    .X(_0397_));
 sg13g2_mux2_1 _4448_ (.A0(net132),
    .A1(net730),
    .S(net701),
    .X(_0398_));
 sg13g2_nor2_1 _4449_ (.A(_1844_),
    .B(_1890_),
    .Y(_1894_));
 sg13g2_mux2_1 _4450_ (.A0(net178),
    .A1(net751),
    .S(net700),
    .X(_0399_));
 sg13g2_nor2_1 _4451_ (.A(net409),
    .B(_1894_),
    .Y(_1895_));
 sg13g2_a21oi_1 _4452_ (.A1(net725),
    .A2(_1894_),
    .Y(_0400_),
    .B1(_1895_));
 sg13g2_nor2_1 _4453_ (.A(net176),
    .B(net700),
    .Y(_1896_));
 sg13g2_a21oi_1 _4454_ (.A1(net720),
    .A2(net700),
    .Y(_0401_),
    .B1(_1896_));
 sg13g2_mux2_1 _4455_ (.A0(net118),
    .A1(net746),
    .S(net700),
    .X(_0402_));
 sg13g2_mux2_1 _4456_ (.A0(net369),
    .A1(net743),
    .S(net700),
    .X(_0403_));
 sg13g2_mux2_1 _4457_ (.A0(net272),
    .A1(net740),
    .S(net700),
    .X(_0404_));
 sg13g2_mux2_1 _4458_ (.A0(net286),
    .A1(net735),
    .S(net700),
    .X(_0405_));
 sg13g2_mux2_1 _4459_ (.A0(net352),
    .A1(net732),
    .S(net700),
    .X(_0406_));
 sg13g2_nor2_2 _4460_ (.A(_1852_),
    .B(_1890_),
    .Y(_1897_));
 sg13g2_mux2_1 _4461_ (.A0(net172),
    .A1(net751),
    .S(net699),
    .X(_0407_));
 sg13g2_nor2_1 _4462_ (.A(net235),
    .B(net699),
    .Y(_1898_));
 sg13g2_a21oi_1 _4463_ (.A1(net725),
    .A2(net699),
    .Y(_0408_),
    .B1(_1898_));
 sg13g2_nor2_1 _4464_ (.A(net240),
    .B(net699),
    .Y(_1899_));
 sg13g2_a21oi_1 _4465_ (.A1(net721),
    .A2(net699),
    .Y(_0409_),
    .B1(_1899_));
 sg13g2_mux2_1 _4466_ (.A0(net399),
    .A1(net746),
    .S(net699),
    .X(_0410_));
 sg13g2_mux2_1 _4467_ (.A0(net138),
    .A1(net743),
    .S(_1897_),
    .X(_0411_));
 sg13g2_mux2_1 _4468_ (.A0(net264),
    .A1(net739),
    .S(_1897_),
    .X(_0412_));
 sg13g2_mux2_1 _4469_ (.A0(net269),
    .A1(net735),
    .S(net699),
    .X(_0413_));
 sg13g2_mux2_1 _4470_ (.A0(net539),
    .A1(net730),
    .S(net699),
    .X(_0414_));
 sg13g2_nor3_2 _4471_ (.A(\MemCell.counter[0] ),
    .B(\MemCell.counter[1] ),
    .C(_1890_),
    .Y(_1900_));
 sg13g2_mux2_1 _4472_ (.A0(net181),
    .A1(net752),
    .S(_1900_),
    .X(_0415_));
 sg13g2_nor2_1 _4473_ (.A(net296),
    .B(net698),
    .Y(_1901_));
 sg13g2_a21oi_1 _4474_ (.A1(net727),
    .A2(_1900_),
    .Y(_0416_),
    .B1(_1901_));
 sg13g2_nor2_1 _4475_ (.A(net201),
    .B(net698),
    .Y(_1902_));
 sg13g2_a21oi_1 _4476_ (.A1(net723),
    .A2(net698),
    .Y(_0417_),
    .B1(_1902_));
 sg13g2_mux2_1 _4477_ (.A0(net165),
    .A1(net748),
    .S(net698),
    .X(_0418_));
 sg13g2_mux2_1 _4478_ (.A0(net125),
    .A1(net744),
    .S(net698),
    .X(_0419_));
 sg13g2_mux2_1 _4479_ (.A0(net397),
    .A1(net739),
    .S(net698),
    .X(_0420_));
 sg13g2_mux2_1 _4480_ (.A0(net331),
    .A1(net736),
    .S(net698),
    .X(_0421_));
 sg13g2_mux2_1 _4481_ (.A0(net246),
    .A1(net731),
    .S(net698),
    .X(_0422_));
 sg13g2_o21ai_1 _4482_ (.B1(net421),
    .Y(_0423_),
    .A1(_2373_),
    .A2(_0903_));
 sg13g2_nor2b_1 _4483_ (.A(\MemCell.curr_state[2] ),
    .B_N(_0900_),
    .Y(_1903_));
 sg13g2_nor3_1 _4484_ (.A(_0897_),
    .B(_0899_),
    .C(_1903_),
    .Y(_1904_));
 sg13g2_nor2_1 _4485_ (.A(\MemCell.o_RX_DV ),
    .B(_1904_),
    .Y(_1905_));
 sg13g2_or2_1 _4486_ (.X(_1906_),
    .B(_1905_),
    .A(_1838_));
 sg13g2_nand2_1 _4487_ (.Y(_1907_),
    .A(net729),
    .B(_1905_));
 sg13g2_o21ai_1 _4488_ (.B1(_1907_),
    .Y(_0424_),
    .A1(net729),
    .A2(_1906_));
 sg13g2_nor3_1 _4489_ (.A(_0909_),
    .B(_1856_),
    .C(_1906_),
    .Y(_1908_));
 sg13g2_a21o_1 _4490_ (.A2(_1905_),
    .A1(net577),
    .B1(_1908_),
    .X(_0425_));
 sg13g2_nor2b_2 _4491_ (.A(_1845_),
    .B_N(_1856_),
    .Y(_1909_));
 sg13g2_mux2_1 _4492_ (.A0(net218),
    .A1(net753),
    .S(net711),
    .X(_0426_));
 sg13g2_nor2_1 _4493_ (.A(net315),
    .B(net711),
    .Y(_1910_));
 sg13g2_a21oi_1 _4494_ (.A1(net727),
    .A2(net711),
    .Y(_0427_),
    .B1(_1910_));
 sg13g2_nor2_1 _4495_ (.A(net288),
    .B(net711),
    .Y(_1911_));
 sg13g2_a21oi_1 _4496_ (.A1(net723),
    .A2(net711),
    .Y(_0428_),
    .B1(_1911_));
 sg13g2_mux2_1 _4497_ (.A0(net280),
    .A1(net748),
    .S(net711),
    .X(_0429_));
 sg13g2_mux2_1 _4498_ (.A0(net344),
    .A1(net744),
    .S(net711),
    .X(_0430_));
 sg13g2_mux2_1 _4499_ (.A0(net295),
    .A1(net739),
    .S(_1909_),
    .X(_0431_));
 sg13g2_mux2_1 _4500_ (.A0(net277),
    .A1(net736),
    .S(_1909_),
    .X(_0432_));
 sg13g2_mux2_1 _4501_ (.A0(net345),
    .A1(net731),
    .S(net711),
    .X(_0433_));
 sg13g2_nand2_1 _4502_ (.Y(_1912_),
    .A(_0124_),
    .B(_1587_));
 sg13g2_or2_1 _4503_ (.X(_1913_),
    .B(_1601_),
    .A(\pwm_module.counter2[28] ));
 sg13g2_a22oi_1 _4504_ (.Y(_1914_),
    .B1(_1591_),
    .B2(_0168_),
    .A2(_1589_),
    .A1(_2332_));
 sg13g2_nand3_1 _4505_ (.B(_1913_),
    .C(_1914_),
    .A(_1912_),
    .Y(_1915_));
 sg13g2_a22oi_1 _4506_ (.Y(_1916_),
    .B1(_1599_),
    .B2(_2331_),
    .A2(_1594_),
    .A1(\pwm_module.counter2[26] ));
 sg13g2_a22oi_1 _4507_ (.Y(_1917_),
    .B1(_1595_),
    .B2(_0125_),
    .A2(_1593_),
    .A1(_2330_));
 sg13g2_nand2b_1 _4508_ (.Y(_1918_),
    .B(_1917_),
    .A_N(_1916_));
 sg13g2_nand2_1 _4509_ (.Y(_1919_),
    .A(\pwm_module.counter2[28] ),
    .B(_1601_));
 sg13g2_or2_1 _4510_ (.X(_1920_),
    .B(_1595_),
    .A(_0125_));
 sg13g2_or2_1 _4511_ (.X(_1921_),
    .B(_1602_),
    .A(\pwm_module.counter2[24] ));
 sg13g2_nand2_1 _4512_ (.Y(_1922_),
    .A(_0126_),
    .B(_1598_));
 sg13g2_nand3_1 _4513_ (.B(_1921_),
    .C(_1922_),
    .A(_1917_),
    .Y(_1923_));
 sg13g2_and4_1 _4514_ (.A(_1918_),
    .B(_1919_),
    .C(_1920_),
    .D(_1923_),
    .X(_1924_));
 sg13g2_nor2_1 _4515_ (.A(_0168_),
    .B(_1591_),
    .Y(_1925_));
 sg13g2_nand2_1 _4516_ (.Y(_1926_),
    .A(\pwm_module.counter2[30] ),
    .B(_1590_));
 sg13g2_or2_1 _4517_ (.X(_1927_),
    .B(_1587_),
    .A(_0124_));
 sg13g2_nand2_1 _4518_ (.Y(_1928_),
    .A(_1926_),
    .B(_1927_));
 sg13g2_a21oi_1 _4519_ (.A1(_1914_),
    .A2(_1928_),
    .Y(_1929_),
    .B1(_1925_));
 sg13g2_o21ai_1 _4520_ (.B1(_1929_),
    .Y(_1930_),
    .A1(_1915_),
    .A2(_1924_));
 sg13g2_nand2_1 _4521_ (.Y(_1931_),
    .A(\pwm_module.counter2[24] ),
    .B(_1602_));
 sg13g2_nand3b_1 _4522_ (.B(_1931_),
    .C(_1916_),
    .Y(_1932_),
    .A_N(_1925_));
 sg13g2_nand4_1 _4523_ (.B(_1920_),
    .C(_1926_),
    .A(_1919_),
    .Y(_1933_),
    .D(_1927_));
 sg13g2_nor4_2 _4524_ (.A(_1915_),
    .B(_1923_),
    .C(_1932_),
    .Y(_1934_),
    .D(_1933_));
 sg13g2_a22oi_1 _4525_ (.Y(_1935_),
    .B1(_1624_),
    .B2(_2327_),
    .A2(_1622_),
    .A1(_0127_));
 sg13g2_a22oi_1 _4526_ (.Y(_1936_),
    .B1(_1631_),
    .B2(_0129_),
    .A2(_1616_),
    .A1(_0128_));
 sg13g2_a22oi_1 _4527_ (.Y(_1937_),
    .B1(_1625_),
    .B2(\pwm_module.counter2[22] ),
    .A2(_1617_),
    .A1(_2328_));
 sg13g2_nand2b_1 _4528_ (.Y(_1938_),
    .B(_1937_),
    .A_N(_1936_));
 sg13g2_a22oi_1 _4529_ (.Y(_1939_),
    .B1(_1935_),
    .B2(_1938_),
    .A2(_1623_),
    .A1(_2326_));
 sg13g2_nor2_1 _4530_ (.A(\pwm_module.counter2[18] ),
    .B(_1641_),
    .Y(_1940_));
 sg13g2_a21o_1 _4531_ (.A2(_1637_),
    .A1(_0130_),
    .B1(_1940_),
    .X(_1941_));
 sg13g2_nand3b_1 _4532_ (.B(\MemCell.counter_value[17] ),
    .C(_0131_),
    .Y(_1942_),
    .A_N(net792));
 sg13g2_o21ai_1 _4533_ (.B1(_1942_),
    .Y(_1943_),
    .A1(\pwm_module.counter2[16] ),
    .A2(_1619_));
 sg13g2_a22oi_1 _4534_ (.Y(_1944_),
    .B1(_1641_),
    .B2(\pwm_module.counter2[18] ),
    .A2(_1628_),
    .A1(_2324_));
 sg13g2_a221oi_1 _4535_ (.B2(_1944_),
    .C1(_1940_),
    .B1(_1943_),
    .A1(_0130_),
    .Y(_1945_),
    .A2(_1637_));
 sg13g2_a22oi_1 _4536_ (.Y(_1946_),
    .B1(_1632_),
    .B2(_2329_),
    .A2(_1623_),
    .A1(_2326_));
 sg13g2_nand4_1 _4537_ (.B(_1936_),
    .C(_1937_),
    .A(_1935_),
    .Y(_1947_),
    .D(_1946_));
 sg13g2_nor2_1 _4538_ (.A(_0130_),
    .B(_1637_),
    .Y(_1948_));
 sg13g2_nand2b_1 _4539_ (.Y(_1949_),
    .B(_1944_),
    .A_N(_1948_));
 sg13g2_nor3_1 _4540_ (.A(_1945_),
    .B(_1947_),
    .C(_1948_),
    .Y(_1950_));
 sg13g2_a22oi_1 _4541_ (.Y(_1951_),
    .B1(_1650_),
    .B2(_2321_),
    .A2(_1648_),
    .A1(_0132_));
 sg13g2_inv_1 _4542_ (.Y(_1952_),
    .A(_1951_));
 sg13g2_or2_1 _4543_ (.X(_1953_),
    .B(_1648_),
    .A(_0132_));
 sg13g2_nand2_1 _4544_ (.Y(_1954_),
    .A(\pwm_module.counter2[14] ),
    .B(_1651_));
 sg13g2_nor2_1 _4545_ (.A(_0133_),
    .B(_1655_),
    .Y(_1955_));
 sg13g2_nand3_1 _4546_ (.B(_1953_),
    .C(_1954_),
    .A(_1951_),
    .Y(_1956_));
 sg13g2_a22oi_1 _4547_ (.Y(_1957_),
    .B1(_1658_),
    .B2(_0134_),
    .A2(_1655_),
    .A1(_0133_));
 sg13g2_o21ai_1 _4548_ (.B1(_1957_),
    .Y(_1958_),
    .A1(_0134_),
    .A2(_1658_));
 sg13g2_nor3_1 _4549_ (.A(_1955_),
    .B(_1956_),
    .C(_1958_),
    .Y(_1959_));
 sg13g2_xnor2_1 _4550_ (.Y(_1960_),
    .A(_0136_),
    .B(_1660_));
 sg13g2_and2_1 _4551_ (.A(_0135_),
    .B(_1662_),
    .X(_1961_));
 sg13g2_nand2_1 _4552_ (.Y(_1962_),
    .A(_0135_),
    .B(_1662_));
 sg13g2_or2_1 _4553_ (.X(_1963_),
    .B(_1662_),
    .A(_0135_));
 sg13g2_or2_1 _4554_ (.X(_1964_),
    .B(_1666_),
    .A(_0137_));
 sg13g2_nand4_1 _4555_ (.B(_1962_),
    .C(_1963_),
    .A(_1960_),
    .Y(_1965_),
    .D(_1964_));
 sg13g2_and2_1 _4556_ (.A(\pwm_module.counter2[8] ),
    .B(_1668_),
    .X(_1966_));
 sg13g2_nor2_1 _4557_ (.A(\pwm_module.counter2[8] ),
    .B(_1668_),
    .Y(_1967_));
 sg13g2_a21oi_1 _4558_ (.A1(_0137_),
    .A2(_1666_),
    .Y(_1968_),
    .B1(_1967_));
 sg13g2_nor4_1 _4559_ (.A(_1955_),
    .B(_1956_),
    .C(_1958_),
    .D(_1966_),
    .Y(_1969_));
 sg13g2_nand3b_1 _4560_ (.B(_1968_),
    .C(_1969_),
    .Y(_1970_),
    .A_N(_1965_));
 sg13g2_nor2_1 _4561_ (.A(\pwm_module.counter2[2] ),
    .B(_1693_),
    .Y(_1971_));
 sg13g2_a21oi_1 _4562_ (.A1(_0142_),
    .A2(_1691_),
    .Y(_1972_),
    .B1(_1971_));
 sg13g2_and2_1 _4563_ (.A(\pwm_module.counter2[2] ),
    .B(_1693_),
    .X(_1973_));
 sg13g2_nor2_1 _4564_ (.A(\pwm_module.counter2[1] ),
    .B(_1695_),
    .Y(_1974_));
 sg13g2_and2_1 _4565_ (.A(\pwm_module.counter2[1] ),
    .B(_1695_),
    .X(_1975_));
 sg13g2_nand2_1 _4566_ (.Y(_1976_),
    .A(\pwm_module.counter2[1] ),
    .B(_1695_));
 sg13g2_nand2_1 _4567_ (.Y(_1977_),
    .A(\pwm_module.counter2[0] ),
    .B(_1698_));
 sg13g2_nand2b_1 _4568_ (.Y(_1978_),
    .B(_1977_),
    .A_N(_1974_));
 sg13g2_a21oi_1 _4569_ (.A1(_1976_),
    .A2(_1977_),
    .Y(_1979_),
    .B1(_1974_));
 sg13g2_o21ai_1 _4570_ (.B1(_1972_),
    .Y(_1980_),
    .A1(_1973_),
    .A2(_1979_));
 sg13g2_a22oi_1 _4571_ (.Y(_1981_),
    .B1(_1686_),
    .B2(\pwm_module.counter2[5] ),
    .A2(_1683_),
    .A1(_0139_));
 sg13g2_nand2b_1 _4572_ (.Y(_1982_),
    .B(_1682_),
    .A_N(_0139_));
 sg13g2_nand2_1 _4573_ (.Y(_1983_),
    .A(\pwm_module.counter2[7] ),
    .B(_1680_));
 sg13g2_or2_1 _4574_ (.X(_1984_),
    .B(_1680_),
    .A(\pwm_module.counter2[7] ));
 sg13g2_nand4_1 _4575_ (.B(_1982_),
    .C(_1983_),
    .A(_1981_),
    .Y(_1985_),
    .D(_1984_));
 sg13g2_a22oi_1 _4576_ (.Y(_1986_),
    .B1(_1690_),
    .B2(_2320_),
    .A2(_1687_),
    .A1(_2319_));
 sg13g2_nand2b_1 _4577_ (.Y(_1987_),
    .B(\pwm_module.counter2[4] ),
    .A_N(_1690_));
 sg13g2_or2_1 _4578_ (.X(_1988_),
    .B(_1691_),
    .A(_0142_));
 sg13g2_nand3_1 _4579_ (.B(_1987_),
    .C(_1988_),
    .A(_1986_),
    .Y(_1989_));
 sg13g2_nand2_1 _4580_ (.Y(_1990_),
    .A(_1986_),
    .B(_1987_));
 sg13g2_nor2_1 _4581_ (.A(_1985_),
    .B(_1989_),
    .Y(_1991_));
 sg13g2_nor2_1 _4582_ (.A(_1985_),
    .B(_1986_),
    .Y(_1992_));
 sg13g2_o21ai_1 _4583_ (.B1(_1984_),
    .Y(_1993_),
    .A1(\pwm_module.counter2[6] ),
    .A2(_1682_));
 sg13g2_a221oi_1 _4584_ (.B2(_1983_),
    .C1(_1992_),
    .B1(_1993_),
    .A1(_1980_),
    .Y(_1994_),
    .A2(_1991_));
 sg13g2_nor2_1 _4585_ (.A(\pwm_module.counter2[10] ),
    .B(_1660_),
    .Y(_1995_));
 sg13g2_a21oi_1 _4586_ (.A1(_1963_),
    .A2(_1995_),
    .Y(_1996_),
    .B1(_1961_));
 sg13g2_o21ai_1 _4587_ (.B1(_1996_),
    .Y(_1997_),
    .A1(_1965_),
    .A2(_1968_));
 sg13g2_nor3_1 _4588_ (.A(_1955_),
    .B(_1956_),
    .C(_1957_),
    .Y(_1998_));
 sg13g2_a221oi_1 _4589_ (.B2(_1997_),
    .C1(_1998_),
    .B1(_1959_),
    .A1(_1952_),
    .Y(_1999_),
    .A2(_1953_));
 sg13g2_o21ai_1 _4590_ (.B1(_1999_),
    .Y(_2000_),
    .A1(_1970_),
    .A2(_1994_));
 sg13g2_a21o_1 _4591_ (.A2(_1619_),
    .A1(\pwm_module.counter2[16] ),
    .B1(_1943_),
    .X(_2001_));
 sg13g2_nor4_1 _4592_ (.A(_1941_),
    .B(_1947_),
    .C(_1949_),
    .D(_2001_),
    .Y(_2002_));
 sg13g2_o21ai_1 _4593_ (.B1(_1934_),
    .Y(_2003_),
    .A1(_1939_),
    .A2(_1950_));
 sg13g2_and2_1 _4594_ (.A(_1934_),
    .B(_2002_),
    .X(_2004_));
 sg13g2_nand2_1 _4595_ (.Y(_2005_),
    .A(_1930_),
    .B(_2003_));
 sg13g2_a21oi_1 _4596_ (.A1(_2000_),
    .A2(_2004_),
    .Y(_2006_),
    .B1(_2005_));
 sg13g2_o21ai_1 _4597_ (.B1(_1988_),
    .Y(_2007_),
    .A1(\pwm_module.counter2[0] ),
    .A2(_1698_));
 sg13g2_nor2_1 _4598_ (.A(_1973_),
    .B(_2007_),
    .Y(_2008_));
 sg13g2_nor4_1 _4599_ (.A(_1975_),
    .B(_1978_),
    .C(_1985_),
    .D(_1990_),
    .Y(_2009_));
 sg13g2_nand4_1 _4600_ (.B(_2004_),
    .C(_2008_),
    .A(_1972_),
    .Y(_2010_),
    .D(_2009_));
 sg13g2_o21ai_1 _4601_ (.B1(_2396_),
    .Y(_2011_),
    .A1(_1970_),
    .A2(_2010_));
 sg13g2_nor2_2 _4602_ (.A(_2006_),
    .B(_2011_),
    .Y(_2012_));
 sg13g2_nand2b_1 _4603_ (.Y(_2013_),
    .B(_2012_),
    .A_N(net685));
 sg13g2_nor2_1 _4604_ (.A(_2317_),
    .B(net688),
    .Y(_2014_));
 sg13g2_a21oi_1 _4605_ (.A1(_2317_),
    .A2(net652),
    .Y(_0434_),
    .B1(_2014_));
 sg13g2_nor2_2 _4606_ (.A(net680),
    .B(_2012_),
    .Y(_2015_));
 sg13g2_nand3b_1 _4607_ (.B(\pwm_module.counter2[1] ),
    .C(\pwm_module.counter2[0] ),
    .Y(_2016_),
    .A_N(net688));
 sg13g2_xnor2_1 _4608_ (.Y(_2017_),
    .A(net495),
    .B(_2014_));
 sg13g2_nor2_1 _4609_ (.A(_2015_),
    .B(net496),
    .Y(_0435_));
 sg13g2_xnor2_1 _4610_ (.Y(_2018_),
    .A(net573),
    .B(_2016_));
 sg13g2_nand3_1 _4611_ (.B(\pwm_module.counter2[1] ),
    .C(\pwm_module.counter2[2] ),
    .A(\pwm_module.counter2[0] ),
    .Y(_2019_));
 sg13g2_nor2b_1 _4612_ (.A(_2015_),
    .B_N(net574),
    .Y(_0436_));
 sg13g2_nand2_1 _4613_ (.Y(_2020_),
    .A(net75),
    .B(net688));
 sg13g2_xnor2_1 _4614_ (.Y(_2021_),
    .A(_0142_),
    .B(_2019_));
 sg13g2_o21ai_1 _4615_ (.B1(_2020_),
    .Y(_0437_),
    .A1(net651),
    .A2(_2021_));
 sg13g2_and4_1 _4616_ (.A(\pwm_module.counter2[0] ),
    .B(\pwm_module.counter2[1] ),
    .C(\pwm_module.counter2[3] ),
    .D(\pwm_module.counter2[2] ),
    .X(_2022_));
 sg13g2_nor2b_1 _4617_ (.A(net688),
    .B_N(_2022_),
    .Y(_2023_));
 sg13g2_xnor2_1 _4618_ (.Y(_2024_),
    .A(net470),
    .B(_2023_));
 sg13g2_nand2_1 _4619_ (.Y(_2025_),
    .A(\pwm_module.counter2[4] ),
    .B(_2022_));
 sg13g2_nor2_1 _4620_ (.A(_2015_),
    .B(_2024_),
    .Y(_0438_));
 sg13g2_nand2_1 _4621_ (.Y(_2026_),
    .A(net341),
    .B(net688));
 sg13g2_xnor2_1 _4622_ (.Y(_2027_),
    .A(_0140_),
    .B(_2025_));
 sg13g2_o21ai_1 _4623_ (.B1(_2026_),
    .Y(_0439_),
    .A1(net651),
    .A2(_2027_));
 sg13g2_nand2_1 _4624_ (.Y(_2028_),
    .A(net260),
    .B(net687));
 sg13g2_nand3_1 _4625_ (.B(\pwm_module.counter2[4] ),
    .C(_2022_),
    .A(\pwm_module.counter2[5] ),
    .Y(_2029_));
 sg13g2_nor2_1 _4626_ (.A(_0139_),
    .B(_2029_),
    .Y(_2030_));
 sg13g2_xnor2_1 _4627_ (.Y(_2031_),
    .A(_0139_),
    .B(_2029_));
 sg13g2_o21ai_1 _4628_ (.B1(_2028_),
    .Y(_0440_),
    .A1(net651),
    .A2(_2031_));
 sg13g2_nand2_1 _4629_ (.Y(_2032_),
    .A(net216),
    .B(net687));
 sg13g2_xor2_1 _4630_ (.B(_2030_),
    .A(_0138_),
    .X(_2033_));
 sg13g2_o21ai_1 _4631_ (.B1(_2032_),
    .Y(_0441_),
    .A1(net651),
    .A2(_2033_));
 sg13g2_nand2_2 _4632_ (.Y(_2034_),
    .A(\pwm_module.counter2[7] ),
    .B(\pwm_module.counter2[6] ));
 sg13g2_nor2_2 _4633_ (.A(_2029_),
    .B(_2034_),
    .Y(_2035_));
 sg13g2_nor2b_1 _4634_ (.A(net686),
    .B_N(_2035_),
    .Y(_2036_));
 sg13g2_xnor2_1 _4635_ (.Y(_2037_),
    .A(net531),
    .B(_2036_));
 sg13g2_nand2_1 _4636_ (.Y(_2038_),
    .A(\pwm_module.counter2[8] ),
    .B(_2035_));
 sg13g2_nor2_1 _4637_ (.A(_2015_),
    .B(_2037_),
    .Y(_0442_));
 sg13g2_nand2_1 _4638_ (.Y(_2039_),
    .A(net147),
    .B(net686));
 sg13g2_xnor2_1 _4639_ (.Y(_2040_),
    .A(_0137_),
    .B(_2038_));
 sg13g2_o21ai_1 _4640_ (.B1(_2039_),
    .Y(_0443_),
    .A1(net651),
    .A2(_2040_));
 sg13g2_nand2_1 _4641_ (.Y(_2041_),
    .A(net300),
    .B(net686));
 sg13g2_nand3_1 _4642_ (.B(\pwm_module.counter2[8] ),
    .C(_2035_),
    .A(net147),
    .Y(_2042_));
 sg13g2_nor2_1 _4643_ (.A(_0136_),
    .B(_2042_),
    .Y(_2043_));
 sg13g2_xnor2_1 _4644_ (.Y(_2044_),
    .A(_0136_),
    .B(_2042_));
 sg13g2_o21ai_1 _4645_ (.B1(_2041_),
    .Y(_0444_),
    .A1(net652),
    .A2(_2044_));
 sg13g2_nand2_1 _4646_ (.Y(_2045_),
    .A(net77),
    .B(net686));
 sg13g2_xor2_1 _4647_ (.B(_2043_),
    .A(_0135_),
    .X(_2046_));
 sg13g2_o21ai_1 _4648_ (.B1(_2045_),
    .Y(_0445_),
    .A1(net652),
    .A2(_2046_));
 sg13g2_nand2_1 _4649_ (.Y(_2047_),
    .A(net93),
    .B(net687));
 sg13g2_nand4_1 _4650_ (.B(\pwm_module.counter2[10] ),
    .C(\pwm_module.counter2[9] ),
    .A(net77),
    .Y(_2048_),
    .D(\pwm_module.counter2[8] ));
 sg13g2_nor3_1 _4651_ (.A(_2029_),
    .B(_2034_),
    .C(_2048_),
    .Y(_2049_));
 sg13g2_nand2b_1 _4652_ (.Y(_2050_),
    .B(_2049_),
    .A_N(_0134_));
 sg13g2_xor2_1 _4653_ (.B(_2049_),
    .A(_0134_),
    .X(_2051_));
 sg13g2_o21ai_1 _4654_ (.B1(_2047_),
    .Y(_0446_),
    .A1(net651),
    .A2(_2051_));
 sg13g2_nand2_1 _4655_ (.Y(_2052_),
    .A(net127),
    .B(net687));
 sg13g2_xnor2_1 _4656_ (.Y(_2053_),
    .A(_0133_),
    .B(_2050_));
 sg13g2_o21ai_1 _4657_ (.B1(_2052_),
    .Y(_0447_),
    .A1(net651),
    .A2(_2053_));
 sg13g2_nand2_1 _4658_ (.Y(_2054_),
    .A(\pwm_module.counter2[13] ),
    .B(\pwm_module.counter2[12] ));
 sg13g2_nor4_2 _4659_ (.A(_2029_),
    .B(_2034_),
    .C(_2048_),
    .Y(_2055_),
    .D(_2054_));
 sg13g2_nor2b_1 _4660_ (.A(net686),
    .B_N(_2055_),
    .Y(_2056_));
 sg13g2_xnor2_1 _4661_ (.Y(_2057_),
    .A(net520),
    .B(_2056_));
 sg13g2_and2_1 _4662_ (.A(\pwm_module.counter2[14] ),
    .B(_2055_),
    .X(_2058_));
 sg13g2_nor2_1 _4663_ (.A(_2015_),
    .B(net521),
    .Y(_0448_));
 sg13g2_nand2_1 _4664_ (.Y(_2059_),
    .A(net46),
    .B(net685));
 sg13g2_xor2_1 _4665_ (.B(_2058_),
    .A(_0132_),
    .X(_2060_));
 sg13g2_o21ai_1 _4666_ (.B1(_2059_),
    .Y(_0449_),
    .A1(net651),
    .A2(_2060_));
 sg13g2_and3_2 _4667_ (.X(_2061_),
    .A(net46),
    .B(\pwm_module.counter2[14] ),
    .C(_2055_));
 sg13g2_nand2b_1 _4668_ (.Y(_2062_),
    .B(_2061_),
    .A_N(net686));
 sg13g2_nand2_1 _4669_ (.Y(_2063_),
    .A(\pwm_module.counter2[16] ),
    .B(_2061_));
 sg13g2_a21oi_1 _4670_ (.A1(_2012_),
    .A2(_2063_),
    .Y(_2064_),
    .B1(net685));
 sg13g2_a21oi_1 _4671_ (.A1(_2325_),
    .A2(_2062_),
    .Y(_0450_),
    .B1(_2064_));
 sg13g2_nand2_1 _4672_ (.Y(_2065_),
    .A(net89),
    .B(net685));
 sg13g2_xnor2_1 _4673_ (.Y(_2066_),
    .A(_0131_),
    .B(_2063_));
 sg13g2_o21ai_1 _4674_ (.B1(_2065_),
    .Y(_0451_),
    .A1(net652),
    .A2(_2066_));
 sg13g2_nor3_1 _4675_ (.A(_2323_),
    .B(net685),
    .C(_2063_),
    .Y(_2067_));
 sg13g2_and2_1 _4676_ (.A(\pwm_module.counter2[17] ),
    .B(\pwm_module.counter2[16] ),
    .X(_2068_));
 sg13g2_nor2_1 _4677_ (.A(net519),
    .B(_2067_),
    .Y(_2069_));
 sg13g2_nand4_1 _4678_ (.B(net89),
    .C(\pwm_module.counter2[16] ),
    .A(\pwm_module.counter2[18] ),
    .Y(_2070_),
    .D(_2061_));
 sg13g2_a21oi_1 _4679_ (.A1(_2012_),
    .A2(_2070_),
    .Y(_2071_),
    .B1(net685));
 sg13g2_nor2_1 _4680_ (.A(_2069_),
    .B(_2071_),
    .Y(_0452_));
 sg13g2_nand2_1 _4681_ (.Y(_2072_),
    .A(net64),
    .B(net685));
 sg13g2_xnor2_1 _4682_ (.Y(_2073_),
    .A(_0130_),
    .B(_2070_));
 sg13g2_o21ai_1 _4683_ (.B1(_2072_),
    .Y(_0453_),
    .A1(net650),
    .A2(_2073_));
 sg13g2_nand2_1 _4684_ (.Y(_2074_),
    .A(net303),
    .B(net680));
 sg13g2_nand4_1 _4685_ (.B(\pwm_module.counter2[18] ),
    .C(_2061_),
    .A(\pwm_module.counter2[19] ),
    .Y(_2075_),
    .D(_2068_));
 sg13g2_nor2_1 _4686_ (.A(_0129_),
    .B(_2075_),
    .Y(_2076_));
 sg13g2_xnor2_1 _4687_ (.Y(_2077_),
    .A(_0129_),
    .B(_2075_));
 sg13g2_o21ai_1 _4688_ (.B1(_2074_),
    .Y(_0454_),
    .A1(net650),
    .A2(_2077_));
 sg13g2_nand2_1 _4689_ (.Y(_2078_),
    .A(net209),
    .B(net680));
 sg13g2_xnor2_1 _4690_ (.Y(_2079_),
    .A(_2328_),
    .B(_2076_));
 sg13g2_o21ai_1 _4691_ (.B1(_2078_),
    .Y(_0455_),
    .A1(net650),
    .A2(_2079_));
 sg13g2_nand2_1 _4692_ (.Y(_2080_),
    .A(net209),
    .B(net303));
 sg13g2_nor2_1 _4693_ (.A(_2075_),
    .B(_2080_),
    .Y(_2081_));
 sg13g2_nand2b_1 _4694_ (.Y(_2082_),
    .B(_2081_),
    .A_N(net688));
 sg13g2_nand2_1 _4695_ (.Y(_2083_),
    .A(net481),
    .B(_2081_));
 sg13g2_a21oi_1 _4696_ (.A1(_2012_),
    .A2(_2083_),
    .Y(_2084_),
    .B1(net688));
 sg13g2_a21oi_1 _4697_ (.A1(_2327_),
    .A2(_2082_),
    .Y(_0456_),
    .B1(_2084_));
 sg13g2_nand2_1 _4698_ (.Y(_2085_),
    .A(net62),
    .B(net685));
 sg13g2_xnor2_1 _4699_ (.Y(_2086_),
    .A(_0127_),
    .B(_2083_));
 sg13g2_o21ai_1 _4700_ (.B1(_2085_),
    .Y(_0457_),
    .A1(net650),
    .A2(_2086_));
 sg13g2_nand4_1 _4701_ (.B(\pwm_module.counter2[22] ),
    .C(\pwm_module.counter2[21] ),
    .A(\pwm_module.counter2[23] ),
    .Y(_2087_),
    .D(\pwm_module.counter2[20] ));
 sg13g2_nor2_1 _4702_ (.A(_2075_),
    .B(_2087_),
    .Y(_2088_));
 sg13g2_nor2b_1 _4703_ (.A(net680),
    .B_N(_2088_),
    .Y(_2089_));
 sg13g2_xnor2_1 _4704_ (.Y(_2090_),
    .A(net546),
    .B(_2089_));
 sg13g2_nand2_1 _4705_ (.Y(_2091_),
    .A(\pwm_module.counter2[24] ),
    .B(_2088_));
 sg13g2_nor2_1 _4706_ (.A(_2015_),
    .B(_2090_),
    .Y(_0458_));
 sg13g2_nand2_1 _4707_ (.Y(_2092_),
    .A(net91),
    .B(net680));
 sg13g2_xnor2_1 _4708_ (.Y(_2093_),
    .A(_0126_),
    .B(_2091_));
 sg13g2_o21ai_1 _4709_ (.B1(_2092_),
    .Y(_0459_),
    .A1(net650),
    .A2(_2093_));
 sg13g2_nand3_1 _4710_ (.B(net580),
    .C(_2088_),
    .A(net91),
    .Y(_2094_));
 sg13g2_or2_1 _4711_ (.X(_2095_),
    .B(_2094_),
    .A(net681));
 sg13g2_or2_1 _4712_ (.X(_2096_),
    .B(_2094_),
    .A(_2330_));
 sg13g2_a21oi_1 _4713_ (.A1(_2012_),
    .A2(_2096_),
    .Y(_2097_),
    .B1(net680));
 sg13g2_a21oi_1 _4714_ (.A1(_2330_),
    .A2(_2095_),
    .Y(_0460_),
    .B1(_2097_));
 sg13g2_nand2_1 _4715_ (.Y(_2098_),
    .A(net66),
    .B(net681));
 sg13g2_xnor2_1 _4716_ (.Y(_2099_),
    .A(_0125_),
    .B(_2096_));
 sg13g2_o21ai_1 _4717_ (.B1(_2098_),
    .Y(_0461_),
    .A1(net650),
    .A2(_2099_));
 sg13g2_nand4_1 _4718_ (.B(\pwm_module.counter2[26] ),
    .C(\pwm_module.counter2[25] ),
    .A(net66),
    .Y(_2100_),
    .D(\pwm_module.counter2[24] ));
 sg13g2_nor3_1 _4719_ (.A(_2075_),
    .B(_2087_),
    .C(_2100_),
    .Y(_2101_));
 sg13g2_nor2b_1 _4720_ (.A(net680),
    .B_N(_2101_),
    .Y(_2102_));
 sg13g2_xnor2_1 _4721_ (.Y(_2103_),
    .A(net499),
    .B(_2102_));
 sg13g2_and2_1 _4722_ (.A(\pwm_module.counter2[28] ),
    .B(_2101_),
    .X(_2104_));
 sg13g2_nor2_1 _4723_ (.A(_2015_),
    .B(net500),
    .Y(_0462_));
 sg13g2_nand2_1 _4724_ (.Y(_2105_),
    .A(net85),
    .B(net681));
 sg13g2_xor2_1 _4725_ (.B(_2104_),
    .A(_0124_),
    .X(_2106_));
 sg13g2_o21ai_1 _4726_ (.B1(_2105_),
    .Y(_0463_),
    .A1(net650),
    .A2(_2106_));
 sg13g2_nand3b_1 _4727_ (.B(_2104_),
    .C(net85),
    .Y(_2107_),
    .A_N(net681));
 sg13g2_nand3_1 _4728_ (.B(net85),
    .C(_2104_),
    .A(net184),
    .Y(_2108_));
 sg13g2_a21oi_1 _4729_ (.A1(_2012_),
    .A2(_2108_),
    .Y(_2109_),
    .B1(net680));
 sg13g2_a21oi_1 _4730_ (.A1(_2332_),
    .A2(_2107_),
    .Y(_0464_),
    .B1(_2109_));
 sg13g2_nand2_1 _4731_ (.Y(_2110_),
    .A(net48),
    .B(net681));
 sg13g2_xnor2_1 _4732_ (.Y(_2111_),
    .A(_0168_),
    .B(_2108_));
 sg13g2_o21ai_1 _4733_ (.B1(_2110_),
    .Y(_0465_),
    .A1(net650),
    .A2(_2111_));
 sg13g2_nor2_2 _4734_ (.A(_0910_),
    .B(_1845_),
    .Y(_2112_));
 sg13g2_mux2_1 _4735_ (.A0(net173),
    .A1(net750),
    .S(net710),
    .X(_0466_));
 sg13g2_nor2_1 _4736_ (.A(net167),
    .B(net710),
    .Y(_2113_));
 sg13g2_a21oi_1 _4737_ (.A1(net724),
    .A2(net710),
    .Y(_0467_),
    .B1(_2113_));
 sg13g2_nor2_1 _4738_ (.A(net124),
    .B(net710),
    .Y(_2114_));
 sg13g2_a21oi_1 _4739_ (.A1(net720),
    .A2(net710),
    .Y(_0468_),
    .B1(_2114_));
 sg13g2_mux2_1 _4740_ (.A0(net206),
    .A1(net746),
    .S(net710),
    .X(_0469_));
 sg13g2_mux2_1 _4741_ (.A0(net168),
    .A1(net742),
    .S(net710),
    .X(_0470_));
 sg13g2_mux2_1 _4742_ (.A0(net113),
    .A1(net738),
    .S(_2112_),
    .X(_0471_));
 sg13g2_mux2_1 _4743_ (.A0(net140),
    .A1(net734),
    .S(_2112_),
    .X(_0472_));
 sg13g2_mux2_1 _4744_ (.A0(net336),
    .A1(net730),
    .S(net710),
    .X(_0473_));
 sg13g2_nor2_1 _4745_ (.A(_0103_),
    .B(_1587_),
    .Y(_2115_));
 sg13g2_nor2_1 _4746_ (.A(_0202_),
    .B(_1591_),
    .Y(_2116_));
 sg13g2_nand2_1 _4747_ (.Y(_2117_),
    .A(_0202_),
    .B(_1591_));
 sg13g2_xnor2_1 _4748_ (.Y(_2118_),
    .A(\pwm_module.counter1[30] ),
    .B(_1589_));
 sg13g2_nand3b_1 _4749_ (.B(_2117_),
    .C(_2118_),
    .Y(_2119_),
    .A_N(_2116_));
 sg13g2_nor2_1 _4750_ (.A(_2115_),
    .B(_2119_),
    .Y(_2120_));
 sg13g2_nand2_1 _4751_ (.Y(_2121_),
    .A(_0103_),
    .B(_1587_));
 sg13g2_o21ai_1 _4752_ (.B1(_2121_),
    .Y(_2122_),
    .A1(\pwm_module.counter1[28] ),
    .A2(_1601_));
 sg13g2_and2_1 _4753_ (.A(\pwm_module.counter1[28] ),
    .B(_1601_),
    .X(_2123_));
 sg13g2_nor4_2 _4754_ (.A(_2115_),
    .B(_2119_),
    .C(_2122_),
    .Y(_2124_),
    .D(_2123_));
 sg13g2_nor2_1 _4755_ (.A(_0104_),
    .B(_1595_),
    .Y(_2125_));
 sg13g2_a22oi_1 _4756_ (.Y(_2126_),
    .B1(_1599_),
    .B2(_2359_),
    .A2(_1594_),
    .A1(\pwm_module.counter1[26] ));
 sg13g2_nand2b_1 _4757_ (.Y(_2127_),
    .B(_2126_),
    .A_N(_2125_));
 sg13g2_nor2_1 _4758_ (.A(\pwm_module.counter1[24] ),
    .B(_1602_),
    .Y(_2128_));
 sg13g2_a21oi_1 _4759_ (.A1(_0105_),
    .A2(_1598_),
    .Y(_2129_),
    .B1(_2128_));
 sg13g2_a22oi_1 _4760_ (.Y(_2130_),
    .B1(_1595_),
    .B2(_0104_),
    .A2(_1593_),
    .A1(_2358_));
 sg13g2_a21oi_1 _4761_ (.A1(\pwm_module.counter1[24] ),
    .A2(_1602_),
    .Y(_2131_),
    .B1(_2127_));
 sg13g2_nand4_1 _4762_ (.B(_2129_),
    .C(_2130_),
    .A(_2124_),
    .Y(_2132_),
    .D(_2131_));
 sg13g2_inv_1 _4763_ (.Y(_2133_),
    .A(_2132_));
 sg13g2_nor2_1 _4764_ (.A(_0106_),
    .B(_1622_),
    .Y(_2134_));
 sg13g2_a221oi_1 _4765_ (.B2(\pwm_module.counter1[22] ),
    .C1(_2134_),
    .B1(_1625_),
    .A1(_2361_),
    .Y(_2135_),
    .A2(_1617_));
 sg13g2_a22oi_1 _4766_ (.Y(_2136_),
    .B1(_1624_),
    .B2(_2360_),
    .A2(_1622_),
    .A1(_0106_));
 sg13g2_a22oi_1 _4767_ (.Y(_2137_),
    .B1(_1631_),
    .B2(_0108_),
    .A2(_1616_),
    .A1(_0107_));
 sg13g2_nand2b_1 _4768_ (.Y(_2138_),
    .B(_1632_),
    .A_N(_0108_));
 sg13g2_nand4_1 _4769_ (.B(_2136_),
    .C(_2137_),
    .A(_2135_),
    .Y(_2139_),
    .D(_2138_));
 sg13g2_nor2_1 _4770_ (.A(\pwm_module.counter1[18] ),
    .B(_1641_),
    .Y(_2140_));
 sg13g2_a21oi_1 _4771_ (.A1(_0109_),
    .A2(_1637_),
    .Y(_2141_),
    .B1(_2140_));
 sg13g2_or2_1 _4772_ (.X(_2142_),
    .B(_1637_),
    .A(_0109_));
 sg13g2_nand2_1 _4773_ (.Y(_2143_),
    .A(\pwm_module.counter1[16] ),
    .B(_1619_));
 sg13g2_nor2_1 _4774_ (.A(\pwm_module.counter1[16] ),
    .B(_1619_),
    .Y(_2144_));
 sg13g2_a21oi_1 _4775_ (.A1(_0110_),
    .A2(_1627_),
    .Y(_2145_),
    .B1(_2144_));
 sg13g2_nand2_1 _4776_ (.Y(_2146_),
    .A(\pwm_module.counter1[18] ),
    .B(_1641_));
 sg13g2_o21ai_1 _4777_ (.B1(_2146_),
    .Y(_2147_),
    .A1(_0110_),
    .A2(_1627_));
 sg13g2_nand4_1 _4778_ (.B(_2142_),
    .C(_2143_),
    .A(_2141_),
    .Y(_2148_),
    .D(_2145_));
 sg13g2_or3_1 _4779_ (.A(_2139_),
    .B(_2147_),
    .C(_2148_),
    .X(_2149_));
 sg13g2_nor2_1 _4780_ (.A(_2132_),
    .B(_2149_),
    .Y(_2150_));
 sg13g2_a22oi_1 _4781_ (.Y(_2151_),
    .B1(_1658_),
    .B2(_0113_),
    .A2(_1655_),
    .A1(_0112_));
 sg13g2_nand3b_1 _4782_ (.B(\MemCell.counter_value[15] ),
    .C(_0111_),
    .Y(_2152_),
    .A_N(net795));
 sg13g2_o21ai_1 _4783_ (.B1(_2152_),
    .Y(_2153_),
    .A1(\pwm_module.counter1[14] ),
    .A2(_1651_));
 sg13g2_or2_1 _4784_ (.X(_2154_),
    .B(_1648_),
    .A(_0111_));
 sg13g2_a22oi_1 _4785_ (.Y(_2155_),
    .B1(_1656_),
    .B2(_2363_),
    .A2(_1651_),
    .A1(\pwm_module.counter1[14] ));
 sg13g2_nand3b_1 _4786_ (.B(_2154_),
    .C(_2155_),
    .Y(_2156_),
    .A_N(_2153_));
 sg13g2_nor2_1 _4787_ (.A(_2151_),
    .B(_2156_),
    .Y(_2157_));
 sg13g2_o21ai_1 _4788_ (.B1(_2151_),
    .Y(_2158_),
    .A1(_0113_),
    .A2(_1658_));
 sg13g2_nor2_1 _4789_ (.A(_2156_),
    .B(_2158_),
    .Y(_2159_));
 sg13g2_and2_1 _4790_ (.A(_0114_),
    .B(_1662_),
    .X(_2160_));
 sg13g2_nand2_1 _4791_ (.Y(_2161_),
    .A(_0114_),
    .B(_1662_));
 sg13g2_nor2_1 _4792_ (.A(_0114_),
    .B(_1662_),
    .Y(_2162_));
 sg13g2_or2_1 _4793_ (.X(_2163_),
    .B(_1660_),
    .A(\pwm_module.counter1[10] ));
 sg13g2_a21oi_1 _4794_ (.A1(_2161_),
    .A2(_2163_),
    .Y(_2164_),
    .B1(_2162_));
 sg13g2_nand2_1 _4795_ (.Y(_2165_),
    .A(_0116_),
    .B(_1666_));
 sg13g2_o21ai_1 _4796_ (.B1(_2165_),
    .Y(_2166_),
    .A1(\pwm_module.counter1[8] ),
    .A2(_1668_));
 sg13g2_nor2_1 _4797_ (.A(_0116_),
    .B(_1666_),
    .Y(_2167_));
 sg13g2_xor2_1 _4798_ (.B(_1660_),
    .A(_0115_),
    .X(_2168_));
 sg13g2_nor4_1 _4799_ (.A(_2160_),
    .B(_2162_),
    .C(_2167_),
    .D(_2168_),
    .Y(_2169_));
 sg13g2_a21o_1 _4800_ (.A2(_2169_),
    .A1(_2166_),
    .B1(_2164_),
    .X(_2170_));
 sg13g2_a221oi_1 _4801_ (.B2(_2170_),
    .C1(_2157_),
    .B1(_2159_),
    .A1(_2153_),
    .Y(_2171_),
    .A2(_2154_));
 sg13g2_nor2_1 _4802_ (.A(\pwm_module.counter1[2] ),
    .B(_1693_),
    .Y(_2172_));
 sg13g2_a21oi_1 _4803_ (.A1(_0121_),
    .A2(_1691_),
    .Y(_2173_),
    .B1(_2172_));
 sg13g2_and2_1 _4804_ (.A(\pwm_module.counter1[2] ),
    .B(_1693_),
    .X(_2174_));
 sg13g2_nor2_1 _4805_ (.A(\pwm_module.counter1[1] ),
    .B(_1695_),
    .Y(_2175_));
 sg13g2_nand2_1 _4806_ (.Y(_2176_),
    .A(net728),
    .B(_1698_));
 sg13g2_xnor2_1 _4807_ (.Y(_2177_),
    .A(_2368_),
    .B(_1695_));
 sg13g2_a21oi_1 _4808_ (.A1(_2176_),
    .A2(_2177_),
    .Y(_2178_),
    .B1(_2175_));
 sg13g2_o21ai_1 _4809_ (.B1(_2173_),
    .Y(_2179_),
    .A1(_2174_),
    .A2(_2178_));
 sg13g2_nand2b_1 _4810_ (.Y(_2180_),
    .B(_1682_),
    .A_N(_0118_));
 sg13g2_nand2_1 _4811_ (.Y(_2181_),
    .A(\pwm_module.counter1[7] ),
    .B(_1680_));
 sg13g2_or2_1 _4812_ (.X(_2182_),
    .B(_1680_),
    .A(\pwm_module.counter1[7] ));
 sg13g2_a22oi_1 _4813_ (.Y(_2183_),
    .B1(_1686_),
    .B2(\pwm_module.counter1[5] ),
    .A2(_1683_),
    .A1(_0118_));
 sg13g2_nand4_1 _4814_ (.B(_2181_),
    .C(_2182_),
    .A(_2180_),
    .Y(_2184_),
    .D(_2183_));
 sg13g2_nand2_1 _4815_ (.Y(_2185_),
    .A(_2367_),
    .B(_1690_));
 sg13g2_o21ai_1 _4816_ (.B1(_2185_),
    .Y(_2186_),
    .A1(\pwm_module.counter1[5] ),
    .A2(_1686_));
 sg13g2_nor2_1 _4817_ (.A(_2367_),
    .B(_1690_),
    .Y(_2187_));
 sg13g2_nor2_1 _4818_ (.A(_0121_),
    .B(_1691_),
    .Y(_2188_));
 sg13g2_nor4_1 _4819_ (.A(_2184_),
    .B(_2186_),
    .C(_2187_),
    .D(_2188_),
    .Y(_2189_));
 sg13g2_nor2b_1 _4820_ (.A(_2184_),
    .B_N(_2186_),
    .Y(_2190_));
 sg13g2_o21ai_1 _4821_ (.B1(_2182_),
    .Y(_2191_),
    .A1(\pwm_module.counter1[6] ),
    .A2(_1682_));
 sg13g2_a221oi_1 _4822_ (.B2(_2181_),
    .C1(_2190_),
    .B1(_2191_),
    .A1(_2179_),
    .Y(_2192_),
    .A2(_2189_));
 sg13g2_a21oi_1 _4823_ (.A1(\pwm_module.counter1[8] ),
    .A2(_1668_),
    .Y(_2193_),
    .B1(_2166_));
 sg13g2_nand3_1 _4824_ (.B(_2169_),
    .C(_2193_),
    .A(_2159_),
    .Y(_2194_));
 sg13g2_o21ai_1 _4825_ (.B1(_2171_),
    .Y(_2195_),
    .A1(_2192_),
    .A2(_2194_));
 sg13g2_o21ai_1 _4826_ (.B1(_2141_),
    .Y(_2196_),
    .A1(_2145_),
    .A2(_2147_));
 sg13g2_nand3b_1 _4827_ (.B(_2142_),
    .C(_2196_),
    .Y(_2197_),
    .A_N(_2139_));
 sg13g2_nand2b_1 _4828_ (.Y(_2198_),
    .B(_2135_),
    .A_N(_2137_));
 sg13g2_o21ai_1 _4829_ (.B1(_2198_),
    .Y(_2199_),
    .A1(_2134_),
    .A2(_2136_));
 sg13g2_nand2b_1 _4830_ (.Y(_2200_),
    .B(_2197_),
    .A_N(_2199_));
 sg13g2_nor3_1 _4831_ (.A(\pwm_module.counter1[30] ),
    .B(_1590_),
    .C(_2116_),
    .Y(_2201_));
 sg13g2_a221oi_1 _4832_ (.B2(_2122_),
    .C1(_2201_),
    .B1(_2120_),
    .A1(_0202_),
    .Y(_2202_),
    .A2(_1591_));
 sg13g2_nor2_1 _4833_ (.A(_2125_),
    .B(_2130_),
    .Y(_2203_));
 sg13g2_nor2_1 _4834_ (.A(_2127_),
    .B(_2129_),
    .Y(_2204_));
 sg13g2_o21ai_1 _4835_ (.B1(_2124_),
    .Y(_2205_),
    .A1(_2203_),
    .A2(_2204_));
 sg13g2_nand2_2 _4836_ (.Y(_2206_),
    .A(_2202_),
    .B(_2205_));
 sg13g2_a221oi_1 _4837_ (.B2(_2133_),
    .C1(_2206_),
    .B1(_2200_),
    .A1(_2150_),
    .Y(_2207_),
    .A2(_2195_));
 sg13g2_nor2_1 _4838_ (.A(net728),
    .B(_1698_),
    .Y(_2208_));
 sg13g2_nor3_1 _4839_ (.A(_2174_),
    .B(_2188_),
    .C(_2208_),
    .Y(_2209_));
 sg13g2_nand4_1 _4840_ (.B(_2176_),
    .C(_2177_),
    .A(_2173_),
    .Y(_2210_),
    .D(_2209_));
 sg13g2_or4_1 _4841_ (.A(_2184_),
    .B(_2186_),
    .C(_2187_),
    .D(_2210_),
    .X(_2211_));
 sg13g2_nor4_1 _4842_ (.A(_2132_),
    .B(_2149_),
    .C(_2194_),
    .D(_2211_),
    .Y(_2212_));
 sg13g2_nor3_1 _4843_ (.A(_2395_),
    .B(_2207_),
    .C(_2212_),
    .Y(_2213_));
 sg13g2_nand2_2 _4844_ (.Y(_2214_),
    .A(net677),
    .B(net657));
 sg13g2_a21oi_1 _4845_ (.A1(net676),
    .A2(net657),
    .Y(_2215_),
    .B1(net728));
 sg13g2_a21oi_1 _4846_ (.A1(net728),
    .A2(net676),
    .Y(_0474_),
    .B1(_2215_));
 sg13g2_nand2_1 _4847_ (.Y(_2216_),
    .A(net551),
    .B(net728));
 sg13g2_or2_1 _4848_ (.X(_2217_),
    .B(net728),
    .A(net551));
 sg13g2_nand4_1 _4849_ (.B(net656),
    .C(_2216_),
    .A(net676),
    .Y(_2218_),
    .D(_2217_));
 sg13g2_o21ai_1 _4850_ (.B1(_2218_),
    .Y(_0475_),
    .A1(_2368_),
    .A2(net676));
 sg13g2_nand3_1 _4851_ (.B(net697),
    .C(net694),
    .A(net533),
    .Y(_2219_));
 sg13g2_nand3_1 _4852_ (.B(\pwm_module.counter1[1] ),
    .C(net728),
    .A(\pwm_module.counter1[2] ),
    .Y(_2220_));
 sg13g2_xor2_1 _4853_ (.B(_2216_),
    .A(net533),
    .X(_2221_));
 sg13g2_o21ai_1 _4854_ (.B1(_2219_),
    .Y(_0476_),
    .A1(net648),
    .A2(_2221_));
 sg13g2_xor2_1 _4855_ (.B(_2220_),
    .A(_0121_),
    .X(_2222_));
 sg13g2_nand3_1 _4856_ (.B(net656),
    .C(_2222_),
    .A(net676),
    .Y(_2223_));
 sg13g2_o21ai_1 _4857_ (.B1(_2223_),
    .Y(_0477_),
    .A1(_2390_),
    .A2(net676));
 sg13g2_nand4_1 _4858_ (.B(\pwm_module.counter1[1] ),
    .C(net728),
    .A(\pwm_module.counter1[2] ),
    .Y(_2224_),
    .D(net152));
 sg13g2_nor2_1 _4859_ (.A(_2367_),
    .B(_2224_),
    .Y(_2225_));
 sg13g2_xnor2_1 _4860_ (.Y(_2226_),
    .A(net441),
    .B(_2224_));
 sg13g2_nand3_1 _4861_ (.B(net656),
    .C(_2226_),
    .A(net676),
    .Y(_2227_));
 sg13g2_o21ai_1 _4862_ (.B1(_2227_),
    .Y(_0478_),
    .A1(_2367_),
    .A2(net677));
 sg13g2_xnor2_1 _4863_ (.Y(_2228_),
    .A(_0119_),
    .B(_2225_));
 sg13g2_nand3_1 _4864_ (.B(net656),
    .C(_2228_),
    .A(net676),
    .Y(_2229_));
 sg13g2_o21ai_1 _4865_ (.B1(_2229_),
    .Y(_0479_),
    .A1(_2366_),
    .A2(net677));
 sg13g2_nand3_1 _4866_ (.B(net697),
    .C(net694),
    .A(net254),
    .Y(_2230_));
 sg13g2_nor3_2 _4867_ (.A(_2366_),
    .B(_2367_),
    .C(_2224_),
    .Y(_2231_));
 sg13g2_nor2b_1 _4868_ (.A(_0118_),
    .B_N(_2231_),
    .Y(_2232_));
 sg13g2_xor2_1 _4869_ (.B(_2231_),
    .A(_0118_),
    .X(_2233_));
 sg13g2_o21ai_1 _4870_ (.B1(_2230_),
    .Y(_0480_),
    .A1(_2214_),
    .A2(_2233_));
 sg13g2_nand3_1 _4871_ (.B(net697),
    .C(net694),
    .A(net233),
    .Y(_2234_));
 sg13g2_xor2_1 _4872_ (.B(_2232_),
    .A(_0117_),
    .X(_2235_));
 sg13g2_o21ai_1 _4873_ (.B1(_2234_),
    .Y(_0481_),
    .A1(_2214_),
    .A2(_2235_));
 sg13g2_and2_1 _4874_ (.A(\pwm_module.counter1[6] ),
    .B(\pwm_module.counter1[7] ),
    .X(_2236_));
 sg13g2_and2_1 _4875_ (.A(_2231_),
    .B(_2236_),
    .X(_2237_));
 sg13g2_or2_1 _4876_ (.X(_2238_),
    .B(_2237_),
    .A(net549));
 sg13g2_nand2_1 _4877_ (.Y(_2239_),
    .A(\pwm_module.counter1[8] ),
    .B(_2237_));
 sg13g2_nand4_1 _4878_ (.B(net656),
    .C(_2238_),
    .A(net677),
    .Y(_2240_),
    .D(_2239_));
 sg13g2_o21ai_1 _4879_ (.B1(_2240_),
    .Y(_0482_),
    .A1(_2364_),
    .A2(net677));
 sg13g2_nand3_1 _4880_ (.B(net695),
    .C(net692),
    .A(net109),
    .Y(_2241_));
 sg13g2_xnor2_1 _4881_ (.Y(_2242_),
    .A(_0116_),
    .B(_2239_));
 sg13g2_o21ai_1 _4882_ (.B1(_2241_),
    .Y(_0483_),
    .A1(_2214_),
    .A2(_2242_));
 sg13g2_nand3_1 _4883_ (.B(net695),
    .C(net692),
    .A(net359),
    .Y(_2243_));
 sg13g2_nand4_1 _4884_ (.B(\pwm_module.counter1[8] ),
    .C(_2231_),
    .A(\pwm_module.counter1[9] ),
    .Y(_2244_),
    .D(_2236_));
 sg13g2_nor2_1 _4885_ (.A(_0115_),
    .B(_2244_),
    .Y(_2245_));
 sg13g2_xnor2_1 _4886_ (.Y(_2246_),
    .A(_0115_),
    .B(_2244_));
 sg13g2_o21ai_1 _4887_ (.B1(_2243_),
    .Y(_0484_),
    .A1(net648),
    .A2(_2246_));
 sg13g2_nand3_1 _4888_ (.B(net695),
    .C(net692),
    .A(net87),
    .Y(_2247_));
 sg13g2_xor2_1 _4889_ (.B(_2245_),
    .A(_0114_),
    .X(_2248_));
 sg13g2_o21ai_1 _4890_ (.B1(_2247_),
    .Y(_0485_),
    .A1(net648),
    .A2(_2248_));
 sg13g2_nand3_1 _4891_ (.B(net695),
    .C(net692),
    .A(net194),
    .Y(_2249_));
 sg13g2_nand2_1 _4892_ (.Y(_2250_),
    .A(net359),
    .B(net87));
 sg13g2_nor2_1 _4893_ (.A(_2244_),
    .B(_2250_),
    .Y(_2251_));
 sg13g2_nor3_1 _4894_ (.A(_0113_),
    .B(_2244_),
    .C(_2250_),
    .Y(_2252_));
 sg13g2_xor2_1 _4895_ (.B(_2251_),
    .A(_0113_),
    .X(_2253_));
 sg13g2_o21ai_1 _4896_ (.B1(_2249_),
    .Y(_0486_),
    .A1(net648),
    .A2(_2253_));
 sg13g2_nand3_1 _4897_ (.B(net695),
    .C(net692),
    .A(net120),
    .Y(_2254_));
 sg13g2_xnor2_1 _4898_ (.Y(_2255_),
    .A(_2363_),
    .B(_2252_));
 sg13g2_o21ai_1 _4899_ (.B1(_2254_),
    .Y(_0487_),
    .A1(net648),
    .A2(_2255_));
 sg13g2_nand2_1 _4900_ (.Y(_2256_),
    .A(net120),
    .B(net194));
 sg13g2_nor3_2 _4901_ (.A(_2244_),
    .B(_2250_),
    .C(_2256_),
    .Y(_2257_));
 sg13g2_a21oi_1 _4902_ (.A1(net674),
    .A2(_2257_),
    .Y(_2258_),
    .B1(net414));
 sg13g2_nand2_1 _4903_ (.Y(_2259_),
    .A(\pwm_module.counter1[14] ),
    .B(_2257_));
 sg13g2_nand2_1 _4904_ (.Y(_2260_),
    .A(net656),
    .B(_2259_));
 sg13g2_a21oi_1 _4905_ (.A1(net674),
    .A2(_2260_),
    .Y(_0488_),
    .B1(_2258_));
 sg13g2_nand3_1 _4906_ (.B(net695),
    .C(net692),
    .A(net106),
    .Y(_2261_));
 sg13g2_xnor2_1 _4907_ (.Y(_2262_),
    .A(_0111_),
    .B(_2259_));
 sg13g2_o21ai_1 _4908_ (.B1(_2261_),
    .Y(_0489_),
    .A1(net648),
    .A2(_2262_));
 sg13g2_and3_1 _4909_ (.X(_2263_),
    .A(\pwm_module.counter1[14] ),
    .B(net106),
    .C(_2257_));
 sg13g2_nand3_1 _4910_ (.B(\pwm_module.counter1[15] ),
    .C(_2257_),
    .A(\pwm_module.counter1[14] ),
    .Y(_2264_));
 sg13g2_nand2_1 _4911_ (.Y(_2265_),
    .A(\pwm_module.counter1[16] ),
    .B(_2263_));
 sg13g2_nand2_1 _4912_ (.Y(_2266_),
    .A(net656),
    .B(_2265_));
 sg13g2_a21oi_1 _4913_ (.A1(net674),
    .A2(_2263_),
    .Y(_2267_),
    .B1(net467));
 sg13g2_a21oi_1 _4914_ (.A1(net674),
    .A2(_2266_),
    .Y(_0490_),
    .B1(net468));
 sg13g2_nand3_1 _4915_ (.B(net695),
    .C(net692),
    .A(net95),
    .Y(_2268_));
 sg13g2_xnor2_1 _4916_ (.Y(_2269_),
    .A(_0110_),
    .B(_2265_));
 sg13g2_o21ai_1 _4917_ (.B1(_2268_),
    .Y(_0491_),
    .A1(net648),
    .A2(_2269_));
 sg13g2_and3_1 _4918_ (.X(_2270_),
    .A(\pwm_module.counter1[16] ),
    .B(net95),
    .C(_2263_));
 sg13g2_a21oi_1 _4919_ (.A1(net674),
    .A2(_2270_),
    .Y(_2271_),
    .B1(net491));
 sg13g2_nand2_1 _4920_ (.Y(_2272_),
    .A(\pwm_module.counter1[18] ),
    .B(_2270_));
 sg13g2_nand2_1 _4921_ (.Y(_2273_),
    .A(net656),
    .B(_2272_));
 sg13g2_a21oi_1 _4922_ (.A1(net674),
    .A2(_2273_),
    .Y(_0492_),
    .B1(_2271_));
 sg13g2_nand3_1 _4923_ (.B(net695),
    .C(net692),
    .A(net68),
    .Y(_2274_));
 sg13g2_xnor2_1 _4924_ (.Y(_2275_),
    .A(_0109_),
    .B(_2272_));
 sg13g2_o21ai_1 _4925_ (.B1(_2274_),
    .Y(_0493_),
    .A1(net648),
    .A2(_2275_));
 sg13g2_nand3_1 _4926_ (.B(net696),
    .C(net693),
    .A(net229),
    .Y(_2276_));
 sg13g2_nand4_1 _4927_ (.B(\pwm_module.counter1[16] ),
    .C(net68),
    .A(\pwm_module.counter1[18] ),
    .Y(_2277_),
    .D(net95));
 sg13g2_nor2_1 _4928_ (.A(_2264_),
    .B(_2277_),
    .Y(_2278_));
 sg13g2_or2_1 _4929_ (.X(_2279_),
    .B(_2277_),
    .A(_2264_));
 sg13g2_xnor2_1 _4930_ (.Y(_2280_),
    .A(net334),
    .B(_2279_));
 sg13g2_o21ai_1 _4931_ (.B1(_2276_),
    .Y(_0494_),
    .A1(net649),
    .A2(_2280_));
 sg13g2_nand3_1 _4932_ (.B(net696),
    .C(net693),
    .A(net212),
    .Y(_2281_));
 sg13g2_nor2_1 _4933_ (.A(_0108_),
    .B(_2279_),
    .Y(_2282_));
 sg13g2_xnor2_1 _4934_ (.Y(_2283_),
    .A(_2361_),
    .B(_2282_));
 sg13g2_o21ai_1 _4935_ (.B1(_2281_),
    .Y(_0495_),
    .A1(net649),
    .A2(_2283_));
 sg13g2_nand4_1 _4936_ (.B(net229),
    .C(net674),
    .A(net212),
    .Y(_2284_),
    .D(_2278_));
 sg13g2_nand3_1 _4937_ (.B(net212),
    .C(\pwm_module.counter1[20] ),
    .A(\pwm_module.counter1[22] ),
    .Y(_2285_));
 sg13g2_nor2_1 _4938_ (.A(_2279_),
    .B(_2285_),
    .Y(_2286_));
 sg13g2_nand2b_1 _4939_ (.Y(_2287_),
    .B(net657),
    .A_N(_2286_));
 sg13g2_a22oi_1 _4940_ (.Y(_0496_),
    .B1(_2287_),
    .B2(net674),
    .A2(net230),
    .A1(_2360_));
 sg13g2_nand3_1 _4941_ (.B(net696),
    .C(net693),
    .A(net58),
    .Y(_2288_));
 sg13g2_xor2_1 _4942_ (.B(_2286_),
    .A(_0106_),
    .X(_2289_));
 sg13g2_o21ai_1 _4943_ (.B1(_2288_),
    .Y(_0497_),
    .A1(net649),
    .A2(_2289_));
 sg13g2_nor4_2 _4944_ (.A(_2391_),
    .B(_2264_),
    .C(_2277_),
    .Y(_2290_),
    .D(_2285_));
 sg13g2_a21oi_1 _4945_ (.A1(net671),
    .A2(_2290_),
    .Y(_2291_),
    .B1(net445));
 sg13g2_and2_1 _4946_ (.A(\pwm_module.counter1[24] ),
    .B(_2290_),
    .X(_2292_));
 sg13g2_nand2b_1 _4947_ (.Y(_2293_),
    .B(net657),
    .A_N(_2292_));
 sg13g2_a21oi_1 _4948_ (.A1(net671),
    .A2(_2293_),
    .Y(_0498_),
    .B1(net446));
 sg13g2_nand3_1 _4949_ (.B(net696),
    .C(net693),
    .A(net162),
    .Y(_2294_));
 sg13g2_xnor2_1 _4950_ (.Y(_2295_),
    .A(_2359_),
    .B(_2292_));
 sg13g2_o21ai_1 _4951_ (.B1(_2294_),
    .Y(_0499_),
    .A1(net649),
    .A2(_2295_));
 sg13g2_nand3_1 _4952_ (.B(net671),
    .C(_2292_),
    .A(net162),
    .Y(_2296_));
 sg13g2_nand3_1 _4953_ (.B(net162),
    .C(_2292_),
    .A(net390),
    .Y(_2297_));
 sg13g2_nand2_1 _4954_ (.Y(_2298_),
    .A(net657),
    .B(_2297_));
 sg13g2_a22oi_1 _4955_ (.Y(_0500_),
    .B1(_2298_),
    .B2(net671),
    .A2(_2296_),
    .A1(_2358_));
 sg13g2_nand3_1 _4956_ (.B(net696),
    .C(net693),
    .A(net83),
    .Y(_2299_));
 sg13g2_xnor2_1 _4957_ (.Y(_2300_),
    .A(_0104_),
    .B(_2297_));
 sg13g2_o21ai_1 _4958_ (.B1(_2299_),
    .Y(_0501_),
    .A1(net649),
    .A2(_2300_));
 sg13g2_and4_1 _4959_ (.A(\pwm_module.counter1[26] ),
    .B(\pwm_module.counter1[24] ),
    .C(\pwm_module.counter1[27] ),
    .D(\pwm_module.counter1[25] ),
    .X(_2301_));
 sg13g2_and2_1 _4960_ (.A(_2290_),
    .B(_2301_),
    .X(_2302_));
 sg13g2_a21oi_1 _4961_ (.A1(net671),
    .A2(_2302_),
    .Y(_2303_),
    .B1(net506));
 sg13g2_nand2_1 _4962_ (.Y(_2304_),
    .A(\pwm_module.counter1[28] ),
    .B(_2302_));
 sg13g2_nand2_1 _4963_ (.Y(_2305_),
    .A(net657),
    .B(_2304_));
 sg13g2_a21oi_1 _4964_ (.A1(net671),
    .A2(_2305_),
    .Y(_0502_),
    .B1(_2303_));
 sg13g2_nand3_1 _4965_ (.B(net696),
    .C(net693),
    .A(net159),
    .Y(_2306_));
 sg13g2_xnor2_1 _4966_ (.Y(_2307_),
    .A(_0103_),
    .B(_2304_));
 sg13g2_o21ai_1 _4967_ (.B1(_2306_),
    .Y(_0503_),
    .A1(net649),
    .A2(_2307_));
 sg13g2_nand4_1 _4968_ (.B(net159),
    .C(net671),
    .A(\pwm_module.counter1[28] ),
    .Y(_2308_),
    .D(_2302_));
 sg13g2_nand4_1 _4969_ (.B(\pwm_module.counter1[28] ),
    .C(net159),
    .A(\pwm_module.counter1[30] ),
    .Y(_2309_),
    .D(_2302_));
 sg13g2_nand2_1 _4970_ (.Y(_2310_),
    .A(net657),
    .B(_2309_));
 sg13g2_a22oi_1 _4971_ (.Y(_0504_),
    .B1(_2310_),
    .B2(net671),
    .A2(_2308_),
    .A1(_2357_));
 sg13g2_nand3_1 _4972_ (.B(net696),
    .C(net693),
    .A(net38),
    .Y(_2311_));
 sg13g2_xnor2_1 _4973_ (.Y(_2312_),
    .A(_0202_),
    .B(_2309_));
 sg13g2_o21ai_1 _4974_ (.B1(_2311_),
    .Y(_0505_),
    .A1(net649),
    .A2(_2312_));
 sg13g2_inv_1 _4975_ (.Y(_0220_),
    .A(net763));
 sg13g2_inv_1 _4976_ (.Y(_0221_),
    .A(net763));
 sg13g2_inv_1 _4977_ (.Y(_0222_),
    .A(net763));
 sg13g2_dfrbp_1 _4978_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net859),
    .D(net1),
    .Q_N(_2620_),
    .Q(reg_ui0));
 sg13g2_dfrbp_1 _4979_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net859),
    .D(net2),
    .Q_N(_0166_),
    .Q(reg_ui1));
 sg13g2_dfrbp_1 _4980_ (.CLK(net766),
    .RESET_B(_0219_),
    .D(_2398_),
    .Q_N(_2398_),
    .Q(\spi_module.r_RX_Bit_Count[0] ));
 sg13g2_dfrbp_1 _4981_ (.CLK(net766),
    .RESET_B(_0220_),
    .D(_0100_),
    .Q_N(_2619_),
    .Q(\spi_module.r_RX_Bit_Count[1] ));
 sg13g2_dfrbp_1 _4982_ (.CLK(net766),
    .RESET_B(_0221_),
    .D(_0101_),
    .Q_N(_2618_),
    .Q(\spi_module.r_RX_Bit_Count[2] ));
 sg13g2_dfrbp_1 _4983_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net797),
    .D(_0223_),
    .Q_N(_0165_),
    .Q(\pwm_module.counter0[0] ));
 sg13g2_dfrbp_1 _4984_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net797),
    .D(_0224_),
    .Q_N(_0164_),
    .Q(\pwm_module.counter0[1] ));
 sg13g2_dfrbp_1 _4985_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net797),
    .D(_0225_),
    .Q_N(_2617_),
    .Q(\pwm_module.counter0[2] ));
 sg13g2_dfrbp_1 _4986_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net797),
    .D(net61),
    .Q_N(_0163_),
    .Q(\pwm_module.counter0[3] ));
 sg13g2_dfrbp_1 _4987_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net797),
    .D(_0227_),
    .Q_N(_0162_),
    .Q(\pwm_module.counter0[4] ));
 sg13g2_dfrbp_1 _4988_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net800),
    .D(net253),
    .Q_N(_0161_),
    .Q(\pwm_module.counter0[5] ));
 sg13g2_dfrbp_1 _4989_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net799),
    .D(net291),
    .Q_N(_0160_),
    .Q(\pwm_module.counter0[6] ));
 sg13g2_dfrbp_1 _4990_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net799),
    .D(net266),
    .Q_N(_0159_),
    .Q(\pwm_module.counter0[7] ));
 sg13g2_dfrbp_1 _4991_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net799),
    .D(_0231_),
    .Q_N(_2616_),
    .Q(\pwm_module.counter0[8] ));
 sg13g2_dfrbp_1 _4992_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net798),
    .D(net368),
    .Q_N(_0158_),
    .Q(\pwm_module.counter0[9] ));
 sg13g2_dfrbp_1 _4993_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net798),
    .D(net456),
    .Q_N(_0157_),
    .Q(\pwm_module.counter0[10] ));
 sg13g2_dfrbp_1 _4994_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net798),
    .D(net98),
    .Q_N(_0156_),
    .Q(\pwm_module.counter0[11] ));
 sg13g2_dfrbp_1 _4995_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net799),
    .D(net199),
    .Q_N(_0155_),
    .Q(\pwm_module.counter0[12] ));
 sg13g2_dfrbp_1 _4996_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net798),
    .D(net435),
    .Q_N(_0154_),
    .Q(\pwm_module.counter0[13] ));
 sg13g2_dfrbp_1 _4997_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net799),
    .D(net555),
    .Q_N(_2615_),
    .Q(\pwm_module.counter0[14] ));
 sg13g2_dfrbp_1 _4998_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net799),
    .D(net71),
    .Q_N(_0153_),
    .Q(\pwm_module.counter0[15] ));
 sg13g2_dfrbp_1 _4999_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net802),
    .D(_0239_),
    .Q_N(_2614_),
    .Q(\pwm_module.counter0[16] ));
 sg13g2_dfrbp_1 _5000_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net802),
    .D(net248),
    .Q_N(_0152_),
    .Q(\pwm_module.counter0[17] ));
 sg13g2_dfrbp_1 _5001_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net800),
    .D(_0241_),
    .Q_N(_2613_),
    .Q(\pwm_module.counter0[18] ));
 sg13g2_dfrbp_1 _5002_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net802),
    .D(net53),
    .Q_N(_0151_),
    .Q(\pwm_module.counter0[19] ));
 sg13g2_dfrbp_1 _5003_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net801),
    .D(net237),
    .Q_N(_0150_),
    .Q(\pwm_module.counter0[20] ));
 sg13g2_dfrbp_1 _5004_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net801),
    .D(net426),
    .Q_N(_0149_),
    .Q(\pwm_module.counter0[21] ));
 sg13g2_dfrbp_1 _5005_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net802),
    .D(net536),
    .Q_N(_2612_),
    .Q(\pwm_module.counter0[22] ));
 sg13g2_dfrbp_1 _5006_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net801),
    .D(net51),
    .Q_N(_0148_),
    .Q(\pwm_module.counter0[23] ));
 sg13g2_dfrbp_1 _5007_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net813),
    .D(_0247_),
    .Q_N(_2611_),
    .Q(\pwm_module.counter0[24] ));
 sg13g2_dfrbp_1 _5008_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net813),
    .D(net401),
    .Q_N(_0147_),
    .Q(\pwm_module.counter0[25] ));
 sg13g2_dfrbp_1 _5009_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net813),
    .D(net553),
    .Q_N(_2610_),
    .Q(\pwm_module.counter0[26] ));
 sg13g2_dfrbp_1 _5010_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net812),
    .D(net73),
    .Q_N(_0146_),
    .Q(\pwm_module.counter0[27] ));
 sg13g2_dfrbp_1 _5011_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net814),
    .D(_0251_),
    .Q_N(_2609_),
    .Q(\pwm_module.counter0[28] ));
 sg13g2_dfrbp_1 _5012_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net813),
    .D(net327),
    .Q_N(_0145_),
    .Q(\pwm_module.counter0[29] ));
 sg13g2_dfrbp_1 _5013_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net813),
    .D(net484),
    .Q_N(_2608_),
    .Q(\pwm_module.counter0[30] ));
 sg13g2_dfrbp_1 _5014_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net812),
    .D(net45),
    .Q_N(_0167_),
    .Q(\pwm_module.counter0[31] ));
 sg13g2_dfrbp_1 _5015_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net837),
    .D(net35),
    .Q_N(_2621_),
    .Q(\spi_module.r3_RX_Done ));
 sg13g2_dfrbp_1 _5016_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net840),
    .D(net718),
    .Q_N(_2607_),
    .Q(\MemCell.o_RX_DV ));
 sg13g2_dfrbp_1 _5017_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net840),
    .D(_0255_),
    .Q_N(_2606_),
    .Q(\MemCell.o_RX_Byte[0] ));
 sg13g2_dfrbp_1 _5018_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net840),
    .D(_0256_),
    .Q_N(_2605_),
    .Q(\MemCell.o_RX_Byte[1] ));
 sg13g2_dfrbp_1 _5019_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net840),
    .D(_0257_),
    .Q_N(_2604_),
    .Q(\MemCell.o_RX_Byte[2] ));
 sg13g2_dfrbp_1 _5020_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net843),
    .D(_0258_),
    .Q_N(_2603_),
    .Q(\MemCell.o_RX_Byte[3] ));
 sg13g2_dfrbp_1 _5021_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net843),
    .D(_0259_),
    .Q_N(_2602_),
    .Q(\MemCell.o_RX_Byte[4] ));
 sg13g2_dfrbp_1 _5022_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net843),
    .D(_0260_),
    .Q_N(_2601_),
    .Q(\MemCell.o_RX_Byte[5] ));
 sg13g2_dfrbp_1 _5023_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net837),
    .D(_0261_),
    .Q_N(_2600_),
    .Q(\MemCell.o_RX_Byte[6] ));
 sg13g2_dfrbp_1 _5024_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net837),
    .D(_0262_),
    .Q_N(_2599_),
    .Q(\MemCell.o_RX_Byte[7] ));
 sg13g2_dfrbp_1 _5025_ (.CLK(net767),
    .RESET_B(net29),
    .D(_0263_),
    .Q_N(_2598_),
    .Q(\spi_module.r_Temp_RX_Byte[0] ));
 sg13g2_dfrbp_1 _5026_ (.CLK(net767),
    .RESET_B(net28),
    .D(_0264_),
    .Q_N(_2597_),
    .Q(\spi_module.r_Temp_RX_Byte[1] ));
 sg13g2_dfrbp_1 _5027_ (.CLK(net766),
    .RESET_B(net27),
    .D(_0265_),
    .Q_N(_2596_),
    .Q(\spi_module.r_Temp_RX_Byte[2] ));
 sg13g2_dfrbp_1 _5028_ (.CLK(net765),
    .RESET_B(net26),
    .D(_0266_),
    .Q_N(_2595_),
    .Q(\spi_module.r_Temp_RX_Byte[3] ));
 sg13g2_dfrbp_1 _5029_ (.CLK(net765),
    .RESET_B(net25),
    .D(_0267_),
    .Q_N(_2594_),
    .Q(\spi_module.r_Temp_RX_Byte[4] ));
 sg13g2_dfrbp_1 _5030_ (.CLK(net765),
    .RESET_B(net24),
    .D(_0268_),
    .Q_N(_2593_),
    .Q(\spi_module.r_Temp_RX_Byte[5] ));
 sg13g2_dfrbp_1 _5031_ (.CLK(net765),
    .RESET_B(net15),
    .D(_0269_),
    .Q_N(_2622_),
    .Q(\spi_module.r_Temp_RX_Byte[6] ));
 sg13g2_dfrbp_1 _5032_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net837),
    .D(\spi_module.r_RX_Done ),
    .Q_N(_2592_),
    .Q(\spi_module.r2_RX_Done ));
 sg13g2_dfrbp_1 _5033_ (.CLK(net767),
    .RESET_B(net23),
    .D(_0270_),
    .Q_N(_2591_),
    .Q(\spi_module.r_RX_Byte[0] ));
 sg13g2_dfrbp_1 _5034_ (.CLK(net767),
    .RESET_B(net22),
    .D(_0271_),
    .Q_N(_2590_),
    .Q(\spi_module.r_RX_Byte[1] ));
 sg13g2_dfrbp_1 _5035_ (.CLK(net767),
    .RESET_B(net21),
    .D(_0272_),
    .Q_N(_2589_),
    .Q(\spi_module.r_RX_Byte[2] ));
 sg13g2_dfrbp_1 _5036_ (.CLK(net767),
    .RESET_B(net20),
    .D(_0273_),
    .Q_N(_2588_),
    .Q(\spi_module.r_RX_Byte[3] ));
 sg13g2_dfrbp_1 _5037_ (.CLK(net765),
    .RESET_B(net19),
    .D(_0274_),
    .Q_N(_2587_),
    .Q(\spi_module.r_RX_Byte[4] ));
 sg13g2_dfrbp_1 _5038_ (.CLK(net765),
    .RESET_B(net18),
    .D(_0275_),
    .Q_N(_2586_),
    .Q(\spi_module.r_RX_Byte[5] ));
 sg13g2_dfrbp_1 _5039_ (.CLK(net765),
    .RESET_B(net17),
    .D(_0276_),
    .Q_N(_2585_),
    .Q(\spi_module.r_RX_Byte[6] ));
 sg13g2_dfrbp_1 _5040_ (.CLK(net765),
    .RESET_B(net16),
    .D(_0277_),
    .Q_N(_2584_),
    .Q(\spi_module.r_RX_Byte[7] ));
 sg13g2_dfrbp_1 _5041_ (.CLK(net766),
    .RESET_B(_0222_),
    .D(_0278_),
    .Q_N(_2583_),
    .Q(\spi_module.r_RX_Done ));
 sg13g2_dfrbp_1 _5042_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net823),
    .D(_0279_),
    .Q_N(_2582_),
    .Q(\MemCell.dc2_reg[3][0] ));
 sg13g2_dfrbp_1 _5043_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net822),
    .D(_0280_),
    .Q_N(_2581_),
    .Q(\MemCell.dc2_reg[3][1] ));
 sg13g2_dfrbp_1 _5044_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net822),
    .D(_0281_),
    .Q_N(_2580_),
    .Q(\MemCell.dc2_reg[3][2] ));
 sg13g2_dfrbp_1 _5045_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net823),
    .D(_0282_),
    .Q_N(_2579_),
    .Q(\MemCell.dc2_reg[3][3] ));
 sg13g2_dfrbp_1 _5046_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net823),
    .D(_0283_),
    .Q_N(_2578_),
    .Q(\MemCell.dc2_reg[3][4] ));
 sg13g2_dfrbp_1 _5047_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net823),
    .D(_0284_),
    .Q_N(_2577_),
    .Q(\MemCell.dc2_reg[3][5] ));
 sg13g2_dfrbp_1 _5048_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net822),
    .D(_0285_),
    .Q_N(_2576_),
    .Q(\MemCell.dc2_reg[3][6] ));
 sg13g2_dfrbp_1 _5049_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net822),
    .D(_0286_),
    .Q_N(_2575_),
    .Q(\MemCell.dc2_reg[3][7] ));
 sg13g2_dfrbp_1 _5050_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net805),
    .D(_0287_),
    .Q_N(_2574_),
    .Q(\MemCell.dc3_reg[2][0] ));
 sg13g2_dfrbp_1 _5051_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net805),
    .D(_0288_),
    .Q_N(_2573_),
    .Q(\MemCell.dc3_reg[2][1] ));
 sg13g2_dfrbp_1 _5052_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net805),
    .D(_0289_),
    .Q_N(_2572_),
    .Q(\MemCell.dc3_reg[2][2] ));
 sg13g2_dfrbp_1 _5053_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net805),
    .D(_0290_),
    .Q_N(_2571_),
    .Q(\MemCell.dc3_reg[2][3] ));
 sg13g2_dfrbp_1 _5054_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net805),
    .D(net117),
    .Q_N(_2570_),
    .Q(\MemCell.dc3_reg[2][4] ));
 sg13g2_dfrbp_1 _5055_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net805),
    .D(_0292_),
    .Q_N(_2569_),
    .Q(\MemCell.dc3_reg[2][5] ));
 sg13g2_dfrbp_1 _5056_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net805),
    .D(_0293_),
    .Q_N(_2568_),
    .Q(\MemCell.dc3_reg[2][6] ));
 sg13g2_dfrbp_1 _5057_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net805),
    .D(_0294_),
    .Q_N(_2567_),
    .Q(\MemCell.dc3_reg[2][7] ));
 sg13g2_dfrbp_1 _5058_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net845),
    .D(_0295_),
    .Q_N(_2566_),
    .Q(\MemCell.dc2_reg[2][0] ));
 sg13g2_dfrbp_1 _5059_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net845),
    .D(_0296_),
    .Q_N(_2565_),
    .Q(\MemCell.dc2_reg[2][1] ));
 sg13g2_dfrbp_1 _5060_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net846),
    .D(_0297_),
    .Q_N(_2564_),
    .Q(\MemCell.dc2_reg[2][2] ));
 sg13g2_dfrbp_1 _5061_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net845),
    .D(_0298_),
    .Q_N(_2563_),
    .Q(\MemCell.dc2_reg[2][3] ));
 sg13g2_dfrbp_1 _5062_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net846),
    .D(_0299_),
    .Q_N(_2562_),
    .Q(\MemCell.dc2_reg[2][4] ));
 sg13g2_dfrbp_1 _5063_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net845),
    .D(_0300_),
    .Q_N(_2561_),
    .Q(\MemCell.dc2_reg[2][5] ));
 sg13g2_dfrbp_1 _5064_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net845),
    .D(_0301_),
    .Q_N(_2560_),
    .Q(\MemCell.dc2_reg[2][6] ));
 sg13g2_dfrbp_1 _5065_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net845),
    .D(_0302_),
    .Q_N(_2559_),
    .Q(\MemCell.dc2_reg[2][7] ));
 sg13g2_dfrbp_1 _5066_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net854),
    .D(_0303_),
    .Q_N(_2558_),
    .Q(\MemCell.dc2_reg[1][0] ));
 sg13g2_dfrbp_1 _5067_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net848),
    .D(_0304_),
    .Q_N(_2557_),
    .Q(\MemCell.dc2_reg[1][1] ));
 sg13g2_dfrbp_1 _5068_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net847),
    .D(_0305_),
    .Q_N(_2556_),
    .Q(\MemCell.dc2_reg[1][2] ));
 sg13g2_dfrbp_1 _5069_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net848),
    .D(_0306_),
    .Q_N(_2555_),
    .Q(\MemCell.dc2_reg[1][3] ));
 sg13g2_dfrbp_1 _5070_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net855),
    .D(_0307_),
    .Q_N(_2554_),
    .Q(\MemCell.dc2_reg[1][4] ));
 sg13g2_dfrbp_1 _5071_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net847),
    .D(_0308_),
    .Q_N(_2553_),
    .Q(\MemCell.dc2_reg[1][5] ));
 sg13g2_dfrbp_1 _5072_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net855),
    .D(_0309_),
    .Q_N(_2552_),
    .Q(\MemCell.dc2_reg[1][6] ));
 sg13g2_dfrbp_1 _5073_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net847),
    .D(_0310_),
    .Q_N(_2551_),
    .Q(\MemCell.dc2_reg[1][7] ));
 sg13g2_dfrbp_1 _5074_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net857),
    .D(_0311_),
    .Q_N(_2550_),
    .Q(\MemCell.dc2_reg[0][0] ));
 sg13g2_dfrbp_1 _5075_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net856),
    .D(_0312_),
    .Q_N(_2549_),
    .Q(\MemCell.dc2_reg[0][1] ));
 sg13g2_dfrbp_1 _5076_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net856),
    .D(_0313_),
    .Q_N(_2548_),
    .Q(\MemCell.dc2_reg[0][2] ));
 sg13g2_dfrbp_1 _5077_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net857),
    .D(net356),
    .Q_N(_2547_),
    .Q(\MemCell.dc2_reg[0][3] ));
 sg13g2_dfrbp_1 _5078_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net857),
    .D(_0315_),
    .Q_N(_2546_),
    .Q(\MemCell.dc2_reg[0][4] ));
 sg13g2_dfrbp_1 _5079_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net855),
    .D(_0316_),
    .Q_N(_2545_),
    .Q(\MemCell.dc2_reg[0][5] ));
 sg13g2_dfrbp_1 _5080_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net854),
    .D(_0317_),
    .Q_N(_2544_),
    .Q(\MemCell.dc2_reg[0][6] ));
 sg13g2_dfrbp_1 _5081_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net855),
    .D(_0318_),
    .Q_N(_2543_),
    .Q(\MemCell.dc2_reg[0][7] ));
 sg13g2_dfrbp_1 _5082_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net811),
    .D(_0319_),
    .Q_N(_2542_),
    .Q(\MemCell.dc1_reg[3][0] ));
 sg13g2_dfrbp_1 _5083_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net811),
    .D(_0320_),
    .Q_N(_2541_),
    .Q(\MemCell.dc1_reg[3][1] ));
 sg13g2_dfrbp_1 _5084_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net811),
    .D(_0321_),
    .Q_N(_2540_),
    .Q(\MemCell.dc1_reg[3][2] ));
 sg13g2_dfrbp_1 _5085_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net811),
    .D(_0322_),
    .Q_N(_2539_),
    .Q(\MemCell.dc1_reg[3][3] ));
 sg13g2_dfrbp_1 _5086_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net811),
    .D(_0323_),
    .Q_N(_2538_),
    .Q(\MemCell.dc1_reg[3][4] ));
 sg13g2_dfrbp_1 _5087_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net811),
    .D(_0324_),
    .Q_N(_2537_),
    .Q(\MemCell.dc1_reg[3][5] ));
 sg13g2_dfrbp_1 _5088_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net811),
    .D(_0325_),
    .Q_N(_2536_),
    .Q(\MemCell.dc1_reg[3][6] ));
 sg13g2_dfrbp_1 _5089_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net811),
    .D(_0326_),
    .Q_N(_2535_),
    .Q(\MemCell.dc1_reg[3][7] ));
 sg13g2_dfrbp_1 _5090_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net800),
    .D(_0327_),
    .Q_N(_2534_),
    .Q(\MemCell.dc1_reg[2][0] ));
 sg13g2_dfrbp_1 _5091_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net800),
    .D(_0328_),
    .Q_N(_2533_),
    .Q(\MemCell.dc1_reg[2][1] ));
 sg13g2_dfrbp_1 _5092_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net800),
    .D(_0329_),
    .Q_N(_2532_),
    .Q(\MemCell.dc1_reg[2][2] ));
 sg13g2_dfrbp_1 _5093_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net800),
    .D(_0330_),
    .Q_N(_2531_),
    .Q(\MemCell.dc1_reg[2][3] ));
 sg13g2_dfrbp_1 _5094_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net801),
    .D(_0331_),
    .Q_N(_2530_),
    .Q(\MemCell.dc1_reg[2][4] ));
 sg13g2_dfrbp_1 _5095_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net801),
    .D(net347),
    .Q_N(_2529_),
    .Q(\MemCell.dc1_reg[2][5] ));
 sg13g2_dfrbp_1 _5096_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net801),
    .D(_0333_),
    .Q_N(_2528_),
    .Q(\MemCell.dc1_reg[2][6] ));
 sg13g2_dfrbp_1 _5097_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net801),
    .D(net279),
    .Q_N(_2527_),
    .Q(\MemCell.dc1_reg[2][7] ));
 sg13g2_dfrbp_1 _5098_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net798),
    .D(_0335_),
    .Q_N(_2526_),
    .Q(\MemCell.dc1_reg[1][0] ));
 sg13g2_dfrbp_1 _5099_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net798),
    .D(_0336_),
    .Q_N(_2525_),
    .Q(\MemCell.dc1_reg[1][1] ));
 sg13g2_dfrbp_1 _5100_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net798),
    .D(_0337_),
    .Q_N(_2524_),
    .Q(\MemCell.dc1_reg[1][2] ));
 sg13g2_dfrbp_1 _5101_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net798),
    .D(_0338_),
    .Q_N(_2523_),
    .Q(\MemCell.dc1_reg[1][3] ));
 sg13g2_dfrbp_1 _5102_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net796),
    .D(_0339_),
    .Q_N(_2522_),
    .Q(\MemCell.dc1_reg[1][4] ));
 sg13g2_dfrbp_1 _5103_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net796),
    .D(_0340_),
    .Q_N(_2521_),
    .Q(\MemCell.dc1_reg[1][5] ));
 sg13g2_dfrbp_1 _5104_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net796),
    .D(_0341_),
    .Q_N(_2520_),
    .Q(\MemCell.dc1_reg[1][6] ));
 sg13g2_dfrbp_1 _5105_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net796),
    .D(_0342_),
    .Q_N(_2519_),
    .Q(\MemCell.dc1_reg[1][7] ));
 sg13g2_dfrbp_1 _5106_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net796),
    .D(_0343_),
    .Q_N(_2518_),
    .Q(\MemCell.dc1_reg[0][0] ));
 sg13g2_dfrbp_1 _5107_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net796),
    .D(_0344_),
    .Q_N(_2517_),
    .Q(\MemCell.dc1_reg[0][1] ));
 sg13g2_dfrbp_1 _5108_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net796),
    .D(_0345_),
    .Q_N(_2516_),
    .Q(\MemCell.dc1_reg[0][2] ));
 sg13g2_dfrbp_1 _5109_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net796),
    .D(_0346_),
    .Q_N(_2515_),
    .Q(\MemCell.dc1_reg[0][3] ));
 sg13g2_dfrbp_1 _5110_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net800),
    .D(_0347_),
    .Q_N(_2514_),
    .Q(\MemCell.dc1_reg[0][4] ));
 sg13g2_dfrbp_1 _5111_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net800),
    .D(_0348_),
    .Q_N(_2513_),
    .Q(\MemCell.dc1_reg[0][5] ));
 sg13g2_dfrbp_1 _5112_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net797),
    .D(_0349_),
    .Q_N(_2512_),
    .Q(\MemCell.dc1_reg[0][6] ));
 sg13g2_dfrbp_1 _5113_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net797),
    .D(_0350_),
    .Q_N(_2511_),
    .Q(\MemCell.dc1_reg[0][7] ));
 sg13g2_dfrbp_1 _5114_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net854),
    .D(_0351_),
    .Q_N(_2510_),
    .Q(\MemCell.prescale_reg[3][0] ));
 sg13g2_dfrbp_1 _5115_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net854),
    .D(_0352_),
    .Q_N(_2509_),
    .Q(\MemCell.prescale_reg[3][1] ));
 sg13g2_dfrbp_1 _5116_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net854),
    .D(_0353_),
    .Q_N(_2508_),
    .Q(\MemCell.prescale_reg[3][2] ));
 sg13g2_dfrbp_1 _5117_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net854),
    .D(_0354_),
    .Q_N(_2507_),
    .Q(\MemCell.prescale_reg[3][3] ));
 sg13g2_dfrbp_1 _5118_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net856),
    .D(_0355_),
    .Q_N(_2506_),
    .Q(\MemCell.prescale_reg[3][4] ));
 sg13g2_dfrbp_1 _5119_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net857),
    .D(_0356_),
    .Q_N(_2505_),
    .Q(\MemCell.prescale_reg[3][5] ));
 sg13g2_dfrbp_1 _5120_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net857),
    .D(_0357_),
    .Q_N(_2504_),
    .Q(\MemCell.prescale_reg[3][6] ));
 sg13g2_dfrbp_1 _5121_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net857),
    .D(_0358_),
    .Q_N(_2503_),
    .Q(\MemCell.prescale_reg[3][7] ));
 sg13g2_dfrbp_1 _5122_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net846),
    .D(_0359_),
    .Q_N(_2502_),
    .Q(\MemCell.prescale_reg[2][0] ));
 sg13g2_dfrbp_1 _5123_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net846),
    .D(_0360_),
    .Q_N(_2501_),
    .Q(\MemCell.prescale_reg[2][1] ));
 sg13g2_dfrbp_1 _5124_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net846),
    .D(_0361_),
    .Q_N(_2500_),
    .Q(\MemCell.prescale_reg[2][2] ));
 sg13g2_dfrbp_1 _5125_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net849),
    .D(_0362_),
    .Q_N(_2499_),
    .Q(\MemCell.prescale_reg[2][3] ));
 sg13g2_dfrbp_1 _5126_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net847),
    .D(_0363_),
    .Q_N(_2498_),
    .Q(\MemCell.prescale_reg[2][4] ));
 sg13g2_dfrbp_1 _5127_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net847),
    .D(_0364_),
    .Q_N(_2497_),
    .Q(\MemCell.prescale_reg[2][5] ));
 sg13g2_dfrbp_1 _5128_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net851),
    .D(_0365_),
    .Q_N(_2496_),
    .Q(\MemCell.prescale_reg[2][6] ));
 sg13g2_dfrbp_1 _5129_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net847),
    .D(_0366_),
    .Q_N(_2495_),
    .Q(\MemCell.prescale_reg[2][7] ));
 sg13g2_dfrbp_1 _5130_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net830),
    .D(_0367_),
    .Q_N(_2494_),
    .Q(\MemCell.dc3_reg[1][0] ));
 sg13g2_dfrbp_1 _5131_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net830),
    .D(_0368_),
    .Q_N(_2493_),
    .Q(\MemCell.dc3_reg[1][1] ));
 sg13g2_dfrbp_1 _5132_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net830),
    .D(_0369_),
    .Q_N(_2492_),
    .Q(\MemCell.dc3_reg[1][2] ));
 sg13g2_dfrbp_1 _5133_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net830),
    .D(_0370_),
    .Q_N(_2491_),
    .Q(\MemCell.dc3_reg[1][3] ));
 sg13g2_dfrbp_1 _5134_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net832),
    .D(_0371_),
    .Q_N(_2490_),
    .Q(\MemCell.dc3_reg[1][4] ));
 sg13g2_dfrbp_1 _5135_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net832),
    .D(_0372_),
    .Q_N(_2489_),
    .Q(\MemCell.dc3_reg[1][5] ));
 sg13g2_dfrbp_1 _5136_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net832),
    .D(_0373_),
    .Q_N(_2488_),
    .Q(\MemCell.dc3_reg[1][6] ));
 sg13g2_dfrbp_1 _5137_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net832),
    .D(_0374_),
    .Q_N(_2487_),
    .Q(\MemCell.dc3_reg[1][7] ));
 sg13g2_dfrbp_1 _5138_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net821),
    .D(_0375_),
    .Q_N(_2486_),
    .Q(\MemCell.prescale_reg[1][0] ));
 sg13g2_dfrbp_1 _5139_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net821),
    .D(_0376_),
    .Q_N(_2485_),
    .Q(\MemCell.prescale_reg[1][1] ));
 sg13g2_dfrbp_1 _5140_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net821),
    .D(_0377_),
    .Q_N(_2484_),
    .Q(\MemCell.prescale_reg[1][2] ));
 sg13g2_dfrbp_1 _5141_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net821),
    .D(_0378_),
    .Q_N(_2483_),
    .Q(\MemCell.prescale_reg[1][3] ));
 sg13g2_dfrbp_1 _5142_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net823),
    .D(net438),
    .Q_N(_2482_),
    .Q(\MemCell.prescale_reg[1][4] ));
 sg13g2_dfrbp_1 _5143_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net823),
    .D(_0380_),
    .Q_N(_2481_),
    .Q(\MemCell.prescale_reg[1][5] ));
 sg13g2_dfrbp_1 _5144_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net827),
    .D(net396),
    .Q_N(_2480_),
    .Q(\MemCell.prescale_reg[1][6] ));
 sg13g2_dfrbp_1 _5145_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net827),
    .D(net349),
    .Q_N(_2479_),
    .Q(\MemCell.prescale_reg[1][7] ));
 sg13g2_dfrbp_1 _5146_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net812),
    .D(_0383_),
    .Q_N(_2478_),
    .Q(\MemCell.prescale_reg[0][0] ));
 sg13g2_dfrbp_1 _5147_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net812),
    .D(_0384_),
    .Q_N(_2477_),
    .Q(\MemCell.prescale_reg[0][1] ));
 sg13g2_dfrbp_1 _5148_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net812),
    .D(_0385_),
    .Q_N(_2476_),
    .Q(\MemCell.prescale_reg[0][2] ));
 sg13g2_dfrbp_1 _5149_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net816),
    .D(_0386_),
    .Q_N(_2475_),
    .Q(\MemCell.prescale_reg[0][3] ));
 sg13g2_dfrbp_1 _5150_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net814),
    .D(_0387_),
    .Q_N(_2474_),
    .Q(\MemCell.prescale_reg[0][4] ));
 sg13g2_dfrbp_1 _5151_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net814),
    .D(_0388_),
    .Q_N(_2473_),
    .Q(\MemCell.prescale_reg[0][5] ));
 sg13g2_dfrbp_1 _5152_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net814),
    .D(_0389_),
    .Q_N(_2472_),
    .Q(\MemCell.prescale_reg[0][6] ));
 sg13g2_dfrbp_1 _5153_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net813),
    .D(_0390_),
    .Q_N(_2471_),
    .Q(\MemCell.prescale_reg[0][7] ));
 sg13g2_dfrbp_1 _5154_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net808),
    .D(_0391_),
    .Q_N(_2470_),
    .Q(\MemCell.counter_value[24] ));
 sg13g2_dfrbp_1 _5155_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net809),
    .D(_0392_),
    .Q_N(_2469_),
    .Q(\MemCell.counter_value[25] ));
 sg13g2_dfrbp_1 _5156_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net809),
    .D(_0393_),
    .Q_N(_2468_),
    .Q(\MemCell.counter_value[26] ));
 sg13g2_dfrbp_1 _5157_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net808),
    .D(_0394_),
    .Q_N(_2467_),
    .Q(\MemCell.counter_value[27] ));
 sg13g2_dfrbp_1 _5158_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net820),
    .D(_0395_),
    .Q_N(_2466_),
    .Q(\MemCell.counter_value[28] ));
 sg13g2_dfrbp_1 _5159_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net820),
    .D(_0396_),
    .Q_N(_2465_),
    .Q(\MemCell.counter_value[29] ));
 sg13g2_dfrbp_1 _5160_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net820),
    .D(_0397_),
    .Q_N(_2464_),
    .Q(\MemCell.counter_value[30] ));
 sg13g2_dfrbp_1 _5161_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net820),
    .D(_0398_),
    .Q_N(_2463_),
    .Q(\MemCell.counter_value[31] ));
 sg13g2_dfrbp_1 _5162_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net808),
    .D(_0399_),
    .Q_N(_2462_),
    .Q(\MemCell.counter_value[16] ));
 sg13g2_dfrbp_1 _5163_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net809),
    .D(_0400_),
    .Q_N(_2461_),
    .Q(\MemCell.counter_value[17] ));
 sg13g2_dfrbp_1 _5164_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net808),
    .D(_0401_),
    .Q_N(_2460_),
    .Q(\MemCell.counter_value[18] ));
 sg13g2_dfrbp_1 _5165_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net808),
    .D(_0402_),
    .Q_N(_2459_),
    .Q(\MemCell.counter_value[19] ));
 sg13g2_dfrbp_1 _5166_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net809),
    .D(_0403_),
    .Q_N(_2458_),
    .Q(\MemCell.counter_value[20] ));
 sg13g2_dfrbp_1 _5167_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net809),
    .D(_0404_),
    .Q_N(_2457_),
    .Q(\MemCell.counter_value[21] ));
 sg13g2_dfrbp_1 _5168_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net809),
    .D(_0405_),
    .Q_N(_2456_),
    .Q(\MemCell.counter_value[22] ));
 sg13g2_dfrbp_1 _5169_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net809),
    .D(_0406_),
    .Q_N(_2455_),
    .Q(\MemCell.counter_value[23] ));
 sg13g2_dfrbp_1 _5170_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net807),
    .D(_0407_),
    .Q_N(_2454_),
    .Q(\MemCell.counter_value[8] ));
 sg13g2_dfrbp_1 _5171_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net807),
    .D(_0408_),
    .Q_N(_2453_),
    .Q(\MemCell.counter_value[9] ));
 sg13g2_dfrbp_1 _5172_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net807),
    .D(_0409_),
    .Q_N(_2452_),
    .Q(\MemCell.counter_value[10] ));
 sg13g2_dfrbp_1 _5173_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net807),
    .D(_0410_),
    .Q_N(_2451_),
    .Q(\MemCell.counter_value[11] ));
 sg13g2_dfrbp_1 _5174_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net835),
    .D(_0411_),
    .Q_N(_2450_),
    .Q(\MemCell.counter_value[12] ));
 sg13g2_dfrbp_1 _5175_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net835),
    .D(_0412_),
    .Q_N(_2449_),
    .Q(\MemCell.counter_value[13] ));
 sg13g2_dfrbp_1 _5176_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net834),
    .D(_0413_),
    .Q_N(_2448_),
    .Q(\MemCell.counter_value[14] ));
 sg13g2_dfrbp_1 _5177_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net807),
    .D(_0414_),
    .Q_N(_2447_),
    .Q(\MemCell.counter_value[15] ));
 sg13g2_dfrbp_1 _5178_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net838),
    .D(net182),
    .Q_N(_2446_),
    .Q(\MemCell.counter_value[0] ));
 sg13g2_dfrbp_1 _5179_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net838),
    .D(net297),
    .Q_N(_2445_),
    .Q(\MemCell.counter_value[1] ));
 sg13g2_dfrbp_1 _5180_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net838),
    .D(net202),
    .Q_N(_2444_),
    .Q(\MemCell.counter_value[2] ));
 sg13g2_dfrbp_1 _5181_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net838),
    .D(_0418_),
    .Q_N(_2443_),
    .Q(\MemCell.counter_value[3] ));
 sg13g2_dfrbp_1 _5182_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net838),
    .D(_0419_),
    .Q_N(_2442_),
    .Q(\MemCell.counter_value[4] ));
 sg13g2_dfrbp_1 _5183_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net838),
    .D(_0420_),
    .Q_N(_2441_),
    .Q(\MemCell.counter_value[5] ));
 sg13g2_dfrbp_1 _5184_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net838),
    .D(_0421_),
    .Q_N(_2440_),
    .Q(\MemCell.counter_value[6] ));
 sg13g2_dfrbp_1 _5185_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net838),
    .D(_0422_),
    .Q_N(_2439_),
    .Q(\MemCell.counter_value[7] ));
 sg13g2_dfrbp_1 _5186_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net856),
    .D(net422),
    .Q_N(_2438_),
    .Q(\MemCell.enable_pwm ));
 sg13g2_dfrbp_1 _5187_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net840),
    .D(_0424_),
    .Q_N(_2437_),
    .Q(\MemCell.counter[0] ));
 sg13g2_dfrbp_1 _5188_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net840),
    .D(_0425_),
    .Q_N(_2436_),
    .Q(\MemCell.counter[1] ));
 sg13g2_dfrbp_1 _5189_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net836),
    .D(net219),
    .Q_N(_2435_),
    .Q(\MemCell.dc3_reg[0][0] ));
 sg13g2_dfrbp_1 _5190_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net836),
    .D(net316),
    .Q_N(_2434_),
    .Q(\MemCell.dc3_reg[0][1] ));
 sg13g2_dfrbp_1 _5191_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net836),
    .D(net289),
    .Q_N(_2433_),
    .Q(\MemCell.dc3_reg[0][2] ));
 sg13g2_dfrbp_1 _5192_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net836),
    .D(_0429_),
    .Q_N(_2432_),
    .Q(\MemCell.dc3_reg[0][3] ));
 sg13g2_dfrbp_1 _5193_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net836),
    .D(_0430_),
    .Q_N(_2431_),
    .Q(\MemCell.dc3_reg[0][4] ));
 sg13g2_dfrbp_1 _5194_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net836),
    .D(_0431_),
    .Q_N(_2430_),
    .Q(\MemCell.dc3_reg[0][5] ));
 sg13g2_dfrbp_1 _5195_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net836),
    .D(_0432_),
    .Q_N(_2429_),
    .Q(\MemCell.dc3_reg[0][6] ));
 sg13g2_dfrbp_1 _5196_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net836),
    .D(_0433_),
    .Q_N(_2623_),
    .Q(\MemCell.dc3_reg[0][7] ));
 sg13g2_dfrbp_1 _5197_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net841),
    .D(net560),
    .Q_N(_2624_),
    .Q(\MemCell.curr_state[0] ));
 sg13g2_dfrbp_1 _5198_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net841),
    .D(\MemCell.next_state[1] ),
    .Q_N(_2625_),
    .Q(\MemCell.curr_state[1] ));
 sg13g2_dfrbp_1 _5199_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net840),
    .D(\MemCell.next_state[2] ),
    .Q_N(_0144_),
    .Q(\MemCell.curr_state[2] ));
 sg13g2_dfrbp_1 _5200_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net832),
    .D(_0434_),
    .Q_N(_2428_),
    .Q(\pwm_module.counter2[0] ));
 sg13g2_dfrbp_1 _5201_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net832),
    .D(_0435_),
    .Q_N(_0143_),
    .Q(\pwm_module.counter2[1] ));
 sg13g2_dfrbp_1 _5202_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net837),
    .D(_0436_),
    .Q_N(_2427_),
    .Q(\pwm_module.counter2[2] ));
 sg13g2_dfrbp_1 _5203_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net833),
    .D(net76),
    .Q_N(_0142_),
    .Q(\pwm_module.counter2[3] ));
 sg13g2_dfrbp_1 _5204_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net837),
    .D(_0438_),
    .Q_N(_0141_),
    .Q(\pwm_module.counter2[4] ));
 sg13g2_dfrbp_1 _5205_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net837),
    .D(net342),
    .Q_N(_0140_),
    .Q(\pwm_module.counter2[5] ));
 sg13g2_dfrbp_1 _5206_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net832),
    .D(net261),
    .Q_N(_0139_),
    .Q(\pwm_module.counter2[6] ));
 sg13g2_dfrbp_1 _5207_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net832),
    .D(net217),
    .Q_N(_0138_),
    .Q(\pwm_module.counter2[7] ));
 sg13g2_dfrbp_1 _5208_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net830),
    .D(_0442_),
    .Q_N(_2426_),
    .Q(\pwm_module.counter2[8] ));
 sg13g2_dfrbp_1 _5209_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net830),
    .D(net148),
    .Q_N(_0137_),
    .Q(\pwm_module.counter2[9] ));
 sg13g2_dfrbp_1 _5210_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net830),
    .D(net301),
    .Q_N(_0136_),
    .Q(\pwm_module.counter2[10] ));
 sg13g2_dfrbp_1 _5211_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net830),
    .D(net78),
    .Q_N(_0135_),
    .Q(\pwm_module.counter2[11] ));
 sg13g2_dfrbp_1 _5212_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net831),
    .D(net94),
    .Q_N(_0134_),
    .Q(\pwm_module.counter2[12] ));
 sg13g2_dfrbp_1 _5213_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net831),
    .D(net128),
    .Q_N(_0133_),
    .Q(\pwm_module.counter2[13] ));
 sg13g2_dfrbp_1 _5214_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net831),
    .D(_0448_),
    .Q_N(_2425_),
    .Q(\pwm_module.counter2[14] ));
 sg13g2_dfrbp_1 _5215_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net831),
    .D(net47),
    .Q_N(_0132_),
    .Q(\pwm_module.counter2[15] ));
 sg13g2_dfrbp_1 _5216_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net834),
    .D(_0450_),
    .Q_N(_2424_),
    .Q(\pwm_module.counter2[16] ));
 sg13g2_dfrbp_1 _5217_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net831),
    .D(net90),
    .Q_N(_0131_),
    .Q(\pwm_module.counter2[17] ));
 sg13g2_dfrbp_1 _5218_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net834),
    .D(_0452_),
    .Q_N(_2423_),
    .Q(\pwm_module.counter2[18] ));
 sg13g2_dfrbp_1 _5219_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net831),
    .D(net65),
    .Q_N(_0130_),
    .Q(\pwm_module.counter2[19] ));
 sg13g2_dfrbp_1 _5220_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net810),
    .D(net304),
    .Q_N(_0129_),
    .Q(\pwm_module.counter2[20] ));
 sg13g2_dfrbp_1 _5221_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net810),
    .D(net210),
    .Q_N(_0128_),
    .Q(\pwm_module.counter2[21] ));
 sg13g2_dfrbp_1 _5222_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net834),
    .D(net482),
    .Q_N(_2422_),
    .Q(\pwm_module.counter2[22] ));
 sg13g2_dfrbp_1 _5223_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net810),
    .D(net63),
    .Q_N(_0127_),
    .Q(\pwm_module.counter2[23] ));
 sg13g2_dfrbp_1 _5224_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net806),
    .D(_0458_),
    .Q_N(_2421_),
    .Q(\pwm_module.counter2[24] ));
 sg13g2_dfrbp_1 _5225_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net806),
    .D(net92),
    .Q_N(_0126_),
    .Q(\pwm_module.counter2[25] ));
 sg13g2_dfrbp_1 _5226_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net807),
    .D(_0460_),
    .Q_N(_2420_),
    .Q(\pwm_module.counter2[26] ));
 sg13g2_dfrbp_1 _5227_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net808),
    .D(net67),
    .Q_N(_0125_),
    .Q(\pwm_module.counter2[27] ));
 sg13g2_dfrbp_1 _5228_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net806),
    .D(_0462_),
    .Q_N(_2419_),
    .Q(\pwm_module.counter2[28] ));
 sg13g2_dfrbp_1 _5229_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net808),
    .D(net86),
    .Q_N(_0124_),
    .Q(\pwm_module.counter2[29] ));
 sg13g2_dfrbp_1 _5230_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net807),
    .D(net185),
    .Q_N(_2418_),
    .Q(\pwm_module.counter2[30] ));
 sg13g2_dfrbp_1 _5231_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net807),
    .D(net49),
    .Q_N(_0168_),
    .Q(\pwm_module.counter2[31] ));
 sg13g2_dfrbp_1 _5232_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net816),
    .D(_0032_),
    .Q_N(_2626_),
    .Q(\pwm_module.prescaler1[0] ));
 sg13g2_dfrbp_1 _5233_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net816),
    .D(_0043_),
    .Q_N(_2627_),
    .Q(\pwm_module.prescaler1[1] ));
 sg13g2_dfrbp_1 _5234_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net816),
    .D(_0054_),
    .Q_N(_2628_),
    .Q(\pwm_module.prescaler1[2] ));
 sg13g2_dfrbp_1 _5235_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net816),
    .D(_0057_),
    .Q_N(_0169_),
    .Q(\pwm_module.prescaler1[3] ));
 sg13g2_dfrbp_1 _5236_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net817),
    .D(_0058_),
    .Q_N(_2629_),
    .Q(\pwm_module.prescaler1[4] ));
 sg13g2_dfrbp_1 _5237_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net816),
    .D(_0059_),
    .Q_N(_0170_),
    .Q(\pwm_module.prescaler1[5] ));
 sg13g2_dfrbp_1 _5238_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net818),
    .D(_0060_),
    .Q_N(_2630_),
    .Q(\pwm_module.prescaler1[6] ));
 sg13g2_dfrbp_1 _5239_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net818),
    .D(_0061_),
    .Q_N(_0171_),
    .Q(\pwm_module.prescaler1[7] ));
 sg13g2_dfrbp_1 _5240_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net818),
    .D(_0062_),
    .Q_N(_2631_),
    .Q(\pwm_module.prescaler1[8] ));
 sg13g2_dfrbp_1 _5241_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net818),
    .D(_0063_),
    .Q_N(_0172_),
    .Q(\pwm_module.prescaler1[9] ));
 sg13g2_dfrbp_1 _5242_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net826),
    .D(_0033_),
    .Q_N(_2632_),
    .Q(\pwm_module.prescaler1[10] ));
 sg13g2_dfrbp_1 _5243_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net825),
    .D(_0034_),
    .Q_N(_0173_),
    .Q(\pwm_module.prescaler1[11] ));
 sg13g2_dfrbp_1 _5244_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net828),
    .D(_0035_),
    .Q_N(_0174_),
    .Q(\pwm_module.prescaler1[12] ));
 sg13g2_dfrbp_1 _5245_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net827),
    .D(_0036_),
    .Q_N(_0175_),
    .Q(\pwm_module.prescaler1[13] ));
 sg13g2_dfrbp_1 _5246_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net828),
    .D(_0037_),
    .Q_N(_2633_),
    .Q(\pwm_module.prescaler1[14] ));
 sg13g2_dfrbp_1 _5247_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net828),
    .D(_0038_),
    .Q_N(_0176_),
    .Q(\pwm_module.prescaler1[15] ));
 sg13g2_dfrbp_1 _5248_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net850),
    .D(_0039_),
    .Q_N(_2634_),
    .Q(\pwm_module.prescaler1[16] ));
 sg13g2_dfrbp_1 _5249_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net850),
    .D(_0040_),
    .Q_N(_0177_),
    .Q(\pwm_module.prescaler1[17] ));
 sg13g2_dfrbp_1 _5250_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net850),
    .D(_0041_),
    .Q_N(_2635_),
    .Q(\pwm_module.prescaler1[18] ));
 sg13g2_dfrbp_1 _5251_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net849),
    .D(_0042_),
    .Q_N(_0178_),
    .Q(\pwm_module.prescaler1[19] ));
 sg13g2_dfrbp_1 _5252_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net852),
    .D(_0044_),
    .Q_N(_0179_),
    .Q(\pwm_module.prescaler1[20] ));
 sg13g2_dfrbp_1 _5253_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net852),
    .D(_0045_),
    .Q_N(_0180_),
    .Q(\pwm_module.prescaler1[21] ));
 sg13g2_dfrbp_1 _5254_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net851),
    .D(_0046_),
    .Q_N(_2636_),
    .Q(\pwm_module.prescaler1[22] ));
 sg13g2_dfrbp_1 _5255_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net852),
    .D(_0047_),
    .Q_N(_0181_),
    .Q(\pwm_module.prescaler1[23] ));
 sg13g2_dfrbp_1 _5256_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net860),
    .D(_0048_),
    .Q_N(_2637_),
    .Q(\pwm_module.prescaler1[24] ));
 sg13g2_dfrbp_1 _5257_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net860),
    .D(_0049_),
    .Q_N(_0182_),
    .Q(\pwm_module.prescaler1[25] ));
 sg13g2_dfrbp_1 _5258_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net860),
    .D(_0050_),
    .Q_N(_2638_),
    .Q(\pwm_module.prescaler1[26] ));
 sg13g2_dfrbp_1 _5259_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net860),
    .D(_0051_),
    .Q_N(_0183_),
    .Q(\pwm_module.prescaler1[27] ));
 sg13g2_dfrbp_1 _5260_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net860),
    .D(net444),
    .Q_N(_2639_),
    .Q(\pwm_module.prescaler1[28] ));
 sg13g2_dfrbp_1 _5261_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net860),
    .D(net101),
    .Q_N(_0184_),
    .Q(\pwm_module.prescaler1[29] ));
 sg13g2_dfrbp_1 _5262_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net860),
    .D(net82),
    .Q_N(_2640_),
    .Q(\pwm_module.prescaler1[30] ));
 sg13g2_dfrbp_1 _5263_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net860),
    .D(_0056_),
    .Q_N(_0185_),
    .Q(\pwm_module.prescaler1[31] ));
 sg13g2_dfrbp_1 _5264_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net856),
    .D(_0097_),
    .Q_N(_2641_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _5265_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net856),
    .D(_0096_),
    .Q_N(_2642_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _5266_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net812),
    .D(_0064_),
    .Q_N(_2643_),
    .Q(\pwm_module.prescaler2[0] ));
 sg13g2_dfrbp_1 _5267_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net812),
    .D(_0075_),
    .Q_N(_2644_),
    .Q(\pwm_module.prescaler2[1] ));
 sg13g2_dfrbp_1 _5268_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net815),
    .D(_0086_),
    .Q_N(_2645_),
    .Q(\pwm_module.prescaler2[2] ));
 sg13g2_dfrbp_1 _5269_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net816),
    .D(_0089_),
    .Q_N(_0186_),
    .Q(\pwm_module.prescaler2[3] ));
 sg13g2_dfrbp_1 _5270_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net818),
    .D(_0090_),
    .Q_N(_2646_),
    .Q(\pwm_module.prescaler2[4] ));
 sg13g2_dfrbp_1 _5271_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net818),
    .D(_0091_),
    .Q_N(_0187_),
    .Q(\pwm_module.prescaler2[5] ));
 sg13g2_dfrbp_1 _5272_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net818),
    .D(_0092_),
    .Q_N(_2647_),
    .Q(\pwm_module.prescaler2[6] ));
 sg13g2_dfrbp_1 _5273_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net813),
    .D(_0093_),
    .Q_N(_0188_),
    .Q(\pwm_module.prescaler2[7] ));
 sg13g2_dfrbp_1 _5274_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net813),
    .D(_0094_),
    .Q_N(_2648_),
    .Q(\pwm_module.prescaler2[8] ));
 sg13g2_dfrbp_1 _5275_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net825),
    .D(_0095_),
    .Q_N(_0189_),
    .Q(\pwm_module.prescaler2[9] ));
 sg13g2_dfrbp_1 _5276_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net825),
    .D(net545),
    .Q_N(_2649_),
    .Q(\pwm_module.prescaler2[10] ));
 sg13g2_dfrbp_1 _5277_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net825),
    .D(_0066_),
    .Q_N(_0190_),
    .Q(\pwm_module.prescaler2[11] ));
 sg13g2_dfrbp_1 _5278_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net825),
    .D(net37),
    .Q_N(_0191_),
    .Q(\pwm_module.prescaler2[12] ));
 sg13g2_dfrbp_1 _5279_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net825),
    .D(_0068_),
    .Q_N(_0192_),
    .Q(\pwm_module.prescaler2[13] ));
 sg13g2_dfrbp_1 _5280_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net827),
    .D(_0069_),
    .Q_N(_2650_),
    .Q(\pwm_module.prescaler2[14] ));
 sg13g2_dfrbp_1 _5281_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net827),
    .D(net41),
    .Q_N(_0193_),
    .Q(\pwm_module.prescaler2[15] ));
 sg13g2_dfrbp_1 _5282_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net827),
    .D(_0071_),
    .Q_N(_2651_),
    .Q(\pwm_module.prescaler2[16] ));
 sg13g2_dfrbp_1 _5283_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net849),
    .D(net43),
    .Q_N(_0194_),
    .Q(\pwm_module.prescaler2[17] ));
 sg13g2_dfrbp_1 _5284_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net849),
    .D(_0073_),
    .Q_N(_2652_),
    .Q(\pwm_module.prescaler2[18] ));
 sg13g2_dfrbp_1 _5285_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net849),
    .D(_0074_),
    .Q_N(_0195_),
    .Q(\pwm_module.prescaler2[19] ));
 sg13g2_dfrbp_1 _5286_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net851),
    .D(_0076_),
    .Q_N(_0196_),
    .Q(\pwm_module.prescaler2[20] ));
 sg13g2_dfrbp_1 _5287_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net851),
    .D(_0077_),
    .Q_N(_0197_),
    .Q(\pwm_module.prescaler2[21] ));
 sg13g2_dfrbp_1 _5288_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net851),
    .D(net511),
    .Q_N(_2653_),
    .Q(\pwm_module.prescaler2[22] ));
 sg13g2_dfrbp_1 _5289_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net851),
    .D(net55),
    .Q_N(_0198_),
    .Q(\pwm_module.prescaler2[23] ));
 sg13g2_dfrbp_1 _5290_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net861),
    .D(net411),
    .Q_N(_2654_),
    .Q(\pwm_module.prescaler2[24] ));
 sg13g2_dfrbp_1 _5291_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net861),
    .D(_0081_),
    .Q_N(_0199_),
    .Q(\pwm_module.prescaler2[25] ));
 sg13g2_dfrbp_1 _5292_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net861),
    .D(_0082_),
    .Q_N(_2655_),
    .Q(\pwm_module.prescaler2[26] ));
 sg13g2_dfrbp_1 _5293_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net861),
    .D(net245),
    .Q_N(_0200_),
    .Q(\pwm_module.prescaler2[27] ));
 sg13g2_dfrbp_1 _5294_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net859),
    .D(_0084_),
    .Q_N(_2656_),
    .Q(\pwm_module.prescaler2[28] ));
 sg13g2_dfrbp_1 _5295_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net862),
    .D(net57),
    .Q_N(_0201_),
    .Q(\pwm_module.prescaler2[29] ));
 sg13g2_dfrbp_1 _5296_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net862),
    .D(net518),
    .Q_N(_2657_),
    .Q(\pwm_module.prescaler2[30] ));
 sg13g2_dfrbp_1 _5297_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net859),
    .D(_0088_),
    .Q_N(_0123_),
    .Q(\pwm_module.prescaler2[31] ));
 sg13g2_dfrbp_1 _5298_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net804),
    .D(_0466_),
    .Q_N(_2417_),
    .Q(\MemCell.dc3_reg[3][0] ));
 sg13g2_dfrbp_1 _5299_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net804),
    .D(_0467_),
    .Q_N(_2416_),
    .Q(\MemCell.dc3_reg[3][1] ));
 sg13g2_dfrbp_1 _5300_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net804),
    .D(_0468_),
    .Q_N(_2415_),
    .Q(\MemCell.dc3_reg[3][2] ));
 sg13g2_dfrbp_1 _5301_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net804),
    .D(_0469_),
    .Q_N(_2414_),
    .Q(\MemCell.dc3_reg[3][3] ));
 sg13g2_dfrbp_1 _5302_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net804),
    .D(_0470_),
    .Q_N(_2413_),
    .Q(\MemCell.dc3_reg[3][4] ));
 sg13g2_dfrbp_1 _5303_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net804),
    .D(_0471_),
    .Q_N(_2412_),
    .Q(\MemCell.dc3_reg[3][5] ));
 sg13g2_dfrbp_1 _5304_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net804),
    .D(_0472_),
    .Q_N(_2411_),
    .Q(\MemCell.dc3_reg[3][6] ));
 sg13g2_dfrbp_1 _5305_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net804),
    .D(_0473_),
    .Q_N(_2658_),
    .Q(\MemCell.dc3_reg[3][7] ));
 sg13g2_dfrbp_1 _5306_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net840),
    .D(_0098_),
    .Q_N(_2410_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _5307_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net856),
    .D(_0474_),
    .Q_N(_2409_),
    .Q(\pwm_module.counter1[0] ));
 sg13g2_dfrbp_1 _5308_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net841),
    .D(_0475_),
    .Q_N(_0122_),
    .Q(\pwm_module.counter1[1] ));
 sg13g2_dfrbp_1 _5309_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net839),
    .D(_0476_),
    .Q_N(_2408_),
    .Q(\pwm_module.counter1[2] ));
 sg13g2_dfrbp_1 _5310_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net841),
    .D(net153),
    .Q_N(_0121_),
    .Q(\pwm_module.counter1[3] ));
 sg13g2_dfrbp_1 _5311_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net856),
    .D(_0478_),
    .Q_N(_0120_),
    .Q(\pwm_module.counter1[4] ));
 sg13g2_dfrbp_1 _5312_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net854),
    .D(net478),
    .Q_N(_0119_),
    .Q(\pwm_module.counter1[5] ));
 sg13g2_dfrbp_1 _5313_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net839),
    .D(net255),
    .Q_N(_0118_),
    .Q(\pwm_module.counter1[6] ));
 sg13g2_dfrbp_1 _5314_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net839),
    .D(net234),
    .Q_N(_0117_),
    .Q(\pwm_module.counter1[7] ));
 sg13g2_dfrbp_1 _5315_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net854),
    .D(net550),
    .Q_N(_2407_),
    .Q(\pwm_module.counter1[8] ));
 sg13g2_dfrbp_1 _5316_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net839),
    .D(net110),
    .Q_N(_0116_),
    .Q(\pwm_module.counter1[9] ));
 sg13g2_dfrbp_1 _5317_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net835),
    .D(net360),
    .Q_N(_0115_),
    .Q(\pwm_module.counter1[10] ));
 sg13g2_dfrbp_1 _5318_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net835),
    .D(net88),
    .Q_N(_0114_),
    .Q(\pwm_module.counter1[11] ));
 sg13g2_dfrbp_1 _5319_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net835),
    .D(net195),
    .Q_N(_0113_),
    .Q(\pwm_module.counter1[12] ));
 sg13g2_dfrbp_1 _5320_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net835),
    .D(net121),
    .Q_N(_0112_),
    .Q(\pwm_module.counter1[13] ));
 sg13g2_dfrbp_1 _5321_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net835),
    .D(_0488_),
    .Q_N(_2406_),
    .Q(\pwm_module.counter1[14] ));
 sg13g2_dfrbp_1 _5322_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net835),
    .D(net107),
    .Q_N(_0111_),
    .Q(\pwm_module.counter1[15] ));
 sg13g2_dfrbp_1 _5323_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net847),
    .D(_0490_),
    .Q_N(_2405_),
    .Q(\pwm_module.counter1[16] ));
 sg13g2_dfrbp_1 _5324_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net834),
    .D(net96),
    .Q_N(_0110_),
    .Q(\pwm_module.counter1[17] ));
 sg13g2_dfrbp_1 _5325_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net847),
    .D(_0492_),
    .Q_N(_2404_),
    .Q(\pwm_module.counter1[18] ));
 sg13g2_dfrbp_1 _5326_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net834),
    .D(net69),
    .Q_N(_0109_),
    .Q(\pwm_module.counter1[19] ));
 sg13g2_dfrbp_1 _5327_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net834),
    .D(_0494_),
    .Q_N(_0108_),
    .Q(\pwm_module.counter1[20] ));
 sg13g2_dfrbp_1 _5328_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net834),
    .D(net213),
    .Q_N(_0107_),
    .Q(\pwm_module.counter1[21] ));
 sg13g2_dfrbp_1 _5329_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net845),
    .D(net231),
    .Q_N(_2403_),
    .Q(\pwm_module.counter1[22] ));
 sg13g2_dfrbp_1 _5330_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net845),
    .D(net59),
    .Q_N(_0106_),
    .Q(\pwm_module.counter1[23] ));
 sg13g2_dfrbp_1 _5331_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net822),
    .D(_0498_),
    .Q_N(_2402_),
    .Q(\pwm_module.counter1[24] ));
 sg13g2_dfrbp_1 _5332_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net822),
    .D(net163),
    .Q_N(_0105_),
    .Q(\pwm_module.counter1[25] ));
 sg13g2_dfrbp_1 _5333_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net822),
    .D(_0500_),
    .Q_N(_2401_),
    .Q(\pwm_module.counter1[26] ));
 sg13g2_dfrbp_1 _5334_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net822),
    .D(net84),
    .Q_N(_0104_),
    .Q(\pwm_module.counter1[27] ));
 sg13g2_dfrbp_1 _5335_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net820),
    .D(_0502_),
    .Q_N(_2400_),
    .Q(\pwm_module.counter1[28] ));
 sg13g2_dfrbp_1 _5336_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net820),
    .D(net160),
    .Q_N(_0103_),
    .Q(\pwm_module.counter1[29] ));
 sg13g2_dfrbp_1 _5337_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net820),
    .D(net309),
    .Q_N(_2399_),
    .Q(\pwm_module.counter1[30] ));
 sg13g2_dfrbp_1 _5338_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net820),
    .D(net39),
    .Q_N(_0202_),
    .Q(\pwm_module.counter1[31] ));
 sg13g2_dfrbp_1 _5339_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net817),
    .D(_0000_),
    .Q_N(_2659_),
    .Q(\pwm_module.prescaler0[0] ));
 sg13g2_dfrbp_1 _5340_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net817),
    .D(_0011_),
    .Q_N(_2660_),
    .Q(\pwm_module.prescaler0[1] ));
 sg13g2_dfrbp_1 _5341_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net817),
    .D(_0022_),
    .Q_N(_2661_),
    .Q(\pwm_module.prescaler0[2] ));
 sg13g2_dfrbp_1 _5342_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net817),
    .D(_0025_),
    .Q_N(_0203_),
    .Q(\pwm_module.prescaler0[3] ));
 sg13g2_dfrbp_1 _5343_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net817),
    .D(net319),
    .Q_N(_2662_),
    .Q(\pwm_module.prescaler0[4] ));
 sg13g2_dfrbp_1 _5344_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net816),
    .D(_0027_),
    .Q_N(_0204_),
    .Q(\pwm_module.prescaler0[5] ));
 sg13g2_dfrbp_1 _5345_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net818),
    .D(net276),
    .Q_N(_2663_),
    .Q(\pwm_module.prescaler0[6] ));
 sg13g2_dfrbp_1 _5346_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net819),
    .D(_0029_),
    .Q_N(_0205_),
    .Q(\pwm_module.prescaler0[7] ));
 sg13g2_dfrbp_1 _5347_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net826),
    .D(_0030_),
    .Q_N(_2664_),
    .Q(\pwm_module.prescaler0[8] ));
 sg13g2_dfrbp_1 _5348_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net826),
    .D(_0031_),
    .Q_N(_0206_),
    .Q(\pwm_module.prescaler0[9] ));
 sg13g2_dfrbp_1 _5349_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net826),
    .D(net461),
    .Q_N(_2665_),
    .Q(\pwm_module.prescaler0[10] ));
 sg13g2_dfrbp_1 _5350_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net826),
    .D(_0002_),
    .Q_N(_0207_),
    .Q(\pwm_module.prescaler0[11] ));
 sg13g2_dfrbp_1 _5351_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net825),
    .D(_0003_),
    .Q_N(_2666_),
    .Q(\pwm_module.prescaler0[12] ));
 sg13g2_dfrbp_1 _5352_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net825),
    .D(_0004_),
    .Q_N(_0208_),
    .Q(\pwm_module.prescaler0[13] ));
 sg13g2_dfrbp_1 _5353_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net827),
    .D(net406),
    .Q_N(_2667_),
    .Q(\pwm_module.prescaler0[14] ));
 sg13g2_dfrbp_1 _5354_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net827),
    .D(_0006_),
    .Q_N(_0209_),
    .Q(\pwm_module.prescaler0[15] ));
 sg13g2_dfrbp_1 _5355_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net850),
    .D(net378),
    .Q_N(_2668_),
    .Q(\pwm_module.prescaler0[16] ));
 sg13g2_dfrbp_1 _5356_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net849),
    .D(_0008_),
    .Q_N(_0210_),
    .Q(\pwm_module.prescaler0[17] ));
 sg13g2_dfrbp_1 _5357_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net849),
    .D(_0009_),
    .Q_N(_2669_),
    .Q(\pwm_module.prescaler0[18] ));
 sg13g2_dfrbp_1 _5358_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net849),
    .D(_0010_),
    .Q_N(_0211_),
    .Q(\pwm_module.prescaler0[19] ));
 sg13g2_dfrbp_1 _5359_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net851),
    .D(_0012_),
    .Q_N(_0212_),
    .Q(\pwm_module.prescaler0[20] ));
 sg13g2_dfrbp_1 _5360_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net851),
    .D(_0013_),
    .Q_N(_0213_),
    .Q(\pwm_module.prescaler0[21] ));
 sg13g2_dfrbp_1 _5361_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net852),
    .D(_0014_),
    .Q_N(_2670_),
    .Q(\pwm_module.prescaler0[22] ));
 sg13g2_dfrbp_1 _5362_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net852),
    .D(_0015_),
    .Q_N(_0214_),
    .Q(\pwm_module.prescaler0[23] ));
 sg13g2_dfrbp_1 _5363_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net861),
    .D(_0016_),
    .Q_N(_2671_),
    .Q(\pwm_module.prescaler0[24] ));
 sg13g2_dfrbp_1 _5364_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net861),
    .D(_0017_),
    .Q_N(_0215_),
    .Q(\pwm_module.prescaler0[25] ));
 sg13g2_dfrbp_1 _5365_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net861),
    .D(net488),
    .Q_N(_0216_),
    .Q(\pwm_module.prescaler0[26] ));
 sg13g2_dfrbp_1 _5366_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net861),
    .D(_0019_),
    .Q_N(_0217_),
    .Q(\pwm_module.prescaler0[27] ));
 sg13g2_dfrbp_1 _5367_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net859),
    .D(_0020_),
    .Q_N(_2672_),
    .Q(\pwm_module.prescaler0[28] ));
 sg13g2_dfrbp_1 _5368_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net859),
    .D(_0021_),
    .Q_N(_0218_),
    .Q(\pwm_module.prescaler0[29] ));
 sg13g2_dfrbp_1 _5369_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net859),
    .D(_0023_),
    .Q_N(_2673_),
    .Q(\pwm_module.prescaler0[30] ));
 sg13g2_dfrbp_1 _5370_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net859),
    .D(_0024_),
    .Q_N(_0102_),
    .Q(\pwm_module.prescaler0[31] ));
 sg13g2_tiehi _5040__16 (.L_HI(net16));
 sg13g2_tiehi _5039__17 (.L_HI(net17));
 sg13g2_tiehi _5038__18 (.L_HI(net18));
 sg13g2_tiehi _5037__19 (.L_HI(net19));
 sg13g2_tiehi _5036__20 (.L_HI(net20));
 sg13g2_tiehi _5035__21 (.L_HI(net21));
 sg13g2_tiehi _5034__22 (.L_HI(net22));
 sg13g2_tiehi _5033__23 (.L_HI(net23));
 sg13g2_tiehi _5030__24 (.L_HI(net24));
 sg13g2_tiehi _5029__25 (.L_HI(net25));
 sg13g2_tiehi _5028__26 (.L_HI(net26));
 sg13g2_tiehi _5027__27 (.L_HI(net27));
 sg13g2_tiehi _5026__28 (.L_HI(net28));
 sg13g2_tiehi _5025__29 (.L_HI(net29));
 sg13g2_tiehi tt_um_pwm_block_30 (.L_HI(net30));
 sg13g2_tiehi tt_um_pwm_block_31 (.L_HI(net31));
 sg13g2_tiehi tt_um_pwm_block_32 (.L_HI(net32));
 sg13g2_tiehi tt_um_pwm_block_33 (.L_HI(net33));
 sg13g2_tiehi tt_um_pwm_block_34 (.L_HI(net34));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_pwm_block_7 (.L_LO(net7));
 sg13g2_tielo tt_um_pwm_block_8 (.L_LO(net8));
 sg13g2_tielo tt_um_pwm_block_9 (.L_LO(net9));
 sg13g2_tielo tt_um_pwm_block_10 (.L_LO(net10));
 sg13g2_tielo tt_um_pwm_block_11 (.L_LO(net11));
 sg13g2_tielo tt_um_pwm_block_12 (.L_LO(net12));
 sg13g2_tielo tt_um_pwm_block_13 (.L_LO(net13));
 sg13g2_tielo tt_um_pwm_block_14 (.L_LO(net14));
 sg13g2_tiehi _5031__15 (.L_HI(net15));
 sg13g2_buf_1 _5400_ (.A(\MemCell.enable_pwm ),
    .X(uio_out[0]));
 sg13g2_ebufn_4 _5401_ (.A(reg_ui0),
    .TE_B(_2397_),
    .Z(uio_out[3]));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(net649));
 sg13g2_buf_4 fanout649 (.X(net649),
    .A(_2214_));
 sg13g2_buf_2 fanout650 (.A(net652),
    .X(net650));
 sg13g2_buf_4 fanout651 (.X(net651),
    .A(net652));
 sg13g2_buf_2 fanout652 (.A(_2013_),
    .X(net652));
 sg13g2_buf_4 fanout653 (.X(net653),
    .A(net654));
 sg13g2_buf_2 fanout654 (.A(_1737_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_1737_),
    .X(net655));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(net657));
 sg13g2_buf_4 fanout657 (.X(net657),
    .A(_2213_));
 sg13g2_buf_2 fanout658 (.A(net659),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(net662),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_4 fanout661 (.X(net661),
    .A(net662));
 sg13g2_buf_2 fanout662 (.A(_1497_),
    .X(net662));
 sg13g2_buf_4 fanout663 (.X(net663),
    .A(net664));
 sg13g2_buf_2 fanout664 (.A(_1497_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(net667),
    .X(net665));
 sg13g2_buf_1 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_4 fanout668 (.X(net668),
    .A(net669));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(_1496_));
 sg13g2_buf_2 fanout670 (.A(net673),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(net673),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_0656_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(net679),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(net679),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(net677),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(net679),
    .X(net678));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(_0656_));
 sg13g2_buf_2 fanout680 (.A(net684),
    .X(net680));
 sg13g2_buf_1 fanout681 (.A(net684),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(net684),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(net684),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(net691),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(net686),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(net688),
    .X(net687));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(net691));
 sg13g2_buf_4 fanout689 (.X(net689),
    .A(net691));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(net691));
 sg13g2_buf_4 fanout691 (.X(net691),
    .A(_0816_));
 sg13g2_buf_2 fanout692 (.A(net694),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_0655_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_0655_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(net697),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_0650_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_0650_),
    .X(net697));
 sg13g2_buf_4 fanout698 (.X(net698),
    .A(_1900_));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(_1897_));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(_1894_));
 sg13g2_buf_2 fanout701 (.A(_1891_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(_1887_),
    .X(net702));
 sg13g2_buf_4 fanout703 (.X(net703),
    .A(_1884_));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(_1877_));
 sg13g2_buf_4 fanout705 (.X(net705),
    .A(_1874_));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(_1857_));
 sg13g2_buf_2 fanout707 (.A(_1853_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_1849_),
    .X(net708));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(_1841_));
 sg13g2_buf_2 fanout710 (.A(_2112_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_1909_),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(_1880_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_1870_),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(_1867_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_1864_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_1861_),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(_1846_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_0099_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_0510_),
    .X(net719));
 sg13g2_buf_4 fanout720 (.X(net720),
    .A(net723));
 sg13g2_buf_2 fanout721 (.A(net723),
    .X(net721));
 sg13g2_buf_8 fanout722 (.A(net723),
    .X(net722));
 sg13g2_buf_4 fanout723 (.X(net723),
    .A(_2345_));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(net727));
 sg13g2_buf_2 fanout725 (.A(net727),
    .X(net725));
 sg13g2_buf_8 fanout726 (.A(net727),
    .X(net726));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(_2344_));
 sg13g2_buf_2 fanout728 (.A(net557),
    .X(net728));
 sg13g2_buf_4 fanout729 (.X(net729),
    .A(net556));
 sg13g2_buf_8 fanout730 (.A(net733),
    .X(net730));
 sg13g2_buf_4 fanout731 (.X(net731),
    .A(net733));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(net733));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(\MemCell.o_RX_Byte[7] ));
 sg13g2_buf_8 fanout734 (.A(net737),
    .X(net734));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(net737));
 sg13g2_buf_2 fanout736 (.A(net737),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(\MemCell.o_RX_Byte[6] ),
    .X(net737));
 sg13g2_buf_8 fanout738 (.A(net741),
    .X(net738));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(net741));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(net741));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(\MemCell.o_RX_Byte[5] ));
 sg13g2_buf_8 fanout742 (.A(net745),
    .X(net742));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(net745));
 sg13g2_buf_2 fanout744 (.A(net745),
    .X(net744));
 sg13g2_buf_4 fanout745 (.X(net745),
    .A(\MemCell.o_RX_Byte[4] ));
 sg13g2_buf_4 fanout746 (.X(net746),
    .A(net749));
 sg13g2_buf_2 fanout747 (.A(net749),
    .X(net747));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(net749));
 sg13g2_buf_4 fanout749 (.X(net749),
    .A(\MemCell.o_RX_Byte[3] ));
 sg13g2_buf_8 fanout750 (.A(net753),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(net753),
    .X(net751));
 sg13g2_buf_8 fanout752 (.A(net753),
    .X(net752));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(net507));
 sg13g2_buf_2 fanout754 (.A(net79),
    .X(net754));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(_2370_));
 sg13g2_buf_2 fanout756 (.A(_2370_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(net760),
    .X(net757));
 sg13g2_buf_1 fanout758 (.A(net760),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(net760),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_2356_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_2347_),
    .X(net761));
 sg13g2_buf_1 fanout762 (.A(_2347_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(net764),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(uio_in[7]),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(net767),
    .X(net765));
 sg13g2_buf_1 fanout766 (.A(net767),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(uio_in[4]),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(ui_in[6]),
    .X(net768));
 sg13g2_buf_1 fanout769 (.A(ui_in[6]),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(net771),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(ui_in[6]),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(net773),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(net774),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(ui_in[5]),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(net777),
    .X(net775));
 sg13g2_buf_1 fanout776 (.A(net777),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(net3),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(net780),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(net787),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(net782),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(net787),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(net784),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(net787),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(net787),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(ui_in[3]));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(net789));
 sg13g2_buf_2 fanout789 (.A(net793),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(net791));
 sg13g2_buf_1 fanout791 (.A(net793),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(net793),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(ui_in[2]),
    .X(net793));
 sg13g2_buf_4 fanout794 (.X(net794),
    .A(ui_in[2]));
 sg13g2_buf_2 fanout795 (.A(ui_in[2]),
    .X(net795));
 sg13g2_buf_4 fanout796 (.X(net796),
    .A(net803));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(net803));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(net799));
 sg13g2_buf_4 fanout799 (.X(net799),
    .A(net803));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(net802));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(net802));
 sg13g2_buf_2 fanout802 (.A(net803),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(net864),
    .X(net803));
 sg13g2_buf_4 fanout804 (.X(net804),
    .A(net806));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(net806));
 sg13g2_buf_2 fanout806 (.A(net810),
    .X(net806));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(net808));
 sg13g2_buf_4 fanout808 (.X(net808),
    .A(net809));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(net810));
 sg13g2_buf_2 fanout810 (.A(net864),
    .X(net810));
 sg13g2_buf_4 fanout811 (.X(net811),
    .A(net812));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(net815));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(net815));
 sg13g2_buf_2 fanout814 (.A(net815),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(net829),
    .X(net815));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(net819));
 sg13g2_buf_4 fanout817 (.X(net817),
    .A(net819));
 sg13g2_buf_4 fanout818 (.X(net818),
    .A(net819));
 sg13g2_buf_2 fanout819 (.A(net829),
    .X(net819));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(net824));
 sg13g2_buf_2 fanout821 (.A(net824),
    .X(net821));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(net824));
 sg13g2_buf_4 fanout823 (.X(net823),
    .A(net824));
 sg13g2_buf_2 fanout824 (.A(net829),
    .X(net824));
 sg13g2_buf_4 fanout825 (.X(net825),
    .A(net828));
 sg13g2_buf_2 fanout826 (.A(net828),
    .X(net826));
 sg13g2_buf_4 fanout827 (.X(net827),
    .A(net828));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(net829));
 sg13g2_buf_2 fanout829 (.A(net864),
    .X(net829));
 sg13g2_buf_4 fanout830 (.X(net830),
    .A(net833));
 sg13g2_buf_4 fanout831 (.X(net831),
    .A(net833));
 sg13g2_buf_4 fanout832 (.X(net832),
    .A(net833));
 sg13g2_buf_2 fanout833 (.A(net844),
    .X(net833));
 sg13g2_buf_4 fanout834 (.X(net834),
    .A(net844));
 sg13g2_buf_4 fanout835 (.X(net835),
    .A(net844));
 sg13g2_buf_4 fanout836 (.X(net836),
    .A(net837));
 sg13g2_buf_4 fanout837 (.X(net837),
    .A(net843));
 sg13g2_buf_4 fanout838 (.X(net838),
    .A(net842));
 sg13g2_buf_2 fanout839 (.A(net842),
    .X(net839));
 sg13g2_buf_4 fanout840 (.X(net840),
    .A(net842));
 sg13g2_buf_2 fanout841 (.A(net842),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(net843),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(net844),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(net864),
    .X(net844));
 sg13g2_buf_4 fanout845 (.X(net845),
    .A(net848));
 sg13g2_buf_2 fanout846 (.A(net848),
    .X(net846));
 sg13g2_buf_4 fanout847 (.X(net847),
    .A(net848));
 sg13g2_buf_2 fanout848 (.A(net863),
    .X(net848));
 sg13g2_buf_4 fanout849 (.X(net849),
    .A(net853));
 sg13g2_buf_2 fanout850 (.A(net853),
    .X(net850));
 sg13g2_buf_4 fanout851 (.X(net851),
    .A(net853));
 sg13g2_buf_2 fanout852 (.A(net853),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(net863),
    .X(net853));
 sg13g2_buf_4 fanout854 (.X(net854),
    .A(net858));
 sg13g2_buf_2 fanout855 (.A(net858),
    .X(net855));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(net858));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(net858));
 sg13g2_buf_2 fanout858 (.A(net863),
    .X(net858));
 sg13g2_buf_4 fanout859 (.X(net859),
    .A(net862));
 sg13g2_buf_4 fanout860 (.X(net860),
    .A(net862));
 sg13g2_buf_4 fanout861 (.X(net861),
    .A(net863));
 sg13g2_buf_2 fanout862 (.A(net863),
    .X(net862));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(net864));
 sg13g2_buf_4 fanout864 (.X(net864),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[4]));
 sg13g2_buf_2 input4 (.A(ui_in[7]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[6]),
    .X(net5));
 sg13g2_tielo tt_um_pwm_block_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_44_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_43_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_35_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_31_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_7_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_17_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_13_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_21_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\spi_module.r2_RX_Done ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0191_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0067_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold4 (.A(\pwm_module.counter1[31] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0505_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0193_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0070_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0194_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0072_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold10 (.A(\pwm_module.counter0[31] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0254_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold12 (.A(\pwm_module.counter2[15] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0449_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold14 (.A(\pwm_module.counter2[31] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0465_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold16 (.A(\pwm_module.counter0[23] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0246_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold18 (.A(\pwm_module.counter0[19] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0242_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0198_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0079_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0201_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0085_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold24 (.A(\pwm_module.counter1[23] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0497_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold26 (.A(\pwm_module.counter0[3] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0226_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold28 (.A(\pwm_module.counter2[23] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0457_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold30 (.A(\pwm_module.counter2[19] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0453_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold32 (.A(\pwm_module.counter2[27] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0461_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold34 (.A(\pwm_module.counter1[19] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0493_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold36 (.A(\pwm_module.counter0[15] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0238_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold38 (.A(\pwm_module.counter0[27] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0250_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold40 (.A(\MemCell.prescale_reg[2][2] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold41 (.A(\pwm_module.counter2[3] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0437_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold43 (.A(\pwm_module.counter2[11] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0445_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold45 (.A(\pwm_module.counter0[0] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold46 (.A(\pwm_module.prescaler1[29] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0703_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0055_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold49 (.A(\pwm_module.counter1[27] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0501_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold51 (.A(\pwm_module.counter2[29] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0463_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold53 (.A(\pwm_module.counter1[11] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0485_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold55 (.A(\pwm_module.counter2[17] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0451_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold57 (.A(\pwm_module.counter2[25] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0459_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold59 (.A(\pwm_module.counter2[12] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0446_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold61 (.A(\pwm_module.counter1[17] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0491_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold63 (.A(\pwm_module.counter0[11] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0234_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold65 (.A(\MemCell.dc3_reg[1][1] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0184_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0053_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold68 (.A(\pwm_module.counter0[4] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold69 (.A(\MemCell.prescale_reg[1][2] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold70 (.A(\MemCell.dc3_reg[2][1] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold71 (.A(\MemCell.dc1_reg[3][1] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold72 (.A(\pwm_module.counter1[15] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0489_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold74 (.A(\MemCell.prescale_reg[0][1] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold75 (.A(\pwm_module.counter1[9] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0483_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0171_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold78 (.A(_1572_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold79 (.A(\MemCell.dc3_reg[3][5] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold80 (.A(\MemCell.dc1_reg[1][2] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold81 (.A(\MemCell.dc1_reg[2][3] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold82 (.A(\MemCell.dc3_reg[2][4] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0291_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold84 (.A(\MemCell.counter_value[19] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold85 (.A(\MemCell.dc2_reg[1][3] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold86 (.A(\pwm_module.counter1[13] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0487_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0178_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0676_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold90 (.A(\MemCell.dc3_reg[3][2] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold91 (.A(\MemCell.counter_value[4] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold92 (.A(\MemCell.dc1_reg[3][3] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold93 (.A(\pwm_module.counter2[13] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0447_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0208_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold96 (.A(_1522_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold97 (.A(\MemCell.dc2_reg[3][5] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold98 (.A(\MemCell.counter_value[31] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold99 (.A(\MemCell.dc3_reg[2][0] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold100 (.A(\MemCell.dc1_reg[0][2] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold101 (.A(\MemCell.dc3_reg[1][5] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold102 (.A(\MemCell.dc3_reg[2][7] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold103 (.A(\MemCell.dc3_reg[2][5] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold104 (.A(\MemCell.counter_value[12] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold105 (.A(\MemCell.dc1_reg[0][0] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold106 (.A(\MemCell.dc3_reg[3][6] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold107 (.A(\MemCell.dc1_reg[1][0] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0176_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold109 (.A(_1584_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold110 (.A(\MemCell.dc3_reg[1][4] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold111 (.A(\MemCell.dc1_reg[1][4] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold112 (.A(\MemCell.dc2_reg[3][4] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold113 (.A(\pwm_module.counter2[9] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0443_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold115 (.A(\MemCell.dc2_reg[0][1] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold116 (.A(\MemCell.dc3_reg[1][2] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold117 (.A(\MemCell.dc1_reg[2][0] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold118 (.A(\pwm_module.counter1[3] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0477_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold120 (.A(\MemCell.dc2_reg[3][7] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold121 (.A(\MemCell.dc2_reg[2][2] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold122 (.A(\MemCell.counter_value[28] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold123 (.A(\MemCell.dc1_reg[2][2] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold124 (.A(\MemCell.dc2_reg[3][2] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold125 (.A(\pwm_module.counter1[29] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0503_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold127 (.A(\MemCell.dc1_reg[3][5] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold128 (.A(\pwm_module.counter1[25] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0499_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold130 (.A(\MemCell.dc3_reg[2][6] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold131 (.A(\MemCell.counter_value[3] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold132 (.A(\MemCell.dc3_reg[1][7] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold133 (.A(\MemCell.dc3_reg[3][1] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold134 (.A(\MemCell.dc3_reg[3][4] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold135 (.A(\MemCell.dc1_reg[0][5] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold136 (.A(\MemCell.dc2_reg[1][7] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold137 (.A(\MemCell.dc2_reg[2][5] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold138 (.A(\MemCell.counter_value[8] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold139 (.A(\MemCell.dc3_reg[3][0] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold140 (.A(\MemCell.dc2_reg[2][4] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold141 (.A(\MemCell.dc2_reg[3][6] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold142 (.A(\MemCell.counter_value[18] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold143 (.A(\MemCell.dc2_reg[1][6] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold144 (.A(\MemCell.counter_value[16] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0172_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold146 (.A(_1575_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold147 (.A(\MemCell.counter_value[0] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0415_),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold149 (.A(\MemCell.prescale_reg[0][2] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold150 (.A(\pwm_module.counter2[30] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0464_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold152 (.A(\MemCell.dc1_reg[1][5] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0213_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold154 (.A(_1541_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold155 (.A(\MemCell.dc3_reg[2][3] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0175_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold157 (.A(_1581_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0181_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0686_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold160 (.A(\pwm_module.counter1[12] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0486_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold162 (.A(\MemCell.dc2_reg[2][0] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold163 (.A(\MemCell.dc3_reg[1][6] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0155_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0235_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold166 (.A(\MemCell.dc1_reg[3][0] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold167 (.A(\MemCell.counter_value[2] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0417_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold169 (.A(\MemCell.dc2_reg[1][4] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0210_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold171 (.A(_1532_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold172 (.A(\MemCell.dc3_reg[3][3] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold173 (.A(\MemCell.dc2_reg[0][2] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold174 (.A(\MemCell.counter_value[29] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold175 (.A(\pwm_module.counter2[21] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0455_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold177 (.A(\MemCell.dc3_reg[2][2] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold178 (.A(\pwm_module.counter1[21] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0495_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold180 (.A(\MemCell.dc1_reg[3][4] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold181 (.A(\MemCell.dc2_reg[3][0] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold182 (.A(\pwm_module.counter2[7] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0441_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold184 (.A(\MemCell.dc3_reg[0][0] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0426_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold186 (.A(\MemCell.dc1_reg[1][6] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold187 (.A(\MemCell.dc1_reg[3][6] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold188 (.A(\pwm_module.prescaler0[2] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold189 (.A(_1500_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold190 (.A(\MemCell.prescale_reg[3][2] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold191 (.A(\MemCell.dc1_reg[2][4] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold192 (.A(\pwm_module.prescaler1[2] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold193 (.A(_1565_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold194 (.A(\MemCell.dc2_reg[1][2] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold195 (.A(\pwm_module.counter1[20] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold196 (.A(_2284_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0496_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold198 (.A(\MemCell.dc1_reg[2][6] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold199 (.A(\pwm_module.counter1[7] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0481_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold201 (.A(\MemCell.counter_value[9] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0150_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0243_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold204 (.A(\pwm_module.prescaler0[0] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold205 (.A(\MemCell.dc1_reg[0][3] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold206 (.A(\MemCell.counter_value[10] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold207 (.A(\MemCell.dc1_reg[0][6] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold208 (.A(\pwm_module.prescaler2[6] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0827_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0200_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0083_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold212 (.A(\MemCell.counter_value[7] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold213 (.A(\pwm_module.counter0[17] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0240_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold215 (.A(\MemCell.counter_value[27] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0203_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold217 (.A(_1501_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold218 (.A(\pwm_module.counter0[5] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0228_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold220 (.A(\pwm_module.counter1[6] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0480_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold222 (.A(\MemCell.dc1_reg[3][2] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0205_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold224 (.A(_1508_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold225 (.A(\MemCell.dc1_reg[0][7] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold226 (.A(\pwm_module.counter2[6] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0440_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold228 (.A(\MemCell.dc2_reg[1][5] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0209_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold230 (.A(\MemCell.counter_value[13] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold231 (.A(\pwm_module.counter0[7] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0230_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0173_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold234 (.A(_1578_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold235 (.A(\MemCell.counter_value[14] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0204_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold237 (.A(_1504_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold238 (.A(\MemCell.counter_value[21] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold239 (.A(\MemCell.prescale_reg[3][7] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold240 (.A(\pwm_module.prescaler0[5] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold241 (.A(_1506_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0028_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold243 (.A(\MemCell.dc3_reg[0][6] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold244 (.A(\MemCell.dc1_reg[2][7] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0334_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold246 (.A(\MemCell.dc3_reg[0][3] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold247 (.A(\MemCell.prescale_reg[3][6] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold248 (.A(\MemCell.counter_value[24] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold249 (.A(\pwm_module.prescaler2[0] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold250 (.A(\MemCell.dc3_reg[1][3] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold251 (.A(\MemCell.dc1_reg[1][7] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold252 (.A(\MemCell.counter_value[22] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold253 (.A(\MemCell.dc2_reg[1][0] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold254 (.A(\MemCell.dc3_reg[0][2] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0428_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold256 (.A(\pwm_module.counter0[6] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0229_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0215_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold259 (.A(_1550_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold260 (.A(\MemCell.dc2_reg[2][3] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold261 (.A(\MemCell.dc3_reg[0][5] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold262 (.A(\MemCell.counter_value[1] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0416_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold264 (.A(\MemCell.counter_value[30] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold265 (.A(\MemCell.dc1_reg[1][3] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold266 (.A(\pwm_module.counter2[10] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0444_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold268 (.A(\MemCell.prescale_reg[3][5] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold269 (.A(\pwm_module.counter2[20] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0454_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0214_),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold272 (.A(_1546_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold273 (.A(\MemCell.dc1_reg[2][1] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold274 (.A(\pwm_module.counter1[30] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0504_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold276 (.A(\MemCell.prescale_reg[3][1] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold277 (.A(\MemCell.dc2_reg[2][7] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0206_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold279 (.A(_1513_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold280 (.A(\MemCell.prescale_reg[2][0] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold281 (.A(\MemCell.dc3_reg[0][1] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0427_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold283 (.A(\pwm_module.prescaler0[4] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold284 (.A(_1503_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0026_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold286 (.A(\MemCell.prescale_reg[2][7] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold287 (.A(\MemCell.prescale_reg[2][1] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold288 (.A(\MemCell.dc2_reg[2][1] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold289 (.A(\MemCell.prescale_reg[0][4] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0211_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold291 (.A(_1536_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold292 (.A(\pwm_module.counter0[29] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0252_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold294 (.A(\pwm_module.prescaler0[17] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold295 (.A(_1533_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold296 (.A(\MemCell.dc2_reg[0][6] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold297 (.A(\MemCell.counter_value[6] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold298 (.A(\MemCell.dc2_reg[1][1] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold299 (.A(_0207_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0108_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold301 (.A(\MemCell.prescale_reg[1][0] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold302 (.A(\MemCell.dc3_reg[3][7] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold303 (.A(\MemCell.dc3_reg[1][0] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0174_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold305 (.A(_1580_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold306 (.A(\MemCell.prescale_reg[2][4] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold307 (.A(\pwm_module.counter2[5] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0439_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold309 (.A(\MemCell.counter_value[25] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold310 (.A(\MemCell.dc3_reg[0][4] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold311 (.A(\MemCell.dc3_reg[0][7] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold312 (.A(\MemCell.dc1_reg[2][5] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0332_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold314 (.A(\MemCell.prescale_reg[1][7] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0382_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold316 (.A(\MemCell.dc1_reg[0][1] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold317 (.A(\MemCell.counter_value[26] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold318 (.A(\MemCell.counter_value[23] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0212_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold320 (.A(_1539_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold321 (.A(\MemCell.dc2_reg[0][3] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0314_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold323 (.A(\pwm_module.prescaler1[0] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold324 (.A(\MemCell.dc1_reg[0][4] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold325 (.A(\pwm_module.counter1[10] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold326 (.A(_0484_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold327 (.A(\MemCell.dc2_reg[3][3] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold328 (.A(\MemCell.dc2_reg[0][0] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold329 (.A(\MemCell.dc2_reg[2][6] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold330 (.A(\MemCell.dc2_reg[0][5] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold331 (.A(\MemCell.prescale_reg[3][3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold332 (.A(\MemCell.prescale_reg[1][1] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold333 (.A(\pwm_module.counter0[9] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0232_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold335 (.A(\MemCell.counter_value[20] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold336 (.A(\MemCell.dc1_reg[1][1] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold337 (.A(\MemCell.prescale_reg[2][5] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold338 (.A(\MemCell.dc2_reg[3][1] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold339 (.A(\MemCell.prescale_reg[0][5] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold340 (.A(\MemCell.dc2_reg[0][7] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold341 (.A(\spi_module.r3_RX_Done ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold342 (.A(\pwm_module.prescaler0[16] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold343 (.A(_1531_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0007_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0177_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold346 (.A(_1586_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold347 (.A(\pwm_module.prescaler0[30] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold348 (.A(_1561_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold349 (.A(\MemCell.prescale_reg[3][4] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold350 (.A(_0197_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0865_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold352 (.A(\MemCell.prescale_reg[0][7] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold353 (.A(\MemCell.prescale_reg[3][0] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0183_),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0696_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold356 (.A(\pwm_module.counter1[26] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0180_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0681_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0185_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0707_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold361 (.A(\MemCell.prescale_reg[1][6] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0381_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold363 (.A(\MemCell.counter_value[5] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold364 (.A(\MemCell.dc1_reg[3][7] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold365 (.A(\MemCell.counter_value[11] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold366 (.A(\pwm_module.counter0[25] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0248_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0187_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold369 (.A(\MemCell.prescale_reg[0][6] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0188_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold371 (.A(\pwm_module.prescaler0[14] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0005_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0179_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0679_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold375 (.A(\MemCell.counter_value[17] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold376 (.A(\pwm_module.prescaler2[24] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold377 (.A(_0080_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold378 (.A(\pwm_module.prescaler2[4] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0823_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold380 (.A(\pwm_module.counter1[14] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold381 (.A(\MemCell.o_RX_Byte[1] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0218_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold383 (.A(\pwm_module.prescaler0[28] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold384 (.A(_1557_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold385 (.A(\MemCell.dc2_reg[0][4] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold386 (.A(\MemCell.curr_state[2] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0901_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0423_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0169_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold390 (.A(_1566_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold391 (.A(\pwm_module.counter0[21] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0244_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0186_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0821_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold395 (.A(\MemCell.prescale_reg[0][0] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold396 (.A(\pwm_module.prescaler0[1] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0189_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0835_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold399 (.A(\MemCell.prescale_reg[1][5] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold400 (.A(\pwm_module.counter0[13] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0236_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold402 (.A(\MemCell.prescale_reg[2][6] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold403 (.A(\MemCell.prescale_reg[1][4] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0379_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold405 (.A(\pwm_module.prescaler1[10] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold406 (.A(_1577_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold407 (.A(\pwm_module.counter1[4] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold408 (.A(\pwm_module.prescaler1[28] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0699_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0052_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold411 (.A(\pwm_module.counter1[24] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold412 (.A(_2291_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0170_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold414 (.A(_1569_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold415 (.A(\pwm_module.prescaler1[6] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold416 (.A(_1571_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold417 (.A(\pwm_module.prescaler1[22] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0685_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold419 (.A(\pwm_module.prescaler1[24] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0690_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold421 (.A(\pwm_module.counter0[10] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold422 (.A(_0233_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold423 (.A(\pwm_module.prescaler1[14] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold424 (.A(_1583_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold425 (.A(\pwm_module.prescaler0[9] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold426 (.A(_1514_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0001_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold428 (.A(\MemCell.prescale_reg[2][3] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold429 (.A(\MemCell.prescale_reg[0][3] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0182_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold431 (.A(\pwm_module.prescaler1[18] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0675_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold433 (.A(\pwm_module.counter1[16] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold434 (.A(_2267_),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold435 (.A(\pwm_module.prescaler1[16] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold436 (.A(\pwm_module.counter2[4] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold437 (.A(\MemCell.prescale_reg[1][3] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold438 (.A(\pwm_module.prescaler1[8] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold439 (.A(_1574_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold440 (.A(_0192_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0845_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold442 (.A(\pwm_module.prescaler1[1] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold443 (.A(\pwm_module.counter1[5] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0479_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold445 (.A(\pwm_module.counter0[18] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold446 (.A(_1792_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold447 (.A(\pwm_module.counter2[22] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0456_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold449 (.A(\pwm_module.counter0[30] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0253_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold451 (.A(\pwm_module.counter0[1] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0216_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold453 (.A(_1553_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0018_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold455 (.A(\pwm_module.prescaler0[12] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold456 (.A(_1521_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold457 (.A(\pwm_module.counter1[18] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0190_),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold459 (.A(_0840_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold460 (.A(\pwm_module.counter0[8] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold461 (.A(\pwm_module.counter2[1] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold462 (.A(_2017_),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0196_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0864_),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold465 (.A(\pwm_module.counter2[28] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold466 (.A(_2103_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold467 (.A(\pwm_module.prescaler1[4] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold468 (.A(_1568_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold469 (.A(_0123_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold470 (.A(_0888_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold471 (.A(\pwm_module.counter2[0] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold472 (.A(\pwm_module.counter1[28] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold473 (.A(\MemCell.o_RX_Byte[0] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold474 (.A(\pwm_module.prescaler2[21] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0866_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0868_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold477 (.A(_0078_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0199_),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0195_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0860_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold481 (.A(\pwm_module.prescaler2[29] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0885_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0886_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0087_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold485 (.A(\pwm_module.counter2[18] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold486 (.A(\pwm_module.counter2[14] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold487 (.A(_2057_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold488 (.A(\pwm_module.counter2[26] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold489 (.A(\pwm_module.prescaler0[8] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold490 (.A(_1512_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold491 (.A(\pwm_module.counter0[16] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold492 (.A(_0217_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold493 (.A(\pwm_module.counter0[2] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold494 (.A(\pwm_module.counter2[16] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold495 (.A(\pwm_module.prescaler1[26] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold496 (.A(_0695_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold497 (.A(\pwm_module.counter2[8] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0102_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold499 (.A(\pwm_module.counter1[2] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold500 (.A(\pwm_module.counter0[20] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold501 (.A(_1805_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold502 (.A(_0245_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold503 (.A(\pwm_module.counter0[28] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold504 (.A(_1824_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold505 (.A(\MemCell.counter_value[15] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold506 (.A(\pwm_module.prescaler2[15] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold507 (.A(_0853_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold508 (.A(_0854_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold509 (.A(\pwm_module.prescaler2[9] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold510 (.A(_0838_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold511 (.A(_0065_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold512 (.A(\pwm_module.counter2[24] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold513 (.A(\pwm_module.prescaler2[2] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold514 (.A(_0819_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold515 (.A(\pwm_module.counter1[8] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0482_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold517 (.A(\pwm_module.counter1[1] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold518 (.A(\pwm_module.counter0[26] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold519 (.A(_0249_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold520 (.A(\pwm_module.counter0[14] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold521 (.A(_0237_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold522 (.A(\MemCell.counter[0] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold523 (.A(\pwm_module.counter1[0] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold524 (.A(_0144_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold525 (.A(\MemCell.o_RX_Byte[2] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold526 (.A(\MemCell.next_state[0] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold527 (.A(\pwm_module.prescaler2[1] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold528 (.A(\pwm_module.prescaler0[24] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold529 (.A(_1548_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold530 (.A(\pwm_module.counter0[24] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold531 (.A(\pwm_module.prescaler0[22] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold532 (.A(_1544_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold533 (.A(\pwm_module.prescaler2[14] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold534 (.A(_0849_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold535 (.A(\pwm_module.prescaler2[8] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold536 (.A(\pwm_module.prescaler2[18] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0858_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold538 (.A(\pwm_module.prescaler2[26] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold539 (.A(\pwm_module.counter2[2] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold540 (.A(_2018_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold541 (.A(\pwm_module.prescaler2[28] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold542 (.A(_0883_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold543 (.A(\MemCell.counter[1] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold544 (.A(\pwm_module.prescaler2[14] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold545 (.A(\pwm_module.prescaler1[0] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold546 (.A(\pwm_module.counter2[24] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold547 (.A(\pwm_module.prescaler0[0] ),
    .X(net581));
 sg13g2_antennanp ANTENNA_1 (.A(_0096_));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(_0096_));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(_0096_));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_fill_2 FILLER_0_42 ();
 sg13g2_fill_2 FILLER_0_53 ();
 sg13g2_fill_2 FILLER_0_72 ();
 sg13g2_fill_1 FILLER_0_74 ();
 sg13g2_fill_1 FILLER_0_89 ();
 sg13g2_decap_4 FILLER_0_155 ();
 sg13g2_fill_2 FILLER_0_159 ();
 sg13g2_decap_4 FILLER_0_175 ();
 sg13g2_decap_4 FILLER_0_189 ();
 sg13g2_fill_1 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_0_229 ();
 sg13g2_decap_4 FILLER_0_236 ();
 sg13g2_fill_2 FILLER_0_240 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_fill_1 FILLER_0_262 ();
 sg13g2_fill_2 FILLER_0_271 ();
 sg13g2_fill_1 FILLER_0_273 ();
 sg13g2_fill_2 FILLER_0_286 ();
 sg13g2_fill_1 FILLER_0_288 ();
 sg13g2_fill_2 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_fill_2 FILLER_1_14 ();
 sg13g2_fill_2 FILLER_1_68 ();
 sg13g2_fill_1 FILLER_1_70 ();
 sg13g2_fill_2 FILLER_1_97 ();
 sg13g2_fill_2 FILLER_1_135 ();
 sg13g2_fill_1 FILLER_1_137 ();
 sg13g2_fill_2 FILLER_1_164 ();
 sg13g2_fill_1 FILLER_1_166 ();
 sg13g2_fill_2 FILLER_1_177 ();
 sg13g2_fill_1 FILLER_1_179 ();
 sg13g2_decap_4 FILLER_1_206 ();
 sg13g2_fill_1 FILLER_1_288 ();
 sg13g2_fill_2 FILLER_1_298 ();
 sg13g2_fill_1 FILLER_1_309 ();
 sg13g2_fill_2 FILLER_1_319 ();
 sg13g2_fill_1 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_4 FILLER_2_28 ();
 sg13g2_fill_2 FILLER_2_110 ();
 sg13g2_fill_1 FILLER_2_169 ();
 sg13g2_fill_2 FILLER_2_206 ();
 sg13g2_fill_1 FILLER_2_208 ();
 sg13g2_fill_1 FILLER_2_219 ();
 sg13g2_fill_2 FILLER_2_244 ();
 sg13g2_fill_1 FILLER_2_324 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_4 FILLER_3_14 ();
 sg13g2_fill_2 FILLER_3_18 ();
 sg13g2_fill_1 FILLER_3_65 ();
 sg13g2_fill_1 FILLER_3_97 ();
 sg13g2_decap_4 FILLER_3_133 ();
 sg13g2_fill_1 FILLER_3_163 ();
 sg13g2_fill_1 FILLER_3_208 ();
 sg13g2_decap_8 FILLER_3_229 ();
 sg13g2_fill_1 FILLER_3_236 ();
 sg13g2_fill_2 FILLER_3_242 ();
 sg13g2_fill_1 FILLER_3_254 ();
 sg13g2_fill_2 FILLER_3_303 ();
 sg13g2_fill_2 FILLER_3_351 ();
 sg13g2_fill_1 FILLER_3_375 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_fill_2 FILLER_4_14 ();
 sg13g2_fill_1 FILLER_4_16 ();
 sg13g2_fill_2 FILLER_4_44 ();
 sg13g2_fill_1 FILLER_4_68 ();
 sg13g2_fill_2 FILLER_4_103 ();
 sg13g2_fill_2 FILLER_4_137 ();
 sg13g2_fill_2 FILLER_4_170 ();
 sg13g2_fill_1 FILLER_4_202 ();
 sg13g2_fill_1 FILLER_4_261 ();
 sg13g2_fill_2 FILLER_4_295 ();
 sg13g2_fill_1 FILLER_4_297 ();
 sg13g2_fill_1 FILLER_4_353 ();
 sg13g2_fill_2 FILLER_4_380 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_2 ();
 sg13g2_fill_2 FILLER_5_29 ();
 sg13g2_fill_2 FILLER_5_59 ();
 sg13g2_fill_2 FILLER_5_73 ();
 sg13g2_fill_2 FILLER_5_136 ();
 sg13g2_fill_2 FILLER_5_144 ();
 sg13g2_fill_1 FILLER_5_146 ();
 sg13g2_fill_1 FILLER_5_170 ();
 sg13g2_decap_4 FILLER_5_234 ();
 sg13g2_fill_1 FILLER_5_238 ();
 sg13g2_fill_2 FILLER_5_360 ();
 sg13g2_fill_1 FILLER_5_362 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_2 ();
 sg13g2_fill_1 FILLER_6_61 ();
 sg13g2_fill_2 FILLER_6_88 ();
 sg13g2_fill_2 FILLER_6_106 ();
 sg13g2_fill_1 FILLER_6_108 ();
 sg13g2_fill_2 FILLER_6_154 ();
 sg13g2_fill_2 FILLER_6_175 ();
 sg13g2_fill_2 FILLER_6_186 ();
 sg13g2_fill_2 FILLER_6_199 ();
 sg13g2_fill_2 FILLER_6_236 ();
 sg13g2_fill_2 FILLER_6_257 ();
 sg13g2_fill_1 FILLER_6_264 ();
 sg13g2_fill_1 FILLER_6_291 ();
 sg13g2_fill_1 FILLER_6_339 ();
 sg13g2_fill_2 FILLER_6_356 ();
 sg13g2_fill_1 FILLER_6_358 ();
 sg13g2_fill_2 FILLER_6_364 ();
 sg13g2_fill_1 FILLER_6_366 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_4 ();
 sg13g2_fill_2 FILLER_7_68 ();
 sg13g2_fill_1 FILLER_7_70 ();
 sg13g2_fill_1 FILLER_7_84 ();
 sg13g2_fill_2 FILLER_7_89 ();
 sg13g2_fill_2 FILLER_7_95 ();
 sg13g2_fill_1 FILLER_7_97 ();
 sg13g2_fill_2 FILLER_7_121 ();
 sg13g2_fill_2 FILLER_7_189 ();
 sg13g2_fill_2 FILLER_7_214 ();
 sg13g2_fill_1 FILLER_7_216 ();
 sg13g2_fill_1 FILLER_7_243 ();
 sg13g2_fill_2 FILLER_7_248 ();
 sg13g2_fill_2 FILLER_7_290 ();
 sg13g2_fill_1 FILLER_7_292 ();
 sg13g2_fill_2 FILLER_7_354 ();
 sg13g2_fill_1 FILLER_7_356 ();
 sg13g2_fill_2 FILLER_7_366 ();
 sg13g2_fill_1 FILLER_7_368 ();
 sg13g2_fill_2 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_14 ();
 sg13g2_fill_1 FILLER_8_55 ();
 sg13g2_fill_1 FILLER_8_69 ();
 sg13g2_fill_2 FILLER_8_95 ();
 sg13g2_fill_1 FILLER_8_124 ();
 sg13g2_fill_1 FILLER_8_140 ();
 sg13g2_fill_1 FILLER_8_146 ();
 sg13g2_fill_2 FILLER_8_213 ();
 sg13g2_fill_2 FILLER_8_220 ();
 sg13g2_fill_2 FILLER_8_231 ();
 sg13g2_fill_1 FILLER_8_233 ();
 sg13g2_fill_2 FILLER_8_253 ();
 sg13g2_fill_1 FILLER_8_255 ();
 sg13g2_fill_1 FILLER_8_315 ();
 sg13g2_fill_2 FILLER_8_327 ();
 sg13g2_fill_1 FILLER_8_329 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_14 ();
 sg13g2_fill_1 FILLER_9_18 ();
 sg13g2_fill_2 FILLER_9_125 ();
 sg13g2_decap_8 FILLER_9_137 ();
 sg13g2_fill_1 FILLER_9_144 ();
 sg13g2_fill_1 FILLER_9_171 ();
 sg13g2_fill_2 FILLER_9_209 ();
 sg13g2_fill_2 FILLER_9_252 ();
 sg13g2_fill_2 FILLER_9_262 ();
 sg13g2_fill_1 FILLER_9_264 ();
 sg13g2_fill_1 FILLER_9_269 ();
 sg13g2_fill_1 FILLER_9_278 ();
 sg13g2_fill_1 FILLER_9_296 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_fill_1 FILLER_9_338 ();
 sg13g2_fill_1 FILLER_9_361 ();
 sg13g2_fill_2 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_4 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_91 ();
 sg13g2_fill_1 FILLER_10_93 ();
 sg13g2_decap_8 FILLER_10_152 ();
 sg13g2_fill_2 FILLER_10_159 ();
 sg13g2_decap_8 FILLER_10_169 ();
 sg13g2_decap_4 FILLER_10_176 ();
 sg13g2_fill_2 FILLER_10_184 ();
 sg13g2_fill_1 FILLER_10_186 ();
 sg13g2_fill_2 FILLER_10_214 ();
 sg13g2_fill_1 FILLER_10_216 ();
 sg13g2_fill_2 FILLER_10_222 ();
 sg13g2_fill_1 FILLER_10_224 ();
 sg13g2_fill_1 FILLER_10_293 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_4 FILLER_11_14 ();
 sg13g2_fill_1 FILLER_11_27 ();
 sg13g2_fill_1 FILLER_11_84 ();
 sg13g2_fill_2 FILLER_11_102 ();
 sg13g2_fill_1 FILLER_11_104 ();
 sg13g2_fill_2 FILLER_11_168 ();
 sg13g2_fill_1 FILLER_11_170 ();
 sg13g2_fill_2 FILLER_11_220 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_fill_1 FILLER_11_238 ();
 sg13g2_fill_1 FILLER_11_270 ();
 sg13g2_fill_1 FILLER_11_321 ();
 sg13g2_fill_1 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_11 ();
 sg13g2_fill_2 FILLER_12_59 ();
 sg13g2_fill_1 FILLER_12_61 ();
 sg13g2_fill_1 FILLER_12_72 ();
 sg13g2_fill_1 FILLER_12_194 ();
 sg13g2_fill_2 FILLER_12_226 ();
 sg13g2_fill_2 FILLER_12_236 ();
 sg13g2_fill_1 FILLER_12_238 ();
 sg13g2_fill_2 FILLER_12_257 ();
 sg13g2_fill_1 FILLER_12_358 ();
 sg13g2_fill_1 FILLER_12_395 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_fill_1 FILLER_13_44 ();
 sg13g2_fill_2 FILLER_13_60 ();
 sg13g2_fill_2 FILLER_13_70 ();
 sg13g2_fill_1 FILLER_13_72 ();
 sg13g2_fill_2 FILLER_13_87 ();
 sg13g2_fill_1 FILLER_13_89 ();
 sg13g2_fill_1 FILLER_13_138 ();
 sg13g2_fill_1 FILLER_13_200 ();
 sg13g2_fill_1 FILLER_13_330 ();
 sg13g2_fill_1 FILLER_13_341 ();
 sg13g2_fill_1 FILLER_13_386 ();
 sg13g2_fill_2 FILLER_13_396 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_1 FILLER_14_29 ();
 sg13g2_fill_2 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_86 ();
 sg13g2_fill_1 FILLER_14_120 ();
 sg13g2_fill_2 FILLER_14_135 ();
 sg13g2_fill_1 FILLER_14_156 ();
 sg13g2_fill_2 FILLER_14_171 ();
 sg13g2_fill_1 FILLER_14_173 ();
 sg13g2_fill_1 FILLER_14_265 ();
 sg13g2_fill_1 FILLER_14_301 ();
 sg13g2_fill_2 FILLER_14_316 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_fill_2 FILLER_14_366 ();
 sg13g2_fill_1 FILLER_14_381 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_54 ();
 sg13g2_fill_1 FILLER_15_56 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_106 ();
 sg13g2_fill_1 FILLER_15_108 ();
 sg13g2_fill_1 FILLER_15_118 ();
 sg13g2_fill_2 FILLER_15_134 ();
 sg13g2_fill_1 FILLER_15_136 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_fill_2 FILLER_15_215 ();
 sg13g2_fill_2 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_285 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_fill_1 FILLER_15_349 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_97 ();
 sg13g2_fill_2 FILLER_16_109 ();
 sg13g2_fill_1 FILLER_16_111 ();
 sg13g2_fill_2 FILLER_16_127 ();
 sg13g2_fill_2 FILLER_16_169 ();
 sg13g2_fill_2 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_fill_2 FILLER_16_253 ();
 sg13g2_fill_2 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_fill_1 FILLER_16_307 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_fill_1 FILLER_16_371 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_23 ();
 sg13g2_fill_2 FILLER_17_121 ();
 sg13g2_fill_2 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_164 ();
 sg13g2_decap_4 FILLER_17_210 ();
 sg13g2_fill_2 FILLER_17_214 ();
 sg13g2_fill_2 FILLER_17_234 ();
 sg13g2_fill_1 FILLER_17_236 ();
 sg13g2_fill_2 FILLER_17_337 ();
 sg13g2_fill_1 FILLER_17_339 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_114 ();
 sg13g2_fill_1 FILLER_18_130 ();
 sg13g2_fill_2 FILLER_18_153 ();
 sg13g2_fill_1 FILLER_18_164 ();
 sg13g2_decap_8 FILLER_18_190 ();
 sg13g2_decap_4 FILLER_18_197 ();
 sg13g2_fill_1 FILLER_18_205 ();
 sg13g2_decap_4 FILLER_18_212 ();
 sg13g2_fill_1 FILLER_18_216 ();
 sg13g2_decap_4 FILLER_18_291 ();
 sg13g2_fill_1 FILLER_18_295 ();
 sg13g2_fill_2 FILLER_18_371 ();
 sg13g2_fill_1 FILLER_18_373 ();
 sg13g2_fill_2 FILLER_18_390 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_11 ();
 sg13g2_fill_1 FILLER_19_26 ();
 sg13g2_decap_8 FILLER_19_90 ();
 sg13g2_fill_1 FILLER_19_112 ();
 sg13g2_fill_2 FILLER_19_155 ();
 sg13g2_fill_1 FILLER_19_191 ();
 sg13g2_fill_1 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_282 ();
 sg13g2_fill_1 FILLER_19_309 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_fill_2 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_19_384 ();
 sg13g2_fill_2 FILLER_19_398 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_27 ();
 sg13g2_fill_1 FILLER_20_29 ();
 sg13g2_fill_2 FILLER_20_40 ();
 sg13g2_fill_1 FILLER_20_42 ();
 sg13g2_fill_2 FILLER_20_78 ();
 sg13g2_fill_1 FILLER_20_80 ();
 sg13g2_decap_4 FILLER_20_86 ();
 sg13g2_fill_1 FILLER_20_94 ();
 sg13g2_decap_8 FILLER_20_99 ();
 sg13g2_decap_8 FILLER_20_106 ();
 sg13g2_decap_8 FILLER_20_138 ();
 sg13g2_fill_2 FILLER_20_145 ();
 sg13g2_fill_1 FILLER_20_230 ();
 sg13g2_fill_2 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_decap_4 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_273 ();
 sg13g2_fill_1 FILLER_20_279 ();
 sg13g2_decap_4 FILLER_20_295 ();
 sg13g2_fill_1 FILLER_20_299 ();
 sg13g2_fill_1 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_37 ();
 sg13g2_decap_4 FILLER_21_64 ();
 sg13g2_fill_1 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_fill_2 FILLER_21_126 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_decap_4 FILLER_21_136 ();
 sg13g2_decap_4 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_2 FILLER_21_172 ();
 sg13g2_fill_1 FILLER_21_195 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_220 ();
 sg13g2_fill_1 FILLER_21_227 ();
 sg13g2_fill_2 FILLER_21_234 ();
 sg13g2_fill_1 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_357 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_decap_4 FILLER_22_128 ();
 sg13g2_fill_2 FILLER_22_132 ();
 sg13g2_decap_4 FILLER_22_143 ();
 sg13g2_fill_2 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_fill_1 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_188 ();
 sg13g2_decap_8 FILLER_22_195 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_decap_8 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_219 ();
 sg13g2_fill_1 FILLER_22_221 ();
 sg13g2_fill_1 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_398 ();
 sg13g2_decap_4 FILLER_23_55 ();
 sg13g2_fill_2 FILLER_23_68 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_100 ();
 sg13g2_decap_4 FILLER_23_161 ();
 sg13g2_fill_1 FILLER_23_165 ();
 sg13g2_decap_4 FILLER_23_175 ();
 sg13g2_fill_1 FILLER_23_179 ();
 sg13g2_decap_4 FILLER_23_193 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_fill_1 FILLER_23_207 ();
 sg13g2_fill_1 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_346 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_16 ();
 sg13g2_fill_2 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_37 ();
 sg13g2_decap_8 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_4 FILLER_24_74 ();
 sg13g2_fill_1 FILLER_24_78 ();
 sg13g2_fill_2 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_111 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_decap_4 FILLER_24_117 ();
 sg13g2_fill_1 FILLER_24_143 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_fill_1 FILLER_24_254 ();
 sg13g2_fill_2 FILLER_24_264 ();
 sg13g2_fill_1 FILLER_24_266 ();
 sg13g2_fill_1 FILLER_24_302 ();
 sg13g2_fill_2 FILLER_24_335 ();
 sg13g2_fill_1 FILLER_24_359 ();
 sg13g2_fill_1 FILLER_25_26 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_53 ();
 sg13g2_fill_2 FILLER_25_219 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_363 ();
 sg13g2_fill_1 FILLER_25_375 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_2 FILLER_26_45 ();
 sg13g2_fill_1 FILLER_26_47 ();
 sg13g2_fill_1 FILLER_26_72 ();
 sg13g2_fill_1 FILLER_26_99 ();
 sg13g2_fill_2 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_220 ();
 sg13g2_fill_2 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_279 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_363 ();
 sg13g2_fill_2 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_39 ();
 sg13g2_fill_1 FILLER_27_41 ();
 sg13g2_fill_1 FILLER_27_86 ();
 sg13g2_fill_1 FILLER_27_145 ();
 sg13g2_fill_2 FILLER_27_152 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_fill_1 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_294 ();
 sg13g2_fill_2 FILLER_27_318 ();
 sg13g2_fill_1 FILLER_27_336 ();
 sg13g2_fill_2 FILLER_27_375 ();
 sg13g2_fill_2 FILLER_28_51 ();
 sg13g2_fill_2 FILLER_28_76 ();
 sg13g2_fill_2 FILLER_28_97 ();
 sg13g2_fill_2 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_123 ();
 sg13g2_fill_2 FILLER_28_152 ();
 sg13g2_fill_2 FILLER_28_249 ();
 sg13g2_fill_1 FILLER_28_251 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_2 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_fill_1 FILLER_28_355 ();
 sg13g2_fill_2 FILLER_29_46 ();
 sg13g2_fill_1 FILLER_29_53 ();
 sg13g2_fill_2 FILLER_29_83 ();
 sg13g2_fill_1 FILLER_29_85 ();
 sg13g2_fill_1 FILLER_29_124 ();
 sg13g2_decap_8 FILLER_29_138 ();
 sg13g2_decap_8 FILLER_29_145 ();
 sg13g2_decap_4 FILLER_29_156 ();
 sg13g2_fill_1 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_166 ();
 sg13g2_fill_1 FILLER_29_185 ();
 sg13g2_fill_1 FILLER_29_206 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_15 ();
 sg13g2_fill_2 FILLER_30_55 ();
 sg13g2_fill_1 FILLER_30_98 ();
 sg13g2_decap_4 FILLER_30_140 ();
 sg13g2_decap_4 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_173 ();
 sg13g2_fill_2 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_fill_2 FILLER_30_361 ();
 sg13g2_fill_2 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_15 ();
 sg13g2_fill_2 FILLER_31_22 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_134 ();
 sg13g2_fill_2 FILLER_31_171 ();
 sg13g2_decap_4 FILLER_31_187 ();
 sg13g2_fill_2 FILLER_31_191 ();
 sg13g2_fill_2 FILLER_31_202 ();
 sg13g2_fill_2 FILLER_31_229 ();
 sg13g2_fill_1 FILLER_31_231 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_291 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_2 FILLER_32_40 ();
 sg13g2_fill_1 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_111 ();
 sg13g2_fill_2 FILLER_32_131 ();
 sg13g2_fill_1 FILLER_32_177 ();
 sg13g2_decap_4 FILLER_32_239 ();
 sg13g2_fill_1 FILLER_32_257 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_fill_1 FILLER_32_282 ();
 sg13g2_fill_1 FILLER_32_329 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_fill_1 FILLER_32_375 ();
 sg13g2_fill_1 FILLER_32_398 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_fill_1 FILLER_33_47 ();
 sg13g2_fill_2 FILLER_33_74 ();
 sg13g2_fill_2 FILLER_33_90 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_204 ();
 sg13g2_fill_1 FILLER_33_249 ();
 sg13g2_fill_2 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_fill_2 FILLER_33_328 ();
 sg13g2_fill_1 FILLER_33_339 ();
 sg13g2_fill_2 FILLER_33_356 ();
 sg13g2_fill_1 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_34_60 ();
 sg13g2_fill_1 FILLER_34_62 ();
 sg13g2_fill_1 FILLER_34_87 ();
 sg13g2_fill_1 FILLER_34_92 ();
 sg13g2_decap_4 FILLER_34_99 ();
 sg13g2_fill_1 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_207 ();
 sg13g2_fill_1 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_336 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_fill_2 FILLER_35_40 ();
 sg13g2_fill_1 FILLER_35_47 ();
 sg13g2_decap_8 FILLER_35_66 ();
 sg13g2_fill_1 FILLER_35_73 ();
 sg13g2_decap_8 FILLER_35_92 ();
 sg13g2_fill_1 FILLER_35_99 ();
 sg13g2_fill_2 FILLER_35_155 ();
 sg13g2_fill_2 FILLER_35_179 ();
 sg13g2_fill_2 FILLER_35_207 ();
 sg13g2_fill_2 FILLER_35_237 ();
 sg13g2_fill_1 FILLER_35_239 ();
 sg13g2_fill_1 FILLER_35_272 ();
 sg13g2_fill_2 FILLER_35_283 ();
 sg13g2_fill_1 FILLER_35_294 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_358 ();
 sg13g2_fill_1 FILLER_35_360 ();
 sg13g2_fill_2 FILLER_35_366 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_11 ();
 sg13g2_fill_1 FILLER_36_13 ();
 sg13g2_fill_2 FILLER_36_35 ();
 sg13g2_fill_1 FILLER_36_69 ();
 sg13g2_decap_4 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_109 ();
 sg13g2_decap_4 FILLER_36_116 ();
 sg13g2_fill_2 FILLER_36_125 ();
 sg13g2_fill_2 FILLER_36_145 ();
 sg13g2_fill_1 FILLER_36_155 ();
 sg13g2_decap_4 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_193 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_4 FILLER_36_224 ();
 sg13g2_fill_1 FILLER_36_228 ();
 sg13g2_fill_2 FILLER_36_234 ();
 sg13g2_fill_1 FILLER_36_236 ();
 sg13g2_decap_8 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_35 ();
 sg13g2_fill_1 FILLER_37_41 ();
 sg13g2_fill_1 FILLER_37_109 ();
 sg13g2_fill_2 FILLER_37_115 ();
 sg13g2_fill_2 FILLER_37_124 ();
 sg13g2_fill_2 FILLER_37_136 ();
 sg13g2_decap_8 FILLER_37_185 ();
 sg13g2_decap_4 FILLER_37_192 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_211 ();
 sg13g2_fill_1 FILLER_37_218 ();
 sg13g2_decap_8 FILLER_37_237 ();
 sg13g2_decap_4 FILLER_37_244 ();
 sg13g2_decap_8 FILLER_37_253 ();
 sg13g2_fill_2 FILLER_37_318 ();
 sg13g2_fill_1 FILLER_38_91 ();
 sg13g2_fill_2 FILLER_38_123 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_150 ();
 sg13g2_fill_2 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_181 ();
 sg13g2_fill_2 FILLER_38_188 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_fill_2 FILLER_38_342 ();
 sg13g2_fill_1 FILLER_38_344 ();
 sg13g2_fill_2 FILLER_38_383 ();
 sg13g2_fill_1 FILLER_38_385 ();
 sg13g2_fill_2 FILLER_38_394 ();
 sg13g2_fill_1 FILLER_39_45 ();
 sg13g2_fill_2 FILLER_39_61 ();
 sg13g2_fill_2 FILLER_39_68 ();
 sg13g2_fill_2 FILLER_39_119 ();
 sg13g2_fill_1 FILLER_39_136 ();
 sg13g2_fill_1 FILLER_39_149 ();
 sg13g2_fill_1 FILLER_39_155 ();
 sg13g2_fill_2 FILLER_39_188 ();
 sg13g2_decap_8 FILLER_39_221 ();
 sg13g2_fill_2 FILLER_39_289 ();
 sg13g2_fill_1 FILLER_39_291 ();
 sg13g2_fill_2 FILLER_39_318 ();
 sg13g2_fill_1 FILLER_39_351 ();
 sg13g2_fill_2 FILLER_39_380 ();
 sg13g2_fill_1 FILLER_39_382 ();
 sg13g2_fill_2 FILLER_40_26 ();
 sg13g2_fill_1 FILLER_40_57 ();
 sg13g2_decap_4 FILLER_40_62 ();
 sg13g2_fill_2 FILLER_40_66 ();
 sg13g2_decap_8 FILLER_40_72 ();
 sg13g2_fill_1 FILLER_40_79 ();
 sg13g2_fill_1 FILLER_40_93 ();
 sg13g2_fill_1 FILLER_40_107 ();
 sg13g2_fill_1 FILLER_40_134 ();
 sg13g2_fill_1 FILLER_40_176 ();
 sg13g2_fill_1 FILLER_40_235 ();
 sg13g2_fill_1 FILLER_40_246 ();
 sg13g2_fill_2 FILLER_40_257 ();
 sg13g2_fill_1 FILLER_40_259 ();
 sg13g2_fill_1 FILLER_40_275 ();
 sg13g2_decap_4 FILLER_40_289 ();
 sg13g2_fill_2 FILLER_40_293 ();
 sg13g2_fill_2 FILLER_40_393 ();
 sg13g2_decap_4 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_4 ();
 sg13g2_fill_1 FILLER_41_32 ();
 sg13g2_fill_1 FILLER_41_43 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_fill_1 FILLER_41_77 ();
 sg13g2_fill_2 FILLER_41_83 ();
 sg13g2_fill_1 FILLER_41_93 ();
 sg13g2_decap_8 FILLER_41_109 ();
 sg13g2_decap_8 FILLER_41_116 ();
 sg13g2_decap_4 FILLER_41_123 ();
 sg13g2_fill_2 FILLER_41_136 ();
 sg13g2_fill_2 FILLER_41_141 ();
 sg13g2_fill_1 FILLER_41_143 ();
 sg13g2_fill_2 FILLER_41_156 ();
 sg13g2_fill_1 FILLER_41_158 ();
 sg13g2_fill_1 FILLER_41_166 ();
 sg13g2_fill_1 FILLER_41_210 ();
 sg13g2_fill_1 FILLER_41_246 ();
 sg13g2_fill_1 FILLER_41_256 ();
 sg13g2_fill_1 FILLER_41_263 ();
 sg13g2_decap_8 FILLER_41_278 ();
 sg13g2_fill_1 FILLER_41_285 ();
 sg13g2_fill_2 FILLER_41_312 ();
 sg13g2_fill_2 FILLER_41_355 ();
 sg13g2_fill_1 FILLER_41_388 ();
 sg13g2_fill_1 FILLER_41_398 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_4 FILLER_42_14 ();
 sg13g2_fill_2 FILLER_42_18 ();
 sg13g2_decap_4 FILLER_42_29 ();
 sg13g2_fill_2 FILLER_42_33 ();
 sg13g2_fill_2 FILLER_42_117 ();
 sg13g2_fill_1 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_124 ();
 sg13g2_fill_1 FILLER_42_131 ();
 sg13g2_fill_1 FILLER_42_165 ();
 sg13g2_decap_4 FILLER_42_171 ();
 sg13g2_fill_2 FILLER_42_175 ();
 sg13g2_fill_2 FILLER_42_182 ();
 sg13g2_fill_1 FILLER_42_184 ();
 sg13g2_fill_2 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_230 ();
 sg13g2_fill_2 FILLER_42_237 ();
 sg13g2_fill_1 FILLER_42_239 ();
 sg13g2_fill_2 FILLER_42_257 ();
 sg13g2_fill_1 FILLER_42_259 ();
 sg13g2_fill_2 FILLER_42_293 ();
 sg13g2_fill_1 FILLER_42_295 ();
 sg13g2_fill_2 FILLER_42_348 ();
 sg13g2_fill_1 FILLER_42_350 ();
 sg13g2_fill_1 FILLER_42_382 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_4 FILLER_43_21 ();
 sg13g2_fill_2 FILLER_43_25 ();
 sg13g2_fill_1 FILLER_43_148 ();
 sg13g2_fill_2 FILLER_43_259 ();
 sg13g2_fill_2 FILLER_43_302 ();
 sg13g2_fill_1 FILLER_43_312 ();
 sg13g2_fill_1 FILLER_43_365 ();
 sg13g2_fill_2 FILLER_43_375 ();
 sg13g2_fill_2 FILLER_43_386 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_41 ();
 sg13g2_fill_2 FILLER_44_92 ();
 sg13g2_fill_2 FILLER_44_121 ();
 sg13g2_fill_1 FILLER_44_142 ();
 sg13g2_decap_8 FILLER_44_151 ();
 sg13g2_decap_8 FILLER_44_158 ();
 sg13g2_fill_1 FILLER_44_165 ();
 sg13g2_decap_4 FILLER_44_201 ();
 sg13g2_fill_1 FILLER_44_224 ();
 sg13g2_fill_1 FILLER_44_234 ();
 sg13g2_fill_2 FILLER_44_296 ();
 sg13g2_fill_1 FILLER_44_321 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_104 ();
 sg13g2_decap_8 FILLER_45_137 ();
 sg13g2_fill_2 FILLER_45_144 ();
 sg13g2_decap_4 FILLER_45_172 ();
 sg13g2_fill_1 FILLER_45_190 ();
 sg13g2_decap_8 FILLER_45_199 ();
 sg13g2_fill_2 FILLER_45_264 ();
 sg13g2_fill_1 FILLER_45_266 ();
 sg13g2_fill_2 FILLER_45_281 ();
 sg13g2_fill_2 FILLER_45_373 ();
 sg13g2_fill_2 FILLER_46_41 ();
 sg13g2_fill_1 FILLER_46_63 ();
 sg13g2_fill_2 FILLER_46_98 ();
 sg13g2_fill_2 FILLER_46_136 ();
 sg13g2_decap_8 FILLER_46_170 ();
 sg13g2_decap_8 FILLER_46_177 ();
 sg13g2_fill_1 FILLER_46_184 ();
 sg13g2_decap_8 FILLER_46_220 ();
 sg13g2_decap_4 FILLER_46_227 ();
 sg13g2_fill_1 FILLER_46_231 ();
 sg13g2_fill_2 FILLER_46_251 ();
 sg13g2_fill_2 FILLER_46_279 ();
 sg13g2_fill_1 FILLER_46_281 ();
 sg13g2_fill_2 FILLER_46_318 ();
 sg13g2_fill_1 FILLER_46_343 ();
 sg13g2_fill_2 FILLER_46_352 ();
 sg13g2_fill_2 FILLER_47_36 ();
 sg13g2_fill_1 FILLER_47_38 ();
 sg13g2_fill_2 FILLER_47_54 ();
 sg13g2_fill_1 FILLER_47_56 ();
 sg13g2_fill_2 FILLER_47_102 ();
 sg13g2_fill_2 FILLER_47_114 ();
 sg13g2_fill_1 FILLER_47_116 ();
 sg13g2_decap_4 FILLER_47_126 ();
 sg13g2_decap_4 FILLER_47_139 ();
 sg13g2_fill_2 FILLER_47_207 ();
 sg13g2_fill_1 FILLER_47_209 ();
 sg13g2_fill_2 FILLER_47_230 ();
 sg13g2_fill_2 FILLER_47_250 ();
 sg13g2_fill_2 FILLER_47_396 ();
 sg13g2_fill_1 FILLER_47_398 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_fill_2 FILLER_48_26 ();
 sg13g2_fill_2 FILLER_48_97 ();
 sg13g2_fill_1 FILLER_48_115 ();
 sg13g2_fill_1 FILLER_48_127 ();
 sg13g2_fill_2 FILLER_48_134 ();
 sg13g2_fill_1 FILLER_48_152 ();
 sg13g2_fill_2 FILLER_48_174 ();
 sg13g2_fill_1 FILLER_48_176 ();
 sg13g2_fill_2 FILLER_48_205 ();
 sg13g2_fill_1 FILLER_48_207 ();
 sg13g2_fill_2 FILLER_48_234 ();
 sg13g2_decap_8 FILLER_48_250 ();
 sg13g2_fill_1 FILLER_48_266 ();
 sg13g2_fill_2 FILLER_48_332 ();
 sg13g2_fill_2 FILLER_48_348 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_2 ();
 sg13g2_fill_1 FILLER_49_62 ();
 sg13g2_fill_1 FILLER_49_99 ();
 sg13g2_fill_1 FILLER_49_106 ();
 sg13g2_fill_2 FILLER_49_115 ();
 sg13g2_fill_1 FILLER_49_117 ();
 sg13g2_fill_2 FILLER_49_161 ();
 sg13g2_decap_4 FILLER_49_234 ();
 sg13g2_fill_2 FILLER_49_238 ();
 sg13g2_fill_1 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_286 ();
 sg13g2_fill_2 FILLER_49_293 ();
 sg13g2_fill_2 FILLER_49_299 ();
 sg13g2_fill_2 FILLER_49_316 ();
 sg13g2_fill_1 FILLER_49_328 ();
 sg13g2_fill_1 FILLER_49_344 ();
 sg13g2_fill_1 FILLER_49_355 ();
 sg13g2_fill_1 FILLER_49_361 ();
 sg13g2_fill_1 FILLER_49_372 ();
 sg13g2_fill_2 FILLER_50_63 ();
 sg13g2_fill_1 FILLER_50_102 ();
 sg13g2_fill_1 FILLER_50_155 ();
 sg13g2_fill_2 FILLER_50_180 ();
 sg13g2_decap_8 FILLER_50_229 ();
 sg13g2_fill_1 FILLER_50_342 ();
 sg13g2_fill_1 FILLER_50_348 ();
 sg13g2_fill_1 FILLER_50_357 ();
 sg13g2_fill_2 FILLER_51_66 ();
 sg13g2_fill_2 FILLER_51_108 ();
 sg13g2_fill_1 FILLER_51_110 ();
 sg13g2_decap_8 FILLER_51_130 ();
 sg13g2_decap_4 FILLER_51_142 ();
 sg13g2_fill_1 FILLER_51_177 ();
 sg13g2_fill_2 FILLER_51_209 ();
 sg13g2_fill_2 FILLER_51_219 ();
 sg13g2_fill_1 FILLER_51_221 ();
 sg13g2_fill_1 FILLER_51_310 ();
 sg13g2_fill_2 FILLER_51_318 ();
 sg13g2_fill_2 FILLER_51_324 ();
 sg13g2_fill_1 FILLER_51_330 ();
 sg13g2_fill_1 FILLER_51_355 ();
 sg13g2_fill_2 FILLER_51_367 ();
 sg13g2_fill_2 FILLER_52_64 ();
 sg13g2_fill_2 FILLER_52_110 ();
 sg13g2_fill_1 FILLER_52_112 ();
 sg13g2_fill_2 FILLER_52_122 ();
 sg13g2_decap_4 FILLER_52_130 ();
 sg13g2_fill_1 FILLER_52_134 ();
 sg13g2_fill_1 FILLER_52_145 ();
 sg13g2_fill_1 FILLER_52_182 ();
 sg13g2_decap_4 FILLER_52_209 ();
 sg13g2_fill_2 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_313 ();
 sg13g2_fill_2 FILLER_52_326 ();
 sg13g2_fill_2 FILLER_52_333 ();
 sg13g2_fill_2 FILLER_52_340 ();
 sg13g2_fill_2 FILLER_52_381 ();
 sg13g2_fill_1 FILLER_53_55 ();
 sg13g2_fill_2 FILLER_53_75 ();
 sg13g2_fill_1 FILLER_53_180 ();
 sg13g2_fill_2 FILLER_53_194 ();
 sg13g2_fill_1 FILLER_53_222 ();
 sg13g2_decap_8 FILLER_53_229 ();
 sg13g2_decap_8 FILLER_53_236 ();
 sg13g2_fill_2 FILLER_53_243 ();
 sg13g2_fill_2 FILLER_53_254 ();
 sg13g2_fill_2 FILLER_53_270 ();
 sg13g2_fill_1 FILLER_53_272 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_7 ();
 sg13g2_fill_1 FILLER_54_9 ();
 sg13g2_fill_1 FILLER_54_22 ();
 sg13g2_fill_2 FILLER_54_37 ();
 sg13g2_fill_1 FILLER_54_52 ();
 sg13g2_decap_8 FILLER_54_122 ();
 sg13g2_fill_2 FILLER_54_179 ();
 sg13g2_fill_1 FILLER_54_195 ();
 sg13g2_decap_4 FILLER_54_223 ();
 sg13g2_fill_2 FILLER_54_227 ();
 sg13g2_decap_8 FILLER_54_232 ();
 sg13g2_decap_4 FILLER_54_239 ();
 sg13g2_fill_2 FILLER_54_264 ();
 sg13g2_fill_1 FILLER_54_266 ();
 sg13g2_fill_2 FILLER_54_361 ();
 sg13g2_fill_1 FILLER_54_368 ();
 sg13g2_fill_2 FILLER_54_380 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_16 ();
 sg13g2_fill_1 FILLER_55_35 ();
 sg13g2_fill_1 FILLER_55_51 ();
 sg13g2_fill_1 FILLER_55_60 ();
 sg13g2_fill_2 FILLER_55_70 ();
 sg13g2_fill_1 FILLER_55_72 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_decap_4 FILLER_55_118 ();
 sg13g2_fill_2 FILLER_55_135 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_fill_1 FILLER_55_162 ();
 sg13g2_fill_2 FILLER_55_180 ();
 sg13g2_fill_1 FILLER_55_182 ();
 sg13g2_decap_8 FILLER_55_210 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_fill_1 FILLER_55_237 ();
 sg13g2_fill_2 FILLER_55_249 ();
 sg13g2_fill_2 FILLER_55_281 ();
 sg13g2_fill_1 FILLER_55_325 ();
 sg13g2_fill_2 FILLER_55_339 ();
 sg13g2_fill_2 FILLER_56_99 ();
 sg13g2_fill_1 FILLER_56_101 ();
 sg13g2_fill_1 FILLER_56_127 ();
 sg13g2_decap_8 FILLER_56_136 ();
 sg13g2_decap_8 FILLER_56_143 ();
 sg13g2_fill_1 FILLER_56_150 ();
 sg13g2_fill_2 FILLER_56_181 ();
 sg13g2_fill_1 FILLER_56_183 ();
 sg13g2_fill_2 FILLER_56_203 ();
 sg13g2_fill_1 FILLER_56_205 ();
 sg13g2_fill_1 FILLER_56_218 ();
 sg13g2_fill_2 FILLER_56_237 ();
 sg13g2_fill_2 FILLER_56_256 ();
 sg13g2_fill_2 FILLER_56_289 ();
 sg13g2_fill_2 FILLER_56_381 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_4 ();
 sg13g2_fill_1 FILLER_57_67 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_fill_2 FILLER_57_185 ();
 sg13g2_fill_2 FILLER_57_314 ();
 sg13g2_fill_2 FILLER_57_349 ();
 sg13g2_fill_1 FILLER_57_382 ();
 sg13g2_fill_2 FILLER_58_105 ();
 sg13g2_fill_1 FILLER_58_123 ();
 sg13g2_fill_1 FILLER_58_150 ();
 sg13g2_decap_4 FILLER_58_165 ();
 sg13g2_fill_1 FILLER_58_169 ();
 sg13g2_fill_1 FILLER_58_178 ();
 sg13g2_fill_2 FILLER_58_280 ();
 sg13g2_fill_2 FILLER_58_294 ();
 sg13g2_fill_2 FILLER_58_353 ();
 sg13g2_fill_1 FILLER_58_391 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_2 FILLER_59_45 ();
 sg13g2_fill_2 FILLER_59_63 ();
 sg13g2_fill_1 FILLER_59_95 ();
 sg13g2_fill_1 FILLER_59_120 ();
 sg13g2_fill_1 FILLER_59_213 ();
 sg13g2_fill_2 FILLER_59_218 ();
 sg13g2_fill_1 FILLER_59_220 ();
 sg13g2_fill_1 FILLER_59_233 ();
 sg13g2_fill_2 FILLER_59_243 ();
 sg13g2_fill_2 FILLER_59_289 ();
 sg13g2_fill_2 FILLER_59_322 ();
 sg13g2_fill_2 FILLER_59_351 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_fill_2 FILLER_60_23 ();
 sg13g2_fill_1 FILLER_60_44 ();
 sg13g2_fill_1 FILLER_60_50 ();
 sg13g2_fill_2 FILLER_60_103 ();
 sg13g2_fill_2 FILLER_60_121 ();
 sg13g2_fill_1 FILLER_60_123 ();
 sg13g2_fill_1 FILLER_60_130 ();
 sg13g2_fill_1 FILLER_60_141 ();
 sg13g2_fill_2 FILLER_60_152 ();
 sg13g2_fill_1 FILLER_60_154 ();
 sg13g2_fill_2 FILLER_60_207 ();
 sg13g2_fill_1 FILLER_60_209 ();
 sg13g2_fill_1 FILLER_60_218 ();
 sg13g2_fill_1 FILLER_60_239 ();
 sg13g2_fill_2 FILLER_60_250 ();
 sg13g2_fill_2 FILLER_60_315 ();
 sg13g2_fill_1 FILLER_60_317 ();
 sg13g2_fill_2 FILLER_60_327 ();
 sg13g2_fill_2 FILLER_60_338 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_25 ();
 sg13g2_fill_2 FILLER_61_32 ();
 sg13g2_fill_1 FILLER_61_34 ();
 sg13g2_fill_2 FILLER_61_47 ();
 sg13g2_fill_1 FILLER_61_49 ();
 sg13g2_fill_2 FILLER_61_55 ();
 sg13g2_fill_1 FILLER_61_82 ();
 sg13g2_fill_2 FILLER_61_114 ();
 sg13g2_fill_1 FILLER_61_116 ();
 sg13g2_fill_2 FILLER_61_130 ();
 sg13g2_fill_1 FILLER_61_132 ();
 sg13g2_fill_2 FILLER_61_149 ();
 sg13g2_fill_2 FILLER_61_193 ();
 sg13g2_decap_4 FILLER_61_208 ();
 sg13g2_fill_2 FILLER_61_229 ();
 sg13g2_fill_1 FILLER_61_238 ();
 sg13g2_fill_1 FILLER_61_304 ();
 sg13g2_fill_1 FILLER_61_314 ();
 sg13g2_fill_1 FILLER_61_342 ();
 sg13g2_fill_2 FILLER_61_351 ();
 sg13g2_fill_2 FILLER_61_361 ();
 sg13g2_fill_2 FILLER_62_45 ();
 sg13g2_fill_1 FILLER_62_89 ();
 sg13g2_fill_2 FILLER_62_175 ();
 sg13g2_fill_1 FILLER_62_177 ();
 sg13g2_fill_2 FILLER_62_229 ();
 sg13g2_fill_2 FILLER_62_281 ();
 sg13g2_fill_1 FILLER_62_283 ();
 sg13g2_fill_2 FILLER_62_360 ();
 sg13g2_fill_2 FILLER_62_388 ();
 sg13g2_fill_1 FILLER_62_399 ();
 sg13g2_fill_2 FILLER_63_68 ();
 sg13g2_fill_2 FILLER_63_169 ();
 sg13g2_fill_1 FILLER_63_171 ();
 sg13g2_fill_2 FILLER_63_279 ();
 sg13g2_fill_1 FILLER_64_60 ();
 sg13g2_fill_2 FILLER_64_79 ();
 sg13g2_fill_2 FILLER_64_117 ();
 sg13g2_fill_2 FILLER_64_124 ();
 sg13g2_decap_8 FILLER_64_137 ();
 sg13g2_fill_1 FILLER_64_144 ();
 sg13g2_fill_1 FILLER_64_155 ();
 sg13g2_fill_2 FILLER_64_186 ();
 sg13g2_fill_2 FILLER_64_193 ();
 sg13g2_fill_1 FILLER_64_195 ();
 sg13g2_decap_4 FILLER_64_211 ();
 sg13g2_decap_4 FILLER_64_259 ();
 sg13g2_fill_1 FILLER_64_263 ();
 sg13g2_fill_1 FILLER_64_310 ();
 sg13g2_fill_1 FILLER_64_343 ();
 sg13g2_fill_1 FILLER_64_382 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_fill_1 FILLER_65_14 ();
 sg13g2_fill_2 FILLER_65_97 ();
 sg13g2_fill_2 FILLER_65_107 ();
 sg13g2_fill_1 FILLER_65_114 ();
 sg13g2_fill_2 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_132 ();
 sg13g2_fill_2 FILLER_65_149 ();
 sg13g2_fill_2 FILLER_65_165 ();
 sg13g2_fill_1 FILLER_65_167 ();
 sg13g2_fill_1 FILLER_65_233 ();
 sg13g2_decap_4 FILLER_65_242 ();
 sg13g2_fill_1 FILLER_65_246 ();
 sg13g2_decap_4 FILLER_65_252 ();
 sg13g2_fill_2 FILLER_65_338 ();
 sg13g2_fill_2 FILLER_65_361 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_fill_1 FILLER_66_21 ();
 sg13g2_fill_2 FILLER_66_32 ();
 sg13g2_fill_1 FILLER_66_34 ();
 sg13g2_fill_1 FILLER_66_109 ();
 sg13g2_fill_1 FILLER_66_128 ();
 sg13g2_fill_1 FILLER_66_132 ();
 sg13g2_fill_2 FILLER_66_166 ();
 sg13g2_fill_1 FILLER_66_181 ();
 sg13g2_fill_2 FILLER_66_248 ();
 sg13g2_fill_1 FILLER_66_250 ();
 sg13g2_fill_1 FILLER_66_264 ();
 sg13g2_fill_1 FILLER_66_274 ();
 sg13g2_fill_2 FILLER_66_311 ();
 sg13g2_fill_2 FILLER_66_340 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_41 ();
 sg13g2_fill_1 FILLER_67_43 ();
 sg13g2_decap_8 FILLER_67_58 ();
 sg13g2_decap_4 FILLER_67_65 ();
 sg13g2_fill_1 FILLER_67_69 ();
 sg13g2_fill_1 FILLER_67_83 ();
 sg13g2_fill_1 FILLER_67_202 ();
 sg13g2_fill_2 FILLER_67_221 ();
 sg13g2_fill_2 FILLER_67_294 ();
 sg13g2_fill_2 FILLER_67_315 ();
 sg13g2_fill_1 FILLER_67_322 ();
 sg13g2_fill_2 FILLER_67_363 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_decap_4 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_68 ();
 sg13g2_fill_2 FILLER_68_75 ();
 sg13g2_fill_2 FILLER_68_87 ();
 sg13g2_fill_1 FILLER_68_89 ();
 sg13g2_fill_1 FILLER_68_142 ();
 sg13g2_fill_1 FILLER_68_160 ();
 sg13g2_fill_1 FILLER_68_210 ();
 sg13g2_fill_2 FILLER_68_220 ();
 sg13g2_fill_1 FILLER_68_280 ();
 sg13g2_fill_1 FILLER_68_325 ();
 sg13g2_fill_1 FILLER_68_342 ();
 sg13g2_fill_2 FILLER_68_392 ();
 sg13g2_decap_4 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_4 ();
 sg13g2_fill_1 FILLER_69_43 ();
 sg13g2_decap_4 FILLER_69_70 ();
 sg13g2_decap_4 FILLER_69_84 ();
 sg13g2_fill_1 FILLER_69_88 ();
 sg13g2_fill_1 FILLER_69_115 ();
 sg13g2_fill_1 FILLER_69_174 ();
 sg13g2_fill_1 FILLER_69_188 ();
 sg13g2_fill_2 FILLER_69_194 ();
 sg13g2_fill_2 FILLER_69_280 ();
 sg13g2_fill_2 FILLER_69_292 ();
 sg13g2_fill_2 FILLER_69_304 ();
 sg13g2_fill_2 FILLER_69_338 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_4 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_24 ();
 sg13g2_fill_2 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_84 ();
 sg13g2_fill_2 FILLER_70_112 ();
 sg13g2_fill_1 FILLER_70_114 ();
 sg13g2_decap_4 FILLER_70_123 ();
 sg13g2_fill_2 FILLER_70_127 ();
 sg13g2_fill_2 FILLER_70_164 ();
 sg13g2_fill_2 FILLER_70_246 ();
 sg13g2_fill_2 FILLER_70_324 ();
 sg13g2_fill_1 FILLER_70_342 ();
 sg13g2_fill_2 FILLER_70_381 ();
 sg13g2_decap_4 FILLER_71_0 ();
 sg13g2_decap_4 FILLER_71_30 ();
 sg13g2_fill_1 FILLER_71_34 ();
 sg13g2_fill_1 FILLER_71_48 ();
 sg13g2_decap_8 FILLER_71_53 ();
 sg13g2_fill_2 FILLER_71_60 ();
 sg13g2_fill_1 FILLER_71_62 ();
 sg13g2_decap_8 FILLER_71_94 ();
 sg13g2_decap_8 FILLER_71_101 ();
 sg13g2_decap_4 FILLER_71_108 ();
 sg13g2_decap_4 FILLER_71_117 ();
 sg13g2_decap_4 FILLER_71_143 ();
 sg13g2_fill_1 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_152 ();
 sg13g2_fill_2 FILLER_71_159 ();
 sg13g2_fill_1 FILLER_71_161 ();
 sg13g2_fill_2 FILLER_71_168 ();
 sg13g2_fill_1 FILLER_71_170 ();
 sg13g2_fill_1 FILLER_71_179 ();
 sg13g2_fill_2 FILLER_71_200 ();
 sg13g2_fill_2 FILLER_71_224 ();
 sg13g2_fill_1 FILLER_71_245 ();
 sg13g2_fill_1 FILLER_71_267 ();
 sg13g2_fill_2 FILLER_71_327 ();
 sg13g2_fill_1 FILLER_71_382 ();
 sg13g2_decap_4 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_30 ();
 sg13g2_fill_2 FILLER_72_99 ();
 sg13g2_decap_8 FILLER_72_127 ();
 sg13g2_decap_4 FILLER_72_134 ();
 sg13g2_fill_1 FILLER_72_138 ();
 sg13g2_decap_4 FILLER_72_148 ();
 sg13g2_fill_1 FILLER_72_160 ();
 sg13g2_decap_8 FILLER_72_175 ();
 sg13g2_fill_2 FILLER_72_182 ();
 sg13g2_fill_2 FILLER_72_200 ();
 sg13g2_fill_1 FILLER_72_202 ();
 sg13g2_fill_2 FILLER_72_217 ();
 sg13g2_fill_1 FILLER_72_219 ();
 sg13g2_fill_2 FILLER_72_229 ();
 sg13g2_fill_2 FILLER_72_314 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_4 ();
 sg13g2_decap_4 FILLER_73_24 ();
 sg13g2_fill_2 FILLER_73_28 ();
 sg13g2_fill_2 FILLER_73_76 ();
 sg13g2_fill_2 FILLER_73_154 ();
 sg13g2_decap_4 FILLER_73_174 ();
 sg13g2_fill_1 FILLER_73_178 ();
 sg13g2_fill_1 FILLER_73_250 ();
 sg13g2_fill_1 FILLER_73_256 ();
 sg13g2_fill_1 FILLER_73_266 ();
 sg13g2_fill_1 FILLER_73_323 ();
 sg13g2_fill_2 FILLER_73_350 ();
 sg13g2_fill_1 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_74_29 ();
 sg13g2_fill_2 FILLER_74_36 ();
 sg13g2_fill_1 FILLER_74_38 ();
 sg13g2_decap_8 FILLER_74_44 ();
 sg13g2_decap_8 FILLER_74_51 ();
 sg13g2_decap_8 FILLER_74_58 ();
 sg13g2_fill_2 FILLER_74_74 ();
 sg13g2_decap_4 FILLER_74_80 ();
 sg13g2_fill_2 FILLER_74_110 ();
 sg13g2_fill_1 FILLER_74_120 ();
 sg13g2_fill_1 FILLER_74_224 ();
 sg13g2_fill_2 FILLER_74_239 ();
 sg13g2_fill_1 FILLER_74_241 ();
 sg13g2_fill_2 FILLER_74_323 ();
 sg13g2_fill_1 FILLER_74_336 ();
 sg13g2_fill_2 FILLER_74_342 ();
 sg13g2_fill_2 FILLER_74_387 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_4 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_4 ();
 sg13g2_decap_4 FILLER_75_61 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_fill_1 FILLER_75_112 ();
 sg13g2_fill_1 FILLER_75_339 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_fill_2 FILLER_76_21 ();
 sg13g2_decap_4 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_50 ();
 sg13g2_fill_2 FILLER_76_57 ();
 sg13g2_decap_4 FILLER_76_69 ();
 sg13g2_fill_2 FILLER_76_73 ();
 sg13g2_fill_2 FILLER_76_79 ();
 sg13g2_decap_8 FILLER_76_100 ();
 sg13g2_fill_1 FILLER_76_107 ();
 sg13g2_fill_1 FILLER_76_138 ();
 sg13g2_fill_2 FILLER_76_155 ();
 sg13g2_fill_1 FILLER_76_203 ();
 sg13g2_fill_1 FILLER_76_218 ();
 sg13g2_fill_2 FILLER_76_224 ();
 sg13g2_fill_1 FILLER_76_272 ();
 sg13g2_fill_1 FILLER_76_333 ();
 sg13g2_fill_1 FILLER_77_26 ();
 sg13g2_fill_2 FILLER_77_38 ();
 sg13g2_decap_4 FILLER_77_76 ();
 sg13g2_fill_1 FILLER_77_80 ();
 sg13g2_fill_1 FILLER_77_117 ();
 sg13g2_fill_1 FILLER_77_122 ();
 sg13g2_fill_1 FILLER_77_213 ();
 sg13g2_fill_1 FILLER_77_231 ();
 sg13g2_fill_2 FILLER_77_262 ();
 sg13g2_fill_2 FILLER_78_161 ();
 sg13g2_fill_1 FILLER_78_163 ();
 sg13g2_fill_2 FILLER_78_195 ();
 sg13g2_fill_1 FILLER_78_319 ();
 sg13g2_decap_4 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_23 ();
 sg13g2_fill_1 FILLER_79_29 ();
 sg13g2_fill_1 FILLER_79_91 ();
 sg13g2_fill_1 FILLER_79_135 ();
 sg13g2_fill_2 FILLER_79_169 ();
 sg13g2_fill_1 FILLER_79_171 ();
 sg13g2_fill_2 FILLER_79_237 ();
 sg13g2_fill_2 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_fill_1 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_40 ();
 sg13g2_decap_4 FILLER_80_47 ();
 sg13g2_fill_1 FILLER_80_51 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_fill_2 FILLER_80_125 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_fill_1 FILLER_80_132 ();
 sg13g2_fill_2 FILLER_80_193 ();
 sg13g2_fill_2 FILLER_80_226 ();
 sg13g2_fill_1 FILLER_80_228 ();
 sg13g2_fill_2 FILLER_80_252 ();
 sg13g2_fill_2 FILLER_80_272 ();
 sg13g2_fill_2 FILLER_80_294 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_351 ();
 assign uio_oe[0] = net30;
 assign uio_oe[1] = net31;
 assign uio_oe[2] = net32;
 assign uio_oe[3] = net33;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net34;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[1] = net9;
 assign uio_out[2] = net10;
 assign uio_out[4] = net11;
 assign uio_out[5] = net12;
 assign uio_out[6] = net13;
 assign uio_out[7] = net14;
endmodule
