module tt_um_ds_comp_adc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire \cic_a.decim_cnt[0] ;
 wire \cic_a.decim_cnt[1] ;
 wire \cic_a.decim_cnt[2] ;
 wire \cic_a.decim_cnt[3] ;
 wire \cic_a.decim_cnt[4] ;
 wire \cic_a.decim_cnt[5] ;
 wire \cic_a.decim_cnt[6] ;
 wire \cic_a.decim_cnt[7] ;
 wire \cic_a.delay[0][0] ;
 wire \cic_a.delay[0][10] ;
 wire \cic_a.delay[0][11] ;
 wire \cic_a.delay[0][12] ;
 wire \cic_a.delay[0][1] ;
 wire \cic_a.delay[0][2] ;
 wire \cic_a.delay[0][3] ;
 wire \cic_a.delay[0][4] ;
 wire \cic_a.delay[0][5] ;
 wire \cic_a.delay[0][6] ;
 wire \cic_a.delay[0][7] ;
 wire \cic_a.delay[0][8] ;
 wire \cic_a.delay[0][9] ;
 wire \cic_a.delay[1][0] ;
 wire \cic_a.delay[1][10] ;
 wire \cic_a.delay[1][11] ;
 wire \cic_a.delay[1][12] ;
 wire \cic_a.delay[1][1] ;
 wire \cic_a.delay[1][2] ;
 wire \cic_a.delay[1][3] ;
 wire \cic_a.delay[1][4] ;
 wire \cic_a.delay[1][5] ;
 wire \cic_a.delay[1][6] ;
 wire \cic_a.delay[1][7] ;
 wire \cic_a.delay[1][8] ;
 wire \cic_a.delay[1][9] ;
 wire \cic_a.filtered_out[0] ;
 wire \cic_a.filtered_out[10] ;
 wire \cic_a.filtered_out[11] ;
 wire \cic_a.filtered_out[12] ;
 wire \cic_a.filtered_out[1] ;
 wire \cic_a.filtered_out[2] ;
 wire \cic_a.filtered_out[3] ;
 wire \cic_a.filtered_out[4] ;
 wire \cic_a.filtered_out[5] ;
 wire \cic_a.filtered_out[6] ;
 wire \cic_a.filtered_out[7] ;
 wire \cic_a.filtered_out[8] ;
 wire \cic_a.filtered_out[9] ;
 wire \cic_a.integrator[0][0] ;
 wire \cic_a.integrator[0][10] ;
 wire \cic_a.integrator[0][11] ;
 wire \cic_a.integrator[0][12] ;
 wire \cic_a.integrator[0][1] ;
 wire \cic_a.integrator[0][2] ;
 wire \cic_a.integrator[0][3] ;
 wire \cic_a.integrator[0][4] ;
 wire \cic_a.integrator[0][5] ;
 wire \cic_a.integrator[0][6] ;
 wire \cic_a.integrator[0][7] ;
 wire \cic_a.integrator[0][8] ;
 wire \cic_a.integrator[0][9] ;
 wire \cic_a.integrator[1][0] ;
 wire \cic_a.integrator[1][10] ;
 wire \cic_a.integrator[1][11] ;
 wire \cic_a.integrator[1][12] ;
 wire \cic_a.integrator[1][1] ;
 wire \cic_a.integrator[1][2] ;
 wire \cic_a.integrator[1][3] ;
 wire \cic_a.integrator[1][4] ;
 wire \cic_a.integrator[1][5] ;
 wire \cic_a.integrator[1][6] ;
 wire \cic_a.integrator[1][7] ;
 wire \cic_a.integrator[1][8] ;
 wire \cic_a.integrator[1][9] ;
 wire \cic_a.pdm_in ;
 wire \cic_a.temp_comb[0][0] ;
 wire \cic_a.temp_comb[0][10] ;
 wire \cic_a.temp_comb[0][11] ;
 wire \cic_a.temp_comb[0][12] ;
 wire \cic_a.temp_comb[0][1] ;
 wire \cic_a.temp_comb[0][2] ;
 wire \cic_a.temp_comb[0][3] ;
 wire \cic_a.temp_comb[0][4] ;
 wire \cic_a.temp_comb[0][5] ;
 wire \cic_a.temp_comb[0][6] ;
 wire \cic_a.temp_comb[0][7] ;
 wire \cic_a.temp_comb[0][8] ;
 wire \cic_a.temp_comb[0][9] ;
 wire \cic_a.temp_comb[1][0] ;
 wire \cic_a.temp_comb[1][10] ;
 wire \cic_a.temp_comb[1][11] ;
 wire \cic_a.temp_comb[1][12] ;
 wire \cic_a.temp_comb[1][1] ;
 wire \cic_a.temp_comb[1][2] ;
 wire \cic_a.temp_comb[1][3] ;
 wire \cic_a.temp_comb[1][4] ;
 wire \cic_a.temp_comb[1][5] ;
 wire \cic_a.temp_comb[1][6] ;
 wire \cic_a.temp_comb[1][7] ;
 wire \cic_a.temp_comb[1][8] ;
 wire \cic_a.temp_comb[1][9] ;
 wire \cic_a.temp_delay[0][0] ;
 wire \cic_a.temp_delay[0][10] ;
 wire \cic_a.temp_delay[0][11] ;
 wire \cic_a.temp_delay[0][12] ;
 wire \cic_a.temp_delay[0][1] ;
 wire \cic_a.temp_delay[0][2] ;
 wire \cic_a.temp_delay[0][3] ;
 wire \cic_a.temp_delay[0][4] ;
 wire \cic_a.temp_delay[0][5] ;
 wire \cic_a.temp_delay[0][6] ;
 wire \cic_a.temp_delay[0][7] ;
 wire \cic_a.temp_delay[0][8] ;
 wire \cic_a.temp_delay[0][9] ;
 wire \cic_a.temp_delay[1][0] ;
 wire \cic_a.temp_delay[1][10] ;
 wire \cic_a.temp_delay[1][11] ;
 wire \cic_a.temp_delay[1][12] ;
 wire \cic_a.temp_delay[1][1] ;
 wire \cic_a.temp_delay[1][2] ;
 wire \cic_a.temp_delay[1][3] ;
 wire \cic_a.temp_delay[1][4] ;
 wire \cic_a.temp_delay[1][5] ;
 wire \cic_a.temp_delay[1][6] ;
 wire \cic_a.temp_delay[1][7] ;
 wire \cic_a.temp_delay[1][8] ;
 wire \cic_a.temp_delay[1][9] ;
 wire \cic_b.decim_cnt[0] ;
 wire \cic_b.decim_cnt[1] ;
 wire \cic_b.decim_cnt[2] ;
 wire \cic_b.decim_cnt[3] ;
 wire \cic_b.decim_cnt[4] ;
 wire \cic_b.decim_cnt[5] ;
 wire \cic_b.decim_cnt[6] ;
 wire \cic_b.decim_cnt[7] ;
 wire \cic_b.delay[0][0] ;
 wire \cic_b.delay[0][10] ;
 wire \cic_b.delay[0][11] ;
 wire \cic_b.delay[0][12] ;
 wire \cic_b.delay[0][1] ;
 wire \cic_b.delay[0][2] ;
 wire \cic_b.delay[0][3] ;
 wire \cic_b.delay[0][4] ;
 wire \cic_b.delay[0][5] ;
 wire \cic_b.delay[0][6] ;
 wire \cic_b.delay[0][7] ;
 wire \cic_b.delay[0][8] ;
 wire \cic_b.delay[0][9] ;
 wire \cic_b.delay[1][0] ;
 wire \cic_b.delay[1][10] ;
 wire \cic_b.delay[1][11] ;
 wire \cic_b.delay[1][12] ;
 wire \cic_b.delay[1][1] ;
 wire \cic_b.delay[1][2] ;
 wire \cic_b.delay[1][3] ;
 wire \cic_b.delay[1][4] ;
 wire \cic_b.delay[1][5] ;
 wire \cic_b.delay[1][6] ;
 wire \cic_b.delay[1][7] ;
 wire \cic_b.delay[1][8] ;
 wire \cic_b.delay[1][9] ;
 wire \cic_b.filtered_out[0] ;
 wire \cic_b.filtered_out[10] ;
 wire \cic_b.filtered_out[11] ;
 wire \cic_b.filtered_out[12] ;
 wire \cic_b.filtered_out[1] ;
 wire \cic_b.filtered_out[2] ;
 wire \cic_b.filtered_out[3] ;
 wire \cic_b.filtered_out[4] ;
 wire \cic_b.filtered_out[5] ;
 wire \cic_b.filtered_out[6] ;
 wire \cic_b.filtered_out[7] ;
 wire \cic_b.filtered_out[8] ;
 wire \cic_b.filtered_out[9] ;
 wire \cic_b.integrator[0][0] ;
 wire \cic_b.integrator[0][10] ;
 wire \cic_b.integrator[0][11] ;
 wire \cic_b.integrator[0][12] ;
 wire \cic_b.integrator[0][1] ;
 wire \cic_b.integrator[0][2] ;
 wire \cic_b.integrator[0][3] ;
 wire \cic_b.integrator[0][4] ;
 wire \cic_b.integrator[0][5] ;
 wire \cic_b.integrator[0][6] ;
 wire \cic_b.integrator[0][7] ;
 wire \cic_b.integrator[0][8] ;
 wire \cic_b.integrator[0][9] ;
 wire \cic_b.integrator[1][0] ;
 wire \cic_b.integrator[1][10] ;
 wire \cic_b.integrator[1][11] ;
 wire \cic_b.integrator[1][12] ;
 wire \cic_b.integrator[1][1] ;
 wire \cic_b.integrator[1][2] ;
 wire \cic_b.integrator[1][3] ;
 wire \cic_b.integrator[1][4] ;
 wire \cic_b.integrator[1][5] ;
 wire \cic_b.integrator[1][6] ;
 wire \cic_b.integrator[1][7] ;
 wire \cic_b.integrator[1][8] ;
 wire \cic_b.integrator[1][9] ;
 wire \cic_b.pdm_in ;
 wire \cic_b.temp_comb[0][0] ;
 wire \cic_b.temp_comb[0][10] ;
 wire \cic_b.temp_comb[0][11] ;
 wire \cic_b.temp_comb[0][12] ;
 wire \cic_b.temp_comb[0][1] ;
 wire \cic_b.temp_comb[0][2] ;
 wire \cic_b.temp_comb[0][3] ;
 wire \cic_b.temp_comb[0][4] ;
 wire \cic_b.temp_comb[0][5] ;
 wire \cic_b.temp_comb[0][6] ;
 wire \cic_b.temp_comb[0][7] ;
 wire \cic_b.temp_comb[0][8] ;
 wire \cic_b.temp_comb[0][9] ;
 wire \cic_b.temp_comb[1][0] ;
 wire \cic_b.temp_comb[1][10] ;
 wire \cic_b.temp_comb[1][11] ;
 wire \cic_b.temp_comb[1][12] ;
 wire \cic_b.temp_comb[1][1] ;
 wire \cic_b.temp_comb[1][2] ;
 wire \cic_b.temp_comb[1][3] ;
 wire \cic_b.temp_comb[1][4] ;
 wire \cic_b.temp_comb[1][5] ;
 wire \cic_b.temp_comb[1][6] ;
 wire \cic_b.temp_comb[1][7] ;
 wire \cic_b.temp_comb[1][8] ;
 wire \cic_b.temp_comb[1][9] ;
 wire \cic_b.temp_delay[0][0] ;
 wire \cic_b.temp_delay[0][10] ;
 wire \cic_b.temp_delay[0][11] ;
 wire \cic_b.temp_delay[0][12] ;
 wire \cic_b.temp_delay[0][1] ;
 wire \cic_b.temp_delay[0][2] ;
 wire \cic_b.temp_delay[0][3] ;
 wire \cic_b.temp_delay[0][4] ;
 wire \cic_b.temp_delay[0][5] ;
 wire \cic_b.temp_delay[0][6] ;
 wire \cic_b.temp_delay[0][7] ;
 wire \cic_b.temp_delay[0][8] ;
 wire \cic_b.temp_delay[0][9] ;
 wire \cic_b.temp_delay[1][0] ;
 wire \cic_b.temp_delay[1][10] ;
 wire \cic_b.temp_delay[1][11] ;
 wire \cic_b.temp_delay[1][12] ;
 wire \cic_b.temp_delay[1][1] ;
 wire \cic_b.temp_delay[1][2] ;
 wire \cic_b.temp_delay[1][3] ;
 wire \cic_b.temp_delay[1][4] ;
 wire \cic_b.temp_delay[1][5] ;
 wire \cic_b.temp_delay[1][6] ;
 wire \cic_b.temp_delay[1][7] ;
 wire \cic_b.temp_delay[1][8] ;
 wire \cic_b.temp_delay[1][9] ;
 wire pdm_a;
 wire pdm_b;
 wire \serializer_a.bit_cnt[0] ;
 wire \serializer_a.bit_cnt[1] ;
 wire \serializer_a.bit_cnt[2] ;
 wire \serializer_a.bit_cnt[3] ;
 wire \serializer_a.sending ;
 wire \serializer_a.serial_out ;
 wire \serializer_a.shift_reg[0] ;
 wire \serializer_a.shift_reg[10] ;
 wire \serializer_a.shift_reg[11] ;
 wire \serializer_a.shift_reg[1] ;
 wire \serializer_a.shift_reg[2] ;
 wire \serializer_a.shift_reg[3] ;
 wire \serializer_a.shift_reg[4] ;
 wire \serializer_a.shift_reg[5] ;
 wire \serializer_a.shift_reg[6] ;
 wire \serializer_a.shift_reg[7] ;
 wire \serializer_a.shift_reg[8] ;
 wire \serializer_a.shift_reg[9] ;
 wire \serializer_a.valid ;
 wire \serializer_ab_subtr.bit_cnt[0] ;
 wire \serializer_ab_subtr.bit_cnt[1] ;
 wire \serializer_ab_subtr.bit_cnt[2] ;
 wire \serializer_ab_subtr.bit_cnt[3] ;
 wire \serializer_ab_subtr.sending ;
 wire \serializer_ab_subtr.serial_out ;
 wire \serializer_ab_subtr.shift_reg[0] ;
 wire \serializer_ab_subtr.shift_reg[10] ;
 wire \serializer_ab_subtr.shift_reg[11] ;
 wire \serializer_ab_subtr.shift_reg[1] ;
 wire \serializer_ab_subtr.shift_reg[2] ;
 wire \serializer_ab_subtr.shift_reg[3] ;
 wire \serializer_ab_subtr.shift_reg[4] ;
 wire \serializer_ab_subtr.shift_reg[5] ;
 wire \serializer_ab_subtr.shift_reg[6] ;
 wire \serializer_ab_subtr.shift_reg[7] ;
 wire \serializer_ab_subtr.shift_reg[8] ;
 wire \serializer_ab_subtr.shift_reg[9] ;
 wire \serializer_ab_subtr.valid ;
 wire \serializer_b.bit_cnt[0] ;
 wire \serializer_b.bit_cnt[1] ;
 wire \serializer_b.bit_cnt[2] ;
 wire \serializer_b.bit_cnt[3] ;
 wire \serializer_b.sending ;
 wire \serializer_b.serial_out ;
 wire \serializer_b.shift_reg[0] ;
 wire \serializer_b.shift_reg[10] ;
 wire \serializer_b.shift_reg[11] ;
 wire \serializer_b.shift_reg[1] ;
 wire \serializer_b.shift_reg[2] ;
 wire \serializer_b.shift_reg[3] ;
 wire \serializer_b.shift_reg[4] ;
 wire \serializer_b.shift_reg[5] ;
 wire \serializer_b.shift_reg[6] ;
 wire \serializer_b.shift_reg[7] ;
 wire \serializer_b.shift_reg[8] ;
 wire \serializer_b.shift_reg[9] ;
 wire \serializer_b.valid ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_leaf_0_clk;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;

 sg13g2_inv_1 _1270_ (.Y(_0077_),
    .A(net2));
 sg13g2_inv_1 _1271_ (.Y(_0076_),
    .A(net1));
 sg13g2_inv_1 _1272_ (.Y(_0000_),
    .A(net24));
 sg13g2_inv_1 _1273_ (.Y(_0689_),
    .A(\cic_a.decim_cnt[3] ));
 sg13g2_inv_1 _1274_ (.Y(_0008_),
    .A(net23));
 sg13g2_inv_1 _1275_ (.Y(_0690_),
    .A(\cic_b.decim_cnt[3] ));
 sg13g2_inv_1 _1276_ (.Y(_0691_),
    .A(net106));
 sg13g2_inv_1 _1277_ (.Y(_0692_),
    .A(net71));
 sg13g2_inv_1 _1278_ (.Y(_0693_),
    .A(\cic_a.filtered_out[4] ));
 sg13g2_inv_1 _1279_ (.Y(_0694_),
    .A(net25));
 sg13g2_inv_1 _1280_ (.Y(_0695_),
    .A(net533));
 sg13g2_inv_1 _1281_ (.Y(_0696_),
    .A(net117));
 sg13g2_inv_1 _1282_ (.Y(_0697_),
    .A(net64));
 sg13g2_inv_1 _1283_ (.Y(_0698_),
    .A(net189));
 sg13g2_inv_1 _1284_ (.Y(_0699_),
    .A(net131));
 sg13g2_inv_1 _1285_ (.Y(_0700_),
    .A(net27));
 sg13g2_inv_1 _1286_ (.Y(_0701_),
    .A(\cic_b.filtered_out[3] ));
 sg13g2_inv_1 _1287_ (.Y(_0702_),
    .A(\cic_b.filtered_out[4] ));
 sg13g2_inv_1 _1288_ (.Y(_0703_),
    .A(net119));
 sg13g2_inv_1 _1289_ (.Y(_0704_),
    .A(net149));
 sg13g2_inv_1 _1290_ (.Y(_0705_),
    .A(net221));
 sg13g2_inv_1 _1291_ (.Y(_0706_),
    .A(net122));
 sg13g2_inv_1 _1292_ (.Y(_0707_),
    .A(net506));
 sg13g2_inv_1 _1293_ (.Y(_0708_),
    .A(net246));
 sg13g2_inv_1 _1294_ (.Y(_0709_),
    .A(net134));
 sg13g2_inv_1 _1295_ (.Y(_0710_),
    .A(net219));
 sg13g2_inv_1 _1296_ (.Y(pdm_a),
    .A(\cic_a.pdm_in ));
 sg13g2_inv_1 _1297_ (.Y(pdm_b),
    .A(\cic_b.pdm_in ));
 sg13g2_inv_1 _1298_ (.Y(_0711_),
    .A(\cic_a.temp_comb[0][9] ));
 sg13g2_inv_1 _1299_ (.Y(_0712_),
    .A(net200));
 sg13g2_inv_1 _1300_ (.Y(_0713_),
    .A(net228));
 sg13g2_inv_1 _1301_ (.Y(_0714_),
    .A(\cic_a.integrator[0][6] ));
 sg13g2_inv_1 _1302_ (.Y(_0715_),
    .A(net542));
 sg13g2_inv_1 _1303_ (.Y(_0716_),
    .A(\cic_a.integrator[1][9] ));
 sg13g2_inv_1 _1304_ (.Y(_0717_),
    .A(\cic_b.delay[0][5] ));
 sg13g2_inv_1 _1305_ (.Y(_0718_),
    .A(net90));
 sg13g2_inv_1 _1306_ (.Y(_0719_),
    .A(\cic_b.delay[0][9] ));
 sg13g2_inv_1 _1307_ (.Y(_0720_),
    .A(\cic_b.temp_comb[0][5] ));
 sg13g2_inv_1 _1308_ (.Y(_0721_),
    .A(net251));
 sg13g2_inv_1 _1309_ (.Y(_0722_),
    .A(\cic_b.temp_comb[0][9] ));
 sg13g2_inv_1 _1310_ (.Y(_0723_),
    .A(net213));
 sg13g2_inv_1 _1311_ (.Y(_0724_),
    .A(net483));
 sg13g2_inv_1 _1312_ (.Y(_0725_),
    .A(\cic_b.integrator[0][6] ));
 sg13g2_inv_1 _1313_ (.Y(_0726_),
    .A(\cic_b.integrator[0][9] ));
 sg13g2_inv_1 _1314_ (.Y(_0727_),
    .A(\cic_a.delay[0][5] ));
 sg13g2_inv_1 _1315_ (.Y(_0728_),
    .A(net83));
 sg13g2_inv_1 _1316_ (.Y(_0729_),
    .A(net120));
 sg13g2_nor2b_1 _1317_ (.A(net411),
    .B_N(net3),
    .Y(_0017_));
 sg13g2_nand2b_2 _1318_ (.Y(_0730_),
    .B(net3),
    .A_N(net405));
 sg13g2_inv_2 _1319_ (.Y(_0019_),
    .A(net402));
 sg13g2_nor2b_1 _1320_ (.A(net572),
    .B_N(net3),
    .Y(_0021_));
 sg13g2_xor2_1 _1321_ (.B(net24),
    .A(net108),
    .X(_0001_));
 sg13g2_nand3_1 _1322_ (.B(net24),
    .C(net561),
    .A(net108),
    .Y(_0731_));
 sg13g2_a21o_1 _1323_ (.A2(net24),
    .A1(net108),
    .B1(net561),
    .X(_0732_));
 sg13g2_and2_1 _1324_ (.A(_0731_),
    .B(_0732_),
    .X(_0002_));
 sg13g2_nor2_1 _1325_ (.A(_0689_),
    .B(_0731_),
    .Y(_0733_));
 sg13g2_xnor2_1 _1326_ (.Y(_0003_),
    .A(net49),
    .B(_0731_));
 sg13g2_and2_2 _1327_ (.A(net35),
    .B(_0733_),
    .X(_0734_));
 sg13g2_xor2_1 _1328_ (.B(_0733_),
    .A(net35),
    .X(_0004_));
 sg13g2_nor3_2 _1329_ (.A(\cic_a.decim_cnt[5] ),
    .B(net177),
    .C(net340),
    .Y(_0735_));
 sg13g2_xnor2_1 _1330_ (.Y(_0736_),
    .A(net556),
    .B(_0734_));
 sg13g2_nor2_1 _1331_ (.A(net341),
    .B(_0736_),
    .Y(_0005_));
 sg13g2_nand3_1 _1332_ (.B(net340),
    .C(_0734_),
    .A(net556),
    .Y(_0737_));
 sg13g2_a21o_1 _1333_ (.A2(_0734_),
    .A1(net556),
    .B1(net340),
    .X(_0738_));
 sg13g2_and2_1 _1334_ (.A(_0737_),
    .B(_0738_),
    .X(_0006_));
 sg13g2_xnor2_1 _1335_ (.Y(_0007_),
    .A(net177),
    .B(_0737_));
 sg13g2_xor2_1 _1336_ (.B(net23),
    .A(net91),
    .X(_0009_));
 sg13g2_nand3_1 _1337_ (.B(net23),
    .C(net563),
    .A(net91),
    .Y(_0739_));
 sg13g2_a21o_1 _1338_ (.A2(net23),
    .A1(net91),
    .B1(net563),
    .X(_0740_));
 sg13g2_and2_1 _1339_ (.A(_0739_),
    .B(_0740_),
    .X(_0010_));
 sg13g2_nor2_1 _1340_ (.A(_0690_),
    .B(_0739_),
    .Y(_0741_));
 sg13g2_xnor2_1 _1341_ (.Y(_0011_),
    .A(net53),
    .B(_0739_));
 sg13g2_and2_1 _1342_ (.A(net29),
    .B(_0741_),
    .X(_0742_));
 sg13g2_xor2_1 _1343_ (.B(_0741_),
    .A(net29),
    .X(_0012_));
 sg13g2_nor3_1 _1344_ (.A(net547),
    .B(net57),
    .C(\cic_b.decim_cnt[6] ),
    .Y(_0743_));
 sg13g2_xnor2_1 _1345_ (.Y(_0744_),
    .A(net547),
    .B(_0742_));
 sg13g2_nor2_1 _1346_ (.A(_0743_),
    .B(_0744_),
    .Y(_0013_));
 sg13g2_nand3_1 _1347_ (.B(net568),
    .C(_0742_),
    .A(net547),
    .Y(_0745_));
 sg13g2_a21o_1 _1348_ (.A2(_0742_),
    .A1(net547),
    .B1(net568),
    .X(_0746_));
 sg13g2_and2_1 _1349_ (.A(_0745_),
    .B(_0746_),
    .X(_0014_));
 sg13g2_xnor2_1 _1350_ (.Y(_0015_),
    .A(net57),
    .B(_0745_));
 sg13g2_nand2_1 _1351_ (.Y(_0747_),
    .A(net514),
    .B(net566));
 sg13g2_nand2_1 _1352_ (.Y(_0748_),
    .A(net607),
    .B(\cic_a.integrator[1][1] ));
 sg13g2_nor2_1 _1353_ (.A(\cic_a.integrator[0][1] ),
    .B(\cic_a.integrator[1][1] ),
    .Y(_0749_));
 sg13g2_xor2_1 _1354_ (.B(net282),
    .A(\cic_a.integrator[0][1] ),
    .X(_0750_));
 sg13g2_xnor2_1 _1355_ (.Y(_0039_),
    .A(_0747_),
    .B(_0750_));
 sg13g2_and2_1 _1356_ (.A(net228),
    .B(net581),
    .X(_0751_));
 sg13g2_or2_1 _1357_ (.X(_0752_),
    .B(\cic_a.integrator[1][2] ),
    .A(net228));
 sg13g2_nand2b_1 _1358_ (.Y(_0753_),
    .B(_0752_),
    .A_N(_0751_));
 sg13g2_o21ai_1 _1359_ (.B1(_0748_),
    .Y(_0754_),
    .A1(_0747_),
    .A2(_0749_));
 sg13g2_xnor2_1 _1360_ (.Y(_0040_),
    .A(_0753_),
    .B(_0754_));
 sg13g2_a21oi_2 _1361_ (.B1(_0751_),
    .Y(_0755_),
    .A2(_0754_),
    .A1(_0752_));
 sg13g2_nand2_1 _1362_ (.Y(_0756_),
    .A(\cic_a.integrator[0][3] ),
    .B(\cic_a.integrator[1][3] ));
 sg13g2_xnor2_1 _1363_ (.Y(_0757_),
    .A(net562),
    .B(net300));
 sg13g2_xor2_1 _1364_ (.B(_0757_),
    .A(_0755_),
    .X(_0041_));
 sg13g2_nand2_1 _1365_ (.Y(_0758_),
    .A(net580),
    .B(\cic_a.integrator[1][4] ));
 sg13g2_xor2_1 _1366_ (.B(\cic_a.integrator[1][4] ),
    .A(net604),
    .X(_0759_));
 sg13g2_o21ai_1 _1367_ (.B1(_0756_),
    .Y(_0760_),
    .A1(_0755_),
    .A2(_0757_));
 sg13g2_nand2_1 _1368_ (.Y(_0761_),
    .A(_0759_),
    .B(_0760_));
 sg13g2_xor2_1 _1369_ (.B(_0760_),
    .A(net605),
    .X(_0042_));
 sg13g2_nor2_1 _1370_ (.A(net590),
    .B(\cic_a.integrator[1][5] ),
    .Y(_0762_));
 sg13g2_nand2_1 _1371_ (.Y(_0763_),
    .A(net590),
    .B(\cic_a.integrator[1][5] ));
 sg13g2_nor2b_1 _1372_ (.A(_0762_),
    .B_N(_0763_),
    .Y(_0764_));
 sg13g2_nand2_1 _1373_ (.Y(_0765_),
    .A(_0758_),
    .B(_0761_));
 sg13g2_xor2_1 _1374_ (.B(_0765_),
    .A(_0764_),
    .X(_0043_));
 sg13g2_nand2_1 _1375_ (.Y(_0766_),
    .A(\cic_a.integrator[0][6] ),
    .B(\cic_a.integrator[1][6] ));
 sg13g2_nor2_1 _1376_ (.A(\cic_a.integrator[0][6] ),
    .B(\cic_a.integrator[1][6] ),
    .Y(_0767_));
 sg13g2_xor2_1 _1377_ (.B(net328),
    .A(net552),
    .X(_0768_));
 sg13g2_nand3_1 _1378_ (.B(_0760_),
    .C(_0764_),
    .A(_0759_),
    .Y(_0769_));
 sg13g2_o21ai_1 _1379_ (.B1(_0763_),
    .Y(_0770_),
    .A1(_0758_),
    .A2(_0762_));
 sg13g2_nor2b_1 _1380_ (.A(_0770_),
    .B_N(_0769_),
    .Y(_0771_));
 sg13g2_xnor2_1 _1381_ (.Y(_0044_),
    .A(_0768_),
    .B(_0771_));
 sg13g2_nor2_1 _1382_ (.A(net602),
    .B(\cic_a.integrator[1][7] ),
    .Y(_0772_));
 sg13g2_nand2_1 _1383_ (.Y(_0773_),
    .A(net602),
    .B(net336));
 sg13g2_nand2b_1 _1384_ (.Y(_0774_),
    .B(_0773_),
    .A_N(_0772_));
 sg13g2_o21ai_1 _1385_ (.B1(_0766_),
    .Y(_0775_),
    .A1(_0767_),
    .A2(_0771_));
 sg13g2_xnor2_1 _1386_ (.Y(_0045_),
    .A(_0774_),
    .B(_0775_));
 sg13g2_o21ai_1 _1387_ (.B1(_0773_),
    .Y(_0776_),
    .A1(_0766_),
    .A2(_0772_));
 sg13g2_nor2_1 _1388_ (.A(_0770_),
    .B(_0776_),
    .Y(_0777_));
 sg13g2_a221oi_1 _1389_ (.B2(_0769_),
    .C1(_0772_),
    .B1(_0777_),
    .A1(_0767_),
    .Y(_0778_),
    .A2(_0773_));
 sg13g2_nand2_1 _1390_ (.Y(_0779_),
    .A(\cic_a.integrator[0][8] ),
    .B(\cic_a.integrator[1][8] ));
 sg13g2_xor2_1 _1391_ (.B(net599),
    .A(net582),
    .X(_0780_));
 sg13g2_inv_1 _1392_ (.Y(_0781_),
    .A(_0780_));
 sg13g2_nand2_1 _1393_ (.Y(_0782_),
    .A(_0778_),
    .B(_0780_));
 sg13g2_xnor2_1 _1394_ (.Y(_0046_),
    .A(_0778_),
    .B(_0781_));
 sg13g2_xnor2_1 _1395_ (.Y(_0783_),
    .A(net542),
    .B(net578));
 sg13g2_nand2_1 _1396_ (.Y(_0784_),
    .A(_0779_),
    .B(_0782_));
 sg13g2_xnor2_1 _1397_ (.Y(_0047_),
    .A(_0783_),
    .B(_0784_));
 sg13g2_nor2_1 _1398_ (.A(_0781_),
    .B(_0783_),
    .Y(_0785_));
 sg13g2_a21oi_1 _1399_ (.A1(_0715_),
    .A2(_0716_),
    .Y(_0786_),
    .B1(_0779_));
 sg13g2_a221oi_1 _1400_ (.B2(_0785_),
    .C1(_0786_),
    .B1(_0778_),
    .A1(\cic_a.integrator[0][9] ),
    .Y(_0787_),
    .A2(\cic_a.integrator[1][9] ));
 sg13g2_nand2_1 _1401_ (.Y(_0788_),
    .A(net545),
    .B(\cic_a.integrator[1][10] ));
 sg13g2_xnor2_1 _1402_ (.Y(_0789_),
    .A(net545),
    .B(net594));
 sg13g2_xor2_1 _1403_ (.B(_0789_),
    .A(_0787_),
    .X(_0036_));
 sg13g2_nor2_1 _1404_ (.A(\cic_a.integrator[0][11] ),
    .B(\cic_a.integrator[1][11] ),
    .Y(_0790_));
 sg13g2_xnor2_1 _1405_ (.Y(_0791_),
    .A(net584),
    .B(net592));
 sg13g2_o21ai_1 _1406_ (.B1(_0788_),
    .Y(_0792_),
    .A1(_0787_),
    .A2(_0789_));
 sg13g2_xnor2_1 _1407_ (.Y(_0037_),
    .A(_0791_),
    .B(_0792_));
 sg13g2_or2_1 _1408_ (.X(_0793_),
    .B(_0791_),
    .A(_0789_));
 sg13g2_nor2_1 _1409_ (.A(_0788_),
    .B(_0790_),
    .Y(_0794_));
 sg13g2_a21oi_1 _1410_ (.A1(\cic_a.integrator[0][11] ),
    .A2(\cic_a.integrator[1][11] ),
    .Y(_0795_),
    .B1(_0794_));
 sg13g2_o21ai_1 _1411_ (.B1(_0795_),
    .Y(_0796_),
    .A1(_0787_),
    .A2(_0793_));
 sg13g2_xnor2_1 _1412_ (.Y(_0797_),
    .A(net139),
    .B(net564));
 sg13g2_xnor2_1 _1413_ (.Y(_0038_),
    .A(_0796_),
    .B(_0797_));
 sg13g2_xor2_1 _1414_ (.B(\cic_a.integrator[0][0] ),
    .A(net514),
    .X(_0035_));
 sg13g2_nand2_1 _1415_ (.Y(_0798_),
    .A(net570),
    .B(net525));
 sg13g2_nand2_1 _1416_ (.Y(_0799_),
    .A(\cic_b.integrator[1][1] ),
    .B(\cic_b.integrator[0][1] ));
 sg13g2_nor2_1 _1417_ (.A(\cic_b.integrator[1][1] ),
    .B(\cic_b.integrator[0][1] ),
    .Y(_0800_));
 sg13g2_xor2_1 _1418_ (.B(\cic_b.integrator[0][1] ),
    .A(net513),
    .X(_0801_));
 sg13g2_xnor2_1 _1419_ (.Y(_0065_),
    .A(_0798_),
    .B(_0801_));
 sg13g2_and2_1 _1420_ (.A(net532),
    .B(net483),
    .X(_0802_));
 sg13g2_or2_1 _1421_ (.X(_0803_),
    .B(net608),
    .A(\cic_b.integrator[1][2] ));
 sg13g2_nand2b_1 _1422_ (.Y(_0804_),
    .B(net609),
    .A_N(_0802_));
 sg13g2_o21ai_1 _1423_ (.B1(_0799_),
    .Y(_0805_),
    .A1(_0798_),
    .A2(_0800_));
 sg13g2_xnor2_1 _1424_ (.Y(_0066_),
    .A(_0804_),
    .B(_0805_));
 sg13g2_a21oi_2 _1425_ (.B1(_0802_),
    .Y(_0806_),
    .A2(_0805_),
    .A1(_0803_));
 sg13g2_nand2_1 _1426_ (.Y(_0807_),
    .A(\cic_b.integrator[1][3] ),
    .B(net596));
 sg13g2_xnor2_1 _1427_ (.Y(_0808_),
    .A(net588),
    .B(net560));
 sg13g2_xor2_1 _1428_ (.B(_0808_),
    .A(_0806_),
    .X(_0067_));
 sg13g2_nand2_1 _1429_ (.Y(_0809_),
    .A(net346),
    .B(net583));
 sg13g2_xor2_1 _1430_ (.B(net583),
    .A(\cic_b.integrator[1][4] ),
    .X(_0810_));
 sg13g2_o21ai_1 _1431_ (.B1(net597),
    .Y(_0811_),
    .A1(_0806_),
    .A2(_0808_));
 sg13g2_nand2_1 _1432_ (.Y(_0812_),
    .A(_0810_),
    .B(_0811_));
 sg13g2_xor2_1 _1433_ (.B(_0811_),
    .A(_0810_),
    .X(_0068_));
 sg13g2_nor2_1 _1434_ (.A(\cic_b.integrator[1][5] ),
    .B(net585),
    .Y(_0813_));
 sg13g2_nand2_1 _1435_ (.Y(_0814_),
    .A(\cic_b.integrator[1][5] ),
    .B(\cic_b.integrator[0][5] ));
 sg13g2_nor2b_1 _1436_ (.A(_0813_),
    .B_N(net586),
    .Y(_0815_));
 sg13g2_nand2_1 _1437_ (.Y(_0816_),
    .A(_0809_),
    .B(_0812_));
 sg13g2_xor2_1 _1438_ (.B(_0816_),
    .A(_0815_),
    .X(_0069_));
 sg13g2_nand2_1 _1439_ (.Y(_0817_),
    .A(\cic_b.integrator[1][6] ),
    .B(net549));
 sg13g2_nor2_1 _1440_ (.A(\cic_b.integrator[1][6] ),
    .B(net600),
    .Y(_0818_));
 sg13g2_xor2_1 _1441_ (.B(net549),
    .A(net238),
    .X(_0819_));
 sg13g2_nand3_1 _1442_ (.B(_0811_),
    .C(_0815_),
    .A(_0810_),
    .Y(_0820_));
 sg13g2_o21ai_1 _1443_ (.B1(_0814_),
    .Y(_0821_),
    .A1(_0809_),
    .A2(_0813_));
 sg13g2_nor2b_1 _1444_ (.A(_0821_),
    .B_N(_0820_),
    .Y(_0822_));
 sg13g2_xnor2_1 _1445_ (.Y(_0070_),
    .A(_0819_),
    .B(_0822_));
 sg13g2_nor2_1 _1446_ (.A(\cic_b.integrator[1][7] ),
    .B(\cic_b.integrator[0][7] ),
    .Y(_0823_));
 sg13g2_nand2_1 _1447_ (.Y(_0824_),
    .A(net306),
    .B(net587));
 sg13g2_nand2b_1 _1448_ (.Y(_0825_),
    .B(_0824_),
    .A_N(_0823_));
 sg13g2_o21ai_1 _1449_ (.B1(_0817_),
    .Y(_0826_),
    .A1(_0818_),
    .A2(_0822_));
 sg13g2_xnor2_1 _1450_ (.Y(_0071_),
    .A(_0825_),
    .B(net601));
 sg13g2_o21ai_1 _1451_ (.B1(_0824_),
    .Y(_0827_),
    .A1(_0817_),
    .A2(_0823_));
 sg13g2_nor2_1 _1452_ (.A(_0821_),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_a221oi_1 _1453_ (.B2(_0820_),
    .C1(_0823_),
    .B1(_0828_),
    .A1(_0818_),
    .Y(_0829_),
    .A2(_0824_));
 sg13g2_nand2_1 _1454_ (.Y(_0830_),
    .A(net471),
    .B(net575));
 sg13g2_xor2_1 _1455_ (.B(net575),
    .A(net471),
    .X(_0831_));
 sg13g2_inv_1 _1456_ (.Y(_0832_),
    .A(_0831_));
 sg13g2_nand2_1 _1457_ (.Y(_0833_),
    .A(_0829_),
    .B(_0831_));
 sg13g2_xnor2_1 _1458_ (.Y(_0072_),
    .A(_0829_),
    .B(_0832_));
 sg13g2_xnor2_1 _1459_ (.Y(_0834_),
    .A(net90),
    .B(net508));
 sg13g2_nand2_1 _1460_ (.Y(_0835_),
    .A(_0830_),
    .B(_0833_));
 sg13g2_xnor2_1 _1461_ (.Y(_0073_),
    .A(_0834_),
    .B(_0835_));
 sg13g2_nor2_1 _1462_ (.A(_0832_),
    .B(_0834_),
    .Y(_0836_));
 sg13g2_a21oi_1 _1463_ (.A1(_0718_),
    .A2(_0726_),
    .Y(_0837_),
    .B1(_0830_));
 sg13g2_a221oi_1 _1464_ (.B2(_0836_),
    .C1(_0837_),
    .B1(_0829_),
    .A1(\cic_b.integrator[1][9] ),
    .Y(_0838_),
    .A2(net512));
 sg13g2_nand2_1 _1465_ (.Y(_0839_),
    .A(net478),
    .B(net20));
 sg13g2_xnor2_1 _1466_ (.Y(_0840_),
    .A(net478),
    .B(net20));
 sg13g2_xor2_1 _1467_ (.B(_0840_),
    .A(_0838_),
    .X(_0062_));
 sg13g2_nor2_1 _1468_ (.A(\cic_b.integrator[1][11] ),
    .B(\cic_b.integrator[0][11] ),
    .Y(_0841_));
 sg13g2_xnor2_1 _1469_ (.Y(_0842_),
    .A(net518),
    .B(net113));
 sg13g2_o21ai_1 _1470_ (.B1(_0839_),
    .Y(_0843_),
    .A1(_0838_),
    .A2(_0840_));
 sg13g2_xnor2_1 _1471_ (.Y(_0063_),
    .A(_0842_),
    .B(_0843_));
 sg13g2_or2_1 _1472_ (.X(_0844_),
    .B(_0842_),
    .A(_0840_));
 sg13g2_nor2_1 _1473_ (.A(_0839_),
    .B(_0841_),
    .Y(_0845_));
 sg13g2_a21oi_1 _1474_ (.A1(net518),
    .A2(net113),
    .Y(_0846_),
    .B1(_0845_));
 sg13g2_o21ai_1 _1475_ (.B1(_0846_),
    .Y(_0847_),
    .A1(_0838_),
    .A2(_0844_));
 sg13g2_xnor2_1 _1476_ (.Y(_0848_),
    .A(\cic_b.integrator[1][12] ),
    .B(net557));
 sg13g2_xnor2_1 _1477_ (.Y(_0064_),
    .A(_0847_),
    .B(net558));
 sg13g2_xor2_1 _1478_ (.B(net525),
    .A(\cic_b.integrator[1][0] ),
    .X(_0061_));
 sg13g2_nand3_1 _1479_ (.B(\cic_a.integrator[0][1] ),
    .C(\cic_a.integrator[0][0] ),
    .A(net31),
    .Y(_0849_));
 sg13g2_a21o_1 _1480_ (.A2(net566),
    .A1(net31),
    .B1(net577),
    .X(_0850_));
 sg13g2_and2_1 _1481_ (.A(_0849_),
    .B(_0850_),
    .X(_0026_));
 sg13g2_nor2_2 _1482_ (.A(_0713_),
    .B(_0849_),
    .Y(_0851_));
 sg13g2_xnor2_1 _1483_ (.Y(_0027_),
    .A(net228),
    .B(_0849_));
 sg13g2_xor2_1 _1484_ (.B(_0851_),
    .A(net562),
    .X(_0028_));
 sg13g2_nand3_1 _1485_ (.B(net580),
    .C(_0851_),
    .A(net562),
    .Y(_0852_));
 sg13g2_a21o_1 _1486_ (.A2(_0851_),
    .A1(net562),
    .B1(net580),
    .X(_0853_));
 sg13g2_and2_1 _1487_ (.A(_0852_),
    .B(_0853_),
    .X(_0029_));
 sg13g2_nand4_1 _1488_ (.B(\cic_a.integrator[0][4] ),
    .C(net500),
    .A(\cic_a.integrator[0][3] ),
    .Y(_0854_),
    .D(_0851_));
 sg13g2_xnor2_1 _1489_ (.Y(_0030_),
    .A(net500),
    .B(_0852_));
 sg13g2_nor2_2 _1490_ (.A(_0714_),
    .B(_0854_),
    .Y(_0855_));
 sg13g2_xnor2_1 _1491_ (.Y(_0031_),
    .A(net552),
    .B(_0854_));
 sg13g2_xor2_1 _1492_ (.B(_0855_),
    .A(net534),
    .X(_0032_));
 sg13g2_nand3_1 _1493_ (.B(net582),
    .C(_0855_),
    .A(net534),
    .Y(_0856_));
 sg13g2_a21o_1 _1494_ (.A2(_0855_),
    .A1(net534),
    .B1(net582),
    .X(_0857_));
 sg13g2_and2_1 _1495_ (.A(_0856_),
    .B(_0857_),
    .X(_0033_));
 sg13g2_nor2_2 _1496_ (.A(_0715_),
    .B(_0856_),
    .Y(_0858_));
 sg13g2_xnor2_1 _1497_ (.Y(_0034_),
    .A(net542),
    .B(_0856_));
 sg13g2_xor2_1 _1498_ (.B(_0858_),
    .A(net545),
    .X(_0023_));
 sg13g2_nand3_1 _1499_ (.B(net584),
    .C(_0858_),
    .A(net545),
    .Y(_0859_));
 sg13g2_a21o_1 _1500_ (.A2(_0858_),
    .A1(net545),
    .B1(net584),
    .X(_0860_));
 sg13g2_and2_1 _1501_ (.A(_0859_),
    .B(_0860_),
    .X(_0024_));
 sg13g2_xnor2_1 _1502_ (.Y(_0025_),
    .A(net139),
    .B(_0859_));
 sg13g2_xor2_1 _1503_ (.B(\cic_a.integrator[0][0] ),
    .A(net31),
    .X(_0022_));
 sg13g2_nor2_2 _1504_ (.A(net3),
    .B(net411),
    .Y(_0861_));
 sg13g2_inv_1 _1505_ (.Y(_0862_),
    .A(_0861_));
 sg13g2_o21ai_1 _1506_ (.B1(net411),
    .Y(_0863_),
    .A1(net96),
    .A2(net105));
 sg13g2_nand4_1 _1507_ (.B(net161),
    .C(net55),
    .A(net412),
    .Y(_0864_),
    .D(_0863_));
 sg13g2_and2_1 _1508_ (.A(_0862_),
    .B(_0864_),
    .X(_0016_));
 sg13g2_nor2_2 _1509_ (.A(net3),
    .B(\serializer_b.sending ),
    .Y(_0865_));
 sg13g2_inv_1 _1510_ (.Y(_0866_),
    .A(_0865_));
 sg13g2_o21ai_1 _1511_ (.B1(net408),
    .Y(_0867_),
    .A1(\serializer_b.bit_cnt[0] ),
    .A2(net68));
 sg13g2_nand4_1 _1512_ (.B(net74),
    .C(net39),
    .A(net408),
    .Y(_0868_),
    .D(_0867_));
 sg13g2_and2_1 _1513_ (.A(net396),
    .B(_0868_),
    .X(_0020_));
 sg13g2_nor2_1 _1514_ (.A(net3),
    .B(net406),
    .Y(_0869_));
 sg13g2_or2_2 _1515_ (.X(_0870_),
    .B(net405),
    .A(net3));
 sg13g2_o21ai_1 _1516_ (.B1(net405),
    .Y(_0871_),
    .A1(net110),
    .A2(net166));
 sg13g2_nand4_1 _1517_ (.B(net51),
    .C(net46),
    .A(net405),
    .Y(_0872_),
    .D(_0871_));
 sg13g2_and2_1 _1518_ (.A(_0870_),
    .B(_0872_),
    .X(_0018_));
 sg13g2_xor2_1 _1519_ (.B(\cic_b.integrator[0][0] ),
    .A(net33),
    .X(_0048_));
 sg13g2_nand3_1 _1520_ (.B(\cic_b.integrator[0][1] ),
    .C(\cic_b.integrator[0][0] ),
    .A(net33),
    .Y(_0873_));
 sg13g2_a21o_1 _1521_ (.A2(net525),
    .A1(net33),
    .B1(net573),
    .X(_0874_));
 sg13g2_and2_1 _1522_ (.A(_0873_),
    .B(_0874_),
    .X(_0052_));
 sg13g2_nor2_2 _1523_ (.A(_0724_),
    .B(_0873_),
    .Y(_0875_));
 sg13g2_xnor2_1 _1524_ (.Y(_0053_),
    .A(net483),
    .B(_0873_));
 sg13g2_xor2_1 _1525_ (.B(_0875_),
    .A(net560),
    .X(_0054_));
 sg13g2_nand3_1 _1526_ (.B(net583),
    .C(_0875_),
    .A(net560),
    .Y(_0876_));
 sg13g2_a21o_1 _1527_ (.A2(_0875_),
    .A1(net560),
    .B1(net583),
    .X(_0877_));
 sg13g2_and2_1 _1528_ (.A(_0876_),
    .B(_0877_),
    .X(_0055_));
 sg13g2_nand4_1 _1529_ (.B(\cic_b.integrator[0][4] ),
    .C(net520),
    .A(\cic_b.integrator[0][3] ),
    .Y(_0878_),
    .D(_0875_));
 sg13g2_xnor2_1 _1530_ (.Y(_0056_),
    .A(net520),
    .B(_0876_));
 sg13g2_nor2_2 _1531_ (.A(_0725_),
    .B(_0878_),
    .Y(_0879_));
 sg13g2_xnor2_1 _1532_ (.Y(_0057_),
    .A(net549),
    .B(_0878_));
 sg13g2_xor2_1 _1533_ (.B(_0879_),
    .A(net536),
    .X(_0058_));
 sg13g2_nand3_1 _1534_ (.B(net575),
    .C(_0879_),
    .A(\cic_b.integrator[0][7] ),
    .Y(_0880_));
 sg13g2_a21o_1 _1535_ (.A2(_0879_),
    .A1(net536),
    .B1(net575),
    .X(_0881_));
 sg13g2_and2_1 _1536_ (.A(_0880_),
    .B(_0881_),
    .X(_0059_));
 sg13g2_nor2_2 _1537_ (.A(_0726_),
    .B(_0880_),
    .Y(_0882_));
 sg13g2_xnor2_1 _1538_ (.Y(_0060_),
    .A(net508),
    .B(_0880_));
 sg13g2_xor2_1 _1539_ (.B(_0882_),
    .A(net20),
    .X(_0049_));
 sg13g2_nand3_1 _1540_ (.B(\cic_b.integrator[0][11] ),
    .C(_0882_),
    .A(net20),
    .Y(_0883_));
 sg13g2_a21o_1 _1541_ (.A2(_0882_),
    .A1(net20),
    .B1(net113),
    .X(_0884_));
 sg13g2_and2_1 _1542_ (.A(net21),
    .B(_0884_),
    .X(_0050_));
 sg13g2_xnor2_1 _1543_ (.Y(_0051_),
    .A(\cic_b.integrator[0][12] ),
    .B(net21));
 sg13g2_and2_2 _1544_ (.A(_0734_),
    .B(_0735_),
    .X(_0885_));
 sg13g2_nand2_1 _1545_ (.Y(_0886_),
    .A(_0734_),
    .B(_0735_));
 sg13g2_mux2_1 _1546_ (.A0(net255),
    .A1(\cic_a.temp_delay[0][0] ),
    .S(net392),
    .X(_0078_));
 sg13g2_mux2_1 _1547_ (.A0(\cic_a.delay[0][1] ),
    .A1(net203),
    .S(net395),
    .X(_0079_));
 sg13g2_mux2_1 _1548_ (.A0(net337),
    .A1(net285),
    .S(net388),
    .X(_0080_));
 sg13g2_mux2_1 _1549_ (.A0(\cic_a.delay[0][3] ),
    .A1(net242),
    .S(net388),
    .X(_0081_));
 sg13g2_mux2_1 _1550_ (.A0(net470),
    .A1(net329),
    .S(net386),
    .X(_0082_));
 sg13g2_nor2_1 _1551_ (.A(net66),
    .B(net376),
    .Y(_0887_));
 sg13g2_a21oi_1 _1552_ (.A1(_0727_),
    .A2(net376),
    .Y(_0083_),
    .B1(_0887_));
 sg13g2_mux2_1 _1553_ (.A0(\cic_a.delay[0][6] ),
    .A1(net196),
    .S(net386),
    .X(_0084_));
 sg13g2_mux2_1 _1554_ (.A0(\cic_a.delay[0][7] ),
    .A1(net173),
    .S(net386),
    .X(_0085_));
 sg13g2_mux2_1 _1555_ (.A0(net175),
    .A1(\cic_a.temp_delay[0][8] ),
    .S(net385),
    .X(_0086_));
 sg13g2_mux2_1 _1556_ (.A0(net287),
    .A1(net92),
    .S(net385),
    .X(_0087_));
 sg13g2_mux2_1 _1557_ (.A0(net332),
    .A1(net313),
    .S(net383),
    .X(_0088_));
 sg13g2_mux2_1 _1558_ (.A0(net335),
    .A1(net244),
    .S(net383),
    .X(_0089_));
 sg13g2_mux2_1 _1559_ (.A0(net169),
    .A1(\cic_a.temp_delay[0][12] ),
    .S(net383),
    .X(_0090_));
 sg13g2_nand2b_2 _1560_ (.Y(_0888_),
    .B(net255),
    .A_N(\cic_a.integrator[1][0] ));
 sg13g2_nand2b_1 _1561_ (.Y(_0889_),
    .B(net514),
    .A_N(net522));
 sg13g2_a21oi_2 _1562_ (.B1(net382),
    .Y(_0890_),
    .A2(_0889_),
    .A1(_0888_));
 sg13g2_a21o_1 _1563_ (.A2(net381),
    .A1(net502),
    .B1(_0890_),
    .X(_0091_));
 sg13g2_nor2_1 _1564_ (.A(net527),
    .B(net394),
    .Y(_0891_));
 sg13g2_nor2b_1 _1565_ (.A(\cic_a.delay[0][1] ),
    .B_N(\cic_a.integrator[1][1] ),
    .Y(_0892_));
 sg13g2_xnor2_1 _1566_ (.Y(_0893_),
    .A(\cic_a.integrator[1][1] ),
    .B(\cic_a.delay[0][1] ));
 sg13g2_xnor2_1 _1567_ (.Y(_0894_),
    .A(_0888_),
    .B(_0893_));
 sg13g2_a21oi_1 _1568_ (.A1(net392),
    .A2(_0894_),
    .Y(_0092_),
    .B1(_0891_));
 sg13g2_nor2_1 _1569_ (.A(net554),
    .B(net392),
    .Y(_0895_));
 sg13g2_nand2b_1 _1570_ (.Y(_0896_),
    .B(\cic_a.integrator[1][2] ),
    .A_N(\cic_a.delay[0][2] ));
 sg13g2_xor2_1 _1571_ (.B(\cic_a.delay[0][2] ),
    .A(\cic_a.integrator[1][2] ),
    .X(_0897_));
 sg13g2_a21oi_2 _1572_ (.B1(_0892_),
    .Y(_0898_),
    .A2(_0893_),
    .A1(_0888_));
 sg13g2_xnor2_1 _1573_ (.Y(_0899_),
    .A(_0897_),
    .B(_0898_));
 sg13g2_a21oi_1 _1574_ (.A1(net392),
    .A2(_0899_),
    .Y(_0093_),
    .B1(_0895_));
 sg13g2_nor2_1 _1575_ (.A(net538),
    .B(net392),
    .Y(_0900_));
 sg13g2_nor2b_1 _1576_ (.A(\cic_a.delay[0][3] ),
    .B_N(\cic_a.integrator[1][3] ),
    .Y(_0901_));
 sg13g2_nand2b_1 _1577_ (.Y(_0902_),
    .B(\cic_a.delay[0][3] ),
    .A_N(\cic_a.integrator[1][3] ));
 sg13g2_nor2b_1 _1578_ (.A(_0901_),
    .B_N(_0902_),
    .Y(_0903_));
 sg13g2_o21ai_1 _1579_ (.B1(_0896_),
    .Y(_0904_),
    .A1(_0897_),
    .A2(_0898_));
 sg13g2_xnor2_1 _1580_ (.Y(_0905_),
    .A(_0903_),
    .B(_0904_));
 sg13g2_a21oi_1 _1581_ (.A1(net392),
    .A2(_0905_),
    .Y(_0094_),
    .B1(_0900_));
 sg13g2_nand2_1 _1582_ (.Y(_0906_),
    .A(net505),
    .B(net378));
 sg13g2_a21oi_2 _1583_ (.B1(_0901_),
    .Y(_0907_),
    .A2(_0904_),
    .A1(_0902_));
 sg13g2_nor2b_1 _1584_ (.A(\cic_a.delay[0][4] ),
    .B_N(\cic_a.integrator[1][4] ),
    .Y(_0908_));
 sg13g2_xor2_1 _1585_ (.B(\cic_a.delay[0][4] ),
    .A(\cic_a.integrator[1][4] ),
    .X(_0909_));
 sg13g2_nor2_1 _1586_ (.A(_0907_),
    .B(_0909_),
    .Y(_0910_));
 sg13g2_a21o_1 _1587_ (.A2(_0909_),
    .A1(_0907_),
    .B1(net378),
    .X(_0911_));
 sg13g2_o21ai_1 _1588_ (.B1(_0906_),
    .Y(_0095_),
    .A1(_0910_),
    .A2(_0911_));
 sg13g2_nand2_1 _1589_ (.Y(_0912_),
    .A(net530),
    .B(net378));
 sg13g2_nor2_1 _1590_ (.A(\cic_a.integrator[1][5] ),
    .B(_0727_),
    .Y(_0913_));
 sg13g2_xor2_1 _1591_ (.B(\cic_a.delay[0][5] ),
    .A(\cic_a.integrator[1][5] ),
    .X(_0914_));
 sg13g2_nor2_1 _1592_ (.A(_0908_),
    .B(_0910_),
    .Y(_0915_));
 sg13g2_xnor2_1 _1593_ (.Y(_0916_),
    .A(_0914_),
    .B(_0915_));
 sg13g2_o21ai_1 _1594_ (.B1(_0912_),
    .Y(_0096_),
    .A1(net378),
    .A2(_0916_));
 sg13g2_nor2_1 _1595_ (.A(net546),
    .B(net388),
    .Y(_0917_));
 sg13g2_nor2b_1 _1596_ (.A(\cic_a.delay[0][6] ),
    .B_N(\cic_a.integrator[1][6] ),
    .Y(_0918_));
 sg13g2_xnor2_1 _1597_ (.Y(_0919_),
    .A(\cic_a.integrator[1][6] ),
    .B(\cic_a.delay[0][6] ));
 sg13g2_a21oi_1 _1598_ (.A1(\cic_a.integrator[1][5] ),
    .A2(_0727_),
    .Y(_0920_),
    .B1(_0908_));
 sg13g2_o21ai_1 _1599_ (.B1(_0920_),
    .Y(_0921_),
    .A1(_0907_),
    .A2(_0909_));
 sg13g2_nor2b_1 _1600_ (.A(_0913_),
    .B_N(_0921_),
    .Y(_0922_));
 sg13g2_xnor2_1 _1601_ (.Y(_0923_),
    .A(_0919_),
    .B(_0922_));
 sg13g2_a21oi_1 _1602_ (.A1(net386),
    .A2(_0923_),
    .Y(_0097_),
    .B1(_0917_));
 sg13g2_nor2b_1 _1603_ (.A(\cic_a.delay[0][7] ),
    .B_N(\cic_a.integrator[1][7] ),
    .Y(_0924_));
 sg13g2_nand2b_1 _1604_ (.Y(_0925_),
    .B(\cic_a.delay[0][7] ),
    .A_N(\cic_a.integrator[1][7] ));
 sg13g2_nor2b_1 _1605_ (.A(_0924_),
    .B_N(_0925_),
    .Y(_0926_));
 sg13g2_a21oi_1 _1606_ (.A1(_0919_),
    .A2(_0922_),
    .Y(_0927_),
    .B1(_0918_));
 sg13g2_xnor2_1 _1607_ (.Y(_0928_),
    .A(_0926_),
    .B(_0927_));
 sg13g2_mux2_1 _1608_ (.A0(net519),
    .A1(_0928_),
    .S(net386),
    .X(_0098_));
 sg13g2_nor2_1 _1609_ (.A(net539),
    .B(net385),
    .Y(_0929_));
 sg13g2_nand3b_1 _1610_ (.B(_0925_),
    .C(_0919_),
    .Y(_0930_),
    .A_N(_0924_));
 sg13g2_or3_1 _1611_ (.A(_0909_),
    .B(_0914_),
    .C(_0930_),
    .X(_0931_));
 sg13g2_a21oi_1 _1612_ (.A1(_0918_),
    .A2(_0925_),
    .Y(_0932_),
    .B1(_0924_));
 sg13g2_or3_1 _1613_ (.A(_0913_),
    .B(_0920_),
    .C(_0930_),
    .X(_0933_));
 sg13g2_and2_1 _1614_ (.A(_0932_),
    .B(_0933_),
    .X(_0934_));
 sg13g2_o21ai_1 _1615_ (.B1(_0934_),
    .Y(_0935_),
    .A1(_0907_),
    .A2(_0931_));
 sg13g2_nor2b_1 _1616_ (.A(\cic_a.delay[0][8] ),
    .B_N(\cic_a.integrator[1][8] ),
    .Y(_0936_));
 sg13g2_nor2b_1 _1617_ (.A(\cic_a.integrator[1][8] ),
    .B_N(\cic_a.delay[0][8] ),
    .Y(_0937_));
 sg13g2_nor2_1 _1618_ (.A(_0936_),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_xnor2_1 _1619_ (.Y(_0939_),
    .A(_0935_),
    .B(_0938_));
 sg13g2_a21oi_1 _1620_ (.A1(net384),
    .A2(_0939_),
    .Y(_0099_),
    .B1(_0929_));
 sg13g2_nor2_1 _1621_ (.A(net551),
    .B(net384),
    .Y(_0940_));
 sg13g2_nor2_1 _1622_ (.A(_0716_),
    .B(\cic_a.delay[0][9] ),
    .Y(_0941_));
 sg13g2_nand2_1 _1623_ (.Y(_0942_),
    .A(_0716_),
    .B(\cic_a.delay[0][9] ));
 sg13g2_nand2b_1 _1624_ (.Y(_0943_),
    .B(_0942_),
    .A_N(_0941_));
 sg13g2_a21oi_1 _1625_ (.A1(_0935_),
    .A2(_0938_),
    .Y(_0944_),
    .B1(_0936_));
 sg13g2_xnor2_1 _1626_ (.Y(_0945_),
    .A(_0943_),
    .B(_0944_));
 sg13g2_a21oi_1 _1627_ (.A1(net384),
    .A2(_0945_),
    .Y(_0100_),
    .B1(_0940_));
 sg13g2_nor2b_1 _1628_ (.A(\cic_a.delay[0][10] ),
    .B_N(\cic_a.integrator[1][10] ),
    .Y(_0946_));
 sg13g2_xnor2_1 _1629_ (.Y(_0947_),
    .A(\cic_a.integrator[1][10] ),
    .B(\cic_a.delay[0][10] ));
 sg13g2_inv_1 _1630_ (.Y(_0948_),
    .A(_0947_));
 sg13g2_a21o_1 _1631_ (.A2(_0942_),
    .A1(_0936_),
    .B1(_0941_),
    .X(_0949_));
 sg13g2_nor3_1 _1632_ (.A(_0936_),
    .B(_0937_),
    .C(_0943_),
    .Y(_0950_));
 sg13g2_a21o_1 _1633_ (.A2(_0950_),
    .A1(_0935_),
    .B1(_0949_),
    .X(_0951_));
 sg13g2_o21ai_1 _1634_ (.B1(net383),
    .Y(_0952_),
    .A1(_0947_),
    .A2(_0951_));
 sg13g2_a21oi_1 _1635_ (.A1(_0947_),
    .A2(_0951_),
    .Y(_0953_),
    .B1(_0952_));
 sg13g2_a21o_1 _1636_ (.A2(net375),
    .A1(net516),
    .B1(_0953_),
    .X(_0101_));
 sg13g2_nor2_1 _1637_ (.A(net476),
    .B(net384),
    .Y(_0954_));
 sg13g2_nor2b_1 _1638_ (.A(\cic_a.delay[0][11] ),
    .B_N(\cic_a.integrator[1][11] ),
    .Y(_0955_));
 sg13g2_nand2b_1 _1639_ (.Y(_0956_),
    .B(\cic_a.delay[0][11] ),
    .A_N(\cic_a.integrator[1][11] ));
 sg13g2_nand2b_1 _1640_ (.Y(_0957_),
    .B(_0956_),
    .A_N(_0955_));
 sg13g2_a21oi_1 _1641_ (.A1(_0947_),
    .A2(_0951_),
    .Y(_0958_),
    .B1(_0946_));
 sg13g2_xnor2_1 _1642_ (.Y(_0959_),
    .A(_0957_),
    .B(_0958_));
 sg13g2_a21oi_1 _1643_ (.A1(net384),
    .A2(_0959_),
    .Y(_0102_),
    .B1(_0954_));
 sg13g2_nor2_1 _1644_ (.A(net198),
    .B(net383),
    .Y(_0960_));
 sg13g2_nor2_1 _1645_ (.A(_0948_),
    .B(_0957_),
    .Y(_0961_));
 sg13g2_a221oi_1 _1646_ (.B2(_0951_),
    .C1(_0955_),
    .B1(_0961_),
    .A1(_0946_),
    .Y(_0962_),
    .A2(_0956_));
 sg13g2_xor2_1 _1647_ (.B(net169),
    .A(\cic_a.integrator[1][12] ),
    .X(_0311_));
 sg13g2_xnor2_1 _1648_ (.Y(_0312_),
    .A(_0962_),
    .B(_0311_));
 sg13g2_a21oi_1 _1649_ (.A1(net383),
    .A2(_0312_),
    .Y(_0103_),
    .B1(_0960_));
 sg13g2_mux2_1 _1650_ (.A0(net241),
    .A1(net99),
    .S(net393),
    .X(_0104_));
 sg13g2_mux2_1 _1651_ (.A0(net331),
    .A1(net194),
    .S(net393),
    .X(_0105_));
 sg13g2_mux2_1 _1652_ (.A0(net129),
    .A1(net109),
    .S(net393),
    .X(_0106_));
 sg13g2_mux2_1 _1653_ (.A0(net289),
    .A1(net162),
    .S(net393),
    .X(_0107_));
 sg13g2_nor2_1 _1654_ (.A(net126),
    .B(net381),
    .Y(_0313_));
 sg13g2_a21oi_1 _1655_ (.A1(_0693_),
    .A2(net381),
    .Y(_0108_),
    .B1(_0313_));
 sg13g2_mux2_1 _1656_ (.A0(net345),
    .A1(net61),
    .S(net391),
    .X(_0109_));
 sg13g2_mux2_1 _1657_ (.A0(net477),
    .A1(net128),
    .S(net390),
    .X(_0110_));
 sg13g2_nor2_1 _1658_ (.A(net148),
    .B(net380),
    .Y(_0314_));
 sg13g2_a21oi_1 _1659_ (.A1(_0695_),
    .A2(net381),
    .Y(_0111_),
    .B1(_0314_));
 sg13g2_mux2_1 _1660_ (.A0(net141),
    .A1(net517),
    .S(net390),
    .X(_0112_));
 sg13g2_mux2_1 _1661_ (.A0(net317),
    .A1(net59),
    .S(net390),
    .X(_0113_));
 sg13g2_mux2_1 _1662_ (.A0(net273),
    .A1(net191),
    .S(net388),
    .X(_0114_));
 sg13g2_mux2_1 _1663_ (.A0(net252),
    .A1(net60),
    .S(net390),
    .X(_0115_));
 sg13g2_mux2_1 _1664_ (.A0(net301),
    .A1(net103),
    .S(net387),
    .X(_0116_));
 sg13g2_mux2_1 _1665_ (.A0(\cic_a.delay[1][0] ),
    .A1(net291),
    .S(net393),
    .X(_0117_));
 sg13g2_mux2_1 _1666_ (.A0(net472),
    .A1(net257),
    .S(net394),
    .X(_0118_));
 sg13g2_mux2_1 _1667_ (.A0(net473),
    .A1(net259),
    .S(net394),
    .X(_0119_));
 sg13g2_mux2_1 _1668_ (.A0(net299),
    .A1(net234),
    .S(net392),
    .X(_0120_));
 sg13g2_mux2_1 _1669_ (.A0(net288),
    .A1(net263),
    .S(net389),
    .X(_0121_));
 sg13g2_mux2_1 _1670_ (.A0(net278),
    .A1(net267),
    .S(net389),
    .X(_0122_));
 sg13g2_mux2_1 _1671_ (.A0(net324),
    .A1(net303),
    .S(net387),
    .X(_0123_));
 sg13g2_mux2_1 _1672_ (.A0(net157),
    .A1(\cic_a.temp_delay[1][7] ),
    .S(net388),
    .X(_0124_));
 sg13g2_mux2_1 _1673_ (.A0(net265),
    .A1(\cic_a.temp_delay[1][8] ),
    .S(net387),
    .X(_0125_));
 sg13g2_nor2_1 _1674_ (.A(net85),
    .B(net377),
    .Y(_0315_));
 sg13g2_a21oi_1 _1675_ (.A1(_0712_),
    .A2(net377),
    .Y(_0126_),
    .B1(_0315_));
 sg13g2_mux2_1 _1676_ (.A0(net215),
    .A1(\cic_a.temp_delay[1][10] ),
    .S(net384),
    .X(_0127_));
 sg13g2_mux2_1 _1677_ (.A0(net319),
    .A1(\cic_a.temp_delay[1][11] ),
    .S(net384),
    .X(_0128_));
 sg13g2_mux2_1 _1678_ (.A0(net236),
    .A1(\cic_a.temp_delay[1][12] ),
    .S(net384),
    .X(_0129_));
 sg13g2_nor2_1 _1679_ (.A(net99),
    .B(net395),
    .Y(_0316_));
 sg13g2_nor2b_1 _1680_ (.A(\cic_a.temp_comb[0][0] ),
    .B_N(\cic_a.delay[1][0] ),
    .Y(_0317_));
 sg13g2_xnor2_1 _1681_ (.Y(_0318_),
    .A(\cic_a.temp_comb[0][0] ),
    .B(\cic_a.delay[1][0] ));
 sg13g2_a21oi_1 _1682_ (.A1(net393),
    .A2(_0318_),
    .Y(_0130_),
    .B1(_0316_));
 sg13g2_nor2_1 _1683_ (.A(net194),
    .B(net393),
    .Y(_0319_));
 sg13g2_nand2b_1 _1684_ (.Y(_0320_),
    .B(\cic_a.temp_comb[0][1] ),
    .A_N(\cic_a.delay[1][1] ));
 sg13g2_xor2_1 _1685_ (.B(\cic_a.delay[1][1] ),
    .A(\cic_a.temp_comb[0][1] ),
    .X(_0321_));
 sg13g2_xnor2_1 _1686_ (.Y(_0322_),
    .A(_0317_),
    .B(_0321_));
 sg13g2_a21oi_1 _1687_ (.A1(net394),
    .A2(_0322_),
    .Y(_0131_),
    .B1(_0319_));
 sg13g2_nor2_1 _1688_ (.A(net109),
    .B(net393),
    .Y(_0323_));
 sg13g2_nor2b_1 _1689_ (.A(\cic_a.delay[1][2] ),
    .B_N(\cic_a.temp_comb[0][2] ),
    .Y(_0324_));
 sg13g2_xnor2_1 _1690_ (.Y(_0325_),
    .A(\cic_a.temp_comb[0][2] ),
    .B(\cic_a.delay[1][2] ));
 sg13g2_o21ai_1 _1691_ (.B1(_0320_),
    .Y(_0326_),
    .A1(_0317_),
    .A2(_0321_));
 sg13g2_xnor2_1 _1692_ (.Y(_0327_),
    .A(_0325_),
    .B(_0326_));
 sg13g2_a21oi_1 _1693_ (.A1(net394),
    .A2(_0327_),
    .Y(_0132_),
    .B1(_0323_));
 sg13g2_nor2_1 _1694_ (.A(net162),
    .B(net394),
    .Y(_0328_));
 sg13g2_nand2b_1 _1695_ (.Y(_0329_),
    .B(\cic_a.temp_comb[0][3] ),
    .A_N(\cic_a.delay[1][3] ));
 sg13g2_xor2_1 _1696_ (.B(\cic_a.delay[1][3] ),
    .A(\cic_a.temp_comb[0][3] ),
    .X(_0330_));
 sg13g2_a21oi_2 _1697_ (.B1(_0324_),
    .Y(_0331_),
    .A2(_0326_),
    .A1(_0325_));
 sg13g2_xnor2_1 _1698_ (.Y(_0332_),
    .A(_0330_),
    .B(_0331_));
 sg13g2_a21oi_1 _1699_ (.A1(net394),
    .A2(_0332_),
    .Y(_0133_),
    .B1(_0328_));
 sg13g2_nor2_1 _1700_ (.A(net126),
    .B(net390),
    .Y(_0333_));
 sg13g2_o21ai_1 _1701_ (.B1(_0329_),
    .Y(_0334_),
    .A1(_0330_),
    .A2(_0331_));
 sg13g2_nor2b_1 _1702_ (.A(\cic_a.delay[1][4] ),
    .B_N(\cic_a.temp_comb[0][4] ),
    .Y(_0335_));
 sg13g2_xnor2_1 _1703_ (.Y(_0336_),
    .A(\cic_a.temp_comb[0][4] ),
    .B(\cic_a.delay[1][4] ));
 sg13g2_xnor2_1 _1704_ (.Y(_0337_),
    .A(_0334_),
    .B(_0336_));
 sg13g2_a21oi_1 _1705_ (.A1(net390),
    .A2(_0337_),
    .Y(_0134_),
    .B1(_0333_));
 sg13g2_nand2b_1 _1706_ (.Y(_0338_),
    .B(\cic_a.delay[1][5] ),
    .A_N(\cic_a.temp_comb[0][5] ));
 sg13g2_nor2b_1 _1707_ (.A(\cic_a.delay[1][5] ),
    .B_N(\cic_a.temp_comb[0][5] ),
    .Y(_0339_));
 sg13g2_xor2_1 _1708_ (.B(net611),
    .A(\cic_a.temp_comb[0][5] ),
    .X(_0340_));
 sg13g2_a21oi_1 _1709_ (.A1(_0334_),
    .A2(_0336_),
    .Y(_0341_),
    .B1(_0335_));
 sg13g2_xnor2_1 _1710_ (.Y(_0342_),
    .A(_0340_),
    .B(_0341_));
 sg13g2_nand2_1 _1711_ (.Y(_0343_),
    .A(net61),
    .B(net380));
 sg13g2_o21ai_1 _1712_ (.B1(_0343_),
    .Y(_0135_),
    .A1(net380),
    .A2(_0342_));
 sg13g2_nor2_1 _1713_ (.A(net128),
    .B(net390),
    .Y(_0344_));
 sg13g2_nand2b_1 _1714_ (.Y(_0345_),
    .B(\cic_a.temp_comb[0][6] ),
    .A_N(\cic_a.delay[1][6] ));
 sg13g2_xor2_1 _1715_ (.B(\cic_a.delay[1][6] ),
    .A(\cic_a.temp_comb[0][6] ),
    .X(_0346_));
 sg13g2_nand3b_1 _1716_ (.B(_0336_),
    .C(_0338_),
    .Y(_0347_),
    .A_N(_0339_));
 sg13g2_inv_1 _1717_ (.Y(_0348_),
    .A(_0347_));
 sg13g2_a21o_1 _1718_ (.A2(_0338_),
    .A1(_0335_),
    .B1(_0339_),
    .X(_0349_));
 sg13g2_a21oi_1 _1719_ (.A1(_0334_),
    .A2(_0348_),
    .Y(_0350_),
    .B1(_0349_));
 sg13g2_xnor2_1 _1720_ (.Y(_0351_),
    .A(_0346_),
    .B(_0350_));
 sg13g2_a21oi_1 _1721_ (.A1(net391),
    .A2(_0351_),
    .Y(_0136_),
    .B1(_0344_));
 sg13g2_nor2_1 _1722_ (.A(net148),
    .B(net391),
    .Y(_0352_));
 sg13g2_nor2b_1 _1723_ (.A(\cic_a.temp_comb[0][7] ),
    .B_N(\cic_a.delay[1][7] ),
    .Y(_0353_));
 sg13g2_nand2b_1 _1724_ (.Y(_0354_),
    .B(\cic_a.temp_comb[0][7] ),
    .A_N(\cic_a.delay[1][7] ));
 sg13g2_nand2b_1 _1725_ (.Y(_0355_),
    .B(_0354_),
    .A_N(_0353_));
 sg13g2_o21ai_1 _1726_ (.B1(_0345_),
    .Y(_0356_),
    .A1(_0346_),
    .A2(_0350_));
 sg13g2_xor2_1 _1727_ (.B(_0356_),
    .A(_0355_),
    .X(_0357_));
 sg13g2_a21oi_1 _1728_ (.A1(net390),
    .A2(_0357_),
    .Y(_0137_),
    .B1(_0352_));
 sg13g2_nor2_1 _1729_ (.A(net517),
    .B(net388),
    .Y(_0358_));
 sg13g2_nand2b_1 _1730_ (.Y(_0359_),
    .B(\cic_a.temp_comb[0][8] ),
    .A_N(\cic_a.delay[1][8] ));
 sg13g2_xor2_1 _1731_ (.B(\cic_a.delay[1][8] ),
    .A(\cic_a.temp_comb[0][8] ),
    .X(_0360_));
 sg13g2_o21ai_1 _1732_ (.B1(_0354_),
    .Y(_0361_),
    .A1(_0345_),
    .A2(_0353_));
 sg13g2_nor2_1 _1733_ (.A(_0346_),
    .B(_0355_),
    .Y(_0362_));
 sg13g2_nor3_1 _1734_ (.A(_0346_),
    .B(_0347_),
    .C(_0355_),
    .Y(_0363_));
 sg13g2_a221oi_1 _1735_ (.B2(_0334_),
    .C1(_0361_),
    .B1(_0363_),
    .A1(_0349_),
    .Y(_0364_),
    .A2(_0362_));
 sg13g2_xnor2_1 _1736_ (.Y(_0365_),
    .A(_0360_),
    .B(_0364_));
 sg13g2_a21oi_1 _1737_ (.A1(net388),
    .A2(_0365_),
    .Y(_0138_),
    .B1(_0358_));
 sg13g2_xnor2_1 _1738_ (.Y(_0366_),
    .A(\cic_a.temp_comb[0][9] ),
    .B(net613));
 sg13g2_o21ai_1 _1739_ (.B1(_0359_),
    .Y(_0367_),
    .A1(_0360_),
    .A2(_0364_));
 sg13g2_xnor2_1 _1740_ (.Y(_0368_),
    .A(_0366_),
    .B(_0367_));
 sg13g2_nand2_1 _1741_ (.Y(_0369_),
    .A(net59),
    .B(net380));
 sg13g2_o21ai_1 _1742_ (.B1(_0369_),
    .Y(_0139_),
    .A1(net380),
    .A2(_0368_));
 sg13g2_nand2b_1 _1743_ (.Y(_0370_),
    .B(_0366_),
    .A_N(_0360_));
 sg13g2_a21oi_1 _1744_ (.A1(_0711_),
    .A2(\cic_a.delay[1][9] ),
    .Y(_0371_),
    .B1(_0359_));
 sg13g2_a21oi_1 _1745_ (.A1(\cic_a.temp_comb[0][9] ),
    .A2(_0712_),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_o21ai_1 _1746_ (.B1(_0372_),
    .Y(_0373_),
    .A1(_0364_),
    .A2(_0370_));
 sg13g2_nor2b_1 _1747_ (.A(\cic_a.delay[1][10] ),
    .B_N(\cic_a.temp_comb[0][10] ),
    .Y(_0374_));
 sg13g2_nor2b_1 _1748_ (.A(\cic_a.temp_comb[0][10] ),
    .B_N(\cic_a.delay[1][10] ),
    .Y(_0375_));
 sg13g2_nor2_1 _1749_ (.A(_0374_),
    .B(_0375_),
    .Y(_0376_));
 sg13g2_o21ai_1 _1750_ (.B1(net387),
    .Y(_0377_),
    .A1(_0373_),
    .A2(_0376_));
 sg13g2_a21oi_1 _1751_ (.A1(_0373_),
    .A2(_0376_),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_a21o_1 _1752_ (.A2(net377),
    .A1(net191),
    .B1(_0378_),
    .X(_0140_));
 sg13g2_nor2b_1 _1753_ (.A(\cic_a.delay[1][11] ),
    .B_N(\cic_a.temp_comb[0][11] ),
    .Y(_0379_));
 sg13g2_nand2b_1 _1754_ (.Y(_0380_),
    .B(\cic_a.delay[1][11] ),
    .A_N(\cic_a.temp_comb[0][11] ));
 sg13g2_nand2b_1 _1755_ (.Y(_0381_),
    .B(_0380_),
    .A_N(_0379_));
 sg13g2_a21oi_1 _1756_ (.A1(_0373_),
    .A2(_0376_),
    .Y(_0382_),
    .B1(_0374_));
 sg13g2_xnor2_1 _1757_ (.Y(_0383_),
    .A(_0381_),
    .B(_0382_));
 sg13g2_nand2_1 _1758_ (.Y(_0384_),
    .A(net60),
    .B(net380));
 sg13g2_o21ai_1 _1759_ (.B1(_0384_),
    .Y(_0141_),
    .A1(net377),
    .A2(_0383_));
 sg13g2_nor2_1 _1760_ (.A(net103),
    .B(net387),
    .Y(_0385_));
 sg13g2_nor3_1 _1761_ (.A(_0374_),
    .B(_0375_),
    .C(_0381_),
    .Y(_0386_));
 sg13g2_a221oi_1 _1762_ (.B2(_0373_),
    .C1(_0379_),
    .B1(_0386_),
    .A1(_0374_),
    .Y(_0387_),
    .A2(_0380_));
 sg13g2_xor2_1 _1763_ (.B(\cic_a.delay[1][12] ),
    .A(\cic_a.temp_comb[0][12] ),
    .X(_0388_));
 sg13g2_xnor2_1 _1764_ (.Y(_0389_),
    .A(_0387_),
    .B(_0388_));
 sg13g2_a21oi_1 _1765_ (.A1(net387),
    .A2(_0389_),
    .Y(_0142_),
    .B1(_0385_));
 sg13g2_mux2_1 _1766_ (.A0(\cic_a.integrator[1][0] ),
    .A1(net271),
    .S(net381),
    .X(_0143_));
 sg13g2_mux2_1 _1767_ (.A0(net282),
    .A1(net203),
    .S(net380),
    .X(_0144_));
 sg13g2_mux2_1 _1768_ (.A0(\cic_a.integrator[1][2] ),
    .A1(net285),
    .S(net382),
    .X(_0145_));
 sg13g2_mux2_1 _1769_ (.A0(net300),
    .A1(net242),
    .S(net378),
    .X(_0146_));
 sg13g2_mux2_1 _1770_ (.A0(\cic_a.integrator[1][4] ),
    .A1(net329),
    .S(net375),
    .X(_0147_));
 sg13g2_mux2_1 _1771_ (.A0(net491),
    .A1(net66),
    .S(net375),
    .X(_0148_));
 sg13g2_mux2_1 _1772_ (.A0(net328),
    .A1(net196),
    .S(net376),
    .X(_0149_));
 sg13g2_mux2_1 _1773_ (.A0(net336),
    .A1(net173),
    .S(net376),
    .X(_0150_));
 sg13g2_mux2_1 _1774_ (.A0(\cic_a.integrator[1][8] ),
    .A1(net468),
    .S(net375),
    .X(_0151_));
 sg13g2_nor2_1 _1775_ (.A(net92),
    .B(net383),
    .Y(_0390_));
 sg13g2_a21oi_1 _1776_ (.A1(_0716_),
    .A2(net383),
    .Y(_0152_),
    .B1(_0390_));
 sg13g2_mux2_1 _1777_ (.A0(\cic_a.integrator[1][10] ),
    .A1(net313),
    .S(net375),
    .X(_0153_));
 sg13g2_mux2_1 _1778_ (.A0(\cic_a.integrator[1][11] ),
    .A1(net244),
    .S(net375),
    .X(_0154_));
 sg13g2_mux2_1 _1779_ (.A0(\cic_a.integrator[1][12] ),
    .A1(net481),
    .S(net375),
    .X(_0155_));
 sg13g2_and2_1 _1780_ (.A(_0742_),
    .B(_0743_),
    .X(_0391_));
 sg13g2_nand2_1 _1781_ (.Y(_0392_),
    .A(_0742_),
    .B(_0743_));
 sg13g2_mux2_1 _1782_ (.A0(net205),
    .A1(\cic_b.temp_delay[0][0] ),
    .S(net373),
    .X(_0156_));
 sg13g2_mux2_1 _1783_ (.A0(net315),
    .A1(\cic_b.temp_delay[0][1] ),
    .S(net373),
    .X(_0157_));
 sg13g2_mux2_1 _1784_ (.A0(net226),
    .A1(\cic_b.temp_delay[0][2] ),
    .S(net370),
    .X(_0158_));
 sg13g2_mux2_1 _1785_ (.A0(net295),
    .A1(\cic_b.temp_delay[0][3] ),
    .S(net367),
    .X(_0159_));
 sg13g2_mux2_1 _1786_ (.A0(\cic_b.delay[0][4] ),
    .A1(net217),
    .S(net367),
    .X(_0160_));
 sg13g2_nor2_1 _1787_ (.A(net146),
    .B(net355),
    .Y(_0393_));
 sg13g2_a21oi_1 _1788_ (.A1(_0717_),
    .A2(net355),
    .Y(_0161_),
    .B1(_0393_));
 sg13g2_mux2_1 _1789_ (.A0(\cic_b.delay[0][6] ),
    .A1(net223),
    .S(net363),
    .X(_0162_));
 sg13g2_mux2_1 _1790_ (.A0(\cic_b.delay[0][7] ),
    .A1(net230),
    .S(net363),
    .X(_0163_));
 sg13g2_mux2_1 _1791_ (.A0(\cic_b.delay[0][8] ),
    .A1(net101),
    .S(net361),
    .X(_0164_));
 sg13g2_nor2_1 _1792_ (.A(net87),
    .B(net352),
    .Y(_0394_));
 sg13g2_a21oi_1 _1793_ (.A1(_0719_),
    .A2(net352),
    .Y(_0165_),
    .B1(_0394_));
 sg13g2_mux2_1 _1794_ (.A0(\cic_b.delay[0][10] ),
    .A1(net248),
    .S(net361),
    .X(_0166_));
 sg13g2_mux2_1 _1795_ (.A0(net209),
    .A1(\cic_b.temp_delay[0][11] ),
    .S(net361),
    .X(_0167_));
 sg13g2_mux2_1 _1796_ (.A0(net192),
    .A1(\cic_b.temp_delay[0][12] ),
    .S(net361),
    .X(_0168_));
 sg13g2_nand2b_2 _1797_ (.Y(_0395_),
    .B(net205),
    .A_N(\cic_b.integrator[1][0] ));
 sg13g2_nand2b_1 _1798_ (.Y(_0396_),
    .B(\cic_b.integrator[1][0] ),
    .A_N(net205));
 sg13g2_a21oi_1 _1799_ (.A1(_0395_),
    .A2(_0396_),
    .Y(_0397_),
    .B1(net357));
 sg13g2_a21o_1 _1800_ (.A2(net357),
    .A1(net528),
    .B1(_0397_),
    .X(_0169_));
 sg13g2_nor2_1 _1801_ (.A(net318),
    .B(net370),
    .Y(_0398_));
 sg13g2_nor2b_1 _1802_ (.A(\cic_b.delay[0][1] ),
    .B_N(\cic_b.integrator[1][1] ),
    .Y(_0399_));
 sg13g2_xnor2_1 _1803_ (.Y(_0400_),
    .A(\cic_b.integrator[1][1] ),
    .B(net315));
 sg13g2_xnor2_1 _1804_ (.Y(_0401_),
    .A(_0395_),
    .B(_0400_));
 sg13g2_a21oi_1 _1805_ (.A1(net373),
    .A2(_0401_),
    .Y(_0170_),
    .B1(_0398_));
 sg13g2_nor2_1 _1806_ (.A(net277),
    .B(net370),
    .Y(_0402_));
 sg13g2_nor2b_1 _1807_ (.A(net485),
    .B_N(\cic_b.integrator[1][2] ),
    .Y(_0403_));
 sg13g2_nand2b_1 _1808_ (.Y(_0404_),
    .B(net226),
    .A_N(\cic_b.integrator[1][2] ));
 sg13g2_nor2b_1 _1809_ (.A(_0403_),
    .B_N(_0404_),
    .Y(_0405_));
 sg13g2_a21o_1 _1810_ (.A2(_0400_),
    .A1(_0395_),
    .B1(_0399_),
    .X(_0406_));
 sg13g2_xnor2_1 _1811_ (.Y(_0407_),
    .A(_0405_),
    .B(_0406_));
 sg13g2_a21oi_1 _1812_ (.A1(net370),
    .A2(_0407_),
    .Y(_0171_),
    .B1(_0402_));
 sg13g2_nor2_1 _1813_ (.A(net344),
    .B(net367),
    .Y(_0408_));
 sg13g2_nand2b_1 _1814_ (.Y(_0409_),
    .B(\cic_b.integrator[1][3] ),
    .A_N(\cic_b.delay[0][3] ));
 sg13g2_xor2_1 _1815_ (.B(net295),
    .A(\cic_b.integrator[1][3] ),
    .X(_0410_));
 sg13g2_a21oi_2 _1816_ (.B1(_0403_),
    .Y(_0411_),
    .A2(_0406_),
    .A1(_0404_));
 sg13g2_xnor2_1 _1817_ (.Y(_0412_),
    .A(_0410_),
    .B(_0411_));
 sg13g2_a21oi_1 _1818_ (.A1(net367),
    .A2(_0412_),
    .Y(_0172_),
    .B1(_0408_));
 sg13g2_nor2_1 _1819_ (.A(net511),
    .B(net367),
    .Y(_0413_));
 sg13g2_o21ai_1 _1820_ (.B1(_0409_),
    .Y(_0414_),
    .A1(_0410_),
    .A2(_0411_));
 sg13g2_nor2b_1 _1821_ (.A(\cic_b.delay[0][4] ),
    .B_N(\cic_b.integrator[1][4] ),
    .Y(_0415_));
 sg13g2_xnor2_1 _1822_ (.Y(_0416_),
    .A(\cic_b.integrator[1][4] ),
    .B(\cic_b.delay[0][4] ));
 sg13g2_nand2_1 _1823_ (.Y(_0417_),
    .A(_0414_),
    .B(_0416_));
 sg13g2_xnor2_1 _1824_ (.Y(_0418_),
    .A(_0414_),
    .B(_0416_));
 sg13g2_a21oi_1 _1825_ (.A1(net367),
    .A2(_0418_),
    .Y(_0173_),
    .B1(_0413_));
 sg13g2_nor2_1 _1826_ (.A(\cic_b.integrator[1][5] ),
    .B(_0717_),
    .Y(_0419_));
 sg13g2_xor2_1 _1827_ (.B(\cic_b.delay[0][5] ),
    .A(\cic_b.integrator[1][5] ),
    .X(_0420_));
 sg13g2_a21oi_1 _1828_ (.A1(_0414_),
    .A2(_0416_),
    .Y(_0421_),
    .B1(_0415_));
 sg13g2_xnor2_1 _1829_ (.Y(_0422_),
    .A(_0420_),
    .B(_0421_));
 sg13g2_nor2_1 _1830_ (.A(net540),
    .B(net367),
    .Y(_0423_));
 sg13g2_a21oi_1 _1831_ (.A1(net367),
    .A2(_0422_),
    .Y(_0174_),
    .B1(_0423_));
 sg13g2_nor2_1 _1832_ (.A(net544),
    .B(net366),
    .Y(_0424_));
 sg13g2_nor2b_1 _1833_ (.A(\cic_b.delay[0][6] ),
    .B_N(\cic_b.integrator[1][6] ),
    .Y(_0425_));
 sg13g2_nand2b_1 _1834_ (.Y(_0426_),
    .B(\cic_b.delay[0][6] ),
    .A_N(\cic_b.integrator[1][6] ));
 sg13g2_xor2_1 _1835_ (.B(\cic_b.delay[0][6] ),
    .A(\cic_b.integrator[1][6] ),
    .X(_0427_));
 sg13g2_a21oi_1 _1836_ (.A1(\cic_b.integrator[1][5] ),
    .A2(_0717_),
    .Y(_0428_),
    .B1(_0415_));
 sg13g2_a21oi_1 _1837_ (.A1(_0417_),
    .A2(_0428_),
    .Y(_0429_),
    .B1(_0419_));
 sg13g2_xor2_1 _1838_ (.B(_0429_),
    .A(_0427_),
    .X(_0430_));
 sg13g2_a21oi_1 _1839_ (.A1(net363),
    .A2(_0430_),
    .Y(_0175_),
    .B1(_0424_));
 sg13g2_nor2_1 _1840_ (.A(net496),
    .B(net363),
    .Y(_0431_));
 sg13g2_nand2b_1 _1841_ (.Y(_0432_),
    .B(\cic_b.delay[0][7] ),
    .A_N(\cic_b.integrator[1][7] ));
 sg13g2_nor2b_1 _1842_ (.A(\cic_b.delay[0][7] ),
    .B_N(\cic_b.integrator[1][7] ),
    .Y(_0433_));
 sg13g2_xor2_1 _1843_ (.B(\cic_b.delay[0][7] ),
    .A(\cic_b.integrator[1][7] ),
    .X(_0434_));
 sg13g2_a21oi_1 _1844_ (.A1(_0426_),
    .A2(_0429_),
    .Y(_0435_),
    .B1(_0425_));
 sg13g2_xnor2_1 _1845_ (.Y(_0436_),
    .A(_0434_),
    .B(_0435_));
 sg13g2_a21oi_1 _1846_ (.A1(net363),
    .A2(_0436_),
    .Y(_0176_),
    .B1(_0431_));
 sg13g2_nor2_1 _1847_ (.A(net312),
    .B(net363),
    .Y(_0437_));
 sg13g2_nor2_1 _1848_ (.A(_0427_),
    .B(_0434_),
    .Y(_0438_));
 sg13g2_nand2_1 _1849_ (.Y(_0439_),
    .A(_0416_),
    .B(_0438_));
 sg13g2_nor2_1 _1850_ (.A(_0420_),
    .B(_0439_),
    .Y(_0440_));
 sg13g2_nor2_1 _1851_ (.A(_0419_),
    .B(_0428_),
    .Y(_0441_));
 sg13g2_a21o_1 _1852_ (.A2(_0432_),
    .A1(_0425_),
    .B1(_0433_),
    .X(_0442_));
 sg13g2_a221oi_1 _1853_ (.B2(_0438_),
    .C1(_0442_),
    .B1(_0441_),
    .A1(_0414_),
    .Y(_0443_),
    .A2(_0440_));
 sg13g2_nand2b_1 _1854_ (.Y(_0444_),
    .B(\cic_b.integrator[1][8] ),
    .A_N(\cic_b.delay[0][8] ));
 sg13g2_xor2_1 _1855_ (.B(net498),
    .A(\cic_b.integrator[1][8] ),
    .X(_0445_));
 sg13g2_xnor2_1 _1856_ (.Y(_0446_),
    .A(_0443_),
    .B(_0445_));
 sg13g2_a21oi_1 _1857_ (.A1(net363),
    .A2(_0446_),
    .Y(_0177_),
    .B1(_0437_));
 sg13g2_xor2_1 _1858_ (.B(\cic_b.delay[0][9] ),
    .A(\cic_b.integrator[1][9] ),
    .X(_0447_));
 sg13g2_o21ai_1 _1859_ (.B1(_0444_),
    .Y(_0448_),
    .A1(_0443_),
    .A2(_0445_));
 sg13g2_xor2_1 _1860_ (.B(_0448_),
    .A(_0447_),
    .X(_0449_));
 sg13g2_nand2_1 _1861_ (.Y(_0450_),
    .A(net474),
    .B(net354));
 sg13g2_o21ai_1 _1862_ (.B1(_0450_),
    .Y(_0178_),
    .A1(net353),
    .A2(_0449_));
 sg13g2_nor2_1 _1863_ (.A(net214),
    .B(net362),
    .Y(_0451_));
 sg13g2_nor2b_1 _1864_ (.A(\cic_b.delay[0][10] ),
    .B_N(\cic_b.integrator[1][10] ),
    .Y(_0452_));
 sg13g2_xnor2_1 _1865_ (.Y(_0453_),
    .A(\cic_b.integrator[1][10] ),
    .B(\cic_b.delay[0][10] ));
 sg13g2_inv_1 _1866_ (.Y(_0454_),
    .A(_0453_));
 sg13g2_a21oi_1 _1867_ (.A1(_0718_),
    .A2(\cic_b.delay[0][9] ),
    .Y(_0455_),
    .B1(_0444_));
 sg13g2_a21oi_1 _1868_ (.A1(\cic_b.integrator[1][9] ),
    .A2(_0719_),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_or2_1 _1869_ (.X(_0457_),
    .B(_0447_),
    .A(_0445_));
 sg13g2_o21ai_1 _1870_ (.B1(_0456_),
    .Y(_0458_),
    .A1(_0443_),
    .A2(_0457_));
 sg13g2_xnor2_1 _1871_ (.Y(_0459_),
    .A(_0453_),
    .B(_0458_));
 sg13g2_a21oi_1 _1872_ (.A1(net361),
    .A2(_0459_),
    .Y(_0179_),
    .B1(_0451_));
 sg13g2_nor2_1 _1873_ (.A(net201),
    .B(net360),
    .Y(_0460_));
 sg13g2_nor2b_1 _1874_ (.A(\cic_b.delay[0][11] ),
    .B_N(\cic_b.integrator[1][11] ),
    .Y(_0461_));
 sg13g2_nand2b_1 _1875_ (.Y(_0462_),
    .B(\cic_b.delay[0][11] ),
    .A_N(\cic_b.integrator[1][11] ));
 sg13g2_nand2b_1 _1876_ (.Y(_0463_),
    .B(_0462_),
    .A_N(_0461_));
 sg13g2_a21oi_1 _1877_ (.A1(_0453_),
    .A2(_0458_),
    .Y(_0464_),
    .B1(_0452_));
 sg13g2_xnor2_1 _1878_ (.Y(_0465_),
    .A(_0463_),
    .B(_0464_));
 sg13g2_a21oi_1 _1879_ (.A1(net360),
    .A2(_0465_),
    .Y(_0180_),
    .B1(_0460_));
 sg13g2_nor2_1 _1880_ (.A(net207),
    .B(net360),
    .Y(_0466_));
 sg13g2_nor2_1 _1881_ (.A(_0454_),
    .B(_0463_),
    .Y(_0467_));
 sg13g2_a221oi_1 _1882_ (.B2(_0458_),
    .C1(_0461_),
    .B1(_0467_),
    .A1(_0452_),
    .Y(_0468_),
    .A2(_0462_));
 sg13g2_xor2_1 _1883_ (.B(net192),
    .A(\cic_b.integrator[1][12] ),
    .X(_0469_));
 sg13g2_xnor2_1 _1884_ (.Y(_0470_),
    .A(_0468_),
    .B(_0469_));
 sg13g2_a21oi_1 _1885_ (.A1(net361),
    .A2(_0470_),
    .Y(_0181_),
    .B1(_0466_));
 sg13g2_mux2_1 _1886_ (.A0(net181),
    .A1(net137),
    .S(net371),
    .X(_0182_));
 sg13g2_mux2_1 _1887_ (.A0(net225),
    .A1(net142),
    .S(net372),
    .X(_0183_));
 sg13g2_mux2_1 _1888_ (.A0(net144),
    .A1(net114),
    .S(net371),
    .X(_0184_));
 sg13g2_nor2_1 _1889_ (.A(net78),
    .B(net358),
    .Y(_0471_));
 sg13g2_a21oi_1 _1890_ (.A1(_0701_),
    .A2(net358),
    .Y(_0185_),
    .B1(_0471_));
 sg13g2_nor2_1 _1891_ (.A(net94),
    .B(net356),
    .Y(_0472_));
 sg13g2_a21oi_1 _1892_ (.A1(_0702_),
    .A2(net356),
    .Y(_0186_),
    .B1(_0472_));
 sg13g2_nor2_1 _1893_ (.A(net89),
    .B(net355),
    .Y(_0473_));
 sg13g2_a21oi_1 _1894_ (.A1(_0703_),
    .A2(net355),
    .Y(_0187_),
    .B1(_0473_));
 sg13g2_mux2_1 _1895_ (.A0(net302),
    .A1(net136),
    .S(net369),
    .X(_0188_));
 sg13g2_mux2_1 _1896_ (.A0(net284),
    .A1(net48),
    .S(net369),
    .X(_0189_));
 sg13g2_mux2_1 _1897_ (.A0(net250),
    .A1(net124),
    .S(net365),
    .X(_0190_));
 sg13g2_mux2_1 _1898_ (.A0(net495),
    .A1(net44),
    .S(net365),
    .X(_0191_));
 sg13g2_mux2_1 _1899_ (.A0(net325),
    .A1(net133),
    .S(net364),
    .X(_0192_));
 sg13g2_mux2_1 _1900_ (.A0(net488),
    .A1(net185),
    .S(net364),
    .X(_0193_));
 sg13g2_mux2_1 _1901_ (.A0(net305),
    .A1(net283),
    .S(net360),
    .X(_0194_));
 sg13g2_mux2_1 _1902_ (.A0(net253),
    .A1(\cic_b.temp_delay[1][0] ),
    .S(net370),
    .X(_0195_));
 sg13g2_mux2_1 _1903_ (.A0(\cic_b.delay[1][1] ),
    .A1(net261),
    .S(net370),
    .X(_0196_));
 sg13g2_mux2_1 _1904_ (.A0(\cic_b.delay[1][2] ),
    .A1(net275),
    .S(net370),
    .X(_0197_));
 sg13g2_mux2_1 _1905_ (.A0(net111),
    .A1(net321),
    .S(net370),
    .X(_0198_));
 sg13g2_mux2_1 _1906_ (.A0(net130),
    .A1(net486),
    .S(net369),
    .X(_0199_));
 sg13g2_nor2_1 _1907_ (.A(net153),
    .B(net356),
    .Y(_0474_));
 sg13g2_a21oi_1 _1908_ (.A1(_0721_),
    .A2(net356),
    .Y(_0200_),
    .B1(_0474_));
 sg13g2_mux2_1 _1909_ (.A0(net326),
    .A1(\cic_b.temp_delay[1][6] ),
    .S(net365),
    .X(_0201_));
 sg13g2_mux2_1 _1910_ (.A0(net239),
    .A1(\cic_b.temp_delay[1][7] ),
    .S(net363),
    .X(_0202_));
 sg13g2_mux2_1 _1911_ (.A0(\cic_b.delay[1][8] ),
    .A1(net310),
    .S(net364),
    .X(_0203_));
 sg13g2_nor2_1 _1912_ (.A(net97),
    .B(net354),
    .Y(_0475_));
 sg13g2_a21oi_1 _1913_ (.A1(_0723_),
    .A2(net354),
    .Y(_0204_),
    .B1(_0475_));
 sg13g2_mux2_1 _1914_ (.A0(net179),
    .A1(\cic_b.temp_delay[1][10] ),
    .S(net362),
    .X(_0205_));
 sg13g2_mux2_1 _1915_ (.A0(net211),
    .A1(\cic_b.temp_delay[1][11] ),
    .S(net362),
    .X(_0206_));
 sg13g2_mux2_1 _1916_ (.A0(net171),
    .A1(\cic_b.temp_delay[1][12] ),
    .S(net360),
    .X(_0207_));
 sg13g2_nor2_1 _1917_ (.A(net137),
    .B(net371),
    .Y(_0476_));
 sg13g2_nor2b_1 _1918_ (.A(\cic_b.temp_comb[0][0] ),
    .B_N(\cic_b.delay[1][0] ),
    .Y(_0477_));
 sg13g2_xnor2_1 _1919_ (.Y(_0478_),
    .A(\cic_b.temp_comb[0][0] ),
    .B(\cic_b.delay[1][0] ));
 sg13g2_a21oi_1 _1920_ (.A1(net371),
    .A2(_0478_),
    .Y(_0208_),
    .B1(_0476_));
 sg13g2_nor2_1 _1921_ (.A(net142),
    .B(net371),
    .Y(_0479_));
 sg13g2_nand2b_1 _1922_ (.Y(_0480_),
    .B(\cic_b.temp_comb[0][1] ),
    .A_N(\cic_b.delay[1][1] ));
 sg13g2_xor2_1 _1923_ (.B(\cic_b.delay[1][1] ),
    .A(\cic_b.temp_comb[0][1] ),
    .X(_0481_));
 sg13g2_xnor2_1 _1924_ (.Y(_0482_),
    .A(_0477_),
    .B(_0481_));
 sg13g2_a21oi_1 _1925_ (.A1(net371),
    .A2(_0482_),
    .Y(_0209_),
    .B1(_0479_));
 sg13g2_nor2_1 _1926_ (.A(net114),
    .B(net371),
    .Y(_0483_));
 sg13g2_nor2b_1 _1927_ (.A(\cic_b.delay[1][2] ),
    .B_N(\cic_b.temp_comb[0][2] ),
    .Y(_0484_));
 sg13g2_xnor2_1 _1928_ (.Y(_0485_),
    .A(\cic_b.temp_comb[0][2] ),
    .B(\cic_b.delay[1][2] ));
 sg13g2_o21ai_1 _1929_ (.B1(_0480_),
    .Y(_0486_),
    .A1(_0477_),
    .A2(_0481_));
 sg13g2_xnor2_1 _1930_ (.Y(_0487_),
    .A(_0485_),
    .B(_0486_));
 sg13g2_a21oi_1 _1931_ (.A1(net371),
    .A2(_0487_),
    .Y(_0210_),
    .B1(_0483_));
 sg13g2_nor2_1 _1932_ (.A(net78),
    .B(net372),
    .Y(_0488_));
 sg13g2_nand2b_1 _1933_ (.Y(_0489_),
    .B(\cic_b.temp_comb[0][3] ),
    .A_N(\cic_b.delay[1][3] ));
 sg13g2_xor2_1 _1934_ (.B(net111),
    .A(\cic_b.temp_comb[0][3] ),
    .X(_0490_));
 sg13g2_a21oi_2 _1935_ (.B1(_0484_),
    .Y(_0491_),
    .A2(_0486_),
    .A1(_0485_));
 sg13g2_xnor2_1 _1936_ (.Y(_0492_),
    .A(_0490_),
    .B(_0491_));
 sg13g2_a21oi_1 _1937_ (.A1(net372),
    .A2(net112),
    .Y(_0211_),
    .B1(_0488_));
 sg13g2_o21ai_1 _1938_ (.B1(_0489_),
    .Y(_0493_),
    .A1(_0490_),
    .A2(_0491_));
 sg13g2_nor2b_1 _1939_ (.A(\cic_b.delay[1][4] ),
    .B_N(\cic_b.temp_comb[0][4] ),
    .Y(_0494_));
 sg13g2_xor2_1 _1940_ (.B(\cic_b.delay[1][4] ),
    .A(\cic_b.temp_comb[0][4] ),
    .X(_0495_));
 sg13g2_nor2b_1 _1941_ (.A(_0495_),
    .B_N(_0493_),
    .Y(_0496_));
 sg13g2_nor2_1 _1942_ (.A(net94),
    .B(net368),
    .Y(_0497_));
 sg13g2_xor2_1 _1943_ (.B(_0495_),
    .A(_0493_),
    .X(_0498_));
 sg13g2_a21oi_1 _1944_ (.A1(net368),
    .A2(_0498_),
    .Y(_0212_),
    .B1(_0497_));
 sg13g2_nor2_1 _1945_ (.A(net89),
    .B(net368),
    .Y(_0499_));
 sg13g2_xor2_1 _1946_ (.B(net614),
    .A(\cic_b.temp_comb[0][5] ),
    .X(_0500_));
 sg13g2_nor2_1 _1947_ (.A(_0494_),
    .B(_0496_),
    .Y(_0501_));
 sg13g2_xnor2_1 _1948_ (.Y(_0502_),
    .A(_0500_),
    .B(_0501_));
 sg13g2_a21oi_1 _1949_ (.A1(net368),
    .A2(_0502_),
    .Y(_0213_),
    .B1(_0499_));
 sg13g2_nor2_1 _1950_ (.A(net136),
    .B(net368),
    .Y(_0503_));
 sg13g2_nand2b_1 _1951_ (.Y(_0504_),
    .B(net612),
    .A_N(\cic_b.delay[1][6] ));
 sg13g2_xor2_1 _1952_ (.B(\cic_b.delay[1][6] ),
    .A(\cic_b.temp_comb[0][6] ),
    .X(_0505_));
 sg13g2_or2_1 _1953_ (.X(_0506_),
    .B(_0500_),
    .A(_0495_));
 sg13g2_inv_1 _1954_ (.Y(_0507_),
    .A(_0506_));
 sg13g2_a21oi_1 _1955_ (.A1(\cic_b.temp_comb[0][5] ),
    .A2(_0721_),
    .Y(_0508_),
    .B1(_0494_));
 sg13g2_a21oi_1 _1956_ (.A1(_0720_),
    .A2(\cic_b.delay[1][5] ),
    .Y(_0509_),
    .B1(_0508_));
 sg13g2_a21oi_1 _1957_ (.A1(_0493_),
    .A2(_0507_),
    .Y(_0510_),
    .B1(_0509_));
 sg13g2_xnor2_1 _1958_ (.Y(_0511_),
    .A(_0505_),
    .B(_0510_));
 sg13g2_a21oi_1 _1959_ (.A1(net368),
    .A2(_0511_),
    .Y(_0214_),
    .B1(_0503_));
 sg13g2_nor2b_1 _1960_ (.A(\cic_b.temp_comb[0][7] ),
    .B_N(\cic_b.delay[1][7] ),
    .Y(_0512_));
 sg13g2_nand2b_1 _1961_ (.Y(_0513_),
    .B(\cic_b.temp_comb[0][7] ),
    .A_N(\cic_b.delay[1][7] ));
 sg13g2_nand2b_1 _1962_ (.Y(_0514_),
    .B(_0513_),
    .A_N(_0512_));
 sg13g2_o21ai_1 _1963_ (.B1(_0504_),
    .Y(_0515_),
    .A1(_0505_),
    .A2(_0510_));
 sg13g2_xor2_1 _1964_ (.B(_0515_),
    .A(_0514_),
    .X(_0516_));
 sg13g2_nand2_1 _1965_ (.Y(_0517_),
    .A(net48),
    .B(net356));
 sg13g2_o21ai_1 _1966_ (.B1(_0517_),
    .Y(_0215_),
    .A1(net356),
    .A2(_0516_));
 sg13g2_nor2_1 _1967_ (.A(net124),
    .B(net365),
    .Y(_0518_));
 sg13g2_nand2b_1 _1968_ (.Y(_0519_),
    .B(\cic_b.temp_comb[0][8] ),
    .A_N(\cic_b.delay[1][8] ));
 sg13g2_xor2_1 _1969_ (.B(\cic_b.delay[1][8] ),
    .A(\cic_b.temp_comb[0][8] ),
    .X(_0520_));
 sg13g2_o21ai_1 _1970_ (.B1(_0513_),
    .Y(_0521_),
    .A1(_0504_),
    .A2(_0512_));
 sg13g2_nor2_1 _1971_ (.A(_0505_),
    .B(_0514_),
    .Y(_0522_));
 sg13g2_nor3_1 _1972_ (.A(_0505_),
    .B(_0506_),
    .C(_0514_),
    .Y(_0523_));
 sg13g2_a221oi_1 _1973_ (.B2(_0493_),
    .C1(_0521_),
    .B1(_0523_),
    .A1(_0509_),
    .Y(_0524_),
    .A2(_0522_));
 sg13g2_xnor2_1 _1974_ (.Y(_0525_),
    .A(_0520_),
    .B(_0524_));
 sg13g2_a21oi_1 _1975_ (.A1(net365),
    .A2(_0525_),
    .Y(_0216_),
    .B1(_0518_));
 sg13g2_xnor2_1 _1976_ (.Y(_0526_),
    .A(\cic_b.temp_comb[0][9] ),
    .B(\cic_b.delay[1][9] ));
 sg13g2_o21ai_1 _1977_ (.B1(_0519_),
    .Y(_0527_),
    .A1(_0520_),
    .A2(_0524_));
 sg13g2_xnor2_1 _1978_ (.Y(_0528_),
    .A(_0526_),
    .B(_0527_));
 sg13g2_nand2_1 _1979_ (.Y(_0529_),
    .A(net44),
    .B(net353));
 sg13g2_o21ai_1 _1980_ (.B1(_0529_),
    .Y(_0217_),
    .A1(net353),
    .A2(_0528_));
 sg13g2_nor2_1 _1981_ (.A(net133),
    .B(net364),
    .Y(_0530_));
 sg13g2_nand2b_1 _1982_ (.Y(_0531_),
    .B(_0526_),
    .A_N(_0520_));
 sg13g2_a21oi_1 _1983_ (.A1(_0722_),
    .A2(\cic_b.delay[1][9] ),
    .Y(_0532_),
    .B1(_0519_));
 sg13g2_a21oi_1 _1984_ (.A1(\cic_b.temp_comb[0][9] ),
    .A2(_0723_),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_o21ai_1 _1985_ (.B1(_0533_),
    .Y(_0534_),
    .A1(_0524_),
    .A2(_0531_));
 sg13g2_nor2b_1 _1986_ (.A(\cic_b.delay[1][10] ),
    .B_N(\cic_b.temp_comb[0][10] ),
    .Y(_0535_));
 sg13g2_nor2b_1 _1987_ (.A(\cic_b.temp_comb[0][10] ),
    .B_N(\cic_b.delay[1][10] ),
    .Y(_0536_));
 sg13g2_nor2_1 _1988_ (.A(_0535_),
    .B(_0536_),
    .Y(_0537_));
 sg13g2_xnor2_1 _1989_ (.Y(_0538_),
    .A(_0534_),
    .B(_0537_));
 sg13g2_a21oi_1 _1990_ (.A1(net364),
    .A2(_0538_),
    .Y(_0218_),
    .B1(_0530_));
 sg13g2_nor2_1 _1991_ (.A(net185),
    .B(net364),
    .Y(_0539_));
 sg13g2_nor2b_1 _1992_ (.A(net211),
    .B_N(\cic_b.temp_comb[0][11] ),
    .Y(_0540_));
 sg13g2_nand2b_1 _1993_ (.Y(_0541_),
    .B(\cic_b.delay[1][11] ),
    .A_N(\cic_b.temp_comb[0][11] ));
 sg13g2_nand2b_1 _1994_ (.Y(_0542_),
    .B(_0541_),
    .A_N(_0540_));
 sg13g2_a21oi_1 _1995_ (.A1(_0534_),
    .A2(_0537_),
    .Y(_0543_),
    .B1(_0535_));
 sg13g2_xnor2_1 _1996_ (.Y(_0544_),
    .A(_0542_),
    .B(_0543_));
 sg13g2_a21oi_1 _1997_ (.A1(net360),
    .A2(_0544_),
    .Y(_0219_),
    .B1(_0539_));
 sg13g2_nor2_1 _1998_ (.A(net283),
    .B(net360),
    .Y(_0545_));
 sg13g2_nor3_1 _1999_ (.A(_0535_),
    .B(_0536_),
    .C(_0542_),
    .Y(_0546_));
 sg13g2_a221oi_1 _2000_ (.B2(_0534_),
    .C1(_0540_),
    .B1(_0546_),
    .A1(_0535_),
    .Y(_0547_),
    .A2(_0541_));
 sg13g2_xor2_1 _2001_ (.B(net171),
    .A(net207),
    .X(_0548_));
 sg13g2_xnor2_1 _2002_ (.Y(_0549_),
    .A(_0547_),
    .B(_0548_));
 sg13g2_a21oi_1 _2003_ (.A1(net360),
    .A2(_0549_),
    .Y(_0220_),
    .B1(_0545_));
 sg13g2_mux2_1 _2004_ (.A0(net502),
    .A1(net291),
    .S(net381),
    .X(_0221_));
 sg13g2_mux2_1 _2005_ (.A0(\cic_a.temp_comb[0][1] ),
    .A1(net257),
    .S(net381),
    .X(_0222_));
 sg13g2_mux2_1 _2006_ (.A0(\cic_a.temp_comb[0][2] ),
    .A1(net259),
    .S(net381),
    .X(_0223_));
 sg13g2_mux2_1 _2007_ (.A0(\cic_a.temp_comb[0][3] ),
    .A1(net234),
    .S(net382),
    .X(_0224_));
 sg13g2_mux2_1 _2008_ (.A0(\cic_a.temp_comb[0][4] ),
    .A1(net263),
    .S(net380),
    .X(_0225_));
 sg13g2_mux2_1 _2009_ (.A0(\cic_a.temp_comb[0][5] ),
    .A1(net267),
    .S(net382),
    .X(_0226_));
 sg13g2_mux2_1 _2010_ (.A0(\cic_a.temp_comb[0][6] ),
    .A1(net303),
    .S(net377),
    .X(_0227_));
 sg13g2_mux2_1 _2011_ (.A0(\cic_a.temp_comb[0][7] ),
    .A1(net479),
    .S(net378),
    .X(_0228_));
 sg13g2_mux2_1 _2012_ (.A0(\cic_a.temp_comb[0][8] ),
    .A1(net342),
    .S(net377),
    .X(_0229_));
 sg13g2_nor2_1 _2013_ (.A(net85),
    .B(net387),
    .Y(_0550_));
 sg13g2_a21oi_1 _2014_ (.A1(_0711_),
    .A2(net387),
    .Y(_0230_),
    .B1(_0550_));
 sg13g2_mux2_1 _2015_ (.A0(\cic_a.temp_comb[0][10] ),
    .A1(net269),
    .S(net377),
    .X(_0231_));
 sg13g2_mux2_1 _2016_ (.A0(net476),
    .A1(net499),
    .S(net377),
    .X(_0232_));
 sg13g2_mux2_1 _2017_ (.A0(net198),
    .A1(net274),
    .S(net375),
    .X(_0233_));
 sg13g2_mux2_1 _2018_ (.A0(\cic_b.integrator[1][0] ),
    .A1(net297),
    .S(net357),
    .X(_0234_));
 sg13g2_mux2_1 _2019_ (.A0(\cic_b.integrator[1][1] ),
    .A1(net338),
    .S(net358),
    .X(_0235_));
 sg13g2_mux2_1 _2020_ (.A0(\cic_b.integrator[1][2] ),
    .A1(net333),
    .S(net357),
    .X(_0236_));
 sg13g2_mux2_1 _2021_ (.A0(\cic_b.integrator[1][3] ),
    .A1(net322),
    .S(net355),
    .X(_0237_));
 sg13g2_mux2_1 _2022_ (.A0(net346),
    .A1(net217),
    .S(net355),
    .X(_0238_));
 sg13g2_mux2_1 _2023_ (.A0(net492),
    .A1(net146),
    .S(net355),
    .X(_0239_));
 sg13g2_mux2_1 _2024_ (.A0(net238),
    .A1(net223),
    .S(net353),
    .X(_0240_));
 sg13g2_mux2_1 _2025_ (.A0(net306),
    .A1(net230),
    .S(net353),
    .X(_0241_));
 sg13g2_mux2_1 _2026_ (.A0(net471),
    .A1(net101),
    .S(net352),
    .X(_0242_));
 sg13g2_nor2_1 _2027_ (.A(net87),
    .B(net361),
    .Y(_0551_));
 sg13g2_a21oi_1 _2028_ (.A1(_0718_),
    .A2(net361),
    .Y(_0243_),
    .B1(_0551_));
 sg13g2_mux2_1 _2029_ (.A0(net478),
    .A1(net248),
    .S(net352),
    .X(_0244_));
 sg13g2_mux2_1 _2030_ (.A0(\cic_b.integrator[1][11] ),
    .A1(net293),
    .S(net352),
    .X(_0245_));
 sg13g2_mux2_1 _2031_ (.A0(\cic_b.integrator[1][12] ),
    .A1(net232),
    .S(net352),
    .X(_0246_));
 sg13g2_a22oi_1 _2032_ (.Y(_0552_),
    .B1(_0861_),
    .B2(net37),
    .A2(net404),
    .A1(\cic_a.filtered_out[0] ));
 sg13g2_inv_1 _2033_ (.Y(_0247_),
    .A(net38));
 sg13g2_a22oi_1 _2034_ (.Y(_0553_),
    .B1(\cic_a.filtered_out[1] ),
    .B2(net404),
    .A2(net37),
    .A1(net411));
 sg13g2_o21ai_1 _2035_ (.B1(_0553_),
    .Y(_0248_),
    .A1(_0691_),
    .A2(_0862_));
 sg13g2_a22oi_1 _2036_ (.Y(_0554_),
    .B1(net129),
    .B2(net404),
    .A2(net106),
    .A1(net411));
 sg13g2_o21ai_1 _2037_ (.B1(_0554_),
    .Y(_0249_),
    .A1(_0692_),
    .A2(_0862_));
 sg13g2_nand2_1 _2038_ (.Y(_0555_),
    .A(net412),
    .B(net71));
 sg13g2_a22oi_1 _2039_ (.Y(_0556_),
    .B1(_0861_),
    .B2(\serializer_a.shift_reg[3] ),
    .A2(net404),
    .A1(\cic_a.filtered_out[3] ));
 sg13g2_nand2_1 _2040_ (.Y(_0250_),
    .A(net72),
    .B(_0556_));
 sg13g2_a22oi_1 _2041_ (.Y(_0557_),
    .B1(\cic_a.filtered_out[4] ),
    .B2(net403),
    .A2(net115),
    .A1(net410));
 sg13g2_o21ai_1 _2042_ (.B1(net116),
    .Y(_0251_),
    .A1(_0694_),
    .A2(net397));
 sg13g2_nand2_1 _2043_ (.Y(_0558_),
    .A(net410),
    .B(net25));
 sg13g2_a22oi_1 _2044_ (.Y(_0559_),
    .B1(_0861_),
    .B2(\serializer_a.shift_reg[5] ),
    .A2(net403),
    .A1(\cic_a.filtered_out[5] ));
 sg13g2_nand2_1 _2045_ (.Y(_0252_),
    .A(_0558_),
    .B(_0559_));
 sg13g2_nand2_1 _2046_ (.Y(_0560_),
    .A(net410),
    .B(net164));
 sg13g2_a22oi_1 _2047_ (.Y(_0561_),
    .B1(_0861_),
    .B2(\serializer_a.shift_reg[6] ),
    .A2(net403),
    .A1(\cic_a.filtered_out[6] ));
 sg13g2_nand2_1 _2048_ (.Y(_0253_),
    .A(_0560_),
    .B(_0561_));
 sg13g2_a22oi_1 _2049_ (.Y(_0562_),
    .B1(\cic_a.filtered_out[7] ),
    .B2(net403),
    .A2(\serializer_a.shift_reg[6] ),
    .A1(net410));
 sg13g2_o21ai_1 _2050_ (.B1(_0562_),
    .Y(_0254_),
    .A1(_0696_),
    .A2(net397));
 sg13g2_a22oi_1 _2051_ (.Y(_0563_),
    .B1(net141),
    .B2(net403),
    .A2(net117),
    .A1(net410));
 sg13g2_o21ai_1 _2052_ (.B1(_0563_),
    .Y(_0255_),
    .A1(_0697_),
    .A2(net397));
 sg13g2_nand2_1 _2053_ (.Y(_0564_),
    .A(net410),
    .B(net64));
 sg13g2_a22oi_1 _2054_ (.Y(_0565_),
    .B1(_0861_),
    .B2(\serializer_a.shift_reg[9] ),
    .A2(net403),
    .A1(\cic_a.filtered_out[9] ));
 sg13g2_nand2_1 _2055_ (.Y(_0256_),
    .A(_0564_),
    .B(_0565_));
 sg13g2_a22oi_1 _2056_ (.Y(_0566_),
    .B1(\cic_a.filtered_out[10] ),
    .B2(net403),
    .A2(\serializer_a.shift_reg[9] ),
    .A1(net410));
 sg13g2_o21ai_1 _2057_ (.B1(_0566_),
    .Y(_0257_),
    .A1(_0698_),
    .A2(net397));
 sg13g2_a22oi_1 _2058_ (.Y(_0567_),
    .B1(\cic_a.filtered_out[11] ),
    .B2(net403),
    .A2(\serializer_a.shift_reg[10] ),
    .A1(net410));
 sg13g2_o21ai_1 _2059_ (.B1(_0567_),
    .Y(_0258_),
    .A1(_0699_),
    .A2(net397));
 sg13g2_a22oi_1 _2060_ (.Y(_0568_),
    .B1(\cic_a.filtered_out[12] ),
    .B2(net404),
    .A2(\serializer_a.shift_reg[11] ),
    .A1(net411));
 sg13g2_o21ai_1 _2061_ (.B1(_0568_),
    .Y(_0259_),
    .A1(_0728_),
    .A2(net397));
 sg13g2_mux2_1 _2062_ (.A0(\cic_b.temp_comb[0][0] ),
    .A1(net308),
    .S(net357),
    .X(_0260_));
 sg13g2_mux2_1 _2063_ (.A0(net318),
    .A1(net261),
    .S(net357),
    .X(_0261_));
 sg13g2_mux2_1 _2064_ (.A0(net277),
    .A1(net275),
    .S(net357),
    .X(_0262_));
 sg13g2_mux2_1 _2065_ (.A0(net344),
    .A1(net321),
    .S(net357),
    .X(_0263_));
 sg13g2_mux2_1 _2066_ (.A0(\cic_b.temp_comb[0][4] ),
    .A1(net486),
    .S(net355),
    .X(_0264_));
 sg13g2_nor2_1 _2067_ (.A(net153),
    .B(net368),
    .Y(_0569_));
 sg13g2_a21oi_1 _2068_ (.A1(_0720_),
    .A2(net368),
    .Y(_0265_),
    .B1(_0569_));
 sg13g2_mux2_1 _2069_ (.A0(\cic_b.temp_comb[0][6] ),
    .A1(net348),
    .S(net353),
    .X(_0266_));
 sg13g2_mux2_1 _2070_ (.A0(\cic_b.temp_comb[0][7] ),
    .A1(net493),
    .S(net353),
    .X(_0267_));
 sg13g2_mux2_1 _2071_ (.A0(net312),
    .A1(net310),
    .S(net353),
    .X(_0268_));
 sg13g2_nor2_1 _2072_ (.A(net97),
    .B(net364),
    .Y(_0570_));
 sg13g2_a21oi_1 _2073_ (.A1(_0722_),
    .A2(net364),
    .Y(_0269_),
    .B1(_0570_));
 sg13g2_mux2_1 _2074_ (.A0(net214),
    .A1(net290),
    .S(net352),
    .X(_0270_));
 sg13g2_mux2_1 _2075_ (.A0(net201),
    .A1(net347),
    .S(net352),
    .X(_0271_));
 sg13g2_mux2_1 _2076_ (.A0(net207),
    .A1(net510),
    .S(net354),
    .X(_0272_));
 sg13g2_a22oi_1 _2077_ (.Y(_0571_),
    .B1(_0865_),
    .B2(net62),
    .A2(net401),
    .A1(\cic_b.filtered_out[0] ));
 sg13g2_inv_1 _2078_ (.Y(_0273_),
    .A(net63));
 sg13g2_nand2_1 _2079_ (.Y(_0572_),
    .A(net408),
    .B(net62));
 sg13g2_a22oi_1 _2080_ (.Y(_0573_),
    .B1(_0865_),
    .B2(net81),
    .A2(net401),
    .A1(\cic_b.filtered_out[1] ));
 sg13g2_nand2_1 _2081_ (.Y(_0274_),
    .A(_0572_),
    .B(net82));
 sg13g2_a22oi_1 _2082_ (.Y(_0574_),
    .B1(net144),
    .B2(net401),
    .A2(net81),
    .A1(\serializer_b.sending ));
 sg13g2_o21ai_1 _2083_ (.B1(net145),
    .Y(_0275_),
    .A1(_0700_),
    .A2(_0866_));
 sg13g2_nand2_1 _2084_ (.Y(_0575_),
    .A(net408),
    .B(net27));
 sg13g2_a22oi_1 _2085_ (.Y(_0576_),
    .B1(_0865_),
    .B2(\serializer_b.shift_reg[3] ),
    .A2(net401),
    .A1(\cic_b.filtered_out[3] ));
 sg13g2_nand2_1 _2086_ (.Y(_0276_),
    .A(_0575_),
    .B(_0576_));
 sg13g2_nand2_1 _2087_ (.Y(_0577_),
    .A(net408),
    .B(net76));
 sg13g2_a22oi_1 _2088_ (.Y(_0578_),
    .B1(_0865_),
    .B2(net41),
    .A2(net400),
    .A1(\cic_b.filtered_out[4] ));
 sg13g2_nand2_1 _2089_ (.Y(_0277_),
    .A(_0577_),
    .B(_0578_));
 sg13g2_nand2_1 _2090_ (.Y(_0579_),
    .A(net409),
    .B(net41));
 sg13g2_a22oi_1 _2091_ (.Y(_0580_),
    .B1(_0865_),
    .B2(\serializer_b.shift_reg[5] ),
    .A2(net400),
    .A1(\cic_b.filtered_out[5] ));
 sg13g2_nand2_1 _2092_ (.Y(_0278_),
    .A(net42),
    .B(_0580_));
 sg13g2_a22oi_1 _2093_ (.Y(_0581_),
    .B1(\cic_b.filtered_out[6] ),
    .B2(net400),
    .A2(\serializer_b.shift_reg[5] ),
    .A1(net409));
 sg13g2_o21ai_1 _2094_ (.B1(_0581_),
    .Y(_0279_),
    .A1(_0704_),
    .A2(net396));
 sg13g2_a22oi_1 _2095_ (.Y(_0582_),
    .B1(\cic_b.filtered_out[7] ),
    .B2(net400),
    .A2(net149),
    .A1(net409));
 sg13g2_o21ai_1 _2096_ (.B1(_0582_),
    .Y(_0280_),
    .A1(_0705_),
    .A2(net396));
 sg13g2_a22oi_1 _2097_ (.Y(_0583_),
    .B1(\cic_b.filtered_out[8] ),
    .B2(net400),
    .A2(\serializer_b.shift_reg[7] ),
    .A1(net409));
 sg13g2_o21ai_1 _2098_ (.B1(_0583_),
    .Y(_0281_),
    .A1(_0706_),
    .A2(net396));
 sg13g2_a22oi_1 _2099_ (.Y(_0584_),
    .B1(net495),
    .B2(net400),
    .A2(net122),
    .A1(net409));
 sg13g2_o21ai_1 _2100_ (.B1(_0584_),
    .Y(_0282_),
    .A1(_0707_),
    .A2(net396));
 sg13g2_a22oi_1 _2101_ (.Y(_0585_),
    .B1(\cic_b.filtered_out[10] ),
    .B2(net400),
    .A2(\serializer_b.shift_reg[9] ),
    .A1(net409));
 sg13g2_o21ai_1 _2102_ (.B1(_0585_),
    .Y(_0283_),
    .A1(_0708_),
    .A2(net396));
 sg13g2_a22oi_1 _2103_ (.Y(_0586_),
    .B1(\cic_b.filtered_out[11] ),
    .B2(net400),
    .A2(\serializer_b.shift_reg[10] ),
    .A1(net409));
 sg13g2_o21ai_1 _2104_ (.B1(_0586_),
    .Y(_0284_),
    .A1(_0709_),
    .A2(net396));
 sg13g2_a22oi_1 _2105_ (.Y(_0587_),
    .B1(\cic_b.filtered_out[12] ),
    .B2(net401),
    .A2(\serializer_b.shift_reg[11] ),
    .A1(net408));
 sg13g2_o21ai_1 _2106_ (.B1(_0587_),
    .Y(_0285_),
    .A1(_0729_),
    .A2(net396));
 sg13g2_nor2_1 _2107_ (.A(net405),
    .B(net110),
    .Y(_0588_));
 sg13g2_a21oi_1 _2108_ (.A1(net110),
    .A2(_0870_),
    .Y(_0286_),
    .B1(_0588_));
 sg13g2_nand2_1 _2109_ (.Y(_0589_),
    .A(net166),
    .B(net399));
 sg13g2_and2_1 _2110_ (.A(net110),
    .B(net166),
    .X(_0590_));
 sg13g2_o21ai_1 _2111_ (.B1(_0589_),
    .Y(_0287_),
    .A1(_0871_),
    .A2(_0590_));
 sg13g2_nand3_1 _2112_ (.B(net51),
    .C(_0590_),
    .A(net405),
    .Y(_0591_));
 sg13g2_nand2_1 _2113_ (.Y(_0592_),
    .A(net402),
    .B(_0591_));
 sg13g2_a21oi_1 _2114_ (.A1(_0870_),
    .A2(_0590_),
    .Y(_0593_),
    .B1(net51));
 sg13g2_nor2_1 _2115_ (.A(_0592_),
    .B(net52),
    .Y(_0288_));
 sg13g2_nor2b_1 _2116_ (.A(net46),
    .B_N(_0591_),
    .Y(_0594_));
 sg13g2_a21oi_1 _2117_ (.A1(net46),
    .A2(_0592_),
    .Y(_0289_),
    .B1(_0594_));
 sg13g2_nor2_1 _2118_ (.A(net408),
    .B(net80),
    .Y(_0595_));
 sg13g2_a21oi_1 _2119_ (.A1(net80),
    .A2(_0866_),
    .Y(_0290_),
    .B1(_0595_));
 sg13g2_nand2_1 _2120_ (.Y(_0596_),
    .A(net68),
    .B(_0865_));
 sg13g2_and2_1 _2121_ (.A(\serializer_b.bit_cnt[0] ),
    .B(net68),
    .X(_0597_));
 sg13g2_o21ai_1 _2122_ (.B1(net69),
    .Y(_0291_),
    .A1(_0867_),
    .A2(_0597_));
 sg13g2_nand3_1 _2123_ (.B(net74),
    .C(_0597_),
    .A(net408),
    .Y(_0598_));
 sg13g2_nand2b_1 _2124_ (.Y(_0599_),
    .B(_0598_),
    .A_N(net401));
 sg13g2_a21oi_1 _2125_ (.A1(_0866_),
    .A2(_0597_),
    .Y(_0600_),
    .B1(net74));
 sg13g2_nor2_1 _2126_ (.A(_0599_),
    .B(net75),
    .Y(_0292_));
 sg13g2_nor2b_1 _2127_ (.A(net39),
    .B_N(_0598_),
    .Y(_0601_));
 sg13g2_a21oi_1 _2128_ (.A1(net39),
    .A2(_0599_),
    .Y(_0293_),
    .B1(_0601_));
 sg13g2_nor2b_2 _2129_ (.A(net241),
    .B_N(net181),
    .Y(_0602_));
 sg13g2_nor2b_1 _2130_ (.A(net181),
    .B_N(\cic_a.filtered_out[0] ),
    .Y(_0603_));
 sg13g2_o21ai_1 _2131_ (.B1(_0019_),
    .Y(_0604_),
    .A1(_0602_),
    .A2(_0603_));
 sg13g2_o21ai_1 _2132_ (.B1(_0604_),
    .Y(_0294_),
    .A1(_0710_),
    .A2(_0870_));
 sg13g2_nand2b_1 _2133_ (.Y(_0605_),
    .B(\cic_a.filtered_out[1] ),
    .A_N(\cic_b.filtered_out[1] ));
 sg13g2_xor2_1 _2134_ (.B(net225),
    .A(\cic_a.filtered_out[1] ),
    .X(_0606_));
 sg13g2_xnor2_1 _2135_ (.Y(_0607_),
    .A(_0602_),
    .B(_0606_));
 sg13g2_nor2_1 _2136_ (.A(net307),
    .B(_0870_),
    .Y(_0608_));
 sg13g2_a221oi_1 _2137_ (.B2(_0607_),
    .C1(_0608_),
    .B1(_0019_),
    .A1(net405),
    .Y(_0295_),
    .A2(_0710_));
 sg13g2_nor2b_1 _2138_ (.A(\cic_b.filtered_out[2] ),
    .B_N(\cic_a.filtered_out[2] ),
    .Y(_0609_));
 sg13g2_nand2b_1 _2139_ (.Y(_0610_),
    .B(\cic_b.filtered_out[2] ),
    .A_N(\cic_a.filtered_out[2] ));
 sg13g2_nor2b_1 _2140_ (.A(_0609_),
    .B_N(_0610_),
    .Y(_0611_));
 sg13g2_o21ai_1 _2141_ (.B1(_0605_),
    .Y(_0612_),
    .A1(_0602_),
    .A2(_0606_));
 sg13g2_xnor2_1 _2142_ (.Y(_0613_),
    .A(_0611_),
    .B(_0612_));
 sg13g2_a22oi_1 _2143_ (.Y(_0614_),
    .B1(net155),
    .B2(net399),
    .A2(\serializer_ab_subtr.shift_reg[1] ),
    .A1(net406));
 sg13g2_o21ai_1 _2144_ (.B1(net156),
    .Y(_0296_),
    .A1(_0730_),
    .A2(_0613_));
 sg13g2_a21oi_1 _2145_ (.A1(_0610_),
    .A2(_0612_),
    .Y(_0615_),
    .B1(_0609_));
 sg13g2_nor2_1 _2146_ (.A(\cic_a.filtered_out[3] ),
    .B(_0701_),
    .Y(_0616_));
 sg13g2_xor2_1 _2147_ (.B(\cic_b.filtered_out[3] ),
    .A(\cic_a.filtered_out[3] ),
    .X(_0617_));
 sg13g2_xnor2_1 _2148_ (.Y(_0618_),
    .A(_0615_),
    .B(_0617_));
 sg13g2_a22oi_1 _2149_ (.Y(_0619_),
    .B1(net279),
    .B2(net399),
    .A2(net155),
    .A1(net406));
 sg13g2_o21ai_1 _2150_ (.B1(net280),
    .Y(_0297_),
    .A1(_0730_),
    .A2(_0618_));
 sg13g2_xor2_1 _2151_ (.B(\cic_b.filtered_out[4] ),
    .A(\cic_a.filtered_out[4] ),
    .X(_0620_));
 sg13g2_a221oi_1 _2152_ (.B2(_0612_),
    .C1(_0609_),
    .B1(_0611_),
    .A1(\cic_a.filtered_out[3] ),
    .Y(_0621_),
    .A2(_0701_));
 sg13g2_o21ai_1 _2153_ (.B1(_0620_),
    .Y(_0622_),
    .A1(_0616_),
    .A2(_0621_));
 sg13g2_or3_2 _2154_ (.A(_0616_),
    .B(_0620_),
    .C(_0621_),
    .X(_0623_));
 sg13g2_nand3_1 _2155_ (.B(_0622_),
    .C(_0623_),
    .A(_0019_),
    .Y(_0624_));
 sg13g2_a22oi_1 _2156_ (.Y(_0625_),
    .B1(net503),
    .B2(net398),
    .A2(net279),
    .A1(net407));
 sg13g2_nand2_1 _2157_ (.Y(_0298_),
    .A(_0624_),
    .B(net504));
 sg13g2_nor2_1 _2158_ (.A(\cic_a.filtered_out[5] ),
    .B(_0703_),
    .Y(_0626_));
 sg13g2_xnor2_1 _2159_ (.Y(_0627_),
    .A(\cic_a.filtered_out[5] ),
    .B(\cic_b.filtered_out[5] ));
 sg13g2_o21ai_1 _2160_ (.B1(_0623_),
    .Y(_0628_),
    .A1(_0693_),
    .A2(\cic_b.filtered_out[4] ));
 sg13g2_xnor2_1 _2161_ (.Y(_0629_),
    .A(_0627_),
    .B(_0628_));
 sg13g2_a22oi_1 _2162_ (.Y(_0630_),
    .B1(net186),
    .B2(net398),
    .A2(\serializer_ab_subtr.shift_reg[4] ),
    .A1(net407));
 sg13g2_o21ai_1 _2163_ (.B1(net187),
    .Y(_0299_),
    .A1(net402),
    .A2(_0629_));
 sg13g2_nand2b_1 _2164_ (.Y(_0631_),
    .B(\cic_a.filtered_out[6] ),
    .A_N(\cic_b.filtered_out[6] ));
 sg13g2_xnor2_1 _2165_ (.Y(_0632_),
    .A(\cic_a.filtered_out[6] ),
    .B(\cic_b.filtered_out[6] ));
 sg13g2_inv_1 _2166_ (.Y(_0633_),
    .A(_0632_));
 sg13g2_a22oi_1 _2167_ (.Y(_0634_),
    .B1(_0703_),
    .B2(\cic_a.filtered_out[5] ),
    .A2(_0702_),
    .A1(\cic_a.filtered_out[4] ));
 sg13g2_a21oi_1 _2168_ (.A1(_0623_),
    .A2(_0634_),
    .Y(_0635_),
    .B1(_0626_));
 sg13g2_nand2_1 _2169_ (.Y(_0636_),
    .A(_0632_),
    .B(_0635_));
 sg13g2_xnor2_1 _2170_ (.Y(_0637_),
    .A(_0632_),
    .B(_0635_));
 sg13g2_a22oi_1 _2171_ (.Y(_0638_),
    .B1(net167),
    .B2(net398),
    .A2(\serializer_ab_subtr.shift_reg[5] ),
    .A1(net407));
 sg13g2_o21ai_1 _2172_ (.B1(net168),
    .Y(_0300_),
    .A1(net402),
    .A2(_0637_));
 sg13g2_nand2_1 _2173_ (.Y(_0639_),
    .A(_0631_),
    .B(_0636_));
 sg13g2_nand2_1 _2174_ (.Y(_0640_),
    .A(_0695_),
    .B(\cic_b.filtered_out[7] ));
 sg13g2_xor2_1 _2175_ (.B(\cic_b.filtered_out[7] ),
    .A(\cic_a.filtered_out[7] ),
    .X(_0641_));
 sg13g2_xor2_1 _2176_ (.B(_0641_),
    .A(_0639_),
    .X(_0642_));
 sg13g2_a22oi_1 _2177_ (.Y(_0643_),
    .B1(net182),
    .B2(net398),
    .A2(net167),
    .A1(net407));
 sg13g2_o21ai_1 _2178_ (.B1(net183),
    .Y(_0301_),
    .A1(net402),
    .A2(_0642_));
 sg13g2_nor2_1 _2179_ (.A(_0633_),
    .B(_0641_),
    .Y(_0644_));
 sg13g2_nand2_1 _2180_ (.Y(_0645_),
    .A(_0627_),
    .B(_0644_));
 sg13g2_nor2_1 _2181_ (.A(_0626_),
    .B(_0634_),
    .Y(_0646_));
 sg13g2_o21ai_1 _2182_ (.B1(_0631_),
    .Y(_0647_),
    .A1(_0695_),
    .A2(\cic_b.filtered_out[7] ));
 sg13g2_a22oi_1 _2183_ (.Y(_0648_),
    .B1(_0647_),
    .B2(_0640_),
    .A2(_0646_),
    .A1(_0644_));
 sg13g2_o21ai_1 _2184_ (.B1(_0648_),
    .Y(_0649_),
    .A1(_0623_),
    .A2(_0645_));
 sg13g2_nand2b_1 _2185_ (.Y(_0650_),
    .B(\cic_a.filtered_out[8] ),
    .A_N(\cic_b.filtered_out[8] ));
 sg13g2_xnor2_1 _2186_ (.Y(_0651_),
    .A(\cic_a.filtered_out[8] ),
    .B(\cic_b.filtered_out[8] ));
 sg13g2_nand2_1 _2187_ (.Y(_0652_),
    .A(_0649_),
    .B(_0651_));
 sg13g2_nor2_1 _2188_ (.A(_0649_),
    .B(_0651_),
    .Y(_0653_));
 sg13g2_nand2_1 _2189_ (.Y(_0654_),
    .A(_0019_),
    .B(_0652_));
 sg13g2_a22oi_1 _2190_ (.Y(_0655_),
    .B1(net159),
    .B2(net398),
    .A2(\serializer_ab_subtr.shift_reg[7] ),
    .A1(net407));
 sg13g2_o21ai_1 _2191_ (.B1(net160),
    .Y(_0302_),
    .A1(_0653_),
    .A2(_0654_));
 sg13g2_nand2b_1 _2192_ (.Y(_0656_),
    .B(\cic_a.filtered_out[9] ),
    .A_N(\cic_b.filtered_out[9] ));
 sg13g2_nor2b_1 _2193_ (.A(\cic_a.filtered_out[9] ),
    .B_N(\cic_b.filtered_out[9] ),
    .Y(_0657_));
 sg13g2_xnor2_1 _2194_ (.Y(_0658_),
    .A(\cic_a.filtered_out[9] ),
    .B(\cic_b.filtered_out[9] ));
 sg13g2_nand2_1 _2195_ (.Y(_0659_),
    .A(_0650_),
    .B(_0652_));
 sg13g2_xnor2_1 _2196_ (.Y(_0660_),
    .A(_0658_),
    .B(_0659_));
 sg13g2_a22oi_1 _2197_ (.Y(_0661_),
    .B1(net523),
    .B2(net398),
    .A2(net159),
    .A1(net407));
 sg13g2_o21ai_1 _2198_ (.B1(net524),
    .Y(_0303_),
    .A1(net402),
    .A2(_0660_));
 sg13g2_and2_1 _2199_ (.A(_0651_),
    .B(_0658_),
    .X(_0662_));
 sg13g2_o21ai_1 _2200_ (.B1(_0656_),
    .Y(_0663_),
    .A1(_0650_),
    .A2(_0657_));
 sg13g2_a21o_2 _2201_ (.A2(_0662_),
    .A1(_0649_),
    .B1(_0663_),
    .X(_0664_));
 sg13g2_nor2b_1 _2202_ (.A(\cic_b.filtered_out[10] ),
    .B_N(\cic_a.filtered_out[10] ),
    .Y(_0665_));
 sg13g2_xnor2_1 _2203_ (.Y(_0666_),
    .A(\cic_a.filtered_out[10] ),
    .B(\cic_b.filtered_out[10] ));
 sg13g2_inv_1 _2204_ (.Y(_0667_),
    .A(_0666_));
 sg13g2_a21oi_1 _2205_ (.A1(_0664_),
    .A2(_0666_),
    .Y(_0668_),
    .B1(net402));
 sg13g2_o21ai_1 _2206_ (.B1(_0668_),
    .Y(_0669_),
    .A1(_0664_),
    .A2(_0666_));
 sg13g2_a22oi_1 _2207_ (.Y(_0670_),
    .B1(net350),
    .B2(net398),
    .A2(\serializer_ab_subtr.shift_reg[9] ),
    .A1(net407));
 sg13g2_nand2_1 _2208_ (.Y(_0304_),
    .A(_0669_),
    .B(net351));
 sg13g2_nor2b_1 _2209_ (.A(\cic_b.filtered_out[11] ),
    .B_N(\cic_a.filtered_out[11] ),
    .Y(_0671_));
 sg13g2_nand2b_1 _2210_ (.Y(_0672_),
    .B(\cic_b.filtered_out[11] ),
    .A_N(\cic_a.filtered_out[11] ));
 sg13g2_nand2b_1 _2211_ (.Y(_0673_),
    .B(_0672_),
    .A_N(_0671_));
 sg13g2_a21oi_1 _2212_ (.A1(_0664_),
    .A2(_0666_),
    .Y(_0674_),
    .B1(_0665_));
 sg13g2_xnor2_1 _2213_ (.Y(_0675_),
    .A(_0673_),
    .B(_0674_));
 sg13g2_a22oi_1 _2214_ (.Y(_0676_),
    .B1(net489),
    .B2(net398),
    .A2(net350),
    .A1(net407));
 sg13g2_o21ai_1 _2215_ (.B1(net490),
    .Y(_0305_),
    .A1(net402),
    .A2(_0675_));
 sg13g2_nor2_1 _2216_ (.A(_0667_),
    .B(_0673_),
    .Y(_0677_));
 sg13g2_a221oi_1 _2217_ (.B2(_0664_),
    .C1(_0671_),
    .B1(_0677_),
    .A1(_0665_),
    .Y(_0678_),
    .A2(_0672_));
 sg13g2_xor2_1 _2218_ (.B(\cic_b.filtered_out[12] ),
    .A(\cic_a.filtered_out[12] ),
    .X(_0679_));
 sg13g2_xnor2_1 _2219_ (.Y(_0680_),
    .A(_0678_),
    .B(_0679_));
 sg13g2_a22oi_1 _2220_ (.Y(_0681_),
    .B1(net151),
    .B2(net399),
    .A2(\serializer_ab_subtr.shift_reg[11] ),
    .A1(net405));
 sg13g2_o21ai_1 _2221_ (.B1(net152),
    .Y(_0306_),
    .A1(_0730_),
    .A2(_0680_));
 sg13g2_nor2_1 _2222_ (.A(net411),
    .B(net96),
    .Y(_0682_));
 sg13g2_a21oi_1 _2223_ (.A1(net96),
    .A2(net397),
    .Y(_0307_),
    .B1(_0682_));
 sg13g2_nand2_1 _2224_ (.Y(_0683_),
    .A(net105),
    .B(_0861_));
 sg13g2_and2_1 _2225_ (.A(net96),
    .B(net105),
    .X(_0684_));
 sg13g2_o21ai_1 _2226_ (.B1(_0683_),
    .Y(_0308_),
    .A1(_0863_),
    .A2(_0684_));
 sg13g2_nand3_1 _2227_ (.B(net161),
    .C(_0684_),
    .A(net411),
    .Y(_0685_));
 sg13g2_nand2b_1 _2228_ (.Y(_0686_),
    .B(_0685_),
    .A_N(net404));
 sg13g2_a21oi_1 _2229_ (.A1(net397),
    .A2(_0684_),
    .Y(_0687_),
    .B1(net161));
 sg13g2_nor2_1 _2230_ (.A(_0686_),
    .B(_0687_),
    .Y(_0309_));
 sg13g2_nor2b_1 _2231_ (.A(net55),
    .B_N(_0685_),
    .Y(_0688_));
 sg13g2_a21oi_1 _2232_ (.A1(net55),
    .A2(_0686_),
    .Y(_0310_),
    .B1(_0688_));
 sg13g2_dfrbp_1 _2233_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net466),
    .D(_0076_),
    .Q_N(\cic_a.pdm_in ),
    .Q(_0074_));
 sg13g2_dfrbp_1 _2234_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net452),
    .D(_0077_),
    .Q_N(\cic_b.pdm_in ),
    .Q(_0075_));
 sg13g2_dfrbp_1 _2235_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net458),
    .D(net256),
    .Q_N(_1195_),
    .Q(\cic_a.delay[0][0] ));
 sg13g2_dfrbp_1 _2236_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net458),
    .D(net204),
    .Q_N(_1194_),
    .Q(\cic_a.delay[0][1] ));
 sg13g2_dfrbp_1 _2237_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net437),
    .D(_0080_),
    .Q_N(_1193_),
    .Q(\cic_a.delay[0][2] ));
 sg13g2_dfrbp_1 _2238_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net437),
    .D(net243),
    .Q_N(_1192_),
    .Q(\cic_a.delay[0][3] ));
 sg13g2_dfrbp_1 _2239_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net430),
    .D(_0082_),
    .Q_N(_1191_),
    .Q(\cic_a.delay[0][4] ));
 sg13g2_dfrbp_1 _2240_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net430),
    .D(net67),
    .Q_N(_1190_),
    .Q(\cic_a.delay[0][5] ));
 sg13g2_dfrbp_1 _2241_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net430),
    .D(net197),
    .Q_N(_1189_),
    .Q(\cic_a.delay[0][6] ));
 sg13g2_dfrbp_1 _2242_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net430),
    .D(net174),
    .Q_N(_1188_),
    .Q(\cic_a.delay[0][7] ));
 sg13g2_dfrbp_1 _2243_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net428),
    .D(net176),
    .Q_N(_1187_),
    .Q(\cic_a.delay[0][8] ));
 sg13g2_dfrbp_1 _2244_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net425),
    .D(_0087_),
    .Q_N(_1186_),
    .Q(\cic_a.delay[0][9] ));
 sg13g2_dfrbp_1 _2245_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net427),
    .D(_0088_),
    .Q_N(_1185_),
    .Q(\cic_a.delay[0][10] ));
 sg13g2_dfrbp_1 _2246_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net426),
    .D(_0089_),
    .Q_N(_1184_),
    .Q(\cic_a.delay[0][11] ));
 sg13g2_dfrbp_1 _2247_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net426),
    .D(net170),
    .Q_N(_1183_),
    .Q(\cic_a.delay[0][12] ));
 sg13g2_dfrbp_1 _2248_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net460),
    .D(_0091_),
    .Q_N(_1182_),
    .Q(\cic_a.temp_comb[0][0] ));
 sg13g2_dfrbp_1 _2249_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net461),
    .D(_0092_),
    .Q_N(_1181_),
    .Q(\cic_a.temp_comb[0][1] ));
 sg13g2_dfrbp_1 _2250_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net459),
    .D(net555),
    .Q_N(_1180_),
    .Q(\cic_a.temp_comb[0][2] ));
 sg13g2_dfrbp_1 _2251_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net436),
    .D(_0094_),
    .Q_N(_1179_),
    .Q(\cic_a.temp_comb[0][3] ));
 sg13g2_dfrbp_1 _2252_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net435),
    .D(_0095_),
    .Q_N(_1178_),
    .Q(\cic_a.temp_comb[0][4] ));
 sg13g2_dfrbp_1 _2253_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net435),
    .D(net531),
    .Q_N(_1177_),
    .Q(\cic_a.temp_comb[0][5] ));
 sg13g2_dfrbp_1 _2254_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net435),
    .D(_0097_),
    .Q_N(_1176_),
    .Q(\cic_a.temp_comb[0][6] ));
 sg13g2_dfrbp_1 _2255_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net435),
    .D(_0098_),
    .Q_N(_1175_),
    .Q(\cic_a.temp_comb[0][7] ));
 sg13g2_dfrbp_1 _2256_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net427),
    .D(_0099_),
    .Q_N(_1174_),
    .Q(\cic_a.temp_comb[0][8] ));
 sg13g2_dfrbp_1 _2257_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net427),
    .D(_0100_),
    .Q_N(_1173_),
    .Q(\cic_a.temp_comb[0][9] ));
 sg13g2_dfrbp_1 _2258_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net427),
    .D(_0101_),
    .Q_N(_1172_),
    .Q(\cic_a.temp_comb[0][10] ));
 sg13g2_dfrbp_1 _2259_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net427),
    .D(_0102_),
    .Q_N(_1171_),
    .Q(\cic_a.temp_comb[0][11] ));
 sg13g2_dfrbp_1 _2260_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net427),
    .D(net199),
    .Q_N(_1170_),
    .Q(\cic_a.temp_comb[0][12] ));
 sg13g2_dfrbp_1 _2261_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net465),
    .D(_0104_),
    .Q_N(_1169_),
    .Q(\cic_a.filtered_out[0] ));
 sg13g2_dfrbp_1 _2262_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net465),
    .D(_0105_),
    .Q_N(_1168_),
    .Q(\cic_a.filtered_out[1] ));
 sg13g2_dfrbp_1 _2263_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net465),
    .D(_0106_),
    .Q_N(_1167_),
    .Q(\cic_a.filtered_out[2] ));
 sg13g2_dfrbp_1 _2264_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net465),
    .D(_0107_),
    .Q_N(_1166_),
    .Q(\cic_a.filtered_out[3] ));
 sg13g2_dfrbp_1 _2265_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net456),
    .D(net127),
    .Q_N(_1165_),
    .Q(\cic_a.filtered_out[4] ));
 sg13g2_dfrbp_1 _2266_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net459),
    .D(_0109_),
    .Q_N(_1164_),
    .Q(\cic_a.filtered_out[5] ));
 sg13g2_dfrbp_1 _2267_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net457),
    .D(_0110_),
    .Q_N(_1163_),
    .Q(\cic_a.filtered_out[6] ));
 sg13g2_dfrbp_1 _2268_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net457),
    .D(_0111_),
    .Q_N(_1162_),
    .Q(\cic_a.filtered_out[7] ));
 sg13g2_dfrbp_1 _2269_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net457),
    .D(_0112_),
    .Q_N(_1161_),
    .Q(\cic_a.filtered_out[8] ));
 sg13g2_dfrbp_1 _2270_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net433),
    .D(_0113_),
    .Q_N(_1160_),
    .Q(\cic_a.filtered_out[9] ));
 sg13g2_dfrbp_1 _2271_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net433),
    .D(_0114_),
    .Q_N(_1159_),
    .Q(\cic_a.filtered_out[10] ));
 sg13g2_dfrbp_1 _2272_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net433),
    .D(_0115_),
    .Q_N(_1158_),
    .Q(\cic_a.filtered_out[11] ));
 sg13g2_dfrbp_1 _2273_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net433),
    .D(_0116_),
    .Q_N(_1196_),
    .Q(\cic_a.filtered_out[12] ));
 sg13g2_dfrbp_1 _2274_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net458),
    .D(net515),
    .Q_N(_1197_),
    .Q(\cic_a.integrator[1][0] ));
 sg13g2_dfrbp_1 _2275_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net458),
    .D(net567),
    .Q_N(_1198_),
    .Q(\cic_a.integrator[1][1] ));
 sg13g2_dfrbp_1 _2276_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net436),
    .D(_0040_),
    .Q_N(_1199_),
    .Q(\cic_a.integrator[1][2] ));
 sg13g2_dfrbp_1 _2277_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net437),
    .D(_0041_),
    .Q_N(_1200_),
    .Q(\cic_a.integrator[1][3] ));
 sg13g2_dfrbp_1 _2278_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net430),
    .D(net606),
    .Q_N(_1201_),
    .Q(\cic_a.integrator[1][4] ));
 sg13g2_dfrbp_1 _2279_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net429),
    .D(net591),
    .Q_N(_1202_),
    .Q(\cic_a.integrator[1][5] ));
 sg13g2_dfrbp_1 _2280_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net429),
    .D(_0044_),
    .Q_N(_1203_),
    .Q(\cic_a.integrator[1][6] ));
 sg13g2_dfrbp_1 _2281_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net428),
    .D(net603),
    .Q_N(_1204_),
    .Q(\cic_a.integrator[1][7] ));
 sg13g2_dfrbp_1 _2282_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net428),
    .D(_0046_),
    .Q_N(_1205_),
    .Q(\cic_a.integrator[1][8] ));
 sg13g2_dfrbp_1 _2283_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net425),
    .D(net579),
    .Q_N(_1206_),
    .Q(\cic_a.integrator[1][9] ));
 sg13g2_dfrbp_1 _2284_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net425),
    .D(net595),
    .Q_N(_1207_),
    .Q(\cic_a.integrator[1][10] ));
 sg13g2_dfrbp_1 _2285_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net425),
    .D(net593),
    .Q_N(_1208_),
    .Q(\cic_a.integrator[1][11] ));
 sg13g2_dfrbp_1 _2286_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net426),
    .D(net565),
    .Q_N(_1157_),
    .Q(\cic_a.integrator[1][12] ));
 sg13g2_dfrbp_1 _2287_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net465),
    .D(net292),
    .Q_N(_1156_),
    .Q(\cic_a.delay[1][0] ));
 sg13g2_dfrbp_1 _2288_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net460),
    .D(_0118_),
    .Q_N(_1155_),
    .Q(\cic_a.delay[1][1] ));
 sg13g2_dfrbp_1 _2289_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net460),
    .D(_0119_),
    .Q_N(_1154_),
    .Q(\cic_a.delay[1][2] ));
 sg13g2_dfrbp_1 _2290_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net459),
    .D(_0120_),
    .Q_N(_1153_),
    .Q(\cic_a.delay[1][3] ));
 sg13g2_dfrbp_1 _2291_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net436),
    .D(_0121_),
    .Q_N(_1152_),
    .Q(\cic_a.delay[1][4] ));
 sg13g2_dfrbp_1 _2292_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net436),
    .D(_0122_),
    .Q_N(_1151_),
    .Q(\cic_a.delay[1][5] ));
 sg13g2_dfrbp_1 _2293_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net435),
    .D(_0123_),
    .Q_N(_1150_),
    .Q(\cic_a.delay[1][6] ));
 sg13g2_dfrbp_1 _2294_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net435),
    .D(net158),
    .Q_N(_1149_),
    .Q(\cic_a.delay[1][7] ));
 sg13g2_dfrbp_1 _2295_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net434),
    .D(net266),
    .Q_N(_1148_),
    .Q(\cic_a.delay[1][8] ));
 sg13g2_dfrbp_1 _2296_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net434),
    .D(_0126_),
    .Q_N(_1147_),
    .Q(\cic_a.delay[1][9] ));
 sg13g2_dfrbp_1 _2297_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net434),
    .D(net216),
    .Q_N(_1146_),
    .Q(\cic_a.delay[1][10] ));
 sg13g2_dfrbp_1 _2298_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net434),
    .D(net320),
    .Q_N(_1145_),
    .Q(\cic_a.delay[1][11] ));
 sg13g2_dfrbp_1 _2299_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net432),
    .D(net237),
    .Q_N(_1209_),
    .Q(\cic_a.delay[1][12] ));
 sg13g2_dfrbp_1 _2300_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net458),
    .D(net32),
    .Q_N(_1210_),
    .Q(\cic_a.integrator[0][0] ));
 sg13g2_dfrbp_1 _2301_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net458),
    .D(_0026_),
    .Q_N(_1211_),
    .Q(\cic_a.integrator[0][1] ));
 sg13g2_dfrbp_1 _2302_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net436),
    .D(net229),
    .Q_N(_1212_),
    .Q(\cic_a.integrator[0][2] ));
 sg13g2_dfrbp_1 _2303_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net430),
    .D(_0028_),
    .Q_N(_1213_),
    .Q(\cic_a.integrator[0][3] ));
 sg13g2_dfrbp_1 _2304_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net430),
    .D(_0029_),
    .Q_N(_1214_),
    .Q(\cic_a.integrator[0][4] ));
 sg13g2_dfrbp_1 _2305_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net429),
    .D(net501),
    .Q_N(_1215_),
    .Q(\cic_a.integrator[0][5] ));
 sg13g2_dfrbp_1 _2306_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net429),
    .D(net553),
    .Q_N(_1216_),
    .Q(\cic_a.integrator[0][6] ));
 sg13g2_dfrbp_1 _2307_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net428),
    .D(net535),
    .Q_N(_1217_),
    .Q(\cic_a.integrator[0][7] ));
 sg13g2_dfrbp_1 _2308_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net428),
    .D(_0033_),
    .Q_N(_1218_),
    .Q(\cic_a.integrator[0][8] ));
 sg13g2_dfrbp_1 _2309_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net425),
    .D(net543),
    .Q_N(_1219_),
    .Q(\cic_a.integrator[0][9] ));
 sg13g2_dfrbp_1 _2310_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net425),
    .D(_0023_),
    .Q_N(_1220_),
    .Q(\cic_a.integrator[0][10] ));
 sg13g2_dfrbp_1 _2311_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net425),
    .D(_0024_),
    .Q_N(_1221_),
    .Q(\cic_a.integrator[0][11] ));
 sg13g2_dfrbp_1 _2312_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net426),
    .D(net140),
    .Q_N(_1144_),
    .Q(\cic_a.integrator[0][12] ));
 sg13g2_dfrbp_1 _2313_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net466),
    .D(net100),
    .Q_N(_1143_),
    .Q(\cic_a.temp_comb[1][0] ));
 sg13g2_dfrbp_1 _2314_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net465),
    .D(net195),
    .Q_N(_1142_),
    .Q(\cic_a.temp_comb[1][1] ));
 sg13g2_dfrbp_1 _2315_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net465),
    .D(_0132_),
    .Q_N(_1141_),
    .Q(\cic_a.temp_comb[1][2] ));
 sg13g2_dfrbp_1 _2316_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net460),
    .D(net163),
    .Q_N(_1140_),
    .Q(\cic_a.temp_comb[1][3] ));
 sg13g2_dfrbp_1 _2317_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net457),
    .D(_0134_),
    .Q_N(_1139_),
    .Q(\cic_a.temp_comb[1][4] ));
 sg13g2_dfrbp_1 _2318_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net459),
    .D(_0135_),
    .Q_N(_1138_),
    .Q(\cic_a.temp_comb[1][5] ));
 sg13g2_dfrbp_1 _2319_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net438),
    .D(_0136_),
    .Q_N(_1137_),
    .Q(\cic_a.temp_comb[1][6] ));
 sg13g2_dfrbp_1 _2320_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net438),
    .D(_0137_),
    .Q_N(_1136_),
    .Q(\cic_a.temp_comb[1][7] ));
 sg13g2_dfrbp_1 _2321_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net433),
    .D(_0138_),
    .Q_N(_1135_),
    .Q(\cic_a.temp_comb[1][8] ));
 sg13g2_dfrbp_1 _2322_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net433),
    .D(_0139_),
    .Q_N(_1134_),
    .Q(\cic_a.temp_comb[1][9] ));
 sg13g2_dfrbp_1 _2323_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net433),
    .D(_0140_),
    .Q_N(_1133_),
    .Q(\cic_a.temp_comb[1][10] ));
 sg13g2_dfrbp_1 _2324_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net433),
    .D(_0141_),
    .Q_N(_1132_),
    .Q(\cic_a.temp_comb[1][11] ));
 sg13g2_dfrbp_1 _2325_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net434),
    .D(net104),
    .Q_N(_1222_),
    .Q(\cic_a.temp_comb[1][12] ));
 sg13g2_dfrbp_1 _2326_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net416),
    .D(_0000_),
    .Q_N(_1223_),
    .Q(\cic_a.decim_cnt[0] ));
 sg13g2_dfrbp_1 _2327_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net417),
    .D(_0001_),
    .Q_N(_1224_),
    .Q(\cic_a.decim_cnt[1] ));
 sg13g2_dfrbp_1 _2328_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net417),
    .D(_0002_),
    .Q_N(_1225_),
    .Q(\cic_a.decim_cnt[2] ));
 sg13g2_dfrbp_1 _2329_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net417),
    .D(net50),
    .Q_N(_1226_),
    .Q(\cic_a.decim_cnt[3] ));
 sg13g2_dfrbp_1 _2330_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net416),
    .D(net36),
    .Q_N(_1227_),
    .Q(\cic_a.decim_cnt[4] ));
 sg13g2_dfrbp_1 _2331_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net416),
    .D(_0005_),
    .Q_N(_1228_),
    .Q(\cic_a.decim_cnt[5] ));
 sg13g2_dfrbp_1 _2332_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net418),
    .D(_0006_),
    .Q_N(_1229_),
    .Q(\cic_a.decim_cnt[6] ));
 sg13g2_dfrbp_1 _2333_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net418),
    .D(net178),
    .Q_N(_1131_),
    .Q(\cic_a.decim_cnt[7] ));
 sg13g2_dfrbp_1 _2334_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net458),
    .D(net272),
    .Q_N(_1130_),
    .Q(\cic_a.temp_delay[0][0] ));
 sg13g2_dfrbp_1 _2335_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net458),
    .D(_0144_),
    .Q_N(_1129_),
    .Q(\cic_a.temp_delay[0][1] ));
 sg13g2_dfrbp_1 _2336_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net436),
    .D(net286),
    .Q_N(_1128_),
    .Q(\cic_a.temp_delay[0][2] ));
 sg13g2_dfrbp_1 _2337_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net437),
    .D(_0146_),
    .Q_N(_1127_),
    .Q(\cic_a.temp_delay[0][3] ));
 sg13g2_dfrbp_1 _2338_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net430),
    .D(net330),
    .Q_N(_1126_),
    .Q(\cic_a.temp_delay[0][4] ));
 sg13g2_dfrbp_1 _2339_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net431),
    .D(_0148_),
    .Q_N(_1125_),
    .Q(\cic_a.temp_delay[0][5] ));
 sg13g2_dfrbp_1 _2340_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net428),
    .D(_0149_),
    .Q_N(_1124_),
    .Q(\cic_a.temp_delay[0][6] ));
 sg13g2_dfrbp_1 _2341_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net428),
    .D(_0150_),
    .Q_N(_1123_),
    .Q(\cic_a.temp_delay[0][7] ));
 sg13g2_dfrbp_1 _2342_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net428),
    .D(net469),
    .Q_N(_1122_),
    .Q(\cic_a.temp_delay[0][8] ));
 sg13g2_dfrbp_1 _2343_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net425),
    .D(net93),
    .Q_N(_1121_),
    .Q(\cic_a.temp_delay[0][9] ));
 sg13g2_dfrbp_1 _2344_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net426),
    .D(net314),
    .Q_N(_1120_),
    .Q(\cic_a.temp_delay[0][10] ));
 sg13g2_dfrbp_1 _2345_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net426),
    .D(net245),
    .Q_N(_1119_),
    .Q(\cic_a.temp_delay[0][11] ));
 sg13g2_dfrbp_1 _2346_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net426),
    .D(net482),
    .Q_N(_1118_),
    .Q(\cic_a.temp_delay[0][12] ));
 sg13g2_dfrbp_1 _2347_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net448),
    .D(net206),
    .Q_N(_1117_),
    .Q(\cic_b.delay[0][0] ));
 sg13g2_dfrbp_1 _2348_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net448),
    .D(net316),
    .Q_N(_1116_),
    .Q(\cic_b.delay[0][1] ));
 sg13g2_dfrbp_1 _2349_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net447),
    .D(net227),
    .Q_N(_1115_),
    .Q(\cic_b.delay[0][2] ));
 sg13g2_dfrbp_1 _2350_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net441),
    .D(net296),
    .Q_N(_1114_),
    .Q(\cic_b.delay[0][3] ));
 sg13g2_dfrbp_1 _2351_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net440),
    .D(net218),
    .Q_N(_1113_),
    .Q(\cic_b.delay[0][4] ));
 sg13g2_dfrbp_1 _2352_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net440),
    .D(net147),
    .Q_N(_1112_),
    .Q(\cic_b.delay[0][5] ));
 sg13g2_dfrbp_1 _2353_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net424),
    .D(net224),
    .Q_N(_1111_),
    .Q(\cic_b.delay[0][6] ));
 sg13g2_dfrbp_1 _2354_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net419),
    .D(net231),
    .Q_N(_1110_),
    .Q(\cic_b.delay[0][7] ));
 sg13g2_dfrbp_1 _2355_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net420),
    .D(net102),
    .Q_N(_1109_),
    .Q(\cic_b.delay[0][8] ));
 sg13g2_dfrbp_1 _2356_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net420),
    .D(net88),
    .Q_N(_1108_),
    .Q(\cic_b.delay[0][9] ));
 sg13g2_dfrbp_1 _2357_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net413),
    .D(net249),
    .Q_N(_1107_),
    .Q(\cic_b.delay[0][10] ));
 sg13g2_dfrbp_1 _2358_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net414),
    .D(net210),
    .Q_N(_1106_),
    .Q(\cic_b.delay[0][11] ));
 sg13g2_dfrbp_1 _2359_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net413),
    .D(net193),
    .Q_N(_1105_),
    .Q(\cic_b.delay[0][12] ));
 sg13g2_dfrbp_1 _2360_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net449),
    .D(net529),
    .Q_N(_1104_),
    .Q(\cic_b.temp_comb[0][0] ));
 sg13g2_dfrbp_1 _2361_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net449),
    .D(_0170_),
    .Q_N(_1103_),
    .Q(\cic_b.temp_comb[0][1] ));
 sg13g2_dfrbp_1 _2362_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net447),
    .D(_0171_),
    .Q_N(_1102_),
    .Q(\cic_b.temp_comb[0][2] ));
 sg13g2_dfrbp_1 _2363_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net441),
    .D(_0172_),
    .Q_N(_1101_),
    .Q(\cic_b.temp_comb[0][3] ));
 sg13g2_dfrbp_1 _2364_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net442),
    .D(_0173_),
    .Q_N(_1100_),
    .Q(\cic_b.temp_comb[0][4] ));
 sg13g2_dfrbp_1 _2365_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net441),
    .D(net541),
    .Q_N(_1099_),
    .Q(\cic_b.temp_comb[0][5] ));
 sg13g2_dfrbp_1 _2366_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net441),
    .D(_0175_),
    .Q_N(_1098_),
    .Q(\cic_b.temp_comb[0][6] ));
 sg13g2_dfrbp_1 _2367_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net441),
    .D(net497),
    .Q_N(_1097_),
    .Q(\cic_b.temp_comb[0][7] ));
 sg13g2_dfrbp_1 _2368_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net424),
    .D(_0177_),
    .Q_N(_1096_),
    .Q(\cic_b.temp_comb[0][8] ));
 sg13g2_dfrbp_1 _2369_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net421),
    .D(net475),
    .Q_N(_1095_),
    .Q(\cic_b.temp_comb[0][9] ));
 sg13g2_dfrbp_1 _2370_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net422),
    .D(_0179_),
    .Q_N(_1094_),
    .Q(\cic_b.temp_comb[0][10] ));
 sg13g2_dfrbp_1 _2371_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net417),
    .D(net202),
    .Q_N(_1093_),
    .Q(\cic_b.temp_comb[0][11] ));
 sg13g2_dfrbp_1 _2372_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net418),
    .D(net208),
    .Q_N(_1092_),
    .Q(\cic_b.temp_comb[0][12] ));
 sg13g2_dfrbp_1 _2373_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net452),
    .D(_0182_),
    .Q_N(_1091_),
    .Q(\cic_b.filtered_out[0] ));
 sg13g2_dfrbp_1 _2374_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net452),
    .D(_0183_),
    .Q_N(_1090_),
    .Q(\cic_b.filtered_out[1] ));
 sg13g2_dfrbp_1 _2375_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net452),
    .D(_0184_),
    .Q_N(_1089_),
    .Q(\cic_b.filtered_out[2] ));
 sg13g2_dfrbp_1 _2376_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net454),
    .D(net79),
    .Q_N(_1088_),
    .Q(\cic_b.filtered_out[3] ));
 sg13g2_dfrbp_1 _2377_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net443),
    .D(net95),
    .Q_N(_1087_),
    .Q(\cic_b.filtered_out[4] ));
 sg13g2_dfrbp_1 _2378_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net443),
    .D(_0187_),
    .Q_N(_1086_),
    .Q(\cic_b.filtered_out[5] ));
 sg13g2_dfrbp_1 _2379_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net445),
    .D(_0188_),
    .Q_N(_1085_),
    .Q(\cic_b.filtered_out[6] ));
 sg13g2_dfrbp_1 _2380_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net445),
    .D(_0189_),
    .Q_N(_1084_),
    .Q(\cic_b.filtered_out[7] ));
 sg13g2_dfrbp_1 _2381_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net445),
    .D(_0190_),
    .Q_N(_1083_),
    .Q(\cic_b.filtered_out[8] ));
 sg13g2_dfrbp_1 _2382_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net421),
    .D(_0191_),
    .Q_N(_1082_),
    .Q(\cic_b.filtered_out[9] ));
 sg13g2_dfrbp_1 _2383_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net421),
    .D(_0192_),
    .Q_N(_1081_),
    .Q(\cic_b.filtered_out[10] ));
 sg13g2_dfrbp_1 _2384_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net421),
    .D(_0193_),
    .Q_N(_1080_),
    .Q(\cic_b.filtered_out[11] ));
 sg13g2_dfrbp_1 _2385_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net422),
    .D(_0194_),
    .Q_N(_1230_),
    .Q(\cic_b.filtered_out[12] ));
 sg13g2_dfrbp_1 _2386_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net448),
    .D(net526),
    .Q_N(_1231_),
    .Q(\cic_b.integrator[1][0] ));
 sg13g2_dfrbp_1 _2387_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net448),
    .D(net571),
    .Q_N(_1232_),
    .Q(\cic_b.integrator[1][1] ));
 sg13g2_dfrbp_1 _2388_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net447),
    .D(net610),
    .Q_N(_1233_),
    .Q(\cic_b.integrator[1][2] ));
 sg13g2_dfrbp_1 _2389_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net441),
    .D(net589),
    .Q_N(_1234_),
    .Q(\cic_b.integrator[1][3] ));
 sg13g2_dfrbp_1 _2390_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net440),
    .D(net598),
    .Q_N(_1235_),
    .Q(\cic_b.integrator[1][4] ));
 sg13g2_dfrbp_1 _2391_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net440),
    .D(_0069_),
    .Q_N(_1236_),
    .Q(\cic_b.integrator[1][5] ));
 sg13g2_dfrbp_1 _2392_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net419),
    .D(_0070_),
    .Q_N(_1237_),
    .Q(\cic_b.integrator[1][6] ));
 sg13g2_dfrbp_1 _2393_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net419),
    .D(_0071_),
    .Q_N(_1238_),
    .Q(\cic_b.integrator[1][7] ));
 sg13g2_dfrbp_1 _2394_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net420),
    .D(_0072_),
    .Q_N(_1239_),
    .Q(\cic_b.integrator[1][8] ));
 sg13g2_dfrbp_1 _2395_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net420),
    .D(_0073_),
    .Q_N(_1240_),
    .Q(\cic_b.integrator[1][9] ));
 sg13g2_dfrbp_1 _2396_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net413),
    .D(_0062_),
    .Q_N(_1241_),
    .Q(\cic_b.integrator[1][10] ));
 sg13g2_dfrbp_1 _2397_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net413),
    .D(_0063_),
    .Q_N(_1242_),
    .Q(\cic_b.integrator[1][11] ));
 sg13g2_dfrbp_1 _2398_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net413),
    .D(net559),
    .Q_N(_1079_),
    .Q(\cic_b.integrator[1][12] ));
 sg13g2_dfrbp_1 _2399_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net449),
    .D(net254),
    .Q_N(_1078_),
    .Q(\cic_b.delay[1][0] ));
 sg13g2_dfrbp_1 _2400_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net449),
    .D(net262),
    .Q_N(_1077_),
    .Q(\cic_b.delay[1][1] ));
 sg13g2_dfrbp_1 _2401_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net450),
    .D(net276),
    .Q_N(_1076_),
    .Q(\cic_b.delay[1][2] ));
 sg13g2_dfrbp_1 _2402_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net447),
    .D(_0198_),
    .Q_N(_1075_),
    .Q(\cic_b.delay[1][3] ));
 sg13g2_dfrbp_1 _2403_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net442),
    .D(_0199_),
    .Q_N(_1074_),
    .Q(\cic_b.delay[1][4] ));
 sg13g2_dfrbp_1 _2404_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net444),
    .D(_0200_),
    .Q_N(_1073_),
    .Q(\cic_b.delay[1][5] ));
 sg13g2_dfrbp_1 _2405_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net445),
    .D(net327),
    .Q_N(_1072_),
    .Q(\cic_b.delay[1][6] ));
 sg13g2_dfrbp_1 _2406_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net445),
    .D(net240),
    .Q_N(_1071_),
    .Q(\cic_b.delay[1][7] ));
 sg13g2_dfrbp_1 _2407_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net421),
    .D(net311),
    .Q_N(_1070_),
    .Q(\cic_b.delay[1][8] ));
 sg13g2_dfrbp_1 _2408_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net421),
    .D(_0204_),
    .Q_N(_1069_),
    .Q(\cic_b.delay[1][9] ));
 sg13g2_dfrbp_1 _2409_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net422),
    .D(net180),
    .Q_N(_1068_),
    .Q(\cic_b.delay[1][10] ));
 sg13g2_dfrbp_1 _2410_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net422),
    .D(net212),
    .Q_N(_1067_),
    .Q(\cic_b.delay[1][11] ));
 sg13g2_dfrbp_1 _2411_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net417),
    .D(net172),
    .Q_N(_1243_),
    .Q(\cic_b.delay[1][12] ));
 sg13g2_dfrbp_1 _2412_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net448),
    .D(net34),
    .Q_N(_1244_),
    .Q(\cic_b.integrator[0][0] ));
 sg13g2_dfrbp_1 _2413_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net448),
    .D(net574),
    .Q_N(_1245_),
    .Q(\cic_b.integrator[0][1] ));
 sg13g2_dfrbp_1 _2414_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net447),
    .D(net484),
    .Q_N(_1246_),
    .Q(\cic_b.integrator[0][2] ));
 sg13g2_dfrbp_1 _2415_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net442),
    .D(_0054_),
    .Q_N(_1247_),
    .Q(\cic_b.integrator[0][3] ));
 sg13g2_dfrbp_1 _2416_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net440),
    .D(_0055_),
    .Q_N(_1248_),
    .Q(\cic_b.integrator[0][4] ));
 sg13g2_dfrbp_1 _2417_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net440),
    .D(net521),
    .Q_N(_1249_),
    .Q(\cic_b.integrator[0][5] ));
 sg13g2_dfrbp_1 _2418_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net419),
    .D(net550),
    .Q_N(_1250_),
    .Q(\cic_b.integrator[0][6] ));
 sg13g2_dfrbp_1 _2419_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net419),
    .D(net537),
    .Q_N(_1251_),
    .Q(\cic_b.integrator[0][7] ));
 sg13g2_dfrbp_1 _2420_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net420),
    .D(net576),
    .Q_N(_1252_),
    .Q(\cic_b.integrator[0][8] ));
 sg13g2_dfrbp_1 _2421_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net420),
    .D(net509),
    .Q_N(_1253_),
    .Q(\cic_b.integrator[0][9] ));
 sg13g2_dfrbp_1 _2422_ (.CLK(clknet_3_0__leaf_clk),
    .RESET_B(net413),
    .D(_0049_),
    .Q_N(_1254_),
    .Q(\cic_b.integrator[0][10] ));
 sg13g2_dfrbp_1 _2423_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net413),
    .D(_0050_),
    .Q_N(_1255_),
    .Q(\cic_b.integrator[0][11] ));
 sg13g2_dfrbp_1 _2424_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net413),
    .D(net22),
    .Q_N(_1066_),
    .Q(\cic_b.integrator[0][12] ));
 sg13g2_dfrbp_1 _2425_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net453),
    .D(net138),
    .Q_N(_1065_),
    .Q(\cic_b.temp_comb[1][0] ));
 sg13g2_dfrbp_1 _2426_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net453),
    .D(net143),
    .Q_N(_1064_),
    .Q(\cic_b.temp_comb[1][1] ));
 sg13g2_dfrbp_1 _2427_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net453),
    .D(_0210_),
    .Q_N(_1063_),
    .Q(\cic_b.temp_comb[1][2] ));
 sg13g2_dfrbp_1 _2428_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net451),
    .D(_0211_),
    .Q_N(_1062_),
    .Q(\cic_b.temp_comb[1][3] ));
 sg13g2_dfrbp_1 _2429_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net444),
    .D(_0212_),
    .Q_N(_1061_),
    .Q(\cic_b.temp_comb[1][4] ));
 sg13g2_dfrbp_1 _2430_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net444),
    .D(_0213_),
    .Q_N(_1060_),
    .Q(\cic_b.temp_comb[1][5] ));
 sg13g2_dfrbp_1 _2431_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net445),
    .D(_0214_),
    .Q_N(_1059_),
    .Q(\cic_b.temp_comb[1][6] ));
 sg13g2_dfrbp_1 _2432_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net445),
    .D(_0215_),
    .Q_N(_1058_),
    .Q(\cic_b.temp_comb[1][7] ));
 sg13g2_dfrbp_1 _2433_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net423),
    .D(net125),
    .Q_N(_1057_),
    .Q(\cic_b.temp_comb[1][8] ));
 sg13g2_dfrbp_1 _2434_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net423),
    .D(net45),
    .Q_N(_1056_),
    .Q(\cic_b.temp_comb[1][9] ));
 sg13g2_dfrbp_1 _2435_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net423),
    .D(_0218_),
    .Q_N(_1055_),
    .Q(\cic_b.temp_comb[1][10] ));
 sg13g2_dfrbp_1 _2436_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net422),
    .D(_0219_),
    .Q_N(_1054_),
    .Q(\cic_b.temp_comb[1][11] ));
 sg13g2_dfrbp_1 _2437_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net422),
    .D(_0220_),
    .Q_N(_1256_),
    .Q(\cic_b.temp_comb[1][12] ));
 sg13g2_dfrbp_1 _2438_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net416),
    .D(_0008_),
    .Q_N(_1257_),
    .Q(\cic_b.decim_cnt[0] ));
 sg13g2_dfrbp_1 _2439_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net416),
    .D(_0009_),
    .Q_N(_1258_),
    .Q(\cic_b.decim_cnt[1] ));
 sg13g2_dfrbp_1 _2440_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net415),
    .D(_0010_),
    .Q_N(_1259_),
    .Q(\cic_b.decim_cnt[2] ));
 sg13g2_dfrbp_1 _2441_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net415),
    .D(net54),
    .Q_N(_1260_),
    .Q(\cic_b.decim_cnt[3] ));
 sg13g2_dfrbp_1 _2442_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net416),
    .D(net30),
    .Q_N(_1261_),
    .Q(\cic_b.decim_cnt[4] ));
 sg13g2_dfrbp_1 _2443_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net417),
    .D(net548),
    .Q_N(_1262_),
    .Q(\cic_b.decim_cnt[5] ));
 sg13g2_dfrbp_1 _2444_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net416),
    .D(_0014_),
    .Q_N(_1263_),
    .Q(\cic_b.decim_cnt[6] ));
 sg13g2_dfrbp_1 _2445_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net416),
    .D(net58),
    .Q_N(_1053_),
    .Q(\cic_b.decim_cnt[7] ));
 sg13g2_dfrbp_1 _2446_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net460),
    .D(_0221_),
    .Q_N(_1052_),
    .Q(\cic_a.temp_delay[1][0] ));
 sg13g2_dfrbp_1 _2447_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net460),
    .D(net258),
    .Q_N(_1051_),
    .Q(\cic_a.temp_delay[1][1] ));
 sg13g2_dfrbp_1 _2448_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net460),
    .D(net260),
    .Q_N(_1050_),
    .Q(\cic_a.temp_delay[1][2] ));
 sg13g2_dfrbp_1 _2449_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net459),
    .D(net235),
    .Q_N(_1049_),
    .Q(\cic_a.temp_delay[1][3] ));
 sg13g2_dfrbp_1 _2450_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net436),
    .D(net264),
    .Q_N(_1048_),
    .Q(\cic_a.temp_delay[1][4] ));
 sg13g2_dfrbp_1 _2451_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net436),
    .D(net268),
    .Q_N(_1047_),
    .Q(\cic_a.temp_delay[1][5] ));
 sg13g2_dfrbp_1 _2452_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net435),
    .D(net304),
    .Q_N(_1046_),
    .Q(\cic_a.temp_delay[1][6] ));
 sg13g2_dfrbp_1 _2453_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net435),
    .D(net480),
    .Q_N(_1045_),
    .Q(\cic_a.temp_delay[1][7] ));
 sg13g2_dfrbp_1 _2454_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net434),
    .D(net343),
    .Q_N(_1044_),
    .Q(\cic_a.temp_delay[1][8] ));
 sg13g2_dfrbp_1 _2455_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net434),
    .D(net86),
    .Q_N(_1043_),
    .Q(\cic_a.temp_delay[1][9] ));
 sg13g2_dfrbp_1 _2456_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net427),
    .D(net270),
    .Q_N(_1042_),
    .Q(\cic_a.temp_delay[1][10] ));
 sg13g2_dfrbp_1 _2457_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net434),
    .D(_0232_),
    .Q_N(_1041_),
    .Q(\cic_a.temp_delay[1][11] ));
 sg13g2_dfrbp_1 _2458_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net432),
    .D(_0233_),
    .Q_N(_1040_),
    .Q(\cic_a.temp_delay[1][12] ));
 sg13g2_dfrbp_1 _2459_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net448),
    .D(net298),
    .Q_N(_1039_),
    .Q(\cic_b.temp_delay[0][0] ));
 sg13g2_dfrbp_1 _2460_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net448),
    .D(net339),
    .Q_N(_1038_),
    .Q(\cic_b.temp_delay[0][1] ));
 sg13g2_dfrbp_1 _2461_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net447),
    .D(net334),
    .Q_N(_1037_),
    .Q(\cic_b.temp_delay[0][2] ));
 sg13g2_dfrbp_1 _2462_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net441),
    .D(net323),
    .Q_N(_1036_),
    .Q(\cic_b.temp_delay[0][3] ));
 sg13g2_dfrbp_1 _2463_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net440),
    .D(_0238_),
    .Q_N(_1035_),
    .Q(\cic_b.temp_delay[0][4] ));
 sg13g2_dfrbp_1 _2464_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net440),
    .D(_0239_),
    .Q_N(_1034_),
    .Q(\cic_b.temp_delay[0][5] ));
 sg13g2_dfrbp_1 _2465_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net419),
    .D(_0240_),
    .Q_N(_1033_),
    .Q(\cic_b.temp_delay[0][6] ));
 sg13g2_dfrbp_1 _2466_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net419),
    .D(_0241_),
    .Q_N(_1032_),
    .Q(\cic_b.temp_delay[0][7] ));
 sg13g2_dfrbp_1 _2467_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net420),
    .D(_0242_),
    .Q_N(_1031_),
    .Q(\cic_b.temp_delay[0][8] ));
 sg13g2_dfrbp_1 _2468_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net420),
    .D(_0243_),
    .Q_N(_1030_),
    .Q(\cic_b.temp_delay[0][9] ));
 sg13g2_dfrbp_1 _2469_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net414),
    .D(_0244_),
    .Q_N(_1029_),
    .Q(\cic_b.temp_delay[0][10] ));
 sg13g2_dfrbp_1 _2470_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net414),
    .D(net294),
    .Q_N(_1028_),
    .Q(\cic_b.temp_delay[0][11] ));
 sg13g2_dfrbp_1 _2471_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net414),
    .D(net233),
    .Q_N(_1027_),
    .Q(\cic_b.temp_delay[0][12] ));
 sg13g2_dfrbp_1 _2472_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net462),
    .D(_0247_),
    .Q_N(_1026_),
    .Q(\serializer_a.shift_reg[0] ));
 sg13g2_dfrbp_1 _2473_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net462),
    .D(net107),
    .Q_N(_1025_),
    .Q(\serializer_a.shift_reg[1] ));
 sg13g2_dfrbp_1 _2474_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net465),
    .D(_0249_),
    .Q_N(_1024_),
    .Q(\serializer_a.shift_reg[2] ));
 sg13g2_dfrbp_1 _2475_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net462),
    .D(net73),
    .Q_N(_1023_),
    .Q(\serializer_a.shift_reg[3] ));
 sg13g2_dfrbp_1 _2476_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net455),
    .D(_0251_),
    .Q_N(_1022_),
    .Q(\serializer_a.shift_reg[4] ));
 sg13g2_dfrbp_1 _2477_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net460),
    .D(net26),
    .Q_N(_1021_),
    .Q(\serializer_a.shift_reg[5] ));
 sg13g2_dfrbp_1 _2478_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net456),
    .D(net165),
    .Q_N(_1020_),
    .Q(\serializer_a.shift_reg[6] ));
 sg13g2_dfrbp_1 _2479_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net456),
    .D(net118),
    .Q_N(_1019_),
    .Q(\serializer_a.shift_reg[7] ));
 sg13g2_dfrbp_1 _2480_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net455),
    .D(_0255_),
    .Q_N(_1018_),
    .Q(\serializer_a.shift_reg[8] ));
 sg13g2_dfrbp_1 _2481_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net455),
    .D(net65),
    .Q_N(_1017_),
    .Q(\serializer_a.shift_reg[9] ));
 sg13g2_dfrbp_1 _2482_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net456),
    .D(net190),
    .Q_N(_1016_),
    .Q(\serializer_a.shift_reg[10] ));
 sg13g2_dfrbp_1 _2483_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net464),
    .D(net132),
    .Q_N(_1015_),
    .Q(\serializer_a.shift_reg[11] ));
 sg13g2_dfrbp_1 _2484_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net464),
    .D(net84),
    .Q_N(_1264_),
    .Q(\serializer_a.serial_out ));
 sg13g2_dfrbp_1 _2485_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net466),
    .D(_0016_),
    .Q_N(_1014_),
    .Q(\serializer_a.sending ));
 sg13g2_dfrbp_1 _2486_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net449),
    .D(net309),
    .Q_N(_1013_),
    .Q(\cic_b.temp_delay[1][0] ));
 sg13g2_dfrbp_1 _2487_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net449),
    .D(_0261_),
    .Q_N(_1012_),
    .Q(\cic_b.temp_delay[1][1] ));
 sg13g2_dfrbp_1 _2488_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net447),
    .D(_0262_),
    .Q_N(_1011_),
    .Q(\cic_b.temp_delay[1][2] ));
 sg13g2_dfrbp_1 _2489_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net447),
    .D(_0263_),
    .Q_N(_1010_),
    .Q(\cic_b.temp_delay[1][3] ));
 sg13g2_dfrbp_1 _2490_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net442),
    .D(net487),
    .Q_N(_1009_),
    .Q(\cic_b.temp_delay[1][4] ));
 sg13g2_dfrbp_1 _2491_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net444),
    .D(net154),
    .Q_N(_1008_),
    .Q(\cic_b.temp_delay[1][5] ));
 sg13g2_dfrbp_1 _2492_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net445),
    .D(net349),
    .Q_N(_1007_),
    .Q(\cic_b.temp_delay[1][6] ));
 sg13g2_dfrbp_1 _2493_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net419),
    .D(net494),
    .Q_N(_1006_),
    .Q(\cic_b.temp_delay[1][7] ));
 sg13g2_dfrbp_1 _2494_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net421),
    .D(_0268_),
    .Q_N(_1005_),
    .Q(\cic_b.temp_delay[1][8] ));
 sg13g2_dfrbp_1 _2495_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net421),
    .D(net98),
    .Q_N(_1004_),
    .Q(\cic_b.temp_delay[1][9] ));
 sg13g2_dfrbp_1 _2496_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net422),
    .D(_0270_),
    .Q_N(_1003_),
    .Q(\cic_b.temp_delay[1][10] ));
 sg13g2_dfrbp_1 _2497_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net422),
    .D(_0271_),
    .Q_N(_1002_),
    .Q(\cic_b.temp_delay[1][11] ));
 sg13g2_dfrbp_1 _2498_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net417),
    .D(_0272_),
    .Q_N(_1265_),
    .Q(\cic_b.temp_delay[1][12] ));
 sg13g2_dfrbp_1 _2499_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net463),
    .D(net404),
    .Q_N(_1001_),
    .Q(\serializer_a.valid ));
 sg13g2_dfrbp_1 _2500_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net452),
    .D(_0273_),
    .Q_N(_1000_),
    .Q(\serializer_b.shift_reg[0] ));
 sg13g2_dfrbp_1 _2501_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net452),
    .D(_0274_),
    .Q_N(_0999_),
    .Q(\serializer_b.shift_reg[1] ));
 sg13g2_dfrbp_1 _2502_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net451),
    .D(_0275_),
    .Q_N(_0998_),
    .Q(\serializer_b.shift_reg[2] ));
 sg13g2_dfrbp_1 _2503_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net451),
    .D(net28),
    .Q_N(_0997_),
    .Q(\serializer_b.shift_reg[3] ));
 sg13g2_dfrbp_1 _2504_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net443),
    .D(net77),
    .Q_N(_0996_),
    .Q(\serializer_b.shift_reg[4] ));
 sg13g2_dfrbp_1 _2505_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net443),
    .D(net43),
    .Q_N(_0995_),
    .Q(\serializer_b.shift_reg[5] ));
 sg13g2_dfrbp_1 _2506_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net443),
    .D(net150),
    .Q_N(_0994_),
    .Q(\serializer_b.shift_reg[6] ));
 sg13g2_dfrbp_1 _2507_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net443),
    .D(net222),
    .Q_N(_0993_),
    .Q(\serializer_b.shift_reg[7] ));
 sg13g2_dfrbp_1 _2508_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net443),
    .D(net123),
    .Q_N(_0992_),
    .Q(\serializer_b.shift_reg[8] ));
 sg13g2_dfrbp_1 _2509_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net443),
    .D(net507),
    .Q_N(_0991_),
    .Q(\serializer_b.shift_reg[9] ));
 sg13g2_dfrbp_1 _2510_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net444),
    .D(net247),
    .Q_N(_0990_),
    .Q(\serializer_b.shift_reg[10] ));
 sg13g2_dfrbp_1 _2511_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net454),
    .D(net135),
    .Q_N(_0989_),
    .Q(\serializer_b.shift_reg[11] ));
 sg13g2_dfrbp_1 _2512_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net452),
    .D(net121),
    .Q_N(_1266_),
    .Q(\serializer_b.serial_out ));
 sg13g2_dfrbp_1 _2513_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net451),
    .D(_0020_),
    .Q_N(_0988_),
    .Q(\serializer_b.sending ));
 sg13g2_dfrbp_1 _2514_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net463),
    .D(_0286_),
    .Q_N(_0987_),
    .Q(\serializer_ab_subtr.bit_cnt[0] ));
 sg13g2_dfrbp_1 _2515_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net463),
    .D(_0287_),
    .Q_N(_0986_),
    .Q(\serializer_ab_subtr.bit_cnt[1] ));
 sg13g2_dfrbp_1 _2516_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net464),
    .D(_0288_),
    .Q_N(_0985_),
    .Q(\serializer_ab_subtr.bit_cnt[2] ));
 sg13g2_dfrbp_1 _2517_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net463),
    .D(net47),
    .Q_N(_1267_),
    .Q(\serializer_ab_subtr.bit_cnt[3] ));
 sg13g2_dfrbp_1 _2518_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net453),
    .D(net401),
    .Q_N(_0984_),
    .Q(\serializer_b.valid ));
 sg13g2_dfrbp_1 _2519_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net451),
    .D(_0290_),
    .Q_N(_0983_),
    .Q(\serializer_b.bit_cnt[0] ));
 sg13g2_dfrbp_1 _2520_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net451),
    .D(net70),
    .Q_N(_0982_),
    .Q(\serializer_b.bit_cnt[1] ));
 sg13g2_dfrbp_1 _2521_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net451),
    .D(_0292_),
    .Q_N(_0981_),
    .Q(\serializer_b.bit_cnt[2] ));
 sg13g2_dfrbp_1 _2522_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net451),
    .D(net40),
    .Q_N(_0980_),
    .Q(\serializer_b.bit_cnt[3] ));
 sg13g2_dfrbp_1 _2523_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net463),
    .D(net220),
    .Q_N(_0979_),
    .Q(\serializer_ab_subtr.shift_reg[0] ));
 sg13g2_dfrbp_1 _2524_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net463),
    .D(_0295_),
    .Q_N(_0978_),
    .Q(\serializer_ab_subtr.shift_reg[1] ));
 sg13g2_dfrbp_1 _2525_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net462),
    .D(_0296_),
    .Q_N(_0977_),
    .Q(\serializer_ab_subtr.shift_reg[2] ));
 sg13g2_dfrbp_1 _2526_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net462),
    .D(net281),
    .Q_N(_0976_),
    .Q(\serializer_ab_subtr.shift_reg[3] ));
 sg13g2_dfrbp_1 _2527_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net462),
    .D(_0298_),
    .Q_N(_0975_),
    .Q(\serializer_ab_subtr.shift_reg[4] ));
 sg13g2_dfrbp_1 _2528_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net455),
    .D(net188),
    .Q_N(_0974_),
    .Q(\serializer_ab_subtr.shift_reg[5] ));
 sg13g2_dfrbp_1 _2529_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net455),
    .D(_0300_),
    .Q_N(_0973_),
    .Q(\serializer_ab_subtr.shift_reg[6] ));
 sg13g2_dfrbp_1 _2530_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net455),
    .D(net184),
    .Q_N(_0972_),
    .Q(\serializer_ab_subtr.shift_reg[7] ));
 sg13g2_dfrbp_1 _2531_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net455),
    .D(_0302_),
    .Q_N(_0971_),
    .Q(\serializer_ab_subtr.shift_reg[8] ));
 sg13g2_dfrbp_1 _2532_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net455),
    .D(_0303_),
    .Q_N(_0970_),
    .Q(\serializer_ab_subtr.shift_reg[9] ));
 sg13g2_dfrbp_1 _2533_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net462),
    .D(_0304_),
    .Q_N(_0969_),
    .Q(\serializer_ab_subtr.shift_reg[10] ));
 sg13g2_dfrbp_1 _2534_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net462),
    .D(_0305_),
    .Q_N(_0968_),
    .Q(\serializer_ab_subtr.shift_reg[11] ));
 sg13g2_dfrbp_1 _2535_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net463),
    .D(_0306_),
    .Q_N(_1268_),
    .Q(\serializer_ab_subtr.serial_out ));
 sg13g2_dfrbp_1 _2536_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net463),
    .D(_0018_),
    .Q_N(_0967_),
    .Q(\serializer_ab_subtr.sending ));
 sg13g2_dfrbp_1 _2537_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net466),
    .D(_0307_),
    .Q_N(_0966_),
    .Q(\serializer_a.bit_cnt[0] ));
 sg13g2_dfrbp_1 _2538_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net466),
    .D(_0308_),
    .Q_N(_0965_),
    .Q(\serializer_a.bit_cnt[1] ));
 sg13g2_dfrbp_1 _2539_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net466),
    .D(_0309_),
    .Q_N(_0964_),
    .Q(\serializer_a.bit_cnt[2] ));
 sg13g2_dfrbp_1 _2540_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net466),
    .D(net56),
    .Q_N(_1269_),
    .Q(\serializer_a.bit_cnt[3] ));
 sg13g2_dfrbp_1 _2541_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net452),
    .D(_0019_),
    .Q_N(_0963_),
    .Q(\serializer_ab_subtr.valid ));
 sg13g2_tielo tt_um_ds_comp_adc_5 (.L_LO(net5));
 sg13g2_tielo tt_um_ds_comp_adc_6 (.L_LO(net6));
 sg13g2_tielo tt_um_ds_comp_adc_7 (.L_LO(net7));
 sg13g2_tielo tt_um_ds_comp_adc_8 (.L_LO(net8));
 sg13g2_tielo tt_um_ds_comp_adc_9 (.L_LO(net9));
 sg13g2_tielo tt_um_ds_comp_adc_10 (.L_LO(net10));
 sg13g2_tielo tt_um_ds_comp_adc_11 (.L_LO(net11));
 sg13g2_tielo tt_um_ds_comp_adc_12 (.L_LO(net12));
 sg13g2_tielo tt_um_ds_comp_adc_13 (.L_LO(net13));
 sg13g2_tielo tt_um_ds_comp_adc_14 (.L_LO(net14));
 sg13g2_tielo tt_um_ds_comp_adc_15 (.L_LO(net15));
 sg13g2_tielo tt_um_ds_comp_adc_16 (.L_LO(net16));
 sg13g2_tielo tt_um_ds_comp_adc_17 (.L_LO(net17));
 sg13g2_tielo tt_um_ds_comp_adc_18 (.L_LO(net18));
 sg13g2_tielo tt_um_ds_comp_adc_19 (.L_LO(net19));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_2 _2558_ (.A(pdm_a),
    .X(uo_out[0]));
 sg13g2_buf_2 _2559_ (.A(pdm_b),
    .X(uo_out[1]));
 sg13g2_buf_1 _2560_ (.A(\serializer_a.serial_out ),
    .X(uo_out[2]));
 sg13g2_buf_1 _2561_ (.A(\serializer_b.serial_out ),
    .X(uo_out[3]));
 sg13g2_buf_1 _2562_ (.A(\serializer_ab_subtr.serial_out ),
    .X(uo_out[4]));
 sg13g2_buf_1 _2563_ (.A(\serializer_a.valid ),
    .X(uo_out[5]));
 sg13g2_buf_1 _2564_ (.A(\serializer_b.valid ),
    .X(uo_out[6]));
 sg13g2_buf_1 _2565_ (.A(\serializer_ab_subtr.valid ),
    .X(uo_out[7]));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(net354));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(net354));
 sg13g2_buf_2 fanout354 (.A(net359),
    .X(net354));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(net359));
 sg13g2_buf_2 fanout356 (.A(net359),
    .X(net356));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(net358));
 sg13g2_buf_2 fanout358 (.A(net359),
    .X(net358));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(_0392_));
 sg13g2_buf_2 fanout360 (.A(net362),
    .X(net360));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(net374));
 sg13g2_buf_2 fanout362 (.A(net374),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(net366),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(net366),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(net366),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(net374),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(net369),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(net369),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(net374),
    .X(net369));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(net373));
 sg13g2_buf_2 fanout371 (.A(net372),
    .X(net371));
 sg13g2_buf_1 fanout372 (.A(net373),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(net374),
    .X(net373));
 sg13g2_buf_4 fanout374 (.X(net374),
    .A(_0391_));
 sg13g2_buf_4 fanout375 (.X(net375),
    .A(net379));
 sg13g2_buf_2 fanout376 (.A(net379),
    .X(net376));
 sg13g2_buf_4 fanout377 (.X(net377),
    .A(net379));
 sg13g2_buf_2 fanout378 (.A(net379),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_0886_),
    .X(net379));
 sg13g2_buf_4 fanout380 (.X(net380),
    .A(net382));
 sg13g2_buf_4 fanout381 (.X(net381),
    .A(net382));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(_0886_));
 sg13g2_buf_2 fanout383 (.A(net385),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(net385),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(net386),
    .X(net385));
 sg13g2_buf_4 fanout386 (.X(net386),
    .A(net389));
 sg13g2_buf_2 fanout387 (.A(net388),
    .X(net387));
 sg13g2_buf_4 fanout388 (.X(net388),
    .A(net389));
 sg13g2_buf_2 fanout389 (.A(_0885_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(net391),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(net392),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(net395),
    .X(net392));
 sg13g2_buf_4 fanout393 (.X(net393),
    .A(net394));
 sg13g2_buf_2 fanout394 (.A(net395),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_0885_),
    .X(net395));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(_0866_));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(_0862_));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(_0869_));
 sg13g2_buf_2 fanout399 (.A(_0869_),
    .X(net399));
 sg13g2_buf_4 fanout400 (.X(net400),
    .A(net401));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(_0021_));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(_0730_));
 sg13g2_buf_2 fanout403 (.A(net404),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_0017_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(net406),
    .X(net405));
 sg13g2_buf_1 fanout406 (.A(\serializer_ab_subtr.sending ),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(\serializer_ab_subtr.sending ),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(net409),
    .X(net408));
 sg13g2_buf_4 fanout409 (.X(net409),
    .A(\serializer_b.sending ));
 sg13g2_buf_2 fanout410 (.A(net412),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(net412),
    .X(net411));
 sg13g2_buf_1 fanout412 (.A(net569),
    .X(net412));
 sg13g2_buf_4 fanout413 (.X(net413),
    .A(net415));
 sg13g2_buf_2 fanout414 (.A(net415),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(net418),
    .X(net415));
 sg13g2_buf_4 fanout416 (.X(net416),
    .A(net417));
 sg13g2_buf_4 fanout417 (.X(net417),
    .A(net418));
 sg13g2_buf_2 fanout418 (.A(net439),
    .X(net418));
 sg13g2_buf_4 fanout419 (.X(net419),
    .A(net424));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(net424));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(net423));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(net424));
 sg13g2_buf_2 fanout423 (.A(net424),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(net439),
    .X(net424));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(net426));
 sg13g2_buf_4 fanout426 (.X(net426),
    .A(net427));
 sg13g2_buf_4 fanout427 (.X(net427),
    .A(net432));
 sg13g2_buf_4 fanout428 (.X(net428),
    .A(net431));
 sg13g2_buf_2 fanout429 (.A(net431),
    .X(net429));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(net431));
 sg13g2_buf_2 fanout431 (.A(net432),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(net439),
    .X(net432));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(net438));
 sg13g2_buf_4 fanout434 (.X(net434),
    .A(net438));
 sg13g2_buf_4 fanout435 (.X(net435),
    .A(net437));
 sg13g2_buf_4 fanout436 (.X(net436),
    .A(net437));
 sg13g2_buf_4 fanout437 (.X(net437),
    .A(net438));
 sg13g2_buf_2 fanout438 (.A(net439),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(rst_n),
    .X(net439));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(net441));
 sg13g2_buf_4 fanout441 (.X(net441),
    .A(net446));
 sg13g2_buf_2 fanout442 (.A(net446),
    .X(net442));
 sg13g2_buf_4 fanout443 (.X(net443),
    .A(net444));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(net446));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(net446));
 sg13g2_buf_2 fanout446 (.A(net467),
    .X(net446));
 sg13g2_buf_4 fanout447 (.X(net447),
    .A(net450));
 sg13g2_buf_4 fanout448 (.X(net448),
    .A(net450));
 sg13g2_buf_4 fanout449 (.X(net449),
    .A(net450));
 sg13g2_buf_2 fanout450 (.A(net467),
    .X(net450));
 sg13g2_buf_4 fanout451 (.X(net451),
    .A(net454));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(net453));
 sg13g2_buf_2 fanout453 (.A(net454),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(net467),
    .X(net454));
 sg13g2_buf_4 fanout455 (.X(net455),
    .A(net457));
 sg13g2_buf_2 fanout456 (.A(net457),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(net461),
    .X(net457));
 sg13g2_buf_4 fanout458 (.X(net458),
    .A(net459));
 sg13g2_buf_4 fanout459 (.X(net459),
    .A(net461));
 sg13g2_buf_4 fanout460 (.X(net460),
    .A(net461));
 sg13g2_buf_2 fanout461 (.A(net467),
    .X(net461));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(net464));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(net464));
 sg13g2_buf_2 fanout464 (.A(net467),
    .X(net464));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(net466));
 sg13g2_buf_4 fanout466 (.X(net466),
    .A(net467));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_4 input3 (.X(net3),
    .A(ui_in[7]));
 sg13g2_tielo tt_um_ds_comp_adc_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_37_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_18_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\cic_b.integrator[0][10] ),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0883_),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0051_),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold4 (.A(\cic_b.decim_cnt[0] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cic_a.decim_cnt[0] ),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold6 (.A(\serializer_a.shift_reg[4] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0252_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold8 (.A(\serializer_b.shift_reg[2] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0276_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cic_b.decim_cnt[4] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0012_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cic_a.pdm_in ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0022_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold14 (.A(\cic_b.pdm_in ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0048_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold16 (.A(\cic_a.decim_cnt[4] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0004_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold18 (.A(\serializer_a.shift_reg[0] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0552_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold20 (.A(\serializer_b.bit_cnt[3] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0293_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold22 (.A(\serializer_b.shift_reg[4] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0579_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0278_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold25 (.A(\cic_b.temp_comb[1][9] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0217_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold27 (.A(\serializer_ab_subtr.bit_cnt[3] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0289_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold29 (.A(\cic_b.temp_comb[1][7] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold30 (.A(\cic_a.decim_cnt[3] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0003_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold32 (.A(\serializer_ab_subtr.bit_cnt[2] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0593_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cic_b.decim_cnt[3] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0011_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold36 (.A(\serializer_a.bit_cnt[3] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0310_),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold38 (.A(\cic_b.decim_cnt[7] ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0015_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cic_a.temp_comb[1][9] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold41 (.A(\cic_a.temp_comb[1][11] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold42 (.A(\cic_a.temp_comb[1][5] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold43 (.A(\serializer_b.shift_reg[0] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0571_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold45 (.A(\serializer_a.shift_reg[8] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0256_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold47 (.A(\cic_a.temp_delay[0][5] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0083_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold49 (.A(\serializer_b.bit_cnt[1] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0596_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0291_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold52 (.A(\serializer_a.shift_reg[2] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0555_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0250_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold55 (.A(\serializer_b.bit_cnt[2] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0600_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold57 (.A(\serializer_b.shift_reg[3] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0277_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold59 (.A(\cic_b.temp_comb[1][3] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0185_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold61 (.A(\serializer_b.bit_cnt[0] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold62 (.A(\serializer_b.shift_reg[1] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0573_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold64 (.A(\serializer_a.serial_out ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0259_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold66 (.A(\cic_a.temp_delay[1][9] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0230_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold68 (.A(\cic_b.temp_delay[0][9] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0165_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold70 (.A(\cic_b.temp_comb[1][5] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cic_b.integrator[1][9] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold72 (.A(\cic_b.decim_cnt[1] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cic_a.temp_delay[0][9] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0152_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cic_b.temp_comb[1][4] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0186_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold77 (.A(\serializer_a.bit_cnt[0] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold78 (.A(\cic_b.temp_delay[1][9] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0269_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cic_a.temp_comb[1][0] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0130_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold82 (.A(\cic_b.temp_delay[0][8] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0164_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold84 (.A(\cic_a.temp_comb[1][12] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0142_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold86 (.A(\serializer_a.bit_cnt[1] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold87 (.A(\serializer_a.shift_reg[1] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0248_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cic_a.decim_cnt[1] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cic_a.temp_comb[1][2] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold91 (.A(\serializer_ab_subtr.bit_cnt[0] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cic_b.delay[1][3] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0492_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold94 (.A(\cic_b.integrator[0][11] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cic_b.temp_comb[1][2] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold96 (.A(\serializer_a.shift_reg[3] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0557_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold98 (.A(\serializer_a.shift_reg[7] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0254_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cic_b.filtered_out[5] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold101 (.A(\serializer_b.serial_out ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0285_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold103 (.A(\serializer_b.shift_reg[8] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0281_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cic_b.temp_comb[1][8] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0216_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold107 (.A(\cic_a.temp_comb[1][4] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0108_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cic_a.temp_comb[1][6] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cic_a.filtered_out[2] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold111 (.A(\cic_b.delay[1][4] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold112 (.A(\serializer_a.shift_reg[11] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0258_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cic_b.temp_comb[1][10] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold115 (.A(\serializer_b.shift_reg[11] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0284_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold117 (.A(\cic_b.temp_comb[1][6] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cic_b.temp_comb[1][0] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0208_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cic_a.integrator[0][12] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0025_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cic_a.filtered_out[8] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold123 (.A(\cic_b.temp_comb[1][1] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0209_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cic_b.filtered_out[2] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0574_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold127 (.A(\cic_b.temp_delay[0][5] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0161_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold129 (.A(\cic_a.temp_comb[1][7] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold130 (.A(\serializer_b.shift_reg[6] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0279_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold132 (.A(\serializer_ab_subtr.serial_out ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0681_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cic_b.temp_delay[1][5] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0265_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold136 (.A(\serializer_ab_subtr.shift_reg[2] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0614_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold138 (.A(\cic_a.delay[1][7] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0124_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold140 (.A(\serializer_ab_subtr.shift_reg[8] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0655_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold142 (.A(\serializer_a.bit_cnt[2] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cic_a.temp_comb[1][3] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0133_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold145 (.A(\serializer_a.shift_reg[5] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0253_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold147 (.A(\serializer_ab_subtr.bit_cnt[1] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold148 (.A(\serializer_ab_subtr.shift_reg[6] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0638_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold150 (.A(\cic_a.delay[0][12] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0090_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cic_b.delay[1][12] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0207_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cic_a.temp_delay[0][7] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0085_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold156 (.A(\cic_a.delay[0][8] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0086_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold158 (.A(\cic_a.decim_cnt[7] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0007_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold160 (.A(\cic_b.delay[1][10] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0205_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold162 (.A(\cic_b.filtered_out[0] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold163 (.A(\serializer_ab_subtr.shift_reg[7] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0643_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0301_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold166 (.A(\cic_b.temp_comb[1][11] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold167 (.A(\serializer_ab_subtr.shift_reg[5] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0630_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0299_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold170 (.A(\serializer_a.shift_reg[10] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0257_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold172 (.A(\cic_a.temp_comb[1][10] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cic_b.delay[0][12] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0168_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold175 (.A(\cic_a.temp_comb[1][1] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0131_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold177 (.A(\cic_a.temp_delay[0][6] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0084_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold179 (.A(\cic_a.temp_comb[0][12] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0103_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold181 (.A(\cic_a.delay[1][9] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cic_b.temp_comb[0][11] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0180_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold184 (.A(\cic_a.temp_delay[0][1] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0079_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold186 (.A(\cic_b.delay[0][0] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0156_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold188 (.A(\cic_b.temp_comb[0][12] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0181_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold190 (.A(\cic_b.delay[0][11] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0167_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold192 (.A(\cic_b.delay[1][11] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0206_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold194 (.A(\cic_b.delay[1][9] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold195 (.A(\cic_b.temp_comb[0][10] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold196 (.A(\cic_a.delay[1][10] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0127_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold198 (.A(\cic_b.temp_delay[0][4] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0160_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold200 (.A(\serializer_ab_subtr.shift_reg[0] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0294_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold202 (.A(\serializer_b.shift_reg[7] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0280_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold204 (.A(\cic_b.temp_delay[0][6] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0162_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold206 (.A(\cic_b.filtered_out[1] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold207 (.A(\cic_b.delay[0][2] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0158_),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold209 (.A(\cic_a.integrator[0][2] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0027_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold211 (.A(\cic_b.temp_delay[0][7] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0163_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold213 (.A(\cic_b.temp_delay[0][12] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0246_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold215 (.A(\cic_a.temp_delay[1][3] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0224_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold217 (.A(\cic_a.delay[1][12] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0129_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold219 (.A(\cic_b.integrator[1][6] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold220 (.A(\cic_b.delay[1][7] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0202_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold222 (.A(\cic_a.filtered_out[0] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold223 (.A(\cic_a.temp_delay[0][3] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0081_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold225 (.A(\cic_a.temp_delay[0][11] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0154_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold227 (.A(\serializer_b.shift_reg[10] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0283_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold229 (.A(\cic_b.temp_delay[0][10] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0166_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold231 (.A(\cic_b.filtered_out[8] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold232 (.A(\cic_b.delay[1][5] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold233 (.A(\cic_a.filtered_out[11] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold234 (.A(\cic_b.delay[1][0] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0195_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold236 (.A(\cic_a.delay[0][0] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0078_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold238 (.A(\cic_a.temp_delay[1][1] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold239 (.A(_0222_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold240 (.A(\cic_a.temp_delay[1][2] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0223_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold242 (.A(\cic_b.temp_delay[1][1] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0196_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold244 (.A(\cic_a.temp_delay[1][4] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0225_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold246 (.A(\cic_a.delay[1][8] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0125_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold248 (.A(\cic_a.temp_delay[1][5] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0226_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold250 (.A(\cic_a.temp_delay[1][10] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0231_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold252 (.A(\cic_a.temp_delay[0][0] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0143_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold254 (.A(\cic_a.filtered_out[10] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold255 (.A(\cic_a.temp_delay[1][12] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold256 (.A(\cic_b.temp_delay[1][2] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0197_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold258 (.A(\cic_b.temp_comb[0][2] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold259 (.A(\cic_a.delay[1][5] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold260 (.A(\serializer_ab_subtr.shift_reg[3] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0619_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0297_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold263 (.A(\cic_a.integrator[1][1] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold264 (.A(\cic_b.temp_comb[1][12] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold265 (.A(\cic_b.filtered_out[7] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold266 (.A(\cic_a.temp_delay[0][2] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0145_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold268 (.A(\cic_a.delay[0][9] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold269 (.A(\cic_a.delay[1][4] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold270 (.A(\cic_a.filtered_out[3] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold271 (.A(\cic_b.temp_delay[1][10] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold272 (.A(\cic_a.temp_delay[1][0] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0117_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold274 (.A(\cic_b.temp_delay[0][11] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0245_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold276 (.A(\cic_b.delay[0][3] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0159_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold278 (.A(\cic_b.temp_delay[0][0] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0234_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold280 (.A(\cic_a.delay[1][3] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold281 (.A(\cic_a.integrator[1][3] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold282 (.A(\cic_a.filtered_out[12] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold283 (.A(\cic_b.filtered_out[6] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold284 (.A(\cic_a.temp_delay[1][6] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0227_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold286 (.A(\cic_b.filtered_out[12] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold287 (.A(\cic_b.integrator[1][7] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold288 (.A(\serializer_ab_subtr.shift_reg[1] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold289 (.A(\cic_b.temp_delay[1][0] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0260_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold291 (.A(\cic_b.temp_delay[1][8] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0203_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold293 (.A(\cic_b.temp_comb[0][8] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold294 (.A(\cic_a.temp_delay[0][10] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold295 (.A(_0153_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold296 (.A(\cic_b.delay[0][1] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0157_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold298 (.A(\cic_a.filtered_out[9] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold299 (.A(\cic_b.temp_comb[0][1] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold300 (.A(\cic_a.delay[1][11] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0128_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold302 (.A(\cic_b.temp_delay[1][3] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold303 (.A(\cic_b.temp_delay[0][3] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0237_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold305 (.A(\cic_a.delay[1][6] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold306 (.A(\cic_b.filtered_out[10] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold307 (.A(\cic_b.delay[1][6] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0201_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold309 (.A(\cic_a.integrator[1][6] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold310 (.A(\cic_a.temp_delay[0][4] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0147_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold312 (.A(\cic_a.filtered_out[1] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold313 (.A(\cic_a.delay[0][10] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold314 (.A(\cic_b.temp_delay[0][2] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0236_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold316 (.A(\cic_a.delay[0][11] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold317 (.A(\cic_a.integrator[1][7] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold318 (.A(\cic_a.delay[0][2] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold319 (.A(\cic_b.temp_delay[0][1] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0235_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold321 (.A(\cic_a.decim_cnt[6] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0735_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold323 (.A(\cic_a.temp_delay[1][8] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0229_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold325 (.A(\cic_b.temp_comb[0][3] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold326 (.A(\cic_a.filtered_out[5] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold327 (.A(\cic_b.integrator[1][4] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold328 (.A(\cic_b.temp_delay[1][11] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold329 (.A(\cic_b.temp_delay[1][6] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0266_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold331 (.A(\serializer_ab_subtr.shift_reg[10] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0670_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold333 (.A(\cic_a.temp_delay[0][8] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0151_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold335 (.A(\cic_a.delay[0][4] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold336 (.A(\cic_b.integrator[1][8] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold337 (.A(\cic_a.delay[1][1] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold338 (.A(\cic_a.delay[1][2] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold339 (.A(\cic_b.temp_comb[0][9] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0178_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold341 (.A(\cic_a.temp_comb[0][11] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold342 (.A(\cic_a.filtered_out[6] ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold343 (.A(\cic_b.integrator[1][10] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold344 (.A(\cic_a.temp_delay[1][7] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0228_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold346 (.A(\cic_a.temp_delay[0][12] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0155_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold348 (.A(\cic_b.integrator[0][2] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0053_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold350 (.A(\cic_b.delay[0][2] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold351 (.A(\cic_b.temp_delay[1][4] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0264_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold353 (.A(\cic_b.filtered_out[11] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold354 (.A(\serializer_ab_subtr.shift_reg[11] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0676_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold356 (.A(\cic_a.integrator[1][5] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold357 (.A(\cic_b.integrator[1][5] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold358 (.A(\cic_b.temp_delay[1][7] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0267_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold360 (.A(\cic_b.filtered_out[9] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold361 (.A(\cic_b.temp_comb[0][7] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0176_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold363 (.A(\cic_b.delay[0][8] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold364 (.A(\cic_a.temp_delay[1][11] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold365 (.A(\cic_a.integrator[0][5] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0030_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold367 (.A(\cic_a.temp_comb[0][0] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold368 (.A(\serializer_ab_subtr.shift_reg[4] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0625_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold370 (.A(\cic_a.temp_comb[0][4] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold371 (.A(\serializer_b.shift_reg[9] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0282_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold373 (.A(\cic_b.integrator[0][9] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0060_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold375 (.A(\cic_b.temp_delay[1][12] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold376 (.A(\cic_b.temp_comb[0][4] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold377 (.A(\cic_b.integrator[0][9] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold378 (.A(\cic_b.integrator[1][1] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold379 (.A(\cic_a.integrator[1][0] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0035_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold381 (.A(\cic_a.temp_comb[0][10] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold382 (.A(\cic_a.temp_comb[1][8] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold383 (.A(\cic_b.integrator[1][11] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold384 (.A(\cic_a.temp_comb[0][7] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold385 (.A(\cic_b.integrator[0][5] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0056_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold387 (.A(\cic_a.delay[0][0] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold388 (.A(\serializer_ab_subtr.shift_reg[9] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0661_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold390 (.A(\cic_b.integrator[0][0] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0061_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold392 (.A(\cic_a.temp_comb[0][1] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold393 (.A(\cic_b.temp_comb[0][0] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0169_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold395 (.A(\cic_a.temp_comb[0][5] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0096_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold397 (.A(\cic_b.integrator[1][2] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold398 (.A(\cic_a.filtered_out[7] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold399 (.A(\cic_a.integrator[0][7] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0032_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold401 (.A(\cic_b.integrator[0][7] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0058_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold403 (.A(\cic_a.temp_comb[0][3] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold404 (.A(\cic_a.temp_comb[0][8] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold405 (.A(\cic_b.temp_comb[0][5] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0174_),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold407 (.A(\cic_a.integrator[0][9] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0034_),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold409 (.A(\cic_b.temp_comb[0][6] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold410 (.A(\cic_a.integrator[0][10] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold411 (.A(\cic_a.temp_comb[0][6] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold412 (.A(\cic_b.decim_cnt[5] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0013_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold414 (.A(\cic_b.integrator[0][6] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0057_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold416 (.A(\cic_a.temp_comb[0][9] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold417 (.A(\cic_a.integrator[0][6] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0031_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold419 (.A(\cic_a.temp_comb[0][2] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0093_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold421 (.A(\cic_a.decim_cnt[5] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold422 (.A(\cic_b.integrator[0][12] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0848_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold424 (.A(_0064_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold425 (.A(\cic_b.integrator[0][3] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold426 (.A(\cic_a.decim_cnt[2] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold427 (.A(\cic_a.integrator[0][3] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold428 (.A(\cic_b.decim_cnt[2] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold429 (.A(\cic_a.integrator[1][12] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0038_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold431 (.A(\cic_a.integrator[0][0] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0039_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold433 (.A(\cic_b.decim_cnt[6] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold434 (.A(\serializer_a.sending ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold435 (.A(\cic_b.integrator[1][0] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0065_),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold437 (.A(\serializer_b.sending ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold438 (.A(\cic_b.integrator[0][1] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0052_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold440 (.A(\cic_b.integrator[0][8] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0059_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold442 (.A(\cic_a.integrator[0][1] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold443 (.A(\cic_a.integrator[1][9] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0047_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold445 (.A(\cic_a.integrator[0][4] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold446 (.A(\cic_a.integrator[1][2] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold447 (.A(\cic_a.integrator[0][8] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold448 (.A(\cic_b.integrator[0][4] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold449 (.A(\cic_a.integrator[0][11] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold450 (.A(\cic_b.integrator[0][5] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold451 (.A(_0814_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold452 (.A(\cic_b.integrator[0][7] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold453 (.A(\cic_b.integrator[1][3] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0067_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold455 (.A(\cic_a.integrator[0][5] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0043_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold457 (.A(\cic_a.integrator[1][11] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0037_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold459 (.A(\cic_a.integrator[1][10] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0036_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold461 (.A(\cic_b.integrator[0][3] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold462 (.A(_0807_),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0068_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold464 (.A(\cic_a.integrator[1][8] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold465 (.A(\cic_b.integrator[0][6] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0826_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold467 (.A(\cic_a.integrator[0][7] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0045_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold469 (.A(\cic_a.integrator[0][4] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold470 (.A(_0759_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold471 (.A(_0042_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold472 (.A(\cic_a.integrator[0][1] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold473 (.A(\cic_b.integrator[0][2] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold474 (.A(_0803_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0066_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold476 (.A(\cic_a.delay[1][5] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold477 (.A(\cic_b.temp_comb[0][6] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold478 (.A(\cic_a.delay[1][9] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold479 (.A(\cic_b.delay[1][5] ),
    .X(net614));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_239 ();
 sg13g2_decap_8 FILLER_4_272 ();
 sg13g2_decap_8 FILLER_4_279 ();
 sg13g2_decap_8 FILLER_4_286 ();
 sg13g2_decap_8 FILLER_4_293 ();
 sg13g2_decap_8 FILLER_4_300 ();
 sg13g2_decap_8 FILLER_4_307 ();
 sg13g2_decap_8 FILLER_4_314 ();
 sg13g2_decap_8 FILLER_4_321 ();
 sg13g2_decap_8 FILLER_4_328 ();
 sg13g2_decap_8 FILLER_4_335 ();
 sg13g2_decap_8 FILLER_4_342 ();
 sg13g2_decap_8 FILLER_4_349 ();
 sg13g2_decap_8 FILLER_4_356 ();
 sg13g2_decap_8 FILLER_4_363 ();
 sg13g2_decap_8 FILLER_4_370 ();
 sg13g2_decap_8 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_fill_2 FILLER_5_262 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_4 FILLER_6_189 ();
 sg13g2_fill_1 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_211 ();
 sg13g2_decap_4 FILLER_6_218 ();
 sg13g2_fill_1 FILLER_6_222 ();
 sg13g2_fill_1 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_fill_2 FILLER_6_249 ();
 sg13g2_fill_1 FILLER_6_274 ();
 sg13g2_decap_8 FILLER_6_279 ();
 sg13g2_decap_8 FILLER_6_286 ();
 sg13g2_decap_8 FILLER_6_293 ();
 sg13g2_decap_8 FILLER_6_300 ();
 sg13g2_decap_8 FILLER_6_307 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_8 FILLER_6_370 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_fill_2 FILLER_7_182 ();
 sg13g2_fill_1 FILLER_7_184 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_fill_2 FILLER_7_252 ();
 sg13g2_fill_1 FILLER_7_254 ();
 sg13g2_fill_2 FILLER_7_290 ();
 sg13g2_fill_1 FILLER_7_292 ();
 sg13g2_decap_8 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_decap_8 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_326 ();
 sg13g2_decap_8 FILLER_7_333 ();
 sg13g2_decap_8 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_347 ();
 sg13g2_decap_8 FILLER_7_354 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_fill_2 FILLER_8_182 ();
 sg13g2_fill_1 FILLER_8_184 ();
 sg13g2_decap_4 FILLER_8_227 ();
 sg13g2_fill_2 FILLER_8_263 ();
 sg13g2_fill_1 FILLER_8_265 ();
 sg13g2_fill_2 FILLER_8_279 ();
 sg13g2_fill_1 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_163 ();
 sg13g2_decap_8 FILLER_9_170 ();
 sg13g2_decap_8 FILLER_9_177 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_4 FILLER_10_133 ();
 sg13g2_fill_1 FILLER_10_137 ();
 sg13g2_fill_2 FILLER_10_141 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_decap_8 FILLER_10_170 ();
 sg13g2_decap_8 FILLER_10_177 ();
 sg13g2_decap_8 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_191 ();
 sg13g2_decap_8 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_205 ();
 sg13g2_decap_4 FILLER_10_212 ();
 sg13g2_fill_1 FILLER_10_216 ();
 sg13g2_fill_2 FILLER_10_226 ();
 sg13g2_fill_2 FILLER_10_254 ();
 sg13g2_fill_1 FILLER_10_256 ();
 sg13g2_fill_2 FILLER_10_278 ();
 sg13g2_fill_2 FILLER_10_298 ();
 sg13g2_fill_1 FILLER_10_300 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_4 FILLER_11_126 ();
 sg13g2_fill_1 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_206 ();
 sg13g2_decap_4 FILLER_11_213 ();
 sg13g2_fill_1 FILLER_11_230 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_decap_8 FILLER_11_247 ();
 sg13g2_decap_8 FILLER_11_254 ();
 sg13g2_fill_2 FILLER_11_261 ();
 sg13g2_fill_1 FILLER_11_263 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_decap_4 FILLER_11_274 ();
 sg13g2_fill_2 FILLER_11_286 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_fill_2 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_316 ();
 sg13g2_fill_1 FILLER_11_323 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_fill_2 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_decap_8 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_8 FILLER_11_397 ();
 sg13g2_decap_4 FILLER_11_404 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_fill_1 FILLER_12_145 ();
 sg13g2_fill_2 FILLER_12_155 ();
 sg13g2_fill_1 FILLER_12_157 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_fill_2 FILLER_12_186 ();
 sg13g2_decap_4 FILLER_12_214 ();
 sg13g2_decap_4 FILLER_12_226 ();
 sg13g2_decap_8 FILLER_12_234 ();
 sg13g2_decap_4 FILLER_12_241 ();
 sg13g2_fill_1 FILLER_12_245 ();
 sg13g2_fill_1 FILLER_12_276 ();
 sg13g2_decap_8 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_293 ();
 sg13g2_decap_4 FILLER_12_300 ();
 sg13g2_fill_2 FILLER_12_304 ();
 sg13g2_fill_2 FILLER_12_327 ();
 sg13g2_fill_2 FILLER_12_337 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_4 FILLER_13_35 ();
 sg13g2_fill_1 FILLER_13_39 ();
 sg13g2_decap_8 FILLER_13_66 ();
 sg13g2_decap_8 FILLER_13_73 ();
 sg13g2_decap_8 FILLER_13_94 ();
 sg13g2_decap_8 FILLER_13_101 ();
 sg13g2_decap_8 FILLER_13_108 ();
 sg13g2_fill_1 FILLER_13_141 ();
 sg13g2_decap_8 FILLER_13_176 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_4 FILLER_13_231 ();
 sg13g2_fill_2 FILLER_13_235 ();
 sg13g2_fill_2 FILLER_13_338 ();
 sg13g2_decap_4 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_369 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_397 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_4 FILLER_14_35 ();
 sg13g2_fill_2 FILLER_14_39 ();
 sg13g2_decap_4 FILLER_14_118 ();
 sg13g2_decap_8 FILLER_14_171 ();
 sg13g2_decap_8 FILLER_14_178 ();
 sg13g2_decap_8 FILLER_14_185 ();
 sg13g2_decap_4 FILLER_14_211 ();
 sg13g2_decap_8 FILLER_14_241 ();
 sg13g2_fill_2 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_4 FILLER_15_119 ();
 sg13g2_fill_2 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_142 ();
 sg13g2_decap_8 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_169 ();
 sg13g2_fill_1 FILLER_15_176 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_fill_1 FILLER_15_219 ();
 sg13g2_decap_4 FILLER_15_248 ();
 sg13g2_fill_2 FILLER_15_252 ();
 sg13g2_fill_1 FILLER_15_263 ();
 sg13g2_fill_1 FILLER_15_273 ();
 sg13g2_fill_1 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_4 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_39 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_fill_2 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_112 ();
 sg13g2_fill_2 FILLER_16_122 ();
 sg13g2_fill_1 FILLER_16_129 ();
 sg13g2_fill_2 FILLER_16_138 ();
 sg13g2_fill_1 FILLER_16_140 ();
 sg13g2_fill_2 FILLER_16_180 ();
 sg13g2_fill_1 FILLER_16_182 ();
 sg13g2_fill_1 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_250 ();
 sg13g2_decap_4 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_fill_2 FILLER_16_287 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_355 ();
 sg13g2_decap_8 FILLER_16_362 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_decap_8 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_decap_8 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_404 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_fill_1 FILLER_17_62 ();
 sg13g2_decap_4 FILLER_17_89 ();
 sg13g2_fill_2 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_131 ();
 sg13g2_fill_2 FILLER_17_149 ();
 sg13g2_fill_1 FILLER_17_260 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_fill_1 FILLER_18_235 ();
 sg13g2_fill_2 FILLER_18_255 ();
 sg13g2_fill_1 FILLER_18_257 ();
 sg13g2_fill_1 FILLER_18_262 ();
 sg13g2_decap_4 FILLER_18_276 ();
 sg13g2_fill_1 FILLER_18_280 ();
 sg13g2_fill_2 FILLER_18_299 ();
 sg13g2_fill_1 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_35 ();
 sg13g2_fill_1 FILLER_19_37 ();
 sg13g2_fill_1 FILLER_19_43 ();
 sg13g2_fill_1 FILLER_19_75 ();
 sg13g2_decap_4 FILLER_19_86 ();
 sg13g2_fill_1 FILLER_19_90 ();
 sg13g2_fill_2 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_127 ();
 sg13g2_fill_2 FILLER_19_134 ();
 sg13g2_fill_2 FILLER_19_180 ();
 sg13g2_fill_1 FILLER_19_182 ();
 sg13g2_fill_2 FILLER_19_192 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_fill_1 FILLER_19_217 ();
 sg13g2_fill_2 FILLER_19_228 ();
 sg13g2_fill_1 FILLER_19_230 ();
 sg13g2_decap_4 FILLER_19_244 ();
 sg13g2_fill_2 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_264 ();
 sg13g2_fill_2 FILLER_19_273 ();
 sg13g2_decap_4 FILLER_19_301 ();
 sg13g2_fill_2 FILLER_19_331 ();
 sg13g2_fill_2 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_4 FILLER_20_28 ();
 sg13g2_fill_2 FILLER_20_32 ();
 sg13g2_decap_4 FILLER_20_51 ();
 sg13g2_fill_1 FILLER_20_55 ();
 sg13g2_decap_8 FILLER_20_64 ();
 sg13g2_fill_2 FILLER_20_71 ();
 sg13g2_fill_1 FILLER_20_73 ();
 sg13g2_fill_2 FILLER_20_78 ();
 sg13g2_fill_1 FILLER_20_80 ();
 sg13g2_decap_4 FILLER_20_99 ();
 sg13g2_decap_4 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_124 ();
 sg13g2_decap_8 FILLER_20_131 ();
 sg13g2_decap_8 FILLER_20_138 ();
 sg13g2_decap_8 FILLER_20_145 ();
 sg13g2_decap_8 FILLER_20_152 ();
 sg13g2_decap_8 FILLER_20_159 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_decap_8 FILLER_20_208 ();
 sg13g2_fill_2 FILLER_20_215 ();
 sg13g2_decap_4 FILLER_20_235 ();
 sg13g2_decap_4 FILLER_20_270 ();
 sg13g2_fill_1 FILLER_20_274 ();
 sg13g2_decap_4 FILLER_20_280 ();
 sg13g2_fill_2 FILLER_20_284 ();
 sg13g2_fill_2 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_108 ();
 sg13g2_fill_2 FILLER_21_171 ();
 sg13g2_decap_8 FILLER_21_199 ();
 sg13g2_decap_8 FILLER_21_206 ();
 sg13g2_decap_4 FILLER_21_213 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_278 ();
 sg13g2_fill_2 FILLER_21_285 ();
 sg13g2_decap_8 FILLER_21_310 ();
 sg13g2_decap_8 FILLER_21_317 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_374 ();
 sg13g2_decap_8 FILLER_21_381 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_4 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_61 ();
 sg13g2_decap_4 FILLER_22_68 ();
 sg13g2_decap_4 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_145 ();
 sg13g2_decap_4 FILLER_22_172 ();
 sg13g2_fill_2 FILLER_22_176 ();
 sg13g2_fill_2 FILLER_22_190 ();
 sg13g2_fill_2 FILLER_22_201 ();
 sg13g2_fill_1 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_235 ();
 sg13g2_fill_2 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_95 ();
 sg13g2_fill_1 FILLER_23_97 ();
 sg13g2_fill_1 FILLER_23_111 ();
 sg13g2_fill_2 FILLER_23_161 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_174 ();
 sg13g2_fill_1 FILLER_23_200 ();
 sg13g2_decap_4 FILLER_23_274 ();
 sg13g2_fill_2 FILLER_23_278 ();
 sg13g2_decap_8 FILLER_23_320 ();
 sg13g2_fill_1 FILLER_23_344 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_48 ();
 sg13g2_decap_8 FILLER_24_55 ();
 sg13g2_fill_2 FILLER_24_62 ();
 sg13g2_decap_4 FILLER_24_69 ();
 sg13g2_fill_2 FILLER_24_73 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_104 ();
 sg13g2_decap_4 FILLER_24_111 ();
 sg13g2_fill_1 FILLER_24_115 ();
 sg13g2_decap_4 FILLER_24_144 ();
 sg13g2_fill_2 FILLER_24_148 ();
 sg13g2_fill_2 FILLER_24_159 ();
 sg13g2_fill_2 FILLER_24_208 ();
 sg13g2_fill_1 FILLER_24_210 ();
 sg13g2_fill_2 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_220 ();
 sg13g2_fill_2 FILLER_24_230 ();
 sg13g2_decap_4 FILLER_24_273 ();
 sg13g2_fill_2 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_299 ();
 sg13g2_fill_1 FILLER_24_301 ();
 sg13g2_decap_4 FILLER_24_328 ();
 sg13g2_fill_2 FILLER_24_332 ();
 sg13g2_fill_2 FILLER_24_342 ();
 sg13g2_fill_1 FILLER_24_344 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_4 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_25 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_134 ();
 sg13g2_decap_4 FILLER_25_144 ();
 sg13g2_fill_1 FILLER_25_148 ();
 sg13g2_fill_2 FILLER_25_166 ();
 sg13g2_fill_2 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_decap_4 FILLER_25_193 ();
 sg13g2_fill_1 FILLER_25_197 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_222 ();
 sg13g2_decap_8 FILLER_25_229 ();
 sg13g2_decap_4 FILLER_25_236 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_284 ();
 sg13g2_fill_2 FILLER_25_290 ();
 sg13g2_fill_1 FILLER_25_292 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_4 FILLER_25_330 ();
 sg13g2_fill_2 FILLER_25_334 ();
 sg13g2_decap_4 FILLER_25_345 ();
 sg13g2_fill_2 FILLER_25_349 ();
 sg13g2_decap_8 FILLER_25_360 ();
 sg13g2_decap_8 FILLER_25_367 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_32 ();
 sg13g2_fill_2 FILLER_26_59 ();
 sg13g2_fill_1 FILLER_26_75 ();
 sg13g2_fill_2 FILLER_26_99 ();
 sg13g2_decap_4 FILLER_26_136 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_decap_4 FILLER_26_285 ();
 sg13g2_fill_1 FILLER_26_289 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_300 ();
 sg13g2_decap_4 FILLER_26_307 ();
 sg13g2_fill_1 FILLER_26_311 ();
 sg13g2_decap_4 FILLER_26_331 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_4 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_100 ();
 sg13g2_decap_4 FILLER_27_106 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_2 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_161 ();
 sg13g2_fill_2 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_decap_4 FILLER_27_245 ();
 sg13g2_fill_2 FILLER_27_249 ();
 sg13g2_decap_8 FILLER_27_256 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_fill_2 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_271 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_4 FILLER_27_294 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_361 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_4 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_72 ();
 sg13g2_fill_1 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_134 ();
 sg13g2_fill_2 FILLER_28_144 ();
 sg13g2_fill_2 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_28_153 ();
 sg13g2_fill_2 FILLER_28_159 ();
 sg13g2_decap_4 FILLER_28_171 ();
 sg13g2_fill_2 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_54 ();
 sg13g2_decap_8 FILLER_29_61 ();
 sg13g2_decap_4 FILLER_29_68 ();
 sg13g2_fill_2 FILLER_29_90 ();
 sg13g2_fill_2 FILLER_29_100 ();
 sg13g2_fill_1 FILLER_29_102 ();
 sg13g2_fill_1 FILLER_29_131 ();
 sg13g2_decap_4 FILLER_29_141 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_165 ();
 sg13g2_decap_4 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_185 ();
 sg13g2_fill_2 FILLER_29_209 ();
 sg13g2_decap_4 FILLER_29_220 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_312 ();
 sg13g2_decap_8 FILLER_29_319 ();
 sg13g2_decap_8 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_354 ();
 sg13g2_decap_8 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_368 ();
 sg13g2_decap_8 FILLER_29_375 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_4 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_32 ();
 sg13g2_fill_2 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_100 ();
 sg13g2_fill_2 FILLER_30_148 ();
 sg13g2_decap_8 FILLER_30_163 ();
 sg13g2_decap_8 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_decap_8 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_190 ();
 sg13g2_decap_4 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_fill_2 FILLER_30_215 ();
 sg13g2_fill_1 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_223 ();
 sg13g2_decap_4 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_decap_8 FILLER_30_325 ();
 sg13g2_decap_8 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_4 FILLER_30_346 ();
 sg13g2_decap_8 FILLER_30_359 ();
 sg13g2_decap_8 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_373 ();
 sg13g2_decap_8 FILLER_30_380 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_68 ();
 sg13g2_fill_1 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_97 ();
 sg13g2_fill_1 FILLER_31_99 ();
 sg13g2_fill_1 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_132 ();
 sg13g2_decap_4 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_fill_2 FILLER_31_173 ();
 sg13g2_fill_1 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_213 ();
 sg13g2_decap_4 FILLER_31_224 ();
 sg13g2_fill_1 FILLER_31_247 ();
 sg13g2_fill_2 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_330 ();
 sg13g2_decap_4 FILLER_31_337 ();
 sg13g2_decap_8 FILLER_31_362 ();
 sg13g2_decap_8 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_376 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_4 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_60 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_4 FILLER_32_112 ();
 sg13g2_fill_1 FILLER_32_125 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_fill_1 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_142 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_fill_1 FILLER_32_151 ();
 sg13g2_fill_2 FILLER_32_204 ();
 sg13g2_decap_4 FILLER_32_267 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_fill_2 FILLER_32_326 ();
 sg13g2_fill_1 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_32_377 ();
 sg13g2_decap_8 FILLER_32_384 ();
 sg13g2_decap_8 FILLER_32_391 ();
 sg13g2_decap_8 FILLER_32_398 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_25 ();
 sg13g2_decap_8 FILLER_33_57 ();
 sg13g2_decap_8 FILLER_33_64 ();
 sg13g2_fill_1 FILLER_33_71 ();
 sg13g2_decap_8 FILLER_33_89 ();
 sg13g2_fill_2 FILLER_33_96 ();
 sg13g2_fill_1 FILLER_33_98 ();
 sg13g2_decap_4 FILLER_33_113 ();
 sg13g2_fill_1 FILLER_33_117 ();
 sg13g2_decap_4 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_decap_4 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_182 ();
 sg13g2_fill_2 FILLER_33_193 ();
 sg13g2_fill_2 FILLER_33_213 ();
 sg13g2_fill_1 FILLER_33_215 ();
 sg13g2_fill_2 FILLER_33_294 ();
 sg13g2_fill_1 FILLER_33_300 ();
 sg13g2_decap_4 FILLER_33_318 ();
 sg13g2_fill_2 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_384 ();
 sg13g2_decap_8 FILLER_33_391 ();
 sg13g2_decap_8 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_18 ();
 sg13g2_decap_8 FILLER_34_55 ();
 sg13g2_decap_8 FILLER_34_62 ();
 sg13g2_fill_2 FILLER_34_69 ();
 sg13g2_decap_8 FILLER_34_162 ();
 sg13g2_decap_8 FILLER_34_169 ();
 sg13g2_decap_4 FILLER_34_176 ();
 sg13g2_decap_4 FILLER_34_205 ();
 sg13g2_fill_2 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_decap_4 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_278 ();
 sg13g2_decap_4 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_289 ();
 sg13g2_decap_4 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_365 ();
 sg13g2_decap_8 FILLER_34_372 ();
 sg13g2_decap_8 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_393 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_4 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_107 ();
 sg13g2_fill_1 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_136 ();
 sg13g2_fill_2 FILLER_35_168 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_192 ();
 sg13g2_decap_8 FILLER_35_199 ();
 sg13g2_fill_2 FILLER_35_206 ();
 sg13g2_fill_1 FILLER_35_208 ();
 sg13g2_decap_8 FILLER_35_227 ();
 sg13g2_decap_4 FILLER_35_234 ();
 sg13g2_decap_4 FILLER_35_270 ();
 sg13g2_fill_1 FILLER_35_274 ();
 sg13g2_decap_8 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_decap_8 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_338 ();
 sg13g2_decap_4 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_349 ();
 sg13g2_decap_8 FILLER_35_355 ();
 sg13g2_decap_8 FILLER_35_362 ();
 sg13g2_decap_8 FILLER_35_369 ();
 sg13g2_decap_8 FILLER_35_376 ();
 sg13g2_decap_8 FILLER_35_383 ();
 sg13g2_decap_8 FILLER_35_390 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_55 ();
 sg13g2_fill_2 FILLER_36_86 ();
 sg13g2_decap_8 FILLER_36_114 ();
 sg13g2_fill_2 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_149 ();
 sg13g2_fill_1 FILLER_36_199 ();
 sg13g2_decap_4 FILLER_36_240 ();
 sg13g2_fill_1 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_249 ();
 sg13g2_decap_8 FILLER_36_255 ();
 sg13g2_fill_2 FILLER_36_262 ();
 sg13g2_fill_1 FILLER_36_264 ();
 sg13g2_fill_1 FILLER_36_330 ();
 sg13g2_decap_8 FILLER_36_340 ();
 sg13g2_decap_8 FILLER_36_347 ();
 sg13g2_decap_8 FILLER_36_354 ();
 sg13g2_decap_8 FILLER_36_361 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_21 ();
 sg13g2_decap_4 FILLER_37_61 ();
 sg13g2_fill_1 FILLER_37_65 ();
 sg13g2_decap_4 FILLER_37_85 ();
 sg13g2_fill_2 FILLER_37_89 ();
 sg13g2_fill_2 FILLER_37_135 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_154 ();
 sg13g2_decap_4 FILLER_37_164 ();
 sg13g2_fill_2 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_206 ();
 sg13g2_decap_8 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_decap_4 FILLER_37_240 ();
 sg13g2_decap_8 FILLER_37_249 ();
 sg13g2_fill_1 FILLER_37_302 ();
 sg13g2_fill_2 FILLER_37_347 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_23 ();
 sg13g2_decap_8 FILLER_38_94 ();
 sg13g2_decap_4 FILLER_38_136 ();
 sg13g2_decap_8 FILLER_38_153 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_4 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_fill_1 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_4 FILLER_39_21 ();
 sg13g2_fill_1 FILLER_39_25 ();
 sg13g2_decap_4 FILLER_39_34 ();
 sg13g2_decap_4 FILLER_39_51 ();
 sg13g2_fill_2 FILLER_39_55 ();
 sg13g2_decap_8 FILLER_39_76 ();
 sg13g2_fill_1 FILLER_39_83 ();
 sg13g2_decap_8 FILLER_39_93 ();
 sg13g2_decap_8 FILLER_39_100 ();
 sg13g2_fill_2 FILLER_39_107 ();
 sg13g2_fill_2 FILLER_39_142 ();
 sg13g2_fill_1 FILLER_39_144 ();
 sg13g2_fill_1 FILLER_39_163 ();
 sg13g2_decap_8 FILLER_39_173 ();
 sg13g2_decap_4 FILLER_39_180 ();
 sg13g2_fill_1 FILLER_39_184 ();
 sg13g2_decap_8 FILLER_39_199 ();
 sg13g2_fill_2 FILLER_39_206 ();
 sg13g2_fill_1 FILLER_39_208 ();
 sg13g2_decap_8 FILLER_39_225 ();
 sg13g2_fill_2 FILLER_39_232 ();
 sg13g2_fill_1 FILLER_39_269 ();
 sg13g2_decap_4 FILLER_39_278 ();
 sg13g2_fill_2 FILLER_39_282 ();
 sg13g2_fill_1 FILLER_39_297 ();
 sg13g2_fill_2 FILLER_39_335 ();
 sg13g2_fill_1 FILLER_39_337 ();
 sg13g2_decap_8 FILLER_39_348 ();
 sg13g2_decap_8 FILLER_39_373 ();
 sg13g2_decap_8 FILLER_39_380 ();
 sg13g2_decap_8 FILLER_39_387 ();
 sg13g2_decap_8 FILLER_39_394 ();
 sg13g2_decap_8 FILLER_39_401 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_fill_2 FILLER_40_28 ();
 sg13g2_fill_1 FILLER_40_59 ();
 sg13g2_fill_2 FILLER_40_83 ();
 sg13g2_fill_1 FILLER_40_85 ();
 sg13g2_fill_1 FILLER_40_91 ();
 sg13g2_fill_2 FILLER_40_102 ();
 sg13g2_fill_1 FILLER_40_109 ();
 sg13g2_fill_2 FILLER_40_114 ();
 sg13g2_fill_1 FILLER_40_116 ();
 sg13g2_decap_4 FILLER_40_122 ();
 sg13g2_decap_4 FILLER_40_135 ();
 sg13g2_fill_2 FILLER_40_147 ();
 sg13g2_fill_1 FILLER_40_175 ();
 sg13g2_fill_2 FILLER_40_228 ();
 sg13g2_fill_2 FILLER_40_240 ();
 sg13g2_fill_1 FILLER_40_242 ();
 sg13g2_fill_2 FILLER_40_248 ();
 sg13g2_decap_4 FILLER_40_258 ();
 sg13g2_fill_1 FILLER_40_262 ();
 sg13g2_decap_8 FILLER_40_272 ();
 sg13g2_fill_1 FILLER_40_279 ();
 sg13g2_fill_2 FILLER_40_288 ();
 sg13g2_fill_2 FILLER_40_305 ();
 sg13g2_fill_1 FILLER_40_307 ();
 sg13g2_decap_4 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_369 ();
 sg13g2_decap_8 FILLER_40_376 ();
 sg13g2_decap_8 FILLER_40_383 ();
 sg13g2_decap_8 FILLER_40_390 ();
 sg13g2_decap_8 FILLER_40_397 ();
 sg13g2_decap_4 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_4 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_18 ();
 sg13g2_decap_4 FILLER_41_77 ();
 sg13g2_fill_1 FILLER_41_116 ();
 sg13g2_fill_2 FILLER_41_132 ();
 sg13g2_decap_4 FILLER_41_184 ();
 sg13g2_fill_2 FILLER_41_188 ();
 sg13g2_decap_8 FILLER_41_264 ();
 sg13g2_decap_8 FILLER_41_271 ();
 sg13g2_decap_4 FILLER_41_278 ();
 sg13g2_fill_2 FILLER_41_299 ();
 sg13g2_fill_2 FILLER_41_308 ();
 sg13g2_fill_1 FILLER_41_310 ();
 sg13g2_decap_8 FILLER_41_355 ();
 sg13g2_decap_8 FILLER_41_362 ();
 sg13g2_decap_8 FILLER_41_369 ();
 sg13g2_decap_8 FILLER_41_376 ();
 sg13g2_decap_8 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_4 FILLER_42_21 ();
 sg13g2_fill_2 FILLER_42_25 ();
 sg13g2_fill_2 FILLER_42_66 ();
 sg13g2_fill_1 FILLER_42_68 ();
 sg13g2_fill_2 FILLER_42_85 ();
 sg13g2_fill_2 FILLER_42_96 ();
 sg13g2_fill_1 FILLER_42_98 ();
 sg13g2_decap_4 FILLER_42_151 ();
 sg13g2_fill_2 FILLER_42_155 ();
 sg13g2_decap_4 FILLER_42_209 ();
 sg13g2_fill_2 FILLER_42_241 ();
 sg13g2_fill_1 FILLER_42_243 ();
 sg13g2_fill_1 FILLER_42_363 ();
 sg13g2_decap_8 FILLER_42_373 ();
 sg13g2_decap_8 FILLER_42_380 ();
 sg13g2_decap_8 FILLER_42_387 ();
 sg13g2_decap_8 FILLER_42_394 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_4 FILLER_43_28 ();
 sg13g2_fill_1 FILLER_43_32 ();
 sg13g2_decap_8 FILLER_43_45 ();
 sg13g2_decap_8 FILLER_43_52 ();
 sg13g2_fill_2 FILLER_43_59 ();
 sg13g2_fill_2 FILLER_43_114 ();
 sg13g2_fill_2 FILLER_43_125 ();
 sg13g2_fill_2 FILLER_43_163 ();
 sg13g2_fill_1 FILLER_43_165 ();
 sg13g2_decap_4 FILLER_43_175 ();
 sg13g2_fill_1 FILLER_43_179 ();
 sg13g2_decap_4 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_4 FILLER_43_210 ();
 sg13g2_decap_4 FILLER_43_250 ();
 sg13g2_fill_1 FILLER_43_254 ();
 sg13g2_decap_8 FILLER_43_291 ();
 sg13g2_fill_2 FILLER_43_298 ();
 sg13g2_fill_1 FILLER_43_300 ();
 sg13g2_fill_1 FILLER_43_309 ();
 sg13g2_decap_4 FILLER_43_343 ();
 sg13g2_fill_1 FILLER_43_347 ();
 sg13g2_decap_8 FILLER_43_374 ();
 sg13g2_decap_8 FILLER_43_381 ();
 sg13g2_decap_8 FILLER_43_388 ();
 sg13g2_decap_8 FILLER_43_395 ();
 sg13g2_decap_8 FILLER_43_402 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_4 FILLER_44_56 ();
 sg13g2_fill_2 FILLER_44_60 ();
 sg13g2_decap_8 FILLER_44_66 ();
 sg13g2_decap_4 FILLER_44_73 ();
 sg13g2_fill_2 FILLER_44_112 ();
 sg13g2_decap_4 FILLER_44_128 ();
 sg13g2_fill_1 FILLER_44_132 ();
 sg13g2_fill_2 FILLER_44_160 ();
 sg13g2_fill_1 FILLER_44_162 ();
 sg13g2_decap_4 FILLER_44_168 ();
 sg13g2_fill_2 FILLER_44_190 ();
 sg13g2_decap_4 FILLER_44_201 ();
 sg13g2_fill_2 FILLER_44_205 ();
 sg13g2_decap_8 FILLER_44_212 ();
 sg13g2_fill_1 FILLER_44_219 ();
 sg13g2_decap_4 FILLER_44_265 ();
 sg13g2_decap_8 FILLER_44_286 ();
 sg13g2_decap_8 FILLER_44_293 ();
 sg13g2_decap_8 FILLER_44_300 ();
 sg13g2_fill_2 FILLER_44_307 ();
 sg13g2_decap_8 FILLER_44_314 ();
 sg13g2_decap_8 FILLER_44_326 ();
 sg13g2_decap_8 FILLER_44_333 ();
 sg13g2_decap_8 FILLER_44_340 ();
 sg13g2_decap_8 FILLER_44_347 ();
 sg13g2_fill_1 FILLER_44_354 ();
 sg13g2_decap_8 FILLER_44_366 ();
 sg13g2_decap_8 FILLER_44_373 ();
 sg13g2_decap_8 FILLER_44_380 ();
 sg13g2_decap_8 FILLER_44_387 ();
 sg13g2_decap_8 FILLER_44_394 ();
 sg13g2_decap_8 FILLER_44_401 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_4 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_37 ();
 sg13g2_decap_8 FILLER_45_44 ();
 sg13g2_decap_4 FILLER_45_51 ();
 sg13g2_fill_2 FILLER_45_55 ();
 sg13g2_fill_2 FILLER_45_62 ();
 sg13g2_fill_1 FILLER_45_64 ();
 sg13g2_fill_2 FILLER_45_70 ();
 sg13g2_fill_1 FILLER_45_72 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_fill_2 FILLER_45_84 ();
 sg13g2_fill_1 FILLER_45_86 ();
 sg13g2_decap_4 FILLER_45_117 ();
 sg13g2_decap_8 FILLER_45_139 ();
 sg13g2_decap_8 FILLER_45_146 ();
 sg13g2_decap_4 FILLER_45_153 ();
 sg13g2_fill_1 FILLER_45_157 ();
 sg13g2_fill_2 FILLER_45_162 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_fill_1 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_258 ();
 sg13g2_fill_1 FILLER_45_265 ();
 sg13g2_decap_8 FILLER_45_279 ();
 sg13g2_decap_8 FILLER_45_286 ();
 sg13g2_fill_2 FILLER_45_293 ();
 sg13g2_decap_8 FILLER_45_303 ();
 sg13g2_fill_2 FILLER_45_310 ();
 sg13g2_fill_1 FILLER_45_312 ();
 sg13g2_fill_2 FILLER_45_326 ();
 sg13g2_fill_1 FILLER_45_328 ();
 sg13g2_decap_4 FILLER_45_337 ();
 sg13g2_fill_1 FILLER_45_349 ();
 sg13g2_decap_8 FILLER_45_368 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_8 FILLER_45_382 ();
 sg13g2_decap_8 FILLER_45_389 ();
 sg13g2_decap_8 FILLER_45_396 ();
 sg13g2_decap_4 FILLER_45_403 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_fill_1 FILLER_46_38 ();
 sg13g2_decap_8 FILLER_46_89 ();
 sg13g2_decap_4 FILLER_46_96 ();
 sg13g2_fill_1 FILLER_46_100 ();
 sg13g2_decap_4 FILLER_46_110 ();
 sg13g2_decap_4 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_229 ();
 sg13g2_fill_2 FILLER_46_236 ();
 sg13g2_fill_1 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_248 ();
 sg13g2_fill_1 FILLER_46_255 ();
 sg13g2_decap_4 FILLER_46_275 ();
 sg13g2_decap_4 FILLER_46_284 ();
 sg13g2_fill_2 FILLER_46_316 ();
 sg13g2_decap_4 FILLER_46_344 ();
 sg13g2_decap_8 FILLER_46_383 ();
 sg13g2_decap_8 FILLER_46_390 ();
 sg13g2_decap_8 FILLER_46_397 ();
 sg13g2_decap_4 FILLER_46_404 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_4 FILLER_47_14 ();
 sg13g2_fill_2 FILLER_47_18 ();
 sg13g2_fill_2 FILLER_47_50 ();
 sg13g2_fill_1 FILLER_47_52 ();
 sg13g2_decap_8 FILLER_47_100 ();
 sg13g2_fill_2 FILLER_47_117 ();
 sg13g2_fill_2 FILLER_47_135 ();
 sg13g2_fill_1 FILLER_47_137 ();
 sg13g2_decap_8 FILLER_47_221 ();
 sg13g2_decap_8 FILLER_47_228 ();
 sg13g2_decap_8 FILLER_47_235 ();
 sg13g2_fill_2 FILLER_47_242 ();
 sg13g2_fill_1 FILLER_47_280 ();
 sg13g2_decap_4 FILLER_47_286 ();
 sg13g2_fill_2 FILLER_47_351 ();
 sg13g2_fill_1 FILLER_47_353 ();
 sg13g2_decap_8 FILLER_47_362 ();
 sg13g2_decap_8 FILLER_47_369 ();
 sg13g2_decap_8 FILLER_47_376 ();
 sg13g2_decap_8 FILLER_47_383 ();
 sg13g2_decap_8 FILLER_47_390 ();
 sg13g2_decap_8 FILLER_47_397 ();
 sg13g2_decap_4 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_fill_1 FILLER_48_21 ();
 sg13g2_decap_4 FILLER_48_44 ();
 sg13g2_fill_1 FILLER_48_48 ();
 sg13g2_fill_1 FILLER_48_59 ();
 sg13g2_fill_2 FILLER_48_78 ();
 sg13g2_decap_8 FILLER_48_88 ();
 sg13g2_fill_1 FILLER_48_95 ();
 sg13g2_decap_4 FILLER_48_105 ();
 sg13g2_fill_1 FILLER_48_109 ();
 sg13g2_fill_2 FILLER_48_122 ();
 sg13g2_decap_8 FILLER_48_137 ();
 sg13g2_fill_2 FILLER_48_158 ();
 sg13g2_fill_1 FILLER_48_160 ();
 sg13g2_fill_1 FILLER_48_179 ();
 sg13g2_decap_8 FILLER_48_195 ();
 sg13g2_decap_4 FILLER_48_202 ();
 sg13g2_fill_2 FILLER_48_206 ();
 sg13g2_decap_4 FILLER_48_216 ();
 sg13g2_fill_1 FILLER_48_220 ();
 sg13g2_decap_8 FILLER_48_236 ();
 sg13g2_decap_4 FILLER_48_243 ();
 sg13g2_decap_8 FILLER_48_338 ();
 sg13g2_decap_4 FILLER_48_345 ();
 sg13g2_decap_8 FILLER_48_354 ();
 sg13g2_decap_8 FILLER_48_361 ();
 sg13g2_decap_8 FILLER_48_368 ();
 sg13g2_decap_8 FILLER_48_375 ();
 sg13g2_decap_8 FILLER_48_382 ();
 sg13g2_decap_8 FILLER_48_389 ();
 sg13g2_decap_8 FILLER_48_396 ();
 sg13g2_decap_4 FILLER_48_403 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_4 FILLER_49_21 ();
 sg13g2_fill_2 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_44 ();
 sg13g2_fill_1 FILLER_49_51 ();
 sg13g2_decap_8 FILLER_49_69 ();
 sg13g2_fill_2 FILLER_49_76 ();
 sg13g2_fill_2 FILLER_49_83 ();
 sg13g2_decap_4 FILLER_49_165 ();
 sg13g2_decap_4 FILLER_49_191 ();
 sg13g2_fill_2 FILLER_49_195 ();
 sg13g2_fill_1 FILLER_49_207 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_fill_2 FILLER_49_266 ();
 sg13g2_decap_4 FILLER_49_273 ();
 sg13g2_fill_1 FILLER_49_277 ();
 sg13g2_decap_4 FILLER_49_282 ();
 sg13g2_fill_2 FILLER_49_286 ();
 sg13g2_decap_4 FILLER_49_314 ();
 sg13g2_fill_2 FILLER_49_318 ();
 sg13g2_fill_2 FILLER_49_325 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_4 FILLER_50_21 ();
 sg13g2_fill_2 FILLER_50_25 ();
 sg13g2_decap_8 FILLER_50_61 ();
 sg13g2_fill_2 FILLER_50_68 ();
 sg13g2_decap_8 FILLER_50_83 ();
 sg13g2_decap_8 FILLER_50_99 ();
 sg13g2_decap_8 FILLER_50_106 ();
 sg13g2_decap_8 FILLER_50_113 ();
 sg13g2_decap_8 FILLER_50_120 ();
 sg13g2_decap_4 FILLER_50_127 ();
 sg13g2_fill_2 FILLER_50_131 ();
 sg13g2_fill_1 FILLER_50_142 ();
 sg13g2_fill_2 FILLER_50_195 ();
 sg13g2_fill_2 FILLER_50_205 ();
 sg13g2_decap_8 FILLER_50_265 ();
 sg13g2_fill_1 FILLER_50_272 ();
 sg13g2_decap_8 FILLER_50_282 ();
 sg13g2_decap_8 FILLER_50_289 ();
 sg13g2_fill_2 FILLER_50_296 ();
 sg13g2_fill_1 FILLER_50_298 ();
 sg13g2_decap_8 FILLER_50_304 ();
 sg13g2_fill_2 FILLER_50_311 ();
 sg13g2_decap_8 FILLER_50_318 ();
 sg13g2_fill_2 FILLER_50_325 ();
 sg13g2_decap_8 FILLER_50_375 ();
 sg13g2_decap_8 FILLER_50_382 ();
 sg13g2_decap_8 FILLER_50_389 ();
 sg13g2_decap_8 FILLER_50_396 ();
 sg13g2_decap_4 FILLER_50_403 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_4 FILLER_51_21 ();
 sg13g2_fill_2 FILLER_51_30 ();
 sg13g2_fill_1 FILLER_51_32 ();
 sg13g2_fill_1 FILLER_51_46 ();
 sg13g2_decap_4 FILLER_51_73 ();
 sg13g2_fill_1 FILLER_51_77 ();
 sg13g2_fill_2 FILLER_51_86 ();
 sg13g2_fill_1 FILLER_51_88 ();
 sg13g2_fill_2 FILLER_51_117 ();
 sg13g2_fill_1 FILLER_51_127 ();
 sg13g2_fill_1 FILLER_51_137 ();
 sg13g2_decap_4 FILLER_51_142 ();
 sg13g2_fill_1 FILLER_51_146 ();
 sg13g2_fill_2 FILLER_51_157 ();
 sg13g2_fill_1 FILLER_51_159 ();
 sg13g2_decap_8 FILLER_51_169 ();
 sg13g2_fill_2 FILLER_51_199 ();
 sg13g2_fill_2 FILLER_51_218 ();
 sg13g2_fill_1 FILLER_51_246 ();
 sg13g2_decap_8 FILLER_51_276 ();
 sg13g2_decap_8 FILLER_51_283 ();
 sg13g2_decap_4 FILLER_51_290 ();
 sg13g2_fill_1 FILLER_51_294 ();
 sg13g2_decap_8 FILLER_51_303 ();
 sg13g2_decap_8 FILLER_51_310 ();
 sg13g2_decap_4 FILLER_51_317 ();
 sg13g2_fill_2 FILLER_51_321 ();
 sg13g2_decap_8 FILLER_51_385 ();
 sg13g2_decap_8 FILLER_51_392 ();
 sg13g2_decap_8 FILLER_51_399 ();
 sg13g2_fill_2 FILLER_51_406 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_14 ();
 sg13g2_fill_1 FILLER_52_18 ();
 sg13g2_decap_8 FILLER_52_45 ();
 sg13g2_fill_1 FILLER_52_52 ();
 sg13g2_fill_2 FILLER_52_79 ();
 sg13g2_fill_2 FILLER_52_112 ();
 sg13g2_fill_1 FILLER_52_114 ();
 sg13g2_decap_8 FILLER_52_150 ();
 sg13g2_decap_4 FILLER_52_157 ();
 sg13g2_fill_1 FILLER_52_161 ();
 sg13g2_fill_1 FILLER_52_176 ();
 sg13g2_fill_2 FILLER_52_188 ();
 sg13g2_fill_1 FILLER_52_190 ();
 sg13g2_decap_4 FILLER_52_279 ();
 sg13g2_fill_1 FILLER_52_288 ();
 sg13g2_fill_2 FILLER_52_331 ();
 sg13g2_decap_8 FILLER_52_351 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_fill_2 FILLER_52_406 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_7 ();
 sg13g2_decap_4 FILLER_53_46 ();
 sg13g2_fill_1 FILLER_53_50 ();
 sg13g2_fill_2 FILLER_53_61 ();
 sg13g2_fill_1 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_74 ();
 sg13g2_fill_2 FILLER_53_117 ();
 sg13g2_decap_4 FILLER_53_185 ();
 sg13g2_fill_2 FILLER_53_189 ();
 sg13g2_fill_1 FILLER_53_195 ();
 sg13g2_fill_2 FILLER_53_213 ();
 sg13g2_fill_1 FILLER_53_233 ();
 sg13g2_decap_4 FILLER_53_243 ();
 sg13g2_fill_2 FILLER_53_247 ();
 sg13g2_fill_1 FILLER_53_254 ();
 sg13g2_fill_1 FILLER_53_291 ();
 sg13g2_fill_2 FILLER_53_327 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_fill_2 FILLER_53_373 ();
 sg13g2_decap_8 FILLER_53_384 ();
 sg13g2_decap_8 FILLER_53_391 ();
 sg13g2_decap_8 FILLER_53_398 ();
 sg13g2_decap_4 FILLER_53_405 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_11 ();
 sg13g2_fill_1 FILLER_54_48 ();
 sg13g2_fill_2 FILLER_54_67 ();
 sg13g2_decap_8 FILLER_54_148 ();
 sg13g2_decap_4 FILLER_54_155 ();
 sg13g2_fill_1 FILLER_54_159 ();
 sg13g2_fill_2 FILLER_54_168 ();
 sg13g2_fill_1 FILLER_54_170 ();
 sg13g2_fill_2 FILLER_54_179 ();
 sg13g2_decap_8 FILLER_54_190 ();
 sg13g2_decap_4 FILLER_54_206 ();
 sg13g2_fill_2 FILLER_54_210 ();
 sg13g2_decap_4 FILLER_54_295 ();
 sg13g2_fill_1 FILLER_54_328 ();
 sg13g2_fill_1 FILLER_54_353 ();
 sg13g2_fill_1 FILLER_54_367 ();
 sg13g2_decap_8 FILLER_54_377 ();
 sg13g2_decap_8 FILLER_54_384 ();
 sg13g2_decap_8 FILLER_54_391 ();
 sg13g2_decap_8 FILLER_54_398 ();
 sg13g2_decap_4 FILLER_54_405 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_4 FILLER_55_21 ();
 sg13g2_fill_2 FILLER_55_35 ();
 sg13g2_fill_1 FILLER_55_51 ();
 sg13g2_decap_8 FILLER_55_62 ();
 sg13g2_decap_4 FILLER_55_69 ();
 sg13g2_decap_8 FILLER_55_78 ();
 sg13g2_decap_8 FILLER_55_85 ();
 sg13g2_decap_4 FILLER_55_92 ();
 sg13g2_fill_1 FILLER_55_96 ();
 sg13g2_fill_2 FILLER_55_106 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_fill_2 FILLER_55_151 ();
 sg13g2_decap_4 FILLER_55_179 ();
 sg13g2_decap_4 FILLER_55_186 ();
 sg13g2_fill_1 FILLER_55_190 ();
 sg13g2_fill_1 FILLER_55_201 ();
 sg13g2_decap_4 FILLER_55_215 ();
 sg13g2_fill_1 FILLER_55_219 ();
 sg13g2_decap_8 FILLER_55_240 ();
 sg13g2_fill_1 FILLER_55_247 ();
 sg13g2_fill_1 FILLER_55_284 ();
 sg13g2_fill_2 FILLER_55_294 ();
 sg13g2_fill_2 FILLER_55_305 ();
 sg13g2_decap_4 FILLER_55_335 ();
 sg13g2_decap_8 FILLER_55_379 ();
 sg13g2_decap_8 FILLER_55_386 ();
 sg13g2_decap_8 FILLER_55_393 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_fill_2 FILLER_56_14 ();
 sg13g2_fill_1 FILLER_56_16 ();
 sg13g2_decap_4 FILLER_56_99 ();
 sg13g2_fill_1 FILLER_56_103 ();
 sg13g2_decap_8 FILLER_56_109 ();
 sg13g2_decap_8 FILLER_56_116 ();
 sg13g2_decap_8 FILLER_56_123 ();
 sg13g2_decap_8 FILLER_56_130 ();
 sg13g2_fill_1 FILLER_56_178 ();
 sg13g2_decap_8 FILLER_56_199 ();
 sg13g2_decap_4 FILLER_56_206 ();
 sg13g2_fill_2 FILLER_56_210 ();
 sg13g2_decap_4 FILLER_56_256 ();
 sg13g2_fill_2 FILLER_56_260 ();
 sg13g2_decap_4 FILLER_56_283 ();
 sg13g2_fill_1 FILLER_56_287 ();
 sg13g2_decap_4 FILLER_56_292 ();
 sg13g2_fill_1 FILLER_56_296 ();
 sg13g2_decap_4 FILLER_56_349 ();
 sg13g2_decap_8 FILLER_56_388 ();
 sg13g2_decap_8 FILLER_56_395 ();
 sg13g2_decap_8 FILLER_56_402 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_21 ();
 sg13g2_fill_1 FILLER_57_97 ();
 sg13g2_fill_2 FILLER_57_111 ();
 sg13g2_fill_1 FILLER_57_113 ();
 sg13g2_fill_1 FILLER_57_122 ();
 sg13g2_fill_2 FILLER_57_149 ();
 sg13g2_fill_1 FILLER_57_151 ();
 sg13g2_fill_2 FILLER_57_169 ();
 sg13g2_fill_1 FILLER_57_171 ();
 sg13g2_decap_8 FILLER_57_187 ();
 sg13g2_decap_8 FILLER_57_194 ();
 sg13g2_decap_8 FILLER_57_204 ();
 sg13g2_decap_4 FILLER_57_211 ();
 sg13g2_fill_2 FILLER_57_215 ();
 sg13g2_decap_8 FILLER_57_226 ();
 sg13g2_decap_4 FILLER_57_233 ();
 sg13g2_fill_1 FILLER_57_237 ();
 sg13g2_fill_2 FILLER_57_262 ();
 sg13g2_fill_1 FILLER_57_264 ();
 sg13g2_fill_2 FILLER_57_306 ();
 sg13g2_decap_8 FILLER_57_387 ();
 sg13g2_decap_8 FILLER_57_394 ();
 sg13g2_decap_8 FILLER_57_401 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_fill_1 FILLER_58_21 ();
 sg13g2_fill_2 FILLER_58_48 ();
 sg13g2_decap_4 FILLER_58_59 ();
 sg13g2_fill_2 FILLER_58_63 ();
 sg13g2_fill_2 FILLER_58_75 ();
 sg13g2_fill_2 FILLER_58_112 ();
 sg13g2_fill_1 FILLER_58_114 ();
 sg13g2_decap_4 FILLER_58_162 ();
 sg13g2_fill_2 FILLER_58_166 ();
 sg13g2_fill_1 FILLER_58_203 ();
 sg13g2_decap_4 FILLER_58_231 ();
 sg13g2_fill_1 FILLER_58_235 ();
 sg13g2_fill_1 FILLER_58_293 ();
 sg13g2_fill_2 FILLER_58_343 ();
 sg13g2_fill_1 FILLER_58_345 ();
 sg13g2_decap_8 FILLER_58_380 ();
 sg13g2_decap_8 FILLER_58_387 ();
 sg13g2_decap_8 FILLER_58_394 ();
 sg13g2_decap_8 FILLER_58_401 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_fill_2 FILLER_59_21 ();
 sg13g2_decap_4 FILLER_59_48 ();
 sg13g2_decap_4 FILLER_59_61 ();
 sg13g2_fill_1 FILLER_59_65 ();
 sg13g2_decap_8 FILLER_59_83 ();
 sg13g2_decap_8 FILLER_59_90 ();
 sg13g2_decap_4 FILLER_59_97 ();
 sg13g2_fill_2 FILLER_59_101 ();
 sg13g2_fill_2 FILLER_59_117 ();
 sg13g2_fill_1 FILLER_59_119 ();
 sg13g2_fill_2 FILLER_59_138 ();
 sg13g2_decap_8 FILLER_59_153 ();
 sg13g2_decap_4 FILLER_59_160 ();
 sg13g2_fill_1 FILLER_59_164 ();
 sg13g2_decap_8 FILLER_59_236 ();
 sg13g2_decap_4 FILLER_59_243 ();
 sg13g2_fill_1 FILLER_59_275 ();
 sg13g2_decap_4 FILLER_59_302 ();
 sg13g2_fill_1 FILLER_59_306 ();
 sg13g2_fill_1 FILLER_59_316 ();
 sg13g2_decap_4 FILLER_59_321 ();
 sg13g2_decap_8 FILLER_59_378 ();
 sg13g2_decap_8 FILLER_59_385 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_399 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_fill_2 FILLER_60_21 ();
 sg13g2_fill_2 FILLER_60_46 ();
 sg13g2_decap_4 FILLER_60_83 ();
 sg13g2_fill_2 FILLER_60_87 ();
 sg13g2_decap_8 FILLER_60_99 ();
 sg13g2_decap_8 FILLER_60_106 ();
 sg13g2_fill_2 FILLER_60_113 ();
 sg13g2_decap_8 FILLER_60_129 ();
 sg13g2_fill_2 FILLER_60_136 ();
 sg13g2_decap_8 FILLER_60_142 ();
 sg13g2_decap_4 FILLER_60_149 ();
 sg13g2_fill_2 FILLER_60_153 ();
 sg13g2_fill_1 FILLER_60_164 ();
 sg13g2_fill_2 FILLER_60_170 ();
 sg13g2_decap_4 FILLER_60_184 ();
 sg13g2_fill_2 FILLER_60_201 ();
 sg13g2_fill_1 FILLER_60_203 ();
 sg13g2_fill_1 FILLER_60_218 ();
 sg13g2_fill_2 FILLER_60_260 ();
 sg13g2_fill_1 FILLER_60_262 ();
 sg13g2_decap_8 FILLER_60_294 ();
 sg13g2_decap_4 FILLER_60_301 ();
 sg13g2_decap_4 FILLER_60_310 ();
 sg13g2_fill_1 FILLER_60_314 ();
 sg13g2_fill_1 FILLER_60_324 ();
 sg13g2_decap_8 FILLER_60_330 ();
 sg13g2_decap_8 FILLER_60_337 ();
 sg13g2_decap_8 FILLER_60_344 ();
 sg13g2_decap_8 FILLER_60_359 ();
 sg13g2_decap_8 FILLER_60_366 ();
 sg13g2_decap_8 FILLER_60_373 ();
 sg13g2_decap_8 FILLER_60_380 ();
 sg13g2_decap_8 FILLER_60_387 ();
 sg13g2_decap_8 FILLER_60_394 ();
 sg13g2_decap_8 FILLER_60_401 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_4 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_11 ();
 sg13g2_decap_4 FILLER_61_113 ();
 sg13g2_decap_4 FILLER_61_122 ();
 sg13g2_fill_2 FILLER_61_136 ();
 sg13g2_decap_4 FILLER_61_209 ();
 sg13g2_fill_2 FILLER_61_244 ();
 sg13g2_fill_1 FILLER_61_246 ();
 sg13g2_fill_1 FILLER_61_329 ();
 sg13g2_decap_8 FILLER_61_356 ();
 sg13g2_decap_8 FILLER_61_363 ();
 sg13g2_decap_8 FILLER_61_370 ();
 sg13g2_decap_8 FILLER_61_377 ();
 sg13g2_decap_8 FILLER_61_384 ();
 sg13g2_decap_8 FILLER_61_391 ();
 sg13g2_decap_8 FILLER_61_398 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_fill_1 FILLER_62_54 ();
 sg13g2_fill_2 FILLER_62_65 ();
 sg13g2_fill_2 FILLER_62_77 ();
 sg13g2_decap_4 FILLER_62_88 ();
 sg13g2_fill_1 FILLER_62_92 ();
 sg13g2_decap_8 FILLER_62_150 ();
 sg13g2_decap_8 FILLER_62_157 ();
 sg13g2_fill_2 FILLER_62_164 ();
 sg13g2_decap_8 FILLER_62_195 ();
 sg13g2_decap_4 FILLER_62_210 ();
 sg13g2_fill_2 FILLER_62_214 ();
 sg13g2_decap_4 FILLER_62_231 ();
 sg13g2_decap_8 FILLER_62_244 ();
 sg13g2_decap_8 FILLER_62_251 ();
 sg13g2_decap_8 FILLER_62_289 ();
 sg13g2_decap_4 FILLER_62_296 ();
 sg13g2_fill_2 FILLER_62_309 ();
 sg13g2_fill_1 FILLER_62_311 ();
 sg13g2_decap_8 FILLER_62_356 ();
 sg13g2_decap_8 FILLER_62_363 ();
 sg13g2_decap_8 FILLER_62_370 ();
 sg13g2_decap_8 FILLER_62_377 ();
 sg13g2_decap_8 FILLER_62_384 ();
 sg13g2_decap_8 FILLER_62_391 ();
 sg13g2_decap_8 FILLER_62_398 ();
 sg13g2_decap_4 FILLER_62_405 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_48 ();
 sg13g2_decap_4 FILLER_63_55 ();
 sg13g2_fill_1 FILLER_63_59 ();
 sg13g2_decap_4 FILLER_63_92 ();
 sg13g2_fill_1 FILLER_63_106 ();
 sg13g2_fill_2 FILLER_63_125 ();
 sg13g2_fill_2 FILLER_63_162 ();
 sg13g2_fill_1 FILLER_63_164 ();
 sg13g2_decap_8 FILLER_63_236 ();
 sg13g2_fill_1 FILLER_63_243 ();
 sg13g2_fill_2 FILLER_63_263 ();
 sg13g2_fill_2 FILLER_63_284 ();
 sg13g2_fill_1 FILLER_63_286 ();
 sg13g2_fill_2 FILLER_63_313 ();
 sg13g2_fill_1 FILLER_63_323 ();
 sg13g2_decap_8 FILLER_63_352 ();
 sg13g2_decap_8 FILLER_63_359 ();
 sg13g2_decap_8 FILLER_63_366 ();
 sg13g2_decap_8 FILLER_63_373 ();
 sg13g2_decap_8 FILLER_63_380 ();
 sg13g2_decap_8 FILLER_63_387 ();
 sg13g2_decap_8 FILLER_63_394 ();
 sg13g2_decap_8 FILLER_63_401 ();
 sg13g2_fill_1 FILLER_63_408 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_4 FILLER_64_28 ();
 sg13g2_fill_2 FILLER_64_32 ();
 sg13g2_fill_1 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_48 ();
 sg13g2_decap_8 FILLER_64_55 ();
 sg13g2_fill_2 FILLER_64_62 ();
 sg13g2_decap_8 FILLER_64_99 ();
 sg13g2_decap_4 FILLER_64_106 ();
 sg13g2_fill_2 FILLER_64_135 ();
 sg13g2_decap_8 FILLER_64_146 ();
 sg13g2_fill_1 FILLER_64_192 ();
 sg13g2_fill_2 FILLER_64_207 ();
 sg13g2_fill_1 FILLER_64_209 ();
 sg13g2_decap_4 FILLER_64_214 ();
 sg13g2_fill_1 FILLER_64_218 ();
 sg13g2_fill_1 FILLER_64_228 ();
 sg13g2_fill_2 FILLER_64_319 ();
 sg13g2_fill_1 FILLER_64_321 ();
 sg13g2_decap_8 FILLER_64_331 ();
 sg13g2_decap_4 FILLER_64_338 ();
 sg13g2_decap_8 FILLER_64_351 ();
 sg13g2_decap_8 FILLER_64_358 ();
 sg13g2_decap_8 FILLER_64_365 ();
 sg13g2_decap_8 FILLER_64_372 ();
 sg13g2_decap_8 FILLER_64_379 ();
 sg13g2_decap_8 FILLER_64_386 ();
 sg13g2_decap_8 FILLER_64_393 ();
 sg13g2_decap_8 FILLER_64_400 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_4 FILLER_65_28 ();
 sg13g2_fill_2 FILLER_65_32 ();
 sg13g2_fill_1 FILLER_65_64 ();
 sg13g2_fill_2 FILLER_65_73 ();
 sg13g2_fill_1 FILLER_65_75 ();
 sg13g2_fill_2 FILLER_65_81 ();
 sg13g2_fill_1 FILLER_65_114 ();
 sg13g2_fill_1 FILLER_65_125 ();
 sg13g2_fill_2 FILLER_65_130 ();
 sg13g2_fill_1 FILLER_65_141 ();
 sg13g2_decap_8 FILLER_65_150 ();
 sg13g2_fill_2 FILLER_65_157 ();
 sg13g2_decap_8 FILLER_65_172 ();
 sg13g2_fill_1 FILLER_65_202 ();
 sg13g2_decap_8 FILLER_65_207 ();
 sg13g2_decap_8 FILLER_65_214 ();
 sg13g2_fill_1 FILLER_65_221 ();
 sg13g2_fill_2 FILLER_65_228 ();
 sg13g2_fill_2 FILLER_65_283 ();
 sg13g2_fill_1 FILLER_65_285 ();
 sg13g2_decap_8 FILLER_65_305 ();
 sg13g2_fill_2 FILLER_65_312 ();
 sg13g2_fill_2 FILLER_65_327 ();
 sg13g2_decap_8 FILLER_65_355 ();
 sg13g2_decap_8 FILLER_65_362 ();
 sg13g2_decap_8 FILLER_65_369 ();
 sg13g2_decap_8 FILLER_65_376 ();
 sg13g2_decap_8 FILLER_65_383 ();
 sg13g2_decap_8 FILLER_65_390 ();
 sg13g2_decap_8 FILLER_65_397 ();
 sg13g2_decap_4 FILLER_65_404 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_4 FILLER_66_14 ();
 sg13g2_fill_2 FILLER_66_18 ();
 sg13g2_fill_1 FILLER_66_128 ();
 sg13g2_decap_8 FILLER_66_156 ();
 sg13g2_fill_1 FILLER_66_163 ();
 sg13g2_decap_8 FILLER_66_177 ();
 sg13g2_decap_4 FILLER_66_184 ();
 sg13g2_fill_1 FILLER_66_188 ();
 sg13g2_fill_2 FILLER_66_207 ();
 sg13g2_fill_1 FILLER_66_209 ();
 sg13g2_fill_2 FILLER_66_236 ();
 sg13g2_fill_1 FILLER_66_295 ();
 sg13g2_decap_4 FILLER_66_306 ();
 sg13g2_decap_8 FILLER_66_354 ();
 sg13g2_decap_8 FILLER_66_361 ();
 sg13g2_decap_8 FILLER_66_368 ();
 sg13g2_decap_8 FILLER_66_375 ();
 sg13g2_decap_8 FILLER_66_382 ();
 sg13g2_decap_8 FILLER_66_389 ();
 sg13g2_decap_8 FILLER_66_396 ();
 sg13g2_decap_4 FILLER_66_403 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_fill_2 FILLER_67_21 ();
 sg13g2_decap_4 FILLER_67_49 ();
 sg13g2_fill_1 FILLER_67_72 ();
 sg13g2_fill_2 FILLER_67_90 ();
 sg13g2_fill_2 FILLER_67_160 ();
 sg13g2_fill_2 FILLER_67_258 ();
 sg13g2_fill_2 FILLER_67_269 ();
 sg13g2_fill_1 FILLER_67_271 ();
 sg13g2_fill_2 FILLER_67_307 ();
 sg13g2_fill_1 FILLER_67_314 ();
 sg13g2_decap_8 FILLER_67_356 ();
 sg13g2_decap_8 FILLER_67_363 ();
 sg13g2_decap_8 FILLER_67_370 ();
 sg13g2_decap_8 FILLER_67_377 ();
 sg13g2_decap_8 FILLER_67_384 ();
 sg13g2_decap_8 FILLER_67_391 ();
 sg13g2_decap_8 FILLER_67_398 ();
 sg13g2_decap_4 FILLER_67_405 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_4 FILLER_68_14 ();
 sg13g2_fill_2 FILLER_68_18 ();
 sg13g2_decap_4 FILLER_68_34 ();
 sg13g2_decap_8 FILLER_68_52 ();
 sg13g2_decap_4 FILLER_68_59 ();
 sg13g2_fill_2 FILLER_68_63 ();
 sg13g2_decap_4 FILLER_68_87 ();
 sg13g2_fill_2 FILLER_68_91 ();
 sg13g2_fill_2 FILLER_68_101 ();
 sg13g2_fill_1 FILLER_68_112 ();
 sg13g2_fill_1 FILLER_68_130 ();
 sg13g2_decap_8 FILLER_68_186 ();
 sg13g2_fill_1 FILLER_68_254 ();
 sg13g2_decap_8 FILLER_68_332 ();
 sg13g2_fill_2 FILLER_68_339 ();
 sg13g2_decap_8 FILLER_68_350 ();
 sg13g2_decap_8 FILLER_68_357 ();
 sg13g2_decap_8 FILLER_68_364 ();
 sg13g2_decap_8 FILLER_68_371 ();
 sg13g2_decap_8 FILLER_68_378 ();
 sg13g2_decap_8 FILLER_68_385 ();
 sg13g2_decap_8 FILLER_68_392 ();
 sg13g2_decap_8 FILLER_68_399 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_fill_1 FILLER_69_21 ();
 sg13g2_fill_1 FILLER_69_44 ();
 sg13g2_decap_4 FILLER_69_96 ();
 sg13g2_fill_2 FILLER_69_100 ();
 sg13g2_decap_8 FILLER_69_111 ();
 sg13g2_fill_2 FILLER_69_126 ();
 sg13g2_fill_1 FILLER_69_128 ();
 sg13g2_fill_1 FILLER_69_171 ();
 sg13g2_fill_1 FILLER_69_214 ();
 sg13g2_fill_1 FILLER_69_220 ();
 sg13g2_decap_4 FILLER_69_258 ();
 sg13g2_decap_4 FILLER_69_270 ();
 sg13g2_decap_8 FILLER_69_292 ();
 sg13g2_decap_4 FILLER_69_299 ();
 sg13g2_fill_2 FILLER_69_316 ();
 sg13g2_decap_8 FILLER_69_356 ();
 sg13g2_decap_8 FILLER_69_363 ();
 sg13g2_decap_8 FILLER_69_370 ();
 sg13g2_decap_8 FILLER_69_377 ();
 sg13g2_decap_8 FILLER_69_384 ();
 sg13g2_decap_8 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_69_398 ();
 sg13g2_decap_4 FILLER_69_405 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_14 ();
 sg13g2_fill_2 FILLER_70_49 ();
 sg13g2_decap_4 FILLER_70_86 ();
 sg13g2_fill_1 FILLER_70_90 ();
 sg13g2_decap_4 FILLER_70_104 ();
 sg13g2_fill_1 FILLER_70_108 ();
 sg13g2_decap_4 FILLER_70_114 ();
 sg13g2_fill_1 FILLER_70_123 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_4 FILLER_70_144 ();
 sg13g2_decap_8 FILLER_70_162 ();
 sg13g2_fill_1 FILLER_70_174 ();
 sg13g2_decap_8 FILLER_70_189 ();
 sg13g2_decap_8 FILLER_70_201 ();
 sg13g2_fill_1 FILLER_70_208 ();
 sg13g2_decap_4 FILLER_70_214 ();
 sg13g2_fill_1 FILLER_70_218 ();
 sg13g2_decap_8 FILLER_70_238 ();
 sg13g2_decap_8 FILLER_70_245 ();
 sg13g2_fill_2 FILLER_70_252 ();
 sg13g2_fill_1 FILLER_70_254 ();
 sg13g2_decap_8 FILLER_70_286 ();
 sg13g2_decap_8 FILLER_70_293 ();
 sg13g2_fill_1 FILLER_70_300 ();
 sg13g2_decap_8 FILLER_70_353 ();
 sg13g2_decap_8 FILLER_70_360 ();
 sg13g2_decap_8 FILLER_70_367 ();
 sg13g2_decap_8 FILLER_70_374 ();
 sg13g2_decap_8 FILLER_70_381 ();
 sg13g2_decap_8 FILLER_70_388 ();
 sg13g2_decap_8 FILLER_70_395 ();
 sg13g2_decap_8 FILLER_70_402 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_fill_1 FILLER_71_21 ();
 sg13g2_fill_1 FILLER_71_74 ();
 sg13g2_fill_2 FILLER_71_128 ();
 sg13g2_fill_1 FILLER_71_130 ();
 sg13g2_decap_8 FILLER_71_175 ();
 sg13g2_decap_8 FILLER_71_182 ();
 sg13g2_fill_1 FILLER_71_189 ();
 sg13g2_fill_1 FILLER_71_241 ();
 sg13g2_fill_1 FILLER_71_250 ();
 sg13g2_fill_1 FILLER_71_257 ();
 sg13g2_fill_1 FILLER_71_276 ();
 sg13g2_fill_1 FILLER_71_337 ();
 sg13g2_decap_8 FILLER_71_356 ();
 sg13g2_decap_8 FILLER_71_363 ();
 sg13g2_decap_8 FILLER_71_370 ();
 sg13g2_decap_8 FILLER_71_377 ();
 sg13g2_decap_8 FILLER_71_384 ();
 sg13g2_decap_8 FILLER_71_391 ();
 sg13g2_decap_8 FILLER_71_398 ();
 sg13g2_decap_4 FILLER_71_405 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_fill_2 FILLER_72_69 ();
 sg13g2_fill_1 FILLER_72_71 ();
 sg13g2_fill_2 FILLER_72_118 ();
 sg13g2_fill_1 FILLER_72_120 ();
 sg13g2_fill_1 FILLER_72_130 ();
 sg13g2_fill_1 FILLER_72_189 ();
 sg13g2_fill_2 FILLER_72_198 ();
 sg13g2_decap_8 FILLER_72_208 ();
 sg13g2_decap_4 FILLER_72_215 ();
 sg13g2_fill_2 FILLER_72_219 ();
 sg13g2_decap_8 FILLER_72_309 ();
 sg13g2_fill_2 FILLER_72_316 ();
 sg13g2_decap_8 FILLER_72_335 ();
 sg13g2_decap_8 FILLER_72_342 ();
 sg13g2_decap_8 FILLER_72_349 ();
 sg13g2_decap_8 FILLER_72_356 ();
 sg13g2_decap_8 FILLER_72_363 ();
 sg13g2_decap_8 FILLER_72_370 ();
 sg13g2_decap_8 FILLER_72_377 ();
 sg13g2_decap_8 FILLER_72_384 ();
 sg13g2_decap_8 FILLER_72_391 ();
 sg13g2_decap_8 FILLER_72_398 ();
 sg13g2_decap_4 FILLER_72_405 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_fill_2 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_52 ();
 sg13g2_decap_8 FILLER_73_59 ();
 sg13g2_decap_8 FILLER_73_66 ();
 sg13g2_decap_8 FILLER_73_73 ();
 sg13g2_decap_4 FILLER_73_80 ();
 sg13g2_fill_2 FILLER_73_110 ();
 sg13g2_fill_2 FILLER_73_156 ();
 sg13g2_fill_1 FILLER_73_158 ();
 sg13g2_fill_2 FILLER_73_195 ();
 sg13g2_fill_1 FILLER_73_197 ();
 sg13g2_decap_8 FILLER_73_229 ();
 sg13g2_decap_4 FILLER_73_236 ();
 sg13g2_fill_2 FILLER_73_240 ();
 sg13g2_fill_2 FILLER_73_262 ();
 sg13g2_fill_1 FILLER_73_281 ();
 sg13g2_decap_8 FILLER_73_304 ();
 sg13g2_decap_4 FILLER_73_311 ();
 sg13g2_fill_1 FILLER_73_315 ();
 sg13g2_decap_8 FILLER_73_334 ();
 sg13g2_decap_8 FILLER_73_341 ();
 sg13g2_decap_8 FILLER_73_348 ();
 sg13g2_decap_8 FILLER_73_355 ();
 sg13g2_decap_8 FILLER_73_362 ();
 sg13g2_decap_8 FILLER_73_369 ();
 sg13g2_decap_8 FILLER_73_376 ();
 sg13g2_decap_8 FILLER_73_383 ();
 sg13g2_decap_8 FILLER_73_390 ();
 sg13g2_decap_8 FILLER_73_397 ();
 sg13g2_decap_4 FILLER_73_404 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_4 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_65 ();
 sg13g2_decap_8 FILLER_74_107 ();
 sg13g2_fill_1 FILLER_74_171 ();
 sg13g2_fill_1 FILLER_74_215 ();
 sg13g2_fill_1 FILLER_74_225 ();
 sg13g2_decap_8 FILLER_74_249 ();
 sg13g2_fill_2 FILLER_74_256 ();
 sg13g2_fill_1 FILLER_74_258 ();
 sg13g2_fill_2 FILLER_74_262 ();
 sg13g2_fill_1 FILLER_74_278 ();
 sg13g2_decap_4 FILLER_74_296 ();
 sg13g2_fill_2 FILLER_74_300 ();
 sg13g2_decap_8 FILLER_74_347 ();
 sg13g2_decap_8 FILLER_74_354 ();
 sg13g2_decap_8 FILLER_74_361 ();
 sg13g2_decap_8 FILLER_74_368 ();
 sg13g2_decap_8 FILLER_74_375 ();
 sg13g2_decap_8 FILLER_74_382 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_4 FILLER_75_35 ();
 sg13g2_fill_2 FILLER_75_39 ();
 sg13g2_decap_8 FILLER_75_107 ();
 sg13g2_decap_8 FILLER_75_114 ();
 sg13g2_decap_8 FILLER_75_121 ();
 sg13g2_decap_8 FILLER_75_128 ();
 sg13g2_fill_1 FILLER_75_212 ();
 sg13g2_fill_1 FILLER_75_261 ();
 sg13g2_decap_8 FILLER_75_325 ();
 sg13g2_decap_8 FILLER_75_332 ();
 sg13g2_decap_8 FILLER_75_339 ();
 sg13g2_decap_8 FILLER_75_346 ();
 sg13g2_decap_8 FILLER_75_353 ();
 sg13g2_decap_8 FILLER_75_360 ();
 sg13g2_decap_8 FILLER_75_367 ();
 sg13g2_decap_8 FILLER_75_374 ();
 sg13g2_decap_8 FILLER_75_381 ();
 sg13g2_decap_8 FILLER_75_388 ();
 sg13g2_decap_8 FILLER_75_395 ();
 sg13g2_decap_8 FILLER_75_402 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_4 FILLER_76_35 ();
 sg13g2_fill_2 FILLER_76_39 ();
 sg13g2_decap_4 FILLER_76_69 ();
 sg13g2_fill_2 FILLER_76_73 ();
 sg13g2_decap_8 FILLER_76_132 ();
 sg13g2_fill_2 FILLER_76_139 ();
 sg13g2_fill_1 FILLER_76_141 ();
 sg13g2_decap_4 FILLER_76_152 ();
 sg13g2_decap_4 FILLER_76_173 ();
 sg13g2_fill_1 FILLER_76_177 ();
 sg13g2_fill_2 FILLER_76_266 ();
 sg13g2_fill_1 FILLER_76_268 ();
 sg13g2_decap_4 FILLER_76_298 ();
 sg13g2_fill_1 FILLER_76_302 ();
 sg13g2_decap_8 FILLER_76_312 ();
 sg13g2_decap_8 FILLER_76_319 ();
 sg13g2_decap_8 FILLER_76_326 ();
 sg13g2_decap_8 FILLER_76_333 ();
 sg13g2_decap_8 FILLER_76_340 ();
 sg13g2_decap_8 FILLER_76_347 ();
 sg13g2_decap_8 FILLER_76_354 ();
 sg13g2_decap_8 FILLER_76_361 ();
 sg13g2_decap_8 FILLER_76_368 ();
 sg13g2_decap_8 FILLER_76_375 ();
 sg13g2_decap_8 FILLER_76_382 ();
 sg13g2_decap_8 FILLER_76_389 ();
 sg13g2_decap_8 FILLER_76_396 ();
 sg13g2_decap_4 FILLER_76_403 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_4 FILLER_77_49 ();
 sg13g2_fill_2 FILLER_77_53 ();
 sg13g2_decap_4 FILLER_77_145 ();
 sg13g2_fill_2 FILLER_77_149 ();
 sg13g2_fill_2 FILLER_77_186 ();
 sg13g2_fill_1 FILLER_77_193 ();
 sg13g2_fill_2 FILLER_77_225 ();
 sg13g2_fill_1 FILLER_77_227 ();
 sg13g2_fill_2 FILLER_77_289 ();
 sg13g2_fill_1 FILLER_77_291 ();
 sg13g2_decap_8 FILLER_77_306 ();
 sg13g2_decap_8 FILLER_77_313 ();
 sg13g2_decap_8 FILLER_77_320 ();
 sg13g2_decap_8 FILLER_77_327 ();
 sg13g2_decap_8 FILLER_77_334 ();
 sg13g2_decap_8 FILLER_77_341 ();
 sg13g2_decap_8 FILLER_77_348 ();
 sg13g2_decap_8 FILLER_77_355 ();
 sg13g2_decap_8 FILLER_77_362 ();
 sg13g2_decap_8 FILLER_77_369 ();
 sg13g2_decap_8 FILLER_77_376 ();
 sg13g2_decap_8 FILLER_77_383 ();
 sg13g2_decap_8 FILLER_77_390 ();
 sg13g2_decap_8 FILLER_77_397 ();
 sg13g2_decap_4 FILLER_77_404 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_fill_2 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_79 ();
 sg13g2_fill_2 FILLER_78_115 ();
 sg13g2_decap_4 FILLER_78_148 ();
 sg13g2_fill_2 FILLER_78_152 ();
 sg13g2_decap_8 FILLER_78_180 ();
 sg13g2_decap_8 FILLER_78_187 ();
 sg13g2_decap_4 FILLER_78_194 ();
 sg13g2_fill_1 FILLER_78_198 ();
 sg13g2_decap_4 FILLER_78_225 ();
 sg13g2_fill_2 FILLER_78_264 ();
 sg13g2_decap_8 FILLER_78_306 ();
 sg13g2_decap_8 FILLER_78_313 ();
 sg13g2_decap_8 FILLER_78_320 ();
 sg13g2_decap_8 FILLER_78_327 ();
 sg13g2_decap_8 FILLER_78_334 ();
 sg13g2_decap_8 FILLER_78_341 ();
 sg13g2_decap_8 FILLER_78_348 ();
 sg13g2_decap_8 FILLER_78_355 ();
 sg13g2_decap_8 FILLER_78_362 ();
 sg13g2_decap_8 FILLER_78_369 ();
 sg13g2_decap_8 FILLER_78_376 ();
 sg13g2_decap_8 FILLER_78_383 ();
 sg13g2_decap_8 FILLER_78_390 ();
 sg13g2_decap_8 FILLER_78_397 ();
 sg13g2_decap_4 FILLER_78_404 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_fill_2 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_102 ();
 sg13g2_decap_8 FILLER_79_109 ();
 sg13g2_fill_1 FILLER_79_116 ();
 sg13g2_decap_8 FILLER_79_158 ();
 sg13g2_decap_8 FILLER_79_165 ();
 sg13g2_decap_4 FILLER_79_172 ();
 sg13g2_fill_2 FILLER_79_176 ();
 sg13g2_decap_8 FILLER_79_208 ();
 sg13g2_fill_2 FILLER_79_215 ();
 sg13g2_decap_4 FILLER_79_257 ();
 sg13g2_fill_1 FILLER_79_261 ();
 sg13g2_fill_1 FILLER_79_275 ();
 sg13g2_decap_8 FILLER_79_302 ();
 sg13g2_decap_8 FILLER_79_309 ();
 sg13g2_decap_8 FILLER_79_316 ();
 sg13g2_decap_8 FILLER_79_323 ();
 sg13g2_decap_8 FILLER_79_330 ();
 sg13g2_decap_8 FILLER_79_337 ();
 sg13g2_decap_8 FILLER_79_344 ();
 sg13g2_decap_8 FILLER_79_351 ();
 sg13g2_decap_8 FILLER_79_358 ();
 sg13g2_decap_8 FILLER_79_365 ();
 sg13g2_decap_8 FILLER_79_372 ();
 sg13g2_decap_8 FILLER_79_379 ();
 sg13g2_decap_8 FILLER_79_386 ();
 sg13g2_decap_8 FILLER_79_393 ();
 sg13g2_decap_8 FILLER_79_400 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_fill_2 FILLER_80_136 ();
 sg13g2_fill_1 FILLER_80_138 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_fill_2 FILLER_80_222 ();
 sg13g2_fill_1 FILLER_80_224 ();
 sg13g2_decap_8 FILLER_80_235 ();
 sg13g2_decap_8 FILLER_80_242 ();
 sg13g2_decap_8 FILLER_80_249 ();
 sg13g2_decap_8 FILLER_80_256 ();
 sg13g2_decap_8 FILLER_80_263 ();
 sg13g2_decap_8 FILLER_80_270 ();
 sg13g2_decap_8 FILLER_80_277 ();
 sg13g2_decap_8 FILLER_80_284 ();
 sg13g2_decap_8 FILLER_80_291 ();
 sg13g2_decap_8 FILLER_80_298 ();
 sg13g2_decap_8 FILLER_80_305 ();
 sg13g2_decap_8 FILLER_80_320 ();
 sg13g2_decap_8 FILLER_80_327 ();
 sg13g2_decap_8 FILLER_80_334 ();
 sg13g2_decap_8 FILLER_80_341 ();
 sg13g2_decap_8 FILLER_80_348 ();
 sg13g2_decap_4 FILLER_80_355 ();
 sg13g2_fill_1 FILLER_80_359 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_379 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_fill_2 FILLER_80_407 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
endmodule
