module tt_um_dpi_adexp (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire clknet_leaf_0_clk;
 wire \core.V[0] ;
 wire \core.V[10] ;
 wire \core.V[11] ;
 wire \core.V[12] ;
 wire \core.V[13] ;
 wire \core.V[14] ;
 wire \core.V[15] ;
 wire \core.V[1] ;
 wire \core.V[2] ;
 wire \core.V[3] ;
 wire \core.V[4] ;
 wire \core.V[5] ;
 wire \core.V[6] ;
 wire \core.V[7] ;
 wire \core.V[8] ;
 wire \core.V[9] ;
 wire \core.V_threshold[10] ;
 wire \core.V_threshold[11] ;
 wire \core.V_threshold[12] ;
 wire \core.V_threshold[13] ;
 wire \core.V_threshold[14] ;
 wire \core.V_threshold[15] ;
 wire \core.V_threshold[8] ;
 wire \core.V_threshold[9] ;
 wire \core.byte_acc[0] ;
 wire \core.byte_acc[1] ;
 wire \core.byte_acc[2] ;
 wire \core.byte_acc[3] ;
 wire \core.byte_acc[4] ;
 wire \core.byte_acc[5] ;
 wire \core.byte_acc[6] ;
 wire \core.byte_acc[7] ;
 wire \core.capacitance[10] ;
 wire \core.capacitance[11] ;
 wire \core.capacitance[12] ;
 wire \core.capacitance[13] ;
 wire \core.capacitance[14] ;
 wire \core.capacitance[15] ;
 wire \core.capacitance[8] ;
 wire \core.capacitance[9] ;
 wire \core.compute_state[0] ;
 wire \core.compute_state[1] ;
 wire \core.compute_state[2] ;
 wire \core.compute_state[3] ;
 wire \core.compute_state[4] ;
 wire \core.compute_state[5] ;
 wire \core.compute_state[6] ;
 wire \core.dV[0] ;
 wire \core.dV[10] ;
 wire \core.dV[11] ;
 wire \core.dV[12] ;
 wire \core.dV[13] ;
 wire \core.dV[14] ;
 wire \core.dV[15] ;
 wire \core.dV[1] ;
 wire \core.dV[2] ;
 wire \core.dV[3] ;
 wire \core.dV[4] ;
 wire \core.dV[5] ;
 wire \core.dV[6] ;
 wire \core.dV[7] ;
 wire \core.dV[8] ;
 wire \core.dV[9] ;
 wire \core.delta_t[10] ;
 wire \core.delta_t[11] ;
 wire \core.delta_t[12] ;
 wire \core.delta_t[13] ;
 wire \core.delta_t[14] ;
 wire \core.delta_t[15] ;
 wire \core.delta_t[8] ;
 wire \core.delta_t[9] ;
 wire \core.drive_current[10] ;
 wire \core.drive_current[11] ;
 wire \core.drive_current[12] ;
 wire \core.drive_current[13] ;
 wire \core.drive_current[14] ;
 wire \core.drive_current[15] ;
 wire \core.drive_current[3] ;
 wire \core.drive_current[4] ;
 wire \core.drive_current[5] ;
 wire \core.drive_current[6] ;
 wire \core.drive_current[7] ;
 wire \core.drive_current[8] ;
 wire \core.drive_current[9] ;
 wire \core.dw[0] ;
 wire \core.dw[10] ;
 wire \core.dw[11] ;
 wire \core.dw[12] ;
 wire \core.dw[13] ;
 wire \core.dw[14] ;
 wire \core.dw[15] ;
 wire \core.dw[1] ;
 wire \core.dw[2] ;
 wire \core.dw[3] ;
 wire \core.dw[4] ;
 wire \core.dw[5] ;
 wire \core.dw[6] ;
 wire \core.dw[7] ;
 wire \core.dw[8] ;
 wire \core.dw[9] ;
 wire \core.exp_term[10] ;
 wire \core.exp_term[11] ;
 wire \core.exp_term[12] ;
 wire \core.exp_term[13] ;
 wire \core.exp_term[14] ;
 wire \core.exp_term[15] ;
 wire \core.exp_term[1] ;
 wire \core.exp_term[2] ;
 wire \core.exp_term[3] ;
 wire \core.exp_term[4] ;
 wire \core.exp_term[5] ;
 wire \core.exp_term[6] ;
 wire \core.exp_term[7] ;
 wire \core.exp_term[8] ;
 wire \core.exp_term[9] ;
 wire \core.ibias[10] ;
 wire \core.ibias[11] ;
 wire \core.ibias[12] ;
 wire \core.ibias[13] ;
 wire \core.ibias[14] ;
 wire \core.ibias[15] ;
 wire \core.ibias[8] ;
 wire \core.ibias[9] ;
 wire \core.leak_current[10] ;
 wire \core.leak_current[11] ;
 wire \core.leak_current[12] ;
 wire \core.leak_current[13] ;
 wire \core.leak_current[14] ;
 wire \core.leak_current[15] ;
 wire \core.leak_current[1] ;
 wire \core.leak_current[2] ;
 wire \core.leak_current[3] ;
 wire \core.leak_current[4] ;
 wire \core.leak_current[5] ;
 wire \core.leak_current[6] ;
 wire \core.leak_current[7] ;
 wire \core.leak_current[8] ;
 wire \core.leak_current[9] ;
 wire \core.load_prev ;
 wire \core.lstate[0] ;
 wire \core.lstate[1] ;
 wire \core.lstate[2] ;
 wire \core.nibble_cnt ;
 wire \core.param_a[10] ;
 wire \core.param_a[11] ;
 wire \core.param_a[12] ;
 wire \core.param_a[13] ;
 wire \core.param_a[14] ;
 wire \core.param_a[15] ;
 wire \core.param_a[8] ;
 wire \core.param_a[9] ;
 wire \core.param_b[10] ;
 wire \core.param_b[11] ;
 wire \core.param_b[12] ;
 wire \core.param_b[13] ;
 wire \core.param_b[14] ;
 wire \core.param_b[15] ;
 wire \core.param_b[8] ;
 wire \core.param_b[9] ;
 wire \core.param_idx[0] ;
 wire \core.param_idx[1] ;
 wire \core.param_idx[2] ;
 wire \core.params[0][0] ;
 wire \core.params[0][1] ;
 wire \core.params[0][2] ;
 wire \core.params[0][3] ;
 wire \core.params[0][4] ;
 wire \core.params[0][5] ;
 wire \core.params[0][6] ;
 wire \core.params[0][7] ;
 wire \core.params[1][0] ;
 wire \core.params[1][1] ;
 wire \core.params[1][2] ;
 wire \core.params[1][3] ;
 wire \core.params[1][4] ;
 wire \core.params[1][5] ;
 wire \core.params[1][6] ;
 wire \core.params[1][7] ;
 wire \core.params[2][0] ;
 wire \core.params[2][1] ;
 wire \core.params[2][2] ;
 wire \core.params[2][3] ;
 wire \core.params[2][4] ;
 wire \core.params[2][5] ;
 wire \core.params[2][6] ;
 wire \core.params[2][7] ;
 wire \core.params[3][0] ;
 wire \core.params[3][1] ;
 wire \core.params[3][2] ;
 wire \core.params[3][3] ;
 wire \core.params[3][4] ;
 wire \core.params[3][5] ;
 wire \core.params[3][6] ;
 wire \core.params[3][7] ;
 wire \core.params[5][0] ;
 wire \core.params[5][1] ;
 wire \core.params[5][2] ;
 wire \core.params[5][3] ;
 wire \core.params[5][4] ;
 wire \core.params[5][5] ;
 wire \core.params[5][6] ;
 wire \core.params[5][7] ;
 wire \core.params[6][0] ;
 wire \core.params[6][1] ;
 wire \core.params[6][2] ;
 wire \core.params[6][3] ;
 wire \core.params[6][4] ;
 wire \core.params[6][5] ;
 wire \core.params[6][6] ;
 wire \core.params[6][7] ;
 wire \core.params[7][0] ;
 wire \core.params[7][1] ;
 wire \core.params[7][2] ;
 wire \core.params[7][3] ;
 wire \core.params[7][4] ;
 wire \core.params[7][5] ;
 wire \core.params[7][6] ;
 wire \core.params[7][7] ;
 wire \core.r_ready ;
 wire \core.spike_reg ;
 wire \core.tau_w[10] ;
 wire \core.tau_w[11] ;
 wire \core.tau_w[12] ;
 wire \core.tau_w[13] ;
 wire \core.tau_w[14] ;
 wire \core.tau_w[15] ;
 wire \core.tau_w[8] ;
 wire \core.tau_w[9] ;
 wire \core.temp_q[0] ;
 wire \core.temp_q[10] ;
 wire \core.temp_q[11] ;
 wire \core.temp_q[12] ;
 wire \core.temp_q[13] ;
 wire \core.temp_q[14] ;
 wire \core.temp_q[15] ;
 wire \core.temp_q[1] ;
 wire \core.temp_q[2] ;
 wire \core.temp_q[3] ;
 wire \core.temp_q[4] ;
 wire \core.temp_q[5] ;
 wire \core.temp_q[6] ;
 wire \core.temp_q[7] ;
 wire \core.temp_q[8] ;
 wire \core.temp_q[9] ;
 wire \core.vm8_reg[2] ;
 wire \core.vm8_reg[3] ;
 wire \core.vm8_reg[4] ;
 wire \core.vm8_reg[5] ;
 wire \core.vm8_reg[6] ;
 wire \core.vm8_reg[7] ;
 wire \core.w8_reg[2] ;
 wire \core.w8_reg[3] ;
 wire \core.w8_reg[4] ;
 wire \core.w8_reg[5] ;
 wire \core.w8_reg[6] ;
 wire \core.w8_reg[7] ;
 wire \core.w[0] ;
 wire \core.w[10] ;
 wire \core.w[11] ;
 wire \core.w[12] ;
 wire \core.w[13] ;
 wire \core.w[14] ;
 wire \core.w[15] ;
 wire \core.w[1] ;
 wire \core.w[2] ;
 wire \core.w[3] ;
 wire \core.w[4] ;
 wire \core.w[5] ;
 wire \core.w[6] ;
 wire \core.w[7] ;
 wire \core.w[8] ;
 wire \core.w[9] ;
 wire \core.watchdog_cnt[0] ;
 wire \core.watchdog_cnt[10] ;
 wire \core.watchdog_cnt[11] ;
 wire \core.watchdog_cnt[1] ;
 wire \core.watchdog_cnt[2] ;
 wire \core.watchdog_cnt[3] ;
 wire \core.watchdog_cnt[4] ;
 wire \core.watchdog_cnt[5] ;
 wire \core.watchdog_cnt[6] ;
 wire \core.watchdog_cnt[7] ;
 wire \core.watchdog_cnt[8] ;
 wire \core.watchdog_cnt[9] ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;

 sg13g2_inv_4 _3373_ (.A(\core.byte_acc[7] ),
    .Y(_2622_));
 sg13g2_inv_2 _3374_ (.Y(_2623_),
    .A(\core.byte_acc[6] ));
 sg13g2_inv_1 _3375_ (.Y(_2624_),
    .A(\core.byte_acc[5] ));
 sg13g2_inv_2 _3376_ (.Y(_2625_),
    .A(net454));
 sg13g2_inv_2 _3377_ (.Y(_2626_),
    .A(\core.byte_acc[2] ));
 sg13g2_inv_2 _3378_ (.Y(_2627_),
    .A(\core.byte_acc[1] ));
 sg13g2_inv_1 _3379_ (.Y(_2628_),
    .A(\core.byte_acc[0] ));
 sg13g2_inv_2 _3380_ (.Y(_2629_),
    .A(net862));
 sg13g2_inv_1 _3381_ (.Y(_2630_),
    .A(net678));
 sg13g2_inv_1 _3382_ (.Y(_2631_),
    .A(net883));
 sg13g2_inv_1 _3383_ (.Y(_2632_),
    .A(\core.V_threshold[15] ));
 sg13g2_inv_4 _3384_ (.A(net691),
    .Y(_2633_));
 sg13g2_inv_1 _3385_ (.Y(_2634_),
    .A(net806));
 sg13g2_inv_1 _3386_ (.Y(_2635_),
    .A(net374));
 sg13g2_inv_1 _3387_ (.Y(_2636_),
    .A(net380));
 sg13g2_inv_1 _3388_ (.Y(_2637_),
    .A(net328));
 sg13g2_inv_1 _3389_ (.Y(_2638_),
    .A(net816));
 sg13g2_inv_1 _3390_ (.Y(_2639_),
    .A(net475));
 sg13g2_inv_1 _3391_ (.Y(_2640_),
    .A(net769));
 sg13g2_inv_1 _3392_ (.Y(_2641_),
    .A(net376));
 sg13g2_inv_1 _3393_ (.Y(_2642_),
    .A(net781));
 sg13g2_inv_1 _3394_ (.Y(_2643_),
    .A(net382));
 sg13g2_inv_1 _3395_ (.Y(_2644_),
    .A(net350));
 sg13g2_inv_1 _3396_ (.Y(_2645_),
    .A(net530));
 sg13g2_inv_1 _3397_ (.Y(_2646_),
    .A(net517));
 sg13g2_inv_1 _3398_ (.Y(_2647_),
    .A(net511));
 sg13g2_inv_1 _3399_ (.Y(_2648_),
    .A(net541));
 sg13g2_inv_1 _3400_ (.Y(_2649_),
    .A(net764));
 sg13g2_inv_1 _3401_ (.Y(_2650_),
    .A(\core.temp_q[15] ));
 sg13g2_inv_1 _3402_ (.Y(_2651_),
    .A(\core.temp_q[9] ));
 sg13g2_inv_1 _3403_ (.Y(_2652_),
    .A(\core.temp_q[8] ));
 sg13g2_inv_1 _3404_ (.Y(_2653_),
    .A(net309));
 sg13g2_inv_1 _3405_ (.Y(_2654_),
    .A(net417));
 sg13g2_inv_1 _3406_ (.Y(_2655_),
    .A(net388));
 sg13g2_inv_1 _3407_ (.Y(_2656_),
    .A(net340));
 sg13g2_inv_1 _3408_ (.Y(_2657_),
    .A(net370));
 sg13g2_inv_1 _3409_ (.Y(_2658_),
    .A(net372));
 sg13g2_inv_1 _3410_ (.Y(_2659_),
    .A(net807));
 sg13g2_inv_1 _3411_ (.Y(_2660_),
    .A(net447));
 sg13g2_inv_1 _3412_ (.Y(_2661_),
    .A(net683));
 sg13g2_inv_2 _3413_ (.Y(_2662_),
    .A(net320));
 sg13g2_inv_1 _3414_ (.Y(_2663_),
    .A(net386));
 sg13g2_inv_2 _3415_ (.Y(_2664_),
    .A(net438));
 sg13g2_inv_2 _3416_ (.Y(_2665_),
    .A(net394));
 sg13g2_inv_1 _3417_ (.Y(_2666_),
    .A(net826));
 sg13g2_inv_1 _3418_ (.Y(_2667_),
    .A(net474));
 sg13g2_inv_1 _3419_ (.Y(_2668_),
    .A(net824));
 sg13g2_inv_1 _3420_ (.Y(_2669_),
    .A(net507));
 sg13g2_inv_1 _3421_ (.Y(_2670_),
    .A(net844));
 sg13g2_inv_1 _3422_ (.Y(_2671_),
    .A(net505));
 sg13g2_inv_1 _3423_ (.Y(_2672_),
    .A(net808));
 sg13g2_inv_1 _3424_ (.Y(_2673_),
    .A(net422));
 sg13g2_inv_1 _3425_ (.Y(_2674_),
    .A(\core.param_a[15] ));
 sg13g2_inv_1 _3426_ (.Y(_2675_),
    .A(net413));
 sg13g2_inv_1 _3427_ (.Y(_2676_),
    .A(net399));
 sg13g2_inv_1 _3428_ (.Y(_2677_),
    .A(net338));
 sg13g2_inv_1 _3429_ (.Y(_2678_),
    .A(net322));
 sg13g2_inv_1 _3430_ (.Y(_2679_),
    .A(net359));
 sg13g2_inv_1 _3431_ (.Y(_2680_),
    .A(net470));
 sg13g2_inv_1 _3432_ (.Y(_2681_),
    .A(net716));
 sg13g2_inv_1 _3433_ (.Y(_2682_),
    .A(net401));
 sg13g2_inv_1 _3434_ (.Y(_2683_),
    .A(net500));
 sg13g2_inv_1 _3435_ (.Y(_2684_),
    .A(net773));
 sg13g2_inv_1 _3436_ (.Y(_2685_),
    .A(net410));
 sg13g2_inv_1 _3437_ (.Y(_2686_),
    .A(net497));
 sg13g2_inv_1 _3438_ (.Y(_2687_),
    .A(net443));
 sg13g2_inv_1 _3439_ (.Y(_2688_),
    .A(net332));
 sg13g2_inv_1 _3440_ (.Y(_2689_),
    .A(net486));
 sg13g2_inv_1 _3441_ (.Y(_2690_),
    .A(net455));
 sg13g2_inv_1 _3442_ (.Y(_2691_),
    .A(net366));
 sg13g2_inv_1 _3443_ (.Y(_2692_),
    .A(net334));
 sg13g2_inv_1 _3444_ (.Y(_2693_),
    .A(net326));
 sg13g2_inv_1 _3445_ (.Y(_2694_),
    .A(net342));
 sg13g2_inv_1 _3446_ (.Y(_2695_),
    .A(net436));
 sg13g2_inv_2 _3447_ (.Y(_2696_),
    .A(net525));
 sg13g2_inv_1 _3448_ (.Y(_2697_),
    .A(net547));
 sg13g2_inv_1 _3449_ (.Y(_2698_),
    .A(net415));
 sg13g2_inv_1 _3450_ (.Y(_2699_),
    .A(net336));
 sg13g2_inv_1 _3451_ (.Y(_2700_),
    .A(net795));
 sg13g2_inv_1 _3452_ (.Y(_2701_),
    .A(net449));
 sg13g2_inv_1 _3453_ (.Y(_2702_),
    .A(net356));
 sg13g2_inv_1 _3454_ (.Y(_2703_),
    .A(net361));
 sg13g2_inv_1 _3455_ (.Y(_2704_),
    .A(net364));
 sg13g2_inv_1 _3456_ (.Y(_2705_),
    .A(\core.tau_w[15] ));
 sg13g2_inv_1 _3457_ (.Y(_2706_),
    .A(net476));
 sg13g2_inv_1 _3458_ (.Y(_2707_),
    .A(net553));
 sg13g2_inv_1 _3459_ (.Y(_2708_),
    .A(net459));
 sg13g2_inv_1 _3460_ (.Y(_2709_),
    .A(net809));
 sg13g2_inv_1 _3461_ (.Y(_2710_),
    .A(net445));
 sg13g2_inv_1 _3462_ (.Y(_2711_),
    .A(net378));
 sg13g2_inv_1 _3463_ (.Y(_2712_),
    .A(net346));
 sg13g2_inv_1 _3464_ (.Y(_2713_),
    .A(net390));
 sg13g2_inv_1 _3465_ (.Y(_2714_),
    .A(net406));
 sg13g2_inv_1 _3466_ (.Y(_2715_),
    .A(net368));
 sg13g2_inv_1 _3467_ (.Y(_2716_),
    .A(net352));
 sg13g2_inv_1 _3468_ (.Y(_2717_),
    .A(net430));
 sg13g2_inv_1 _3469_ (.Y(_2718_),
    .A(net324));
 sg13g2_inv_1 _3470_ (.Y(_2719_),
    .A(\core.lstate[2] ));
 sg13g2_inv_4 _3471_ (.A(net749),
    .Y(_2720_));
 sg13g2_inv_1 _3472_ (.Y(_2721_),
    .A(net739));
 sg13g2_inv_1 _3473_ (.Y(_2722_),
    .A(\core.watchdog_cnt[8] ));
 sg13g2_inv_1 _3474_ (.Y(_2723_),
    .A(\core.watchdog_cnt[5] ));
 sg13g2_inv_1 _3475_ (.Y(_2724_),
    .A(net392));
 sg13g2_inv_1 _3476_ (.Y(_2725_),
    .A(_0008_));
 sg13g2_inv_1 _3477_ (.Y(_2726_),
    .A(_0019_));
 sg13g2_inv_1 _3478_ (.Y(_2727_),
    .A(_0026_));
 sg13g2_inv_1 _3479_ (.Y(_2728_),
    .A(_0025_));
 sg13g2_inv_1 _3480_ (.Y(_2729_),
    .A(_0027_));
 sg13g2_inv_1 _3481_ (.Y(_2730_),
    .A(_0031_));
 sg13g2_inv_1 _3482_ (.Y(_2731_),
    .A(_0032_));
 sg13g2_inv_1 _3483_ (.Y(_2732_),
    .A(_0034_));
 sg13g2_inv_1 _3484_ (.Y(_2733_),
    .A(_0033_));
 sg13g2_inv_1 _3485_ (.Y(_2734_),
    .A(_0035_));
 sg13g2_inv_1 _3486_ (.Y(_2735_),
    .A(net463));
 sg13g2_nand2_2 _3487_ (.Y(_2736_),
    .A(net745),
    .B(net739));
 sg13g2_or3_1 _3488_ (.A(\core.delta_t[10] ),
    .B(\core.delta_t[9] ),
    .C(\core.delta_t[8] ),
    .X(_2737_));
 sg13g2_or2_1 _3489_ (.X(_2738_),
    .B(_2737_),
    .A(\core.delta_t[11] ));
 sg13g2_or2_1 _3490_ (.X(_2739_),
    .B(_2738_),
    .A(\core.delta_t[12] ));
 sg13g2_nor2_1 _3491_ (.A(\core.delta_t[13] ),
    .B(_2739_),
    .Y(_2740_));
 sg13g2_nor4_2 _3492_ (.A(net681),
    .B(\core.delta_t[14] ),
    .C(\core.delta_t[13] ),
    .Y(_2741_),
    .D(_2739_));
 sg13g2_a21oi_1 _3493_ (.A1(\core.compute_state[4] ),
    .A2(_2741_),
    .Y(_2742_),
    .B1(net408));
 sg13g2_nor2_1 _3494_ (.A(_2736_),
    .B(net409),
    .Y(_0006_));
 sg13g2_nor2_2 _3495_ (.A(net850),
    .B(_2736_),
    .Y(_2743_));
 sg13g2_inv_1 _3496_ (.Y(_0005_),
    .A(_2743_));
 sg13g2_nand2_1 _3497_ (.Y(_2744_),
    .A(\core.w8_reg[2] ),
    .B(net741));
 sg13g2_o21ai_1 _3498_ (.B1(_2744_),
    .Y(uo_out[1]),
    .A1(_2648_),
    .A2(net741));
 sg13g2_nand2_1 _3499_ (.Y(_2745_),
    .A(\core.w8_reg[3] ),
    .B(net1));
 sg13g2_o21ai_1 _3500_ (.B1(_2745_),
    .Y(uo_out[2]),
    .A1(_2647_),
    .A2(net741));
 sg13g2_nand2_1 _3501_ (.Y(_2746_),
    .A(\core.w8_reg[4] ),
    .B(net1));
 sg13g2_o21ai_1 _3502_ (.B1(_2746_),
    .Y(uo_out[3]),
    .A1(_2646_),
    .A2(net741));
 sg13g2_nand2_1 _3503_ (.Y(_2747_),
    .A(\core.w8_reg[5] ),
    .B(net1));
 sg13g2_o21ai_1 _3504_ (.B1(_2747_),
    .Y(uo_out[4]),
    .A1(_2645_),
    .A2(net741));
 sg13g2_mux2_2 _3505_ (.A0(\core.vm8_reg[6] ),
    .A1(\core.w8_reg[6] ),
    .S(net741),
    .X(uo_out[5]));
 sg13g2_nor2_1 _3506_ (.A(\core.vm8_reg[7] ),
    .B(net741),
    .Y(_2748_));
 sg13g2_a21oi_2 _3507_ (.B1(_2748_),
    .Y(uo_out[6]),
    .A2(net741),
    .A1(_2649_));
 sg13g2_nand2_1 _3508_ (.Y(_2749_),
    .A(net740),
    .B(net857));
 sg13g2_nor2_1 _3509_ (.A(net724),
    .B(net648),
    .Y(_0004_));
 sg13g2_and2_1 _3510_ (.A(net740),
    .B(\core.compute_state[0] ),
    .X(_2750_));
 sg13g2_and2_1 _3511_ (.A(net744),
    .B(net644),
    .X(_0003_));
 sg13g2_nand2_1 _3512_ (.Y(_2751_),
    .A(net740),
    .B(net852));
 sg13g2_nor2_1 _3513_ (.A(net724),
    .B(net640),
    .Y(_0002_));
 sg13g2_nor2b_1 _3514_ (.A(_2741_),
    .B_N(net861),
    .Y(_2752_));
 sg13g2_nand2_1 _3515_ (.Y(_2753_),
    .A(net739),
    .B(_2752_));
 sg13g2_nor2_1 _3516_ (.A(net723),
    .B(_2753_),
    .Y(_0001_));
 sg13g2_and2_1 _3517_ (.A(net739),
    .B(net893),
    .X(_2754_));
 sg13g2_nand2_2 _3518_ (.Y(_2755_),
    .A(net739),
    .B(net791));
 sg13g2_nor2_1 _3519_ (.A(net721),
    .B(_2755_),
    .Y(_0000_));
 sg13g2_nor3_2 _3520_ (.A(\core.lstate[0] ),
    .B(\core.lstate[1] ),
    .C(_2719_),
    .Y(_2756_));
 sg13g2_o21ai_1 _3521_ (.B1(net753),
    .Y(_2757_),
    .A1(net853),
    .A2(_2756_));
 sg13g2_nand2_1 _3522_ (.Y(_2758_),
    .A(\core.lstate[0] ),
    .B(\core.lstate[1] ));
 sg13g2_nand3_1 _3523_ (.B(\core.lstate[1] ),
    .C(net853),
    .A(\core.lstate[0] ),
    .Y(_2759_));
 sg13g2_nor2b_2 _3524_ (.A(\core.load_prev ),
    .B_N(net2),
    .Y(_2760_));
 sg13g2_nand2b_2 _3525_ (.Y(_2761_),
    .B(net2),
    .A_N(\core.load_prev ));
 sg13g2_nand4_1 _3526_ (.B(net4),
    .C(net7),
    .A(net5),
    .Y(_2762_),
    .D(net6));
 sg13g2_nor3_1 _3527_ (.A(_2759_),
    .B(_2761_),
    .C(_2762_),
    .Y(_2763_));
 sg13g2_nand2_1 _3528_ (.Y(_2764_),
    .A(net3),
    .B(_2756_));
 sg13g2_nand4_1 _3529_ (.B(\core.watchdog_cnt[9] ),
    .C(\core.watchdog_cnt[8] ),
    .A(\core.watchdog_cnt[10] ),
    .Y(_2765_),
    .D(\core.watchdog_cnt[11] ));
 sg13g2_o21ai_1 _3530_ (.B1(\core.watchdog_cnt[7] ),
    .Y(_2766_),
    .A1(\core.watchdog_cnt[6] ),
    .A2(\core.watchdog_cnt[5] ));
 sg13g2_nor2_2 _3531_ (.A(_2765_),
    .B(_2766_),
    .Y(_2767_));
 sg13g2_nor3_1 _3532_ (.A(net853),
    .B(_2764_),
    .C(_2767_),
    .Y(_2768_));
 sg13g2_nor2_1 _3533_ (.A(_2763_),
    .B(net854),
    .Y(_2769_));
 sg13g2_nor2_1 _3534_ (.A(_2757_),
    .B(net855),
    .Y(_0058_));
 sg13g2_nand2_1 _3535_ (.Y(_2770_),
    .A(\core.lstate[1] ),
    .B(_0054_));
 sg13g2_nor2_2 _3536_ (.A(\core.lstate[0] ),
    .B(_2770_),
    .Y(_2771_));
 sg13g2_nand2_1 _3537_ (.Y(_2772_),
    .A(net685),
    .B(net684));
 sg13g2_nand2_1 _3538_ (.Y(_2773_),
    .A(net847),
    .B(net685));
 sg13g2_nand3_1 _3539_ (.B(net685),
    .C(net684),
    .A(\core.param_idx[0] ),
    .Y(_2774_));
 sg13g2_nand4_1 _3540_ (.B(net685),
    .C(net684),
    .A(\core.param_idx[0] ),
    .Y(_2775_),
    .D(_2771_));
 sg13g2_nor2b_2 _3541_ (.A(\core.lstate[1] ),
    .B_N(_0054_),
    .Y(_2776_));
 sg13g2_nor2b_1 _3542_ (.A(\core.lstate[0] ),
    .B_N(_2776_),
    .Y(_2777_));
 sg13g2_nand2b_2 _3543_ (.Y(_2778_),
    .B(_2776_),
    .A_N(\core.lstate[0] ));
 sg13g2_nand2_2 _3544_ (.Y(_2779_),
    .A(_2767_),
    .B(_2778_));
 sg13g2_inv_1 _3545_ (.Y(_2780_),
    .A(_2779_));
 sg13g2_and2_1 _3546_ (.A(\core.lstate[0] ),
    .B(_2776_),
    .X(_2781_));
 sg13g2_nand2_1 _3547_ (.Y(_2782_),
    .A(\core.nibble_cnt ),
    .B(_2760_));
 sg13g2_nand4_1 _3548_ (.B(net3),
    .C(_2760_),
    .A(\core.nibble_cnt ),
    .Y(_2783_),
    .D(net631));
 sg13g2_o21ai_1 _3549_ (.B1(_2783_),
    .Y(_2784_),
    .A1(net766),
    .A2(_2780_));
 sg13g2_nand2_1 _3550_ (.Y(_2785_),
    .A(net3),
    .B(_2760_));
 sg13g2_a22oi_1 _3551_ (.Y(_2786_),
    .B1(_2785_),
    .B2(net633),
    .A2(_2781_),
    .A1(net3));
 sg13g2_inv_1 _3552_ (.Y(_2787_),
    .A(_2786_));
 sg13g2_o21ai_1 _3553_ (.B1(_2764_),
    .Y(_2788_),
    .A1(_2759_),
    .A2(_2760_));
 sg13g2_o21ai_1 _3554_ (.B1(net767),
    .Y(_2789_),
    .A1(_2787_),
    .A2(_2788_));
 sg13g2_a21oi_1 _3555_ (.A1(_2775_),
    .A2(_2789_),
    .Y(_0059_),
    .B1(_2757_));
 sg13g2_nand3_1 _3556_ (.B(net631),
    .C(_2782_),
    .A(net3),
    .Y(_2790_));
 sg13g2_nor2_1 _3557_ (.A(net633),
    .B(_2788_),
    .Y(_2791_));
 sg13g2_or2_2 _3558_ (.X(_2792_),
    .B(_2785_),
    .A(_2778_));
 sg13g2_a22oi_1 _3559_ (.Y(_2793_),
    .B1(_2792_),
    .B2(net784),
    .A2(_2791_),
    .A1(_2790_));
 sg13g2_a21oi_1 _3560_ (.A1(_2779_),
    .A2(_2793_),
    .Y(_2794_),
    .B1(_2771_));
 sg13g2_nor2_1 _3561_ (.A(_2757_),
    .B(net785),
    .Y(_0060_));
 sg13g2_nor2_2 _3562_ (.A(net865),
    .B(_2761_),
    .Y(_2795_));
 sg13g2_nand2_1 _3563_ (.Y(_2796_),
    .A(net631),
    .B(_2795_));
 sg13g2_and2_1 _3564_ (.A(_2792_),
    .B(_2796_),
    .X(_2797_));
 sg13g2_and2_1 _3565_ (.A(net4),
    .B(net631),
    .X(_2798_));
 sg13g2_a22oi_1 _3566_ (.Y(_2799_),
    .B1(_2798_),
    .B2(net866),
    .A2(_2797_),
    .A1(net869));
 sg13g2_nor2_1 _3567_ (.A(net736),
    .B(_2799_),
    .Y(_0061_));
 sg13g2_and2_1 _3568_ (.A(net5),
    .B(net631),
    .X(_2800_));
 sg13g2_a22oi_1 _3569_ (.Y(_2801_),
    .B1(_2800_),
    .B2(net866),
    .A2(_2797_),
    .A1(\core.byte_acc[5] ));
 sg13g2_nor2_1 _3570_ (.A(net735),
    .B(net867),
    .Y(_0062_));
 sg13g2_and2_1 _3571_ (.A(net6),
    .B(net631),
    .X(_2802_));
 sg13g2_a22oi_1 _3572_ (.Y(_2803_),
    .B1(_2802_),
    .B2(_2795_),
    .A2(_2797_),
    .A1(net863));
 sg13g2_nor2_1 _3573_ (.A(net736),
    .B(net864),
    .Y(_0063_));
 sg13g2_and2_1 _3574_ (.A(net7),
    .B(net631),
    .X(_2804_));
 sg13g2_a22oi_1 _3575_ (.Y(_2805_),
    .B1(_2804_),
    .B2(_2795_),
    .A2(_2797_),
    .A1(net827));
 sg13g2_nor2_1 _3576_ (.A(net736),
    .B(net828),
    .Y(_0064_));
 sg13g2_and2_1 _3577_ (.A(net755),
    .B(net2),
    .X(_0065_));
 sg13g2_nand2_1 _3578_ (.Y(_2806_),
    .A(net754),
    .B(_2771_));
 sg13g2_or2_1 _3579_ (.X(_2807_),
    .B(_2806_),
    .A(\core.param_idx[0] ));
 sg13g2_nor3_2 _3580_ (.A(net685),
    .B(net684),
    .C(_2807_),
    .Y(_2808_));
 sg13g2_nor2_2 _3581_ (.A(net731),
    .B(_2808_),
    .Y(_2809_));
 sg13g2_a22oi_1 _3582_ (.Y(_2810_),
    .B1(_2809_),
    .B2(net348),
    .A2(net617),
    .A1(\core.byte_acc[0] ));
 sg13g2_inv_1 _3583_ (.Y(_0066_),
    .A(net349));
 sg13g2_a22oi_1 _3584_ (.Y(_0067_),
    .B1(_2809_),
    .B2(_2660_),
    .A2(net617),
    .A1(_2627_));
 sg13g2_a22oi_1 _3585_ (.Y(_2811_),
    .B1(_2809_),
    .B2(net372),
    .A2(net617),
    .A1(\core.byte_acc[2] ));
 sg13g2_inv_1 _3586_ (.Y(_0068_),
    .A(net373));
 sg13g2_a22oi_1 _3587_ (.Y(_2812_),
    .B1(_2809_),
    .B2(net370),
    .A2(net617),
    .A1(\core.byte_acc[3] ));
 sg13g2_inv_1 _3588_ (.Y(_0069_),
    .A(net371));
 sg13g2_a22oi_1 _3589_ (.Y(_2813_),
    .B1(_2809_),
    .B2(net340),
    .A2(net617),
    .A1(\core.byte_acc[4] ));
 sg13g2_inv_1 _3590_ (.Y(_0070_),
    .A(net341));
 sg13g2_a22oi_1 _3591_ (.Y(_2814_),
    .B1(_2809_),
    .B2(net388),
    .A2(net617),
    .A1(\core.byte_acc[5] ));
 sg13g2_inv_1 _3592_ (.Y(_0071_),
    .A(net389));
 sg13g2_a22oi_1 _3593_ (.Y(_2815_),
    .B1(_2809_),
    .B2(net417),
    .A2(net617),
    .A1(\core.byte_acc[6] ));
 sg13g2_inv_1 _3594_ (.Y(_0072_),
    .A(net418));
 sg13g2_a22oi_1 _3595_ (.Y(_0073_),
    .B1(_2809_),
    .B2(_2717_),
    .A2(net617),
    .A1(_2622_));
 sg13g2_o21ai_1 _3596_ (.B1(net752),
    .Y(_2816_),
    .A1(net699),
    .A2(net363));
 sg13g2_a21oi_1 _3597_ (.A1(net699),
    .A2(_2716_),
    .Y(_0074_),
    .B1(_2816_));
 sg13g2_o21ai_1 _3598_ (.B1(net752),
    .Y(_2817_),
    .A1(net704),
    .A2(net396));
 sg13g2_a21oi_1 _3599_ (.A1(net703),
    .A2(_2715_),
    .Y(_0075_),
    .B1(net397));
 sg13g2_a21oi_1 _3600_ (.A1(net703),
    .A2(\core.params[1][2] ),
    .Y(_2818_),
    .B1(net736));
 sg13g2_o21ai_1 _3601_ (.B1(_2818_),
    .Y(_0076_),
    .A1(net703),
    .A2(_2713_));
 sg13g2_o21ai_1 _3602_ (.B1(net752),
    .Y(_2819_),
    .A1(net703),
    .A2(net451));
 sg13g2_a21oi_1 _3603_ (.A1(net703),
    .A2(_2712_),
    .Y(_0077_),
    .B1(_2819_));
 sg13g2_o21ai_1 _3604_ (.B1(net752),
    .Y(_2820_),
    .A1(net698),
    .A2(net452));
 sg13g2_a21oi_1 _3605_ (.A1(net699),
    .A2(_2711_),
    .Y(_0078_),
    .B1(_2820_));
 sg13g2_a21oi_1 _3606_ (.A1(net704),
    .A2(net445),
    .Y(_2821_),
    .B1(net733));
 sg13g2_o21ai_1 _3607_ (.B1(_2821_),
    .Y(_0079_),
    .A1(net699),
    .A2(_2709_));
 sg13g2_a21oi_1 _3608_ (.A1(net703),
    .A2(net459),
    .Y(_2822_),
    .B1(net733));
 sg13g2_o21ai_1 _3609_ (.B1(_2822_),
    .Y(_0080_),
    .A1(net698),
    .A2(_2707_));
 sg13g2_o21ai_1 _3610_ (.B1(net751),
    .Y(_2823_),
    .A1(net698),
    .A2(net518));
 sg13g2_a21oi_1 _3611_ (.A1(net698),
    .A2(_2706_),
    .Y(_0081_),
    .B1(_2823_));
 sg13g2_o21ai_1 _3612_ (.B1(net754),
    .Y(_2824_),
    .A1(net701),
    .A2(net426));
 sg13g2_a21oi_1 _3613_ (.A1(net701),
    .A2(_2704_),
    .Y(_0082_),
    .B1(_2824_));
 sg13g2_o21ai_1 _3614_ (.B1(net754),
    .Y(_2825_),
    .A1(net702),
    .A2(net433));
 sg13g2_a21oi_1 _3615_ (.A1(net702),
    .A2(_2703_),
    .Y(_0083_),
    .B1(_2825_));
 sg13g2_o21ai_1 _3616_ (.B1(net754),
    .Y(_2826_),
    .A1(net702),
    .A2(net442));
 sg13g2_a21oi_1 _3617_ (.A1(net702),
    .A2(_2702_),
    .Y(_0084_),
    .B1(_2826_));
 sg13g2_a21oi_1 _3618_ (.A1(net702),
    .A2(net449),
    .Y(_2827_),
    .B1(net735));
 sg13g2_o21ai_1 _3619_ (.B1(_2827_),
    .Y(_0085_),
    .A1(net702),
    .A2(_2700_));
 sg13g2_o21ai_1 _3620_ (.B1(net754),
    .Y(_2828_),
    .A1(net701),
    .A2(net465));
 sg13g2_a21oi_1 _3621_ (.A1(net701),
    .A2(_2699_),
    .Y(_0086_),
    .B1(_2828_));
 sg13g2_a21oi_1 _3622_ (.A1(net701),
    .A2(net415),
    .Y(_2829_),
    .B1(net735));
 sg13g2_o21ai_1 _3623_ (.B1(_2829_),
    .Y(_0087_),
    .A1(net701),
    .A2(_2697_));
 sg13g2_o21ai_1 _3624_ (.B1(net754),
    .Y(_2830_),
    .A1(_2633_),
    .A2(net354));
 sg13g2_a21oi_1 _3625_ (.A1(_2633_),
    .A2(_2696_),
    .Y(_0088_),
    .B1(_2830_));
 sg13g2_o21ai_1 _3626_ (.B1(net754),
    .Y(_2831_),
    .A1(net701),
    .A2(net466));
 sg13g2_a21oi_1 _3627_ (.A1(net701),
    .A2(_2695_),
    .Y(_0089_),
    .B1(_2831_));
 sg13g2_o21ai_1 _3628_ (.B1(net750),
    .Y(_2832_),
    .A1(net694),
    .A2(net358));
 sg13g2_a21oi_1 _3629_ (.A1(net694),
    .A2(_2694_),
    .Y(_0090_),
    .B1(_2832_));
 sg13g2_o21ai_1 _3630_ (.B1(net750),
    .Y(_2833_),
    .A1(net694),
    .A2(net420));
 sg13g2_a21oi_1 _3631_ (.A1(net694),
    .A2(_2693_),
    .Y(_0091_),
    .B1(_2833_));
 sg13g2_o21ai_1 _3632_ (.B1(net750),
    .Y(_2834_),
    .A1(net693),
    .A2(net434));
 sg13g2_a21oi_1 _3633_ (.A1(net693),
    .A2(_2692_),
    .Y(_0092_),
    .B1(_2834_));
 sg13g2_a21oi_1 _3634_ (.A1(net694),
    .A2(net366),
    .Y(_2835_),
    .B1(net731));
 sg13g2_o21ai_1 _3635_ (.B1(_2835_),
    .Y(_0093_),
    .A1(net694),
    .A2(_2690_));
 sg13g2_o21ai_1 _3636_ (.B1(net756),
    .Y(_2836_),
    .A1(_2633_),
    .A2(net344));
 sg13g2_a21oi_1 _3637_ (.A1(_2633_),
    .A2(_2689_),
    .Y(_0094_),
    .B1(_2836_));
 sg13g2_o21ai_1 _3638_ (.B1(net750),
    .Y(_2837_),
    .A1(net694),
    .A2(net428));
 sg13g2_a21oi_1 _3639_ (.A1(net695),
    .A2(_2688_),
    .Y(_0095_),
    .B1(_2837_));
 sg13g2_a21oi_1 _3640_ (.A1(net693),
    .A2(net443),
    .Y(_2838_),
    .B1(net732));
 sg13g2_o21ai_1 _3641_ (.B1(_2838_),
    .Y(_0096_),
    .A1(net693),
    .A2(_2686_));
 sg13g2_a21oi_1 _3642_ (.A1(net694),
    .A2(net410),
    .Y(_2839_),
    .B1(net731));
 sg13g2_o21ai_1 _3643_ (.B1(_2839_),
    .Y(_0097_),
    .A1(net693),
    .A2(_2684_));
 sg13g2_o21ai_1 _3644_ (.B1(net748),
    .Y(_2840_),
    .A1(net697),
    .A2(net718));
 sg13g2_a21oi_1 _3645_ (.A1(net697),
    .A2(_2683_),
    .Y(_0098_),
    .B1(_2840_));
 sg13g2_a21oi_1 _3646_ (.A1(net700),
    .A2(net401),
    .Y(_2841_),
    .B1(net733));
 sg13g2_o21ai_1 _3647_ (.B1(_2841_),
    .Y(_0099_),
    .A1(net697),
    .A2(_2681_));
 sg13g2_o21ai_1 _3648_ (.B1(net751),
    .Y(_2842_),
    .A1(net697),
    .A2(net713));
 sg13g2_a21oi_1 _3649_ (.A1(net697),
    .A2(_2680_),
    .Y(_0100_),
    .B1(_2842_));
 sg13g2_o21ai_1 _3650_ (.B1(net752),
    .Y(_2843_),
    .A1(net698),
    .A2(net711));
 sg13g2_a21oi_1 _3651_ (.A1(net698),
    .A2(_2679_),
    .Y(_0101_),
    .B1(_2843_));
 sg13g2_o21ai_1 _3652_ (.B1(net752),
    .Y(_2844_),
    .A1(net698),
    .A2(net709));
 sg13g2_a21oi_1 _3653_ (.A1(net698),
    .A2(_2678_),
    .Y(_0102_),
    .B1(_2844_));
 sg13g2_o21ai_1 _3654_ (.B1(net751),
    .Y(_2845_),
    .A1(net700),
    .A2(net707));
 sg13g2_a21oi_1 _3655_ (.A1(net697),
    .A2(_2677_),
    .Y(_0103_),
    .B1(net425));
 sg13g2_o21ai_1 _3656_ (.B1(net751),
    .Y(_2846_),
    .A1(net697),
    .A2(net432));
 sg13g2_a21oi_1 _3657_ (.A1(net697),
    .A2(_2676_),
    .Y(_0104_),
    .B1(_2846_));
 sg13g2_o21ai_1 _3658_ (.B1(net752),
    .Y(_2847_),
    .A1(net703),
    .A2(\core.param_a[15] ));
 sg13g2_a21oi_1 _3659_ (.A1(net703),
    .A2(_2675_),
    .Y(_0105_),
    .B1(_2847_));
 sg13g2_or2_1 _3660_ (.X(_2848_),
    .B(_2806_),
    .A(net313));
 sg13g2_nor2_1 _3661_ (.A(_2772_),
    .B(_2848_),
    .Y(_2849_));
 sg13g2_nor2_2 _3662_ (.A(net732),
    .B(_2849_),
    .Y(_2850_));
 sg13g2_a22oi_1 _3663_ (.Y(_2851_),
    .B1(_2850_),
    .B2(net342),
    .A2(net616),
    .A1(\core.byte_acc[0] ));
 sg13g2_inv_1 _3664_ (.Y(_0106_),
    .A(net343));
 sg13g2_a22oi_1 _3665_ (.Y(_2852_),
    .B1(_2850_),
    .B2(net326),
    .A2(net616),
    .A1(\core.byte_acc[1] ));
 sg13g2_inv_1 _3666_ (.Y(_0107_),
    .A(net327));
 sg13g2_a22oi_1 _3667_ (.Y(_2853_),
    .B1(_2850_),
    .B2(net334),
    .A2(net616),
    .A1(\core.byte_acc[2] ));
 sg13g2_inv_1 _3668_ (.Y(_0108_),
    .A(net335));
 sg13g2_a22oi_1 _3669_ (.Y(_0109_),
    .B1(_2850_),
    .B2(_2691_),
    .A2(net616),
    .A1(_2625_));
 sg13g2_a22oi_1 _3670_ (.Y(_2854_),
    .B1(_2850_),
    .B2(net344),
    .A2(net616),
    .A1(\core.byte_acc[4] ));
 sg13g2_inv_1 _3671_ (.Y(_0110_),
    .A(net345));
 sg13g2_a22oi_1 _3672_ (.Y(_2855_),
    .B1(_2850_),
    .B2(net332),
    .A2(net616),
    .A1(\core.byte_acc[5] ));
 sg13g2_inv_1 _3673_ (.Y(_0111_),
    .A(net333));
 sg13g2_a22oi_1 _3674_ (.Y(_0112_),
    .B1(_2850_),
    .B2(_2687_),
    .A2(net616),
    .A1(_2623_));
 sg13g2_a22oi_1 _3675_ (.Y(_0113_),
    .B1(_2850_),
    .B2(_2685_),
    .A2(net616),
    .A1(_2622_));
 sg13g2_nor2_1 _3676_ (.A(_2772_),
    .B(_2807_),
    .Y(_0335_));
 sg13g2_nor2_2 _3677_ (.A(net731),
    .B(net615),
    .Y(_0336_));
 sg13g2_a22oi_1 _3678_ (.Y(_0114_),
    .B1(_0336_),
    .B2(_2673_),
    .A2(_0335_),
    .A1(_2628_));
 sg13g2_a22oi_1 _3679_ (.Y(_0115_),
    .B1(_0336_),
    .B2(_2671_),
    .A2(net615),
    .A1(_2627_));
 sg13g2_a22oi_1 _3680_ (.Y(_0116_),
    .B1(_0336_),
    .B2(_2669_),
    .A2(net615),
    .A1(_2626_));
 sg13g2_a22oi_1 _3681_ (.Y(_0117_),
    .B1(_0336_),
    .B2(_2667_),
    .A2(net615),
    .A1(_2625_));
 sg13g2_a22oi_1 _3682_ (.Y(_0337_),
    .B1(_0336_),
    .B2(net394),
    .A2(net615),
    .A1(\core.byte_acc[4] ));
 sg13g2_inv_1 _3683_ (.Y(_0118_),
    .A(net395));
 sg13g2_a22oi_1 _3684_ (.Y(_0338_),
    .B1(_0336_),
    .B2(net438),
    .A2(net615),
    .A1(\core.byte_acc[5] ));
 sg13g2_inv_1 _3685_ (.Y(_0119_),
    .A(net439));
 sg13g2_a22oi_1 _3686_ (.Y(_0339_),
    .B1(_0336_),
    .B2(net386),
    .A2(net615),
    .A1(\core.byte_acc[6] ));
 sg13g2_inv_1 _3687_ (.Y(_0120_),
    .A(net387));
 sg13g2_a22oi_1 _3688_ (.Y(_0121_),
    .B1(_0336_),
    .B2(_2718_),
    .A2(net615),
    .A1(_2622_));
 sg13g2_o21ai_1 _3689_ (.B1(_2764_),
    .Y(_0340_),
    .A1(_2756_),
    .A2(_2763_));
 sg13g2_o21ai_1 _3690_ (.B1(net753),
    .Y(_0341_),
    .A1(net876),
    .A2(_0340_));
 sg13g2_a21oi_1 _3691_ (.A1(_2633_),
    .A2(_0340_),
    .Y(_0122_),
    .B1(_0341_));
 sg13g2_nor2_1 _3692_ (.A(_2767_),
    .B(net632),
    .Y(_0342_));
 sg13g2_a21oi_1 _3693_ (.A1(net633),
    .A2(_2785_),
    .Y(_0343_),
    .B1(_2761_));
 sg13g2_nand2_1 _3694_ (.Y(_0344_),
    .A(_2776_),
    .B(_0343_));
 sg13g2_nand2_1 _3695_ (.Y(_0345_),
    .A(net755),
    .B(_0344_));
 sg13g2_nand2_1 _3696_ (.Y(_0346_),
    .A(net860),
    .B(_2778_));
 sg13g2_o21ai_1 _3697_ (.B1(_0346_),
    .Y(_0347_),
    .A1(net860),
    .A2(net622));
 sg13g2_nor2_1 _3698_ (.A(net614),
    .B(_0347_),
    .Y(_0123_));
 sg13g2_nand2_1 _3699_ (.Y(_0348_),
    .A(\core.watchdog_cnt[0] ),
    .B(net812));
 sg13g2_a22oi_1 _3700_ (.Y(_0349_),
    .B1(net622),
    .B2(_0348_),
    .A2(net632),
    .A1(net812));
 sg13g2_nor2_1 _3701_ (.A(\core.watchdog_cnt[0] ),
    .B(net812),
    .Y(_0350_));
 sg13g2_nor3_1 _3702_ (.A(net614),
    .B(_0349_),
    .C(net813),
    .Y(_0124_));
 sg13g2_xor2_1 _3703_ (.B(_0348_),
    .A(_0046_),
    .X(_0351_));
 sg13g2_a22oi_1 _3704_ (.Y(_0352_),
    .B1(net622),
    .B2(_0351_),
    .A2(net632),
    .A1(net536));
 sg13g2_nor2_1 _3705_ (.A(net614),
    .B(net537),
    .Y(_0125_));
 sg13g2_nand3_1 _3706_ (.B(_2779_),
    .C(_0344_),
    .A(net753),
    .Y(_0353_));
 sg13g2_nand4_1 _3707_ (.B(\core.watchdog_cnt[1] ),
    .C(net536),
    .A(\core.watchdog_cnt[0] ),
    .Y(_0354_),
    .D(_2778_));
 sg13g2_nand4_1 _3708_ (.B(net892),
    .C(net536),
    .A(\core.watchdog_cnt[0] ),
    .Y(_0355_),
    .D(net761));
 sg13g2_xor2_1 _3709_ (.B(_0354_),
    .A(net761),
    .X(_0356_));
 sg13g2_nor2_1 _3710_ (.A(_0353_),
    .B(net762),
    .Y(_0126_));
 sg13g2_xor2_1 _3711_ (.B(_0355_),
    .A(_0047_),
    .X(_0357_));
 sg13g2_a22oi_1 _3712_ (.Y(_0358_),
    .B1(net622),
    .B2(_0357_),
    .A2(net632),
    .A1(net463));
 sg13g2_nor2_1 _3713_ (.A(net614),
    .B(net464),
    .Y(_0127_));
 sg13g2_nor3_1 _3714_ (.A(_2735_),
    .B(net632),
    .C(_0355_),
    .Y(_0359_));
 sg13g2_nor3_2 _3715_ (.A(_2723_),
    .B(_2735_),
    .C(_0355_),
    .Y(_0360_));
 sg13g2_xnor2_1 _3716_ (.Y(_0361_),
    .A(net788),
    .B(_0359_));
 sg13g2_nor2_1 _3717_ (.A(_0353_),
    .B(_0361_),
    .Y(_0128_));
 sg13g2_xnor2_1 _3718_ (.Y(_0362_),
    .A(net550),
    .B(_0360_));
 sg13g2_a22oi_1 _3719_ (.Y(_0363_),
    .B1(net622),
    .B2(_0362_),
    .A2(net632),
    .A1(\core.watchdog_cnt[6] ));
 sg13g2_nor2_1 _3720_ (.A(net614),
    .B(net551),
    .Y(_0129_));
 sg13g2_nand3_1 _3721_ (.B(\core.watchdog_cnt[6] ),
    .C(_0360_),
    .A(net480),
    .Y(_0364_));
 sg13g2_a22oi_1 _3722_ (.Y(_0365_),
    .B1(net622),
    .B2(_0364_),
    .A2(net632),
    .A1(net480));
 sg13g2_a21oi_1 _3723_ (.A1(\core.watchdog_cnt[6] ),
    .A2(_0360_),
    .Y(_0366_),
    .B1(net480));
 sg13g2_nor3_1 _3724_ (.A(net614),
    .B(_0365_),
    .C(net481),
    .Y(_0130_));
 sg13g2_xor2_1 _3725_ (.B(_0364_),
    .A(net489),
    .X(_0367_));
 sg13g2_a22oi_1 _3726_ (.Y(_0368_),
    .B1(_0342_),
    .B2(net490),
    .A2(net633),
    .A1(\core.watchdog_cnt[8] ));
 sg13g2_nor2_1 _3727_ (.A(_0345_),
    .B(net491),
    .Y(_0131_));
 sg13g2_nor2_1 _3728_ (.A(_2722_),
    .B(_0364_),
    .Y(_0369_));
 sg13g2_nand2_1 _3729_ (.Y(_0370_),
    .A(net799),
    .B(_0369_));
 sg13g2_a22oi_1 _3730_ (.Y(_0371_),
    .B1(net622),
    .B2(_0370_),
    .A2(net633),
    .A1(net799));
 sg13g2_nor2_1 _3731_ (.A(net799),
    .B(_0369_),
    .Y(_0372_));
 sg13g2_nor3_1 _3732_ (.A(net614),
    .B(_0371_),
    .C(net800),
    .Y(_0132_));
 sg13g2_xor2_1 _3733_ (.B(_0370_),
    .A(_0050_),
    .X(_0373_));
 sg13g2_a22oi_1 _3734_ (.Y(_0374_),
    .B1(net622),
    .B2(_0373_),
    .A2(net632),
    .A1(net483));
 sg13g2_nor2_1 _3735_ (.A(net614),
    .B(net484),
    .Y(_0133_));
 sg13g2_nand4_1 _3736_ (.B(\core.watchdog_cnt[9] ),
    .C(_2778_),
    .A(\core.watchdog_cnt[10] ),
    .Y(_0375_),
    .D(_0369_));
 sg13g2_a21oi_1 _3737_ (.A1(_2724_),
    .A2(_0375_),
    .Y(_0134_),
    .B1(_0353_));
 sg13g2_nand4_1 _3738_ (.B(_2758_),
    .C(_2775_),
    .A(_0054_),
    .Y(_0376_),
    .D(_2786_));
 sg13g2_and2_1 _3739_ (.A(_2779_),
    .B(_0376_),
    .X(_0377_));
 sg13g2_and2_1 _3740_ (.A(_2771_),
    .B(_2774_),
    .X(_0378_));
 sg13g2_a22oi_1 _3741_ (.Y(_0379_),
    .B1(_0378_),
    .B2(net313),
    .A2(_0377_),
    .A1(\core.param_idx[0] ));
 sg13g2_nor2_1 _3742_ (.A(net735),
    .B(net314),
    .Y(_0135_));
 sg13g2_a22oi_1 _3743_ (.Y(_0380_),
    .B1(_0377_),
    .B2(net685),
    .A2(_2773_),
    .A1(_2771_));
 sg13g2_o21ai_1 _3744_ (.B1(net754),
    .Y(_0381_),
    .A1(net847),
    .A2(net685));
 sg13g2_nor2_1 _3745_ (.A(_0380_),
    .B(_0381_),
    .Y(_0136_));
 sg13g2_nand2b_1 _3746_ (.Y(_0382_),
    .B(_2773_),
    .A_N(net684));
 sg13g2_nand2_1 _3747_ (.Y(_0383_),
    .A(_2776_),
    .B(_2786_));
 sg13g2_a22oi_1 _3748_ (.Y(_0384_),
    .B1(_0378_),
    .B2(_0382_),
    .A2(_2779_),
    .A1(net684));
 sg13g2_nand2_1 _3749_ (.Y(_0385_),
    .A(net753),
    .B(_0383_));
 sg13g2_nor2_1 _3750_ (.A(_0384_),
    .B(_0385_),
    .Y(_0137_));
 sg13g2_nand4_1 _3751_ (.B(net317),
    .C(_2760_),
    .A(net3),
    .Y(_0386_),
    .D(net631));
 sg13g2_nand4_1 _3752_ (.B(_2779_),
    .C(_0344_),
    .A(\core.nibble_cnt ),
    .Y(_0387_),
    .D(_0383_));
 sg13g2_a21oi_1 _3753_ (.A1(net318),
    .A2(_0387_),
    .Y(_0138_),
    .B1(net735));
 sg13g2_nand3_1 _3754_ (.B(_2760_),
    .C(_2781_),
    .A(\core.nibble_cnt ),
    .Y(_0388_));
 sg13g2_nand2_1 _3755_ (.Y(_0389_),
    .A(_2792_),
    .B(_0388_));
 sg13g2_a21oi_1 _3756_ (.A1(_2792_),
    .A2(_0388_),
    .Y(_0390_),
    .B1(_2798_));
 sg13g2_o21ai_1 _3757_ (.B1(net753),
    .Y(_0391_),
    .A1(\core.byte_acc[0] ),
    .A2(_0389_));
 sg13g2_nor2_1 _3758_ (.A(_0390_),
    .B(_0391_),
    .Y(_0139_));
 sg13g2_a21oi_1 _3759_ (.A1(_2792_),
    .A2(_0388_),
    .Y(_0392_),
    .B1(_2800_));
 sg13g2_o21ai_1 _3760_ (.B1(net753),
    .Y(_0393_),
    .A1(net874),
    .A2(_0389_));
 sg13g2_nor2_1 _3761_ (.A(_0392_),
    .B(_0393_),
    .Y(_0140_));
 sg13g2_a21oi_1 _3762_ (.A1(_2792_),
    .A2(_0388_),
    .Y(_0394_),
    .B1(_2802_));
 sg13g2_o21ai_1 _3763_ (.B1(net753),
    .Y(_0395_),
    .A1(net798),
    .A2(_0389_));
 sg13g2_nor2_1 _3764_ (.A(_0394_),
    .B(_0395_),
    .Y(_0141_));
 sg13g2_a21oi_1 _3765_ (.A1(_2792_),
    .A2(_0388_),
    .Y(_0396_),
    .B1(_2804_));
 sg13g2_o21ai_1 _3766_ (.B1(net753),
    .Y(_0397_),
    .A1(net454),
    .A2(_0389_));
 sg13g2_nor2_1 _3767_ (.A(_0396_),
    .B(_0397_),
    .Y(_0142_));
 sg13g2_o21ai_1 _3768_ (.B1(net747),
    .Y(_0398_),
    .A1(net829),
    .A2(net643));
 sg13g2_a21oi_1 _3769_ (.A1(_2630_),
    .A2(net643),
    .Y(_0143_),
    .B1(_0398_));
 sg13g2_xnor2_1 _3770_ (.Y(_0399_),
    .A(net676),
    .B(net677));
 sg13g2_inv_1 _3771_ (.Y(_0400_),
    .A(_0399_));
 sg13g2_o21ai_1 _3772_ (.B1(net746),
    .Y(_0401_),
    .A1(net842),
    .A2(net642));
 sg13g2_a21oi_1 _3773_ (.A1(net642),
    .A2(_0399_),
    .Y(_0144_),
    .B1(_0401_));
 sg13g2_nor3_2 _3774_ (.A(net673),
    .B(net676),
    .C(net677),
    .Y(_0402_));
 sg13g2_o21ai_1 _3775_ (.B1(net673),
    .Y(_0403_),
    .A1(net676),
    .A2(net677));
 sg13g2_nor2b_2 _3776_ (.A(_0402_),
    .B_N(_0403_),
    .Y(_0404_));
 sg13g2_nand2_1 _3777_ (.Y(_0405_),
    .A(net677),
    .B(_0404_));
 sg13g2_xnor2_1 _3778_ (.Y(_0406_),
    .A(net677),
    .B(_0404_));
 sg13g2_o21ai_1 _3779_ (.B1(net746),
    .Y(_0407_),
    .A1(net819),
    .A2(net642));
 sg13g2_a21oi_1 _3780_ (.A1(net642),
    .A2(_0406_),
    .Y(_0145_),
    .B1(_0407_));
 sg13g2_nor2_2 _3781_ (.A(net671),
    .B(_0399_),
    .Y(_0408_));
 sg13g2_nor2b_1 _3782_ (.A(net671),
    .B_N(_0402_),
    .Y(_0409_));
 sg13g2_xnor2_1 _3783_ (.Y(_0410_),
    .A(net671),
    .B(_0402_));
 sg13g2_nor2_1 _3784_ (.A(_0400_),
    .B(_0410_),
    .Y(_0411_));
 sg13g2_nor3_2 _3785_ (.A(_0405_),
    .B(_0408_),
    .C(_0411_),
    .Y(_0412_));
 sg13g2_o21ai_1 _3786_ (.B1(_0405_),
    .Y(_0413_),
    .A1(_0408_),
    .A2(_0411_));
 sg13g2_nand2b_1 _3787_ (.Y(_0414_),
    .B(_0413_),
    .A_N(_0412_));
 sg13g2_o21ai_1 _3788_ (.B1(net746),
    .Y(_0415_),
    .A1(net831),
    .A2(net643));
 sg13g2_a21oi_1 _3789_ (.A1(net643),
    .A2(_0414_),
    .Y(_0146_),
    .B1(_0415_));
 sg13g2_nand2b_1 _3790_ (.Y(_0416_),
    .B(_0404_),
    .A_N(net668));
 sg13g2_nor2b_1 _3791_ (.A(net668),
    .B_N(_0409_),
    .Y(_0417_));
 sg13g2_xnor2_1 _3792_ (.Y(_0418_),
    .A(net668),
    .B(_0409_));
 sg13g2_mux2_1 _3793_ (.A0(_0418_),
    .A1(net668),
    .S(_0404_),
    .X(_0419_));
 sg13g2_and2_1 _3794_ (.A(_0408_),
    .B(_0419_),
    .X(_0420_));
 sg13g2_xor2_1 _3795_ (.B(_0419_),
    .A(_0408_),
    .X(_0421_));
 sg13g2_and2_1 _3796_ (.A(_0412_),
    .B(_0421_),
    .X(_0422_));
 sg13g2_xnor2_1 _3797_ (.Y(_0423_),
    .A(_0412_),
    .B(_0421_));
 sg13g2_o21ai_1 _3798_ (.B1(net746),
    .Y(_0424_),
    .A1(net839),
    .A2(net643));
 sg13g2_a21oi_1 _3799_ (.A1(net642),
    .A2(_0423_),
    .Y(_0147_),
    .B1(_0424_));
 sg13g2_nor2b_1 _3800_ (.A(net666),
    .B_N(_0410_),
    .Y(_0425_));
 sg13g2_nor2b_1 _3801_ (.A(net666),
    .B_N(_0417_),
    .Y(_0426_));
 sg13g2_xnor2_1 _3802_ (.Y(_0427_),
    .A(net666),
    .B(_0417_));
 sg13g2_nor2_1 _3803_ (.A(_0410_),
    .B(_0427_),
    .Y(_0428_));
 sg13g2_nor2_1 _3804_ (.A(_0425_),
    .B(_0428_),
    .Y(_0429_));
 sg13g2_nand2b_1 _3805_ (.Y(_0430_),
    .B(_0429_),
    .A_N(_0416_));
 sg13g2_xnor2_1 _3806_ (.Y(_0431_),
    .A(_0416_),
    .B(_0429_));
 sg13g2_o21ai_1 _3807_ (.B1(_0431_),
    .Y(_0432_),
    .A1(_0420_),
    .A2(_0422_));
 sg13g2_or3_1 _3808_ (.A(_0420_),
    .B(_0422_),
    .C(_0431_),
    .X(_0433_));
 sg13g2_nand2_1 _3809_ (.Y(_0434_),
    .A(_0432_),
    .B(_0433_));
 sg13g2_o21ai_1 _3810_ (.B1(net746),
    .Y(_0435_),
    .A1(net815),
    .A2(net642));
 sg13g2_a21oi_1 _3811_ (.A1(net642),
    .A2(_0434_),
    .Y(_0148_),
    .B1(_0435_));
 sg13g2_nor2b_1 _3812_ (.A(net664),
    .B_N(_0418_),
    .Y(_0436_));
 sg13g2_nor2b_1 _3813_ (.A(net664),
    .B_N(_0426_),
    .Y(_0437_));
 sg13g2_xnor2_1 _3814_ (.Y(_0438_),
    .A(net664),
    .B(_0426_));
 sg13g2_nor2_1 _3815_ (.A(_0418_),
    .B(_0438_),
    .Y(_0439_));
 sg13g2_nor2_1 _3816_ (.A(_0436_),
    .B(_0439_),
    .Y(_0440_));
 sg13g2_nand2_1 _3817_ (.Y(_0441_),
    .A(_0425_),
    .B(_0440_));
 sg13g2_xnor2_1 _3818_ (.Y(_0442_),
    .A(_0425_),
    .B(_0440_));
 sg13g2_a21o_1 _3819_ (.A2(_0432_),
    .A1(_0430_),
    .B1(_0442_),
    .X(_0443_));
 sg13g2_nand3_1 _3820_ (.B(_0432_),
    .C(_0442_),
    .A(_0430_),
    .Y(_0444_));
 sg13g2_nand2_1 _3821_ (.Y(_0445_),
    .A(_0443_),
    .B(_0444_));
 sg13g2_o21ai_1 _3822_ (.B1(net742),
    .Y(_0446_),
    .A1(net835),
    .A2(net641));
 sg13g2_a21oi_1 _3823_ (.A1(net642),
    .A2(_0445_),
    .Y(_0149_),
    .B1(_0446_));
 sg13g2_nor2b_1 _3824_ (.A(net662),
    .B_N(_0427_),
    .Y(_0447_));
 sg13g2_nand2b_1 _3825_ (.Y(_0448_),
    .B(_0437_),
    .A_N(net662));
 sg13g2_xnor2_1 _3826_ (.Y(_0449_),
    .A(net662),
    .B(_0437_));
 sg13g2_inv_1 _3827_ (.Y(_0450_),
    .A(_0449_));
 sg13g2_nor2_1 _3828_ (.A(_0427_),
    .B(_0449_),
    .Y(_0451_));
 sg13g2_nor2_1 _3829_ (.A(_0447_),
    .B(_0451_),
    .Y(_0452_));
 sg13g2_nand2_1 _3830_ (.Y(_0453_),
    .A(_0436_),
    .B(_0452_));
 sg13g2_xnor2_1 _3831_ (.Y(_0454_),
    .A(_0436_),
    .B(_0452_));
 sg13g2_a21o_1 _3832_ (.A2(_0443_),
    .A1(_0441_),
    .B1(_0454_),
    .X(_0455_));
 sg13g2_nand3_1 _3833_ (.B(_0443_),
    .C(_0454_),
    .A(_0441_),
    .Y(_0456_));
 sg13g2_nand2_1 _3834_ (.Y(_0457_),
    .A(_0455_),
    .B(_0456_));
 sg13g2_o21ai_1 _3835_ (.B1(net742),
    .Y(_0458_),
    .A1(net821),
    .A2(net641));
 sg13g2_a21oi_1 _3836_ (.A1(net641),
    .A2(_0457_),
    .Y(_0150_),
    .B1(_0458_));
 sg13g2_nor2b_1 _3837_ (.A(net661),
    .B_N(_0438_),
    .Y(_0459_));
 sg13g2_nor2_2 _3838_ (.A(net661),
    .B(_0448_),
    .Y(_0460_));
 sg13g2_xor2_1 _3839_ (.B(_0448_),
    .A(net661),
    .X(_0461_));
 sg13g2_nor2_1 _3840_ (.A(_0438_),
    .B(_0461_),
    .Y(_0462_));
 sg13g2_nor2_1 _3841_ (.A(_0459_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_xnor2_1 _3842_ (.Y(_0464_),
    .A(_0447_),
    .B(_0463_));
 sg13g2_a21oi_1 _3843_ (.A1(_0453_),
    .A2(_0455_),
    .Y(_0465_),
    .B1(_0464_));
 sg13g2_nand3_1 _3844_ (.B(_0455_),
    .C(_0464_),
    .A(_0453_),
    .Y(_0466_));
 sg13g2_nand2b_1 _3845_ (.Y(_0467_),
    .B(_0466_),
    .A_N(_0465_));
 sg13g2_o21ai_1 _3846_ (.B1(net742),
    .Y(_0468_),
    .A1(net820),
    .A2(net641));
 sg13g2_a21oi_1 _3847_ (.A1(net641),
    .A2(_0467_),
    .Y(_0151_),
    .B1(_0468_));
 sg13g2_nor2_1 _3848_ (.A(_0052_),
    .B(_0450_),
    .Y(_0469_));
 sg13g2_xnor2_1 _3849_ (.Y(_0470_),
    .A(_0052_),
    .B(_0460_));
 sg13g2_nor2_1 _3850_ (.A(_0449_),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_nor2_1 _3851_ (.A(_0469_),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_nor2_1 _3852_ (.A(_0459_),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_a21oi_1 _3853_ (.A1(_0447_),
    .A2(_0463_),
    .Y(_0474_),
    .B1(_0465_));
 sg13g2_nand2_1 _3854_ (.Y(_0475_),
    .A(_0459_),
    .B(_0472_));
 sg13g2_and2_1 _3855_ (.A(_0474_),
    .B(_0475_),
    .X(_0476_));
 sg13g2_nand2b_1 _3856_ (.Y(_0477_),
    .B(_0475_),
    .A_N(_0473_));
 sg13g2_xnor2_1 _3857_ (.Y(_0478_),
    .A(_0474_),
    .B(_0477_));
 sg13g2_o21ai_1 _3858_ (.B1(net742),
    .Y(_0479_),
    .A1(net834),
    .A2(net641));
 sg13g2_a21oi_1 _3859_ (.A1(net641),
    .A2(_0478_),
    .Y(_0152_),
    .B1(_0479_));
 sg13g2_nor2b_1 _3860_ (.A(_0460_),
    .B_N(net657),
    .Y(_0480_));
 sg13g2_xnor2_1 _3861_ (.Y(_0481_),
    .A(_0053_),
    .B(_0480_));
 sg13g2_nand2_1 _3862_ (.Y(_0482_),
    .A(_0461_),
    .B(_0481_));
 sg13g2_xnor2_1 _3863_ (.Y(_0483_),
    .A(_0461_),
    .B(_0481_));
 sg13g2_nor3_1 _3864_ (.A(_0052_),
    .B(_0450_),
    .C(_0483_),
    .Y(_0484_));
 sg13g2_xor2_1 _3865_ (.B(_0483_),
    .A(_0469_),
    .X(_0485_));
 sg13g2_nor3_1 _3866_ (.A(_0473_),
    .B(_0476_),
    .C(_0485_),
    .Y(_0486_));
 sg13g2_o21ai_1 _3867_ (.B1(_0485_),
    .Y(_0487_),
    .A1(_0473_),
    .A2(_0476_));
 sg13g2_nand2b_1 _3868_ (.Y(_0488_),
    .B(_0487_),
    .A_N(_0486_));
 sg13g2_o21ai_1 _3869_ (.B1(net742),
    .Y(_0489_),
    .A1(net830),
    .A2(net645));
 sg13g2_a21oi_1 _3870_ (.A1(net641),
    .A2(_0488_),
    .Y(_0153_),
    .B1(_0489_));
 sg13g2_nor2_1 _3871_ (.A(net656),
    .B(_0480_),
    .Y(_0490_));
 sg13g2_xor2_1 _3872_ (.B(_0490_),
    .A(net655),
    .X(_0491_));
 sg13g2_nand2_1 _3873_ (.Y(_0492_),
    .A(_0470_),
    .B(_0491_));
 sg13g2_xnor2_1 _3874_ (.Y(_0493_),
    .A(_0470_),
    .B(_0491_));
 sg13g2_xor2_1 _3875_ (.B(_0493_),
    .A(_0482_),
    .X(_0494_));
 sg13g2_o21ai_1 _3876_ (.B1(_0494_),
    .Y(_0495_),
    .A1(_0484_),
    .A2(_0486_));
 sg13g2_or3_1 _3877_ (.A(_0484_),
    .B(_0486_),
    .C(_0494_),
    .X(_0496_));
 sg13g2_nand2_1 _3878_ (.Y(_0497_),
    .A(_0495_),
    .B(_0496_));
 sg13g2_o21ai_1 _3879_ (.B1(net743),
    .Y(_0498_),
    .A1(net825),
    .A2(net644));
 sg13g2_a21oi_1 _3880_ (.A1(net644),
    .A2(_0497_),
    .Y(_0154_),
    .B1(_0498_));
 sg13g2_o21ai_1 _3881_ (.B1(_0495_),
    .Y(_0499_),
    .A1(_0482_),
    .A2(_0493_));
 sg13g2_a21oi_1 _3882_ (.A1(net657),
    .A2(_0460_),
    .Y(_0500_),
    .B1(_0052_));
 sg13g2_o21ai_1 _3883_ (.B1(net655),
    .Y(_0501_),
    .A1(net656),
    .A2(_0500_));
 sg13g2_inv_1 _3884_ (.Y(_0502_),
    .A(_0501_));
 sg13g2_xor2_1 _3885_ (.B(_0501_),
    .A(net654),
    .X(_0503_));
 sg13g2_and2_1 _3886_ (.A(_0481_),
    .B(_0503_),
    .X(_0504_));
 sg13g2_xor2_1 _3887_ (.B(_0503_),
    .A(_0481_),
    .X(_0505_));
 sg13g2_nand2b_1 _3888_ (.Y(_0506_),
    .B(_0505_),
    .A_N(_0492_));
 sg13g2_xnor2_1 _3889_ (.Y(_0507_),
    .A(_0492_),
    .B(_0505_));
 sg13g2_nand2_1 _3890_ (.Y(_0508_),
    .A(_0499_),
    .B(_0507_));
 sg13g2_xnor2_1 _3891_ (.Y(_0509_),
    .A(_0499_),
    .B(_0507_));
 sg13g2_o21ai_1 _3892_ (.B1(net744),
    .Y(_0510_),
    .A1(net840),
    .A2(net645));
 sg13g2_a21oi_1 _3893_ (.A1(net644),
    .A2(_0509_),
    .Y(_0155_),
    .B1(net841));
 sg13g2_nor2_1 _3894_ (.A(_0021_),
    .B(_0501_),
    .Y(_0511_));
 sg13g2_xnor2_1 _3895_ (.Y(_0512_),
    .A(net653),
    .B(_0511_));
 sg13g2_nand2_1 _3896_ (.Y(_0513_),
    .A(_0491_),
    .B(_0512_));
 sg13g2_xor2_1 _3897_ (.B(_0512_),
    .A(_0491_),
    .X(_0514_));
 sg13g2_xnor2_1 _3898_ (.Y(_0515_),
    .A(_0504_),
    .B(_0514_));
 sg13g2_a21oi_1 _3899_ (.A1(_0506_),
    .A2(_0508_),
    .Y(_0516_),
    .B1(_0515_));
 sg13g2_nand3_1 _3900_ (.B(_0508_),
    .C(_0515_),
    .A(_0506_),
    .Y(_0517_));
 sg13g2_nand2b_1 _3901_ (.Y(_0518_),
    .B(_0517_),
    .A_N(_0516_));
 sg13g2_o21ai_1 _3902_ (.B1(net745),
    .Y(_0519_),
    .A1(net843),
    .A2(net644));
 sg13g2_a21oi_1 _3903_ (.A1(net644),
    .A2(_0518_),
    .Y(_0156_),
    .B1(_0519_));
 sg13g2_o21ai_1 _3904_ (.B1(net744),
    .Y(_0520_),
    .A1(net823),
    .A2(net644));
 sg13g2_a21oi_1 _3905_ (.A1(_0504_),
    .A2(_0514_),
    .Y(_0521_),
    .B1(_0516_));
 sg13g2_o21ai_1 _3906_ (.B1(net653),
    .Y(_0522_),
    .A1(net654),
    .A2(_0502_));
 sg13g2_nand2_1 _3907_ (.Y(_0523_),
    .A(_0503_),
    .B(_0522_));
 sg13g2_xnor2_1 _3908_ (.Y(_0524_),
    .A(_2629_),
    .B(_0523_));
 sg13g2_xnor2_1 _3909_ (.Y(_0525_),
    .A(_0513_),
    .B(_0524_));
 sg13g2_xnor2_1 _3910_ (.Y(_0526_),
    .A(_0521_),
    .B(_0525_));
 sg13g2_a21oi_1 _3911_ (.A1(net644),
    .A2(_0526_),
    .Y(_0157_),
    .B1(_0520_));
 sg13g2_a21oi_1 _3912_ (.A1(net690),
    .A2(net422),
    .Y(_0527_),
    .B1(net731));
 sg13g2_o21ai_1 _3913_ (.B1(_0527_),
    .Y(_0158_),
    .A1(net691),
    .A2(_2672_));
 sg13g2_a21oi_2 _3914_ (.B1(net731),
    .Y(_0528_),
    .A2(net505),
    .A1(net691));
 sg13g2_o21ai_1 _3915_ (.B1(_0528_),
    .Y(_0159_),
    .A1(net686),
    .A2(_2670_));
 sg13g2_a21oi_2 _3916_ (.B1(net728),
    .Y(_0529_),
    .A2(net507),
    .A1(net687));
 sg13g2_o21ai_1 _3917_ (.B1(_0529_),
    .Y(_0160_),
    .A1(net686),
    .A2(_2668_));
 sg13g2_a21oi_2 _3918_ (.B1(net731),
    .Y(_0530_),
    .A2(net474),
    .A1(net691));
 sg13g2_o21ai_1 _3919_ (.B1(_0530_),
    .Y(_0161_),
    .A1(net687),
    .A2(_2666_));
 sg13g2_o21ai_1 _3920_ (.B1(net744),
    .Y(_0531_),
    .A1(net686),
    .A2(net529));
 sg13g2_a21oi_1 _3921_ (.A1(net686),
    .A2(_2665_),
    .Y(_0162_),
    .B1(_0531_));
 sg13g2_o21ai_1 _3922_ (.B1(net744),
    .Y(_0532_),
    .A1(net686),
    .A2(net494));
 sg13g2_a21oi_1 _3923_ (.A1(net686),
    .A2(_2664_),
    .Y(_0163_),
    .B1(_0532_));
 sg13g2_o21ai_1 _3924_ (.B1(net749),
    .Y(_0533_),
    .A1(net690),
    .A2(net412));
 sg13g2_a21oi_1 _3925_ (.A1(net690),
    .A2(_2663_),
    .Y(_0164_),
    .B1(_0533_));
 sg13g2_o21ai_1 _3926_ (.B1(net744),
    .Y(_0534_),
    .A1(net686),
    .A2(\core.ibias[15] ));
 sg13g2_a21oi_1 _3927_ (.A1(net686),
    .A2(_2662_),
    .Y(_0165_),
    .B1(_0534_));
 sg13g2_o21ai_1 _3928_ (.B1(net749),
    .Y(_0535_),
    .A1(_2633_),
    .A2(net348));
 sg13g2_a21oi_1 _3929_ (.A1(_2633_),
    .A2(_2661_),
    .Y(_0166_),
    .B1(_0535_));
 sg13g2_a21oi_1 _3930_ (.A1(net689),
    .A2(net447),
    .Y(_0536_),
    .B1(net731));
 sg13g2_o21ai_1 _3931_ (.B1(_0536_),
    .Y(_0167_),
    .A1(net689),
    .A2(_2659_));
 sg13g2_o21ai_1 _3932_ (.B1(net749),
    .Y(_0537_),
    .A1(net689),
    .A2(net435));
 sg13g2_a21oi_1 _3933_ (.A1(net689),
    .A2(_2658_),
    .Y(_0168_),
    .B1(_0537_));
 sg13g2_o21ai_1 _3934_ (.B1(net749),
    .Y(_0538_),
    .A1(net688),
    .A2(net403));
 sg13g2_a21oi_1 _3935_ (.A1(net688),
    .A2(_2657_),
    .Y(_0169_),
    .B1(_0538_));
 sg13g2_o21ai_1 _3936_ (.B1(net749),
    .Y(_0539_),
    .A1(net688),
    .A2(net498));
 sg13g2_a21oi_1 _3937_ (.A1(net689),
    .A2(_2656_),
    .Y(_0170_),
    .B1(_0539_));
 sg13g2_o21ai_1 _3938_ (.B1(net749),
    .Y(_0540_),
    .A1(net688),
    .A2(net453));
 sg13g2_a21oi_1 _3939_ (.A1(net688),
    .A2(_2655_),
    .Y(_0171_),
    .B1(_0540_));
 sg13g2_o21ai_1 _3940_ (.B1(net749),
    .Y(_0541_),
    .A1(net688),
    .A2(net457));
 sg13g2_a21oi_1 _3941_ (.A1(net688),
    .A2(_2654_),
    .Y(_0172_),
    .B1(_0541_));
 sg13g2_o21ai_1 _3942_ (.B1(net750),
    .Y(_0542_),
    .A1(net689),
    .A2(net681));
 sg13g2_a21oi_1 _3943_ (.A1(net688),
    .A2(_2653_),
    .Y(_0173_),
    .B1(_0542_));
 sg13g2_nand2_1 _3944_ (.Y(_0543_),
    .A(net472),
    .B(net604));
 sg13g2_nand2_1 _3945_ (.Y(_0544_),
    .A(\core.delta_t[13] ),
    .B(_2739_));
 sg13g2_nand3b_1 _3946_ (.B(_0544_),
    .C(net681),
    .Y(_0545_),
    .A_N(_2740_));
 sg13g2_o21ai_1 _3947_ (.B1(_0545_),
    .Y(_0546_),
    .A1(net681),
    .A2(_0014_));
 sg13g2_xnor2_1 _3948_ (.Y(_0547_),
    .A(\core.delta_t[14] ),
    .B(_2740_));
 sg13g2_nand2_1 _3949_ (.Y(_0548_),
    .A(net680),
    .B(_0547_));
 sg13g2_o21ai_1 _3950_ (.B1(_0548_),
    .Y(_0549_),
    .A1(net680),
    .A2(_0015_));
 sg13g2_or2_2 _3951_ (.X(_0550_),
    .B(net594),
    .A(net601));
 sg13g2_nand2_1 _3952_ (.Y(_0551_),
    .A(\core.delta_t[12] ),
    .B(_2738_));
 sg13g2_nand3_1 _3953_ (.B(_2739_),
    .C(_0551_),
    .A(net681),
    .Y(_0552_));
 sg13g2_o21ai_1 _3954_ (.B1(_0552_),
    .Y(_0553_),
    .A1(\core.delta_t[15] ),
    .A2(_0013_));
 sg13g2_and3_1 _3955_ (.X(_0554_),
    .A(net601),
    .B(net594),
    .C(net612));
 sg13g2_and3_1 _3956_ (.X(_0555_),
    .A(net680),
    .B(_0015_),
    .C(_2740_));
 sg13g2_a21oi_1 _3957_ (.A1(net601),
    .A2(net594),
    .Y(_0556_),
    .B1(net609));
 sg13g2_nor2_2 _3958_ (.A(_0554_),
    .B(net610),
    .Y(_0557_));
 sg13g2_or2_2 _3959_ (.X(_0558_),
    .B(net610),
    .A(_0554_));
 sg13g2_and2_2 _3960_ (.A(_0550_),
    .B(_0557_),
    .X(_0559_));
 sg13g2_nand2_2 _3961_ (.Y(_0560_),
    .A(_0550_),
    .B(_0557_));
 sg13g2_nand2b_1 _3962_ (.Y(_0561_),
    .B(net594),
    .A_N(net612));
 sg13g2_a21oi_1 _3963_ (.A1(net601),
    .A2(_0561_),
    .Y(_0562_),
    .B1(net609));
 sg13g2_inv_2 _3964_ (.Y(_0563_),
    .A(net585));
 sg13g2_nor2b_1 _3965_ (.A(net612),
    .B_N(_0550_),
    .Y(_0564_));
 sg13g2_xnor2_1 _3966_ (.Y(_0565_),
    .A(_0556_),
    .B(_0564_));
 sg13g2_nor2_1 _3967_ (.A(_0028_),
    .B(net579),
    .Y(_0566_));
 sg13g2_a21oi_1 _3968_ (.A1(_2729_),
    .A2(net579),
    .Y(_0567_),
    .B1(_0566_));
 sg13g2_nand2_1 _3969_ (.Y(_0568_),
    .A(net584),
    .B(_0567_));
 sg13g2_a21oi_1 _3970_ (.A1(_2728_),
    .A2(net579),
    .Y(_0569_),
    .B1(net584));
 sg13g2_o21ai_1 _3971_ (.B1(_0569_),
    .Y(_0570_),
    .A1(_0026_),
    .A2(net579));
 sg13g2_nand2_1 _3972_ (.Y(_0571_),
    .A(_0568_),
    .B(_0570_));
 sg13g2_nor2_1 _3973_ (.A(net681),
    .B(_0011_),
    .Y(_0572_));
 sg13g2_nand2_1 _3974_ (.Y(_0573_),
    .A(\core.delta_t[11] ),
    .B(_2737_));
 sg13g2_nand3_1 _3975_ (.B(_2738_),
    .C(_0573_),
    .A(net681),
    .Y(_0574_));
 sg13g2_nor2b_2 _3976_ (.A(_0572_),
    .B_N(_0574_),
    .Y(_0575_));
 sg13g2_nand2b_2 _3977_ (.Y(_0576_),
    .B(_0574_),
    .A_N(_0572_));
 sg13g2_o21ai_1 _3978_ (.B1(\core.delta_t[10] ),
    .Y(_0577_),
    .A1(\core.delta_t[9] ),
    .A2(net682));
 sg13g2_nand3_1 _3979_ (.B(_2737_),
    .C(_0577_),
    .A(net680),
    .Y(_0578_));
 sg13g2_o21ai_1 _3980_ (.B1(_0578_),
    .Y(_0579_),
    .A1(net680),
    .A2(_0010_));
 sg13g2_inv_1 _3981_ (.Y(_0580_),
    .A(net621));
 sg13g2_or4_2 _3982_ (.A(\core.delta_t[9] ),
    .B(net682),
    .C(_0576_),
    .D(net621),
    .X(_0581_));
 sg13g2_nor3_1 _3983_ (.A(_0550_),
    .B(net612),
    .C(_0581_),
    .Y(_0582_));
 sg13g2_nor3_2 _3984_ (.A(net602),
    .B(net609),
    .C(_0582_),
    .Y(_0583_));
 sg13g2_or3_2 _3985_ (.A(net602),
    .B(net609),
    .C(_0582_),
    .X(_0584_));
 sg13g2_nand2b_1 _3986_ (.Y(_0585_),
    .B(\core.V_threshold[8] ),
    .A_N(net660));
 sg13g2_xnor2_1 _3987_ (.Y(_0586_),
    .A(net660),
    .B(\core.V_threshold[8] ));
 sg13g2_nor2_1 _3988_ (.A(_0550_),
    .B(net609),
    .Y(_0587_));
 sg13g2_a21oi_1 _3989_ (.A1(_0558_),
    .A2(_0586_),
    .Y(_0588_),
    .B1(_0584_));
 sg13g2_a22oi_1 _3990_ (.Y(_0589_),
    .B1(net583),
    .B2(_0023_),
    .A2(_0571_),
    .A1(_0559_));
 sg13g2_nand2_1 _3991_ (.Y(_0590_),
    .A(_0588_),
    .B(_0589_));
 sg13g2_a21oi_1 _3992_ (.A1(_0543_),
    .A2(_0590_),
    .Y(_0174_),
    .B1(net729));
 sg13g2_nor2_1 _3993_ (.A(_2729_),
    .B(net579),
    .Y(_0591_));
 sg13g2_a21oi_1 _3994_ (.A1(_0026_),
    .A2(net579),
    .Y(_0592_),
    .B1(_0591_));
 sg13g2_mux2_1 _3995_ (.A0(_0586_),
    .A1(_0028_),
    .S(net579),
    .X(_0593_));
 sg13g2_nor2_1 _3996_ (.A(_0563_),
    .B(_0593_),
    .Y(_0594_));
 sg13g2_a21oi_1 _3997_ (.A1(_0563_),
    .A2(_0592_),
    .Y(_0595_),
    .B1(_0594_));
 sg13g2_nor2_1 _3998_ (.A(_0560_),
    .B(_0595_),
    .Y(_0596_));
 sg13g2_nor2b_1 _3999_ (.A(\core.V_threshold[12] ),
    .B_N(net654),
    .Y(_0597_));
 sg13g2_xnor2_1 _4000_ (.Y(_0598_),
    .A(net654),
    .B(\core.V_threshold[12] ));
 sg13g2_xor2_1 _4001_ (.B(\core.V_threshold[11] ),
    .A(\core.V[11] ),
    .X(_0599_));
 sg13g2_nor2b_1 _4002_ (.A(\core.V_threshold[10] ),
    .B_N(net656),
    .Y(_0600_));
 sg13g2_xnor2_1 _4003_ (.Y(_0601_),
    .A(net656),
    .B(\core.V_threshold[10] ));
 sg13g2_nor2b_1 _4004_ (.A(\core.V_threshold[9] ),
    .B_N(net658),
    .Y(_0602_));
 sg13g2_xnor2_1 _4005_ (.Y(_0603_),
    .A(net657),
    .B(\core.V_threshold[9] ));
 sg13g2_a21oi_1 _4006_ (.A1(_0585_),
    .A2(_0603_),
    .Y(_0604_),
    .B1(_0602_));
 sg13g2_inv_1 _4007_ (.Y(_0605_),
    .A(_0604_));
 sg13g2_a21oi_1 _4008_ (.A1(_0601_),
    .A2(_0605_),
    .Y(_0606_),
    .B1(_0600_));
 sg13g2_nor2_1 _4009_ (.A(_0599_),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_a21oi_1 _4010_ (.A1(net655),
    .A2(_2638_),
    .Y(_0608_),
    .B1(_0607_));
 sg13g2_inv_1 _4011_ (.Y(_0609_),
    .A(_0608_));
 sg13g2_xnor2_1 _4012_ (.Y(_0610_),
    .A(_0598_),
    .B(_0608_));
 sg13g2_xnor2_1 _4013_ (.Y(_0611_),
    .A(_0599_),
    .B(_0606_));
 sg13g2_nor2_1 _4014_ (.A(net581),
    .B(_0610_),
    .Y(_0612_));
 sg13g2_a21oi_2 _4015_ (.B1(_0612_),
    .Y(_0613_),
    .A2(_0611_),
    .A1(net580));
 sg13g2_xnor2_1 _4016_ (.Y(_0614_),
    .A(_0601_),
    .B(_0604_));
 sg13g2_xor2_1 _4017_ (.B(_0603_),
    .A(_0585_),
    .X(_0615_));
 sg13g2_mux2_1 _4018_ (.A0(_0614_),
    .A1(_0615_),
    .S(net581),
    .X(_0616_));
 sg13g2_and2_1 _4019_ (.A(_0563_),
    .B(_0616_),
    .X(_0617_));
 sg13g2_a21oi_2 _4020_ (.B1(_0617_),
    .Y(_0618_),
    .A2(_0613_),
    .A1(net585));
 sg13g2_a21oi_1 _4021_ (.A1(_2728_),
    .A2(net583),
    .Y(_0619_),
    .B1(_0596_));
 sg13g2_o21ai_1 _4022_ (.B1(_0619_),
    .Y(_0620_),
    .A1(_0557_),
    .A2(_0618_));
 sg13g2_a22oi_1 _4023_ (.Y(_0621_),
    .B1(_0583_),
    .B2(_0620_),
    .A2(net604),
    .A1(net562));
 sg13g2_nor2_1 _4024_ (.A(net729),
    .B(_0621_),
    .Y(_0175_));
 sg13g2_nor2b_1 _4025_ (.A(\core.V_threshold[13] ),
    .B_N(net653),
    .Y(_0622_));
 sg13g2_xor2_1 _4026_ (.B(\core.V_threshold[13] ),
    .A(\core.V[13] ),
    .X(_0623_));
 sg13g2_a21oi_1 _4027_ (.A1(_0598_),
    .A2(_0609_),
    .Y(_0624_),
    .B1(_0597_));
 sg13g2_nor2_1 _4028_ (.A(_0623_),
    .B(_0624_),
    .Y(_0625_));
 sg13g2_xnor2_1 _4029_ (.Y(_0626_),
    .A(\core.V[14] ),
    .B(\core.V_threshold[14] ));
 sg13g2_o21ai_1 _4030_ (.B1(_0626_),
    .Y(_0627_),
    .A1(_0622_),
    .A2(_0625_));
 sg13g2_or3_1 _4031_ (.A(_0622_),
    .B(_0625_),
    .C(_0626_),
    .X(_0628_));
 sg13g2_and2_1 _4032_ (.A(_0627_),
    .B(_0628_),
    .X(_0629_));
 sg13g2_o21ai_1 _4033_ (.B1(_0627_),
    .Y(_0630_),
    .A1(_2629_),
    .A2(\core.V_threshold[14] ));
 sg13g2_xnor2_1 _4034_ (.Y(_0631_),
    .A(\core.V[15] ),
    .B(\core.V_threshold[15] ));
 sg13g2_xnor2_1 _4035_ (.Y(_0632_),
    .A(_0630_),
    .B(_0631_));
 sg13g2_nor2_1 _4036_ (.A(net581),
    .B(_0632_),
    .Y(_0633_));
 sg13g2_a21oi_1 _4037_ (.A1(net580),
    .A2(_0629_),
    .Y(_0634_),
    .B1(_0633_));
 sg13g2_nand2_1 _4038_ (.Y(_0635_),
    .A(net585),
    .B(_0632_));
 sg13g2_a21oi_1 _4039_ (.A1(_0563_),
    .A2(_0634_),
    .Y(_0636_),
    .B1(_0560_));
 sg13g2_xnor2_1 _4040_ (.Y(_0637_),
    .A(_0623_),
    .B(_0624_));
 sg13g2_nand2_1 _4041_ (.Y(_0638_),
    .A(net580),
    .B(_0610_));
 sg13g2_o21ai_1 _4042_ (.B1(_0638_),
    .Y(_0639_),
    .A1(net580),
    .A2(_0637_));
 sg13g2_nand2_1 _4043_ (.Y(_0640_),
    .A(net585),
    .B(_0639_));
 sg13g2_nor2_1 _4044_ (.A(net580),
    .B(_0611_),
    .Y(_0641_));
 sg13g2_a21oi_1 _4045_ (.A1(net580),
    .A2(_0614_),
    .Y(_0642_),
    .B1(_0641_));
 sg13g2_o21ai_1 _4046_ (.B1(_0640_),
    .Y(_0643_),
    .A1(net585),
    .A2(_0642_));
 sg13g2_a22oi_1 _4047_ (.Y(_0644_),
    .B1(_0643_),
    .B2(_0560_),
    .A2(_0636_),
    .A1(_0635_));
 sg13g2_nor2_1 _4048_ (.A(net581),
    .B(_0615_),
    .Y(_0645_));
 sg13g2_a21oi_1 _4049_ (.A1(net579),
    .A2(_0586_),
    .Y(_0646_),
    .B1(_0645_));
 sg13g2_nor2_1 _4050_ (.A(net584),
    .B(_0567_),
    .Y(_0647_));
 sg13g2_a21oi_1 _4051_ (.A1(net584),
    .A2(_0646_),
    .Y(_0648_),
    .B1(_0647_));
 sg13g2_a22oi_1 _4052_ (.Y(_0649_),
    .B1(_0643_),
    .B2(_0558_),
    .A2(net583),
    .A1(_2727_));
 sg13g2_o21ai_1 _4053_ (.B1(_0649_),
    .Y(_0650_),
    .A1(_0560_),
    .A2(_0648_));
 sg13g2_a22oi_1 _4054_ (.Y(_0651_),
    .B1(_0583_),
    .B2(_0650_),
    .A2(net604),
    .A1(net543));
 sg13g2_nor2_1 _4055_ (.A(net729),
    .B(net544),
    .Y(_0176_));
 sg13g2_nand2_1 _4056_ (.Y(_0652_),
    .A(net580),
    .B(_0637_));
 sg13g2_o21ai_1 _4057_ (.B1(_0652_),
    .Y(_0653_),
    .A1(net580),
    .A2(_0629_));
 sg13g2_inv_1 _4058_ (.Y(_0654_),
    .A(_0653_));
 sg13g2_nor2_1 _4059_ (.A(_0563_),
    .B(_0653_),
    .Y(_0655_));
 sg13g2_a21oi_2 _4060_ (.B1(_0655_),
    .Y(_0656_),
    .A2(_0613_),
    .A1(_0563_));
 sg13g2_nand2_1 _4061_ (.Y(_0657_),
    .A(net584),
    .B(_0616_));
 sg13g2_o21ai_1 _4062_ (.B1(_0657_),
    .Y(_0658_),
    .A1(net584),
    .A2(_0593_));
 sg13g2_inv_1 _4063_ (.Y(_0659_),
    .A(_0658_));
 sg13g2_a22oi_1 _4064_ (.Y(_0660_),
    .B1(_0658_),
    .B2(_0559_),
    .A2(net583),
    .A1(_2729_));
 sg13g2_o21ai_1 _4065_ (.B1(_0660_),
    .Y(_0661_),
    .A1(_0557_),
    .A2(_0656_));
 sg13g2_a22oi_1 _4066_ (.Y(_0662_),
    .B1(_0583_),
    .B2(_0661_),
    .A2(net604),
    .A1(net534));
 sg13g2_nor2_1 _4067_ (.A(net729),
    .B(net535),
    .Y(_0177_));
 sg13g2_o21ai_1 _4068_ (.B1(_0583_),
    .Y(_0663_),
    .A1(_0557_),
    .A2(_0610_));
 sg13g2_nor2_1 _4069_ (.A(net584),
    .B(_0646_),
    .Y(_0664_));
 sg13g2_a21oi_1 _4070_ (.A1(net584),
    .A2(_0642_),
    .Y(_0665_),
    .B1(_0664_));
 sg13g2_inv_1 _4071_ (.Y(_0666_),
    .A(_0665_));
 sg13g2_a221oi_1 _4072_ (.B2(_0559_),
    .C1(_0663_),
    .B1(_0666_),
    .A1(_0571_),
    .Y(_0667_),
    .A2(net583));
 sg13g2_a21oi_1 _4073_ (.A1(net427),
    .A2(net602),
    .Y(_0668_),
    .B1(_0667_));
 sg13g2_nor2_1 _4074_ (.A(net728),
    .B(_0668_),
    .Y(_0178_));
 sg13g2_a21o_1 _4075_ (.A2(_0637_),
    .A1(_0558_),
    .B1(_0584_),
    .X(_0669_));
 sg13g2_a221oi_1 _4076_ (.B2(_0559_),
    .C1(_0669_),
    .B1(_0618_),
    .A1(_0587_),
    .Y(_0670_),
    .A2(_0595_));
 sg13g2_a21oi_1 _4077_ (.A1(net441),
    .A2(net602),
    .Y(_0671_),
    .B1(_0670_));
 sg13g2_nor2_1 _4078_ (.A(net728),
    .B(_0671_),
    .Y(_0179_));
 sg13g2_nand2_1 _4079_ (.Y(_0672_),
    .A(net429),
    .B(net602));
 sg13g2_o21ai_1 _4080_ (.B1(_0583_),
    .Y(_0673_),
    .A1(_0557_),
    .A2(_0629_));
 sg13g2_a21oi_1 _4081_ (.A1(_0587_),
    .A2(_0648_),
    .Y(_0674_),
    .B1(_0673_));
 sg13g2_o21ai_1 _4082_ (.B1(_0674_),
    .Y(_0675_),
    .A1(_0560_),
    .A2(_0643_));
 sg13g2_a21oi_1 _4083_ (.A1(_0672_),
    .A2(_0675_),
    .Y(_0180_),
    .B1(net728));
 sg13g2_nor2_2 _4084_ (.A(_0584_),
    .B(_0632_),
    .Y(_0676_));
 sg13g2_inv_1 _4085_ (.Y(_0677_),
    .A(_0676_));
 sg13g2_a21oi_2 _4086_ (.B1(_0584_),
    .Y(_0678_),
    .A2(_0632_),
    .A1(_0558_));
 sg13g2_inv_1 _4087_ (.Y(_0679_),
    .A(_0678_));
 sg13g2_a22oi_1 _4088_ (.Y(_0680_),
    .B1(_0659_),
    .B2(net583),
    .A2(_0656_),
    .A1(_0559_));
 sg13g2_a22oi_1 _4089_ (.Y(_0681_),
    .B1(_0678_),
    .B2(_0680_),
    .A2(net602),
    .A1(net467));
 sg13g2_nor2_1 _4090_ (.A(net727),
    .B(_0681_),
    .Y(_0181_));
 sg13g2_nor2_1 _4091_ (.A(_0550_),
    .B(_0665_),
    .Y(_0682_));
 sg13g2_o21ai_1 _4092_ (.B1(_0559_),
    .Y(_0683_),
    .A1(_0563_),
    .A2(_0634_));
 sg13g2_a21oi_1 _4093_ (.A1(_0563_),
    .A2(_0639_),
    .Y(_0684_),
    .B1(_0683_));
 sg13g2_o21ai_1 _4094_ (.B1(_0557_),
    .Y(_0685_),
    .A1(_0682_),
    .A2(_0684_));
 sg13g2_a22oi_1 _4095_ (.Y(_0686_),
    .B1(_0678_),
    .B2(_0685_),
    .A2(net602),
    .A1(net458));
 sg13g2_nor2_1 _4096_ (.A(net727),
    .B(_0686_),
    .Y(_0182_));
 sg13g2_o21ai_1 _4097_ (.B1(_0635_),
    .Y(_0687_),
    .A1(net585),
    .A2(_0654_));
 sg13g2_a221oi_1 _4098_ (.B2(_0559_),
    .C1(_0679_),
    .B1(_0687_),
    .A1(net583),
    .Y(_0688_),
    .A2(_0618_));
 sg13g2_a21oi_1 _4099_ (.A1(net763),
    .A2(net604),
    .Y(_0689_),
    .B1(_0688_));
 sg13g2_nor2_1 _4100_ (.A(net729),
    .B(_0689_),
    .Y(_0183_));
 sg13g2_nand2_1 _4101_ (.Y(_0690_),
    .A(_0557_),
    .B(_0644_));
 sg13g2_a22oi_1 _4102_ (.Y(_0691_),
    .B1(_0678_),
    .B2(_0690_),
    .A2(net602),
    .A1(net811));
 sg13g2_nor2_1 _4103_ (.A(net727),
    .B(_0691_),
    .Y(_0184_));
 sg13g2_a22oi_1 _4104_ (.Y(_0692_),
    .B1(_0677_),
    .B2(_0550_),
    .A2(_0656_),
    .A1(net583));
 sg13g2_a22oi_1 _4105_ (.Y(_0693_),
    .B1(_0678_),
    .B2(_0692_),
    .A2(net603),
    .A1(net540));
 sg13g2_nor2_1 _4106_ (.A(net727),
    .B(_0693_),
    .Y(_0185_));
 sg13g2_a21oi_1 _4107_ (.A1(net556),
    .A2(net603),
    .Y(_0694_),
    .B1(_0676_));
 sg13g2_nor2_1 _4108_ (.A(net727),
    .B(_0694_),
    .Y(_0186_));
 sg13g2_a21oi_1 _4109_ (.A1(net770),
    .A2(net603),
    .Y(_0695_),
    .B1(_0676_));
 sg13g2_nor2_1 _4110_ (.A(net727),
    .B(_0695_),
    .Y(_0187_));
 sg13g2_a21oi_1 _4111_ (.A1(net783),
    .A2(net603),
    .Y(_0696_),
    .B1(_0676_));
 sg13g2_nor2_1 _4112_ (.A(net727),
    .B(_0696_),
    .Y(_0188_));
 sg13g2_a21oi_1 _4113_ (.A1(net822),
    .A2(net603),
    .Y(_0697_),
    .B1(_0676_));
 sg13g2_nor2_1 _4114_ (.A(net727),
    .B(_0697_),
    .Y(_0189_));
 sg13g2_and2_1 _4115_ (.A(\core.compute_state[3] ),
    .B(net740),
    .X(_0698_));
 sg13g2_nand2_2 _4116_ (.Y(_0699_),
    .A(net850),
    .B(net739));
 sg13g2_nor2_1 _4117_ (.A(net722),
    .B(_0699_),
    .Y(_0700_));
 sg13g2_nand2_2 _4118_ (.Y(_0701_),
    .A(net751),
    .B(_0698_));
 sg13g2_xnor2_1 _4119_ (.Y(_0702_),
    .A(\core.w[10] ),
    .B(\core.dw[10] ));
 sg13g2_nor2_1 _4120_ (.A(\core.w[9] ),
    .B(\core.dw[9] ),
    .Y(_0703_));
 sg13g2_and2_1 _4121_ (.A(\core.w[7] ),
    .B(\core.dw[7] ),
    .X(_0704_));
 sg13g2_or2_1 _4122_ (.X(_0705_),
    .B(\core.dw[7] ),
    .A(\core.w[7] ));
 sg13g2_nand2b_1 _4123_ (.Y(_0706_),
    .B(_0705_),
    .A_N(_0704_));
 sg13g2_and2_1 _4124_ (.A(\core.w[6] ),
    .B(\core.dw[6] ),
    .X(_0707_));
 sg13g2_nand2_1 _4125_ (.Y(_0708_),
    .A(\core.w[4] ),
    .B(\core.dw[4] ));
 sg13g2_nand2_1 _4126_ (.Y(_0709_),
    .A(\core.w[3] ),
    .B(\core.dw[3] ));
 sg13g2_xnor2_1 _4127_ (.Y(_0710_),
    .A(\core.w[3] ),
    .B(\core.dw[3] ));
 sg13g2_and2_1 _4128_ (.A(\core.w[2] ),
    .B(\core.dw[2] ),
    .X(_0711_));
 sg13g2_nand2_1 _4129_ (.Y(_0712_),
    .A(\core.w[1] ),
    .B(\core.dw[1] ));
 sg13g2_nand2_1 _4130_ (.Y(_0713_),
    .A(\core.w[0] ),
    .B(\core.dw[0] ));
 sg13g2_xnor2_1 _4131_ (.Y(_0714_),
    .A(\core.w[1] ),
    .B(\core.dw[1] ));
 sg13g2_o21ai_1 _4132_ (.B1(_0712_),
    .Y(_0715_),
    .A1(_0713_),
    .A2(_0714_));
 sg13g2_xor2_1 _4133_ (.B(\core.dw[2] ),
    .A(\core.w[2] ),
    .X(_0716_));
 sg13g2_a21oi_1 _4134_ (.A1(_0715_),
    .A2(_0716_),
    .Y(_0717_),
    .B1(_0711_));
 sg13g2_o21ai_1 _4135_ (.B1(_0709_),
    .Y(_0718_),
    .A1(_0710_),
    .A2(_0717_));
 sg13g2_inv_1 _4136_ (.Y(_0719_),
    .A(_0718_));
 sg13g2_xnor2_1 _4137_ (.Y(_0720_),
    .A(\core.w[4] ),
    .B(\core.dw[4] ));
 sg13g2_o21ai_1 _4138_ (.B1(_0708_),
    .Y(_0721_),
    .A1(_0719_),
    .A2(_0720_));
 sg13g2_xnor2_1 _4139_ (.Y(_0722_),
    .A(\core.w[5] ),
    .B(\core.dw[5] ));
 sg13g2_nor2b_1 _4140_ (.A(_0722_),
    .B_N(_0721_),
    .Y(_0723_));
 sg13g2_a21o_1 _4141_ (.A2(\core.dw[5] ),
    .A1(\core.w[5] ),
    .B1(_0723_),
    .X(_0724_));
 sg13g2_or2_1 _4142_ (.X(_0725_),
    .B(\core.dw[6] ),
    .A(\core.w[6] ));
 sg13g2_nand2b_1 _4143_ (.Y(_0726_),
    .B(_0725_),
    .A_N(_0707_));
 sg13g2_a21o_1 _4144_ (.A2(_0725_),
    .A1(_0724_),
    .B1(_0707_),
    .X(_0727_));
 sg13g2_a21o_1 _4145_ (.A2(_0727_),
    .A1(_0705_),
    .B1(_0704_),
    .X(_0728_));
 sg13g2_xor2_1 _4146_ (.B(\core.dw[8] ),
    .A(\core.w[8] ),
    .X(_0729_));
 sg13g2_and2_1 _4147_ (.A(_0728_),
    .B(_0729_),
    .X(_0730_));
 sg13g2_a21oi_1 _4148_ (.A1(\core.w[8] ),
    .A2(\core.dw[8] ),
    .Y(_0731_),
    .B1(_0730_));
 sg13g2_a221oi_1 _4149_ (.B2(\core.w[8] ),
    .C1(_0730_),
    .B1(\core.dw[8] ),
    .A1(\core.w[9] ),
    .Y(_0732_),
    .A2(\core.dw[9] ));
 sg13g2_nor2_1 _4150_ (.A(_0703_),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_nor3_1 _4151_ (.A(_0702_),
    .B(_0703_),
    .C(_0732_),
    .Y(_0734_));
 sg13g2_xnor2_1 _4152_ (.Y(_0735_),
    .A(_0702_),
    .B(_0733_));
 sg13g2_a22oi_1 _4153_ (.Y(_0736_),
    .B1(net629),
    .B2(_0735_),
    .A2(net650),
    .A1(net440));
 sg13g2_inv_1 _4154_ (.Y(_0190_),
    .A(_0736_));
 sg13g2_a21oi_1 _4155_ (.A1(\core.w[10] ),
    .A2(\core.dw[10] ),
    .Y(_0737_),
    .B1(_0734_));
 sg13g2_nand2_1 _4156_ (.Y(_0738_),
    .A(\core.w[11] ),
    .B(\core.dw[11] ));
 sg13g2_nor2_1 _4157_ (.A(\core.w[11] ),
    .B(\core.dw[11] ),
    .Y(_0739_));
 sg13g2_xor2_1 _4158_ (.B(\core.dw[11] ),
    .A(\core.w[11] ),
    .X(_0740_));
 sg13g2_xnor2_1 _4159_ (.Y(_0741_),
    .A(_0737_),
    .B(_0740_));
 sg13g2_a22oi_1 _4160_ (.Y(_0742_),
    .B1(net630),
    .B2(_0741_),
    .A2(net650),
    .A1(net492));
 sg13g2_inv_1 _4161_ (.Y(_0191_),
    .A(_0742_));
 sg13g2_and2_1 _4162_ (.A(\core.w[12] ),
    .B(\core.dw[12] ),
    .X(_0743_));
 sg13g2_xor2_1 _4163_ (.B(\core.dw[12] ),
    .A(\core.w[12] ),
    .X(_0744_));
 sg13g2_o21ai_1 _4164_ (.B1(_0738_),
    .Y(_0745_),
    .A1(_0737_),
    .A2(_0739_));
 sg13g2_xor2_1 _4165_ (.B(_0745_),
    .A(_0744_),
    .X(_0746_));
 sg13g2_a22oi_1 _4166_ (.Y(_0747_),
    .B1(net629),
    .B2(_0746_),
    .A2(net650),
    .A1(net482));
 sg13g2_inv_1 _4167_ (.Y(_0192_),
    .A(_0747_));
 sg13g2_nand2_1 _4168_ (.Y(_0748_),
    .A(net384),
    .B(net650));
 sg13g2_a21o_1 _4169_ (.A2(_0745_),
    .A1(_0744_),
    .B1(_0743_),
    .X(_0749_));
 sg13g2_xor2_1 _4170_ (.B(\core.dw[13] ),
    .A(\core.w[13] ),
    .X(_0750_));
 sg13g2_xnor2_1 _4171_ (.Y(_0751_),
    .A(_0749_),
    .B(_0750_));
 sg13g2_inv_1 _4172_ (.Y(_0752_),
    .A(_0751_));
 sg13g2_o21ai_1 _4173_ (.B1(_0748_),
    .Y(_0193_),
    .A1(_0701_),
    .A2(_0751_));
 sg13g2_nand2_1 _4174_ (.Y(_0753_),
    .A(net419),
    .B(net649));
 sg13g2_nand2_1 _4175_ (.Y(_0754_),
    .A(\core.w[14] ),
    .B(\core.dw[14] ));
 sg13g2_xnor2_1 _4176_ (.Y(_0755_),
    .A(\core.w[14] ),
    .B(\core.dw[14] ));
 sg13g2_a21o_1 _4177_ (.A2(\core.dw[13] ),
    .A1(\core.w[13] ),
    .B1(_0749_),
    .X(_0756_));
 sg13g2_o21ai_1 _4178_ (.B1(_0756_),
    .Y(_0757_),
    .A1(\core.w[13] ),
    .A2(\core.dw[13] ));
 sg13g2_xnor2_1 _4179_ (.Y(_0758_),
    .A(_0755_),
    .B(_0757_));
 sg13g2_o21ai_1 _4180_ (.B1(_0753_),
    .Y(_0194_),
    .A1(net628),
    .A2(_0758_));
 sg13g2_o21ai_1 _4181_ (.B1(_0754_),
    .Y(_0759_),
    .A1(_0755_),
    .A2(_0757_));
 sg13g2_xnor2_1 _4182_ (.Y(_0760_),
    .A(\core.w[15] ),
    .B(\core.dw[15] ));
 sg13g2_xnor2_1 _4183_ (.Y(_0761_),
    .A(_0759_),
    .B(_0760_));
 sg13g2_a22oi_1 _4184_ (.Y(_0195_),
    .B1(net629),
    .B2(_0761_),
    .A2(net649),
    .A1(_2649_));
 sg13g2_and2_1 _4185_ (.A(\core.V[10] ),
    .B(\core.dV[10] ),
    .X(_0762_));
 sg13g2_xor2_1 _4186_ (.B(\core.dV[10] ),
    .A(net656),
    .X(_0763_));
 sg13g2_nor2_1 _4187_ (.A(net657),
    .B(\core.dV[9] ),
    .Y(_0764_));
 sg13g2_and2_1 _4188_ (.A(net660),
    .B(\core.dV[8] ),
    .X(_0765_));
 sg13g2_nand2_1 _4189_ (.Y(_0766_),
    .A(net663),
    .B(\core.dV[7] ));
 sg13g2_xnor2_1 _4190_ (.Y(_0767_),
    .A(net663),
    .B(\core.dV[7] ));
 sg13g2_and2_1 _4191_ (.A(net665),
    .B(\core.dV[6] ),
    .X(_0768_));
 sg13g2_or2_1 _4192_ (.X(_0769_),
    .B(\core.dV[6] ),
    .A(net665));
 sg13g2_nand2b_1 _4193_ (.Y(_0770_),
    .B(_0769_),
    .A_N(_0768_));
 sg13g2_xnor2_1 _4194_ (.Y(_0771_),
    .A(net667),
    .B(\core.dV[5] ));
 sg13g2_nand2_1 _4195_ (.Y(_0772_),
    .A(net669),
    .B(\core.dV[4] ));
 sg13g2_xor2_1 _4196_ (.B(\core.dV[4] ),
    .A(net669),
    .X(_0773_));
 sg13g2_and2_1 _4197_ (.A(net672),
    .B(\core.dV[3] ),
    .X(_0774_));
 sg13g2_nand2_1 _4198_ (.Y(_0775_),
    .A(net674),
    .B(\core.dV[2] ));
 sg13g2_nand2_1 _4199_ (.Y(_0776_),
    .A(net675),
    .B(\core.dV[1] ));
 sg13g2_xor2_1 _4200_ (.B(\core.dV[1] ),
    .A(net675),
    .X(_0777_));
 sg13g2_nand3_1 _4201_ (.B(\core.dV[0] ),
    .C(_0777_),
    .A(net678),
    .Y(_0778_));
 sg13g2_and2_1 _4202_ (.A(_0776_),
    .B(_0778_),
    .X(_0779_));
 sg13g2_xnor2_1 _4203_ (.Y(_0780_),
    .A(net674),
    .B(\core.dV[2] ));
 sg13g2_o21ai_1 _4204_ (.B1(_0775_),
    .Y(_0781_),
    .A1(_0779_),
    .A2(_0780_));
 sg13g2_xor2_1 _4205_ (.B(\core.dV[3] ),
    .A(net672),
    .X(_0782_));
 sg13g2_a21o_1 _4206_ (.A2(_0782_),
    .A1(_0781_),
    .B1(_0774_),
    .X(_0783_));
 sg13g2_nand2_1 _4207_ (.Y(_0784_),
    .A(_0773_),
    .B(_0783_));
 sg13g2_nand2_1 _4208_ (.Y(_0785_),
    .A(_0772_),
    .B(_0784_));
 sg13g2_a21oi_1 _4209_ (.A1(_0772_),
    .A2(_0784_),
    .Y(_0786_),
    .B1(_0771_));
 sg13g2_a21o_1 _4210_ (.A2(\core.dV[5] ),
    .A1(net667),
    .B1(_0786_),
    .X(_0787_));
 sg13g2_a21o_1 _4211_ (.A2(_0787_),
    .A1(_0769_),
    .B1(_0768_),
    .X(_0788_));
 sg13g2_inv_1 _4212_ (.Y(_0789_),
    .A(_0788_));
 sg13g2_o21ai_1 _4213_ (.B1(_0766_),
    .Y(_0790_),
    .A1(_0767_),
    .A2(_0789_));
 sg13g2_xor2_1 _4214_ (.B(\core.dV[8] ),
    .A(net660),
    .X(_0791_));
 sg13g2_a21o_1 _4215_ (.A2(_0791_),
    .A1(_0790_),
    .B1(_0765_),
    .X(_0792_));
 sg13g2_a21oi_1 _4216_ (.A1(net657),
    .A2(\core.dV[9] ),
    .Y(_0793_),
    .B1(_0792_));
 sg13g2_nor2_1 _4217_ (.A(_0764_),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_xnor2_1 _4218_ (.Y(_0795_),
    .A(_0763_),
    .B(_0794_));
 sg13g2_a22oi_1 _4219_ (.Y(_0196_),
    .B1(net629),
    .B2(_0795_),
    .A2(net649),
    .A1(_2648_));
 sg13g2_a21oi_2 _4220_ (.B1(_0762_),
    .Y(_0796_),
    .A2(_0794_),
    .A1(_0763_));
 sg13g2_nand2_1 _4221_ (.Y(_0797_),
    .A(\core.V[11] ),
    .B(\core.dV[11] ));
 sg13g2_nor2_1 _4222_ (.A(net655),
    .B(\core.dV[11] ),
    .Y(_0798_));
 sg13g2_xnor2_1 _4223_ (.Y(_0799_),
    .A(net655),
    .B(\core.dV[11] ));
 sg13g2_xnor2_1 _4224_ (.Y(_0800_),
    .A(_0796_),
    .B(_0799_));
 sg13g2_a22oi_1 _4225_ (.Y(_0197_),
    .B1(net629),
    .B2(_0800_),
    .A2(net649),
    .A1(_2647_));
 sg13g2_and2_1 _4226_ (.A(\core.V[12] ),
    .B(\core.dV[12] ),
    .X(_0801_));
 sg13g2_xor2_1 _4227_ (.B(\core.dV[12] ),
    .A(net654),
    .X(_0802_));
 sg13g2_o21ai_1 _4228_ (.B1(_0797_),
    .Y(_0803_),
    .A1(_0796_),
    .A2(_0798_));
 sg13g2_xnor2_1 _4229_ (.Y(_0804_),
    .A(_0802_),
    .B(_0803_));
 sg13g2_a22oi_1 _4230_ (.Y(_0198_),
    .B1(net629),
    .B2(_0804_),
    .A2(net649),
    .A1(_2646_));
 sg13g2_a21o_1 _4231_ (.A2(_0803_),
    .A1(_0802_),
    .B1(_0801_),
    .X(_0805_));
 sg13g2_xor2_1 _4232_ (.B(\core.dV[13] ),
    .A(net653),
    .X(_0806_));
 sg13g2_xnor2_1 _4233_ (.Y(_0807_),
    .A(_0805_),
    .B(_0806_));
 sg13g2_a22oi_1 _4234_ (.Y(_0199_),
    .B1(net629),
    .B2(_0807_),
    .A2(net649),
    .A1(_2645_));
 sg13g2_nand2_1 _4235_ (.Y(_0808_),
    .A(net330),
    .B(net649));
 sg13g2_nand2_1 _4236_ (.Y(_0809_),
    .A(\core.V[14] ),
    .B(\core.dV[14] ));
 sg13g2_xnor2_1 _4237_ (.Y(_0810_),
    .A(\core.V[14] ),
    .B(\core.dV[14] ));
 sg13g2_a21o_1 _4238_ (.A2(\core.dV[13] ),
    .A1(net653),
    .B1(_0805_),
    .X(_0811_));
 sg13g2_o21ai_1 _4239_ (.B1(_0811_),
    .Y(_0812_),
    .A1(net653),
    .A2(\core.dV[13] ));
 sg13g2_xnor2_1 _4240_ (.Y(_0813_),
    .A(_0810_),
    .B(_0812_));
 sg13g2_o21ai_1 _4241_ (.B1(_0808_),
    .Y(_0200_),
    .A1(_0701_),
    .A2(_0813_));
 sg13g2_o21ai_1 _4242_ (.B1(_0809_),
    .Y(_0814_),
    .A1(_0810_),
    .A2(_0812_));
 sg13g2_xor2_1 _4243_ (.B(\core.dV[15] ),
    .A(\core.V[15] ),
    .X(_0815_));
 sg13g2_xnor2_1 _4244_ (.Y(_0816_),
    .A(_0814_),
    .B(_0815_));
 sg13g2_a22oi_1 _4245_ (.Y(_0817_),
    .B1(net629),
    .B2(_0816_),
    .A2(net649),
    .A1(net405));
 sg13g2_inv_1 _4246_ (.Y(_0201_),
    .A(_0817_));
 sg13g2_nor2_1 _4247_ (.A(\core.tau_w[15] ),
    .B(_0016_),
    .Y(_0818_));
 sg13g2_or3_1 _4248_ (.A(\core.tau_w[11] ),
    .B(\core.tau_w[10] ),
    .C(\core.tau_w[9] ),
    .X(_0819_));
 sg13g2_nor2_2 _4249_ (.A(\core.tau_w[8] ),
    .B(_0819_),
    .Y(_0820_));
 sg13g2_nand2b_1 _4250_ (.Y(_0821_),
    .B(_0820_),
    .A_N(\core.tau_w[12] ));
 sg13g2_xnor2_1 _4251_ (.Y(_0822_),
    .A(\core.tau_w[12] ),
    .B(_0820_));
 sg13g2_a21oi_1 _4252_ (.A1(\core.tau_w[15] ),
    .A2(_0822_),
    .Y(_0823_),
    .B1(_0818_));
 sg13g2_a21oi_1 _4253_ (.A1(_0016_),
    .A2(_0820_),
    .Y(_0824_),
    .B1(_2705_));
 sg13g2_xnor2_1 _4254_ (.Y(_0825_),
    .A(\core.tau_w[13] ),
    .B(_0824_));
 sg13g2_and2_1 _4255_ (.A(_0823_),
    .B(_0825_),
    .X(_0826_));
 sg13g2_or2_1 _4256_ (.X(_0827_),
    .B(_0017_),
    .A(\core.tau_w[15] ));
 sg13g2_o21ai_1 _4257_ (.B1(_0827_),
    .Y(_0828_),
    .A1(_2705_),
    .A2(\core.tau_w[14] ));
 sg13g2_nor3_2 _4258_ (.A(_2705_),
    .B(\core.tau_w[13] ),
    .C(_0821_),
    .Y(_0829_));
 sg13g2_nand2b_1 _4259_ (.Y(_0830_),
    .B(_0829_),
    .A_N(\core.tau_w[14] ));
 sg13g2_o21ai_1 _4260_ (.B1(_0830_),
    .Y(_0831_),
    .A1(_0828_),
    .A2(_0829_));
 sg13g2_inv_1 _4261_ (.Y(_0832_),
    .A(_0831_));
 sg13g2_nand3_1 _4262_ (.B(_0826_),
    .C(_0831_),
    .A(_0820_),
    .Y(_0833_));
 sg13g2_nor4_1 _4263_ (.A(\core.tau_w[14] ),
    .B(\core.tau_w[13] ),
    .C(\core.tau_w[12] ),
    .D(_0819_),
    .Y(_0834_));
 sg13g2_nor3_2 _4264_ (.A(\core.tau_w[15] ),
    .B(net638),
    .C(_0834_),
    .Y(_0835_));
 sg13g2_and2_2 _4265_ (.A(_0833_),
    .B(_0835_),
    .X(_0836_));
 sg13g2_nand2_1 _4266_ (.Y(_0837_),
    .A(_0833_),
    .B(_0835_));
 sg13g2_or2_1 _4267_ (.X(_0838_),
    .B(_0825_),
    .A(_0823_));
 sg13g2_nor2_1 _4268_ (.A(_0831_),
    .B(_0838_),
    .Y(_0839_));
 sg13g2_nand2_2 _4269_ (.Y(_0840_),
    .A(_0017_),
    .B(_0829_));
 sg13g2_nor2b_2 _4270_ (.A(_0839_),
    .B_N(_0840_),
    .Y(_0841_));
 sg13g2_o21ai_1 _4271_ (.B1(_0840_),
    .Y(_0842_),
    .A1(_0831_),
    .A2(_0838_));
 sg13g2_nor2_1 _4272_ (.A(_0825_),
    .B(_0832_),
    .Y(_0843_));
 sg13g2_nand2_1 _4273_ (.Y(_0844_),
    .A(_0838_),
    .B(_0840_));
 sg13g2_nor2_2 _4274_ (.A(_0843_),
    .B(_0844_),
    .Y(_0845_));
 sg13g2_inv_1 _4275_ (.Y(_0846_),
    .A(net582));
 sg13g2_a221oi_1 _4276_ (.B2(_0823_),
    .C1(_0839_),
    .B1(_0843_),
    .A1(_0826_),
    .Y(_0847_),
    .A2(_0832_));
 sg13g2_nor2_1 _4277_ (.A(\core.tau_w[14] ),
    .B(_0840_),
    .Y(_0848_));
 sg13g2_mux2_1 _4278_ (.A0(_0840_),
    .A1(_0848_),
    .S(_0847_),
    .X(_0849_));
 sg13g2_nand2_2 _4279_ (.Y(_0850_),
    .A(net678),
    .B(net710));
 sg13g2_and2_2 _4280_ (.A(net676),
    .B(net708),
    .X(_0851_));
 sg13g2_nor2b_1 _4281_ (.A(_0850_),
    .B_N(_0851_),
    .Y(_0852_));
 sg13g2_nand2b_1 _4282_ (.Y(_0853_),
    .B(_0851_),
    .A_N(_0850_));
 sg13g2_a22oi_1 _4283_ (.Y(_0854_),
    .B1(net710),
    .B2(\core.V[1] ),
    .A2(net708),
    .A1(net679));
 sg13g2_nand3b_1 _4284_ (.B(_0019_),
    .C(_0853_),
    .Y(_0855_),
    .A_N(_0854_));
 sg13g2_nand2_1 _4285_ (.Y(_0856_),
    .A(net673),
    .B(net710));
 sg13g2_nand2_1 _4286_ (.Y(_0857_),
    .A(net679),
    .B(net706));
 sg13g2_nand3_1 _4287_ (.B(net706),
    .C(_0851_),
    .A(net679),
    .Y(_0858_));
 sg13g2_xnor2_1 _4288_ (.Y(_0859_),
    .A(_0851_),
    .B(_0857_));
 sg13g2_nand2b_1 _4289_ (.Y(_0860_),
    .B(_0859_),
    .A_N(_0856_));
 sg13g2_xnor2_1 _4290_ (.Y(_0861_),
    .A(_0856_),
    .B(_0859_));
 sg13g2_nand2_1 _4291_ (.Y(_0862_),
    .A(_0020_),
    .B(_0861_));
 sg13g2_xnor2_1 _4292_ (.Y(_0863_),
    .A(_0020_),
    .B(_0861_));
 sg13g2_nor2_1 _4293_ (.A(_0855_),
    .B(_0863_),
    .Y(_0864_));
 sg13g2_nand2_1 _4294_ (.Y(_0865_),
    .A(net670),
    .B(net712));
 sg13g2_nand2_2 _4295_ (.Y(_0866_),
    .A(net674),
    .B(net712));
 sg13g2_nand2_1 _4296_ (.Y(_0867_),
    .A(net670),
    .B(net714));
 sg13g2_nand2_1 _4297_ (.Y(_0868_),
    .A(net668),
    .B(net717));
 sg13g2_xor2_1 _4298_ (.B(_0867_),
    .A(_0866_),
    .X(_0869_));
 sg13g2_nand2b_1 _4299_ (.Y(_0870_),
    .B(_0869_),
    .A_N(_0868_));
 sg13g2_o21ai_1 _4300_ (.B1(_0870_),
    .Y(_0871_),
    .A1(_0866_),
    .A2(_0867_));
 sg13g2_nand2_1 _4301_ (.Y(_0872_),
    .A(net666),
    .B(net717));
 sg13g2_nand2_1 _4302_ (.Y(_0873_),
    .A(net668),
    .B(net712));
 sg13g2_nand2_1 _4303_ (.Y(_0874_),
    .A(net668),
    .B(net714));
 sg13g2_or2_1 _4304_ (.X(_0875_),
    .B(_0873_),
    .A(_0867_));
 sg13g2_xnor2_1 _4305_ (.Y(_0876_),
    .A(_0865_),
    .B(_0874_));
 sg13g2_xor2_1 _4306_ (.B(_0876_),
    .A(_0872_),
    .X(_0877_));
 sg13g2_and2_1 _4307_ (.A(_0852_),
    .B(_0877_),
    .X(_0878_));
 sg13g2_xnor2_1 _4308_ (.Y(_0879_),
    .A(_0853_),
    .B(_0877_));
 sg13g2_xnor2_1 _4309_ (.Y(_0880_),
    .A(_0871_),
    .B(_0879_));
 sg13g2_xor2_1 _4310_ (.B(_0863_),
    .A(_0855_),
    .X(_0881_));
 sg13g2_nor2b_1 _4311_ (.A(_0880_),
    .B_N(_0881_),
    .Y(_0882_));
 sg13g2_nor2_1 _4312_ (.A(_0864_),
    .B(_0882_),
    .Y(_0883_));
 sg13g2_nand2_1 _4313_ (.Y(_0884_),
    .A(net677),
    .B(net705));
 sg13g2_or2_1 _4314_ (.X(_0885_),
    .B(_0884_),
    .A(\core.w[6] ));
 sg13g2_xor2_1 _4315_ (.B(_0884_),
    .A(\core.w[6] ),
    .X(_0886_));
 sg13g2_and2_1 _4316_ (.A(net670),
    .B(net710),
    .X(_0887_));
 sg13g2_and2_1 _4317_ (.A(net673),
    .B(net706),
    .X(_0888_));
 sg13g2_nand2_1 _4318_ (.Y(_0889_),
    .A(net673),
    .B(net706));
 sg13g2_a22oi_1 _4319_ (.Y(_0890_),
    .B1(net708),
    .B2(net673),
    .A2(net706),
    .A1(net676));
 sg13g2_a21oi_1 _4320_ (.A1(_0851_),
    .A2(_0888_),
    .Y(_0891_),
    .B1(_0890_));
 sg13g2_xor2_1 _4321_ (.B(_0891_),
    .A(_0887_),
    .X(_0892_));
 sg13g2_nand2_1 _4322_ (.Y(_0893_),
    .A(_0886_),
    .B(_0892_));
 sg13g2_xnor2_1 _4323_ (.Y(_0894_),
    .A(_0886_),
    .B(_0892_));
 sg13g2_nor2_1 _4324_ (.A(_0862_),
    .B(_0894_),
    .Y(_0895_));
 sg13g2_xor2_1 _4325_ (.B(_0894_),
    .A(_0862_),
    .X(_0896_));
 sg13g2_o21ai_1 _4326_ (.B1(_0875_),
    .Y(_0897_),
    .A1(_0872_),
    .A2(_0876_));
 sg13g2_and2_1 _4327_ (.A(_0858_),
    .B(_0860_),
    .X(_0898_));
 sg13g2_nand2_1 _4328_ (.Y(_0899_),
    .A(net665),
    .B(net717));
 sg13g2_nand2_1 _4329_ (.Y(_0900_),
    .A(net667),
    .B(net712));
 sg13g2_nand2_1 _4330_ (.Y(_0901_),
    .A(net667),
    .B(net714));
 sg13g2_or2_1 _4331_ (.X(_0902_),
    .B(_0900_),
    .A(_0874_));
 sg13g2_xnor2_1 _4332_ (.Y(_0903_),
    .A(_0873_),
    .B(_0901_));
 sg13g2_xor2_1 _4333_ (.B(_0903_),
    .A(_0899_),
    .X(_0904_));
 sg13g2_nor2b_1 _4334_ (.A(_0898_),
    .B_N(_0904_),
    .Y(_0905_));
 sg13g2_xnor2_1 _4335_ (.Y(_0906_),
    .A(_0898_),
    .B(_0904_));
 sg13g2_xor2_1 _4336_ (.B(_0906_),
    .A(_0897_),
    .X(_0907_));
 sg13g2_xnor2_1 _4337_ (.Y(_0908_),
    .A(_0896_),
    .B(_0907_));
 sg13g2_nor2_1 _4338_ (.A(_0883_),
    .B(_0908_),
    .Y(_0909_));
 sg13g2_a21o_1 _4339_ (.A2(_0879_),
    .A1(_0871_),
    .B1(_0878_),
    .X(_0910_));
 sg13g2_xor2_1 _4340_ (.B(_0908_),
    .A(_0883_),
    .X(_0911_));
 sg13g2_a21oi_1 _4341_ (.A1(_0910_),
    .A2(_0911_),
    .Y(_0912_),
    .B1(_0909_));
 sg13g2_a21o_1 _4342_ (.A2(_0906_),
    .A1(_0897_),
    .B1(_0905_),
    .X(_0913_));
 sg13g2_a21oi_1 _4343_ (.A1(_0896_),
    .A2(_0907_),
    .Y(_0914_),
    .B1(_0895_));
 sg13g2_o21ai_1 _4344_ (.B1(_0902_),
    .Y(_0915_),
    .A1(_0899_),
    .A2(_0903_));
 sg13g2_a22oi_1 _4345_ (.Y(_0916_),
    .B1(_0891_),
    .B2(_0887_),
    .A2(_0888_),
    .A1(_0851_));
 sg13g2_nand2_1 _4346_ (.Y(_0917_),
    .A(net662),
    .B(net717));
 sg13g2_nand2_1 _4347_ (.Y(_0918_),
    .A(net664),
    .B(net712));
 sg13g2_nand2_1 _4348_ (.Y(_0919_),
    .A(net664),
    .B(net714));
 sg13g2_xor2_1 _4349_ (.B(_0919_),
    .A(_0900_),
    .X(_0920_));
 sg13g2_nand2b_1 _4350_ (.Y(_0921_),
    .B(_0920_),
    .A_N(_0917_));
 sg13g2_xnor2_1 _4351_ (.Y(_0922_),
    .A(_0917_),
    .B(_0920_));
 sg13g2_nor2b_1 _4352_ (.A(_0916_),
    .B_N(_0922_),
    .Y(_0923_));
 sg13g2_xnor2_1 _4353_ (.Y(_0924_),
    .A(_0916_),
    .B(_0922_));
 sg13g2_xnor2_1 _4354_ (.Y(_0925_),
    .A(_0915_),
    .B(_0924_));
 sg13g2_nand2_1 _4355_ (.Y(_0926_),
    .A(net669),
    .B(net710));
 sg13g2_nand2_1 _4356_ (.Y(_0927_),
    .A(net670),
    .B(net706));
 sg13g2_nand2_1 _4357_ (.Y(_0928_),
    .A(net670),
    .B(net708));
 sg13g2_xnor2_1 _4358_ (.Y(_0929_),
    .A(_0888_),
    .B(_0928_));
 sg13g2_nand2b_1 _4359_ (.Y(_0930_),
    .B(_0929_),
    .A_N(_0926_));
 sg13g2_xnor2_1 _4360_ (.Y(_0931_),
    .A(_0926_),
    .B(_0929_));
 sg13g2_and2_1 _4361_ (.A(net676),
    .B(net705),
    .X(_0932_));
 sg13g2_nor2_1 _4362_ (.A(net677),
    .B(net651),
    .Y(_0933_));
 sg13g2_nor3_1 _4363_ (.A(net677),
    .B(\core.w[7] ),
    .C(net651),
    .Y(_0934_));
 sg13g2_xnor2_1 _4364_ (.Y(_0935_),
    .A(\core.w[7] ),
    .B(_0933_));
 sg13g2_xor2_1 _4365_ (.B(_0935_),
    .A(_0932_),
    .X(_0936_));
 sg13g2_nor2b_1 _4366_ (.A(_0885_),
    .B_N(_0936_),
    .Y(_0937_));
 sg13g2_xnor2_1 _4367_ (.Y(_0938_),
    .A(_0885_),
    .B(_0936_));
 sg13g2_xnor2_1 _4368_ (.Y(_0939_),
    .A(_0931_),
    .B(_0938_));
 sg13g2_nor2_1 _4369_ (.A(_0893_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_xor2_1 _4370_ (.B(_0939_),
    .A(_0893_),
    .X(_0941_));
 sg13g2_nor2b_1 _4371_ (.A(_0925_),
    .B_N(_0941_),
    .Y(_0942_));
 sg13g2_xnor2_1 _4372_ (.Y(_0943_),
    .A(_0925_),
    .B(_0941_));
 sg13g2_nor2b_1 _4373_ (.A(_0914_),
    .B_N(_0943_),
    .Y(_0944_));
 sg13g2_xnor2_1 _4374_ (.Y(_0945_),
    .A(_0914_),
    .B(_0943_));
 sg13g2_xnor2_1 _4375_ (.Y(_0946_),
    .A(_0913_),
    .B(_0945_));
 sg13g2_nor2_1 _4376_ (.A(_0912_),
    .B(_0946_),
    .Y(_0947_));
 sg13g2_xor2_1 _4377_ (.B(_0946_),
    .A(_0912_),
    .X(_0948_));
 sg13g2_a21oi_1 _4378_ (.A1(\core.param_a[15] ),
    .A2(_0948_),
    .Y(_0949_),
    .B1(_0947_));
 sg13g2_a21oi_1 _4379_ (.A1(_0915_),
    .A2(_0924_),
    .Y(_0950_),
    .B1(_0923_));
 sg13g2_nor2_1 _4380_ (.A(_0940_),
    .B(_0942_),
    .Y(_0951_));
 sg13g2_o21ai_1 _4381_ (.B1(_0921_),
    .Y(_0952_),
    .A1(_0900_),
    .A2(_0919_));
 sg13g2_o21ai_1 _4382_ (.B1(_0930_),
    .Y(_0953_),
    .A1(_0889_),
    .A2(_0928_));
 sg13g2_nand2_1 _4383_ (.Y(_0954_),
    .A(net661),
    .B(net717));
 sg13g2_nand2_1 _4384_ (.Y(_0955_),
    .A(net662),
    .B(net712));
 sg13g2_nand2_1 _4385_ (.Y(_0956_),
    .A(net662),
    .B(net714));
 sg13g2_xor2_1 _4386_ (.B(_0956_),
    .A(_0918_),
    .X(_0957_));
 sg13g2_nand2b_1 _4387_ (.Y(_0958_),
    .B(_0957_),
    .A_N(_0954_));
 sg13g2_xnor2_1 _4388_ (.Y(_0959_),
    .A(_0954_),
    .B(_0957_));
 sg13g2_xnor2_1 _4389_ (.Y(_0960_),
    .A(_0953_),
    .B(_0959_));
 sg13g2_nor2b_1 _4390_ (.A(_0960_),
    .B_N(_0952_),
    .Y(_0961_));
 sg13g2_xor2_1 _4391_ (.B(_0960_),
    .A(_0952_),
    .X(_0962_));
 sg13g2_inv_1 _4392_ (.Y(_0963_),
    .A(_0962_));
 sg13g2_a21oi_1 _4393_ (.A1(_0931_),
    .A2(_0938_),
    .Y(_0964_),
    .B1(_0937_));
 sg13g2_nand2_1 _4394_ (.Y(_0965_),
    .A(net666),
    .B(net710));
 sg13g2_nand2_1 _4395_ (.Y(_0966_),
    .A(net669),
    .B(net706));
 sg13g2_nand2_1 _4396_ (.Y(_0967_),
    .A(net669),
    .B(net708));
 sg13g2_xor2_1 _4397_ (.B(_0967_),
    .A(_0927_),
    .X(_0968_));
 sg13g2_nand2b_1 _4398_ (.Y(_0969_),
    .B(_0968_),
    .A_N(_0965_));
 sg13g2_xnor2_1 _4399_ (.Y(_0970_),
    .A(_0965_),
    .B(_0968_));
 sg13g2_a21oi_1 _4400_ (.A1(_0932_),
    .A2(_0935_),
    .Y(_0971_),
    .B1(_0934_));
 sg13g2_and2_1 _4401_ (.A(net674),
    .B(net705),
    .X(_0972_));
 sg13g2_nor2_1 _4402_ (.A(net676),
    .B(net651),
    .Y(_0973_));
 sg13g2_nor3_1 _4403_ (.A(net676),
    .B(\core.w[8] ),
    .C(net651),
    .Y(_0974_));
 sg13g2_xnor2_1 _4404_ (.Y(_0975_),
    .A(\core.w[8] ),
    .B(_0973_));
 sg13g2_xor2_1 _4405_ (.B(_0975_),
    .A(_0972_),
    .X(_0976_));
 sg13g2_nor2b_1 _4406_ (.A(_0971_),
    .B_N(_0976_),
    .Y(_0977_));
 sg13g2_xnor2_1 _4407_ (.Y(_0978_),
    .A(_0971_),
    .B(_0976_));
 sg13g2_xnor2_1 _4408_ (.Y(_0979_),
    .A(_0970_),
    .B(_0978_));
 sg13g2_nor2_1 _4409_ (.A(_0964_),
    .B(_0979_),
    .Y(_0980_));
 sg13g2_xor2_1 _4410_ (.B(_0979_),
    .A(_0964_),
    .X(_0981_));
 sg13g2_xnor2_1 _4411_ (.Y(_0982_),
    .A(_0962_),
    .B(_0981_));
 sg13g2_o21ai_1 _4412_ (.B1(_0982_),
    .Y(_0983_),
    .A1(_0940_),
    .A2(_0942_));
 sg13g2_xnor2_1 _4413_ (.Y(_0984_),
    .A(_0951_),
    .B(_0982_));
 sg13g2_nand2b_1 _4414_ (.Y(_0985_),
    .B(_0984_),
    .A_N(_0950_));
 sg13g2_xor2_1 _4415_ (.B(_0984_),
    .A(_0950_),
    .X(_0986_));
 sg13g2_a21o_1 _4416_ (.A2(_0945_),
    .A1(_0913_),
    .B1(_0944_),
    .X(_0987_));
 sg13g2_nor2b_1 _4417_ (.A(_0986_),
    .B_N(_0987_),
    .Y(_0988_));
 sg13g2_xor2_1 _4418_ (.B(_0987_),
    .A(_0986_),
    .X(_0989_));
 sg13g2_nor2_1 _4419_ (.A(_0949_),
    .B(_0989_),
    .Y(_0990_));
 sg13g2_xnor2_1 _4420_ (.Y(_0991_),
    .A(_0910_),
    .B(_0911_));
 sg13g2_nor2_1 _4421_ (.A(\core.w[3] ),
    .B(_0850_),
    .Y(_0992_));
 sg13g2_o21ai_1 _4422_ (.B1(_2726_),
    .Y(_0993_),
    .A1(_0852_),
    .A2(_0854_));
 sg13g2_nand2_1 _4423_ (.Y(_0994_),
    .A(_0855_),
    .B(_0993_));
 sg13g2_nor3_1 _4424_ (.A(\core.w[3] ),
    .B(_0850_),
    .C(_0994_),
    .Y(_0995_));
 sg13g2_xor2_1 _4425_ (.B(_0994_),
    .A(_0992_),
    .X(_0996_));
 sg13g2_nand2_1 _4426_ (.Y(_0997_),
    .A(net675),
    .B(net715));
 sg13g2_nor2_1 _4427_ (.A(_0866_),
    .B(_0997_),
    .Y(_0998_));
 sg13g2_nand2_1 _4428_ (.Y(_0999_),
    .A(net670),
    .B(net718));
 sg13g2_a22oi_1 _4429_ (.Y(_1000_),
    .B1(net715),
    .B2(net674),
    .A2(net713),
    .A1(net675));
 sg13g2_or3_1 _4430_ (.A(_0998_),
    .B(_0999_),
    .C(_1000_),
    .X(_1001_));
 sg13g2_nand2b_1 _4431_ (.Y(_1002_),
    .B(_1001_),
    .A_N(_0998_));
 sg13g2_xnor2_1 _4432_ (.Y(_1003_),
    .A(_0868_),
    .B(_0869_));
 sg13g2_nand2_1 _4433_ (.Y(_1004_),
    .A(_1002_),
    .B(_1003_));
 sg13g2_xnor2_1 _4434_ (.Y(_1005_),
    .A(_1002_),
    .B(_1003_));
 sg13g2_nor2_1 _4435_ (.A(_0996_),
    .B(_1005_),
    .Y(_1006_));
 sg13g2_nor2_1 _4436_ (.A(_0995_),
    .B(_1006_),
    .Y(_1007_));
 sg13g2_xnor2_1 _4437_ (.Y(_1008_),
    .A(_0880_),
    .B(_0881_));
 sg13g2_nor2b_1 _4438_ (.A(_1007_),
    .B_N(_1008_),
    .Y(_1009_));
 sg13g2_xnor2_1 _4439_ (.Y(_1010_),
    .A(_1007_),
    .B(_1008_));
 sg13g2_nor2b_1 _4440_ (.A(_1004_),
    .B_N(_1010_),
    .Y(_1011_));
 sg13g2_nor2_1 _4441_ (.A(_1009_),
    .B(_1011_),
    .Y(_1012_));
 sg13g2_xnor2_1 _4442_ (.Y(_1013_),
    .A(\core.param_a[15] ),
    .B(_0948_));
 sg13g2_or3_1 _4443_ (.A(_0991_),
    .B(_1012_),
    .C(_1013_),
    .X(_1014_));
 sg13g2_xor2_1 _4444_ (.B(_0850_),
    .A(\core.w[3] ),
    .X(_1015_));
 sg13g2_and4_1 _4445_ (.A(net675),
    .B(net678),
    .C(net713),
    .D(net715),
    .X(_1016_));
 sg13g2_nand2_1 _4446_ (.Y(_1017_),
    .A(net674),
    .B(net718));
 sg13g2_a22oi_1 _4447_ (.Y(_1018_),
    .B1(net714),
    .B2(net675),
    .A2(net712),
    .A1(net678));
 sg13g2_or3_1 _4448_ (.A(_1016_),
    .B(_1017_),
    .C(_1018_),
    .X(_1019_));
 sg13g2_nand2b_1 _4449_ (.Y(_1020_),
    .B(_1019_),
    .A_N(_1016_));
 sg13g2_o21ai_1 _4450_ (.B1(_0999_),
    .Y(_1021_),
    .A1(_0998_),
    .A2(_1000_));
 sg13g2_nand3_1 _4451_ (.B(_1020_),
    .C(_1021_),
    .A(_1001_),
    .Y(_1022_));
 sg13g2_a21o_1 _4452_ (.A2(_1021_),
    .A1(_1001_),
    .B1(_1020_),
    .X(_1023_));
 sg13g2_nand3_1 _4453_ (.B(_1022_),
    .C(_1023_),
    .A(_1015_),
    .Y(_1024_));
 sg13g2_xor2_1 _4454_ (.B(_1005_),
    .A(_0996_),
    .X(_1025_));
 sg13g2_nand2b_1 _4455_ (.Y(_1026_),
    .B(_1025_),
    .A_N(_1024_));
 sg13g2_xnor2_1 _4456_ (.Y(_1027_),
    .A(_1024_),
    .B(_1025_));
 sg13g2_nand2b_1 _4457_ (.Y(_1028_),
    .B(_1027_),
    .A_N(_1022_));
 sg13g2_nand2_1 _4458_ (.Y(_1029_),
    .A(_1026_),
    .B(_1028_));
 sg13g2_xor2_1 _4459_ (.B(_1010_),
    .A(_1004_),
    .X(_1030_));
 sg13g2_nor2b_1 _4460_ (.A(_1030_),
    .B_N(_1029_),
    .Y(_1031_));
 sg13g2_xor2_1 _4461_ (.B(_1012_),
    .A(_0991_),
    .X(_1032_));
 sg13g2_and2_1 _4462_ (.A(_1031_),
    .B(_1032_),
    .X(_1033_));
 sg13g2_nor3_1 _4463_ (.A(\core.w[2] ),
    .B(\core.w[1] ),
    .C(\core.w[0] ),
    .Y(_1034_));
 sg13g2_nand2_1 _4464_ (.Y(_1035_),
    .A(net678),
    .B(net717));
 sg13g2_nor2_1 _4465_ (.A(_0997_),
    .B(_1035_),
    .Y(_1036_));
 sg13g2_o21ai_1 _4466_ (.B1(_1017_),
    .Y(_1037_),
    .A1(_1016_),
    .A2(_1018_));
 sg13g2_nand3_1 _4467_ (.B(_1036_),
    .C(_1037_),
    .A(_1019_),
    .Y(_1038_));
 sg13g2_inv_1 _4468_ (.Y(_1039_),
    .A(_1038_));
 sg13g2_a21oi_1 _4469_ (.A1(_1019_),
    .A2(_1037_),
    .Y(_1040_),
    .B1(_1036_));
 sg13g2_nor2_1 _4470_ (.A(_1039_),
    .B(_1040_),
    .Y(_1041_));
 sg13g2_o21ai_1 _4471_ (.B1(\core.w[2] ),
    .Y(_1042_),
    .A1(\core.w[1] ),
    .A2(\core.w[0] ));
 sg13g2_nor2b_1 _4472_ (.A(_1034_),
    .B_N(_1042_),
    .Y(_1043_));
 sg13g2_a21oi_1 _4473_ (.A1(_1041_),
    .A2(_1042_),
    .Y(_1044_),
    .B1(_1034_));
 sg13g2_a21o_1 _4474_ (.A2(_1023_),
    .A1(_1022_),
    .B1(_1015_),
    .X(_1045_));
 sg13g2_nand2_1 _4475_ (.Y(_1046_),
    .A(_1024_),
    .B(_1045_));
 sg13g2_nor2_1 _4476_ (.A(_1044_),
    .B(_1046_),
    .Y(_1047_));
 sg13g2_xor2_1 _4477_ (.B(_1046_),
    .A(_1044_),
    .X(_1048_));
 sg13g2_a21oi_1 _4478_ (.A1(_1039_),
    .A2(_1048_),
    .Y(_1049_),
    .B1(_1047_));
 sg13g2_xnor2_1 _4479_ (.Y(_1050_),
    .A(_1022_),
    .B(_1027_));
 sg13g2_nand2b_1 _4480_ (.Y(_1051_),
    .B(_1050_),
    .A_N(_1049_));
 sg13g2_xor2_1 _4481_ (.B(_1030_),
    .A(_1029_),
    .X(_1052_));
 sg13g2_xor2_1 _4482_ (.B(_1050_),
    .A(_1049_),
    .X(_1053_));
 sg13g2_xnor2_1 _4483_ (.Y(_1054_),
    .A(_1039_),
    .B(_1048_));
 sg13g2_xnor2_1 _4484_ (.Y(_1055_),
    .A(\core.w[1] ),
    .B(\core.w[0] ));
 sg13g2_a22oi_1 _4485_ (.Y(_1056_),
    .B1(net717),
    .B2(net675),
    .A2(net715),
    .A1(net678));
 sg13g2_or3_1 _4486_ (.A(_1036_),
    .B(_1055_),
    .C(_1056_),
    .X(_1057_));
 sg13g2_xnor2_1 _4487_ (.Y(_1058_),
    .A(_1041_),
    .B(_1043_));
 sg13g2_or2_1 _4488_ (.X(_1059_),
    .B(_1058_),
    .A(_1057_));
 sg13g2_or2_1 _4489_ (.X(_1060_),
    .B(_1059_),
    .A(_1054_));
 sg13g2_nor2_1 _4490_ (.A(_1053_),
    .B(_1060_),
    .Y(_1061_));
 sg13g2_o21ai_1 _4491_ (.B1(_1055_),
    .Y(_1062_),
    .A1(_1036_),
    .A2(_1056_));
 sg13g2_nor2_1 _4492_ (.A(_0018_),
    .B(_1035_),
    .Y(_1063_));
 sg13g2_nand3_1 _4493_ (.B(_1062_),
    .C(_1063_),
    .A(_1057_),
    .Y(_1064_));
 sg13g2_xor2_1 _4494_ (.B(_1058_),
    .A(_1057_),
    .X(_1065_));
 sg13g2_nand2b_1 _4495_ (.Y(_1066_),
    .B(_1065_),
    .A_N(_1064_));
 sg13g2_or2_1 _4496_ (.X(_1067_),
    .B(_1066_),
    .A(_1054_));
 sg13g2_inv_1 _4497_ (.Y(_1068_),
    .A(_1067_));
 sg13g2_xor2_1 _4498_ (.B(_1060_),
    .A(_1053_),
    .X(_1069_));
 sg13g2_a21o_1 _4499_ (.A2(_1069_),
    .A1(_1068_),
    .B1(_1061_),
    .X(_1070_));
 sg13g2_xor2_1 _4500_ (.B(_1052_),
    .A(_1051_),
    .X(_1071_));
 sg13g2_nand2_1 _4501_ (.Y(_1072_),
    .A(_1070_),
    .B(_1071_));
 sg13g2_o21ai_1 _4502_ (.B1(_1072_),
    .Y(_1073_),
    .A1(_1051_),
    .A2(_1052_));
 sg13g2_or2_1 _4503_ (.X(_1074_),
    .B(_1032_),
    .A(_1031_));
 sg13g2_nand2b_1 _4504_ (.Y(_1075_),
    .B(_1074_),
    .A_N(_1033_));
 sg13g2_a21oi_1 _4505_ (.A1(_1073_),
    .A2(_1074_),
    .Y(_1076_),
    .B1(_1033_));
 sg13g2_o21ai_1 _4506_ (.B1(_1013_),
    .Y(_1077_),
    .A1(_0991_),
    .A2(_1012_));
 sg13g2_nand2_1 _4507_ (.Y(_1078_),
    .A(_1014_),
    .B(_1077_));
 sg13g2_o21ai_1 _4508_ (.B1(_1014_),
    .Y(_1079_),
    .A1(_1076_),
    .A2(_1078_));
 sg13g2_xor2_1 _4509_ (.B(_0989_),
    .A(_0949_),
    .X(_1080_));
 sg13g2_a21oi_1 _4510_ (.A1(_1079_),
    .A2(_1080_),
    .Y(_1081_),
    .B1(_0990_));
 sg13g2_a21oi_1 _4511_ (.A1(_0953_),
    .A2(_0959_),
    .Y(_1082_),
    .B1(_0961_));
 sg13g2_a21oi_1 _4512_ (.A1(_0963_),
    .A2(_0981_),
    .Y(_1083_),
    .B1(_0980_));
 sg13g2_o21ai_1 _4513_ (.B1(_0958_),
    .Y(_1084_),
    .A1(_0918_),
    .A2(_0956_));
 sg13g2_inv_1 _4514_ (.Y(_1085_),
    .A(_1084_));
 sg13g2_o21ai_1 _4515_ (.B1(_0969_),
    .Y(_1086_),
    .A1(_0927_),
    .A2(_0967_));
 sg13g2_nand2b_1 _4516_ (.Y(_1087_),
    .B(net717),
    .A_N(net659));
 sg13g2_nand2_1 _4517_ (.Y(_1088_),
    .A(net661),
    .B(net712));
 sg13g2_nand2_1 _4518_ (.Y(_1089_),
    .A(net661),
    .B(net714));
 sg13g2_xor2_1 _4519_ (.B(_1089_),
    .A(_0955_),
    .X(_1090_));
 sg13g2_nand2b_1 _4520_ (.Y(_1091_),
    .B(_1090_),
    .A_N(_1087_));
 sg13g2_xnor2_1 _4521_ (.Y(_1092_),
    .A(_1087_),
    .B(_1090_));
 sg13g2_nand2_1 _4522_ (.Y(_1093_),
    .A(_1086_),
    .B(_1092_));
 sg13g2_xnor2_1 _4523_ (.Y(_1094_),
    .A(_1086_),
    .B(_1092_));
 sg13g2_xnor2_1 _4524_ (.Y(_1095_),
    .A(_1085_),
    .B(_1094_));
 sg13g2_inv_1 _4525_ (.Y(_1096_),
    .A(_1095_));
 sg13g2_a21oi_1 _4526_ (.A1(_0970_),
    .A2(_0978_),
    .Y(_1097_),
    .B1(_0977_));
 sg13g2_nand2_1 _4527_ (.Y(_1098_),
    .A(net664),
    .B(net710));
 sg13g2_nand2_1 _4528_ (.Y(_1099_),
    .A(net666),
    .B(net706));
 sg13g2_nand2_1 _4529_ (.Y(_1100_),
    .A(net666),
    .B(net708));
 sg13g2_xor2_1 _4530_ (.B(_1100_),
    .A(_0966_),
    .X(_1101_));
 sg13g2_nand2b_1 _4531_ (.Y(_1102_),
    .B(_1101_),
    .A_N(_1098_));
 sg13g2_xnor2_1 _4532_ (.Y(_1103_),
    .A(_1098_),
    .B(_1101_));
 sg13g2_a21oi_1 _4533_ (.A1(_0972_),
    .A2(_0975_),
    .Y(_1104_),
    .B1(_0974_));
 sg13g2_and2_1 _4534_ (.A(net670),
    .B(net705),
    .X(_1105_));
 sg13g2_nor2_1 _4535_ (.A(net673),
    .B(net651),
    .Y(_1106_));
 sg13g2_nor3_1 _4536_ (.A(net673),
    .B(\core.w[9] ),
    .C(net651),
    .Y(_1107_));
 sg13g2_xnor2_1 _4537_ (.Y(_1108_),
    .A(\core.w[9] ),
    .B(_1106_));
 sg13g2_xor2_1 _4538_ (.B(_1108_),
    .A(_1105_),
    .X(_1109_));
 sg13g2_nor2b_1 _4539_ (.A(_1104_),
    .B_N(_1109_),
    .Y(_1110_));
 sg13g2_xnor2_1 _4540_ (.Y(_1111_),
    .A(_1104_),
    .B(_1109_));
 sg13g2_xnor2_1 _4541_ (.Y(_1112_),
    .A(_1103_),
    .B(_1111_));
 sg13g2_nor2_1 _4542_ (.A(_1097_),
    .B(_1112_),
    .Y(_1113_));
 sg13g2_xor2_1 _4543_ (.B(_1112_),
    .A(_1097_),
    .X(_1114_));
 sg13g2_xnor2_1 _4544_ (.Y(_1115_),
    .A(_1095_),
    .B(_1114_));
 sg13g2_nand2b_1 _4545_ (.Y(_1116_),
    .B(_1115_),
    .A_N(_1083_));
 sg13g2_xnor2_1 _4546_ (.Y(_1117_),
    .A(_1083_),
    .B(_1115_));
 sg13g2_nand2b_1 _4547_ (.Y(_1118_),
    .B(_1117_),
    .A_N(_1082_));
 sg13g2_xor2_1 _4548_ (.B(_1117_),
    .A(_1082_),
    .X(_1119_));
 sg13g2_a21oi_2 _4549_ (.B1(_1119_),
    .Y(_1120_),
    .A2(_0985_),
    .A1(_0983_));
 sg13g2_nand3_1 _4550_ (.B(_0985_),
    .C(_1119_),
    .A(_0983_),
    .Y(_1121_));
 sg13g2_nor2b_1 _4551_ (.A(_1120_),
    .B_N(_1121_),
    .Y(_1122_));
 sg13g2_nand2_1 _4552_ (.Y(_1123_),
    .A(_0988_),
    .B(_1122_));
 sg13g2_xnor2_1 _4553_ (.Y(_1124_),
    .A(_0988_),
    .B(_1122_));
 sg13g2_xor2_1 _4554_ (.B(_1124_),
    .A(_1081_),
    .X(_1125_));
 sg13g2_xnor2_1 _4555_ (.Y(_1126_),
    .A(_1079_),
    .B(_1080_));
 sg13g2_nor2_1 _4556_ (.A(net575),
    .B(_1125_),
    .Y(_1127_));
 sg13g2_a21oi_1 _4557_ (.A1(net576),
    .A2(_1126_),
    .Y(_1128_),
    .B1(_1127_));
 sg13g2_o21ai_1 _4558_ (.B1(_1123_),
    .Y(_1129_),
    .A1(_1081_),
    .A2(_1124_));
 sg13g2_o21ai_1 _4559_ (.B1(_1093_),
    .Y(_1130_),
    .A1(_1085_),
    .A2(_1094_));
 sg13g2_a21oi_1 _4560_ (.A1(_1096_),
    .A2(_1114_),
    .Y(_1131_),
    .B1(_1113_));
 sg13g2_a21oi_1 _4561_ (.A1(_1103_),
    .A2(_1111_),
    .Y(_1132_),
    .B1(_1110_));
 sg13g2_nand2_1 _4562_ (.Y(_1133_),
    .A(net662),
    .B(net710));
 sg13g2_nand2_1 _4563_ (.Y(_1134_),
    .A(net664),
    .B(net707));
 sg13g2_nand2_1 _4564_ (.Y(_1135_),
    .A(net664),
    .B(net708));
 sg13g2_xor2_1 _4565_ (.B(_1135_),
    .A(_1099_),
    .X(_1136_));
 sg13g2_nand2b_1 _4566_ (.Y(_1137_),
    .B(_1136_),
    .A_N(_1133_));
 sg13g2_xnor2_1 _4567_ (.Y(_1138_),
    .A(_1133_),
    .B(_1136_));
 sg13g2_a21oi_1 _4568_ (.A1(_1105_),
    .A2(_1108_),
    .Y(_1139_),
    .B1(_1107_));
 sg13g2_and2_1 _4569_ (.A(net668),
    .B(net705),
    .X(_1140_));
 sg13g2_nor2_1 _4570_ (.A(net671),
    .B(net651),
    .Y(_1141_));
 sg13g2_nor3_1 _4571_ (.A(net670),
    .B(\core.w[10] ),
    .C(net651),
    .Y(_1142_));
 sg13g2_xnor2_1 _4572_ (.Y(_1143_),
    .A(\core.w[10] ),
    .B(_1141_));
 sg13g2_xor2_1 _4573_ (.B(_1143_),
    .A(_1140_),
    .X(_1144_));
 sg13g2_nor2b_1 _4574_ (.A(_1139_),
    .B_N(_1144_),
    .Y(_1145_));
 sg13g2_xnor2_1 _4575_ (.Y(_1146_),
    .A(_1139_),
    .B(_1144_));
 sg13g2_xnor2_1 _4576_ (.Y(_1147_),
    .A(_1138_),
    .B(_1146_));
 sg13g2_nor2_1 _4577_ (.A(_1132_),
    .B(_1147_),
    .Y(_1148_));
 sg13g2_xor2_1 _4578_ (.B(_1147_),
    .A(_1132_),
    .X(_1149_));
 sg13g2_o21ai_1 _4579_ (.B1(_1091_),
    .Y(_1150_),
    .A1(_0955_),
    .A2(_1089_));
 sg13g2_inv_1 _4580_ (.Y(_1151_),
    .A(_1150_));
 sg13g2_o21ai_1 _4581_ (.B1(_1102_),
    .Y(_1152_),
    .A1(_0966_),
    .A2(_1100_));
 sg13g2_nor2_1 _4582_ (.A(net656),
    .B(net657),
    .Y(_1153_));
 sg13g2_xnor2_1 _4583_ (.Y(_1154_),
    .A(net656),
    .B(net658));
 sg13g2_nand2_1 _4584_ (.Y(_1155_),
    .A(net718),
    .B(_1154_));
 sg13g2_nand2b_1 _4585_ (.Y(_1156_),
    .B(net713),
    .A_N(net659));
 sg13g2_nand2b_1 _4586_ (.Y(_1157_),
    .B(net714),
    .A_N(net659));
 sg13g2_xor2_1 _4587_ (.B(_1157_),
    .A(_1088_),
    .X(_1158_));
 sg13g2_nand2b_1 _4588_ (.Y(_1159_),
    .B(_1158_),
    .A_N(_1155_));
 sg13g2_xnor2_1 _4589_ (.Y(_1160_),
    .A(_1155_),
    .B(_1158_));
 sg13g2_nand2_1 _4590_ (.Y(_1161_),
    .A(_1152_),
    .B(_1160_));
 sg13g2_xnor2_1 _4591_ (.Y(_1162_),
    .A(_1152_),
    .B(_1160_));
 sg13g2_xnor2_1 _4592_ (.Y(_1163_),
    .A(_1151_),
    .B(_1162_));
 sg13g2_inv_1 _4593_ (.Y(_1164_),
    .A(_1163_));
 sg13g2_xnor2_1 _4594_ (.Y(_1165_),
    .A(_1149_),
    .B(_1164_));
 sg13g2_nor2_1 _4595_ (.A(_1131_),
    .B(_1165_),
    .Y(_1166_));
 sg13g2_xor2_1 _4596_ (.B(_1165_),
    .A(_1131_),
    .X(_1167_));
 sg13g2_xnor2_1 _4597_ (.Y(_1168_),
    .A(_1130_),
    .B(_1167_));
 sg13g2_a21oi_2 _4598_ (.B1(_1168_),
    .Y(_1169_),
    .A2(_1118_),
    .A1(_1116_));
 sg13g2_nand3_1 _4599_ (.B(_1118_),
    .C(_1168_),
    .A(_1116_),
    .Y(_1170_));
 sg13g2_nor2b_1 _4600_ (.A(_1169_),
    .B_N(_1170_),
    .Y(_1171_));
 sg13g2_and2_1 _4601_ (.A(_1120_),
    .B(_1171_),
    .X(_1172_));
 sg13g2_xor2_1 _4602_ (.B(_1171_),
    .A(_1120_),
    .X(_1173_));
 sg13g2_xnor2_1 _4603_ (.Y(_1174_),
    .A(_1129_),
    .B(_1173_));
 sg13g2_a21o_1 _4604_ (.A2(_1173_),
    .A1(_1129_),
    .B1(_1172_),
    .X(_1175_));
 sg13g2_o21ai_1 _4605_ (.B1(_1161_),
    .Y(_1176_),
    .A1(_1151_),
    .A2(_1162_));
 sg13g2_a21oi_1 _4606_ (.A1(_1149_),
    .A2(_1164_),
    .Y(_1177_),
    .B1(_1148_));
 sg13g2_o21ai_1 _4607_ (.B1(_1159_),
    .Y(_1178_),
    .A1(_1088_),
    .A2(_1157_));
 sg13g2_inv_1 _4608_ (.Y(_1179_),
    .A(_1178_));
 sg13g2_o21ai_1 _4609_ (.B1(_1137_),
    .Y(_1180_),
    .A1(_1099_),
    .A2(_1135_));
 sg13g2_nor2b_1 _4610_ (.A(_1153_),
    .B_N(net655),
    .Y(_1181_));
 sg13g2_xnor2_1 _4611_ (.Y(_1182_),
    .A(net655),
    .B(_1153_));
 sg13g2_nand2_2 _4612_ (.Y(_1183_),
    .A(\core.param_a[8] ),
    .B(_1182_));
 sg13g2_nand2_1 _4613_ (.Y(_1184_),
    .A(\core.param_a[10] ),
    .B(_1154_));
 sg13g2_nand2_1 _4614_ (.Y(_1185_),
    .A(net715),
    .B(_1154_));
 sg13g2_xor2_1 _4615_ (.B(_1185_),
    .A(_1156_),
    .X(_1186_));
 sg13g2_nand2b_1 _4616_ (.Y(_1187_),
    .B(_1186_),
    .A_N(_1183_));
 sg13g2_xnor2_1 _4617_ (.Y(_1188_),
    .A(_1183_),
    .B(_1186_));
 sg13g2_nand2_1 _4618_ (.Y(_1189_),
    .A(_1180_),
    .B(_1188_));
 sg13g2_xnor2_1 _4619_ (.Y(_1190_),
    .A(_1180_),
    .B(_1188_));
 sg13g2_xnor2_1 _4620_ (.Y(_1191_),
    .A(_1179_),
    .B(_1190_));
 sg13g2_inv_1 _4621_ (.Y(_1192_),
    .A(_1191_));
 sg13g2_a21oi_1 _4622_ (.A1(_1138_),
    .A2(_1146_),
    .Y(_1193_),
    .B1(_1145_));
 sg13g2_nand2_1 _4623_ (.Y(_1194_),
    .A(net661),
    .B(net711));
 sg13g2_nand2_1 _4624_ (.Y(_1195_),
    .A(net663),
    .B(net707));
 sg13g2_nand2_1 _4625_ (.Y(_1196_),
    .A(net662),
    .B(net708));
 sg13g2_xor2_1 _4626_ (.B(_1196_),
    .A(_1134_),
    .X(_1197_));
 sg13g2_nand2b_1 _4627_ (.Y(_1198_),
    .B(_1197_),
    .A_N(_1194_));
 sg13g2_xnor2_1 _4628_ (.Y(_1199_),
    .A(_1194_),
    .B(_1197_));
 sg13g2_a21oi_2 _4629_ (.B1(_1142_),
    .Y(_1200_),
    .A2(_1143_),
    .A1(_1140_));
 sg13g2_and2_1 _4630_ (.A(net666),
    .B(net705),
    .X(_1201_));
 sg13g2_nor2_1 _4631_ (.A(\core.V[4] ),
    .B(net652),
    .Y(_1202_));
 sg13g2_nor3_1 _4632_ (.A(net669),
    .B(\core.w[11] ),
    .C(net652),
    .Y(_1203_));
 sg13g2_xnor2_1 _4633_ (.Y(_1204_),
    .A(\core.w[11] ),
    .B(_1202_));
 sg13g2_xor2_1 _4634_ (.B(_1204_),
    .A(_1201_),
    .X(_1205_));
 sg13g2_nor2b_1 _4635_ (.A(_1200_),
    .B_N(_1205_),
    .Y(_1206_));
 sg13g2_xnor2_1 _4636_ (.Y(_1207_),
    .A(_1200_),
    .B(_1205_));
 sg13g2_xnor2_1 _4637_ (.Y(_1208_),
    .A(_1199_),
    .B(_1207_));
 sg13g2_nor2_1 _4638_ (.A(_1193_),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_xor2_1 _4639_ (.B(_1208_),
    .A(_1193_),
    .X(_1210_));
 sg13g2_xnor2_1 _4640_ (.Y(_1211_),
    .A(_1191_),
    .B(_1210_));
 sg13g2_nor2b_1 _4641_ (.A(_1177_),
    .B_N(_1211_),
    .Y(_1212_));
 sg13g2_xnor2_1 _4642_ (.Y(_1213_),
    .A(_1177_),
    .B(_1211_));
 sg13g2_xnor2_1 _4643_ (.Y(_1214_),
    .A(_1176_),
    .B(_1213_));
 sg13g2_a21oi_2 _4644_ (.B1(_1166_),
    .Y(_1215_),
    .A2(_1167_),
    .A1(_1130_));
 sg13g2_nor2_2 _4645_ (.A(_1214_),
    .B(_1215_),
    .Y(_1216_));
 sg13g2_inv_1 _4646_ (.Y(_1217_),
    .A(_1216_));
 sg13g2_xor2_1 _4647_ (.B(_1215_),
    .A(_1214_),
    .X(_1218_));
 sg13g2_and2_1 _4648_ (.A(_1169_),
    .B(_1218_),
    .X(_1219_));
 sg13g2_xnor2_1 _4649_ (.Y(_1220_),
    .A(_1169_),
    .B(_1218_));
 sg13g2_inv_1 _4650_ (.Y(_1221_),
    .A(_1220_));
 sg13g2_xnor2_1 _4651_ (.Y(_1222_),
    .A(_1175_),
    .B(_1220_));
 sg13g2_nor2_1 _4652_ (.A(net574),
    .B(_1222_),
    .Y(_1223_));
 sg13g2_a21oi_1 _4653_ (.A1(net576),
    .A2(_1174_),
    .Y(_1224_),
    .B1(_1223_));
 sg13g2_mux2_2 _4654_ (.A0(_1128_),
    .A1(_1224_),
    .S(net582),
    .X(_1225_));
 sg13g2_a21oi_2 _4655_ (.B1(_0842_),
    .Y(_1226_),
    .A2(_0831_),
    .A1(_0825_));
 sg13g2_inv_1 _4656_ (.Y(_1227_),
    .A(_1226_));
 sg13g2_nor2_2 _4657_ (.A(_0842_),
    .B(net586),
    .Y(_1228_));
 sg13g2_nand2_2 _4658_ (.Y(_1229_),
    .A(_0841_),
    .B(_1227_));
 sg13g2_nand2_1 _4659_ (.Y(_1230_),
    .A(_1059_),
    .B(_1066_));
 sg13g2_xnor2_1 _4660_ (.Y(_1231_),
    .A(_1054_),
    .B(_1230_));
 sg13g2_xnor2_1 _4661_ (.Y(_1232_),
    .A(_1064_),
    .B(_1065_));
 sg13g2_mux2_1 _4662_ (.A0(_1231_),
    .A1(_1232_),
    .S(net575),
    .X(_1233_));
 sg13g2_o21ai_1 _4663_ (.B1(_1228_),
    .Y(_1234_),
    .A1(net577),
    .A2(_1233_));
 sg13g2_xnor2_1 _4664_ (.Y(_1235_),
    .A(_1067_),
    .B(_1069_));
 sg13g2_xor2_1 _4665_ (.B(_1071_),
    .A(_1070_),
    .X(_1236_));
 sg13g2_mux2_1 _4666_ (.A0(_1236_),
    .A1(_1235_),
    .S(net574),
    .X(_1237_));
 sg13g2_nor2_1 _4667_ (.A(net582),
    .B(_1237_),
    .Y(_1238_));
 sg13g2_xnor2_1 _4668_ (.Y(_1239_),
    .A(_1076_),
    .B(_1078_));
 sg13g2_xor2_1 _4669_ (.B(_1075_),
    .A(_1073_),
    .X(_1240_));
 sg13g2_mux2_1 _4670_ (.A0(_1239_),
    .A1(_1240_),
    .S(net574),
    .X(_1241_));
 sg13g2_a21oi_2 _4671_ (.B1(_1238_),
    .Y(_1242_),
    .A2(_1241_),
    .A1(net582));
 sg13g2_a22oi_1 _4672_ (.Y(_1243_),
    .B1(net586),
    .B2(_1242_),
    .A2(_1225_),
    .A1(_0842_));
 sg13g2_nand2_1 _4673_ (.Y(_1244_),
    .A(_1234_),
    .B(_1243_));
 sg13g2_a22oi_1 _4674_ (.Y(_1245_),
    .B1(_0836_),
    .B2(_1244_),
    .A2(net638),
    .A1(net549));
 sg13g2_nor2_1 _4675_ (.A(net725),
    .B(_1245_),
    .Y(_0202_));
 sg13g2_a21o_2 _4676_ (.A2(_1221_),
    .A1(_1175_),
    .B1(_1219_),
    .X(_1246_));
 sg13g2_o21ai_1 _4677_ (.B1(_1189_),
    .Y(_1247_),
    .A1(_1179_),
    .A2(_1190_));
 sg13g2_a21oi_1 _4678_ (.A1(_1192_),
    .A2(_1210_),
    .Y(_1248_),
    .B1(_1209_));
 sg13g2_a21oi_1 _4679_ (.A1(_1199_),
    .A2(_1207_),
    .Y(_1249_),
    .B1(_1206_));
 sg13g2_nor2b_1 _4680_ (.A(net659),
    .B_N(net711),
    .Y(_1250_));
 sg13g2_nand2_1 _4681_ (.Y(_1251_),
    .A(net660),
    .B(net709));
 sg13g2_xor2_1 _4682_ (.B(_1251_),
    .A(_1195_),
    .X(_1252_));
 sg13g2_nand2_1 _4683_ (.Y(_1253_),
    .A(_1250_),
    .B(_1252_));
 sg13g2_xnor2_1 _4684_ (.Y(_1254_),
    .A(_1250_),
    .B(_1252_));
 sg13g2_a21oi_1 _4685_ (.A1(_1201_),
    .A2(_1204_),
    .Y(_1255_),
    .B1(_1203_));
 sg13g2_inv_1 _4686_ (.Y(_1256_),
    .A(_1255_));
 sg13g2_and2_1 _4687_ (.A(net665),
    .B(\core.param_a[14] ),
    .X(_1257_));
 sg13g2_nor2_1 _4688_ (.A(net667),
    .B(net652),
    .Y(_1258_));
 sg13g2_nor3_1 _4689_ (.A(net667),
    .B(\core.w[12] ),
    .C(net652),
    .Y(_1259_));
 sg13g2_xnor2_1 _4690_ (.Y(_1260_),
    .A(\core.w[12] ),
    .B(_1258_));
 sg13g2_xor2_1 _4691_ (.B(_1260_),
    .A(_1257_),
    .X(_1261_));
 sg13g2_xnor2_1 _4692_ (.Y(_1262_),
    .A(_1255_),
    .B(_1261_));
 sg13g2_nor2b_1 _4693_ (.A(_1254_),
    .B_N(_1262_),
    .Y(_1263_));
 sg13g2_xnor2_1 _4694_ (.Y(_1264_),
    .A(_1254_),
    .B(_1262_));
 sg13g2_nand2b_1 _4695_ (.Y(_1265_),
    .B(_1264_),
    .A_N(_1249_));
 sg13g2_xnor2_1 _4696_ (.Y(_1266_),
    .A(_1249_),
    .B(_1264_));
 sg13g2_inv_1 _4697_ (.Y(_1267_),
    .A(_1266_));
 sg13g2_o21ai_1 _4698_ (.B1(_1187_),
    .Y(_1268_),
    .A1(_1156_),
    .A2(_1185_));
 sg13g2_o21ai_1 _4699_ (.B1(_1198_),
    .Y(_1269_),
    .A1(_1134_),
    .A2(_1196_));
 sg13g2_xnor2_1 _4700_ (.Y(_1270_),
    .A(_0021_),
    .B(_1181_));
 sg13g2_nand2_1 _4701_ (.Y(_1271_),
    .A(\core.param_a[8] ),
    .B(_1270_));
 sg13g2_nand2_1 _4702_ (.Y(_1272_),
    .A(net713),
    .B(_1182_));
 sg13g2_nand2_1 _4703_ (.Y(_1273_),
    .A(net716),
    .B(_1182_));
 sg13g2_xor2_1 _4704_ (.B(_1273_),
    .A(_1184_),
    .X(_1274_));
 sg13g2_nand2b_1 _4705_ (.Y(_1275_),
    .B(_1274_),
    .A_N(_1271_));
 sg13g2_xnor2_1 _4706_ (.Y(_1276_),
    .A(_1271_),
    .B(_1274_));
 sg13g2_and2_1 _4707_ (.A(_1269_),
    .B(_1276_),
    .X(_1277_));
 sg13g2_xor2_1 _4708_ (.B(_1276_),
    .A(_1269_),
    .X(_1278_));
 sg13g2_xnor2_1 _4709_ (.Y(_1279_),
    .A(_1268_),
    .B(_1278_));
 sg13g2_xor2_1 _4710_ (.B(_1279_),
    .A(_1266_),
    .X(_1280_));
 sg13g2_nor2_1 _4711_ (.A(_1248_),
    .B(_1280_),
    .Y(_1281_));
 sg13g2_xor2_1 _4712_ (.B(_1280_),
    .A(_1248_),
    .X(_1282_));
 sg13g2_xnor2_1 _4713_ (.Y(_1283_),
    .A(_1247_),
    .B(_1282_));
 sg13g2_a21oi_2 _4714_ (.B1(_1212_),
    .Y(_1284_),
    .A2(_1213_),
    .A1(_1176_));
 sg13g2_nor2_1 _4715_ (.A(_1283_),
    .B(_1284_),
    .Y(_1285_));
 sg13g2_inv_1 _4716_ (.Y(_1286_),
    .A(_1285_));
 sg13g2_xnor2_1 _4717_ (.Y(_1287_),
    .A(_1283_),
    .B(_1284_));
 sg13g2_xor2_1 _4718_ (.B(_1287_),
    .A(_1216_),
    .X(_1288_));
 sg13g2_nand2b_1 _4719_ (.Y(_1289_),
    .B(_1246_),
    .A_N(_1288_));
 sg13g2_xor2_1 _4720_ (.B(_1288_),
    .A(_1246_),
    .X(_1290_));
 sg13g2_nand2_1 _4721_ (.Y(_1291_),
    .A(net574),
    .B(_1222_));
 sg13g2_o21ai_1 _4722_ (.B1(_1291_),
    .Y(_1292_),
    .A1(net576),
    .A2(_1290_));
 sg13g2_nand2_1 _4723_ (.Y(_1293_),
    .A(net574),
    .B(_1125_));
 sg13g2_o21ai_1 _4724_ (.B1(_1293_),
    .Y(_1294_),
    .A1(net576),
    .A2(_1174_));
 sg13g2_mux2_1 _4725_ (.A0(_1292_),
    .A1(_1294_),
    .S(net577),
    .X(_1295_));
 sg13g2_nand2_1 _4726_ (.Y(_1296_),
    .A(_0842_),
    .B(_1295_));
 sg13g2_mux2_1 _4727_ (.A0(_1235_),
    .A1(_1231_),
    .S(net575),
    .X(_1297_));
 sg13g2_o21ai_1 _4728_ (.B1(_1228_),
    .Y(_1298_),
    .A1(net577),
    .A2(_1297_));
 sg13g2_nor2_1 _4729_ (.A(net574),
    .B(_1240_),
    .Y(_1299_));
 sg13g2_a21oi_2 _4730_ (.B1(_1299_),
    .Y(_1300_),
    .A2(_1236_),
    .A1(net574));
 sg13g2_nand2_1 _4731_ (.Y(_1301_),
    .A(net578),
    .B(_1300_));
 sg13g2_mux2_1 _4732_ (.A0(_1126_),
    .A1(_1239_),
    .S(net574),
    .X(_1302_));
 sg13g2_nand2_1 _4733_ (.Y(_1303_),
    .A(net582),
    .B(_1302_));
 sg13g2_nand3_1 _4734_ (.B(_1301_),
    .C(_1303_),
    .A(net586),
    .Y(_1304_));
 sg13g2_nand3_1 _4735_ (.B(_1298_),
    .C(_1304_),
    .A(_1296_),
    .Y(_1305_));
 sg13g2_a22oi_1 _4736_ (.Y(_1306_),
    .B1(_0836_),
    .B2(_1305_),
    .A2(net638),
    .A1(net780));
 sg13g2_nor2_1 _4737_ (.A(net724),
    .B(_1306_),
    .Y(_0203_));
 sg13g2_o21ai_1 _4738_ (.B1(_1289_),
    .Y(_1307_),
    .A1(_1217_),
    .A2(_1287_));
 sg13g2_a21oi_1 _4739_ (.A1(_1268_),
    .A2(_1278_),
    .Y(_1308_),
    .B1(_1277_));
 sg13g2_o21ai_1 _4740_ (.B1(_1265_),
    .Y(_1309_),
    .A1(_1267_),
    .A2(_1279_));
 sg13g2_o21ai_1 _4741_ (.B1(_1275_),
    .Y(_1310_),
    .A1(_1184_),
    .A2(_1273_));
 sg13g2_inv_1 _4742_ (.Y(_1311_),
    .A(_1310_));
 sg13g2_o21ai_1 _4743_ (.B1(_1253_),
    .Y(_1312_),
    .A1(_1195_),
    .A2(_1251_));
 sg13g2_and3_1 _4744_ (.X(_1313_),
    .A(net653),
    .B(net654),
    .C(_1181_));
 sg13g2_a21oi_1 _4745_ (.A1(net654),
    .A2(_1181_),
    .Y(_1314_),
    .B1(net653));
 sg13g2_nor2_1 _4746_ (.A(_1313_),
    .B(_1314_),
    .Y(_1315_));
 sg13g2_nand2_1 _4747_ (.Y(_1316_),
    .A(net718),
    .B(_1315_));
 sg13g2_nand2_1 _4748_ (.Y(_1317_),
    .A(net713),
    .B(_1270_));
 sg13g2_nand2_1 _4749_ (.Y(_1318_),
    .A(net716),
    .B(_1270_));
 sg13g2_xor2_1 _4750_ (.B(_1318_),
    .A(_1272_),
    .X(_1319_));
 sg13g2_nand2b_1 _4751_ (.Y(_1320_),
    .B(_1319_),
    .A_N(_1316_));
 sg13g2_xnor2_1 _4752_ (.Y(_1321_),
    .A(_1316_),
    .B(_1319_));
 sg13g2_nand2_1 _4753_ (.Y(_1322_),
    .A(_1312_),
    .B(_1321_));
 sg13g2_xnor2_1 _4754_ (.Y(_1323_),
    .A(_1312_),
    .B(_1321_));
 sg13g2_xnor2_1 _4755_ (.Y(_1324_),
    .A(_1310_),
    .B(_1323_));
 sg13g2_a21oi_1 _4756_ (.A1(_1256_),
    .A2(_1261_),
    .Y(_1325_),
    .B1(_1263_));
 sg13g2_nand2_1 _4757_ (.Y(_1326_),
    .A(net711),
    .B(_1154_));
 sg13g2_nor2b_1 _4758_ (.A(net658),
    .B_N(net707),
    .Y(_1327_));
 sg13g2_nor2b_1 _4759_ (.A(net658),
    .B_N(net709),
    .Y(_1328_));
 sg13g2_nand2b_1 _4760_ (.Y(_1329_),
    .B(_1327_),
    .A_N(_1251_));
 sg13g2_a21o_1 _4761_ (.A2(net707),
    .A1(net660),
    .B1(_1328_),
    .X(_1330_));
 sg13g2_and2_1 _4762_ (.A(_1329_),
    .B(_1330_),
    .X(_1331_));
 sg13g2_nand2b_1 _4763_ (.Y(_1332_),
    .B(_1331_),
    .A_N(_1326_));
 sg13g2_xnor2_1 _4764_ (.Y(_1333_),
    .A(_1326_),
    .B(_1331_));
 sg13g2_a21oi_1 _4765_ (.A1(_1257_),
    .A2(_1260_),
    .Y(_1334_),
    .B1(_1259_));
 sg13g2_and2_1 _4766_ (.A(net663),
    .B(net705),
    .X(_1335_));
 sg13g2_nor2_1 _4767_ (.A(net665),
    .B(net652),
    .Y(_1336_));
 sg13g2_nor3_1 _4768_ (.A(net665),
    .B(\core.w[13] ),
    .C(net652),
    .Y(_1337_));
 sg13g2_xnor2_1 _4769_ (.Y(_1338_),
    .A(\core.w[13] ),
    .B(_1336_));
 sg13g2_xnor2_1 _4770_ (.Y(_1339_),
    .A(_1335_),
    .B(_1338_));
 sg13g2_nor2_1 _4771_ (.A(_1334_),
    .B(_1339_),
    .Y(_1340_));
 sg13g2_xor2_1 _4772_ (.B(_1339_),
    .A(_1334_),
    .X(_1341_));
 sg13g2_xnor2_1 _4773_ (.Y(_1342_),
    .A(_1333_),
    .B(_1341_));
 sg13g2_nor2_1 _4774_ (.A(_1325_),
    .B(_1342_),
    .Y(_1343_));
 sg13g2_xor2_1 _4775_ (.B(_1342_),
    .A(_1325_),
    .X(_1344_));
 sg13g2_xor2_1 _4776_ (.B(_1344_),
    .A(_1324_),
    .X(_1345_));
 sg13g2_nand2_1 _4777_ (.Y(_1346_),
    .A(_1309_),
    .B(_1345_));
 sg13g2_xnor2_1 _4778_ (.Y(_1347_),
    .A(_1309_),
    .B(_1345_));
 sg13g2_xnor2_1 _4779_ (.Y(_1348_),
    .A(_1308_),
    .B(_1347_));
 sg13g2_a21oi_2 _4780_ (.B1(_1281_),
    .Y(_1349_),
    .A2(_1282_),
    .A1(_1247_));
 sg13g2_xnor2_1 _4781_ (.Y(_1350_),
    .A(_1348_),
    .B(_1349_));
 sg13g2_nor2_1 _4782_ (.A(_1286_),
    .B(_1350_),
    .Y(_1351_));
 sg13g2_xnor2_1 _4783_ (.Y(_1352_),
    .A(_1286_),
    .B(_1350_));
 sg13g2_inv_1 _4784_ (.Y(_1353_),
    .A(_1352_));
 sg13g2_xnor2_1 _4785_ (.Y(_1354_),
    .A(_1307_),
    .B(_1353_));
 sg13g2_mux2_1 _4786_ (.A0(_1354_),
    .A1(_1290_),
    .S(net576),
    .X(_1355_));
 sg13g2_nand2_1 _4787_ (.Y(_1356_),
    .A(net577),
    .B(_1224_));
 sg13g2_o21ai_1 _4788_ (.B1(_1356_),
    .Y(_1357_),
    .A1(net578),
    .A2(_1355_));
 sg13g2_o21ai_1 _4789_ (.B1(_1228_),
    .Y(_1358_),
    .A1(net577),
    .A2(_1237_));
 sg13g2_nor2_1 _4790_ (.A(net577),
    .B(_1128_),
    .Y(_1359_));
 sg13g2_a21oi_2 _4791_ (.B1(_1359_),
    .Y(_1360_),
    .A2(_1241_),
    .A1(net577));
 sg13g2_a22oi_1 _4792_ (.Y(_1361_),
    .B1(_1360_),
    .B2(net586),
    .A2(_1357_),
    .A1(_0842_));
 sg13g2_nand2_1 _4793_ (.Y(_1362_),
    .A(_1358_),
    .B(_1361_));
 sg13g2_a22oi_1 _4794_ (.Y(_1363_),
    .B1(_0836_),
    .B2(_1362_),
    .A2(net638),
    .A1(net760));
 sg13g2_nor2_1 _4795_ (.A(net725),
    .B(_1363_),
    .Y(_0204_));
 sg13g2_a21o_1 _4796_ (.A2(_1353_),
    .A1(_1307_),
    .B1(_1351_),
    .X(_1364_));
 sg13g2_o21ai_1 _4797_ (.B1(_1346_),
    .Y(_1365_),
    .A1(_1308_),
    .A2(_1347_));
 sg13g2_o21ai_1 _4798_ (.B1(_1322_),
    .Y(_1366_),
    .A1(_1311_),
    .A2(_1323_));
 sg13g2_a21oi_1 _4799_ (.A1(_1324_),
    .A2(_1344_),
    .Y(_1367_),
    .B1(_1343_));
 sg13g2_a21oi_1 _4800_ (.A1(_1333_),
    .A2(_1341_),
    .Y(_1368_),
    .B1(_1340_));
 sg13g2_nand2_1 _4801_ (.Y(_1369_),
    .A(net711),
    .B(_1182_));
 sg13g2_nand2_1 _4802_ (.Y(_1370_),
    .A(net707),
    .B(_1154_));
 sg13g2_nand3_1 _4803_ (.B(_1154_),
    .C(_1328_),
    .A(net707),
    .Y(_1371_));
 sg13g2_a21o_1 _4804_ (.A2(_1154_),
    .A1(net709),
    .B1(_1327_),
    .X(_1372_));
 sg13g2_and2_1 _4805_ (.A(_1371_),
    .B(_1372_),
    .X(_1373_));
 sg13g2_nand2b_1 _4806_ (.Y(_1374_),
    .B(_1373_),
    .A_N(_1369_));
 sg13g2_xnor2_1 _4807_ (.Y(_1375_),
    .A(_1369_),
    .B(_1373_));
 sg13g2_a21oi_2 _4808_ (.B1(_1337_),
    .Y(_1376_),
    .A2(_1338_),
    .A1(_1335_));
 sg13g2_nand2_1 _4809_ (.Y(_1377_),
    .A(net660),
    .B(\core.param_a[14] ));
 sg13g2_nand2b_1 _4810_ (.Y(_1378_),
    .B(\core.param_a[15] ),
    .A_N(net663));
 sg13g2_xor2_1 _4811_ (.B(_1378_),
    .A(\core.w[14] ),
    .X(_1379_));
 sg13g2_nand2b_1 _4812_ (.Y(_1380_),
    .B(_1379_),
    .A_N(_1377_));
 sg13g2_xor2_1 _4813_ (.B(_1379_),
    .A(_1377_),
    .X(_1381_));
 sg13g2_nor2_1 _4814_ (.A(_1376_),
    .B(_1381_),
    .Y(_1382_));
 sg13g2_xor2_1 _4815_ (.B(_1381_),
    .A(_1376_),
    .X(_1383_));
 sg13g2_xnor2_1 _4816_ (.Y(_1384_),
    .A(_1375_),
    .B(_1383_));
 sg13g2_or2_1 _4817_ (.X(_1385_),
    .B(_1384_),
    .A(_1368_));
 sg13g2_xnor2_1 _4818_ (.Y(_1386_),
    .A(_1368_),
    .B(_1384_));
 sg13g2_o21ai_1 _4819_ (.B1(_1320_),
    .Y(_1387_),
    .A1(_1272_),
    .A2(_1318_));
 sg13g2_nand2_1 _4820_ (.Y(_1388_),
    .A(_1329_),
    .B(_1332_));
 sg13g2_or2_1 _4821_ (.X(_1389_),
    .B(_1313_),
    .A(\core.V[14] ));
 sg13g2_xnor2_1 _4822_ (.Y(_1390_),
    .A(\core.V[14] ),
    .B(_1313_));
 sg13g2_nand2_1 _4823_ (.Y(_1391_),
    .A(net718),
    .B(_1390_));
 sg13g2_nand2_1 _4824_ (.Y(_1392_),
    .A(net716),
    .B(_1315_));
 sg13g2_nand2_1 _4825_ (.Y(_1393_),
    .A(net713),
    .B(_1315_));
 sg13g2_xor2_1 _4826_ (.B(_1392_),
    .A(_1317_),
    .X(_1394_));
 sg13g2_nand2b_1 _4827_ (.Y(_1395_),
    .B(_1394_),
    .A_N(_1391_));
 sg13g2_xnor2_1 _4828_ (.Y(_1396_),
    .A(_1391_),
    .B(_1394_));
 sg13g2_and2_1 _4829_ (.A(_1388_),
    .B(_1396_),
    .X(_1397_));
 sg13g2_xor2_1 _4830_ (.B(_1396_),
    .A(_1388_),
    .X(_1398_));
 sg13g2_xnor2_1 _4831_ (.Y(_1399_),
    .A(_1387_),
    .B(_1398_));
 sg13g2_xnor2_1 _4832_ (.Y(_1400_),
    .A(_1386_),
    .B(_1399_));
 sg13g2_nor2_1 _4833_ (.A(_1367_),
    .B(_1400_),
    .Y(_1401_));
 sg13g2_xor2_1 _4834_ (.B(_1400_),
    .A(_1367_),
    .X(_1402_));
 sg13g2_xor2_1 _4835_ (.B(_1402_),
    .A(_1366_),
    .X(_1403_));
 sg13g2_nand2_1 _4836_ (.Y(_1404_),
    .A(_1365_),
    .B(_1403_));
 sg13g2_xnor2_1 _4837_ (.Y(_1405_),
    .A(_1365_),
    .B(_1403_));
 sg13g2_nor3_1 _4838_ (.A(_1348_),
    .B(_1349_),
    .C(_1405_),
    .Y(_1406_));
 sg13g2_o21ai_1 _4839_ (.B1(_1405_),
    .Y(_1407_),
    .A1(_1348_),
    .A2(_1349_));
 sg13g2_nand2b_1 _4840_ (.Y(_1408_),
    .B(_1407_),
    .A_N(_1406_));
 sg13g2_nor2b_1 _4841_ (.A(_1408_),
    .B_N(_1364_),
    .Y(_1409_));
 sg13g2_xor2_1 _4842_ (.B(_1408_),
    .A(_1364_),
    .X(_1410_));
 sg13g2_mux2_1 _4843_ (.A0(_1410_),
    .A1(_1354_),
    .S(net576),
    .X(_1411_));
 sg13g2_nand2_1 _4844_ (.Y(_1412_),
    .A(net577),
    .B(_1292_));
 sg13g2_o21ai_1 _4845_ (.B1(_1412_),
    .Y(_1413_),
    .A1(net578),
    .A2(_1411_));
 sg13g2_inv_1 _4846_ (.Y(_1414_),
    .A(_1413_));
 sg13g2_nand2b_1 _4847_ (.Y(_1415_),
    .B(net582),
    .A_N(_1300_));
 sg13g2_nand2_1 _4848_ (.Y(_1416_),
    .A(net582),
    .B(_1294_));
 sg13g2_o21ai_1 _4849_ (.B1(_1416_),
    .Y(_1417_),
    .A1(net582),
    .A2(_1302_));
 sg13g2_nor2_1 _4850_ (.A(_1227_),
    .B(_1417_),
    .Y(_1418_));
 sg13g2_a221oi_1 _4851_ (.B2(_1228_),
    .C1(_1418_),
    .B1(_1415_),
    .A1(_0842_),
    .Y(_1419_),
    .A2(_1414_));
 sg13g2_a22oi_1 _4852_ (.Y(_1420_),
    .B1(_0836_),
    .B2(_1419_),
    .A2(net638),
    .A1(net526));
 sg13g2_nor2_1 _4853_ (.A(net725),
    .B(_1420_),
    .Y(_0205_));
 sg13g2_nor2_1 _4854_ (.A(_1406_),
    .B(_1409_),
    .Y(_1421_));
 sg13g2_a21oi_1 _4855_ (.A1(_1366_),
    .A2(_1402_),
    .Y(_1422_),
    .B1(_1401_));
 sg13g2_o21ai_1 _4856_ (.B1(_1385_),
    .Y(_1423_),
    .A1(_1386_),
    .A2(_1399_));
 sg13g2_a21oi_1 _4857_ (.A1(_1387_),
    .A2(_1398_),
    .Y(_1424_),
    .B1(_1397_));
 sg13g2_nand2_1 _4858_ (.Y(_1425_),
    .A(net711),
    .B(_1270_));
 sg13g2_o21ai_1 _4859_ (.B1(_1380_),
    .Y(_1426_),
    .A1(\core.w[14] ),
    .A2(_1378_));
 sg13g2_xnor2_1 _4860_ (.Y(_1427_),
    .A(_1425_),
    .B(_1426_));
 sg13g2_nor2_1 _4861_ (.A(\core.V[8] ),
    .B(net652),
    .Y(_1428_));
 sg13g2_nand2b_1 _4862_ (.Y(_1429_),
    .B(net705),
    .A_N(net658));
 sg13g2_xnor2_1 _4863_ (.Y(_1430_),
    .A(\core.w[15] ),
    .B(_1429_));
 sg13g2_xnor2_1 _4864_ (.Y(_1431_),
    .A(_1428_),
    .B(_1430_));
 sg13g2_nand2_1 _4865_ (.Y(_1432_),
    .A(net709),
    .B(_1182_));
 sg13g2_xor2_1 _4866_ (.B(_1432_),
    .A(_1370_),
    .X(_1433_));
 sg13g2_xnor2_1 _4867_ (.Y(_1434_),
    .A(_1431_),
    .B(_1433_));
 sg13g2_xnor2_1 _4868_ (.Y(_1435_),
    .A(_1427_),
    .B(_1434_));
 sg13g2_o21ai_1 _4869_ (.B1(net718),
    .Y(_1436_),
    .A1(\core.V[15] ),
    .A2(_1389_));
 sg13g2_a21oi_1 _4870_ (.A1(\core.V[15] ),
    .A2(_1389_),
    .Y(_1437_),
    .B1(_1436_));
 sg13g2_nand2_1 _4871_ (.Y(_1438_),
    .A(_1371_),
    .B(_1374_));
 sg13g2_xnor2_1 _4872_ (.Y(_1439_),
    .A(_1437_),
    .B(_1438_));
 sg13g2_a21oi_1 _4873_ (.A1(_1318_),
    .A2(_1395_),
    .Y(_1440_),
    .B1(_1393_));
 sg13g2_a21o_1 _4874_ (.A2(_1395_),
    .A1(_1393_),
    .B1(_1440_),
    .X(_1441_));
 sg13g2_a21oi_1 _4875_ (.A1(_1375_),
    .A2(_1383_),
    .Y(_1442_),
    .B1(_1382_));
 sg13g2_nand2_1 _4876_ (.Y(_1443_),
    .A(net716),
    .B(_1390_));
 sg13g2_xnor2_1 _4877_ (.Y(_1444_),
    .A(_1435_),
    .B(_1442_));
 sg13g2_xnor2_1 _4878_ (.Y(_1445_),
    .A(_1439_),
    .B(_1443_));
 sg13g2_xnor2_1 _4879_ (.Y(_1446_),
    .A(_1444_),
    .B(_1445_));
 sg13g2_xnor2_1 _4880_ (.Y(_1447_),
    .A(_1441_),
    .B(_1446_));
 sg13g2_xnor2_1 _4881_ (.Y(_1448_),
    .A(_1423_),
    .B(_1447_));
 sg13g2_xnor2_1 _4882_ (.Y(_1449_),
    .A(_1424_),
    .B(_1448_));
 sg13g2_xnor2_1 _4883_ (.Y(_1450_),
    .A(_1422_),
    .B(_1449_));
 sg13g2_xnor2_1 _4884_ (.Y(_1451_),
    .A(_1404_),
    .B(_1450_));
 sg13g2_xnor2_1 _4885_ (.Y(_1452_),
    .A(_1421_),
    .B(_1451_));
 sg13g2_mux2_1 _4886_ (.A0(_1452_),
    .A1(_1410_),
    .S(net576),
    .X(_1453_));
 sg13g2_mux2_1 _4887_ (.A0(_1355_),
    .A1(_1453_),
    .S(_0845_),
    .X(_1454_));
 sg13g2_a22oi_1 _4888_ (.Y(_1455_),
    .B1(_1228_),
    .B2(_1242_),
    .A2(net586),
    .A1(_1225_));
 sg13g2_o21ai_1 _4889_ (.B1(_1455_),
    .Y(_1456_),
    .A1(_0841_),
    .A2(_1454_));
 sg13g2_a22oi_1 _4890_ (.Y(_1457_),
    .B1(_0836_),
    .B2(_1456_),
    .A2(net638),
    .A1(net782));
 sg13g2_nor2_1 _4891_ (.A(net725),
    .B(_1457_),
    .Y(_0206_));
 sg13g2_nand2_1 _4892_ (.Y(_1458_),
    .A(_0845_),
    .B(_1452_));
 sg13g2_nand2_1 _4893_ (.Y(_1459_),
    .A(net578),
    .B(_1411_));
 sg13g2_and2_1 _4894_ (.A(_1458_),
    .B(_1459_),
    .X(_1460_));
 sg13g2_and3_1 _4895_ (.X(_1461_),
    .A(_1228_),
    .B(_1301_),
    .C(_1303_));
 sg13g2_a221oi_1 _4896_ (.B2(_0842_),
    .C1(_1461_),
    .B1(_1460_),
    .A1(net586),
    .Y(_1462_),
    .A2(_1295_));
 sg13g2_inv_1 _4897_ (.Y(_1463_),
    .A(_1462_));
 sg13g2_a22oi_1 _4898_ (.Y(_1464_),
    .B1(_0836_),
    .B2(_1463_),
    .A2(net638),
    .A1(net542));
 sg13g2_nor2_1 _4899_ (.A(net725),
    .B(_1464_),
    .Y(_0207_));
 sg13g2_nand2_1 _4900_ (.Y(_1465_),
    .A(net578),
    .B(_1453_));
 sg13g2_nand2_1 _4901_ (.Y(_1466_),
    .A(_1458_),
    .B(_1465_));
 sg13g2_a22oi_1 _4902_ (.Y(_1467_),
    .B1(_1360_),
    .B2(_1228_),
    .A2(_1357_),
    .A1(net586));
 sg13g2_o21ai_1 _4903_ (.B1(_1467_),
    .Y(_1468_),
    .A1(_0841_),
    .A2(_1466_));
 sg13g2_a22oi_1 _4904_ (.Y(_1469_),
    .B1(_0836_),
    .B2(_1468_),
    .A2(net638),
    .A1(net485));
 sg13g2_nor2_1 _4905_ (.A(net734),
    .B(_1469_),
    .Y(_0208_));
 sg13g2_nand2b_2 _4906_ (.Y(_1470_),
    .B(_0836_),
    .A_N(_1452_));
 sg13g2_a21oi_2 _4907_ (.B1(_0837_),
    .Y(_1471_),
    .A2(_1452_),
    .A1(_0842_));
 sg13g2_nor2_1 _4908_ (.A(_1229_),
    .B(_1417_),
    .Y(_1472_));
 sg13g2_a21oi_1 _4909_ (.A1(_1226_),
    .A2(_1414_),
    .Y(_1473_),
    .B1(_1472_));
 sg13g2_a22oi_1 _4910_ (.Y(_1474_),
    .B1(_1471_),
    .B2(_1473_),
    .A2(net639),
    .A1(net757));
 sg13g2_nor2_1 _4911_ (.A(net734),
    .B(_1474_),
    .Y(_0209_));
 sg13g2_nor2_1 _4912_ (.A(_1225_),
    .B(_1229_),
    .Y(_1475_));
 sg13g2_a21oi_1 _4913_ (.A1(_1226_),
    .A2(_1454_),
    .Y(_1476_),
    .B1(_1475_));
 sg13g2_a22oi_1 _4914_ (.Y(_1477_),
    .B1(_1471_),
    .B2(_1476_),
    .A2(net639),
    .A1(net793));
 sg13g2_nor2_1 _4915_ (.A(net734),
    .B(_1477_),
    .Y(_0210_));
 sg13g2_nor2_1 _4916_ (.A(_1227_),
    .B(_1460_),
    .Y(_1478_));
 sg13g2_nor2_1 _4917_ (.A(_1229_),
    .B(_1295_),
    .Y(_1479_));
 sg13g2_nor2_1 _4918_ (.A(_1478_),
    .B(_1479_),
    .Y(_1480_));
 sg13g2_a22oi_1 _4919_ (.Y(_1481_),
    .B1(_1471_),
    .B2(_1480_),
    .A2(net639),
    .A1(net836));
 sg13g2_nor2_1 _4920_ (.A(net734),
    .B(_1481_),
    .Y(_0211_));
 sg13g2_nor2_1 _4921_ (.A(_1229_),
    .B(_1357_),
    .Y(_1482_));
 sg13g2_a21oi_1 _4922_ (.A1(net586),
    .A2(_1466_),
    .Y(_1483_),
    .B1(_1482_));
 sg13g2_a22oi_1 _4923_ (.Y(_1484_),
    .B1(_1471_),
    .B2(_1483_),
    .A2(net639),
    .A1(net552));
 sg13g2_nor2_1 _4924_ (.A(net734),
    .B(_1484_),
    .Y(_0212_));
 sg13g2_nand2_1 _4925_ (.Y(_1485_),
    .A(_1228_),
    .B(_1414_));
 sg13g2_a21oi_1 _4926_ (.A1(_1229_),
    .A2(_1452_),
    .Y(_1486_),
    .B1(_0837_));
 sg13g2_a22oi_1 _4927_ (.Y(_1487_),
    .B1(_1485_),
    .B2(_1486_),
    .A2(net639),
    .A1(net803));
 sg13g2_nor2_1 _4928_ (.A(net734),
    .B(net804),
    .Y(_0213_));
 sg13g2_nand2_1 _4929_ (.Y(_1488_),
    .A(net502),
    .B(net640));
 sg13g2_a21oi_1 _4930_ (.A1(_1470_),
    .A2(net503),
    .Y(_0214_),
    .B1(net733));
 sg13g2_nand2_1 _4931_ (.Y(_1489_),
    .A(net789),
    .B(net640));
 sg13g2_a21oi_1 _4932_ (.A1(_1470_),
    .A2(net790),
    .Y(_0215_),
    .B1(net733));
 sg13g2_nand2_1 _4933_ (.Y(_1490_),
    .A(net758),
    .B(net640));
 sg13g2_a21oi_1 _4934_ (.A1(_1470_),
    .A2(net759),
    .Y(_0216_),
    .B1(net733));
 sg13g2_nand2_1 _4935_ (.Y(_1491_),
    .A(net478),
    .B(net640));
 sg13g2_a21oi_1 _4936_ (.A1(_1470_),
    .A2(net479),
    .Y(_0217_),
    .B1(net733));
 sg13g2_nor3_2 _4937_ (.A(\core.capacitance[11] ),
    .B(\core.capacitance[9] ),
    .C(\core.capacitance[8] ),
    .Y(_1492_));
 sg13g2_nor2b_1 _4938_ (.A(\core.capacitance[10] ),
    .B_N(_1492_),
    .Y(_1493_));
 sg13g2_a21oi_1 _4939_ (.A1(_0030_),
    .A2(_1493_),
    .Y(_1494_),
    .B1(_2684_));
 sg13g2_xnor2_1 _4940_ (.Y(_1495_),
    .A(\core.capacitance[13] ),
    .B(_1494_));
 sg13g2_nor2_1 _4941_ (.A(\core.capacitance[13] ),
    .B(\core.capacitance[12] ),
    .Y(_1496_));
 sg13g2_nand3_1 _4942_ (.B(_1493_),
    .C(_1496_),
    .A(\core.capacitance[15] ),
    .Y(_1497_));
 sg13g2_mux2_1 _4943_ (.A0(_0031_),
    .A1(\core.capacitance[14] ),
    .S(\core.capacitance[15] ),
    .X(_1498_));
 sg13g2_nand2_1 _4944_ (.Y(_1499_),
    .A(_1497_),
    .B(_1498_));
 sg13g2_o21ai_1 _4945_ (.B1(_1499_),
    .Y(_1500_),
    .A1(\core.capacitance[14] ),
    .A2(_1497_));
 sg13g2_and2_2 _4946_ (.A(_1495_),
    .B(_1500_),
    .X(_1501_));
 sg13g2_o21ai_1 _4947_ (.B1(_1494_),
    .Y(_1502_),
    .A1(_0030_),
    .A2(_1493_));
 sg13g2_o21ai_1 _4948_ (.B1(_1502_),
    .Y(_1503_),
    .A1(\core.capacitance[15] ),
    .A2(_2689_));
 sg13g2_inv_1 _4949_ (.Y(_1504_),
    .A(_1503_));
 sg13g2_nor2_1 _4950_ (.A(_2684_),
    .B(_0045_),
    .Y(_1505_));
 sg13g2_a21oi_1 _4951_ (.A1(_2684_),
    .A2(\core.capacitance[10] ),
    .Y(_1506_),
    .B1(_1505_));
 sg13g2_nand4_1 _4952_ (.B(_1501_),
    .C(_1504_),
    .A(_1492_),
    .Y(_1507_),
    .D(_1506_));
 sg13g2_nor2_2 _4953_ (.A(_2730_),
    .B(_1497_),
    .Y(_1508_));
 sg13g2_or2_2 _4954_ (.X(_1509_),
    .B(_1497_),
    .A(_2730_));
 sg13g2_nand4_1 _4955_ (.B(\core.compute_state[1] ),
    .C(_1507_),
    .A(net739),
    .Y(_1510_),
    .D(_1509_));
 sg13g2_inv_1 _4956_ (.Y(_1511_),
    .A(_1510_));
 sg13g2_nor2_1 _4957_ (.A(_1495_),
    .B(_1500_),
    .Y(_1512_));
 sg13g2_and2_2 _4958_ (.A(_1503_),
    .B(_1512_),
    .X(_1513_));
 sg13g2_nor2_2 _4959_ (.A(_1508_),
    .B(_1513_),
    .Y(_1514_));
 sg13g2_nand2b_2 _4960_ (.Y(_1515_),
    .B(_1514_),
    .A_N(_1501_));
 sg13g2_inv_2 _4961_ (.Y(_1516_),
    .A(_1515_));
 sg13g2_nor2_1 _4962_ (.A(_1500_),
    .B(_1503_),
    .Y(_1517_));
 sg13g2_o21ai_1 _4963_ (.B1(_1509_),
    .Y(_1518_),
    .A1(_1495_),
    .A2(_1517_));
 sg13g2_inv_1 _4964_ (.Y(_1519_),
    .A(_1518_));
 sg13g2_nor3_1 _4965_ (.A(_1501_),
    .B(_1503_),
    .C(_1512_),
    .Y(_1520_));
 sg13g2_or2_1 _4966_ (.X(_1521_),
    .B(_1520_),
    .A(_1513_));
 sg13g2_a21oi_1 _4967_ (.A1(_0030_),
    .A2(_1508_),
    .Y(_1522_),
    .B1(_1521_));
 sg13g2_a21o_2 _4968_ (.A2(_1521_),
    .A1(_1508_),
    .B1(_1522_),
    .X(_1523_));
 sg13g2_nand2_1 _4969_ (.Y(_1524_),
    .A(_0036_),
    .B(net573));
 sg13g2_o21ai_1 _4970_ (.B1(_1524_),
    .Y(_1525_),
    .A1(_2734_),
    .A2(net572));
 sg13g2_o21ai_1 _4971_ (.B1(net592),
    .Y(_1526_),
    .A1(_0033_),
    .A2(net573));
 sg13g2_a21oi_1 _4972_ (.A1(_2732_),
    .A2(net572),
    .Y(_1527_),
    .B1(_1526_));
 sg13g2_a21o_1 _4973_ (.A2(_1525_),
    .A1(_1519_),
    .B1(_1527_),
    .X(_1528_));
 sg13g2_and2_1 _4974_ (.A(_1501_),
    .B(_1509_),
    .X(_1529_));
 sg13g2_nor2_1 _4975_ (.A(_0037_),
    .B(_1514_),
    .Y(_1530_));
 sg13g2_a21oi_1 _4976_ (.A1(_2731_),
    .A2(net591),
    .Y(_1531_),
    .B1(_1530_));
 sg13g2_o21ai_1 _4977_ (.B1(_1531_),
    .Y(_1532_),
    .A1(_1515_),
    .A2(_1528_));
 sg13g2_a22oi_1 _4978_ (.Y(_1533_),
    .B1(_1511_),
    .B2(_1532_),
    .A2(net646),
    .A1(net509));
 sg13g2_nor2_1 _4979_ (.A(net726),
    .B(net510),
    .Y(_0218_));
 sg13g2_mux2_1 _4980_ (.A0(_0042_),
    .A1(_0044_),
    .S(net573),
    .X(_1534_));
 sg13g2_nand2_1 _4981_ (.Y(_1535_),
    .A(_1518_),
    .B(_1534_));
 sg13g2_a21oi_1 _4982_ (.A1(_0043_),
    .A2(_1519_),
    .Y(_1536_),
    .B1(_1515_));
 sg13g2_nand2_1 _4983_ (.Y(_1537_),
    .A(_1535_),
    .B(_1536_));
 sg13g2_mux2_1 _4984_ (.A0(_0040_),
    .A1(_0041_),
    .S(net572),
    .X(_1538_));
 sg13g2_mux2_1 _4985_ (.A0(_0038_),
    .A1(_0039_),
    .S(net572),
    .X(_1539_));
 sg13g2_mux2_1 _4986_ (.A0(_1538_),
    .A1(_1539_),
    .S(net592),
    .X(_1540_));
 sg13g2_nor2_1 _4987_ (.A(_1516_),
    .B(_1540_),
    .Y(_1541_));
 sg13g2_mux2_1 _4988_ (.A0(_0036_),
    .A1(_0037_),
    .S(net573),
    .X(_1542_));
 sg13g2_o21ai_1 _4989_ (.B1(net592),
    .Y(_1543_),
    .A1(_0034_),
    .A2(net572));
 sg13g2_a21oi_1 _4990_ (.A1(_2734_),
    .A2(net572),
    .Y(_1544_),
    .B1(_1543_));
 sg13g2_a21o_1 _4991_ (.A2(_1542_),
    .A1(_1519_),
    .B1(_1544_),
    .X(_1545_));
 sg13g2_nor2_1 _4992_ (.A(_1515_),
    .B(_1545_),
    .Y(_1546_));
 sg13g2_a21oi_1 _4993_ (.A1(_2733_),
    .A2(net591),
    .Y(_1547_),
    .B1(_1546_));
 sg13g2_o21ai_1 _4994_ (.B1(_1547_),
    .Y(_1548_),
    .A1(_1514_),
    .A2(_1540_));
 sg13g2_a22oi_1 _4995_ (.Y(_1549_),
    .B1(_1511_),
    .B2(_1548_),
    .A2(net646),
    .A1(net515));
 sg13g2_nor2_1 _4996_ (.A(net726),
    .B(net516),
    .Y(_0219_));
 sg13g2_mux2_1 _4997_ (.A0(_0044_),
    .A1(_0043_),
    .S(net573),
    .X(_1550_));
 sg13g2_nand2_1 _4998_ (.Y(_1551_),
    .A(_1518_),
    .B(_1550_));
 sg13g2_mux2_1 _4999_ (.A0(_0041_),
    .A1(_0042_),
    .S(net573),
    .X(_1552_));
 sg13g2_mux2_1 _5000_ (.A0(_0039_),
    .A1(_0040_),
    .S(net572),
    .X(_1553_));
 sg13g2_mux2_1 _5001_ (.A0(_1552_),
    .A1(_1553_),
    .S(net592),
    .X(_1554_));
 sg13g2_nor2_1 _5002_ (.A(_1516_),
    .B(_1554_),
    .Y(_1555_));
 sg13g2_a21oi_2 _5003_ (.B1(_1555_),
    .Y(_1556_),
    .A2(_1551_),
    .A1(_1536_));
 sg13g2_mux2_1 _5004_ (.A0(_0037_),
    .A1(_0038_),
    .S(net572),
    .X(_1557_));
 sg13g2_mux2_1 _5005_ (.A0(_1525_),
    .A1(_1557_),
    .S(_1519_),
    .X(_1558_));
 sg13g2_nor2_1 _5006_ (.A(_1515_),
    .B(_1558_),
    .Y(_1559_));
 sg13g2_a21oi_1 _5007_ (.A1(_2732_),
    .A2(net591),
    .Y(_1560_),
    .B1(_1559_));
 sg13g2_o21ai_1 _5008_ (.B1(_1560_),
    .Y(_1561_),
    .A1(_1514_),
    .A2(_1556_));
 sg13g2_a22oi_1 _5009_ (.Y(_1562_),
    .B1(_1511_),
    .B2(_1561_),
    .A2(net646),
    .A1(net519));
 sg13g2_nor2_1 _5010_ (.A(net724),
    .B(net520),
    .Y(_0220_));
 sg13g2_mux2_1 _5011_ (.A0(_1534_),
    .A1(_1538_),
    .S(net592),
    .X(_1563_));
 sg13g2_mux2_1 _5012_ (.A0(_1539_),
    .A1(_1542_),
    .S(net592),
    .X(_1564_));
 sg13g2_nor2_1 _5013_ (.A(_1515_),
    .B(_1564_),
    .Y(_1565_));
 sg13g2_a21oi_1 _5014_ (.A1(_2734_),
    .A2(net591),
    .Y(_1566_),
    .B1(_1565_));
 sg13g2_o21ai_1 _5015_ (.B1(_1566_),
    .Y(_1567_),
    .A1(_1514_),
    .A2(_1563_));
 sg13g2_a22oi_1 _5016_ (.Y(_1568_),
    .B1(_1511_),
    .B2(_1567_),
    .A2(net646),
    .A1(net523));
 sg13g2_nor2_1 _5017_ (.A(net724),
    .B(net524),
    .Y(_0221_));
 sg13g2_mux2_1 _5018_ (.A0(_1553_),
    .A1(_1557_),
    .S(net592),
    .X(_1569_));
 sg13g2_a21oi_1 _5019_ (.A1(_0041_),
    .A2(_1513_),
    .Y(_1570_),
    .B1(_1510_));
 sg13g2_a22oi_1 _5020_ (.Y(_1571_),
    .B1(_1569_),
    .B2(_1516_),
    .A2(net591),
    .A1(_1528_));
 sg13g2_a22oi_1 _5021_ (.Y(_1572_),
    .B1(_1570_),
    .B2(_1571_),
    .A2(net646),
    .A1(net545));
 sg13g2_nor2_1 _5022_ (.A(net722),
    .B(net546),
    .Y(_0222_));
 sg13g2_a21oi_1 _5023_ (.A1(_0042_),
    .A2(_1513_),
    .Y(_1573_),
    .B1(_1510_));
 sg13g2_a22oi_1 _5024_ (.Y(_1574_),
    .B1(_1545_),
    .B2(net591),
    .A2(_1540_),
    .A1(_1516_));
 sg13g2_a22oi_1 _5025_ (.Y(_1575_),
    .B1(_1573_),
    .B2(_1574_),
    .A2(net646),
    .A1(net527));
 sg13g2_nor2_1 _5026_ (.A(net721),
    .B(net528),
    .Y(_0223_));
 sg13g2_a21oi_1 _5027_ (.A1(_0044_),
    .A2(_1513_),
    .Y(_1576_),
    .B1(_1510_));
 sg13g2_a22oi_1 _5028_ (.Y(_1577_),
    .B1(_1558_),
    .B2(net591),
    .A2(_1554_),
    .A1(_1516_));
 sg13g2_a22oi_1 _5029_ (.Y(_1578_),
    .B1(_1576_),
    .B2(_1577_),
    .A2(net646),
    .A1(net461));
 sg13g2_nor2_1 _5030_ (.A(net721),
    .B(net462),
    .Y(_0224_));
 sg13g2_nor2_2 _5031_ (.A(_0043_),
    .B(_1510_),
    .Y(_1579_));
 sg13g2_a21oi_2 _5032_ (.B1(_1510_),
    .Y(_1580_),
    .A2(_1513_),
    .A1(_0043_));
 sg13g2_a22oi_1 _5033_ (.Y(_1581_),
    .B1(_1564_),
    .B2(_1529_),
    .A2(_1563_),
    .A1(_1516_));
 sg13g2_a22oi_1 _5034_ (.Y(_1582_),
    .B1(_1580_),
    .B2(_1581_),
    .A2(net646),
    .A1(net538));
 sg13g2_nor2_1 _5035_ (.A(net721),
    .B(net539),
    .Y(_0225_));
 sg13g2_mux2_1 _5036_ (.A0(_1550_),
    .A1(_1552_),
    .S(net592),
    .X(_1583_));
 sg13g2_a22oi_1 _5037_ (.Y(_1584_),
    .B1(_1583_),
    .B2(_1516_),
    .A2(_1569_),
    .A1(_1501_));
 sg13g2_nand2b_1 _5038_ (.Y(_1585_),
    .B(_1514_),
    .A_N(_1584_));
 sg13g2_a22oi_1 _5039_ (.Y(_1586_),
    .B1(_1580_),
    .B2(_1585_),
    .A2(net647),
    .A1(net801));
 sg13g2_nor2_1 _5040_ (.A(net721),
    .B(net802),
    .Y(_0226_));
 sg13g2_nand3b_1 _5041_ (.B(_1514_),
    .C(_1537_),
    .Y(_1587_),
    .A_N(_1541_));
 sg13g2_a22oi_1 _5042_ (.Y(_1588_),
    .B1(_1580_),
    .B2(_1587_),
    .A2(net647),
    .A1(net837));
 sg13g2_nor2_1 _5043_ (.A(net721),
    .B(net838),
    .Y(_0227_));
 sg13g2_nand2_1 _5044_ (.Y(_1589_),
    .A(_1514_),
    .B(_1556_));
 sg13g2_a22oi_1 _5045_ (.Y(_1590_),
    .B1(_1580_),
    .B2(_1589_),
    .A2(net647),
    .A1(net774));
 sg13g2_nor2_1 _5046_ (.A(net721),
    .B(net775),
    .Y(_0228_));
 sg13g2_nor2_1 _5047_ (.A(_1515_),
    .B(_1579_),
    .Y(_1591_));
 sg13g2_a21oi_1 _5048_ (.A1(net591),
    .A2(_1563_),
    .Y(_1592_),
    .B1(_1591_));
 sg13g2_a22oi_1 _5049_ (.Y(_1593_),
    .B1(_1580_),
    .B2(_1592_),
    .A2(net647),
    .A1(net832));
 sg13g2_nor2_1 _5050_ (.A(net721),
    .B(net833),
    .Y(_0229_));
 sg13g2_a21oi_1 _5051_ (.A1(net796),
    .A2(net648),
    .Y(_1594_),
    .B1(_1579_));
 sg13g2_nor2_1 _5052_ (.A(net730),
    .B(net797),
    .Y(_0230_));
 sg13g2_a21oi_1 _5053_ (.A1(net817),
    .A2(net648),
    .Y(_1595_),
    .B1(_1579_));
 sg13g2_nor2_1 _5054_ (.A(net730),
    .B(net818),
    .Y(_0231_));
 sg13g2_a21oi_1 _5055_ (.A1(net558),
    .A2(net648),
    .Y(_1596_),
    .B1(_1579_));
 sg13g2_nor2_1 _5056_ (.A(net730),
    .B(net559),
    .Y(_0232_));
 sg13g2_a21oi_1 _5057_ (.A1(net512),
    .A2(net648),
    .Y(_1597_),
    .B1(_1579_));
 sg13g2_nor2_1 _5058_ (.A(net730),
    .B(net513),
    .Y(_0233_));
 sg13g2_nand2b_1 _5059_ (.Y(_1598_),
    .B(\core.exp_term[1] ),
    .A_N(\core.w[1] ));
 sg13g2_xnor2_1 _5060_ (.Y(_1599_),
    .A(\core.exp_term[1] ),
    .B(\core.w[1] ));
 sg13g2_nand2_1 _5061_ (.Y(_1600_),
    .A(\core.leak_current[1] ),
    .B(_1599_));
 sg13g2_xor2_1 _5062_ (.B(_1599_),
    .A(\core.leak_current[1] ),
    .X(_1601_));
 sg13g2_nand2_1 _5063_ (.Y(_1602_),
    .A(_0018_),
    .B(_1601_));
 sg13g2_nor2b_1 _5064_ (.A(\core.w[2] ),
    .B_N(\core.exp_term[2] ),
    .Y(_1603_));
 sg13g2_xnor2_1 _5065_ (.Y(_1604_),
    .A(\core.exp_term[2] ),
    .B(\core.w[2] ));
 sg13g2_xnor2_1 _5066_ (.Y(_1605_),
    .A(\core.leak_current[2] ),
    .B(_1604_));
 sg13g2_a21oi_2 _5067_ (.B1(_1605_),
    .Y(_1606_),
    .A2(_1600_),
    .A1(_1598_));
 sg13g2_nand3_1 _5068_ (.B(_1600_),
    .C(_1605_),
    .A(_1598_),
    .Y(_1607_));
 sg13g2_nor2b_1 _5069_ (.A(_1606_),
    .B_N(_1607_),
    .Y(_1608_));
 sg13g2_nand2b_1 _5070_ (.Y(_1609_),
    .B(_1608_),
    .A_N(_1602_));
 sg13g2_a21oi_1 _5071_ (.A1(\core.leak_current[2] ),
    .A2(_1604_),
    .Y(_1610_),
    .B1(_1603_));
 sg13g2_nor2b_1 _5072_ (.A(\core.w[3] ),
    .B_N(\core.exp_term[3] ),
    .Y(_1611_));
 sg13g2_xnor2_1 _5073_ (.Y(_1612_),
    .A(\core.exp_term[3] ),
    .B(\core.w[3] ));
 sg13g2_xnor2_1 _5074_ (.Y(_1613_),
    .A(\core.leak_current[3] ),
    .B(_1612_));
 sg13g2_nor2_1 _5075_ (.A(_1610_),
    .B(_1613_),
    .Y(_1614_));
 sg13g2_xor2_1 _5076_ (.B(_1613_),
    .A(_1610_),
    .X(_1615_));
 sg13g2_nand2_1 _5077_ (.Y(_1616_),
    .A(_1606_),
    .B(_1615_));
 sg13g2_xnor2_1 _5078_ (.Y(_1617_),
    .A(_1606_),
    .B(_1615_));
 sg13g2_or2_1 _5079_ (.X(_1618_),
    .B(_1617_),
    .A(_1609_));
 sg13g2_xnor2_1 _5080_ (.Y(_1619_),
    .A(_1609_),
    .B(_1617_));
 sg13g2_o21ai_1 _5081_ (.B1(net747),
    .Y(_1620_),
    .A1(net771),
    .A2(net636));
 sg13g2_a21oi_1 _5082_ (.A1(net636),
    .A2(_1619_),
    .Y(_0234_),
    .B1(_1620_));
 sg13g2_a21oi_1 _5083_ (.A1(\core.leak_current[3] ),
    .A2(_1612_),
    .Y(_1621_),
    .B1(_1611_));
 sg13g2_nor2b_1 _5084_ (.A(\core.w[4] ),
    .B_N(\core.exp_term[4] ),
    .Y(_1622_));
 sg13g2_xnor2_1 _5085_ (.Y(_1623_),
    .A(\core.exp_term[4] ),
    .B(\core.w[4] ));
 sg13g2_xnor2_1 _5086_ (.Y(_1624_),
    .A(\core.leak_current[4] ),
    .B(_1623_));
 sg13g2_nor2_1 _5087_ (.A(_1621_),
    .B(_1624_),
    .Y(_1625_));
 sg13g2_xor2_1 _5088_ (.B(_1624_),
    .A(_1621_),
    .X(_1626_));
 sg13g2_and2_1 _5089_ (.A(_1614_),
    .B(_1626_),
    .X(_1627_));
 sg13g2_xnor2_1 _5090_ (.Y(_1628_),
    .A(_1614_),
    .B(_1626_));
 sg13g2_a21oi_1 _5091_ (.A1(_1616_),
    .A2(_1618_),
    .Y(_1629_),
    .B1(_1628_));
 sg13g2_nand3_1 _5092_ (.B(_1618_),
    .C(_1628_),
    .A(_1616_),
    .Y(_1630_));
 sg13g2_nand2b_1 _5093_ (.Y(_1631_),
    .B(_1630_),
    .A_N(_1629_));
 sg13g2_o21ai_1 _5094_ (.B1(net747),
    .Y(_1632_),
    .A1(net495),
    .A2(net635));
 sg13g2_a21oi_1 _5095_ (.A1(net636),
    .A2(_1631_),
    .Y(_0235_),
    .B1(_1632_));
 sg13g2_a21oi_1 _5096_ (.A1(\core.leak_current[4] ),
    .A2(_1623_),
    .Y(_1633_),
    .B1(_1622_));
 sg13g2_nor2b_1 _5097_ (.A(\core.w[5] ),
    .B_N(\core.exp_term[5] ),
    .Y(_1634_));
 sg13g2_xnor2_1 _5098_ (.Y(_1635_),
    .A(\core.exp_term[5] ),
    .B(\core.w[5] ));
 sg13g2_xnor2_1 _5099_ (.Y(_1636_),
    .A(\core.leak_current[5] ),
    .B(_1635_));
 sg13g2_nor2_1 _5100_ (.A(_1633_),
    .B(_1636_),
    .Y(_1637_));
 sg13g2_xor2_1 _5101_ (.B(_1636_),
    .A(_1633_),
    .X(_1638_));
 sg13g2_nand2_1 _5102_ (.Y(_1639_),
    .A(_1625_),
    .B(_1638_));
 sg13g2_xor2_1 _5103_ (.B(_1638_),
    .A(_1625_),
    .X(_1640_));
 sg13g2_o21ai_1 _5104_ (.B1(_1640_),
    .Y(_1641_),
    .A1(_1627_),
    .A2(_1629_));
 sg13g2_or3_1 _5105_ (.A(_1627_),
    .B(_1629_),
    .C(_1640_),
    .X(_1642_));
 sg13g2_a21oi_1 _5106_ (.A1(_1641_),
    .A2(_1642_),
    .Y(_1643_),
    .B1(_2755_));
 sg13g2_o21ai_1 _5107_ (.B1(net746),
    .Y(_1644_),
    .A1(net554),
    .A2(net636));
 sg13g2_nor2_1 _5108_ (.A(_1643_),
    .B(_1644_),
    .Y(_0236_));
 sg13g2_a21oi_1 _5109_ (.A1(\core.leak_current[5] ),
    .A2(_1635_),
    .Y(_1645_),
    .B1(_1634_));
 sg13g2_nand2b_1 _5110_ (.Y(_1646_),
    .B(\core.exp_term[6] ),
    .A_N(\core.w[6] ));
 sg13g2_xnor2_1 _5111_ (.Y(_1647_),
    .A(\core.exp_term[6] ),
    .B(\core.w[6] ));
 sg13g2_nand2_1 _5112_ (.Y(_1648_),
    .A(\core.leak_current[6] ),
    .B(_1647_));
 sg13g2_xnor2_1 _5113_ (.Y(_1649_),
    .A(\core.leak_current[6] ),
    .B(_1647_));
 sg13g2_nor2_1 _5114_ (.A(_1645_),
    .B(_1649_),
    .Y(_1650_));
 sg13g2_xor2_1 _5115_ (.B(_1649_),
    .A(_1645_),
    .X(_1651_));
 sg13g2_nand2_1 _5116_ (.Y(_1652_),
    .A(_1637_),
    .B(_1651_));
 sg13g2_xnor2_1 _5117_ (.Y(_1653_),
    .A(_1637_),
    .B(_1651_));
 sg13g2_a21o_1 _5118_ (.A2(_1641_),
    .A1(_1639_),
    .B1(_1653_),
    .X(_1654_));
 sg13g2_nand3_1 _5119_ (.B(_1641_),
    .C(_1653_),
    .A(_1639_),
    .Y(_1655_));
 sg13g2_a21oi_1 _5120_ (.A1(_1654_),
    .A2(_1655_),
    .Y(_1656_),
    .B1(_2755_));
 sg13g2_o21ai_1 _5121_ (.B1(net746),
    .Y(_1657_),
    .A1(net566),
    .A2(net636));
 sg13g2_nor2_1 _5122_ (.A(_1656_),
    .B(_1657_),
    .Y(_0237_));
 sg13g2_nor2b_1 _5123_ (.A(\core.w[7] ),
    .B_N(\core.exp_term[7] ),
    .Y(_1658_));
 sg13g2_xnor2_1 _5124_ (.Y(_1659_),
    .A(\core.exp_term[7] ),
    .B(\core.w[7] ));
 sg13g2_xnor2_1 _5125_ (.Y(_1660_),
    .A(\core.leak_current[7] ),
    .B(_1659_));
 sg13g2_a21oi_1 _5126_ (.A1(_1646_),
    .A2(_1648_),
    .Y(_1661_),
    .B1(_1660_));
 sg13g2_inv_1 _5127_ (.Y(_1662_),
    .A(_1661_));
 sg13g2_nand3_1 _5128_ (.B(_1648_),
    .C(_1660_),
    .A(_1646_),
    .Y(_1663_));
 sg13g2_nor2b_1 _5129_ (.A(_1661_),
    .B_N(_1663_),
    .Y(_1664_));
 sg13g2_nand2_1 _5130_ (.Y(_1665_),
    .A(_1650_),
    .B(_1664_));
 sg13g2_xnor2_1 _5131_ (.Y(_1666_),
    .A(_1650_),
    .B(_1664_));
 sg13g2_a21o_1 _5132_ (.A2(_1654_),
    .A1(_1652_),
    .B1(_1666_),
    .X(_1667_));
 sg13g2_nand3_1 _5133_ (.B(_1654_),
    .C(_1666_),
    .A(_1652_),
    .Y(_1668_));
 sg13g2_a21oi_1 _5134_ (.A1(_1667_),
    .A2(_1668_),
    .Y(_1669_),
    .B1(_2755_));
 sg13g2_o21ai_1 _5135_ (.B1(net746),
    .Y(_1670_),
    .A1(net560),
    .A2(net636));
 sg13g2_nor2_1 _5136_ (.A(_1669_),
    .B(_1670_),
    .Y(_0238_));
 sg13g2_a21oi_1 _5137_ (.A1(\core.leak_current[7] ),
    .A2(_1659_),
    .Y(_1671_),
    .B1(_1658_));
 sg13g2_nor2b_1 _5138_ (.A(\core.w[8] ),
    .B_N(\core.ibias[8] ),
    .Y(_1672_));
 sg13g2_xnor2_1 _5139_ (.Y(_1673_),
    .A(\core.w[8] ),
    .B(\core.ibias[8] ));
 sg13g2_xnor2_1 _5140_ (.Y(_1674_),
    .A(\core.exp_term[8] ),
    .B(_1673_));
 sg13g2_nor2_1 _5141_ (.A(_1671_),
    .B(_1674_),
    .Y(_1675_));
 sg13g2_xor2_1 _5142_ (.B(_1674_),
    .A(_1671_),
    .X(_1676_));
 sg13g2_xnor2_1 _5143_ (.Y(_1677_),
    .A(\core.leak_current[8] ),
    .B(_1676_));
 sg13g2_nor2_1 _5144_ (.A(_1662_),
    .B(_1677_),
    .Y(_1678_));
 sg13g2_xnor2_1 _5145_ (.Y(_1679_),
    .A(_1662_),
    .B(_1677_));
 sg13g2_a21oi_1 _5146_ (.A1(_1665_),
    .A2(_1667_),
    .Y(_1680_),
    .B1(_1679_));
 sg13g2_nand3_1 _5147_ (.B(_1667_),
    .C(_1679_),
    .A(_1665_),
    .Y(_1681_));
 sg13g2_nand2b_1 _5148_ (.Y(_1682_),
    .B(_1681_),
    .A_N(_1680_));
 sg13g2_o21ai_1 _5149_ (.B1(net742),
    .Y(_1683_),
    .A1(net499),
    .A2(net636));
 sg13g2_a21oi_1 _5150_ (.A1(net635),
    .A2(_1682_),
    .Y(_0239_),
    .B1(_1683_));
 sg13g2_a21oi_1 _5151_ (.A1(\core.leak_current[8] ),
    .A2(_1676_),
    .Y(_1684_),
    .B1(_1675_));
 sg13g2_a21oi_1 _5152_ (.A1(\core.exp_term[8] ),
    .A2(_1673_),
    .Y(_1685_),
    .B1(_1672_));
 sg13g2_nor2b_1 _5153_ (.A(\core.w[9] ),
    .B_N(\core.ibias[9] ),
    .Y(_1686_));
 sg13g2_xnor2_1 _5154_ (.Y(_1687_),
    .A(\core.w[9] ),
    .B(\core.ibias[9] ));
 sg13g2_xnor2_1 _5155_ (.Y(_1688_),
    .A(\core.exp_term[9] ),
    .B(_1687_));
 sg13g2_nor2_1 _5156_ (.A(_1685_),
    .B(_1688_),
    .Y(_1689_));
 sg13g2_xor2_1 _5157_ (.B(_1688_),
    .A(_1685_),
    .X(_1690_));
 sg13g2_xnor2_1 _5158_ (.Y(_1691_),
    .A(\core.leak_current[9] ),
    .B(_1690_));
 sg13g2_xor2_1 _5159_ (.B(_1691_),
    .A(_1684_),
    .X(_1692_));
 sg13g2_o21ai_1 _5160_ (.B1(_1692_),
    .Y(_1693_),
    .A1(_1678_),
    .A2(_1680_));
 sg13g2_or3_1 _5161_ (.A(_1678_),
    .B(_1680_),
    .C(_1692_),
    .X(_1694_));
 sg13g2_a21oi_1 _5162_ (.A1(_1693_),
    .A2(_1694_),
    .Y(_1695_),
    .B1(_2755_));
 sg13g2_o21ai_1 _5163_ (.B1(net743),
    .Y(_1696_),
    .A1(net563),
    .A2(net635));
 sg13g2_nor2_1 _5164_ (.A(_1695_),
    .B(_1696_),
    .Y(_0240_));
 sg13g2_o21ai_1 _5165_ (.B1(_1693_),
    .Y(_1697_),
    .A1(_1684_),
    .A2(_1691_));
 sg13g2_a21oi_1 _5166_ (.A1(\core.leak_current[9] ),
    .A2(_1690_),
    .Y(_1698_),
    .B1(_1689_));
 sg13g2_a21oi_1 _5167_ (.A1(\core.exp_term[9] ),
    .A2(_1687_),
    .Y(_1699_),
    .B1(_1686_));
 sg13g2_nor2b_1 _5168_ (.A(\core.w[10] ),
    .B_N(\core.ibias[10] ),
    .Y(_1700_));
 sg13g2_xnor2_1 _5169_ (.Y(_1701_),
    .A(\core.w[10] ),
    .B(\core.ibias[10] ));
 sg13g2_xnor2_1 _5170_ (.Y(_1702_),
    .A(\core.exp_term[10] ),
    .B(_1701_));
 sg13g2_nor2_1 _5171_ (.A(_1699_),
    .B(_1702_),
    .Y(_1703_));
 sg13g2_xor2_1 _5172_ (.B(_1702_),
    .A(_1699_),
    .X(_1704_));
 sg13g2_xnor2_1 _5173_ (.Y(_1705_),
    .A(\core.leak_current[10] ),
    .B(_1704_));
 sg13g2_nor2_1 _5174_ (.A(_1698_),
    .B(_1705_),
    .Y(_1706_));
 sg13g2_xor2_1 _5175_ (.B(_1705_),
    .A(_1698_),
    .X(_1707_));
 sg13g2_xnor2_1 _5176_ (.Y(_1708_),
    .A(_1697_),
    .B(_1707_));
 sg13g2_o21ai_1 _5177_ (.B1(net742),
    .Y(_1709_),
    .A1(net493),
    .A2(net635));
 sg13g2_a21oi_1 _5178_ (.A1(net635),
    .A2(_1708_),
    .Y(_0241_),
    .B1(_1709_));
 sg13g2_a21o_1 _5179_ (.A2(_1707_),
    .A1(_1697_),
    .B1(_1706_),
    .X(_1710_));
 sg13g2_a21oi_1 _5180_ (.A1(\core.leak_current[10] ),
    .A2(_1704_),
    .Y(_1711_),
    .B1(_1703_));
 sg13g2_a21oi_1 _5181_ (.A1(\core.exp_term[10] ),
    .A2(_1701_),
    .Y(_1712_),
    .B1(_1700_));
 sg13g2_nor2b_1 _5182_ (.A(\core.w[11] ),
    .B_N(\core.ibias[11] ),
    .Y(_1713_));
 sg13g2_xnor2_1 _5183_ (.Y(_1714_),
    .A(\core.w[11] ),
    .B(\core.ibias[11] ));
 sg13g2_xnor2_1 _5184_ (.Y(_1715_),
    .A(\core.exp_term[11] ),
    .B(_1714_));
 sg13g2_nor2_1 _5185_ (.A(_1712_),
    .B(_1715_),
    .Y(_1716_));
 sg13g2_xor2_1 _5186_ (.B(_1715_),
    .A(_1712_),
    .X(_1717_));
 sg13g2_xnor2_1 _5187_ (.Y(_1718_),
    .A(\core.leak_current[11] ),
    .B(_1717_));
 sg13g2_nor2_1 _5188_ (.A(_1711_),
    .B(_1718_),
    .Y(_1719_));
 sg13g2_xor2_1 _5189_ (.B(_1718_),
    .A(_1711_),
    .X(_1720_));
 sg13g2_and2_1 _5190_ (.A(_1710_),
    .B(_1720_),
    .X(_1721_));
 sg13g2_xnor2_1 _5191_ (.Y(_1722_),
    .A(_1710_),
    .B(_1720_));
 sg13g2_o21ai_1 _5192_ (.B1(net742),
    .Y(_1723_),
    .A1(net772),
    .A2(net635));
 sg13g2_a21oi_1 _5193_ (.A1(net635),
    .A2(_1722_),
    .Y(_0242_),
    .B1(_1723_));
 sg13g2_a21oi_1 _5194_ (.A1(\core.leak_current[11] ),
    .A2(_1717_),
    .Y(_1724_),
    .B1(_1716_));
 sg13g2_a21oi_1 _5195_ (.A1(\core.exp_term[11] ),
    .A2(_1714_),
    .Y(_1725_),
    .B1(_1713_));
 sg13g2_nor2b_1 _5196_ (.A(\core.w[12] ),
    .B_N(\core.ibias[12] ),
    .Y(_1726_));
 sg13g2_xnor2_1 _5197_ (.Y(_1727_),
    .A(\core.w[12] ),
    .B(\core.ibias[12] ));
 sg13g2_xnor2_1 _5198_ (.Y(_1728_),
    .A(\core.exp_term[12] ),
    .B(_1727_));
 sg13g2_or2_1 _5199_ (.X(_1729_),
    .B(_1728_),
    .A(_1725_));
 sg13g2_xor2_1 _5200_ (.B(_1728_),
    .A(_1725_),
    .X(_1730_));
 sg13g2_nand2_1 _5201_ (.Y(_1731_),
    .A(\core.leak_current[12] ),
    .B(_1730_));
 sg13g2_xnor2_1 _5202_ (.Y(_1732_),
    .A(\core.leak_current[12] ),
    .B(_1730_));
 sg13g2_nor2_1 _5203_ (.A(_1724_),
    .B(_1732_),
    .Y(_1733_));
 sg13g2_xor2_1 _5204_ (.B(_1732_),
    .A(_1724_),
    .X(_1734_));
 sg13g2_o21ai_1 _5205_ (.B1(_1734_),
    .Y(_1735_),
    .A1(_1719_),
    .A2(_1721_));
 sg13g2_or3_1 _5206_ (.A(_1719_),
    .B(_1721_),
    .C(_1734_),
    .X(_1736_));
 sg13g2_a21oi_1 _5207_ (.A1(_1735_),
    .A2(_1736_),
    .Y(_1737_),
    .B1(_2755_));
 sg13g2_o21ai_1 _5208_ (.B1(net743),
    .Y(_1738_),
    .A1(net532),
    .A2(net635));
 sg13g2_nor2_1 _5209_ (.A(_1737_),
    .B(_1738_),
    .Y(_0243_));
 sg13g2_o21ai_1 _5210_ (.B1(net743),
    .Y(_1739_),
    .A1(net488),
    .A2(net637));
 sg13g2_nor2b_1 _5211_ (.A(_1733_),
    .B_N(_1735_),
    .Y(_1740_));
 sg13g2_a21oi_1 _5212_ (.A1(\core.exp_term[12] ),
    .A2(_1727_),
    .Y(_1741_),
    .B1(_1726_));
 sg13g2_nor2b_1 _5213_ (.A(\core.w[13] ),
    .B_N(\core.ibias[13] ),
    .Y(_1742_));
 sg13g2_xnor2_1 _5214_ (.Y(_1743_),
    .A(\core.w[13] ),
    .B(\core.ibias[13] ));
 sg13g2_xnor2_1 _5215_ (.Y(_1744_),
    .A(\core.exp_term[13] ),
    .B(_1743_));
 sg13g2_nor2_1 _5216_ (.A(_1741_),
    .B(_1744_),
    .Y(_1745_));
 sg13g2_xor2_1 _5217_ (.B(_1744_),
    .A(_1741_),
    .X(_1746_));
 sg13g2_xnor2_1 _5218_ (.Y(_1747_),
    .A(\core.leak_current[13] ),
    .B(_1746_));
 sg13g2_nand3_1 _5219_ (.B(_1731_),
    .C(_1747_),
    .A(_1729_),
    .Y(_1748_));
 sg13g2_a21oi_1 _5220_ (.A1(_1729_),
    .A2(_1731_),
    .Y(_1749_),
    .B1(_1747_));
 sg13g2_inv_1 _5221_ (.Y(_1750_),
    .A(_1749_));
 sg13g2_nand2_1 _5222_ (.Y(_1751_),
    .A(_1748_),
    .B(_1750_));
 sg13g2_xnor2_1 _5223_ (.Y(_1752_),
    .A(_1740_),
    .B(_1751_));
 sg13g2_a21oi_1 _5224_ (.A1(net637),
    .A2(_1752_),
    .Y(_0244_),
    .B1(_1739_));
 sg13g2_a21oi_1 _5225_ (.A1(\core.leak_current[13] ),
    .A2(_1746_),
    .Y(_1753_),
    .B1(_1745_));
 sg13g2_a21oi_1 _5226_ (.A1(\core.exp_term[13] ),
    .A2(_1743_),
    .Y(_1754_),
    .B1(_1742_));
 sg13g2_nor2b_1 _5227_ (.A(\core.w[14] ),
    .B_N(\core.ibias[14] ),
    .Y(_1755_));
 sg13g2_xnor2_1 _5228_ (.Y(_1756_),
    .A(\core.w[14] ),
    .B(\core.ibias[14] ));
 sg13g2_xnor2_1 _5229_ (.Y(_1757_),
    .A(\core.exp_term[14] ),
    .B(_1756_));
 sg13g2_nor2_1 _5230_ (.A(_1754_),
    .B(_1757_),
    .Y(_1758_));
 sg13g2_xor2_1 _5231_ (.B(_1757_),
    .A(_1754_),
    .X(_1759_));
 sg13g2_xnor2_1 _5232_ (.Y(_1760_),
    .A(\core.leak_current[14] ),
    .B(_1759_));
 sg13g2_xor2_1 _5233_ (.B(_1760_),
    .A(_1753_),
    .X(_1761_));
 sg13g2_nor2b_1 _5234_ (.A(_1740_),
    .B_N(_1748_),
    .Y(_1762_));
 sg13g2_o21ai_1 _5235_ (.B1(_1761_),
    .Y(_1763_),
    .A1(_1749_),
    .A2(_1762_));
 sg13g2_or3_1 _5236_ (.A(_1749_),
    .B(_1761_),
    .C(_1762_),
    .X(_1764_));
 sg13g2_nand2_1 _5237_ (.Y(_1765_),
    .A(_1763_),
    .B(_1764_));
 sg13g2_o21ai_1 _5238_ (.B1(net745),
    .Y(_1766_),
    .A1(net557),
    .A2(net637));
 sg13g2_a21oi_1 _5239_ (.A1(net637),
    .A2(_1765_),
    .Y(_0245_),
    .B1(_1766_));
 sg13g2_o21ai_1 _5240_ (.B1(net745),
    .Y(_1767_),
    .A1(net487),
    .A2(net637));
 sg13g2_o21ai_1 _5241_ (.B1(_1763_),
    .Y(_1768_),
    .A1(_1753_),
    .A2(_1760_));
 sg13g2_a21oi_1 _5242_ (.A1(\core.leak_current[14] ),
    .A2(_1759_),
    .Y(_1769_),
    .B1(_1758_));
 sg13g2_a21oi_1 _5243_ (.A1(\core.exp_term[14] ),
    .A2(_1756_),
    .Y(_1770_),
    .B1(_1755_));
 sg13g2_xnor2_1 _5244_ (.Y(_1771_),
    .A(\core.exp_term[15] ),
    .B(\core.w[15] ));
 sg13g2_xnor2_1 _5245_ (.Y(_1772_),
    .A(\core.ibias[15] ),
    .B(_1771_));
 sg13g2_xnor2_1 _5246_ (.Y(_1773_),
    .A(_1770_),
    .B(_1772_));
 sg13g2_xnor2_1 _5247_ (.Y(_1774_),
    .A(\core.leak_current[15] ),
    .B(_1773_));
 sg13g2_xnor2_1 _5248_ (.Y(_1775_),
    .A(_1769_),
    .B(_1774_));
 sg13g2_xnor2_1 _5249_ (.Y(_1776_),
    .A(_1768_),
    .B(_1775_));
 sg13g2_a21oi_1 _5250_ (.A1(net637),
    .A2(_1776_),
    .Y(_0246_),
    .B1(_1767_));
 sg13g2_o21ai_1 _5251_ (.B1(net750),
    .Y(_1777_),
    .A1(net695),
    .A2(net421));
 sg13g2_a21oi_1 _5252_ (.A1(net695),
    .A2(_2644_),
    .Y(_0247_),
    .B1(_1777_));
 sg13g2_a21oi_1 _5253_ (.A1(net695),
    .A2(net382),
    .Y(_1778_),
    .B1(net732));
 sg13g2_o21ai_1 _5254_ (.B1(_1778_),
    .Y(_0248_),
    .A1(net693),
    .A2(_2642_));
 sg13g2_a21oi_1 _5255_ (.A1(net692),
    .A2(net376),
    .Y(_1779_),
    .B1(net732));
 sg13g2_o21ai_1 _5256_ (.B1(_1779_),
    .Y(_0249_),
    .A1(net692),
    .A2(_2640_));
 sg13g2_a21oi_2 _5257_ (.B1(net732),
    .Y(_1780_),
    .A2(net475),
    .A1(net693));
 sg13g2_o21ai_1 _5258_ (.B1(_1780_),
    .Y(_0250_),
    .A1(net687),
    .A2(_2638_));
 sg13g2_o21ai_1 _5259_ (.B1(net756),
    .Y(_1781_),
    .A1(net692),
    .A2(net398));
 sg13g2_a21oi_1 _5260_ (.A1(net692),
    .A2(_2637_),
    .Y(_0251_),
    .B1(_1781_));
 sg13g2_o21ai_1 _5261_ (.B1(net750),
    .Y(_1782_),
    .A1(net692),
    .A2(net404));
 sg13g2_a21oi_1 _5262_ (.A1(net695),
    .A2(_2636_),
    .Y(_0252_),
    .B1(_1782_));
 sg13g2_a21oi_1 _5263_ (.A1(net692),
    .A2(net374),
    .Y(_1783_),
    .B1(net732));
 sg13g2_o21ai_1 _5264_ (.B1(_1783_),
    .Y(_0253_),
    .A1(net692),
    .A2(_2634_));
 sg13g2_a21oi_1 _5265_ (.A1(net311),
    .A2(net695),
    .Y(_1784_),
    .B1(net732));
 sg13g2_o21ai_1 _5266_ (.B1(_1784_),
    .Y(_0254_),
    .A1(_2632_),
    .A2(net692));
 sg13g2_nor2_1 _5267_ (.A(\core.V_threshold[15] ),
    .B(_0816_),
    .Y(_1785_));
 sg13g2_nand2_1 _5268_ (.Y(_1786_),
    .A(\core.V_threshold[14] ),
    .B(_0813_));
 sg13g2_nand2_1 _5269_ (.Y(_1787_),
    .A(\core.V_threshold[13] ),
    .B(_0807_));
 sg13g2_nor2_1 _5270_ (.A(\core.V_threshold[13] ),
    .B(_0807_),
    .Y(_1788_));
 sg13g2_nand2_1 _5271_ (.Y(_1789_),
    .A(\core.V_threshold[12] ),
    .B(_0804_));
 sg13g2_nor2_1 _5272_ (.A(\core.V_threshold[11] ),
    .B(_0800_),
    .Y(_1790_));
 sg13g2_nor2_1 _5273_ (.A(\core.V_threshold[10] ),
    .B(_0795_),
    .Y(_1791_));
 sg13g2_xor2_1 _5274_ (.B(\core.dV[9] ),
    .A(net657),
    .X(_1792_));
 sg13g2_xnor2_1 _5275_ (.Y(_1793_),
    .A(_0792_),
    .B(_1792_));
 sg13g2_nor2_1 _5276_ (.A(\core.V_threshold[9] ),
    .B(_1793_),
    .Y(_1794_));
 sg13g2_xnor2_1 _5277_ (.Y(_1795_),
    .A(_0790_),
    .B(_0791_));
 sg13g2_xnor2_1 _5278_ (.Y(_1796_),
    .A(_0767_),
    .B(_0788_));
 sg13g2_xnor2_1 _5279_ (.Y(_1797_),
    .A(_0770_),
    .B(_0787_));
 sg13g2_xor2_1 _5280_ (.B(_0785_),
    .A(_0771_),
    .X(_1798_));
 sg13g2_xnor2_1 _5281_ (.Y(_1799_),
    .A(_0773_),
    .B(_0783_));
 sg13g2_xnor2_1 _5282_ (.Y(_1800_),
    .A(_0781_),
    .B(_0782_));
 sg13g2_xor2_1 _5283_ (.B(_0780_),
    .A(_0779_),
    .X(_1801_));
 sg13g2_or2_1 _5284_ (.X(_1802_),
    .B(\core.dV[0] ),
    .A(net678));
 sg13g2_o21ai_1 _5285_ (.B1(_0778_),
    .Y(_1803_),
    .A1(_0777_),
    .A2(_1802_));
 sg13g2_nand4_1 _5286_ (.B(_1799_),
    .C(_1800_),
    .A(_1798_),
    .Y(_1804_),
    .D(_1803_));
 sg13g2_nor4_2 _5287_ (.A(_1796_),
    .B(_1797_),
    .C(_1801_),
    .Y(_1805_),
    .D(_1804_));
 sg13g2_o21ai_1 _5288_ (.B1(_1795_),
    .Y(_1806_),
    .A1(\core.V_threshold[8] ),
    .A2(_1805_));
 sg13g2_nand2_1 _5289_ (.Y(_1807_),
    .A(\core.V_threshold[8] ),
    .B(_1805_));
 sg13g2_a21oi_1 _5290_ (.A1(_1806_),
    .A2(_1807_),
    .Y(_1808_),
    .B1(_1794_));
 sg13g2_a221oi_1 _5291_ (.B2(\core.V_threshold[9] ),
    .C1(_1808_),
    .B1(_1793_),
    .A1(\core.V_threshold[10] ),
    .Y(_1809_),
    .A2(_0795_));
 sg13g2_nor2_1 _5292_ (.A(_1791_),
    .B(_1809_),
    .Y(_1810_));
 sg13g2_a21oi_1 _5293_ (.A1(\core.V_threshold[11] ),
    .A2(_0800_),
    .Y(_1811_),
    .B1(_1810_));
 sg13g2_o21ai_1 _5294_ (.B1(_1789_),
    .Y(_1812_),
    .A1(_1790_),
    .A2(_1811_));
 sg13g2_o21ai_1 _5295_ (.B1(_1812_),
    .Y(_1813_),
    .A1(\core.V_threshold[12] ),
    .A2(_0804_));
 sg13g2_a21oi_1 _5296_ (.A1(_1787_),
    .A2(_1813_),
    .Y(_1814_),
    .B1(_1788_));
 sg13g2_o21ai_1 _5297_ (.B1(_1814_),
    .Y(_1815_),
    .A1(\core.V_threshold[14] ),
    .A2(_0813_));
 sg13g2_a22oi_1 _5298_ (.Y(_1816_),
    .B1(_1786_),
    .B2(_1815_),
    .A2(_0816_),
    .A1(\core.V_threshold[15] ));
 sg13g2_nor2_2 _5299_ (.A(_1785_),
    .B(_1816_),
    .Y(_1817_));
 sg13g2_inv_1 _5300_ (.Y(_1818_),
    .A(net569));
 sg13g2_a22oi_1 _5301_ (.Y(_1819_),
    .B1(net630),
    .B2(_1817_),
    .A2(net650),
    .A1(net468));
 sg13g2_inv_1 _5302_ (.Y(_0255_),
    .A(net469));
 sg13g2_nor2_1 _5303_ (.A(net724),
    .B(net634),
    .Y(_1820_));
 sg13g2_nor3_1 _5304_ (.A(_2631_),
    .B(net725),
    .C(net634),
    .Y(_1821_));
 sg13g2_nand3_1 _5305_ (.B(_0741_),
    .C(_0746_),
    .A(_0735_),
    .Y(_1822_));
 sg13g2_nand4_1 _5306_ (.B(_0758_),
    .C(_0761_),
    .A(_0751_),
    .Y(_1823_),
    .D(_1822_));
 sg13g2_xor2_1 _5307_ (.B(\core.dw[9] ),
    .A(\core.w[9] ),
    .X(_1824_));
 sg13g2_xnor2_1 _5308_ (.Y(_1825_),
    .A(_0731_),
    .B(_1824_));
 sg13g2_xnor2_1 _5309_ (.Y(_1826_),
    .A(_0706_),
    .B(_0727_));
 sg13g2_xnor2_1 _5310_ (.Y(_1827_),
    .A(_0724_),
    .B(_0726_));
 sg13g2_xnor2_1 _5311_ (.Y(_1828_),
    .A(_0721_),
    .B(_0722_));
 sg13g2_xnor2_1 _5312_ (.Y(_1829_),
    .A(_0718_),
    .B(_0720_));
 sg13g2_xnor2_1 _5313_ (.Y(_1830_),
    .A(_0710_),
    .B(_0717_));
 sg13g2_xnor2_1 _5314_ (.Y(_1831_),
    .A(_0715_),
    .B(_0716_));
 sg13g2_xnor2_1 _5315_ (.Y(_1832_),
    .A(\core.w[0] ),
    .B(\core.dw[0] ));
 sg13g2_xnor2_1 _5316_ (.Y(_1833_),
    .A(_0713_),
    .B(_0714_));
 sg13g2_nand4_1 _5317_ (.B(_1831_),
    .C(_1832_),
    .A(_1830_),
    .Y(_1834_),
    .D(_1833_));
 sg13g2_nor4_1 _5318_ (.A(_1827_),
    .B(_1828_),
    .C(_1829_),
    .D(_1834_),
    .Y(_1835_));
 sg13g2_nand2b_1 _5319_ (.Y(_1836_),
    .B(_1835_),
    .A_N(_1826_));
 sg13g2_xor2_1 _5320_ (.B(_0729_),
    .A(_0728_),
    .X(_1837_));
 sg13g2_nand3_1 _5321_ (.B(_1836_),
    .C(_1837_),
    .A(_1825_),
    .Y(_1838_));
 sg13g2_nor4_2 _5322_ (.A(_0751_),
    .B(_0758_),
    .C(_1822_),
    .Y(_1839_),
    .D(_1838_));
 sg13g2_nand2b_2 _5323_ (.Y(_1840_),
    .B(_1839_),
    .A_N(_0761_));
 sg13g2_and2_1 _5324_ (.A(_1823_),
    .B(_1840_),
    .X(_1841_));
 sg13g2_nor2_1 _5325_ (.A(net628),
    .B(_1832_),
    .Y(_1842_));
 sg13g2_a21o_1 _5326_ (.A2(_1842_),
    .A1(net571),
    .B1(_1821_),
    .X(_0256_));
 sg13g2_nor2_1 _5327_ (.A(net628),
    .B(_1833_),
    .Y(_1843_));
 sg13g2_a22oi_1 _5328_ (.Y(_1844_),
    .B1(net571),
    .B2(_1843_),
    .A2(net625),
    .A1(net878));
 sg13g2_inv_1 _5329_ (.Y(_0257_),
    .A(_1844_));
 sg13g2_nor2_1 _5330_ (.A(net628),
    .B(_1831_),
    .Y(_1845_));
 sg13g2_a22oi_1 _5331_ (.Y(_1846_),
    .B1(net571),
    .B2(_1845_),
    .A2(net625),
    .A1(net882));
 sg13g2_inv_1 _5332_ (.Y(_0258_),
    .A(_1846_));
 sg13g2_nor2_1 _5333_ (.A(net628),
    .B(_1830_),
    .Y(_1847_));
 sg13g2_a22oi_1 _5334_ (.Y(_1848_),
    .B1(net571),
    .B2(_1847_),
    .A2(net625),
    .A1(net888));
 sg13g2_inv_1 _5335_ (.Y(_0259_),
    .A(_1848_));
 sg13g2_nand2_1 _5336_ (.Y(_1849_),
    .A(net885),
    .B(net627));
 sg13g2_nand3_1 _5337_ (.B(_1829_),
    .C(net571),
    .A(net630),
    .Y(_1850_));
 sg13g2_nand2_1 _5338_ (.Y(_0260_),
    .A(_1849_),
    .B(_1850_));
 sg13g2_nand2_1 _5339_ (.Y(_1851_),
    .A(net890),
    .B(net627));
 sg13g2_nand3_1 _5340_ (.B(_1828_),
    .C(net571),
    .A(net630),
    .Y(_1852_));
 sg13g2_nand2_1 _5341_ (.Y(_0261_),
    .A(_1851_),
    .B(_1852_));
 sg13g2_nand2_1 _5342_ (.Y(_1853_),
    .A(net875),
    .B(net627));
 sg13g2_nand3_1 _5343_ (.B(_1827_),
    .C(net571),
    .A(net630),
    .Y(_1854_));
 sg13g2_nand2_1 _5344_ (.Y(_0262_),
    .A(_1853_),
    .B(_1854_));
 sg13g2_nand2_1 _5345_ (.Y(_1855_),
    .A(net881),
    .B(net626));
 sg13g2_nand3_1 _5346_ (.B(_1826_),
    .C(net571),
    .A(net630),
    .Y(_1856_));
 sg13g2_nand2_1 _5347_ (.Y(_0263_),
    .A(_1855_),
    .B(_1856_));
 sg13g2_nand2_1 _5348_ (.Y(_1857_),
    .A(\core.param_b[8] ),
    .B(net570));
 sg13g2_xor2_1 _5349_ (.B(_1857_),
    .A(_1837_),
    .X(_1858_));
 sg13g2_and2_1 _5350_ (.A(net630),
    .B(_1823_),
    .X(_1859_));
 sg13g2_inv_1 _5351_ (.Y(_1860_),
    .A(_1859_));
 sg13g2_a21oi_1 _5352_ (.A1(_1840_),
    .A2(_1858_),
    .Y(_1861_),
    .B1(_1860_));
 sg13g2_a21o_1 _5353_ (.A2(net626),
    .A1(\core.w[8] ),
    .B1(_1861_),
    .X(_0264_));
 sg13g2_nand2_1 _5354_ (.Y(_1862_),
    .A(\core.param_b[8] ),
    .B(_1837_));
 sg13g2_nand2_1 _5355_ (.Y(_1863_),
    .A(\core.param_b[9] ),
    .B(_1825_));
 sg13g2_xor2_1 _5356_ (.B(_1825_),
    .A(\core.param_b[9] ),
    .X(_1864_));
 sg13g2_nand2b_1 _5357_ (.Y(_1865_),
    .B(_1864_),
    .A_N(_1862_));
 sg13g2_xnor2_1 _5358_ (.Y(_1866_),
    .A(_1862_),
    .B(_1864_));
 sg13g2_nand2_1 _5359_ (.Y(_1867_),
    .A(net569),
    .B(_1866_));
 sg13g2_nand2_1 _5360_ (.Y(_1868_),
    .A(_1818_),
    .B(_1825_));
 sg13g2_nand3_1 _5361_ (.B(_1867_),
    .C(_1868_),
    .A(_1840_),
    .Y(_1869_));
 sg13g2_a22oi_1 _5362_ (.Y(_1870_),
    .B1(_1859_),
    .B2(_1869_),
    .A2(net626),
    .A1(\core.w[9] ));
 sg13g2_inv_1 _5363_ (.Y(_0265_),
    .A(_1870_));
 sg13g2_xnor2_1 _5364_ (.Y(_1871_),
    .A(\core.param_b[10] ),
    .B(_0735_));
 sg13g2_a21oi_1 _5365_ (.A1(_1863_),
    .A2(_1865_),
    .Y(_1872_),
    .B1(_1871_));
 sg13g2_nand3_1 _5366_ (.B(_1865_),
    .C(_1871_),
    .A(_1863_),
    .Y(_1873_));
 sg13g2_nor2b_1 _5367_ (.A(_1872_),
    .B_N(_1873_),
    .Y(_1874_));
 sg13g2_nand2_1 _5368_ (.Y(_1875_),
    .A(net570),
    .B(_1874_));
 sg13g2_nand2_1 _5369_ (.Y(_1876_),
    .A(net634),
    .B(_1841_));
 sg13g2_a21oi_1 _5370_ (.A1(_0735_),
    .A2(_1818_),
    .Y(_1877_),
    .B1(_1876_));
 sg13g2_nand2_1 _5371_ (.Y(_1878_),
    .A(net891),
    .B(net751));
 sg13g2_a22oi_1 _5372_ (.Y(_0266_),
    .B1(_1878_),
    .B2(net628),
    .A2(_1877_),
    .A1(_1875_));
 sg13g2_nand2_1 _5373_ (.Y(_1879_),
    .A(_0741_),
    .B(_1818_));
 sg13g2_a21oi_1 _5374_ (.A1(\core.param_b[10] ),
    .A2(_0735_),
    .Y(_1880_),
    .B1(_1872_));
 sg13g2_xor2_1 _5375_ (.B(_0741_),
    .A(\core.param_b[11] ),
    .X(_1881_));
 sg13g2_nor2b_1 _5376_ (.A(_1880_),
    .B_N(_1881_),
    .Y(_1882_));
 sg13g2_xnor2_1 _5377_ (.Y(_1883_),
    .A(_1880_),
    .B(_1881_));
 sg13g2_a21oi_1 _5378_ (.A1(net570),
    .A2(_1883_),
    .Y(_1884_),
    .B1(_1876_));
 sg13g2_nand2_1 _5379_ (.Y(_1885_),
    .A(net887),
    .B(net751));
 sg13g2_a22oi_1 _5380_ (.Y(_0267_),
    .B1(_1885_),
    .B2(net628),
    .A2(_1884_),
    .A1(_1879_));
 sg13g2_nand2_1 _5381_ (.Y(_1886_),
    .A(_0746_),
    .B(_1818_));
 sg13g2_a21oi_1 _5382_ (.A1(\core.param_b[11] ),
    .A2(_0741_),
    .Y(_1887_),
    .B1(_1882_));
 sg13g2_xnor2_1 _5383_ (.Y(_1888_),
    .A(\core.param_b[12] ),
    .B(_0746_));
 sg13g2_nor2_1 _5384_ (.A(_1887_),
    .B(_1888_),
    .Y(_1889_));
 sg13g2_xor2_1 _5385_ (.B(_1888_),
    .A(_1887_),
    .X(_1890_));
 sg13g2_a21oi_1 _5386_ (.A1(net569),
    .A2(_1890_),
    .Y(_1891_),
    .B1(_1876_));
 sg13g2_nand2_1 _5387_ (.Y(_1892_),
    .A(net877),
    .B(net751));
 sg13g2_a22oi_1 _5388_ (.Y(_0268_),
    .B1(_1892_),
    .B2(net628),
    .A2(_1891_),
    .A1(_1886_));
 sg13g2_a21oi_1 _5389_ (.A1(\core.param_b[12] ),
    .A2(_0746_),
    .Y(_1893_),
    .B1(_1889_));
 sg13g2_nand2_1 _5390_ (.Y(_1894_),
    .A(\core.param_b[13] ),
    .B(_0752_));
 sg13g2_xor2_1 _5391_ (.B(_0751_),
    .A(\core.param_b[13] ),
    .X(_1895_));
 sg13g2_xor2_1 _5392_ (.B(_1895_),
    .A(_1893_),
    .X(_1896_));
 sg13g2_o21ai_1 _5393_ (.B1(_1840_),
    .Y(_1897_),
    .A1(_0751_),
    .A2(net569));
 sg13g2_a21o_1 _5394_ (.A2(_1896_),
    .A1(net569),
    .B1(_1897_),
    .X(_1898_));
 sg13g2_a22oi_1 _5395_ (.Y(_1899_),
    .B1(_1859_),
    .B2(_1898_),
    .A2(net626),
    .A1(net886));
 sg13g2_inv_1 _5396_ (.Y(_0269_),
    .A(_1899_));
 sg13g2_o21ai_1 _5397_ (.B1(_1894_),
    .Y(_1900_),
    .A1(_1893_),
    .A2(_1895_));
 sg13g2_xnor2_1 _5398_ (.Y(_1901_),
    .A(_2696_),
    .B(_0758_));
 sg13g2_nand2b_1 _5399_ (.Y(_1902_),
    .B(_1900_),
    .A_N(_1901_));
 sg13g2_xnor2_1 _5400_ (.Y(_1903_),
    .A(_1900_),
    .B(_1901_));
 sg13g2_o21ai_1 _5401_ (.B1(_1840_),
    .Y(_1904_),
    .A1(_0758_),
    .A2(net569));
 sg13g2_a21o_1 _5402_ (.A2(_1903_),
    .A1(net569),
    .B1(_1904_),
    .X(_1905_));
 sg13g2_a22oi_1 _5403_ (.Y(_1906_),
    .B1(_1859_),
    .B2(_1905_),
    .A2(net626),
    .A1(net873));
 sg13g2_inv_1 _5404_ (.Y(_0270_),
    .A(_1906_));
 sg13g2_o21ai_1 _5405_ (.B1(_1902_),
    .Y(_1907_),
    .A1(_2696_),
    .A2(_0758_));
 sg13g2_xor2_1 _5406_ (.B(_0761_),
    .A(\core.param_b[15] ),
    .X(_1908_));
 sg13g2_xnor2_1 _5407_ (.Y(_1909_),
    .A(_1907_),
    .B(_1908_));
 sg13g2_nand2_1 _5408_ (.Y(_1910_),
    .A(net569),
    .B(_1909_));
 sg13g2_nor2_1 _5409_ (.A(_1818_),
    .B(_1839_),
    .Y(_1911_));
 sg13g2_o21ai_1 _5410_ (.B1(_1910_),
    .Y(_1912_),
    .A1(_0761_),
    .A2(_1911_));
 sg13g2_nand3_1 _5411_ (.B(_1823_),
    .C(_1912_),
    .A(net634),
    .Y(_1913_));
 sg13g2_o21ai_1 _5412_ (.B1(_1913_),
    .Y(_1914_),
    .A1(net871),
    .A2(net634));
 sg13g2_nor2_1 _5413_ (.A(net733),
    .B(_1914_),
    .Y(_0271_));
 sg13g2_nor3_1 _5414_ (.A(_2630_),
    .B(net726),
    .C(net634),
    .Y(_0272_));
 sg13g2_and2_1 _5415_ (.A(net675),
    .B(net625),
    .X(_0273_));
 sg13g2_and2_1 _5416_ (.A(net674),
    .B(net625),
    .X(_0274_));
 sg13g2_and2_1 _5417_ (.A(net672),
    .B(net626),
    .X(_0275_));
 sg13g2_and2_1 _5418_ (.A(net669),
    .B(net625),
    .X(_0276_));
 sg13g2_and2_1 _5419_ (.A(net667),
    .B(net626),
    .X(_0277_));
 sg13g2_and2_1 _5420_ (.A(net665),
    .B(net625),
    .X(_0278_));
 sg13g2_and2_1 _5421_ (.A(net663),
    .B(net625),
    .X(_0279_));
 sg13g2_a21o_1 _5422_ (.A2(_0699_),
    .A1(net660),
    .B1(net724),
    .X(_0280_));
 sg13g2_a21o_1 _5423_ (.A2(_1793_),
    .A1(_0795_),
    .B1(_0800_),
    .X(_1915_));
 sg13g2_a21oi_1 _5424_ (.A1(_0804_),
    .A2(_1915_),
    .Y(_1916_),
    .B1(_0807_));
 sg13g2_nand3b_1 _5425_ (.B(_0816_),
    .C(_1916_),
    .Y(_1917_),
    .A_N(_0813_));
 sg13g2_nand2_1 _5426_ (.Y(_1918_),
    .A(net634),
    .B(_1917_));
 sg13g2_nand2_1 _5427_ (.Y(_1919_),
    .A(net744),
    .B(_1918_));
 sg13g2_a21o_1 _5428_ (.A2(_0699_),
    .A1(net657),
    .B1(_1919_),
    .X(_0281_));
 sg13g2_o21ai_1 _5429_ (.B1(_1918_),
    .Y(_1920_),
    .A1(net656),
    .A2(net634));
 sg13g2_nand2_1 _5430_ (.Y(_0282_),
    .A(net744),
    .B(_1920_));
 sg13g2_a21o_1 _5431_ (.A2(_0699_),
    .A1(net655),
    .B1(_1919_),
    .X(_0283_));
 sg13g2_a21o_1 _5432_ (.A2(_0699_),
    .A1(net654),
    .B1(net722),
    .X(_0284_));
 sg13g2_nand2b_1 _5433_ (.Y(_0285_),
    .B(net626),
    .A_N(net496));
 sg13g2_a21oi_1 _5434_ (.A1(_2629_),
    .A2(_0699_),
    .Y(_0286_),
    .B1(net722));
 sg13g2_a21o_1 _5435_ (.A2(_0699_),
    .A1(net859),
    .B1(net724),
    .X(_0287_));
 sg13g2_nand2b_1 _5436_ (.Y(_1921_),
    .B(net684),
    .A_N(net685));
 sg13g2_nor2_1 _5437_ (.A(_2848_),
    .B(_1921_),
    .Y(_1922_));
 sg13g2_nor2_2 _5438_ (.A(net732),
    .B(net608),
    .Y(_1923_));
 sg13g2_a22oi_1 _5439_ (.Y(_1924_),
    .B1(_1923_),
    .B2(net350),
    .A2(_1922_),
    .A1(\core.byte_acc[0] ));
 sg13g2_inv_1 _5440_ (.Y(_0288_),
    .A(net351));
 sg13g2_a22oi_1 _5441_ (.Y(_0289_),
    .B1(_1923_),
    .B2(_2643_),
    .A2(net608),
    .A1(_2627_));
 sg13g2_a22oi_1 _5442_ (.Y(_0290_),
    .B1(_1923_),
    .B2(_2641_),
    .A2(net608),
    .A1(_2626_));
 sg13g2_a22oi_1 _5443_ (.Y(_0291_),
    .B1(_1923_),
    .B2(_2639_),
    .A2(net608),
    .A1(_2625_));
 sg13g2_a22oi_1 _5444_ (.Y(_1925_),
    .B1(_1923_),
    .B2(net328),
    .A2(net608),
    .A1(\core.byte_acc[4] ));
 sg13g2_inv_1 _5445_ (.Y(_0292_),
    .A(net329));
 sg13g2_a22oi_1 _5446_ (.Y(_1926_),
    .B1(_1923_),
    .B2(net380),
    .A2(net608),
    .A1(\core.byte_acc[5] ));
 sg13g2_inv_1 _5447_ (.Y(_0293_),
    .A(net381));
 sg13g2_a22oi_1 _5448_ (.Y(_0294_),
    .B1(_1923_),
    .B2(_2635_),
    .A2(net608),
    .A1(_2623_));
 sg13g2_a22oi_1 _5449_ (.Y(_1927_),
    .B1(_1923_),
    .B2(net315),
    .A2(net608),
    .A1(\core.byte_acc[7] ));
 sg13g2_inv_1 _5450_ (.Y(_0295_),
    .A(net316));
 sg13g2_nand2b_1 _5451_ (.Y(_1928_),
    .B(\core.param_idx[1] ),
    .A_N(\core.param_idx[2] ));
 sg13g2_nor2_1 _5452_ (.A(_2848_),
    .B(_1928_),
    .Y(_1929_));
 sg13g2_nor2_2 _5453_ (.A(net735),
    .B(net607),
    .Y(_1930_));
 sg13g2_a22oi_1 _5454_ (.Y(_1931_),
    .B1(_1930_),
    .B2(net364),
    .A2(net607),
    .A1(\core.byte_acc[0] ));
 sg13g2_inv_1 _5455_ (.Y(_0296_),
    .A(net365));
 sg13g2_a22oi_1 _5456_ (.Y(_1932_),
    .B1(_1930_),
    .B2(net361),
    .A2(net607),
    .A1(\core.byte_acc[1] ));
 sg13g2_inv_1 _5457_ (.Y(_0297_),
    .A(net362));
 sg13g2_a22oi_1 _5458_ (.Y(_1933_),
    .B1(_1930_),
    .B2(net356),
    .A2(_1929_),
    .A1(\core.byte_acc[2] ));
 sg13g2_inv_1 _5459_ (.Y(_0298_),
    .A(net357));
 sg13g2_a22oi_1 _5460_ (.Y(_0299_),
    .B1(_1930_),
    .B2(_2701_),
    .A2(net607),
    .A1(_2625_));
 sg13g2_a22oi_1 _5461_ (.Y(_1934_),
    .B1(_1930_),
    .B2(net336),
    .A2(net607),
    .A1(\core.byte_acc[4] ));
 sg13g2_inv_1 _5462_ (.Y(_0300_),
    .A(net337));
 sg13g2_a22oi_1 _5463_ (.Y(_0301_),
    .B1(_1930_),
    .B2(_2698_),
    .A2(net607),
    .A1(_2624_));
 sg13g2_a22oi_1 _5464_ (.Y(_1935_),
    .B1(_1930_),
    .B2(net354),
    .A2(net607),
    .A1(\core.byte_acc[6] ));
 sg13g2_inv_1 _5465_ (.Y(_0302_),
    .A(net355));
 sg13g2_a22oi_1 _5466_ (.Y(_0303_),
    .B1(_1930_),
    .B2(_2695_),
    .A2(net607),
    .A1(_2622_));
 sg13g2_nor2_2 _5467_ (.A(_2807_),
    .B(_1928_),
    .Y(_1936_));
 sg13g2_nor2_2 _5468_ (.A(net735),
    .B(net606),
    .Y(_1937_));
 sg13g2_a22oi_1 _5469_ (.Y(_1938_),
    .B1(_1937_),
    .B2(net500),
    .A2(net606),
    .A1(net521));
 sg13g2_inv_1 _5470_ (.Y(_0304_),
    .A(_1938_));
 sg13g2_a22oi_1 _5471_ (.Y(_0305_),
    .B1(_1937_),
    .B2(_2682_),
    .A2(net606),
    .A1(_2627_));
 sg13g2_a22oi_1 _5472_ (.Y(_1939_),
    .B1(_1937_),
    .B2(net470),
    .A2(net606),
    .A1(net798));
 sg13g2_inv_1 _5473_ (.Y(_0306_),
    .A(_1939_));
 sg13g2_a22oi_1 _5474_ (.Y(_1940_),
    .B1(_1937_),
    .B2(net359),
    .A2(net606),
    .A1(net454));
 sg13g2_inv_1 _5475_ (.Y(_0307_),
    .A(_1940_));
 sg13g2_a22oi_1 _5476_ (.Y(_1941_),
    .B1(_1937_),
    .B2(net322),
    .A2(net606),
    .A1(\core.byte_acc[4] ));
 sg13g2_inv_1 _5477_ (.Y(_0308_),
    .A(net323));
 sg13g2_a22oi_1 _5478_ (.Y(_1942_),
    .B1(_1937_),
    .B2(net338),
    .A2(net606),
    .A1(\core.byte_acc[5] ));
 sg13g2_inv_1 _5479_ (.Y(_0309_),
    .A(net339));
 sg13g2_a22oi_1 _5480_ (.Y(_1943_),
    .B1(_1937_),
    .B2(net399),
    .A2(net606),
    .A1(\core.byte_acc[6] ));
 sg13g2_inv_1 _5481_ (.Y(_0310_),
    .A(net400));
 sg13g2_a22oi_1 _5482_ (.Y(_0311_),
    .B1(_1937_),
    .B2(_2675_),
    .A2(_1936_),
    .A1(_2622_));
 sg13g2_nor3_2 _5483_ (.A(\core.param_idx[1] ),
    .B(net684),
    .C(_2848_),
    .Y(_1944_));
 sg13g2_nor2_2 _5484_ (.A(net735),
    .B(net605),
    .Y(_1945_));
 sg13g2_a22oi_1 _5485_ (.Y(_1946_),
    .B1(_1945_),
    .B2(net352),
    .A2(net605),
    .A1(\core.byte_acc[0] ));
 sg13g2_inv_1 _5486_ (.Y(_0312_),
    .A(net353));
 sg13g2_a22oi_1 _5487_ (.Y(_1947_),
    .B1(_1945_),
    .B2(net368),
    .A2(net605),
    .A1(\core.byte_acc[1] ));
 sg13g2_inv_1 _5488_ (.Y(_0313_),
    .A(net369));
 sg13g2_a22oi_1 _5489_ (.Y(_0314_),
    .B1(_1945_),
    .B2(_2714_),
    .A2(net605),
    .A1(_2626_));
 sg13g2_a22oi_1 _5490_ (.Y(_1948_),
    .B1(_1945_),
    .B2(net346),
    .A2(net605),
    .A1(\core.byte_acc[3] ));
 sg13g2_inv_1 _5491_ (.Y(_0315_),
    .A(net347));
 sg13g2_a22oi_1 _5492_ (.Y(_1949_),
    .B1(_1945_),
    .B2(net378),
    .A2(net605),
    .A1(\core.byte_acc[4] ));
 sg13g2_inv_1 _5493_ (.Y(_0316_),
    .A(net379));
 sg13g2_a22oi_1 _5494_ (.Y(_0317_),
    .B1(_1945_),
    .B2(_2710_),
    .A2(_1944_),
    .A1(_2624_));
 sg13g2_a22oi_1 _5495_ (.Y(_0318_),
    .B1(_1945_),
    .B2(_2708_),
    .A2(net605),
    .A1(_2623_));
 sg13g2_a22oi_1 _5496_ (.Y(_0319_),
    .B1(_1945_),
    .B2(_2706_),
    .A2(net605),
    .A1(_2622_));
 sg13g2_or3_1 _5497_ (.A(_2721_),
    .B(_2742_),
    .C(_2752_),
    .X(_1950_));
 sg13g2_nand2_1 _5498_ (.Y(_1951_),
    .A(\core.temp_q[15] ),
    .B(\core.temp_q[14] ));
 sg13g2_nand4_1 _5499_ (.B(\core.temp_q[12] ),
    .C(\core.temp_q[11] ),
    .A(\core.temp_q[13] ),
    .Y(_1952_),
    .D(\core.temp_q[10] ));
 sg13g2_nor2_1 _5500_ (.A(_1951_),
    .B(_1952_),
    .Y(_1953_));
 sg13g2_nor4_2 _5501_ (.A(\core.temp_q[3] ),
    .B(\core.temp_q[2] ),
    .C(\core.temp_q[1] ),
    .Y(_1954_),
    .D(\core.temp_q[0] ));
 sg13g2_nor4_1 _5502_ (.A(\core.temp_q[7] ),
    .B(\core.temp_q[6] ),
    .C(\core.temp_q[5] ),
    .D(\core.temp_q[4] ),
    .Y(_1955_));
 sg13g2_nand4_1 _5503_ (.B(_2652_),
    .C(_1954_),
    .A(_2651_),
    .Y(_1956_),
    .D(_1955_));
 sg13g2_a21oi_2 _5504_ (.B1(_2650_),
    .Y(_1957_),
    .A2(_1956_),
    .A1(_1953_));
 sg13g2_a21o_2 _5505_ (.A2(_1956_),
    .A1(_1953_),
    .B1(_2650_),
    .X(_1958_));
 sg13g2_nor2_1 _5506_ (.A(\core.temp_q[14] ),
    .B(\core.temp_q[13] ),
    .Y(_1959_));
 sg13g2_nor3_1 _5507_ (.A(\core.temp_q[12] ),
    .B(\core.temp_q[11] ),
    .C(\core.temp_q[10] ),
    .Y(_1960_));
 sg13g2_a21oi_2 _5508_ (.B1(\core.temp_q[15] ),
    .Y(_1961_),
    .A2(_1960_),
    .A1(_1959_));
 sg13g2_a21o_2 _5509_ (.A2(_1960_),
    .A1(_1959_),
    .B1(\core.temp_q[15] ),
    .X(_1962_));
 sg13g2_o21ai_1 _5510_ (.B1(_0008_),
    .Y(_1963_),
    .A1(_1951_),
    .A2(_1952_));
 sg13g2_or3_1 _5511_ (.A(_0008_),
    .B(_1951_),
    .C(_1952_),
    .X(_1964_));
 sg13g2_a21oi_2 _5512_ (.B1(_2652_),
    .Y(_1965_),
    .A2(_1964_),
    .A1(_1963_));
 sg13g2_or2_1 _5513_ (.X(_1966_),
    .B(_1965_),
    .A(_1961_));
 sg13g2_o21ai_1 _5514_ (.B1(_1958_),
    .Y(_1967_),
    .A1(_1961_),
    .A2(_1965_));
 sg13g2_o21ai_1 _5515_ (.B1(_1962_),
    .Y(_1968_),
    .A1(\core.temp_q[10] ),
    .A2(_2725_));
 sg13g2_a21o_1 _5516_ (.A2(_1964_),
    .A1(_1963_),
    .B1(_0007_),
    .X(_1969_));
 sg13g2_and2_1 _5517_ (.A(_1962_),
    .B(_1969_),
    .X(_1970_));
 sg13g2_nand2_1 _5518_ (.Y(_1971_),
    .A(_1962_),
    .B(_1969_));
 sg13g2_a21o_1 _5519_ (.A2(_1964_),
    .A1(_1963_),
    .B1(_2651_),
    .X(_1972_));
 sg13g2_and2_1 _5520_ (.A(_1962_),
    .B(_1972_),
    .X(_1973_));
 sg13g2_a21oi_2 _5521_ (.B1(_1957_),
    .Y(_1974_),
    .A2(_1972_),
    .A1(_1962_));
 sg13g2_a21o_2 _5522_ (.A2(_1972_),
    .A1(_1962_),
    .B1(_1957_),
    .X(_1975_));
 sg13g2_a21o_2 _5523_ (.A2(_1969_),
    .A1(_1962_),
    .B1(_1957_),
    .X(_1976_));
 sg13g2_nand2_1 _5524_ (.Y(_1977_),
    .A(_1971_),
    .B(_1974_));
 sg13g2_nor3_1 _5525_ (.A(_1968_),
    .B(_1970_),
    .C(_1975_),
    .Y(_1978_));
 sg13g2_and2_2 _5526_ (.A(_1958_),
    .B(_1968_),
    .X(_1979_));
 sg13g2_nand2_2 _5527_ (.Y(_1980_),
    .A(_1958_),
    .B(_1968_));
 sg13g2_and3_1 _5528_ (.X(_1981_),
    .A(_1975_),
    .B(_1976_),
    .C(net618));
 sg13g2_nor2_1 _5529_ (.A(_1978_),
    .B(_1981_),
    .Y(_1982_));
 sg13g2_o21ai_1 _5530_ (.B1(_1967_),
    .Y(_1983_),
    .A1(_1978_),
    .A2(_1981_));
 sg13g2_nand2b_1 _5531_ (.Y(_1984_),
    .B(_1973_),
    .A_N(_1967_));
 sg13g2_nand2_1 _5532_ (.Y(_1985_),
    .A(_1970_),
    .B(_1979_));
 sg13g2_or2_2 _5533_ (.X(_1986_),
    .B(_1985_),
    .A(_1984_));
 sg13g2_nand4_1 _5534_ (.B(_1962_),
    .C(_1965_),
    .A(_1958_),
    .Y(_1987_),
    .D(_1969_));
 sg13g2_and2_1 _5535_ (.A(_1973_),
    .B(_1979_),
    .X(_1988_));
 sg13g2_nand2_1 _5536_ (.Y(_1989_),
    .A(_1973_),
    .B(_1979_));
 sg13g2_and2_1 _5537_ (.A(_1983_),
    .B(_1986_),
    .X(_1990_));
 sg13g2_nand2_1 _5538_ (.Y(_1991_),
    .A(net683),
    .B(net590));
 sg13g2_nand3b_1 _5539_ (.B(\core.compute_state[2] ),
    .C(net739),
    .Y(_1992_),
    .A_N(_2752_));
 sg13g2_inv_1 _5540_ (.Y(_1993_),
    .A(net596));
 sg13g2_nor2_1 _5541_ (.A(_1991_),
    .B(net596),
    .Y(_1994_));
 sg13g2_a21oi_1 _5542_ (.A1(net776),
    .A2(net599),
    .Y(_1995_),
    .B1(_1994_));
 sg13g2_nor2_1 _5543_ (.A(net720),
    .B(_1995_),
    .Y(_0320_));
 sg13g2_nor2_1 _5544_ (.A(_1966_),
    .B(_1976_),
    .Y(_1996_));
 sg13g2_or2_1 _5545_ (.X(_1997_),
    .B(_1976_),
    .A(_1966_));
 sg13g2_nand2_1 _5546_ (.Y(_1998_),
    .A(_1975_),
    .B(_1987_));
 sg13g2_nor4_2 _5547_ (.A(_1957_),
    .B(_1961_),
    .C(_1965_),
    .Y(_1999_),
    .D(_1972_));
 sg13g2_nand2_1 _5548_ (.Y(_2000_),
    .A(_1976_),
    .B(_1999_));
 sg13g2_a22oi_1 _5549_ (.Y(_2001_),
    .B1(_1999_),
    .B2(_1976_),
    .A2(_1987_),
    .A1(_1975_));
 sg13g2_o21ai_1 _5550_ (.B1(net618),
    .Y(_2002_),
    .A1(_1996_),
    .A2(_2001_));
 sg13g2_xor2_1 _5551_ (.B(net682),
    .A(\core.delta_t[9] ),
    .X(_2003_));
 sg13g2_nor2_1 _5552_ (.A(net680),
    .B(_0009_),
    .Y(_2004_));
 sg13g2_a21o_1 _5553_ (.A2(_2003_),
    .A1(net680),
    .B1(_2004_),
    .X(_2005_));
 sg13g2_a21oi_2 _5554_ (.B1(_2004_),
    .Y(_2006_),
    .A2(_2003_),
    .A1(net680));
 sg13g2_nand2_1 _5555_ (.Y(_2007_),
    .A(net595),
    .B(net623));
 sg13g2_nand2_1 _5556_ (.Y(_2008_),
    .A(net590),
    .B(net623));
 sg13g2_nor2_1 _5557_ (.A(_1991_),
    .B(_2007_),
    .Y(_2009_));
 sg13g2_a22oi_1 _5558_ (.Y(_2010_),
    .B1(net623),
    .B2(net590),
    .A2(net595),
    .A1(net683));
 sg13g2_or2_1 _5559_ (.X(_2011_),
    .B(_2010_),
    .A(_2009_));
 sg13g2_nor2_1 _5560_ (.A(net596),
    .B(_2011_),
    .Y(_2012_));
 sg13g2_a21oi_1 _5561_ (.A1(net794),
    .A2(net598),
    .Y(_2013_),
    .B1(_2012_));
 sg13g2_nor2_1 _5562_ (.A(net720),
    .B(_2013_),
    .Y(_0321_));
 sg13g2_nand3_1 _5563_ (.B(_1984_),
    .C(_1985_),
    .A(_1977_),
    .Y(_2014_));
 sg13g2_and2_2 _5564_ (.A(_1986_),
    .B(_2014_),
    .X(_2015_));
 sg13g2_nand2_1 _5565_ (.Y(_2016_),
    .A(_1986_),
    .B(_2014_));
 sg13g2_nand2_1 _5566_ (.Y(_2017_),
    .A(net683),
    .B(_2015_));
 sg13g2_nand2_1 _5567_ (.Y(_2018_),
    .A(net620),
    .B(net595));
 sg13g2_nand2_1 _5568_ (.Y(_2019_),
    .A(net620),
    .B(net590));
 sg13g2_or2_1 _5569_ (.X(_2020_),
    .B(_2018_),
    .A(_2008_));
 sg13g2_and2_1 _5570_ (.A(_2007_),
    .B(_2019_),
    .X(_2021_));
 sg13g2_xor2_1 _5571_ (.B(_2019_),
    .A(_2007_),
    .X(_2022_));
 sg13g2_xnor2_1 _5572_ (.Y(_2023_),
    .A(_2017_),
    .B(_2022_));
 sg13g2_nand2_1 _5573_ (.Y(_2024_),
    .A(_2009_),
    .B(_2023_));
 sg13g2_xor2_1 _5574_ (.B(_2023_),
    .A(_2009_),
    .X(_2025_));
 sg13g2_inv_1 _5575_ (.Y(_2026_),
    .A(_2025_));
 sg13g2_nand2b_1 _5576_ (.Y(_2027_),
    .B(_2025_),
    .A_N(_1991_));
 sg13g2_a21o_1 _5577_ (.A2(_2023_),
    .A1(_1993_),
    .B1(_1994_),
    .X(_2028_));
 sg13g2_a22oi_1 _5578_ (.Y(_2029_),
    .B1(_2027_),
    .B2(_2028_),
    .A2(net598),
    .A1(net792));
 sg13g2_nor2_1 _5579_ (.A(net719),
    .B(_2029_),
    .Y(_0322_));
 sg13g2_o21ai_1 _5580_ (.B1(_2020_),
    .Y(_2030_),
    .A1(_2017_),
    .A2(_2021_));
 sg13g2_nand3_1 _5581_ (.B(_1980_),
    .C(_1997_),
    .A(_1974_),
    .Y(_2031_));
 sg13g2_nand2_1 _5582_ (.Y(_2032_),
    .A(_1967_),
    .B(_1976_));
 sg13g2_a21oi_2 _5583_ (.B1(net618),
    .Y(_2033_),
    .A2(_1976_),
    .A1(_1967_));
 sg13g2_o21ai_1 _5584_ (.B1(_2031_),
    .Y(_2034_),
    .A1(_1979_),
    .A2(_1984_));
 sg13g2_a21o_2 _5585_ (.A2(_2033_),
    .A1(_1984_),
    .B1(_2034_),
    .X(_2035_));
 sg13g2_nor2b_1 _5586_ (.A(_0012_),
    .B_N(_2035_),
    .Y(_2036_));
 sg13g2_nand2_1 _5587_ (.Y(_2037_),
    .A(_2030_),
    .B(_2036_));
 sg13g2_xnor2_1 _5588_ (.Y(_2038_),
    .A(_2030_),
    .B(_2036_));
 sg13g2_nor2_2 _5589_ (.A(_2006_),
    .B(_2016_),
    .Y(_2039_));
 sg13g2_nand2_1 _5590_ (.Y(_2040_),
    .A(net619),
    .B(net595));
 sg13g2_nand2_1 _5591_ (.Y(_2041_),
    .A(net619),
    .B(net590));
 sg13g2_nor2_1 _5592_ (.A(_2019_),
    .B(_2040_),
    .Y(_2042_));
 sg13g2_xor2_1 _5593_ (.B(_2041_),
    .A(_2018_),
    .X(_2043_));
 sg13g2_xnor2_1 _5594_ (.Y(_2044_),
    .A(_2039_),
    .B(_2043_));
 sg13g2_nor2_1 _5595_ (.A(_2038_),
    .B(_2044_),
    .Y(_2045_));
 sg13g2_xor2_1 _5596_ (.B(_2044_),
    .A(_2038_),
    .X(_2046_));
 sg13g2_nor2b_1 _5597_ (.A(_2011_),
    .B_N(_2046_),
    .Y(_2047_));
 sg13g2_nor2b_1 _5598_ (.A(_2024_),
    .B_N(_2046_),
    .Y(_2048_));
 sg13g2_xor2_1 _5599_ (.B(_2046_),
    .A(_2024_),
    .X(_2049_));
 sg13g2_inv_1 _5600_ (.Y(_2050_),
    .A(_2049_));
 sg13g2_a21oi_1 _5601_ (.A1(_2011_),
    .A2(_2049_),
    .Y(_2051_),
    .B1(_2047_));
 sg13g2_inv_1 _5602_ (.Y(_2052_),
    .A(_2051_));
 sg13g2_nor2b_1 _5603_ (.A(_2027_),
    .B_N(_2051_),
    .Y(_2053_));
 sg13g2_nand2_1 _5604_ (.Y(_2054_),
    .A(_2027_),
    .B(_2052_));
 sg13g2_nor2_1 _5605_ (.A(net596),
    .B(_2053_),
    .Y(_2055_));
 sg13g2_a22oi_1 _5606_ (.Y(_2056_),
    .B1(_2054_),
    .B2(_2055_),
    .A2(net598),
    .A1(net777));
 sg13g2_nor2_1 _5607_ (.A(net719),
    .B(_2056_),
    .Y(_0323_));
 sg13g2_or2_1 _5608_ (.X(_2057_),
    .B(_2053_),
    .A(_2047_));
 sg13g2_a21oi_1 _5609_ (.A1(_2039_),
    .A2(_2043_),
    .Y(_2058_),
    .B1(_2042_));
 sg13g2_nand2_1 _5610_ (.Y(_2059_),
    .A(net623),
    .B(_2035_));
 sg13g2_nor2_1 _5611_ (.A(_2058_),
    .B(_2059_),
    .Y(_2060_));
 sg13g2_xor2_1 _5612_ (.B(_2059_),
    .A(_2058_),
    .X(_2061_));
 sg13g2_nand2_1 _5613_ (.Y(_2062_),
    .A(net620),
    .B(_2015_));
 sg13g2_nand2_1 _5614_ (.Y(_2063_),
    .A(net613),
    .B(_2002_));
 sg13g2_nand3_1 _5615_ (.B(_1983_),
    .C(_1986_),
    .A(net613),
    .Y(_2064_));
 sg13g2_or2_1 _5616_ (.X(_2065_),
    .B(_2064_),
    .A(_2040_));
 sg13g2_xor2_1 _5617_ (.B(_2064_),
    .A(_2040_),
    .X(_2066_));
 sg13g2_nand2b_1 _5618_ (.Y(_2067_),
    .B(_2066_),
    .A_N(_2062_));
 sg13g2_xor2_1 _5619_ (.B(_2066_),
    .A(_2062_),
    .X(_2068_));
 sg13g2_o21ai_1 _5620_ (.B1(_1967_),
    .Y(_2069_),
    .A1(_0007_),
    .A2(_1975_));
 sg13g2_inv_1 _5621_ (.Y(_2070_),
    .A(_2069_));
 sg13g2_o21ai_1 _5622_ (.B1(_1982_),
    .Y(_2071_),
    .A1(net618),
    .A2(_2070_));
 sg13g2_nor2b_1 _5623_ (.A(_0012_),
    .B_N(_2071_),
    .Y(_2072_));
 sg13g2_nand2b_1 _5624_ (.Y(_2073_),
    .B(_2072_),
    .A_N(_2068_));
 sg13g2_xnor2_1 _5625_ (.Y(_2074_),
    .A(_2068_),
    .B(_2072_));
 sg13g2_nand2_1 _5626_ (.Y(_2075_),
    .A(_2061_),
    .B(_2074_));
 sg13g2_xnor2_1 _5627_ (.Y(_2076_),
    .A(_2061_),
    .B(_2074_));
 sg13g2_or3_1 _5628_ (.A(_2038_),
    .B(_2044_),
    .C(_2076_),
    .X(_2077_));
 sg13g2_xor2_1 _5629_ (.B(_2076_),
    .A(_2045_),
    .X(_2078_));
 sg13g2_xor2_1 _5630_ (.B(_2078_),
    .A(_2037_),
    .X(_2079_));
 sg13g2_nand2_1 _5631_ (.Y(_2080_),
    .A(_2048_),
    .B(_2079_));
 sg13g2_xnor2_1 _5632_ (.Y(_2081_),
    .A(_2048_),
    .B(_2079_));
 sg13g2_nor2_1 _5633_ (.A(_2026_),
    .B(_2081_),
    .Y(_2082_));
 sg13g2_xnor2_1 _5634_ (.Y(_2083_),
    .A(_2025_),
    .B(_2081_));
 sg13g2_and2_1 _5635_ (.A(_2057_),
    .B(_2083_),
    .X(_2084_));
 sg13g2_o21ai_1 _5636_ (.B1(_1993_),
    .Y(_2085_),
    .A1(_2057_),
    .A2(_2083_));
 sg13g2_nor2_1 _5637_ (.A(_2084_),
    .B(_2085_),
    .Y(_2086_));
 sg13g2_a21oi_1 _5638_ (.A1(net805),
    .A2(net598),
    .Y(_2087_),
    .B1(_2086_));
 sg13g2_nor2_1 _5639_ (.A(net719),
    .B(_2087_),
    .Y(_0324_));
 sg13g2_o21ai_1 _5640_ (.B1(_2077_),
    .Y(_2088_),
    .A1(_2037_),
    .A2(_2078_));
 sg13g2_nand2_1 _5641_ (.Y(_2089_),
    .A(net620),
    .B(_2035_));
 sg13g2_a21oi_2 _5642_ (.B1(_2089_),
    .Y(_2090_),
    .A2(_2067_),
    .A1(_2065_));
 sg13g2_nand3_1 _5643_ (.B(_2067_),
    .C(_2089_),
    .A(_2065_),
    .Y(_2091_));
 sg13g2_nor2b_1 _5644_ (.A(_2090_),
    .B_N(_2091_),
    .Y(_2092_));
 sg13g2_nand2_1 _5645_ (.Y(_2093_),
    .A(net623),
    .B(_2071_));
 sg13g2_nand4_1 _5646_ (.B(_1966_),
    .C(_1971_),
    .A(_1958_),
    .Y(_2094_),
    .D(_1974_));
 sg13g2_and3_1 _5647_ (.X(_2095_),
    .A(_2651_),
    .B(_2032_),
    .C(_2094_));
 sg13g2_nand3_1 _5648_ (.B(_2032_),
    .C(_2094_),
    .A(net618),
    .Y(_2096_));
 sg13g2_o21ai_1 _5649_ (.B1(_2096_),
    .Y(_2097_),
    .A1(net618),
    .A2(_2095_));
 sg13g2_nand2_1 _5650_ (.Y(_2098_),
    .A(net683),
    .B(net588));
 sg13g2_nor2_1 _5651_ (.A(_2093_),
    .B(_2098_),
    .Y(_2099_));
 sg13g2_xor2_1 _5652_ (.B(_2098_),
    .A(_2093_),
    .X(_2100_));
 sg13g2_inv_1 _5653_ (.Y(_2101_),
    .A(_2100_));
 sg13g2_nor2_2 _5654_ (.A(_0575_),
    .B(_2016_),
    .Y(_2102_));
 sg13g2_nand2_1 _5655_ (.Y(_2103_),
    .A(net600),
    .B(net595));
 sg13g2_nand3_1 _5656_ (.B(_1983_),
    .C(_1986_),
    .A(net600),
    .Y(_2104_));
 sg13g2_nor2_1 _5657_ (.A(_2064_),
    .B(_2103_),
    .Y(_2105_));
 sg13g2_xor2_1 _5658_ (.B(_2104_),
    .A(_2063_),
    .X(_2106_));
 sg13g2_xnor2_1 _5659_ (.Y(_2107_),
    .A(_2102_),
    .B(_2106_));
 sg13g2_nor2_1 _5660_ (.A(_2101_),
    .B(_2107_),
    .Y(_2108_));
 sg13g2_xor2_1 _5661_ (.B(_2107_),
    .A(_2100_),
    .X(_2109_));
 sg13g2_xor2_1 _5662_ (.B(_2109_),
    .A(_2073_),
    .X(_2110_));
 sg13g2_nand2_1 _5663_ (.Y(_2111_),
    .A(_2092_),
    .B(_2110_));
 sg13g2_xnor2_1 _5664_ (.Y(_2112_),
    .A(_2092_),
    .B(_2110_));
 sg13g2_nor2_1 _5665_ (.A(_2075_),
    .B(_2112_),
    .Y(_2113_));
 sg13g2_xor2_1 _5666_ (.B(_2112_),
    .A(_2075_),
    .X(_2114_));
 sg13g2_xnor2_1 _5667_ (.Y(_2115_),
    .A(_2060_),
    .B(_2114_));
 sg13g2_nand2b_1 _5668_ (.Y(_2116_),
    .B(_2088_),
    .A_N(_2115_));
 sg13g2_xor2_1 _5669_ (.B(_2115_),
    .A(_2088_),
    .X(_2117_));
 sg13g2_or2_1 _5670_ (.X(_2118_),
    .B(_2117_),
    .A(_2049_));
 sg13g2_xor2_1 _5671_ (.B(_2117_),
    .A(_2080_),
    .X(_2119_));
 sg13g2_o21ai_1 _5672_ (.B1(_2118_),
    .Y(_2120_),
    .A1(_2050_),
    .A2(_2119_));
 sg13g2_nor2_1 _5673_ (.A(_2082_),
    .B(_2084_),
    .Y(_2121_));
 sg13g2_or2_1 _5674_ (.X(_2122_),
    .B(_2121_),
    .A(_2120_));
 sg13g2_a21oi_1 _5675_ (.A1(_2120_),
    .A2(_2121_),
    .Y(_2123_),
    .B1(net596));
 sg13g2_a22oi_1 _5676_ (.Y(_2124_),
    .B1(_2122_),
    .B2(_2123_),
    .A2(net598),
    .A1(net787));
 sg13g2_nor2_1 _5677_ (.A(net719),
    .B(_2124_),
    .Y(_0325_));
 sg13g2_nand2_1 _5678_ (.Y(_2125_),
    .A(net531),
    .B(net598));
 sg13g2_o21ai_1 _5679_ (.B1(_2116_),
    .Y(_2126_),
    .A1(_2080_),
    .A2(_2117_));
 sg13g2_a21oi_1 _5680_ (.A1(_2060_),
    .A2(_2114_),
    .Y(_2127_),
    .B1(_2113_));
 sg13g2_and2_1 _5681_ (.A(net613),
    .B(_2015_),
    .X(_2128_));
 sg13g2_nand2_2 _5682_ (.Y(_2129_),
    .A(net593),
    .B(_1990_));
 sg13g2_nor2_1 _5683_ (.A(_2103_),
    .B(_2129_),
    .Y(_2130_));
 sg13g2_xor2_1 _5684_ (.B(_2129_),
    .A(_2103_),
    .X(_2131_));
 sg13g2_xor2_1 _5685_ (.B(_2131_),
    .A(_2128_),
    .X(_2132_));
 sg13g2_nand2_1 _5686_ (.Y(_2133_),
    .A(net620),
    .B(_2071_));
 sg13g2_mux2_1 _5687_ (.A0(_1975_),
    .A1(_1976_),
    .S(_1966_),
    .X(_2134_));
 sg13g2_mux2_2 _5688_ (.A0(_1989_),
    .A1(_1979_),
    .S(_2134_),
    .X(_2135_));
 sg13g2_mux2_2 _5689_ (.A0(_1988_),
    .A1(net618),
    .S(_2134_),
    .X(_2136_));
 sg13g2_nor2_1 _5690_ (.A(_0012_),
    .B(_2136_),
    .Y(_2137_));
 sg13g2_and3_1 _5691_ (.X(_2138_),
    .A(net623),
    .B(net588),
    .C(_2137_));
 sg13g2_a21oi_1 _5692_ (.A1(net623),
    .A2(net588),
    .Y(_2139_),
    .B1(_2137_));
 sg13g2_or3_1 _5693_ (.A(_2133_),
    .B(_2138_),
    .C(_2139_),
    .X(_2140_));
 sg13g2_o21ai_1 _5694_ (.B1(_2133_),
    .Y(_2141_),
    .A1(_2138_),
    .A2(_2139_));
 sg13g2_nand3_1 _5695_ (.B(_2140_),
    .C(_2141_),
    .A(_2099_),
    .Y(_2142_));
 sg13g2_a21o_1 _5696_ (.A2(_2141_),
    .A1(_2140_),
    .B1(_2099_),
    .X(_2143_));
 sg13g2_and2_1 _5697_ (.A(_2142_),
    .B(_2143_),
    .X(_2144_));
 sg13g2_nand3_1 _5698_ (.B(_2142_),
    .C(_2143_),
    .A(_2132_),
    .Y(_2145_));
 sg13g2_a21oi_1 _5699_ (.A1(_2142_),
    .A2(_2143_),
    .Y(_2146_),
    .B1(_2132_));
 sg13g2_xor2_1 _5700_ (.B(_2144_),
    .A(_2132_),
    .X(_2147_));
 sg13g2_nand3b_1 _5701_ (.B(_2108_),
    .C(_2145_),
    .Y(_2148_),
    .A_N(_2146_));
 sg13g2_xnor2_1 _5702_ (.Y(_2149_),
    .A(_2108_),
    .B(_2147_));
 sg13g2_and2_1 _5703_ (.A(net619),
    .B(_2035_),
    .X(_2150_));
 sg13g2_a21oi_1 _5704_ (.A1(_2102_),
    .A2(_2106_),
    .Y(_2151_),
    .B1(_2105_));
 sg13g2_nor3_1 _5705_ (.A(_2073_),
    .B(_2109_),
    .C(_2151_),
    .Y(_2152_));
 sg13g2_o21ai_1 _5706_ (.B1(_2151_),
    .Y(_2153_),
    .A1(_2073_),
    .A2(_2109_));
 sg13g2_nor2b_1 _5707_ (.A(_2152_),
    .B_N(_2153_),
    .Y(_2154_));
 sg13g2_xnor2_1 _5708_ (.Y(_2155_),
    .A(_2150_),
    .B(_2154_));
 sg13g2_nor2_1 _5709_ (.A(_2149_),
    .B(_2155_),
    .Y(_2156_));
 sg13g2_xnor2_1 _5710_ (.Y(_2157_),
    .A(_2149_),
    .B(_2155_));
 sg13g2_nor2_1 _5711_ (.A(_2111_),
    .B(_2157_),
    .Y(_2158_));
 sg13g2_xor2_1 _5712_ (.B(_2157_),
    .A(_2111_),
    .X(_2159_));
 sg13g2_xnor2_1 _5713_ (.Y(_2160_),
    .A(_2090_),
    .B(_2159_));
 sg13g2_nor2_1 _5714_ (.A(_2127_),
    .B(_2160_),
    .Y(_2161_));
 sg13g2_xor2_1 _5715_ (.B(_2160_),
    .A(_2127_),
    .X(_2162_));
 sg13g2_xnor2_1 _5716_ (.Y(_2163_),
    .A(_2126_),
    .B(_2162_));
 sg13g2_or2_1 _5717_ (.X(_2164_),
    .B(_2163_),
    .A(_2081_));
 sg13g2_nand2_1 _5718_ (.Y(_2165_),
    .A(_2081_),
    .B(_2163_));
 sg13g2_and2_1 _5719_ (.A(_2164_),
    .B(_2165_),
    .X(_2166_));
 sg13g2_nand2_1 _5720_ (.Y(_2167_),
    .A(_2118_),
    .B(_2122_));
 sg13g2_nand2_1 _5721_ (.Y(_2168_),
    .A(_2166_),
    .B(_2167_));
 sg13g2_o21ai_1 _5722_ (.B1(_1993_),
    .Y(_2169_),
    .A1(_2166_),
    .A2(_2167_));
 sg13g2_nand2b_1 _5723_ (.Y(_2170_),
    .B(_2168_),
    .A_N(_2169_));
 sg13g2_a21oi_1 _5724_ (.A1(_2125_),
    .A2(_2170_),
    .Y(_0326_),
    .B1(net720));
 sg13g2_a21oi_1 _5725_ (.A1(_2126_),
    .A2(_2162_),
    .Y(_2171_),
    .B1(_2161_));
 sg13g2_a21oi_1 _5726_ (.A1(_2090_),
    .A2(_2159_),
    .Y(_2172_),
    .B1(_2158_));
 sg13g2_a21oi_1 _5727_ (.A1(_2150_),
    .A2(_2153_),
    .Y(_2173_),
    .B1(_2152_));
 sg13g2_nand2_1 _5728_ (.Y(_2174_),
    .A(_2142_),
    .B(_2145_));
 sg13g2_nand2_1 _5729_ (.Y(_2175_),
    .A(net600),
    .B(_2015_));
 sg13g2_inv_1 _5730_ (.Y(_2176_),
    .A(_2175_));
 sg13g2_nand2_1 _5731_ (.Y(_2177_),
    .A(net611),
    .B(net595));
 sg13g2_nor2_1 _5732_ (.A(_2129_),
    .B(_2177_),
    .Y(_2178_));
 sg13g2_nand2_1 _5733_ (.Y(_2179_),
    .A(net611),
    .B(net590));
 sg13g2_a22oi_1 _5734_ (.Y(_2180_),
    .B1(net595),
    .B2(net593),
    .A2(net590),
    .A1(net611));
 sg13g2_nor2_1 _5735_ (.A(_2178_),
    .B(_2180_),
    .Y(_2181_));
 sg13g2_xnor2_1 _5736_ (.Y(_2182_),
    .A(_2176_),
    .B(_2181_));
 sg13g2_nand2b_1 _5737_ (.Y(_2183_),
    .B(_2140_),
    .A_N(_2138_));
 sg13g2_nand2_1 _5738_ (.Y(_2184_),
    .A(net619),
    .B(_2071_));
 sg13g2_nand2_1 _5739_ (.Y(_2185_),
    .A(net620),
    .B(_2135_));
 sg13g2_nand2_1 _5740_ (.Y(_2186_),
    .A(net621),
    .B(net588));
 sg13g2_nor2_1 _5741_ (.A(_2006_),
    .B(_2136_),
    .Y(_2187_));
 sg13g2_nand3_1 _5742_ (.B(net588),
    .C(_2187_),
    .A(net620),
    .Y(_2188_));
 sg13g2_a21oi_1 _5743_ (.A1(net620),
    .A2(net588),
    .Y(_2189_),
    .B1(_2187_));
 sg13g2_xnor2_1 _5744_ (.Y(_2190_),
    .A(_2186_),
    .B(_2187_));
 sg13g2_xnor2_1 _5745_ (.Y(_2191_),
    .A(_2184_),
    .B(_2190_));
 sg13g2_nand2_1 _5746_ (.Y(_2192_),
    .A(_2183_),
    .B(_2191_));
 sg13g2_xnor2_1 _5747_ (.Y(_2193_),
    .A(_2183_),
    .B(_2191_));
 sg13g2_xnor2_1 _5748_ (.Y(_2194_),
    .A(_2182_),
    .B(_2193_));
 sg13g2_nand2b_1 _5749_ (.Y(_2195_),
    .B(_2174_),
    .A_N(_2194_));
 sg13g2_xnor2_1 _5750_ (.Y(_2196_),
    .A(_2174_),
    .B(_2194_));
 sg13g2_a21oi_1 _5751_ (.A1(_1968_),
    .A2(_1974_),
    .Y(_2197_),
    .B1(_1997_));
 sg13g2_a21oi_2 _5752_ (.B1(_2197_),
    .Y(_2198_),
    .A2(_1980_),
    .A1(_1975_));
 sg13g2_nand2_1 _5753_ (.Y(_2199_),
    .A(net683),
    .B(net587));
 sg13g2_nand3_1 _5754_ (.B(_2196_),
    .C(net587),
    .A(net683),
    .Y(_2200_));
 sg13g2_xor2_1 _5755_ (.B(_2199_),
    .A(_2196_),
    .X(_2201_));
 sg13g2_nand2_1 _5756_ (.Y(_2202_),
    .A(net613),
    .B(_2035_));
 sg13g2_a21oi_1 _5757_ (.A1(_2128_),
    .A2(_2131_),
    .Y(_2203_),
    .B1(_2130_));
 sg13g2_nor2_1 _5758_ (.A(_2148_),
    .B(_2203_),
    .Y(_2204_));
 sg13g2_xnor2_1 _5759_ (.Y(_2205_),
    .A(_2148_),
    .B(_2203_));
 sg13g2_nor2_1 _5760_ (.A(_2202_),
    .B(_2205_),
    .Y(_2206_));
 sg13g2_xnor2_1 _5761_ (.Y(_2207_),
    .A(_2202_),
    .B(_2205_));
 sg13g2_nor2_1 _5762_ (.A(_2201_),
    .B(_2207_),
    .Y(_2208_));
 sg13g2_xor2_1 _5763_ (.B(_2207_),
    .A(_2201_),
    .X(_2209_));
 sg13g2_nand2_1 _5764_ (.Y(_2210_),
    .A(_2156_),
    .B(_2209_));
 sg13g2_xnor2_1 _5765_ (.Y(_2211_),
    .A(_2156_),
    .B(_2209_));
 sg13g2_xor2_1 _5766_ (.B(_2211_),
    .A(_2173_),
    .X(_2212_));
 sg13g2_nand2b_1 _5767_ (.Y(_2213_),
    .B(_2212_),
    .A_N(_2172_));
 sg13g2_nor2b_1 _5768_ (.A(_2212_),
    .B_N(_2172_),
    .Y(_2214_));
 sg13g2_xnor2_1 _5769_ (.Y(_2215_),
    .A(_2172_),
    .B(_2212_));
 sg13g2_xnor2_1 _5770_ (.Y(_2216_),
    .A(_2171_),
    .B(_2215_));
 sg13g2_nand2_1 _5771_ (.Y(_2217_),
    .A(_2119_),
    .B(_2216_));
 sg13g2_xor2_1 _5772_ (.B(_2216_),
    .A(_2119_),
    .X(_2218_));
 sg13g2_xnor2_1 _5773_ (.Y(_2219_),
    .A(_2119_),
    .B(_2216_));
 sg13g2_xnor2_1 _5774_ (.Y(_2220_),
    .A(_2164_),
    .B(_2219_));
 sg13g2_nand4_1 _5775_ (.B(_2165_),
    .C(_2167_),
    .A(_2164_),
    .Y(_2221_),
    .D(_2218_));
 sg13g2_a21oi_1 _5776_ (.A1(_2168_),
    .A2(_2220_),
    .Y(_2222_),
    .B1(net596));
 sg13g2_a22oi_1 _5777_ (.Y(_2223_),
    .B1(_2221_),
    .B2(_2222_),
    .A2(net598),
    .A1(net765));
 sg13g2_nor2_1 _5778_ (.A(net719),
    .B(_2223_),
    .Y(_0327_));
 sg13g2_nand2_1 _5779_ (.Y(_2224_),
    .A(net514),
    .B(net598));
 sg13g2_o21ai_1 _5780_ (.B1(_2221_),
    .Y(_2225_),
    .A1(_2164_),
    .A2(_2219_));
 sg13g2_o21ai_1 _5781_ (.B1(_2213_),
    .Y(_2226_),
    .A1(_2171_),
    .A2(_2214_));
 sg13g2_o21ai_1 _5782_ (.B1(_2210_),
    .Y(_2227_),
    .A1(_2173_),
    .A2(_2211_));
 sg13g2_nor2_1 _5783_ (.A(_2204_),
    .B(_2206_),
    .Y(_2228_));
 sg13g2_nand2_1 _5784_ (.Y(_2229_),
    .A(net600),
    .B(_2035_));
 sg13g2_a21oi_1 _5785_ (.A1(_2176_),
    .A2(_2181_),
    .Y(_2230_),
    .B1(_2178_));
 sg13g2_nor2_1 _5786_ (.A(_2195_),
    .B(_2230_),
    .Y(_2231_));
 sg13g2_xnor2_1 _5787_ (.Y(_2232_),
    .A(_2195_),
    .B(_2230_));
 sg13g2_nor2_1 _5788_ (.A(_2229_),
    .B(_2232_),
    .Y(_2233_));
 sg13g2_xnor2_1 _5789_ (.Y(_2234_),
    .A(_2229_),
    .B(_2232_));
 sg13g2_inv_1 _5790_ (.Y(_2235_),
    .A(_2234_));
 sg13g2_o21ai_1 _5791_ (.B1(_2192_),
    .Y(_2236_),
    .A1(_2182_),
    .A2(_2193_));
 sg13g2_o21ai_1 _5792_ (.B1(_2188_),
    .Y(_2237_),
    .A1(_2184_),
    .A2(_2189_));
 sg13g2_nand2_1 _5793_ (.Y(_2238_),
    .A(net613),
    .B(_2071_));
 sg13g2_nand2_1 _5794_ (.Y(_2239_),
    .A(net619),
    .B(_2135_));
 sg13g2_nand2_1 _5795_ (.Y(_2240_),
    .A(net619),
    .B(net588));
 sg13g2_nor2_1 _5796_ (.A(_2186_),
    .B(_2239_),
    .Y(_2241_));
 sg13g2_xnor2_1 _5797_ (.Y(_2242_),
    .A(_2185_),
    .B(_2240_));
 sg13g2_nor2_1 _5798_ (.A(_2238_),
    .B(_2242_),
    .Y(_2243_));
 sg13g2_xor2_1 _5799_ (.B(_2242_),
    .A(_2238_),
    .X(_2244_));
 sg13g2_nand2_1 _5800_ (.Y(_2245_),
    .A(_2237_),
    .B(_2244_));
 sg13g2_xnor2_1 _5801_ (.Y(_2246_),
    .A(_2237_),
    .B(_2244_));
 sg13g2_nand2_1 _5802_ (.Y(_2247_),
    .A(net593),
    .B(_2015_));
 sg13g2_nand2_1 _5803_ (.Y(_2248_),
    .A(_2177_),
    .B(_2179_));
 sg13g2_nand3_1 _5804_ (.B(net590),
    .C(net595),
    .A(net611),
    .Y(_2249_));
 sg13g2_nand2_2 _5805_ (.Y(_2250_),
    .A(_2248_),
    .B(_2249_));
 sg13g2_xnor2_1 _5806_ (.Y(_2251_),
    .A(_2247_),
    .B(_2250_));
 sg13g2_xor2_1 _5807_ (.B(_2251_),
    .A(_2246_),
    .X(_2252_));
 sg13g2_xnor2_1 _5808_ (.Y(_2253_),
    .A(_2236_),
    .B(_2252_));
 sg13g2_o21ai_1 _5809_ (.B1(_1998_),
    .Y(_2254_),
    .A1(_1979_),
    .A2(_1996_));
 sg13g2_inv_1 _5810_ (.Y(_2255_),
    .A(_2254_));
 sg13g2_nor2_2 _5811_ (.A(_2006_),
    .B(_2254_),
    .Y(_2256_));
 sg13g2_nand2_1 _5812_ (.Y(_2257_),
    .A(net624),
    .B(net587));
 sg13g2_nand3_1 _5813_ (.B(_2198_),
    .C(_2256_),
    .A(net682),
    .Y(_2258_));
 sg13g2_o21ai_1 _5814_ (.B1(_2257_),
    .Y(_2259_),
    .A1(_2661_),
    .A2(_2254_));
 sg13g2_nand2_2 _5815_ (.Y(_2260_),
    .A(_2258_),
    .B(_2259_));
 sg13g2_nor2_1 _5816_ (.A(_2253_),
    .B(_2260_),
    .Y(_2261_));
 sg13g2_xor2_1 _5817_ (.B(_2260_),
    .A(_2253_),
    .X(_2262_));
 sg13g2_nor2b_1 _5818_ (.A(_2200_),
    .B_N(_2262_),
    .Y(_2263_));
 sg13g2_xnor2_1 _5819_ (.Y(_2264_),
    .A(_2200_),
    .B(_2262_));
 sg13g2_xnor2_1 _5820_ (.Y(_2265_),
    .A(_2234_),
    .B(_2264_));
 sg13g2_nand2_1 _5821_ (.Y(_2266_),
    .A(_2208_),
    .B(_2265_));
 sg13g2_xnor2_1 _5822_ (.Y(_2267_),
    .A(_2208_),
    .B(_2265_));
 sg13g2_xor2_1 _5823_ (.B(_2267_),
    .A(_2228_),
    .X(_2268_));
 sg13g2_and2_1 _5824_ (.A(_2227_),
    .B(_2268_),
    .X(_2269_));
 sg13g2_or2_1 _5825_ (.X(_2270_),
    .B(_2268_),
    .A(_2227_));
 sg13g2_xor2_1 _5826_ (.B(_2268_),
    .A(_2227_),
    .X(_2271_));
 sg13g2_xnor2_1 _5827_ (.Y(_2272_),
    .A(_2226_),
    .B(_2271_));
 sg13g2_nor2_1 _5828_ (.A(_2163_),
    .B(_2272_),
    .Y(_2273_));
 sg13g2_xor2_1 _5829_ (.B(_2272_),
    .A(_2163_),
    .X(_2274_));
 sg13g2_nor2b_1 _5830_ (.A(_2217_),
    .B_N(_2274_),
    .Y(_2275_));
 sg13g2_xnor2_1 _5831_ (.Y(_2276_),
    .A(_2217_),
    .B(_2274_));
 sg13g2_a21oi_1 _5832_ (.A1(_2225_),
    .A2(_2276_),
    .Y(_2277_),
    .B1(net596));
 sg13g2_o21ai_1 _5833_ (.B1(_2277_),
    .Y(_2278_),
    .A1(_2225_),
    .A2(_2276_));
 sg13g2_a21oi_1 _5834_ (.A1(_2224_),
    .A2(_2278_),
    .Y(_0328_),
    .B1(net719));
 sg13g2_a21o_1 _5835_ (.A2(_2276_),
    .A1(_2225_),
    .B1(_2275_),
    .X(_2279_));
 sg13g2_a21oi_1 _5836_ (.A1(_2226_),
    .A2(_2270_),
    .Y(_2280_),
    .B1(_2269_));
 sg13g2_o21ai_1 _5837_ (.B1(_2266_),
    .Y(_2281_),
    .A1(_2228_),
    .A2(_2267_));
 sg13g2_nor2_1 _5838_ (.A(_2231_),
    .B(_2233_),
    .Y(_2282_));
 sg13g2_a21oi_1 _5839_ (.A1(_2235_),
    .A2(_2264_),
    .Y(_2283_),
    .B1(_2263_));
 sg13g2_o21ai_1 _5840_ (.B1(_2249_),
    .Y(_2284_),
    .A1(_2247_),
    .A2(_2250_));
 sg13g2_a21o_1 _5841_ (.A2(_2252_),
    .A1(_2236_),
    .B1(_2284_),
    .X(_2285_));
 sg13g2_nand2_1 _5842_ (.Y(_2286_),
    .A(net593),
    .B(_2035_));
 sg13g2_nand2b_1 _5843_ (.Y(_2287_),
    .B(_2285_),
    .A_N(_2286_));
 sg13g2_xor2_1 _5844_ (.B(_2286_),
    .A(_2285_),
    .X(_2288_));
 sg13g2_nand2_1 _5845_ (.Y(_2289_),
    .A(net621),
    .B(_2198_));
 sg13g2_o21ai_1 _5846_ (.B1(_1975_),
    .Y(_2290_),
    .A1(_1967_),
    .A2(_1970_));
 sg13g2_nand2_1 _5847_ (.Y(_2291_),
    .A(_1980_),
    .B(_1987_));
 sg13g2_nand2_2 _5848_ (.Y(_2292_),
    .A(_2290_),
    .B(_2291_));
 sg13g2_and2_1 _5849_ (.A(_2290_),
    .B(_2291_),
    .X(_2293_));
 sg13g2_nor2_1 _5850_ (.A(_0012_),
    .B(_2292_),
    .Y(_2294_));
 sg13g2_nand2_1 _5851_ (.Y(_2295_),
    .A(_2256_),
    .B(_2294_));
 sg13g2_xor2_1 _5852_ (.B(_2294_),
    .A(_2256_),
    .X(_2296_));
 sg13g2_nand2b_1 _5853_ (.Y(_2297_),
    .B(_2296_),
    .A_N(_2289_));
 sg13g2_xor2_1 _5854_ (.B(_2296_),
    .A(_2289_),
    .X(_2298_));
 sg13g2_nor2_1 _5855_ (.A(_2258_),
    .B(_2298_),
    .Y(_2299_));
 sg13g2_xor2_1 _5856_ (.B(_2298_),
    .A(_2258_),
    .X(_2300_));
 sg13g2_o21ai_1 _5857_ (.B1(_2245_),
    .Y(_2301_),
    .A1(_2246_),
    .A2(_2251_));
 sg13g2_nand2_1 _5858_ (.Y(_2302_),
    .A(net600),
    .B(_2071_));
 sg13g2_and2_1 _5859_ (.A(net612),
    .B(_2135_),
    .X(_2303_));
 sg13g2_nand2_1 _5860_ (.Y(_2304_),
    .A(net613),
    .B(net589));
 sg13g2_nand3_1 _5861_ (.B(net589),
    .C(_2303_),
    .A(net619),
    .Y(_2305_));
 sg13g2_xnor2_1 _5862_ (.Y(_2306_),
    .A(_2239_),
    .B(_2304_));
 sg13g2_xor2_1 _5863_ (.B(_2306_),
    .A(_2302_),
    .X(_2307_));
 sg13g2_o21ai_1 _5864_ (.B1(_2307_),
    .Y(_2308_),
    .A1(_2241_),
    .A2(_2243_));
 sg13g2_or3_1 _5865_ (.A(_2241_),
    .B(_2243_),
    .C(_2307_),
    .X(_2309_));
 sg13g2_and2_1 _5866_ (.A(net611),
    .B(_2015_),
    .X(_2310_));
 sg13g2_nand2b_1 _5867_ (.Y(_2311_),
    .B(_2310_),
    .A_N(_2250_));
 sg13g2_xnor2_1 _5868_ (.Y(_2312_),
    .A(_2250_),
    .B(_2310_));
 sg13g2_xor2_1 _5869_ (.B(_2310_),
    .A(_2250_),
    .X(_2313_));
 sg13g2_a21o_1 _5870_ (.A2(_2309_),
    .A1(_2308_),
    .B1(_2312_),
    .X(_2314_));
 sg13g2_nand2_1 _5871_ (.Y(_2315_),
    .A(_2301_),
    .B(_2314_));
 sg13g2_xor2_1 _5872_ (.B(_2314_),
    .A(_2301_),
    .X(_2316_));
 sg13g2_nand2_1 _5873_ (.Y(_2317_),
    .A(_2300_),
    .B(_2316_));
 sg13g2_xnor2_1 _5874_ (.Y(_2318_),
    .A(_2300_),
    .B(_2316_));
 sg13g2_or3_1 _5875_ (.A(_2253_),
    .B(_2260_),
    .C(_2318_),
    .X(_2319_));
 sg13g2_xor2_1 _5876_ (.B(_2318_),
    .A(_2261_),
    .X(_2320_));
 sg13g2_xor2_1 _5877_ (.B(_2320_),
    .A(_2288_),
    .X(_2321_));
 sg13g2_nand2b_1 _5878_ (.Y(_2322_),
    .B(_2321_),
    .A_N(_2283_));
 sg13g2_xnor2_1 _5879_ (.Y(_2323_),
    .A(_2283_),
    .B(_2321_));
 sg13g2_nand2b_1 _5880_ (.Y(_2324_),
    .B(_2323_),
    .A_N(_2282_));
 sg13g2_xnor2_1 _5881_ (.Y(_2325_),
    .A(_2282_),
    .B(_2323_));
 sg13g2_nand2_1 _5882_ (.Y(_2326_),
    .A(_2281_),
    .B(_2325_));
 sg13g2_xnor2_1 _5883_ (.Y(_2327_),
    .A(_2281_),
    .B(_2325_));
 sg13g2_xor2_1 _5884_ (.B(_2327_),
    .A(_2280_),
    .X(_2328_));
 sg13g2_nand2_1 _5885_ (.Y(_2329_),
    .A(_2216_),
    .B(_2328_));
 sg13g2_xnor2_1 _5886_ (.Y(_2330_),
    .A(_2216_),
    .B(_2328_));
 sg13g2_nor3_1 _5887_ (.A(_2163_),
    .B(_2272_),
    .C(_2330_),
    .Y(_2331_));
 sg13g2_xnor2_1 _5888_ (.Y(_2332_),
    .A(_2273_),
    .B(_2330_));
 sg13g2_o21ai_1 _5889_ (.B1(_1993_),
    .Y(_2333_),
    .A1(_2279_),
    .A2(_2332_));
 sg13g2_a21oi_1 _5890_ (.A1(_2279_),
    .A2(_2332_),
    .Y(_2334_),
    .B1(_2333_));
 sg13g2_a21oi_1 _5891_ (.A1(net565),
    .A2(net599),
    .Y(_2335_),
    .B1(_2334_));
 sg13g2_nor2_1 _5892_ (.A(net719),
    .B(_2335_),
    .Y(_0329_));
 sg13g2_a21o_1 _5893_ (.A2(_2332_),
    .A1(_2279_),
    .B1(_2331_),
    .X(_2336_));
 sg13g2_o21ai_1 _5894_ (.B1(_2326_),
    .Y(_2337_),
    .A1(_2280_),
    .A2(_2327_));
 sg13g2_nand2_1 _5895_ (.Y(_2338_),
    .A(_2322_),
    .B(_2324_));
 sg13g2_o21ai_1 _5896_ (.B1(_2319_),
    .Y(_2339_),
    .A1(_2288_),
    .A2(_2320_));
 sg13g2_and2_2 _5897_ (.A(net611),
    .B(_2035_),
    .X(_2340_));
 sg13g2_and2_1 _5898_ (.A(_2249_),
    .B(_2311_),
    .X(_2341_));
 sg13g2_nand2_1 _5899_ (.Y(_2342_),
    .A(_2315_),
    .B(_2341_));
 sg13g2_nand2_2 _5900_ (.Y(_2343_),
    .A(_2340_),
    .B(_2342_));
 sg13g2_inv_1 _5901_ (.Y(_2344_),
    .A(_2343_));
 sg13g2_xor2_1 _5902_ (.B(_2342_),
    .A(_2340_),
    .X(_2345_));
 sg13g2_o21ai_1 _5903_ (.B1(_2305_),
    .Y(_2346_),
    .A1(_2302_),
    .A2(_2306_));
 sg13g2_nand2_1 _5904_ (.Y(_2347_),
    .A(net593),
    .B(_2071_));
 sg13g2_nand2_1 _5905_ (.Y(_2348_),
    .A(net601),
    .B(_2135_));
 sg13g2_nand3_1 _5906_ (.B(net589),
    .C(_2303_),
    .A(net600),
    .Y(_2349_));
 sg13g2_a21o_1 _5907_ (.A2(net589),
    .A1(net600),
    .B1(_2303_),
    .X(_2350_));
 sg13g2_nand2_1 _5908_ (.Y(_2351_),
    .A(_2349_),
    .B(_2350_));
 sg13g2_xor2_1 _5909_ (.B(_2351_),
    .A(_2347_),
    .X(_2352_));
 sg13g2_nand2_1 _5910_ (.Y(_2353_),
    .A(_2346_),
    .B(_2352_));
 sg13g2_xnor2_1 _5911_ (.Y(_2354_),
    .A(_2346_),
    .B(_2352_));
 sg13g2_xnor2_1 _5912_ (.Y(_2355_),
    .A(_2312_),
    .B(_2354_));
 sg13g2_xnor2_1 _5913_ (.Y(_2356_),
    .A(_2299_),
    .B(_2355_));
 sg13g2_xnor2_1 _5914_ (.Y(_2357_),
    .A(_2308_),
    .B(_2356_));
 sg13g2_nand2_1 _5915_ (.Y(_2358_),
    .A(_0576_),
    .B(net587));
 sg13g2_nor2_1 _5916_ (.A(_0580_),
    .B(_2292_),
    .Y(_2359_));
 sg13g2_nor2_1 _5917_ (.A(_0580_),
    .B(_2254_),
    .Y(_2360_));
 sg13g2_nand2_1 _5918_ (.Y(_2361_),
    .A(net624),
    .B(_2293_));
 sg13g2_nand2_1 _5919_ (.Y(_2362_),
    .A(_2256_),
    .B(_2359_));
 sg13g2_xnor2_1 _5920_ (.Y(_2363_),
    .A(_2360_),
    .B(_2361_));
 sg13g2_nand2b_1 _5921_ (.Y(_2364_),
    .B(_2363_),
    .A_N(_2358_));
 sg13g2_xor2_1 _5922_ (.B(_2363_),
    .A(_2358_),
    .X(_2365_));
 sg13g2_a21oi_2 _5923_ (.B1(_2365_),
    .Y(_2366_),
    .A2(_2297_),
    .A1(_2295_));
 sg13g2_nand3_1 _5924_ (.B(_2297_),
    .C(_2365_),
    .A(_2295_),
    .Y(_2367_));
 sg13g2_nor2b_1 _5925_ (.A(_2366_),
    .B_N(_2367_),
    .Y(_2368_));
 sg13g2_and2_2 _5926_ (.A(_2069_),
    .B(_2096_),
    .X(_2369_));
 sg13g2_nand3_1 _5927_ (.B(_2368_),
    .C(_2369_),
    .A(net682),
    .Y(_2370_));
 sg13g2_a21o_1 _5928_ (.A2(_2369_),
    .A1(net682),
    .B1(_2368_),
    .X(_2371_));
 sg13g2_nand2_1 _5929_ (.Y(_2372_),
    .A(_2370_),
    .B(_2371_));
 sg13g2_nor2_1 _5930_ (.A(_2357_),
    .B(_2372_),
    .Y(_2373_));
 sg13g2_xnor2_1 _5931_ (.Y(_2374_),
    .A(_2357_),
    .B(_2372_));
 sg13g2_xor2_1 _5932_ (.B(_2374_),
    .A(_2317_),
    .X(_2375_));
 sg13g2_nand2_1 _5933_ (.Y(_2376_),
    .A(_2345_),
    .B(_2375_));
 sg13g2_xor2_1 _5934_ (.B(_2375_),
    .A(_2345_),
    .X(_2377_));
 sg13g2_nand2_1 _5935_ (.Y(_2378_),
    .A(_2339_),
    .B(_2377_));
 sg13g2_xnor2_1 _5936_ (.Y(_2379_),
    .A(_2339_),
    .B(_2377_));
 sg13g2_xor2_1 _5937_ (.B(_2379_),
    .A(_2287_),
    .X(_2380_));
 sg13g2_and2_1 _5938_ (.A(_2338_),
    .B(_2380_),
    .X(_2381_));
 sg13g2_or2_1 _5939_ (.X(_2382_),
    .B(_2380_),
    .A(_2338_));
 sg13g2_xor2_1 _5940_ (.B(_2380_),
    .A(_2338_),
    .X(_2383_));
 sg13g2_xnor2_1 _5941_ (.Y(_2384_),
    .A(_2337_),
    .B(_2383_));
 sg13g2_nor2_1 _5942_ (.A(_2272_),
    .B(_2384_),
    .Y(_2385_));
 sg13g2_xor2_1 _5943_ (.B(_2384_),
    .A(_2272_),
    .X(_2386_));
 sg13g2_nor2b_1 _5944_ (.A(_2329_),
    .B_N(_2386_),
    .Y(_2387_));
 sg13g2_xnor2_1 _5945_ (.Y(_2388_),
    .A(_2329_),
    .B(_2386_));
 sg13g2_nand2_1 _5946_ (.Y(_2389_),
    .A(_2336_),
    .B(_2388_));
 sg13g2_nor2_1 _5947_ (.A(_2336_),
    .B(_2388_),
    .Y(_2390_));
 sg13g2_nor2_1 _5948_ (.A(net596),
    .B(_2390_),
    .Y(_2391_));
 sg13g2_a22oi_1 _5949_ (.Y(_2392_),
    .B1(_2389_),
    .B2(_2391_),
    .A2(net599),
    .A1(net568));
 sg13g2_nor2_1 _5950_ (.A(net719),
    .B(_2392_),
    .Y(_0330_));
 sg13g2_nand2_1 _5951_ (.Y(_2393_),
    .A(net504),
    .B(net599));
 sg13g2_a21o_1 _5952_ (.A2(_2388_),
    .A1(_2336_),
    .B1(_2387_),
    .X(_2394_));
 sg13g2_a21oi_1 _5953_ (.A1(_2337_),
    .A2(_2382_),
    .Y(_2395_),
    .B1(_2381_));
 sg13g2_o21ai_1 _5954_ (.B1(_2378_),
    .Y(_2396_),
    .A1(_2287_),
    .A2(_2379_));
 sg13g2_o21ai_1 _5955_ (.B1(_2376_),
    .Y(_2397_),
    .A1(_2317_),
    .A2(_2374_));
 sg13g2_nand2b_1 _5956_ (.Y(_2398_),
    .B(_2341_),
    .A_N(_2340_));
 sg13g2_a21oi_1 _5957_ (.A1(_2299_),
    .A2(_2355_),
    .Y(_2399_),
    .B1(_2398_));
 sg13g2_o21ai_1 _5958_ (.B1(_2399_),
    .Y(_2400_),
    .A1(_2308_),
    .A2(_2356_));
 sg13g2_and2_1 _5959_ (.A(_2343_),
    .B(_2400_),
    .X(_2401_));
 sg13g2_o21ai_1 _5960_ (.B1(_2353_),
    .Y(_2402_),
    .A1(_2313_),
    .A2(_2354_));
 sg13g2_o21ai_1 _5961_ (.B1(_2349_),
    .Y(_2403_),
    .A1(_2347_),
    .A2(_2351_));
 sg13g2_nand2_2 _5962_ (.Y(_2404_),
    .A(net609),
    .B(_2071_));
 sg13g2_nand2_1 _5963_ (.Y(_2405_),
    .A(net593),
    .B(_2135_));
 sg13g2_nand2_1 _5964_ (.Y(_2406_),
    .A(net594),
    .B(net589));
 sg13g2_xnor2_1 _5965_ (.Y(_2407_),
    .A(_2348_),
    .B(_2406_));
 sg13g2_or2_1 _5966_ (.X(_2408_),
    .B(_2407_),
    .A(_2404_));
 sg13g2_xor2_1 _5967_ (.B(_2407_),
    .A(_2404_),
    .X(_2409_));
 sg13g2_nand2_1 _5968_ (.Y(_2410_),
    .A(_2403_),
    .B(_2409_));
 sg13g2_xnor2_1 _5969_ (.Y(_2411_),
    .A(_2403_),
    .B(_2409_));
 sg13g2_xnor2_1 _5970_ (.Y(_2412_),
    .A(_2312_),
    .B(_2411_));
 sg13g2_xnor2_1 _5971_ (.Y(_2413_),
    .A(_2366_),
    .B(_2412_));
 sg13g2_nor2b_1 _5972_ (.A(_2413_),
    .B_N(_2402_),
    .Y(_2414_));
 sg13g2_xor2_1 _5973_ (.B(_2413_),
    .A(_2402_),
    .X(_2415_));
 sg13g2_inv_1 _5974_ (.Y(_2416_),
    .A(_2415_));
 sg13g2_nand2_1 _5975_ (.Y(_2417_),
    .A(net613),
    .B(net587));
 sg13g2_nor2_2 _5976_ (.A(_0575_),
    .B(_2292_),
    .Y(_2418_));
 sg13g2_nand2_1 _5977_ (.Y(_2419_),
    .A(net619),
    .B(_2255_));
 sg13g2_xor2_1 _5978_ (.B(_2419_),
    .A(_2359_),
    .X(_2420_));
 sg13g2_nor2_1 _5979_ (.A(_2417_),
    .B(_2420_),
    .Y(_2421_));
 sg13g2_xnor2_1 _5980_ (.Y(_2422_),
    .A(_2417_),
    .B(_2420_));
 sg13g2_a21oi_2 _5981_ (.B1(_2422_),
    .Y(_2423_),
    .A2(_2364_),
    .A1(_2362_));
 sg13g2_nand3_1 _5982_ (.B(_2364_),
    .C(_2422_),
    .A(_2362_),
    .Y(_2424_));
 sg13g2_nor2b_1 _5983_ (.A(_2423_),
    .B_N(_2424_),
    .Y(_2425_));
 sg13g2_a21oi_1 _5984_ (.A1(_1971_),
    .A2(_1973_),
    .Y(_2426_),
    .B1(net618));
 sg13g2_nand2_2 _5985_ (.Y(_2427_),
    .A(_2000_),
    .B(_2426_));
 sg13g2_nand2_1 _5986_ (.Y(_2428_),
    .A(net624),
    .B(_2033_));
 sg13g2_nor2_1 _5987_ (.A(_2006_),
    .B(_2427_),
    .Y(_2429_));
 sg13g2_nor2b_1 _5988_ (.A(_0012_),
    .B_N(_2033_),
    .Y(_2430_));
 sg13g2_nand2_2 _5989_ (.Y(_2431_),
    .A(_2429_),
    .B(_2430_));
 sg13g2_nand2_1 _5990_ (.Y(_2432_),
    .A(net624),
    .B(_2369_));
 sg13g2_o21ai_1 _5991_ (.B1(_2432_),
    .Y(_2433_),
    .A1(_0012_),
    .A2(_2427_));
 sg13g2_nand3_1 _5992_ (.B(_2431_),
    .C(_2433_),
    .A(_2425_),
    .Y(_2434_));
 sg13g2_a21o_1 _5993_ (.A2(_2433_),
    .A1(_2431_),
    .B1(_2425_),
    .X(_2435_));
 sg13g2_nand2_1 _5994_ (.Y(_2436_),
    .A(_2434_),
    .B(_2435_));
 sg13g2_nor2_1 _5995_ (.A(_2370_),
    .B(_2436_),
    .Y(_2437_));
 sg13g2_xor2_1 _5996_ (.B(_2436_),
    .A(_2370_),
    .X(_2438_));
 sg13g2_xnor2_1 _5997_ (.Y(_2439_),
    .A(_2415_),
    .B(_2438_));
 sg13g2_and2_1 _5998_ (.A(_2373_),
    .B(_2439_),
    .X(_2440_));
 sg13g2_xor2_1 _5999_ (.B(_2439_),
    .A(_2373_),
    .X(_2441_));
 sg13g2_xnor2_1 _6000_ (.Y(_2442_),
    .A(_2401_),
    .B(_2441_));
 sg13g2_nor2b_1 _6001_ (.A(_2442_),
    .B_N(_2397_),
    .Y(_2443_));
 sg13g2_xnor2_1 _6002_ (.Y(_2444_),
    .A(_2397_),
    .B(_2442_));
 sg13g2_xnor2_1 _6003_ (.Y(_2445_),
    .A(_2343_),
    .B(_2444_));
 sg13g2_nand2_1 _6004_ (.Y(_2446_),
    .A(_2396_),
    .B(_2445_));
 sg13g2_xnor2_1 _6005_ (.Y(_2447_),
    .A(_2396_),
    .B(_2445_));
 sg13g2_xnor2_1 _6006_ (.Y(_2448_),
    .A(_2395_),
    .B(_2447_));
 sg13g2_inv_1 _6007_ (.Y(_2449_),
    .A(_2448_));
 sg13g2_nand2_1 _6008_ (.Y(_2450_),
    .A(_2328_),
    .B(_2449_));
 sg13g2_xor2_1 _6009_ (.B(_2448_),
    .A(_2328_),
    .X(_2451_));
 sg13g2_nor3_1 _6010_ (.A(_2272_),
    .B(_2384_),
    .C(_2451_),
    .Y(_2452_));
 sg13g2_xnor2_1 _6011_ (.Y(_2453_),
    .A(_2385_),
    .B(_2451_));
 sg13g2_a21oi_1 _6012_ (.A1(_2394_),
    .A2(_2453_),
    .Y(_2454_),
    .B1(net597));
 sg13g2_o21ai_1 _6013_ (.B1(_2454_),
    .Y(_2455_),
    .A1(_2394_),
    .A2(_2453_));
 sg13g2_a21oi_1 _6014_ (.A1(_2393_),
    .A2(_2455_),
    .Y(_0331_),
    .B1(net720));
 sg13g2_nand2_1 _6015_ (.Y(_2456_),
    .A(net522),
    .B(net599));
 sg13g2_a21o_1 _6016_ (.A2(_2453_),
    .A1(_2394_),
    .B1(_2452_),
    .X(_2457_));
 sg13g2_o21ai_1 _6017_ (.B1(_2446_),
    .Y(_2458_),
    .A1(_2395_),
    .A2(_2447_));
 sg13g2_a21oi_1 _6018_ (.A1(_2344_),
    .A2(_2444_),
    .Y(_2459_),
    .B1(_2443_));
 sg13g2_a21oi_1 _6019_ (.A1(_2401_),
    .A2(_2441_),
    .Y(_2460_),
    .B1(_2440_));
 sg13g2_a21oi_1 _6020_ (.A1(_2416_),
    .A2(_2438_),
    .Y(_2461_),
    .B1(_2437_));
 sg13g2_o21ai_1 _6021_ (.B1(_2410_),
    .Y(_2462_),
    .A1(_2313_),
    .A2(_2411_));
 sg13g2_inv_1 _6022_ (.Y(_2463_),
    .A(_2462_));
 sg13g2_o21ai_1 _6023_ (.B1(_2408_),
    .Y(_2464_),
    .A1(_2348_),
    .A2(_2406_));
 sg13g2_nand2_1 _6024_ (.Y(_2465_),
    .A(net609),
    .B(net588));
 sg13g2_nor2_1 _6025_ (.A(_2405_),
    .B(_2465_),
    .Y(_2466_));
 sg13g2_nor2_1 _6026_ (.A(_2136_),
    .B(_2465_),
    .Y(_2467_));
 sg13g2_xnor2_1 _6027_ (.Y(_2468_),
    .A(_2405_),
    .B(_2465_));
 sg13g2_nor2_1 _6028_ (.A(_2404_),
    .B(_2468_),
    .Y(_2469_));
 sg13g2_xor2_1 _6029_ (.B(_2468_),
    .A(_2404_),
    .X(_2470_));
 sg13g2_nand2_1 _6030_ (.Y(_2471_),
    .A(_2464_),
    .B(_2470_));
 sg13g2_xnor2_1 _6031_ (.Y(_2472_),
    .A(_2464_),
    .B(_2470_));
 sg13g2_or2_1 _6032_ (.X(_2473_),
    .B(_2472_),
    .A(_2313_));
 sg13g2_xnor2_1 _6033_ (.Y(_2474_),
    .A(_2312_),
    .B(_2472_));
 sg13g2_nand2_1 _6034_ (.Y(_2475_),
    .A(_2423_),
    .B(_2474_));
 sg13g2_xnor2_1 _6035_ (.Y(_2476_),
    .A(_2423_),
    .B(_2474_));
 sg13g2_xnor2_1 _6036_ (.Y(_2477_),
    .A(_2462_),
    .B(_2476_));
 sg13g2_a21oi_1 _6037_ (.A1(_2360_),
    .A2(_2418_),
    .Y(_2478_),
    .B1(_2421_));
 sg13g2_nand2_1 _6038_ (.Y(_2479_),
    .A(net601),
    .B(net587));
 sg13g2_nand2_1 _6039_ (.Y(_2480_),
    .A(net612),
    .B(_2293_));
 sg13g2_nand2_1 _6040_ (.Y(_2481_),
    .A(net612),
    .B(_2255_));
 sg13g2_inv_1 _6041_ (.Y(_2482_),
    .A(_2481_));
 sg13g2_xor2_1 _6042_ (.B(_2481_),
    .A(_2418_),
    .X(_2483_));
 sg13g2_nor2_1 _6043_ (.A(_2479_),
    .B(_2483_),
    .Y(_2484_));
 sg13g2_xnor2_1 _6044_ (.Y(_2485_),
    .A(_2479_),
    .B(_2483_));
 sg13g2_nor2_1 _6045_ (.A(_2431_),
    .B(_2485_),
    .Y(_2486_));
 sg13g2_xnor2_1 _6046_ (.Y(_2487_),
    .A(_2431_),
    .B(_2485_));
 sg13g2_nor2_1 _6047_ (.A(_2478_),
    .B(_2487_),
    .Y(_2488_));
 sg13g2_xor2_1 _6048_ (.B(_2487_),
    .A(_2478_),
    .X(_2489_));
 sg13g2_nand2_1 _6049_ (.Y(_2490_),
    .A(net621),
    .B(_2369_));
 sg13g2_xnor2_1 _6050_ (.Y(_2491_),
    .A(_2429_),
    .B(_2430_));
 sg13g2_xor2_1 _6051_ (.B(_2491_),
    .A(_2490_),
    .X(_2492_));
 sg13g2_nand2_1 _6052_ (.Y(_2493_),
    .A(_2489_),
    .B(_2492_));
 sg13g2_xnor2_1 _6053_ (.Y(_2494_),
    .A(_2489_),
    .B(_2492_));
 sg13g2_nor2_1 _6054_ (.A(_2434_),
    .B(_2494_),
    .Y(_2495_));
 sg13g2_xor2_1 _6055_ (.B(_2494_),
    .A(_2434_),
    .X(_2496_));
 sg13g2_xor2_1 _6056_ (.B(_2496_),
    .A(_2477_),
    .X(_2497_));
 sg13g2_nand2b_1 _6057_ (.Y(_2498_),
    .B(_2497_),
    .A_N(_2461_));
 sg13g2_xnor2_1 _6058_ (.Y(_2499_),
    .A(_2461_),
    .B(_2497_));
 sg13g2_a21oi_1 _6059_ (.A1(_2366_),
    .A2(_2412_),
    .Y(_2500_),
    .B1(_2414_));
 sg13g2_and2_1 _6060_ (.A(_2343_),
    .B(_2398_),
    .X(_2501_));
 sg13g2_nand2b_1 _6061_ (.Y(_2502_),
    .B(_2500_),
    .A_N(_2501_));
 sg13g2_nand2_1 _6062_ (.Y(_2503_),
    .A(_2499_),
    .B(_2502_));
 sg13g2_xor2_1 _6063_ (.B(_2502_),
    .A(_2499_),
    .X(_2504_));
 sg13g2_nor2b_1 _6064_ (.A(_2460_),
    .B_N(_2504_),
    .Y(_2505_));
 sg13g2_xnor2_1 _6065_ (.Y(_2506_),
    .A(_2460_),
    .B(_2504_));
 sg13g2_xnor2_1 _6066_ (.Y(_2507_),
    .A(_2343_),
    .B(_2506_));
 sg13g2_nor2b_1 _6067_ (.A(_2459_),
    .B_N(_2507_),
    .Y(_2508_));
 sg13g2_xnor2_1 _6068_ (.Y(_2509_),
    .A(_2459_),
    .B(_2507_));
 sg13g2_xnor2_1 _6069_ (.Y(_2510_),
    .A(_2458_),
    .B(_2509_));
 sg13g2_nor2_1 _6070_ (.A(_2384_),
    .B(_2510_),
    .Y(_2511_));
 sg13g2_xor2_1 _6071_ (.B(_2510_),
    .A(_2384_),
    .X(_2512_));
 sg13g2_nor2b_1 _6072_ (.A(_2450_),
    .B_N(_2512_),
    .Y(_2513_));
 sg13g2_xnor2_1 _6073_ (.Y(_2514_),
    .A(_2450_),
    .B(_2512_));
 sg13g2_a21oi_1 _6074_ (.A1(_2457_),
    .A2(_2514_),
    .Y(_2515_),
    .B1(net597));
 sg13g2_o21ai_1 _6075_ (.B1(_2515_),
    .Y(_2516_),
    .A1(_2457_),
    .A2(_2514_));
 sg13g2_a21oi_1 _6076_ (.A1(_2456_),
    .A2(_2516_),
    .Y(_0332_),
    .B1(net720));
 sg13g2_a21oi_1 _6077_ (.A1(_2457_),
    .A2(_2514_),
    .Y(_2517_),
    .B1(_2513_));
 sg13g2_a21o_1 _6078_ (.A2(_2509_),
    .A1(_2458_),
    .B1(_2508_),
    .X(_2518_));
 sg13g2_a21o_1 _6079_ (.A2(_2506_),
    .A1(_2344_),
    .B1(_2505_),
    .X(_2519_));
 sg13g2_and2_1 _6080_ (.A(_2498_),
    .B(_2503_),
    .X(_2520_));
 sg13g2_o21ai_1 _6081_ (.B1(_2475_),
    .Y(_2521_),
    .A1(_2463_),
    .A2(_2476_));
 sg13g2_nor2b_1 _6082_ (.A(_2341_),
    .B_N(_2521_),
    .Y(_2522_));
 sg13g2_xnor2_1 _6083_ (.Y(_2523_),
    .A(_2341_),
    .B(_2521_));
 sg13g2_xnor2_1 _6084_ (.Y(_2524_),
    .A(_2340_),
    .B(_2523_));
 sg13g2_a21oi_2 _6085_ (.B1(_2495_),
    .Y(_2525_),
    .A2(_2496_),
    .A1(_2477_));
 sg13g2_nand2_1 _6086_ (.Y(_2526_),
    .A(_2471_),
    .B(_2473_));
 sg13g2_o21ai_1 _6087_ (.B1(net609),
    .Y(_2527_),
    .A1(net589),
    .A2(_2135_));
 sg13g2_nor2_1 _6088_ (.A(_2467_),
    .B(_2527_),
    .Y(_2528_));
 sg13g2_xnor2_1 _6089_ (.Y(_2529_),
    .A(_2404_),
    .B(_2528_));
 sg13g2_nor3_1 _6090_ (.A(_2466_),
    .B(_2469_),
    .C(_2529_),
    .Y(_2530_));
 sg13g2_o21ai_1 _6091_ (.B1(_2529_),
    .Y(_2531_),
    .A1(_2466_),
    .A2(_2469_));
 sg13g2_nor2b_2 _6092_ (.A(_2530_),
    .B_N(_2531_),
    .Y(_2532_));
 sg13g2_xnor2_1 _6093_ (.Y(_2533_),
    .A(_2313_),
    .B(_2532_));
 sg13g2_nor3_1 _6094_ (.A(_2486_),
    .B(_2488_),
    .C(_2533_),
    .Y(_2534_));
 sg13g2_a21o_1 _6095_ (.A2(_2473_),
    .A1(_2471_),
    .B1(_2534_),
    .X(_2535_));
 sg13g2_xnor2_1 _6096_ (.Y(_2536_),
    .A(_2526_),
    .B(_2534_));
 sg13g2_a21oi_2 _6097_ (.B1(_2484_),
    .Y(_2537_),
    .A2(_2482_),
    .A1(_2418_));
 sg13g2_o21ai_1 _6098_ (.B1(_2431_),
    .Y(_2538_),
    .A1(_2490_),
    .A2(_2491_));
 sg13g2_nand2_1 _6099_ (.Y(_2539_),
    .A(net593),
    .B(net587));
 sg13g2_and2_1 _6100_ (.A(net601),
    .B(_2293_),
    .X(_2540_));
 sg13g2_nand2_1 _6101_ (.Y(_2541_),
    .A(net600),
    .B(_2255_));
 sg13g2_xnor2_1 _6102_ (.Y(_2542_),
    .A(_2480_),
    .B(_2541_));
 sg13g2_or2_1 _6103_ (.X(_2543_),
    .B(_2542_),
    .A(_2539_));
 sg13g2_xnor2_1 _6104_ (.Y(_2544_),
    .A(_2539_),
    .B(_2542_));
 sg13g2_nand2b_1 _6105_ (.Y(_2545_),
    .B(_2538_),
    .A_N(_2544_));
 sg13g2_xor2_1 _6106_ (.B(_2544_),
    .A(_2538_),
    .X(_2546_));
 sg13g2_xor2_1 _6107_ (.B(_2546_),
    .A(_2537_),
    .X(_2547_));
 sg13g2_nand2_1 _6108_ (.Y(_2548_),
    .A(_0576_),
    .B(_2369_));
 sg13g2_nand2_1 _6109_ (.Y(_2549_),
    .A(net621),
    .B(_2033_));
 sg13g2_nor2_1 _6110_ (.A(_0580_),
    .B(_2427_),
    .Y(_2550_));
 sg13g2_inv_1 _6111_ (.Y(_2551_),
    .A(_2550_));
 sg13g2_xnor2_1 _6112_ (.Y(_2552_),
    .A(_2428_),
    .B(_2550_));
 sg13g2_nand2b_1 _6113_ (.Y(_2553_),
    .B(_2552_),
    .A_N(_2548_));
 sg13g2_xor2_1 _6114_ (.B(_2552_),
    .A(_2548_),
    .X(_2554_));
 sg13g2_nand3_1 _6115_ (.B(_1979_),
    .C(_2290_),
    .A(net682),
    .Y(_2555_));
 sg13g2_xor2_1 _6116_ (.B(_2555_),
    .A(_2554_),
    .X(_2556_));
 sg13g2_xnor2_1 _6117_ (.Y(_2557_),
    .A(_2547_),
    .B(_2556_));
 sg13g2_nor2_1 _6118_ (.A(_2493_),
    .B(_2557_),
    .Y(_2558_));
 sg13g2_xor2_1 _6119_ (.B(_2557_),
    .A(_2493_),
    .X(_2559_));
 sg13g2_xnor2_1 _6120_ (.Y(_2560_),
    .A(_2536_),
    .B(_2559_));
 sg13g2_xor2_1 _6121_ (.B(_2560_),
    .A(_2525_),
    .X(_2561_));
 sg13g2_nand2b_1 _6122_ (.Y(_2562_),
    .B(_2561_),
    .A_N(_2524_));
 sg13g2_xnor2_1 _6123_ (.Y(_2563_),
    .A(_2524_),
    .B(_2561_));
 sg13g2_nand2b_1 _6124_ (.Y(_2564_),
    .B(_2563_),
    .A_N(_2520_));
 sg13g2_xnor2_1 _6125_ (.Y(_2565_),
    .A(_2520_),
    .B(_2563_));
 sg13g2_nand2_1 _6126_ (.Y(_2566_),
    .A(_2344_),
    .B(_2565_));
 sg13g2_xnor2_1 _6127_ (.Y(_2567_),
    .A(_2343_),
    .B(_2565_));
 sg13g2_and2_1 _6128_ (.A(_2519_),
    .B(_2567_),
    .X(_2568_));
 sg13g2_xnor2_1 _6129_ (.Y(_2569_),
    .A(_2519_),
    .B(_2567_));
 sg13g2_inv_1 _6130_ (.Y(_2570_),
    .A(_2569_));
 sg13g2_xnor2_1 _6131_ (.Y(_2571_),
    .A(_2518_),
    .B(_2570_));
 sg13g2_nor2_1 _6132_ (.A(_2448_),
    .B(_2571_),
    .Y(_2572_));
 sg13g2_xnor2_1 _6133_ (.Y(_2573_),
    .A(_2449_),
    .B(_2571_));
 sg13g2_nand2_1 _6134_ (.Y(_2574_),
    .A(_2511_),
    .B(_2573_));
 sg13g2_xnor2_1 _6135_ (.Y(_2575_),
    .A(_2511_),
    .B(_2573_));
 sg13g2_nor2_1 _6136_ (.A(_2517_),
    .B(_2575_),
    .Y(_2576_));
 sg13g2_nand2_1 _6137_ (.Y(_2577_),
    .A(_2517_),
    .B(_2575_));
 sg13g2_nor2_1 _6138_ (.A(net597),
    .B(_2576_),
    .Y(_2578_));
 sg13g2_a22oi_1 _6139_ (.Y(_2579_),
    .B1(_2577_),
    .B2(_2578_),
    .A2(net599),
    .A1(net548));
 sg13g2_nor2_1 _6140_ (.A(net720),
    .B(_2579_),
    .Y(_0333_));
 sg13g2_nand2_1 _6141_ (.Y(_2580_),
    .A(net456),
    .B(net599));
 sg13g2_o21ai_1 _6142_ (.B1(_2574_),
    .Y(_2581_),
    .A1(_2517_),
    .A2(_2575_));
 sg13g2_a21oi_1 _6143_ (.A1(_2518_),
    .A2(_2570_),
    .Y(_2582_),
    .B1(_2568_));
 sg13g2_and2_1 _6144_ (.A(_2564_),
    .B(_2566_),
    .X(_2583_));
 sg13g2_o21ai_1 _6145_ (.B1(_2562_),
    .Y(_2584_),
    .A1(_2525_),
    .A2(_2560_));
 sg13g2_a21oi_1 _6146_ (.A1(_2340_),
    .A2(_2523_),
    .Y(_2585_),
    .B1(_2522_));
 sg13g2_a21oi_1 _6147_ (.A1(_2536_),
    .A2(_2559_),
    .Y(_2586_),
    .B1(_2558_));
 sg13g2_a22oi_1 _6148_ (.Y(_2587_),
    .B1(_2547_),
    .B2(_2556_),
    .A2(_2532_),
    .A1(_2312_));
 sg13g2_nand2_1 _6149_ (.Y(_2588_),
    .A(_2531_),
    .B(_2587_));
 sg13g2_o21ai_1 _6150_ (.B1(_2313_),
    .Y(_2589_),
    .A1(_2554_),
    .A2(_2555_));
 sg13g2_o21ai_1 _6151_ (.B1(_2545_),
    .Y(_2590_),
    .A1(_2537_),
    .A2(_2546_));
 sg13g2_nand2_1 _6152_ (.Y(_2591_),
    .A(net612),
    .B(_2369_));
 sg13g2_nand3_1 _6153_ (.B(net623),
    .C(_2290_),
    .A(_1979_),
    .Y(_2592_));
 sg13g2_nand3_1 _6154_ (.B(_1968_),
    .C(_1974_),
    .A(net682),
    .Y(_2593_));
 sg13g2_xor2_1 _6155_ (.B(_2593_),
    .A(_2592_),
    .X(_2594_));
 sg13g2_nor2_1 _6156_ (.A(_0575_),
    .B(_2427_),
    .Y(_2595_));
 sg13g2_xnor2_1 _6157_ (.Y(_2596_),
    .A(_2549_),
    .B(_2595_));
 sg13g2_xnor2_1 _6158_ (.Y(_2597_),
    .A(_2594_),
    .B(_2596_));
 sg13g2_xnor2_1 _6159_ (.Y(_2598_),
    .A(_2591_),
    .B(_2597_));
 sg13g2_o21ai_1 _6160_ (.B1(_2553_),
    .Y(_2599_),
    .A1(_2428_),
    .A2(_2551_));
 sg13g2_nand2_1 _6161_ (.Y(_2600_),
    .A(net610),
    .B(net587));
 sg13g2_and2_1 _6162_ (.A(net593),
    .B(_2255_),
    .X(_2601_));
 sg13g2_xnor2_1 _6163_ (.Y(_2602_),
    .A(_2600_),
    .B(_2601_));
 sg13g2_xnor2_1 _6164_ (.Y(_2603_),
    .A(_2540_),
    .B(_2602_));
 sg13g2_xnor2_1 _6165_ (.Y(_2604_),
    .A(_2599_),
    .B(_2603_));
 sg13g2_xnor2_1 _6166_ (.Y(_2605_),
    .A(_2598_),
    .B(_2604_));
 sg13g2_xnor2_1 _6167_ (.Y(_2606_),
    .A(_2590_),
    .B(_2605_));
 sg13g2_xnor2_1 _6168_ (.Y(_2607_),
    .A(_2589_),
    .B(_2606_));
 sg13g2_xnor2_1 _6169_ (.Y(_2608_),
    .A(_2588_),
    .B(_2607_));
 sg13g2_a22oi_1 _6170_ (.Y(_2609_),
    .B1(_2540_),
    .B2(_2482_),
    .A2(_2531_),
    .A1(net610));
 sg13g2_a21oi_1 _6171_ (.A1(_2543_),
    .A2(_2609_),
    .Y(_2610_),
    .B1(_2501_));
 sg13g2_xnor2_1 _6172_ (.Y(_2611_),
    .A(_2535_),
    .B(_2610_));
 sg13g2_xnor2_1 _6173_ (.Y(_2612_),
    .A(_2608_),
    .B(_2611_));
 sg13g2_xnor2_1 _6174_ (.Y(_2613_),
    .A(_2586_),
    .B(_2612_));
 sg13g2_xnor2_1 _6175_ (.Y(_2614_),
    .A(_2585_),
    .B(_2613_));
 sg13g2_xnor2_1 _6176_ (.Y(_2615_),
    .A(_2584_),
    .B(_2614_));
 sg13g2_xnor2_1 _6177_ (.Y(_2616_),
    .A(_2583_),
    .B(_2615_));
 sg13g2_xnor2_1 _6178_ (.Y(_2617_),
    .A(_2510_),
    .B(_2616_));
 sg13g2_xnor2_1 _6179_ (.Y(_2618_),
    .A(_2582_),
    .B(_2617_));
 sg13g2_xnor2_1 _6180_ (.Y(_2619_),
    .A(_2572_),
    .B(_2618_));
 sg13g2_a21oi_1 _6181_ (.A1(_2581_),
    .A2(_2619_),
    .Y(_2620_),
    .B1(net597));
 sg13g2_o21ai_1 _6182_ (.B1(_2620_),
    .Y(_2621_),
    .A1(_2581_),
    .A2(_2619_));
 sg13g2_a21oi_1 _6183_ (.A1(_2580_),
    .A2(_2621_),
    .Y(_0334_),
    .B1(net723));
 sg13g2_dfrbp_1 _6184_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net73),
    .D(net856),
    .Q_N(_0054_),
    .Q(\core.lstate[2] ));
 sg13g2_dfrbp_1 _6185_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net45),
    .D(net768),
    .Q_N(_0057_),
    .Q(\core.lstate[1] ));
 sg13g2_dfrbp_1 _6186_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net44),
    .D(net786),
    .Q_N(_0056_),
    .Q(\core.lstate[0] ));
 sg13g2_dfrbp_1 _6187_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net43),
    .D(_0061_),
    .Q_N(_3081_),
    .Q(\core.byte_acc[4] ));
 sg13g2_dfrbp_1 _6188_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net41),
    .D(_0062_),
    .Q_N(_3080_),
    .Q(\core.byte_acc[5] ));
 sg13g2_dfrbp_1 _6189_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net39),
    .D(_0063_),
    .Q_N(_3079_),
    .Q(\core.byte_acc[6] ));
 sg13g2_dfrbp_1 _6190_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net37),
    .D(_0064_),
    .Q_N(_3078_),
    .Q(\core.byte_acc[7] ));
 sg13g2_dfrbp_1 _6191_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net35),
    .D(_0065_),
    .Q_N(_3077_),
    .Q(\core.load_prev ));
 sg13g2_dfrbp_1 _6192_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net34),
    .D(_0066_),
    .Q_N(_3076_),
    .Q(\core.params[0][0] ));
 sg13g2_dfrbp_1 _6193_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net32),
    .D(net448),
    .Q_N(_3075_),
    .Q(\core.params[0][1] ));
 sg13g2_dfrbp_1 _6194_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net30),
    .D(_0068_),
    .Q_N(_3074_),
    .Q(\core.params[0][2] ));
 sg13g2_dfrbp_1 _6195_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net28),
    .D(_0069_),
    .Q_N(_3073_),
    .Q(\core.params[0][3] ));
 sg13g2_dfrbp_1 _6196_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net26),
    .D(_0070_),
    .Q_N(_3072_),
    .Q(\core.params[0][4] ));
 sg13g2_dfrbp_1 _6197_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net308),
    .D(_0071_),
    .Q_N(_3071_),
    .Q(\core.params[0][5] ));
 sg13g2_dfrbp_1 _6198_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net306),
    .D(_0072_),
    .Q_N(_3070_),
    .Q(\core.params[0][6] ));
 sg13g2_dfrbp_1 _6199_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net304),
    .D(net431),
    .Q_N(_2857_),
    .Q(\core.params[0][7] ));
 sg13g2_dfrbp_1 _6200_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net302),
    .D(_0074_),
    .Q_N(_3069_),
    .Q(\core.tau_w[8] ));
 sg13g2_dfrbp_1 _6201_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net300),
    .D(_0075_),
    .Q_N(_3068_),
    .Q(\core.tau_w[9] ));
 sg13g2_dfrbp_1 _6202_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net298),
    .D(net391),
    .Q_N(_0022_),
    .Q(\core.tau_w[10] ));
 sg13g2_dfrbp_1 _6203_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net296),
    .D(_0077_),
    .Q_N(_3067_),
    .Q(\core.tau_w[11] ));
 sg13g2_dfrbp_1 _6204_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net294),
    .D(_0078_),
    .Q_N(_0016_),
    .Q(\core.tau_w[12] ));
 sg13g2_dfrbp_1 _6205_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net292),
    .D(net810),
    .Q_N(_3066_),
    .Q(\core.tau_w[13] ));
 sg13g2_dfrbp_1 _6206_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net290),
    .D(_0080_),
    .Q_N(_0017_),
    .Q(\core.tau_w[14] ));
 sg13g2_dfrbp_1 _6207_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net288),
    .D(_0081_),
    .Q_N(_3065_),
    .Q(\core.tau_w[15] ));
 sg13g2_dfrbp_1 _6208_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net286),
    .D(_0082_),
    .Q_N(_3064_),
    .Q(\core.param_b[8] ));
 sg13g2_dfrbp_1 _6209_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net284),
    .D(_0083_),
    .Q_N(_3063_),
    .Q(\core.param_b[9] ));
 sg13g2_dfrbp_1 _6210_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net282),
    .D(_0084_),
    .Q_N(_3062_),
    .Q(\core.param_b[10] ));
 sg13g2_dfrbp_1 _6211_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net280),
    .D(_0085_),
    .Q_N(_3061_),
    .Q(\core.param_b[11] ));
 sg13g2_dfrbp_1 _6212_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net278),
    .D(_0086_),
    .Q_N(_3060_),
    .Q(\core.param_b[12] ));
 sg13g2_dfrbp_1 _6213_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net276),
    .D(_0087_),
    .Q_N(_3059_),
    .Q(\core.param_b[13] ));
 sg13g2_dfrbp_1 _6214_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net274),
    .D(_0088_),
    .Q_N(_3058_),
    .Q(\core.param_b[14] ));
 sg13g2_dfrbp_1 _6215_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net272),
    .D(_0089_),
    .Q_N(_3057_),
    .Q(\core.param_b[15] ));
 sg13g2_dfrbp_1 _6216_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net270),
    .D(_0090_),
    .Q_N(_3056_),
    .Q(\core.capacitance[8] ));
 sg13g2_dfrbp_1 _6217_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net268),
    .D(_0091_),
    .Q_N(_3055_),
    .Q(\core.capacitance[9] ));
 sg13g2_dfrbp_1 _6218_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net266),
    .D(_0092_),
    .Q_N(_0045_),
    .Q(\core.capacitance[10] ));
 sg13g2_dfrbp_1 _6219_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net264),
    .D(_0093_),
    .Q_N(_3054_),
    .Q(\core.capacitance[11] ));
 sg13g2_dfrbp_1 _6220_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net262),
    .D(_0094_),
    .Q_N(_0030_),
    .Q(\core.capacitance[12] ));
 sg13g2_dfrbp_1 _6221_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net260),
    .D(_0095_),
    .Q_N(_3053_),
    .Q(\core.capacitance[13] ));
 sg13g2_dfrbp_1 _6222_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net258),
    .D(_0096_),
    .Q_N(_0031_),
    .Q(\core.capacitance[14] ));
 sg13g2_dfrbp_1 _6223_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net256),
    .D(_0097_),
    .Q_N(_3052_),
    .Q(\core.capacitance[15] ));
 sg13g2_dfrbp_1 _6224_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net254),
    .D(net501),
    .Q_N(_3051_),
    .Q(\core.param_a[8] ));
 sg13g2_dfrbp_1 _6225_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net252),
    .D(net779),
    .Q_N(_3050_),
    .Q(\core.param_a[9] ));
 sg13g2_dfrbp_1 _6226_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net250),
    .D(net471),
    .Q_N(_3049_),
    .Q(\core.param_a[10] ));
 sg13g2_dfrbp_1 _6227_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net248),
    .D(net360),
    .Q_N(_3048_),
    .Q(\core.param_a[11] ));
 sg13g2_dfrbp_1 _6228_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net246),
    .D(_0102_),
    .Q_N(_3047_),
    .Q(\core.param_a[12] ));
 sg13g2_dfrbp_1 _6229_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net244),
    .D(_0103_),
    .Q_N(_3046_),
    .Q(\core.param_a[13] ));
 sg13g2_dfrbp_1 _6230_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net242),
    .D(_0104_),
    .Q_N(_3045_),
    .Q(\core.param_a[14] ));
 sg13g2_dfrbp_1 _6231_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net74),
    .D(_0105_),
    .Q_N(_3082_),
    .Q(\core.param_a[15] ));
 sg13g2_dfrbp_1 _6232_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net75),
    .D(_0005_),
    .Q_N(_3083_),
    .Q(\core.compute_state[0] ));
 sg13g2_dfrbp_1 _6233_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net76),
    .D(_0000_),
    .Q_N(_3084_),
    .Q(\core.compute_state[1] ));
 sg13g2_dfrbp_1 _6234_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net77),
    .D(_0001_),
    .Q_N(_3085_),
    .Q(\core.compute_state[2] ));
 sg13g2_dfrbp_1 _6235_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net78),
    .D(_0002_),
    .Q_N(_3086_),
    .Q(\core.compute_state[3] ));
 sg13g2_dfrbp_1 _6236_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net79),
    .D(_0003_),
    .Q_N(_3087_),
    .Q(\core.compute_state[4] ));
 sg13g2_dfrbp_1 _6237_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net285),
    .D(_0004_),
    .Q_N(_3088_),
    .Q(\core.compute_state[5] ));
 sg13g2_dfrbp_1 _6238_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net240),
    .D(_0006_),
    .Q_N(_3044_),
    .Q(\core.compute_state[6] ));
 sg13g2_dfrbp_1 _6239_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net238),
    .D(_0106_),
    .Q_N(_3043_),
    .Q(\core.params[7][0] ));
 sg13g2_dfrbp_1 _6240_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net236),
    .D(_0107_),
    .Q_N(_3042_),
    .Q(\core.params[7][1] ));
 sg13g2_dfrbp_1 _6241_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net234),
    .D(_0108_),
    .Q_N(_3041_),
    .Q(\core.params[7][2] ));
 sg13g2_dfrbp_1 _6242_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net232),
    .D(net367),
    .Q_N(_3040_),
    .Q(\core.params[7][3] ));
 sg13g2_dfrbp_1 _6243_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net230),
    .D(_0110_),
    .Q_N(_3039_),
    .Q(\core.params[7][4] ));
 sg13g2_dfrbp_1 _6244_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net228),
    .D(_0111_),
    .Q_N(_3038_),
    .Q(\core.params[7][5] ));
 sg13g2_dfrbp_1 _6245_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net226),
    .D(net444),
    .Q_N(_3037_),
    .Q(\core.params[7][6] ));
 sg13g2_dfrbp_1 _6246_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net224),
    .D(net411),
    .Q_N(_3036_),
    .Q(\core.params[7][7] ));
 sg13g2_dfrbp_1 _6247_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net223),
    .D(net423),
    .Q_N(_3035_),
    .Q(\core.params[6][0] ));
 sg13g2_dfrbp_1 _6248_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net221),
    .D(net506),
    .Q_N(_3034_),
    .Q(\core.params[6][1] ));
 sg13g2_dfrbp_1 _6249_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net220),
    .D(net508),
    .Q_N(_3033_),
    .Q(\core.params[6][2] ));
 sg13g2_dfrbp_1 _6250_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net218),
    .D(_0117_),
    .Q_N(_3032_),
    .Q(\core.params[6][3] ));
 sg13g2_dfrbp_1 _6251_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net217),
    .D(_0118_),
    .Q_N(_3031_),
    .Q(\core.params[6][4] ));
 sg13g2_dfrbp_1 _6252_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net215),
    .D(_0119_),
    .Q_N(_3030_),
    .Q(\core.params[6][5] ));
 sg13g2_dfrbp_1 _6253_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net213),
    .D(_0120_),
    .Q_N(_3029_),
    .Q(\core.params[6][6] ));
 sg13g2_dfrbp_1 _6254_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net211),
    .D(net325),
    .Q_N(_2858_),
    .Q(\core.params[6][7] ));
 sg13g2_dfrbp_1 _6255_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net209),
    .D(_0122_),
    .Q_N(_3028_),
    .Q(\core.r_ready ));
 sg13g2_dfrbp_1 _6256_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net207),
    .D(_0123_),
    .Q_N(_3027_),
    .Q(\core.watchdog_cnt[0] ));
 sg13g2_dfrbp_1 _6257_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net206),
    .D(net814),
    .Q_N(_3026_),
    .Q(\core.watchdog_cnt[1] ));
 sg13g2_dfrbp_1 _6258_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net205),
    .D(_0125_),
    .Q_N(_0046_),
    .Q(\core.watchdog_cnt[2] ));
 sg13g2_dfrbp_1 _6259_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net204),
    .D(_0126_),
    .Q_N(_3025_),
    .Q(\core.watchdog_cnt[3] ));
 sg13g2_dfrbp_1 _6260_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net203),
    .D(_0127_),
    .Q_N(_0047_),
    .Q(\core.watchdog_cnt[4] ));
 sg13g2_dfrbp_1 _6261_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net202),
    .D(_0128_),
    .Q_N(_3024_),
    .Q(\core.watchdog_cnt[5] ));
 sg13g2_dfrbp_1 _6262_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net201),
    .D(_0129_),
    .Q_N(_0048_),
    .Q(\core.watchdog_cnt[6] ));
 sg13g2_dfrbp_1 _6263_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net200),
    .D(_0130_),
    .Q_N(_3023_),
    .Q(\core.watchdog_cnt[7] ));
 sg13g2_dfrbp_1 _6264_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net199),
    .D(_0131_),
    .Q_N(_0049_),
    .Q(\core.watchdog_cnt[8] ));
 sg13g2_dfrbp_1 _6265_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net198),
    .D(_0132_),
    .Q_N(_3022_),
    .Q(\core.watchdog_cnt[9] ));
 sg13g2_dfrbp_1 _6266_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net197),
    .D(_0133_),
    .Q_N(_0050_),
    .Q(\core.watchdog_cnt[10] ));
 sg13g2_dfrbp_1 _6267_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net196),
    .D(net393),
    .Q_N(_3021_),
    .Q(\core.watchdog_cnt[11] ));
 sg13g2_dfrbp_1 _6268_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net195),
    .D(_0135_),
    .Q_N(_0055_),
    .Q(\core.param_idx[0] ));
 sg13g2_dfrbp_1 _6269_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net194),
    .D(net848),
    .Q_N(_3020_),
    .Q(\core.param_idx[1] ));
 sg13g2_dfrbp_1 _6270_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net193),
    .D(_0137_),
    .Q_N(_3019_),
    .Q(\core.param_idx[2] ));
 sg13g2_dfrbp_1 _6271_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net192),
    .D(net319),
    .Q_N(_0051_),
    .Q(\core.nibble_cnt ));
 sg13g2_dfrbp_1 _6272_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net191),
    .D(_0139_),
    .Q_N(_3018_),
    .Q(\core.byte_acc[0] ));
 sg13g2_dfrbp_1 _6273_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net189),
    .D(_0140_),
    .Q_N(_3017_),
    .Q(\core.byte_acc[1] ));
 sg13g2_dfrbp_1 _6274_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net187),
    .D(_0141_),
    .Q_N(_3016_),
    .Q(\core.byte_acc[2] ));
 sg13g2_dfrbp_1 _6275_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net185),
    .D(_0142_),
    .Q_N(_3015_),
    .Q(\core.byte_acc[3] ));
 sg13g2_dfrbp_1 _6276_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net183),
    .D(_0143_),
    .Q_N(_3014_),
    .Q(\core.leak_current[1] ));
 sg13g2_dfrbp_1 _6277_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net181),
    .D(_0144_),
    .Q_N(_3013_),
    .Q(\core.leak_current[2] ));
 sg13g2_dfrbp_1 _6278_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net179),
    .D(_0145_),
    .Q_N(_3012_),
    .Q(\core.leak_current[3] ));
 sg13g2_dfrbp_1 _6279_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net177),
    .D(_0146_),
    .Q_N(_3011_),
    .Q(\core.leak_current[4] ));
 sg13g2_dfrbp_1 _6280_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net175),
    .D(_0147_),
    .Q_N(_3010_),
    .Q(\core.leak_current[5] ));
 sg13g2_dfrbp_1 _6281_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net173),
    .D(_0148_),
    .Q_N(_3009_),
    .Q(\core.leak_current[6] ));
 sg13g2_dfrbp_1 _6282_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net171),
    .D(_0149_),
    .Q_N(_3008_),
    .Q(\core.leak_current[7] ));
 sg13g2_dfrbp_1 _6283_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net169),
    .D(_0150_),
    .Q_N(_3007_),
    .Q(\core.leak_current[8] ));
 sg13g2_dfrbp_1 _6284_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net167),
    .D(_0151_),
    .Q_N(_3006_),
    .Q(\core.leak_current[9] ));
 sg13g2_dfrbp_1 _6285_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net165),
    .D(_0152_),
    .Q_N(_3005_),
    .Q(\core.leak_current[10] ));
 sg13g2_dfrbp_1 _6286_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net163),
    .D(_0153_),
    .Q_N(_3004_),
    .Q(\core.leak_current[11] ));
 sg13g2_dfrbp_1 _6287_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net161),
    .D(_0154_),
    .Q_N(_3003_),
    .Q(\core.leak_current[12] ));
 sg13g2_dfrbp_1 _6288_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net159),
    .D(_0155_),
    .Q_N(_3002_),
    .Q(\core.leak_current[13] ));
 sg13g2_dfrbp_1 _6289_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net157),
    .D(_0156_),
    .Q_N(_3001_),
    .Q(\core.leak_current[14] ));
 sg13g2_dfrbp_1 _6290_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net155),
    .D(_0157_),
    .Q_N(_3000_),
    .Q(\core.leak_current[15] ));
 sg13g2_dfrbp_1 _6291_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net153),
    .D(_0158_),
    .Q_N(_2999_),
    .Q(\core.ibias[8] ));
 sg13g2_dfrbp_1 _6292_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net151),
    .D(_0159_),
    .Q_N(_2998_),
    .Q(\core.ibias[9] ));
 sg13g2_dfrbp_1 _6293_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net149),
    .D(_0160_),
    .Q_N(_2997_),
    .Q(\core.ibias[10] ));
 sg13g2_dfrbp_1 _6294_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net147),
    .D(_0161_),
    .Q_N(_2996_),
    .Q(\core.ibias[11] ));
 sg13g2_dfrbp_1 _6295_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net145),
    .D(_0162_),
    .Q_N(_2995_),
    .Q(\core.ibias[12] ));
 sg13g2_dfrbp_1 _6296_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net143),
    .D(_0163_),
    .Q_N(_2994_),
    .Q(\core.ibias[13] ));
 sg13g2_dfrbp_1 _6297_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net141),
    .D(_0164_),
    .Q_N(_2993_),
    .Q(\core.ibias[14] ));
 sg13g2_dfrbp_1 _6298_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net140),
    .D(net321),
    .Q_N(_2992_),
    .Q(\core.ibias[15] ));
 sg13g2_dfrbp_1 _6299_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net138),
    .D(_0166_),
    .Q_N(_0012_),
    .Q(\core.delta_t[8] ));
 sg13g2_dfrbp_1 _6300_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net136),
    .D(_0167_),
    .Q_N(_0009_),
    .Q(\core.delta_t[9] ));
 sg13g2_dfrbp_1 _6301_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net134),
    .D(_0168_),
    .Q_N(_0010_),
    .Q(\core.delta_t[10] ));
 sg13g2_dfrbp_1 _6302_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net133),
    .D(_0169_),
    .Q_N(_0011_),
    .Q(\core.delta_t[11] ));
 sg13g2_dfrbp_1 _6303_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net131),
    .D(_0170_),
    .Q_N(_0013_),
    .Q(\core.delta_t[12] ));
 sg13g2_dfrbp_1 _6304_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net129),
    .D(_0171_),
    .Q_N(_0014_),
    .Q(\core.delta_t[13] ));
 sg13g2_dfrbp_1 _6305_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net127),
    .D(_0172_),
    .Q_N(_0015_),
    .Q(\core.delta_t[14] ));
 sg13g2_dfrbp_1 _6306_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net126),
    .D(net310),
    .Q_N(_2991_),
    .Q(\core.delta_t[15] ));
 sg13g2_dfrbp_1 _6307_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net118),
    .D(net473),
    .Q_N(_2990_),
    .Q(\core.temp_q[0] ));
 sg13g2_dfrbp_1 _6308_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net116),
    .D(_0175_),
    .Q_N(_2989_),
    .Q(\core.temp_q[1] ));
 sg13g2_dfrbp_1 _6309_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net114),
    .D(_0176_),
    .Q_N(_2988_),
    .Q(\core.temp_q[2] ));
 sg13g2_dfrbp_1 _6310_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net113),
    .D(_0177_),
    .Q_N(_2987_),
    .Q(\core.temp_q[3] ));
 sg13g2_dfrbp_1 _6311_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net111),
    .D(_0178_),
    .Q_N(_2986_),
    .Q(\core.temp_q[4] ));
 sg13g2_dfrbp_1 _6312_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net109),
    .D(_0179_),
    .Q_N(_2985_),
    .Q(\core.temp_q[5] ));
 sg13g2_dfrbp_1 _6313_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net107),
    .D(_0180_),
    .Q_N(_2984_),
    .Q(\core.temp_q[6] ));
 sg13g2_dfrbp_1 _6314_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net106),
    .D(_0181_),
    .Q_N(_0007_),
    .Q(\core.temp_q[7] ));
 sg13g2_dfrbp_1 _6315_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net104),
    .D(_0182_),
    .Q_N(_2983_),
    .Q(\core.temp_q[8] ));
 sg13g2_dfrbp_1 _6316_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net102),
    .D(_0183_),
    .Q_N(_2982_),
    .Q(\core.temp_q[9] ));
 sg13g2_dfrbp_1 _6317_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net100),
    .D(_0184_),
    .Q_N(_2981_),
    .Q(\core.temp_q[10] ));
 sg13g2_dfrbp_1 _6318_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net99),
    .D(_0185_),
    .Q_N(_2980_),
    .Q(\core.temp_q[11] ));
 sg13g2_dfrbp_1 _6319_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net97),
    .D(_0186_),
    .Q_N(_2979_),
    .Q(\core.temp_q[12] ));
 sg13g2_dfrbp_1 _6320_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net95),
    .D(_0187_),
    .Q_N(_2978_),
    .Q(\core.temp_q[13] ));
 sg13g2_dfrbp_1 _6321_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net93),
    .D(_0188_),
    .Q_N(_2977_),
    .Q(\core.temp_q[14] ));
 sg13g2_dfrbp_1 _6322_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net91),
    .D(_0189_),
    .Q_N(_0008_),
    .Q(\core.temp_q[15] ));
 sg13g2_dfrbp_1 _6323_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net89),
    .D(_0190_),
    .Q_N(_2976_),
    .Q(\core.w8_reg[2] ));
 sg13g2_dfrbp_1 _6324_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net87),
    .D(_0191_),
    .Q_N(_2975_),
    .Q(\core.w8_reg[3] ));
 sg13g2_dfrbp_1 _6325_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net85),
    .D(_0192_),
    .Q_N(_2974_),
    .Q(\core.w8_reg[4] ));
 sg13g2_dfrbp_1 _6326_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net83),
    .D(net385),
    .Q_N(_2973_),
    .Q(\core.w8_reg[5] ));
 sg13g2_dfrbp_1 _6327_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net81),
    .D(_0194_),
    .Q_N(_2972_),
    .Q(\core.w8_reg[6] ));
 sg13g2_dfrbp_1 _6328_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net72),
    .D(_0195_),
    .Q_N(_2971_),
    .Q(\core.w8_reg[7] ));
 sg13g2_dfrbp_1 _6329_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net70),
    .D(_0196_),
    .Q_N(_2970_),
    .Q(\core.vm8_reg[2] ));
 sg13g2_dfrbp_1 _6330_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net68),
    .D(_0197_),
    .Q_N(_2969_),
    .Q(\core.vm8_reg[3] ));
 sg13g2_dfrbp_1 _6331_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net66),
    .D(_0198_),
    .Q_N(_2968_),
    .Q(\core.vm8_reg[4] ));
 sg13g2_dfrbp_1 _6332_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net64),
    .D(_0199_),
    .Q_N(_2967_),
    .Q(\core.vm8_reg[5] ));
 sg13g2_dfrbp_1 _6333_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net62),
    .D(net331),
    .Q_N(_2966_),
    .Q(\core.vm8_reg[6] ));
 sg13g2_dfrbp_1 _6334_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net60),
    .D(_0201_),
    .Q_N(_2965_),
    .Q(\core.vm8_reg[7] ));
 sg13g2_dfrbp_1 _6335_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net58),
    .D(_0202_),
    .Q_N(_2964_),
    .Q(\core.dw[0] ));
 sg13g2_dfrbp_1 _6336_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net56),
    .D(_0203_),
    .Q_N(_2963_),
    .Q(\core.dw[1] ));
 sg13g2_dfrbp_1 _6337_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net54),
    .D(_0204_),
    .Q_N(_2962_),
    .Q(\core.dw[2] ));
 sg13g2_dfrbp_1 _6338_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net52),
    .D(_0205_),
    .Q_N(_2961_),
    .Q(\core.dw[3] ));
 sg13g2_dfrbp_1 _6339_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net50),
    .D(_0206_),
    .Q_N(_2960_),
    .Q(\core.dw[4] ));
 sg13g2_dfrbp_1 _6340_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net48),
    .D(_0207_),
    .Q_N(_2959_),
    .Q(\core.dw[5] ));
 sg13g2_dfrbp_1 _6341_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net46),
    .D(_0208_),
    .Q_N(_2958_),
    .Q(\core.dw[6] ));
 sg13g2_dfrbp_1 _6342_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net40),
    .D(_0209_),
    .Q_N(_2957_),
    .Q(\core.dw[7] ));
 sg13g2_dfrbp_1 _6343_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net36),
    .D(_0210_),
    .Q_N(_2956_),
    .Q(\core.dw[8] ));
 sg13g2_dfrbp_1 _6344_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net31),
    .D(_0211_),
    .Q_N(_2955_),
    .Q(\core.dw[9] ));
 sg13g2_dfrbp_1 _6345_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net27),
    .D(_0212_),
    .Q_N(_2954_),
    .Q(\core.dw[10] ));
 sg13g2_dfrbp_1 _6346_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net307),
    .D(_0213_),
    .Q_N(_2953_),
    .Q(\core.dw[11] ));
 sg13g2_dfrbp_1 _6347_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net303),
    .D(_0214_),
    .Q_N(_2952_),
    .Q(\core.dw[12] ));
 sg13g2_dfrbp_1 _6348_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net299),
    .D(_0215_),
    .Q_N(_2951_),
    .Q(\core.dw[13] ));
 sg13g2_dfrbp_1 _6349_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net295),
    .D(_0216_),
    .Q_N(_2950_),
    .Q(\core.dw[14] ));
 sg13g2_dfrbp_1 _6350_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net291),
    .D(_0217_),
    .Q_N(_2949_),
    .Q(\core.dw[15] ));
 sg13g2_dfrbp_1 _6351_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net287),
    .D(_0218_),
    .Q_N(_2948_),
    .Q(\core.dV[0] ));
 sg13g2_dfrbp_1 _6352_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net283),
    .D(_0219_),
    .Q_N(_2947_),
    .Q(\core.dV[1] ));
 sg13g2_dfrbp_1 _6353_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net279),
    .D(_0220_),
    .Q_N(_2946_),
    .Q(\core.dV[2] ));
 sg13g2_dfrbp_1 _6354_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net275),
    .D(_0221_),
    .Q_N(_2945_),
    .Q(\core.dV[3] ));
 sg13g2_dfrbp_1 _6355_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net271),
    .D(_0222_),
    .Q_N(_2944_),
    .Q(\core.dV[4] ));
 sg13g2_dfrbp_1 _6356_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net267),
    .D(_0223_),
    .Q_N(_2943_),
    .Q(\core.dV[5] ));
 sg13g2_dfrbp_1 _6357_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net263),
    .D(_0224_),
    .Q_N(_2942_),
    .Q(\core.dV[6] ));
 sg13g2_dfrbp_1 _6358_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net259),
    .D(_0225_),
    .Q_N(_2941_),
    .Q(\core.dV[7] ));
 sg13g2_dfrbp_1 _6359_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net255),
    .D(_0226_),
    .Q_N(_2940_),
    .Q(\core.dV[8] ));
 sg13g2_dfrbp_1 _6360_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net251),
    .D(_0227_),
    .Q_N(_2939_),
    .Q(\core.dV[9] ));
 sg13g2_dfrbp_1 _6361_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net247),
    .D(_0228_),
    .Q_N(_2938_),
    .Q(\core.dV[10] ));
 sg13g2_dfrbp_1 _6362_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net243),
    .D(_0229_),
    .Q_N(_2937_),
    .Q(\core.dV[11] ));
 sg13g2_dfrbp_1 _6363_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net239),
    .D(_0230_),
    .Q_N(_2936_),
    .Q(\core.dV[12] ));
 sg13g2_dfrbp_1 _6364_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net235),
    .D(_0231_),
    .Q_N(_2935_),
    .Q(\core.dV[13] ));
 sg13g2_dfrbp_1 _6365_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net231),
    .D(_0232_),
    .Q_N(_2934_),
    .Q(\core.dV[14] ));
 sg13g2_dfrbp_1 _6366_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net227),
    .D(_0233_),
    .Q_N(_2933_),
    .Q(\core.dV[15] ));
 sg13g2_dfrbp_1 _6367_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net214),
    .D(_0234_),
    .Q_N(_0032_),
    .Q(\core.drive_current[3] ));
 sg13g2_dfrbp_1 _6368_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net210),
    .D(_0235_),
    .Q_N(_0033_),
    .Q(\core.drive_current[4] ));
 sg13g2_dfrbp_1 _6369_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net190),
    .D(net555),
    .Q_N(_0034_),
    .Q(\core.drive_current[5] ));
 sg13g2_dfrbp_1 _6370_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net186),
    .D(net567),
    .Q_N(_0035_),
    .Q(\core.drive_current[6] ));
 sg13g2_dfrbp_1 _6371_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net182),
    .D(net561),
    .Q_N(_0036_),
    .Q(\core.drive_current[7] ));
 sg13g2_dfrbp_1 _6372_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net178),
    .D(_0239_),
    .Q_N(_0037_),
    .Q(\core.drive_current[8] ));
 sg13g2_dfrbp_1 _6373_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net174),
    .D(net564),
    .Q_N(_0038_),
    .Q(\core.drive_current[9] ));
 sg13g2_dfrbp_1 _6374_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net170),
    .D(_0241_),
    .Q_N(_0039_),
    .Q(\core.drive_current[10] ));
 sg13g2_dfrbp_1 _6375_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net166),
    .D(_0242_),
    .Q_N(_0040_),
    .Q(\core.drive_current[11] ));
 sg13g2_dfrbp_1 _6376_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net162),
    .D(net533),
    .Q_N(_0041_),
    .Q(\core.drive_current[12] ));
 sg13g2_dfrbp_1 _6377_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net158),
    .D(_0244_),
    .Q_N(_0042_),
    .Q(\core.drive_current[13] ));
 sg13g2_dfrbp_1 _6378_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net154),
    .D(_0245_),
    .Q_N(_0044_),
    .Q(\core.drive_current[14] ));
 sg13g2_dfrbp_1 _6379_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net150),
    .D(_0246_),
    .Q_N(_0043_),
    .Q(\core.drive_current[15] ));
 sg13g2_dfrbp_1 _6380_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net146),
    .D(_0247_),
    .Q_N(_2932_),
    .Q(\core.V_threshold[8] ));
 sg13g2_dfrbp_1 _6381_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net142),
    .D(_0248_),
    .Q_N(_2931_),
    .Q(\core.V_threshold[9] ));
 sg13g2_dfrbp_1 _6382_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net139),
    .D(_0249_),
    .Q_N(_2930_),
    .Q(\core.V_threshold[10] ));
 sg13g2_dfrbp_1 _6383_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net135),
    .D(_0250_),
    .Q_N(_2929_),
    .Q(\core.V_threshold[11] ));
 sg13g2_dfrbp_1 _6384_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net132),
    .D(_0251_),
    .Q_N(_2928_),
    .Q(\core.V_threshold[12] ));
 sg13g2_dfrbp_1 _6385_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net128),
    .D(_0252_),
    .Q_N(_2927_),
    .Q(\core.V_threshold[13] ));
 sg13g2_dfrbp_1 _6386_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net125),
    .D(_0253_),
    .Q_N(_2926_),
    .Q(\core.V_threshold[14] ));
 sg13g2_dfrbp_1 _6387_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net123),
    .D(net312),
    .Q_N(_2925_),
    .Q(\core.V_threshold[15] ));
 sg13g2_dfrbp_1 _6388_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net122),
    .D(_0255_),
    .Q_N(_2924_),
    .Q(\core.spike_reg ));
 sg13g2_dfrbp_1 _6389_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net120),
    .D(net884),
    .Q_N(_0018_),
    .Q(\core.w[0] ));
 sg13g2_dfrbp_1 _6390_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net119),
    .D(_0257_),
    .Q_N(_2923_),
    .Q(\core.w[1] ));
 sg13g2_dfrbp_1 _6391_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net115),
    .D(_0258_),
    .Q_N(_2922_),
    .Q(\core.w[2] ));
 sg13g2_dfrbp_1 _6392_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net112),
    .D(_0259_),
    .Q_N(_2921_),
    .Q(\core.w[3] ));
 sg13g2_dfrbp_1 _6393_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net108),
    .D(_0260_),
    .Q_N(_0019_),
    .Q(\core.w[4] ));
 sg13g2_dfrbp_1 _6394_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net105),
    .D(_0261_),
    .Q_N(_0020_),
    .Q(\core.w[5] ));
 sg13g2_dfrbp_1 _6395_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net101),
    .D(_0262_),
    .Q_N(_2920_),
    .Q(\core.w[6] ));
 sg13g2_dfrbp_1 _6396_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net98),
    .D(_0263_),
    .Q_N(_2919_),
    .Q(\core.w[7] ));
 sg13g2_dfrbp_1 _6397_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net94),
    .D(_0264_),
    .Q_N(_2918_),
    .Q(\core.w[8] ));
 sg13g2_dfrbp_1 _6398_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net90),
    .D(_0265_),
    .Q_N(_2917_),
    .Q(\core.w[9] ));
 sg13g2_dfrbp_1 _6399_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net86),
    .D(_0266_),
    .Q_N(_2916_),
    .Q(\core.w[10] ));
 sg13g2_dfrbp_1 _6400_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net82),
    .D(_0267_),
    .Q_N(_2915_),
    .Q(\core.w[11] ));
 sg13g2_dfrbp_1 _6401_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net71),
    .D(_0268_),
    .Q_N(_2914_),
    .Q(\core.w[12] ));
 sg13g2_dfrbp_1 _6402_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net67),
    .D(_0269_),
    .Q_N(_2913_),
    .Q(\core.w[13] ));
 sg13g2_dfrbp_1 _6403_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net63),
    .D(_0270_),
    .Q_N(_2912_),
    .Q(\core.w[14] ));
 sg13g2_dfrbp_1 _6404_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net59),
    .D(_0271_),
    .Q_N(_2911_),
    .Q(\core.w[15] ));
 sg13g2_dfrbp_1 _6405_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net55),
    .D(_0272_),
    .Q_N(_2910_),
    .Q(\core.V[0] ));
 sg13g2_dfrbp_1 _6406_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net51),
    .D(_0273_),
    .Q_N(_0029_),
    .Q(\core.V[1] ));
 sg13g2_dfrbp_1 _6407_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net47),
    .D(_0274_),
    .Q_N(_0024_),
    .Q(\core.V[2] ));
 sg13g2_dfrbp_1 _6408_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net38),
    .D(_0275_),
    .Q_N(_0023_),
    .Q(\core.V[3] ));
 sg13g2_dfrbp_1 _6409_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net29),
    .D(_0276_),
    .Q_N(_0025_),
    .Q(\core.V[4] ));
 sg13g2_dfrbp_1 _6410_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net305),
    .D(_0277_),
    .Q_N(_0026_),
    .Q(\core.V[5] ));
 sg13g2_dfrbp_1 _6411_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net297),
    .D(_0278_),
    .Q_N(_0027_),
    .Q(\core.V[6] ));
 sg13g2_dfrbp_1 _6412_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net289),
    .D(_0279_),
    .Q_N(_0028_),
    .Q(\core.V[7] ));
 sg13g2_dfrbp_1 _6413_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net281),
    .D(_0280_),
    .Q_N(_2909_),
    .Q(\core.V[8] ));
 sg13g2_dfrbp_1 _6414_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net273),
    .D(_0281_),
    .Q_N(_0052_),
    .Q(\core.V[9] ));
 sg13g2_dfrbp_1 _6415_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net265),
    .D(_0282_),
    .Q_N(_0053_),
    .Q(\core.V[10] ));
 sg13g2_dfrbp_1 _6416_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net257),
    .D(_0283_),
    .Q_N(_2908_),
    .Q(\core.V[11] ));
 sg13g2_dfrbp_1 _6417_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net249),
    .D(_0284_),
    .Q_N(_0021_),
    .Q(\core.V[12] ));
 sg13g2_dfrbp_1 _6418_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net241),
    .D(_0285_),
    .Q_N(_2907_),
    .Q(\core.V[13] ));
 sg13g2_dfrbp_1 _6419_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net233),
    .D(_0286_),
    .Q_N(_2906_),
    .Q(\core.V[14] ));
 sg13g2_dfrbp_1 _6420_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net225),
    .D(_0287_),
    .Q_N(_2905_),
    .Q(\core.V[15] ));
 sg13g2_dfrbp_1 _6421_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net219),
    .D(_0288_),
    .Q_N(_2904_),
    .Q(\core.params[5][0] ));
 sg13g2_dfrbp_1 _6422_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net212),
    .D(net383),
    .Q_N(_2903_),
    .Q(\core.params[5][1] ));
 sg13g2_dfrbp_1 _6423_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net188),
    .D(net377),
    .Q_N(_2902_),
    .Q(\core.params[5][2] ));
 sg13g2_dfrbp_1 _6424_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net180),
    .D(_0291_),
    .Q_N(_2901_),
    .Q(\core.params[5][3] ));
 sg13g2_dfrbp_1 _6425_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net172),
    .D(_0292_),
    .Q_N(_2900_),
    .Q(\core.params[5][4] ));
 sg13g2_dfrbp_1 _6426_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net164),
    .D(_0293_),
    .Q_N(_2899_),
    .Q(\core.params[5][5] ));
 sg13g2_dfrbp_1 _6427_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net156),
    .D(net375),
    .Q_N(_2898_),
    .Q(\core.params[5][6] ));
 sg13g2_dfrbp_1 _6428_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net148),
    .D(_0295_),
    .Q_N(_2856_),
    .Q(\core.params[5][7] ));
 sg13g2_dfrbp_1 _6429_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net92),
    .D(_0296_),
    .Q_N(_2897_),
    .Q(\core.params[3][0] ));
 sg13g2_dfrbp_1 _6430_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net84),
    .D(_0297_),
    .Q_N(_2896_),
    .Q(\core.params[3][1] ));
 sg13g2_dfrbp_1 _6431_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net69),
    .D(_0298_),
    .Q_N(_2895_),
    .Q(\core.params[3][2] ));
 sg13g2_dfrbp_1 _6432_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net61),
    .D(net450),
    .Q_N(_2894_),
    .Q(\core.params[3][3] ));
 sg13g2_dfrbp_1 _6433_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net53),
    .D(_0300_),
    .Q_N(_2893_),
    .Q(\core.params[3][4] ));
 sg13g2_dfrbp_1 _6434_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net42),
    .D(net416),
    .Q_N(_2892_),
    .Q(\core.params[3][5] ));
 sg13g2_dfrbp_1 _6435_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net25),
    .D(_0302_),
    .Q_N(_2891_),
    .Q(\core.params[3][6] ));
 sg13g2_dfrbp_1 _6436_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net293),
    .D(net437),
    .Q_N(_2890_),
    .Q(\core.params[3][7] ));
 sg13g2_dfrbp_1 _6437_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net277),
    .D(_0304_),
    .Q_N(_2889_),
    .Q(\core.params[2][0] ));
 sg13g2_dfrbp_1 _6438_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net261),
    .D(net402),
    .Q_N(_2888_),
    .Q(\core.params[2][1] ));
 sg13g2_dfrbp_1 _6439_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net245),
    .D(_0306_),
    .Q_N(_2887_),
    .Q(\core.params[2][2] ));
 sg13g2_dfrbp_1 _6440_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net229),
    .D(_0307_),
    .Q_N(_2886_),
    .Q(\core.params[2][3] ));
 sg13g2_dfrbp_1 _6441_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net216),
    .D(_0308_),
    .Q_N(_2885_),
    .Q(\core.params[2][4] ));
 sg13g2_dfrbp_1 _6442_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net184),
    .D(_0309_),
    .Q_N(_2884_),
    .Q(\core.params[2][5] ));
 sg13g2_dfrbp_1 _6443_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net168),
    .D(_0310_),
    .Q_N(_2883_),
    .Q(\core.params[2][6] ));
 sg13g2_dfrbp_1 _6444_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net152),
    .D(net414),
    .Q_N(_2882_),
    .Q(\core.params[2][7] ));
 sg13g2_dfrbp_1 _6445_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net137),
    .D(_0312_),
    .Q_N(_2881_),
    .Q(\core.params[1][0] ));
 sg13g2_dfrbp_1 _6446_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net124),
    .D(_0313_),
    .Q_N(_2880_),
    .Q(\core.params[1][1] ));
 sg13g2_dfrbp_1 _6447_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net117),
    .D(net407),
    .Q_N(_2879_),
    .Q(\core.params[1][2] ));
 sg13g2_dfrbp_1 _6448_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net103),
    .D(_0315_),
    .Q_N(_2878_),
    .Q(\core.params[1][3] ));
 sg13g2_dfrbp_1 _6449_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net88),
    .D(_0316_),
    .Q_N(_2877_),
    .Q(\core.params[1][4] ));
 sg13g2_dfrbp_1 _6450_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net65),
    .D(net446),
    .Q_N(_2876_),
    .Q(\core.params[1][5] ));
 sg13g2_dfrbp_1 _6451_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net49),
    .D(net460),
    .Q_N(_2875_),
    .Q(\core.params[1][6] ));
 sg13g2_dfrbp_1 _6452_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net301),
    .D(net477),
    .Q_N(_2874_),
    .Q(\core.params[1][7] ));
 sg13g2_dfrbp_1 _6453_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net269),
    .D(_0320_),
    .Q_N(_2873_),
    .Q(\core.exp_term[1] ));
 sg13g2_dfrbp_1 _6454_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net237),
    .D(_0321_),
    .Q_N(_2872_),
    .Q(\core.exp_term[2] ));
 sg13g2_dfrbp_1 _6455_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net208),
    .D(_0322_),
    .Q_N(_2871_),
    .Q(\core.exp_term[3] ));
 sg13g2_dfrbp_1 _6456_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net160),
    .D(_0323_),
    .Q_N(_2870_),
    .Q(\core.exp_term[4] ));
 sg13g2_dfrbp_1 _6457_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net130),
    .D(_0324_),
    .Q_N(_2869_),
    .Q(\core.exp_term[5] ));
 sg13g2_dfrbp_1 _6458_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net110),
    .D(_0325_),
    .Q_N(_2868_),
    .Q(\core.exp_term[6] ));
 sg13g2_dfrbp_1 _6459_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net80),
    .D(_0326_),
    .Q_N(_2867_),
    .Q(\core.exp_term[7] ));
 sg13g2_dfrbp_1 _6460_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net33),
    .D(_0327_),
    .Q_N(_2866_),
    .Q(\core.exp_term[8] ));
 sg13g2_dfrbp_1 _6461_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net253),
    .D(_0328_),
    .Q_N(_2865_),
    .Q(\core.exp_term[9] ));
 sg13g2_dfrbp_1 _6462_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net176),
    .D(_0329_),
    .Q_N(_2864_),
    .Q(\core.exp_term[10] ));
 sg13g2_dfrbp_1 _6463_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net121),
    .D(_0330_),
    .Q_N(_2863_),
    .Q(\core.exp_term[11] ));
 sg13g2_dfrbp_1 _6464_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net57),
    .D(_0331_),
    .Q_N(_2862_),
    .Q(\core.exp_term[12] ));
 sg13g2_dfrbp_1 _6465_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net222),
    .D(_0332_),
    .Q_N(_2861_),
    .Q(\core.exp_term[13] ));
 sg13g2_dfrbp_1 _6466_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net96),
    .D(_0333_),
    .Q_N(_2860_),
    .Q(\core.exp_term[14] ));
 sg13g2_dfrbp_1 _6467_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net144),
    .D(_0334_),
    .Q_N(_2859_),
    .Q(\core.exp_term[15] ));
 sg13g2_tiehi _6196__26 (.L_HI(net26));
 sg13g2_tiehi _6345__27 (.L_HI(net27));
 sg13g2_tiehi _6195__28 (.L_HI(net28));
 sg13g2_tiehi _6409__29 (.L_HI(net29));
 sg13g2_tiehi _6194__30 (.L_HI(net30));
 sg13g2_tiehi _6344__31 (.L_HI(net31));
 sg13g2_tiehi _6193__32 (.L_HI(net32));
 sg13g2_tiehi _6460__33 (.L_HI(net33));
 sg13g2_tiehi _6192__34 (.L_HI(net34));
 sg13g2_tiehi _6191__35 (.L_HI(net35));
 sg13g2_tiehi _6343__36 (.L_HI(net36));
 sg13g2_tiehi _6190__37 (.L_HI(net37));
 sg13g2_tiehi _6408__38 (.L_HI(net38));
 sg13g2_tiehi _6189__39 (.L_HI(net39));
 sg13g2_tiehi _6342__40 (.L_HI(net40));
 sg13g2_tiehi _6188__41 (.L_HI(net41));
 sg13g2_tiehi _6434__42 (.L_HI(net42));
 sg13g2_tiehi _6187__43 (.L_HI(net43));
 sg13g2_tiehi _6186__44 (.L_HI(net44));
 sg13g2_tiehi _6185__45 (.L_HI(net45));
 sg13g2_tiehi _6341__46 (.L_HI(net46));
 sg13g2_tiehi _6407__47 (.L_HI(net47));
 sg13g2_tiehi _6340__48 (.L_HI(net48));
 sg13g2_tiehi _6451__49 (.L_HI(net49));
 sg13g2_tiehi _6339__50 (.L_HI(net50));
 sg13g2_tiehi _6406__51 (.L_HI(net51));
 sg13g2_tiehi _6338__52 (.L_HI(net52));
 sg13g2_tiehi _6433__53 (.L_HI(net53));
 sg13g2_tiehi _6337__54 (.L_HI(net54));
 sg13g2_tiehi _6405__55 (.L_HI(net55));
 sg13g2_tiehi _6336__56 (.L_HI(net56));
 sg13g2_tiehi _6464__57 (.L_HI(net57));
 sg13g2_tiehi _6335__58 (.L_HI(net58));
 sg13g2_tiehi _6404__59 (.L_HI(net59));
 sg13g2_tiehi _6334__60 (.L_HI(net60));
 sg13g2_tiehi _6432__61 (.L_HI(net61));
 sg13g2_tiehi _6333__62 (.L_HI(net62));
 sg13g2_tiehi _6403__63 (.L_HI(net63));
 sg13g2_tiehi _6332__64 (.L_HI(net64));
 sg13g2_tiehi _6450__65 (.L_HI(net65));
 sg13g2_tiehi _6331__66 (.L_HI(net66));
 sg13g2_tiehi _6402__67 (.L_HI(net67));
 sg13g2_tiehi _6330__68 (.L_HI(net68));
 sg13g2_tiehi _6431__69 (.L_HI(net69));
 sg13g2_tiehi _6329__70 (.L_HI(net70));
 sg13g2_tiehi _6401__71 (.L_HI(net71));
 sg13g2_tiehi _6328__72 (.L_HI(net72));
 sg13g2_tiehi _6184__73 (.L_HI(net73));
 sg13g2_tiehi _6231__74 (.L_HI(net74));
 sg13g2_tiehi _6232__75 (.L_HI(net75));
 sg13g2_tiehi _6233__76 (.L_HI(net76));
 sg13g2_tiehi _6234__77 (.L_HI(net77));
 sg13g2_tiehi _6235__78 (.L_HI(net78));
 sg13g2_tiehi _6236__79 (.L_HI(net79));
 sg13g2_tiehi _6459__80 (.L_HI(net80));
 sg13g2_tiehi _6327__81 (.L_HI(net81));
 sg13g2_tiehi _6400__82 (.L_HI(net82));
 sg13g2_tiehi _6326__83 (.L_HI(net83));
 sg13g2_tiehi _6430__84 (.L_HI(net84));
 sg13g2_tiehi _6325__85 (.L_HI(net85));
 sg13g2_tiehi _6399__86 (.L_HI(net86));
 sg13g2_tiehi _6324__87 (.L_HI(net87));
 sg13g2_tiehi _6449__88 (.L_HI(net88));
 sg13g2_tiehi _6323__89 (.L_HI(net89));
 sg13g2_tiehi _6398__90 (.L_HI(net90));
 sg13g2_tiehi _6322__91 (.L_HI(net91));
 sg13g2_tiehi _6429__92 (.L_HI(net92));
 sg13g2_tiehi _6321__93 (.L_HI(net93));
 sg13g2_tiehi _6397__94 (.L_HI(net94));
 sg13g2_tiehi _6320__95 (.L_HI(net95));
 sg13g2_tiehi _6466__96 (.L_HI(net96));
 sg13g2_tiehi _6319__97 (.L_HI(net97));
 sg13g2_tiehi _6396__98 (.L_HI(net98));
 sg13g2_tiehi _6318__99 (.L_HI(net99));
 sg13g2_tiehi _6317__100 (.L_HI(net100));
 sg13g2_tiehi _6395__101 (.L_HI(net101));
 sg13g2_tiehi _6316__102 (.L_HI(net102));
 sg13g2_tiehi _6448__103 (.L_HI(net103));
 sg13g2_tiehi _6315__104 (.L_HI(net104));
 sg13g2_tiehi _6394__105 (.L_HI(net105));
 sg13g2_tiehi _6314__106 (.L_HI(net106));
 sg13g2_tiehi _6313__107 (.L_HI(net107));
 sg13g2_tiehi _6393__108 (.L_HI(net108));
 sg13g2_tiehi _6312__109 (.L_HI(net109));
 sg13g2_tiehi _6458__110 (.L_HI(net110));
 sg13g2_tiehi _6311__111 (.L_HI(net111));
 sg13g2_tiehi _6392__112 (.L_HI(net112));
 sg13g2_tiehi _6310__113 (.L_HI(net113));
 sg13g2_tiehi _6309__114 (.L_HI(net114));
 sg13g2_tiehi _6391__115 (.L_HI(net115));
 sg13g2_tiehi _6308__116 (.L_HI(net116));
 sg13g2_tiehi _6447__117 (.L_HI(net117));
 sg13g2_tiehi _6307__118 (.L_HI(net118));
 sg13g2_tiehi _6390__119 (.L_HI(net119));
 sg13g2_tiehi _6389__120 (.L_HI(net120));
 sg13g2_tiehi _6463__121 (.L_HI(net121));
 sg13g2_tiehi _6388__122 (.L_HI(net122));
 sg13g2_tiehi _6387__123 (.L_HI(net123));
 sg13g2_tiehi _6446__124 (.L_HI(net124));
 sg13g2_tiehi _6386__125 (.L_HI(net125));
 sg13g2_tiehi _6306__126 (.L_HI(net126));
 sg13g2_tiehi _6305__127 (.L_HI(net127));
 sg13g2_tiehi _6385__128 (.L_HI(net128));
 sg13g2_tiehi _6304__129 (.L_HI(net129));
 sg13g2_tiehi _6457__130 (.L_HI(net130));
 sg13g2_tiehi _6303__131 (.L_HI(net131));
 sg13g2_tiehi _6384__132 (.L_HI(net132));
 sg13g2_tiehi _6302__133 (.L_HI(net133));
 sg13g2_tiehi _6301__134 (.L_HI(net134));
 sg13g2_tiehi _6383__135 (.L_HI(net135));
 sg13g2_tiehi _6300__136 (.L_HI(net136));
 sg13g2_tiehi _6445__137 (.L_HI(net137));
 sg13g2_tiehi _6299__138 (.L_HI(net138));
 sg13g2_tiehi _6382__139 (.L_HI(net139));
 sg13g2_tiehi _6298__140 (.L_HI(net140));
 sg13g2_tiehi _6297__141 (.L_HI(net141));
 sg13g2_tiehi _6381__142 (.L_HI(net142));
 sg13g2_tiehi _6296__143 (.L_HI(net143));
 sg13g2_tiehi _6467__144 (.L_HI(net144));
 sg13g2_tiehi _6295__145 (.L_HI(net145));
 sg13g2_tiehi _6380__146 (.L_HI(net146));
 sg13g2_tiehi _6294__147 (.L_HI(net147));
 sg13g2_tiehi _6428__148 (.L_HI(net148));
 sg13g2_tiehi _6293__149 (.L_HI(net149));
 sg13g2_tiehi _6379__150 (.L_HI(net150));
 sg13g2_tiehi _6292__151 (.L_HI(net151));
 sg13g2_tiehi _6444__152 (.L_HI(net152));
 sg13g2_tiehi _6291__153 (.L_HI(net153));
 sg13g2_tiehi _6378__154 (.L_HI(net154));
 sg13g2_tiehi _6290__155 (.L_HI(net155));
 sg13g2_tiehi _6427__156 (.L_HI(net156));
 sg13g2_tiehi _6289__157 (.L_HI(net157));
 sg13g2_tiehi _6377__158 (.L_HI(net158));
 sg13g2_tiehi _6288__159 (.L_HI(net159));
 sg13g2_tiehi _6456__160 (.L_HI(net160));
 sg13g2_tiehi _6287__161 (.L_HI(net161));
 sg13g2_tiehi _6376__162 (.L_HI(net162));
 sg13g2_tiehi _6286__163 (.L_HI(net163));
 sg13g2_tiehi _6426__164 (.L_HI(net164));
 sg13g2_tiehi _6285__165 (.L_HI(net165));
 sg13g2_tiehi _6375__166 (.L_HI(net166));
 sg13g2_tiehi _6284__167 (.L_HI(net167));
 sg13g2_tiehi _6443__168 (.L_HI(net168));
 sg13g2_tiehi _6283__169 (.L_HI(net169));
 sg13g2_tiehi _6374__170 (.L_HI(net170));
 sg13g2_tiehi _6282__171 (.L_HI(net171));
 sg13g2_tiehi _6425__172 (.L_HI(net172));
 sg13g2_tiehi _6281__173 (.L_HI(net173));
 sg13g2_tiehi _6373__174 (.L_HI(net174));
 sg13g2_tiehi _6280__175 (.L_HI(net175));
 sg13g2_tiehi _6462__176 (.L_HI(net176));
 sg13g2_tiehi _6279__177 (.L_HI(net177));
 sg13g2_tiehi _6372__178 (.L_HI(net178));
 sg13g2_tiehi _6278__179 (.L_HI(net179));
 sg13g2_tiehi _6424__180 (.L_HI(net180));
 sg13g2_tiehi _6277__181 (.L_HI(net181));
 sg13g2_tiehi _6371__182 (.L_HI(net182));
 sg13g2_tiehi _6276__183 (.L_HI(net183));
 sg13g2_tiehi _6442__184 (.L_HI(net184));
 sg13g2_tiehi _6275__185 (.L_HI(net185));
 sg13g2_tiehi _6370__186 (.L_HI(net186));
 sg13g2_tiehi _6274__187 (.L_HI(net187));
 sg13g2_tiehi _6423__188 (.L_HI(net188));
 sg13g2_tiehi _6273__189 (.L_HI(net189));
 sg13g2_tiehi _6369__190 (.L_HI(net190));
 sg13g2_tiehi _6272__191 (.L_HI(net191));
 sg13g2_tiehi _6271__192 (.L_HI(net192));
 sg13g2_tiehi _6270__193 (.L_HI(net193));
 sg13g2_tiehi _6269__194 (.L_HI(net194));
 sg13g2_tiehi _6268__195 (.L_HI(net195));
 sg13g2_tiehi _6267__196 (.L_HI(net196));
 sg13g2_tiehi _6266__197 (.L_HI(net197));
 sg13g2_tiehi _6265__198 (.L_HI(net198));
 sg13g2_tiehi _6264__199 (.L_HI(net199));
 sg13g2_tiehi _6263__200 (.L_HI(net200));
 sg13g2_tiehi _6262__201 (.L_HI(net201));
 sg13g2_tiehi _6261__202 (.L_HI(net202));
 sg13g2_tiehi _6260__203 (.L_HI(net203));
 sg13g2_tiehi _6259__204 (.L_HI(net204));
 sg13g2_tiehi _6258__205 (.L_HI(net205));
 sg13g2_tiehi _6257__206 (.L_HI(net206));
 sg13g2_tiehi _6256__207 (.L_HI(net207));
 sg13g2_tiehi _6455__208 (.L_HI(net208));
 sg13g2_tiehi _6255__209 (.L_HI(net209));
 sg13g2_tiehi _6368__210 (.L_HI(net210));
 sg13g2_tiehi _6254__211 (.L_HI(net211));
 sg13g2_tiehi _6422__212 (.L_HI(net212));
 sg13g2_tiehi _6253__213 (.L_HI(net213));
 sg13g2_tiehi _6367__214 (.L_HI(net214));
 sg13g2_tiehi _6252__215 (.L_HI(net215));
 sg13g2_tiehi _6441__216 (.L_HI(net216));
 sg13g2_tiehi _6251__217 (.L_HI(net217));
 sg13g2_tiehi _6250__218 (.L_HI(net218));
 sg13g2_tiehi _6421__219 (.L_HI(net219));
 sg13g2_tiehi _6249__220 (.L_HI(net220));
 sg13g2_tiehi _6248__221 (.L_HI(net221));
 sg13g2_tiehi _6465__222 (.L_HI(net222));
 sg13g2_tiehi _6247__223 (.L_HI(net223));
 sg13g2_tiehi _6246__224 (.L_HI(net224));
 sg13g2_tiehi _6420__225 (.L_HI(net225));
 sg13g2_tiehi _6245__226 (.L_HI(net226));
 sg13g2_tiehi _6366__227 (.L_HI(net227));
 sg13g2_tiehi _6244__228 (.L_HI(net228));
 sg13g2_tiehi _6440__229 (.L_HI(net229));
 sg13g2_tiehi _6243__230 (.L_HI(net230));
 sg13g2_tiehi _6365__231 (.L_HI(net231));
 sg13g2_tiehi _6242__232 (.L_HI(net232));
 sg13g2_tiehi _6419__233 (.L_HI(net233));
 sg13g2_tiehi _6241__234 (.L_HI(net234));
 sg13g2_tiehi _6364__235 (.L_HI(net235));
 sg13g2_tiehi _6240__236 (.L_HI(net236));
 sg13g2_tiehi _6454__237 (.L_HI(net237));
 sg13g2_tiehi _6239__238 (.L_HI(net238));
 sg13g2_tiehi _6363__239 (.L_HI(net239));
 sg13g2_tiehi _6238__240 (.L_HI(net240));
 sg13g2_tiehi _6418__241 (.L_HI(net241));
 sg13g2_tiehi _6230__242 (.L_HI(net242));
 sg13g2_tiehi _6362__243 (.L_HI(net243));
 sg13g2_tiehi _6229__244 (.L_HI(net244));
 sg13g2_tiehi _6439__245 (.L_HI(net245));
 sg13g2_tiehi _6228__246 (.L_HI(net246));
 sg13g2_tiehi _6361__247 (.L_HI(net247));
 sg13g2_tiehi _6227__248 (.L_HI(net248));
 sg13g2_tiehi _6417__249 (.L_HI(net249));
 sg13g2_tiehi _6226__250 (.L_HI(net250));
 sg13g2_tiehi _6360__251 (.L_HI(net251));
 sg13g2_tiehi _6225__252 (.L_HI(net252));
 sg13g2_tiehi _6461__253 (.L_HI(net253));
 sg13g2_tiehi _6224__254 (.L_HI(net254));
 sg13g2_tiehi _6359__255 (.L_HI(net255));
 sg13g2_tiehi _6223__256 (.L_HI(net256));
 sg13g2_tiehi _6416__257 (.L_HI(net257));
 sg13g2_tiehi _6222__258 (.L_HI(net258));
 sg13g2_tiehi _6358__259 (.L_HI(net259));
 sg13g2_tiehi _6221__260 (.L_HI(net260));
 sg13g2_tiehi _6438__261 (.L_HI(net261));
 sg13g2_tiehi _6220__262 (.L_HI(net262));
 sg13g2_tiehi _6357__263 (.L_HI(net263));
 sg13g2_tiehi _6219__264 (.L_HI(net264));
 sg13g2_tiehi _6415__265 (.L_HI(net265));
 sg13g2_tiehi _6218__266 (.L_HI(net266));
 sg13g2_tiehi _6356__267 (.L_HI(net267));
 sg13g2_tiehi _6217__268 (.L_HI(net268));
 sg13g2_tiehi _6453__269 (.L_HI(net269));
 sg13g2_tiehi _6216__270 (.L_HI(net270));
 sg13g2_tiehi _6355__271 (.L_HI(net271));
 sg13g2_tiehi _6215__272 (.L_HI(net272));
 sg13g2_tiehi _6414__273 (.L_HI(net273));
 sg13g2_tiehi _6214__274 (.L_HI(net274));
 sg13g2_tiehi _6354__275 (.L_HI(net275));
 sg13g2_tiehi _6213__276 (.L_HI(net276));
 sg13g2_tiehi _6437__277 (.L_HI(net277));
 sg13g2_tiehi _6212__278 (.L_HI(net278));
 sg13g2_tiehi _6353__279 (.L_HI(net279));
 sg13g2_tiehi _6211__280 (.L_HI(net280));
 sg13g2_tiehi _6413__281 (.L_HI(net281));
 sg13g2_tiehi _6210__282 (.L_HI(net282));
 sg13g2_tiehi _6352__283 (.L_HI(net283));
 sg13g2_tiehi _6209__284 (.L_HI(net284));
 sg13g2_tiehi _6237__285 (.L_HI(net285));
 sg13g2_tiehi _6208__286 (.L_HI(net286));
 sg13g2_tiehi _6351__287 (.L_HI(net287));
 sg13g2_tiehi _6207__288 (.L_HI(net288));
 sg13g2_tiehi _6412__289 (.L_HI(net289));
 sg13g2_tiehi _6206__290 (.L_HI(net290));
 sg13g2_tiehi _6350__291 (.L_HI(net291));
 sg13g2_tiehi _6205__292 (.L_HI(net292));
 sg13g2_tiehi _6436__293 (.L_HI(net293));
 sg13g2_tiehi _6204__294 (.L_HI(net294));
 sg13g2_tiehi _6349__295 (.L_HI(net295));
 sg13g2_tiehi _6203__296 (.L_HI(net296));
 sg13g2_tiehi _6411__297 (.L_HI(net297));
 sg13g2_tiehi _6202__298 (.L_HI(net298));
 sg13g2_tiehi _6348__299 (.L_HI(net299));
 sg13g2_tiehi _6201__300 (.L_HI(net300));
 sg13g2_tiehi _6452__301 (.L_HI(net301));
 sg13g2_tiehi _6200__302 (.L_HI(net302));
 sg13g2_tiehi _6347__303 (.L_HI(net303));
 sg13g2_tiehi _6199__304 (.L_HI(net304));
 sg13g2_tiehi _6410__305 (.L_HI(net305));
 sg13g2_tiehi _6198__306 (.L_HI(net306));
 sg13g2_tiehi _6346__307 (.L_HI(net307));
 sg13g2_tiehi _6197__308 (.L_HI(net308));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_dpi_adexp_9 (.L_LO(net9));
 sg13g2_tielo tt_um_dpi_adexp_10 (.L_LO(net10));
 sg13g2_tielo tt_um_dpi_adexp_11 (.L_LO(net11));
 sg13g2_tielo tt_um_dpi_adexp_12 (.L_LO(net12));
 sg13g2_tielo tt_um_dpi_adexp_13 (.L_LO(net13));
 sg13g2_tielo tt_um_dpi_adexp_14 (.L_LO(net14));
 sg13g2_tielo tt_um_dpi_adexp_15 (.L_LO(net15));
 sg13g2_tielo tt_um_dpi_adexp_16 (.L_LO(net16));
 sg13g2_tielo tt_um_dpi_adexp_17 (.L_LO(net17));
 sg13g2_tielo tt_um_dpi_adexp_18 (.L_LO(net18));
 sg13g2_tielo tt_um_dpi_adexp_19 (.L_LO(net19));
 sg13g2_tielo tt_um_dpi_adexp_20 (.L_LO(net20));
 sg13g2_tielo tt_um_dpi_adexp_21 (.L_LO(net21));
 sg13g2_tielo tt_um_dpi_adexp_22 (.L_LO(net22));
 sg13g2_tielo tt_um_dpi_adexp_23 (.L_LO(net23));
 sg13g2_tielo tt_um_dpi_adexp_24 (.L_LO(net24));
 sg13g2_tiehi _6435__25 (.L_HI(net25));
 sg13g2_buf_2 _6769_ (.A(\core.spike_reg ),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout569 (.A(net570),
    .X(net569));
 sg13g2_buf_1 fanout570 (.A(_1817_),
    .X(net570));
 sg13g2_buf_4 fanout571 (.X(net571),
    .A(_1841_));
 sg13g2_buf_2 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_1523_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net575),
    .X(net574));
 sg13g2_buf_1 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(_0849_));
 sg13g2_buf_2 fanout577 (.A(_0846_),
    .X(net577));
 sg13g2_buf_1 fanout578 (.A(_0846_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net581),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_0565_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_0845_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_0587_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_0562_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_0562_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_1226_),
    .X(net586));
 sg13g2_buf_4 fanout587 (.X(net587),
    .A(_2198_));
 sg13g2_buf_4 fanout588 (.X(net588),
    .A(_2097_));
 sg13g2_buf_2 fanout589 (.A(_2097_),
    .X(net589));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(_1990_));
 sg13g2_buf_2 fanout591 (.A(_1529_),
    .X(net591));
 sg13g2_buf_4 fanout592 (.X(net592),
    .A(_1518_));
 sg13g2_buf_4 fanout593 (.X(net593),
    .A(_0549_));
 sg13g2_buf_1 fanout594 (.A(_0549_),
    .X(net594));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(_2002_));
 sg13g2_buf_2 fanout596 (.A(_1992_),
    .X(net596));
 sg13g2_buf_1 fanout597 (.A(_1992_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(_1950_));
 sg13g2_buf_4 fanout600 (.X(net600),
    .A(_0546_));
 sg13g2_buf_2 fanout601 (.A(_0546_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(net604),
    .X(net602));
 sg13g2_buf_1 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_2753_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_1944_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_1936_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_1929_),
    .X(net607));
 sg13g2_buf_4 fanout608 (.X(net608),
    .A(_1922_));
 sg13g2_buf_2 fanout609 (.A(net610),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(net611),
    .X(net610));
 sg13g2_buf_4 fanout611 (.X(net611),
    .A(_0555_));
 sg13g2_buf_4 fanout612 (.X(net612),
    .A(net613));
 sg13g2_buf_4 fanout613 (.X(net613),
    .A(_0553_));
 sg13g2_buf_2 fanout614 (.A(_0345_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_0335_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_2849_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_2808_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_1980_),
    .X(net618));
 sg13g2_buf_4 fanout619 (.X(net619),
    .A(_0576_));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(net621));
 sg13g2_buf_4 fanout621 (.X(net621),
    .A(_0579_));
 sg13g2_buf_4 fanout622 (.X(net622),
    .A(_0342_));
 sg13g2_buf_4 fanout623 (.X(net623),
    .A(_2005_));
 sg13g2_buf_1 fanout624 (.A(_2005_),
    .X(net624));
 sg13g2_buf_4 fanout625 (.X(net625),
    .A(net627));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(net627));
 sg13g2_buf_2 fanout627 (.A(_1820_),
    .X(net627));
 sg13g2_buf_4 fanout628 (.X(net628),
    .A(_0701_));
 sg13g2_buf_4 fanout629 (.X(net629),
    .A(net630));
 sg13g2_buf_4 fanout630 (.X(net630),
    .A(_0700_));
 sg13g2_buf_2 fanout631 (.A(_2781_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_2777_),
    .X(net633));
 sg13g2_buf_4 fanout634 (.X(net634),
    .A(_0698_));
 sg13g2_buf_2 fanout635 (.A(net637),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(net637),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_2754_),
    .X(net637));
 sg13g2_buf_4 fanout638 (.X(net638),
    .A(net640));
 sg13g2_buf_1 fanout639 (.A(net640),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_2751_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(net645),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(net643),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net645),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_4 fanout645 (.X(net645),
    .A(_2750_));
 sg13g2_buf_2 fanout646 (.A(net648),
    .X(net646));
 sg13g2_buf_1 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(_2749_));
 sg13g2_buf_2 fanout649 (.A(_2743_),
    .X(net649));
 sg13g2_buf_1 fanout650 (.A(_2743_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_2674_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_2674_),
    .X(net652));
 sg13g2_buf_4 fanout653 (.X(net653),
    .A(\core.V[13] ));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(net872));
 sg13g2_buf_4 fanout655 (.X(net655),
    .A(net880));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(net889));
 sg13g2_buf_2 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(net659),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(\core.V[9] ),
    .X(net659));
 sg13g2_buf_4 fanout660 (.X(net660),
    .A(net661));
 sg13g2_buf_4 fanout661 (.X(net661),
    .A(\core.V[8] ));
 sg13g2_buf_4 fanout662 (.X(net662),
    .A(\core.V[7] ));
 sg13g2_buf_2 fanout663 (.A(net858),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(net665),
    .X(net664));
 sg13g2_buf_4 fanout665 (.X(net665),
    .A(net846));
 sg13g2_buf_4 fanout666 (.X(net666),
    .A(net667));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(net851));
 sg13g2_buf_2 fanout668 (.A(net669),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(net868),
    .X(net669));
 sg13g2_buf_4 fanout670 (.X(net670),
    .A(net671));
 sg13g2_buf_2 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(net849),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(net674),
    .X(net673));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(net845));
 sg13g2_buf_2 fanout675 (.A(net870),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(\core.V[1] ),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(net679),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(net679),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(\core.V[0] ),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(net681),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(\core.delta_t[15] ),
    .X(net681));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(net683));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(\core.delta_t[8] ));
 sg13g2_buf_2 fanout684 (.A(net879),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(\core.param_idx[1] ),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(net696),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(net689),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_1 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(net696),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(net696),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(\core.r_ready ),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(net700),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(net700),
    .X(net698));
 sg13g2_buf_1 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(\core.r_ready ),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(net704),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(net704),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(net704),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(\core.r_ready ),
    .X(net704));
 sg13g2_buf_4 fanout705 (.X(net705),
    .A(\core.param_a[14] ));
 sg13g2_buf_2 fanout706 (.A(net707),
    .X(net706));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(net424));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(\core.param_a[12] ));
 sg13g2_buf_2 fanout709 (.A(\core.param_a[12] ),
    .X(net709));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(net711));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(\core.param_a[11] ));
 sg13g2_buf_2 fanout712 (.A(net713),
    .X(net712));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(\core.param_a[10] ));
 sg13g2_buf_2 fanout714 (.A(net716),
    .X(net714));
 sg13g2_buf_1 fanout715 (.A(net716),
    .X(net715));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(net778));
 sg13g2_buf_2 fanout717 (.A(net718),
    .X(net717));
 sg13g2_buf_4 fanout718 (.X(net718),
    .A(\core.param_a[8] ));
 sg13g2_buf_2 fanout719 (.A(net720),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(net723),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(net722),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(net723),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_2720_),
    .X(net723));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(net726));
 sg13g2_buf_2 fanout725 (.A(net726),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_2720_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(net729),
    .X(net727));
 sg13g2_buf_1 fanout728 (.A(net729),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(net730),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(net738),
    .X(net730));
 sg13g2_buf_4 fanout731 (.X(net731),
    .A(net738));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(net738));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(net737));
 sg13g2_buf_2 fanout734 (.A(net737),
    .X(net734));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(net737));
 sg13g2_buf_2 fanout736 (.A(net737),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(net738),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_2720_),
    .X(net738));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(ui_in[2]));
 sg13g2_buf_2 fanout740 (.A(ui_in[2]),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(net1),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(net743),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(net748),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(net748),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(net748),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(net747),
    .X(net746));
 sg13g2_buf_1 fanout747 (.A(net748),
    .X(net747));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(rst_n));
 sg13g2_buf_4 fanout749 (.X(net749),
    .A(net750));
 sg13g2_buf_4 fanout750 (.X(net750),
    .A(net756));
 sg13g2_buf_4 fanout751 (.X(net751),
    .A(net755));
 sg13g2_buf_2 fanout752 (.A(net755),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(net755),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(net755),
    .X(net754));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(net756));
 sg13g2_buf_2 fanout756 (.A(rst_n),
    .X(net756));
 sg13g2_buf_2 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[0]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[1]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[2]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[3]),
    .X(net7));
 sg13g2_tielo tt_um_dpi_adexp_8 (.L_LO(net8));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload1 (.A(clknet_leaf_34_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_36_clk));
 sg13g2_inv_4 clkload3 (.A(clknet_leaf_38_clk));
 sg13g2_inv_2 clkload4 (.A(clknet_leaf_2_clk));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_29_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_30_clk));
 sg13g2_inv_8 clkload7 (.A(clknet_leaf_31_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_28_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_4_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_5_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_2857_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0173_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold3 (.A(_2856_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0254_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0055_),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0379_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold7 (.A(\core.params[5][7] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold8 (.A(_1927_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0051_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0386_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0138_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold12 (.A(_2858_),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0165_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold14 (.A(\core.params[2][4] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold15 (.A(_1941_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold16 (.A(\core.params[6][7] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0121_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold18 (.A(\core.params[7][1] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold19 (.A(_2852_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold20 (.A(\core.params[5][4] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold21 (.A(_1925_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold22 (.A(\core.vm8_reg[6] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0200_),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold24 (.A(\core.params[7][5] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold25 (.A(_2855_),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold26 (.A(\core.params[7][2] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold27 (.A(_2853_),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold28 (.A(\core.params[3][4] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold29 (.A(_1934_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold30 (.A(\core.params[2][5] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold31 (.A(_1942_),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold32 (.A(\core.params[0][4] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold33 (.A(_2813_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold34 (.A(\core.params[7][0] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold35 (.A(_2851_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold36 (.A(\core.params[7][4] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold37 (.A(_2854_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold38 (.A(\core.params[1][3] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold39 (.A(_1948_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold40 (.A(\core.params[0][0] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold41 (.A(_2810_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold42 (.A(\core.params[5][0] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold43 (.A(_1924_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold44 (.A(\core.params[1][0] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold45 (.A(_1946_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold46 (.A(\core.params[3][6] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold47 (.A(_1935_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold48 (.A(\core.params[3][2] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold49 (.A(_1933_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold50 (.A(\core.capacitance[8] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold51 (.A(\core.params[2][3] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0101_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold53 (.A(\core.params[3][1] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold54 (.A(_1932_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold55 (.A(\core.tau_w[8] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold56 (.A(\core.params[3][0] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold57 (.A(_1931_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold58 (.A(\core.params[7][3] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0109_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold60 (.A(\core.params[1][1] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold61 (.A(_1947_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold62 (.A(\core.params[0][3] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold63 (.A(_2812_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold64 (.A(\core.params[0][2] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold65 (.A(_2811_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold66 (.A(\core.params[5][6] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0294_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold68 (.A(\core.params[5][2] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0290_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold70 (.A(\core.params[1][4] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold71 (.A(_1949_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold72 (.A(\core.params[5][5] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold73 (.A(_1926_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold74 (.A(\core.params[5][1] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0289_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold76 (.A(\core.w8_reg[5] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0193_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold78 (.A(\core.params[6][6] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0339_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold80 (.A(\core.params[0][5] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold81 (.A(_2814_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold82 (.A(\core.tau_w[10] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0076_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold84 (.A(\core.watchdog_cnt[11] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0134_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold86 (.A(\core.params[6][4] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0337_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold88 (.A(\core.tau_w[9] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold89 (.A(_2817_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold90 (.A(\core.V_threshold[12] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold91 (.A(\core.params[2][6] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold92 (.A(_1943_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold93 (.A(\core.params[2][1] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0305_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold95 (.A(\core.delta_t[11] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold96 (.A(\core.V_threshold[13] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold97 (.A(\core.vm8_reg[7] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold98 (.A(\core.params[1][2] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0314_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold100 (.A(\core.compute_state[2] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold101 (.A(_2742_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold102 (.A(\core.params[7][7] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0113_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold104 (.A(\core.ibias[14] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold105 (.A(\core.params[2][7] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0311_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold107 (.A(\core.params[3][5] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0301_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold109 (.A(\core.params[0][6] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold110 (.A(_2815_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold111 (.A(\core.w8_reg[6] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold112 (.A(\core.capacitance[9] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold113 (.A(\core.V_threshold[8] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold114 (.A(\core.params[6][0] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0114_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold116 (.A(\core.param_a[13] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold117 (.A(_2845_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold118 (.A(\core.param_b[8] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold119 (.A(\core.temp_q[4] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold120 (.A(\core.capacitance[13] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold121 (.A(\core.temp_q[6] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold122 (.A(\core.params[0][7] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0073_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold124 (.A(\core.param_a[14] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold125 (.A(\core.param_b[9] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold126 (.A(\core.capacitance[10] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold127 (.A(\core.delta_t[10] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold128 (.A(\core.params[3][7] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0303_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold130 (.A(\core.params[6][5] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0338_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold132 (.A(\core.w8_reg[2] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold133 (.A(\core.temp_q[5] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold134 (.A(\core.param_b[10] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold135 (.A(\core.params[7][6] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0112_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold137 (.A(\core.params[1][5] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0317_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold139 (.A(\core.params[0][1] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0067_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold141 (.A(\core.params[3][3] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0299_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold143 (.A(\core.tau_w[11] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold144 (.A(\core.tau_w[12] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold145 (.A(\core.delta_t[13] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold146 (.A(\core.byte_acc[3] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold147 (.A(\core.capacitance[11] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold148 (.A(\core.exp_term[15] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold149 (.A(\core.delta_t[14] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold150 (.A(\core.temp_q[8] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold151 (.A(\core.params[1][6] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0318_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold153 (.A(\core.dV[6] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold154 (.A(_1578_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold155 (.A(\core.watchdog_cnt[4] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0358_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold157 (.A(\core.param_b[12] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold158 (.A(\core.param_b[15] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold159 (.A(\core.temp_q[7] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold160 (.A(\core.spike_reg ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold161 (.A(_1819_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold162 (.A(\core.params[2][2] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0100_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold164 (.A(\core.temp_q[0] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0174_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold166 (.A(\core.params[6][3] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold167 (.A(\core.params[5][3] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold168 (.A(\core.params[1][7] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0319_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold170 (.A(\core.dw[15] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold171 (.A(_1491_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold172 (.A(\core.watchdog_cnt[7] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0366_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold174 (.A(\core.w8_reg[4] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold175 (.A(\core.watchdog_cnt[10] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0374_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold177 (.A(\core.dw[6] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold178 (.A(\core.capacitance[12] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold179 (.A(\core.drive_current[15] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold180 (.A(\core.drive_current[13] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0049_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0367_),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0368_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold184 (.A(\core.w8_reg[3] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold185 (.A(\core.drive_current[10] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold186 (.A(\core.ibias[13] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold187 (.A(\core.drive_current[4] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold188 (.A(\core.V[13] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold189 (.A(\core.capacitance[14] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold190 (.A(\core.delta_t[12] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold191 (.A(\core.drive_current[8] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold192 (.A(\core.params[2][0] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0098_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold194 (.A(\core.dw[12] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold195 (.A(_1488_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold196 (.A(\core.exp_term[12] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold197 (.A(\core.params[6][1] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0115_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold199 (.A(\core.params[6][2] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0116_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold201 (.A(\core.dV[0] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold202 (.A(_1533_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold203 (.A(\core.vm8_reg[3] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold204 (.A(\core.dV[15] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold205 (.A(_1597_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold206 (.A(\core.exp_term[9] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold207 (.A(\core.dV[1] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold208 (.A(_1549_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold209 (.A(\core.vm8_reg[4] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold210 (.A(\core.tau_w[15] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold211 (.A(\core.dV[2] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold212 (.A(_1562_),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold213 (.A(\core.byte_acc[0] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold214 (.A(\core.exp_term[13] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold215 (.A(\core.dV[3] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold216 (.A(_1568_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold217 (.A(\core.param_b[14] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold218 (.A(\core.dw[3] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold219 (.A(\core.dV[5] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold220 (.A(_1575_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold221 (.A(\core.ibias[12] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold222 (.A(\core.vm8_reg[5] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold223 (.A(\core.exp_term[7] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold224 (.A(\core.drive_current[12] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0243_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold226 (.A(\core.temp_q[3] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0662_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold228 (.A(\core.watchdog_cnt[2] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0352_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold230 (.A(\core.dV[7] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold231 (.A(_1582_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold232 (.A(\core.temp_q[11] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold233 (.A(\core.vm8_reg[2] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold234 (.A(\core.dw[5] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold235 (.A(\core.temp_q[2] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0651_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold237 (.A(\core.dV[4] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold238 (.A(_1572_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold239 (.A(\core.param_b[13] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold240 (.A(\core.exp_term[14] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold241 (.A(\core.dw[0] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0048_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0363_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold244 (.A(\core.dw[10] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold245 (.A(\core.tau_w[14] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold246 (.A(\core.drive_current[5] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0236_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold248 (.A(\core.temp_q[12] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold249 (.A(\core.drive_current[14] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold250 (.A(\core.dV[14] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold251 (.A(_1596_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold252 (.A(\core.drive_current[7] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0238_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold254 (.A(\core.temp_q[1] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold255 (.A(\core.drive_current[9] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0240_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold257 (.A(\core.exp_term[10] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold258 (.A(\core.drive_current[6] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0237_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold260 (.A(\core.exp_term[11] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold261 (.A(\core.dw[7] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold262 (.A(\core.dw[14] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold263 (.A(_1490_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold264 (.A(\core.dw[2] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold265 (.A(\core.watchdog_cnt[3] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0356_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold267 (.A(\core.temp_q[9] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold268 (.A(\core.w8_reg[7] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold269 (.A(\core.exp_term[8] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0057_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold271 (.A(_2784_),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0059_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold273 (.A(\core.V_threshold[10] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold274 (.A(\core.temp_q[13] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold275 (.A(\core.drive_current[3] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold276 (.A(\core.drive_current[11] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold277 (.A(\core.capacitance[15] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold278 (.A(\core.dV[10] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold279 (.A(_1590_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold280 (.A(\core.exp_term[1] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold281 (.A(\core.exp_term[4] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold282 (.A(\core.param_a[9] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0099_),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold284 (.A(\core.dw[1] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold285 (.A(\core.V_threshold[9] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold286 (.A(\core.dw[4] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold287 (.A(\core.temp_q[14] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0056_),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold289 (.A(_2794_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0060_),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold291 (.A(\core.exp_term[6] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold292 (.A(\core.watchdog_cnt[5] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold293 (.A(\core.dw[13] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold294 (.A(_1489_),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold295 (.A(\core.compute_state[6] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold296 (.A(\core.exp_term[3] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold297 (.A(\core.dw[8] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold298 (.A(\core.exp_term[2] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold299 (.A(\core.param_b[11] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold300 (.A(\core.dV[12] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold301 (.A(_1594_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold302 (.A(\core.byte_acc[2] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold303 (.A(\core.watchdog_cnt[9] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0372_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold305 (.A(\core.dV[8] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold306 (.A(_1586_),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold307 (.A(\core.dw[11] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold308 (.A(_1487_),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold309 (.A(\core.exp_term[5] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold310 (.A(\core.V_threshold[14] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold311 (.A(\core.delta_t[9] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold312 (.A(\core.ibias[8] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold313 (.A(\core.tau_w[13] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0079_),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold315 (.A(\core.temp_q[10] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold316 (.A(\core.watchdog_cnt[1] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0350_),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0124_),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold319 (.A(\core.leak_current[6] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold320 (.A(\core.V_threshold[11] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold321 (.A(\core.dV[13] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold322 (.A(_1595_),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold323 (.A(\core.leak_current[3] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold324 (.A(\core.leak_current[9] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold325 (.A(\core.leak_current[8] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold326 (.A(\core.temp_q[15] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold327 (.A(\core.leak_current[15] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold328 (.A(\core.ibias[10] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold329 (.A(\core.leak_current[12] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold330 (.A(\core.ibias[11] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold331 (.A(\core.byte_acc[7] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold332 (.A(_2805_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold333 (.A(\core.leak_current[1] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold334 (.A(\core.leak_current[11] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold335 (.A(\core.leak_current[4] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold336 (.A(\core.dV[11] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold337 (.A(_1593_),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold338 (.A(\core.leak_current[10] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold339 (.A(\core.leak_current[7] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold340 (.A(\core.dw[9] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold341 (.A(\core.dV[9] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold342 (.A(_1588_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold343 (.A(\core.leak_current[5] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold344 (.A(\core.leak_current[13] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0510_),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold346 (.A(\core.leak_current[2] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold347 (.A(\core.leak_current[14] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold348 (.A(\core.ibias[9] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold349 (.A(\core.V[2] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold350 (.A(\core.V[6] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold351 (.A(\core.param_idx[0] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0136_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold353 (.A(\core.V[3] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold354 (.A(\core.compute_state[3] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold355 (.A(\core.V[5] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold356 (.A(\core.compute_state[5] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0054_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold358 (.A(_2768_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold359 (.A(_2769_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0058_),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold361 (.A(\core.compute_state[1] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold362 (.A(\core.V[7] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold363 (.A(\core.V[15] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold364 (.A(\core.watchdog_cnt[0] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold365 (.A(\core.compute_state[4] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold366 (.A(\core.V[14] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold367 (.A(\core.byte_acc[6] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold368 (.A(_2803_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold369 (.A(\core.nibble_cnt ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold370 (.A(_2795_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold371 (.A(_2801_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold372 (.A(\core.V[4] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold373 (.A(\core.byte_acc[4] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold374 (.A(\core.V[1] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold375 (.A(\core.w[15] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold376 (.A(\core.V[12] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold377 (.A(\core.w[14] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold378 (.A(\core.byte_acc[1] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold379 (.A(\core.w[6] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold380 (.A(\core.lstate[0] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold381 (.A(\core.w[12] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold382 (.A(\core.w[1] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold383 (.A(\core.param_idx[2] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold384 (.A(\core.V[11] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold385 (.A(\core.w[7] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold386 (.A(\core.w[2] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold387 (.A(\core.w[0] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0256_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold389 (.A(\core.w[4] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold390 (.A(\core.w[13] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold391 (.A(\core.w[11] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold392 (.A(\core.w[3] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold393 (.A(\core.V[10] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold394 (.A(\core.w[5] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold395 (.A(\core.w[10] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold396 (.A(\core.watchdog_cnt[1] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold397 (.A(\core.compute_state[6] ),
    .X(net893));
 sg13g2_antennanp ANTENNA_1 (.A(_0125_));
 sg13g2_antennanp ANTENNA_2 (.A(_0125_));
 sg13g2_antennanp ANTENNA_3 (.A(_0125_));
 sg13g2_antennanp ANTENNA_4 (.A(_0128_));
 sg13g2_antennanp ANTENNA_5 (.A(_0131_));
 sg13g2_antennanp ANTENNA_6 (.A(_0133_));
 sg13g2_antennanp ANTENNA_7 (.A(_0142_));
 sg13g2_antennanp ANTENNA_8 (.A(clk));
 sg13g2_antennanp ANTENNA_9 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_10 (.A(_0060_));
 sg13g2_antennanp ANTENNA_11 (.A(_0062_));
 sg13g2_antennanp ANTENNA_12 (.A(_0063_));
 sg13g2_antennanp ANTENNA_13 (.A(_0063_));
 sg13g2_antennanp ANTENNA_14 (.A(_0064_));
 sg13g2_antennanp ANTENNA_15 (.A(_0128_));
 sg13g2_antennanp ANTENNA_16 (.A(_0131_));
 sg13g2_antennanp ANTENNA_17 (.A(_0133_));
 sg13g2_antennanp ANTENNA_18 (.A(_0142_));
 sg13g2_antennanp ANTENNA_19 (.A(_0372_));
 sg13g2_antennanp ANTENNA_20 (.A(_2769_));
 sg13g2_antennanp ANTENNA_21 (.A(clk));
 sg13g2_antennanp ANTENNA_22 (.A(uio_in[1]));
 sg13g2_antennanp ANTENNA_23 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_24 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_25 (.A(_0060_));
 sg13g2_antennanp ANTENNA_26 (.A(_0128_));
 sg13g2_antennanp ANTENNA_27 (.A(_0128_));
 sg13g2_antennanp ANTENNA_28 (.A(_0131_));
 sg13g2_antennanp ANTENNA_29 (.A(_0142_));
 sg13g2_antennanp ANTENNA_30 (.A(clk));
 sg13g2_antennanp ANTENNA_31 (.A(ui_in[3]));
 sg13g2_antennanp ANTENNA_32 (.A(uio_in[1]));
 sg13g2_antennanp ANTENNA_33 (.A(uio_in[2]));
 sg13g2_antennanp ANTENNA_34 (.A(uio_in[3]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_67 ();
 sg13g2_decap_8 FILLER_0_78 ();
 sg13g2_decap_4 FILLER_0_85 ();
 sg13g2_decap_4 FILLER_0_97 ();
 sg13g2_fill_2 FILLER_0_101 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_fill_2 FILLER_0_119 ();
 sg13g2_fill_2 FILLER_0_130 ();
 sg13g2_fill_1 FILLER_0_132 ();
 sg13g2_fill_2 FILLER_0_137 ();
 sg13g2_decap_8 FILLER_0_144 ();
 sg13g2_fill_2 FILLER_0_151 ();
 sg13g2_fill_1 FILLER_0_153 ();
 sg13g2_fill_2 FILLER_0_159 ();
 sg13g2_fill_1 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_167 ();
 sg13g2_decap_8 FILLER_0_174 ();
 sg13g2_fill_1 FILLER_0_181 ();
 sg13g2_decap_4 FILLER_0_186 ();
 sg13g2_fill_1 FILLER_0_190 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_fill_2 FILLER_0_212 ();
 sg13g2_decap_8 FILLER_0_218 ();
 sg13g2_decap_4 FILLER_0_225 ();
 sg13g2_fill_2 FILLER_0_229 ();
 sg13g2_fill_1 FILLER_0_236 ();
 sg13g2_decap_8 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_4 FILLER_0_268 ();
 sg13g2_fill_1 FILLER_0_272 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_4 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_293 ();
 sg13g2_decap_4 FILLER_0_300 ();
 sg13g2_fill_1 FILLER_0_304 ();
 sg13g2_decap_4 FILLER_0_308 ();
 sg13g2_fill_1 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_4 FILLER_0_344 ();
 sg13g2_fill_2 FILLER_0_348 ();
 sg13g2_fill_2 FILLER_0_355 ();
 sg13g2_fill_1 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_4 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_4 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_46 ();
 sg13g2_fill_1 FILLER_1_103 ();
 sg13g2_fill_2 FILLER_1_138 ();
 sg13g2_decap_4 FILLER_1_155 ();
 sg13g2_decap_4 FILLER_1_167 ();
 sg13g2_fill_1 FILLER_1_202 ();
 sg13g2_fill_2 FILLER_1_234 ();
 sg13g2_decap_8 FILLER_1_257 ();
 sg13g2_fill_2 FILLER_1_277 ();
 sg13g2_fill_1 FILLER_1_279 ();
 sg13g2_fill_2 FILLER_1_374 ();
 sg13g2_fill_1 FILLER_1_376 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_fill_2 FILLER_2_35 ();
 sg13g2_fill_2 FILLER_2_93 ();
 sg13g2_fill_2 FILLER_2_140 ();
 sg13g2_fill_1 FILLER_2_179 ();
 sg13g2_fill_1 FILLER_2_225 ();
 sg13g2_fill_1 FILLER_2_247 ();
 sg13g2_fill_2 FILLER_2_256 ();
 sg13g2_decap_4 FILLER_2_319 ();
 sg13g2_fill_2 FILLER_2_371 ();
 sg13g2_fill_1 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_4 FILLER_3_28 ();
 sg13g2_fill_2 FILLER_3_104 ();
 sg13g2_fill_2 FILLER_3_119 ();
 sg13g2_fill_1 FILLER_3_187 ();
 sg13g2_fill_1 FILLER_3_229 ();
 sg13g2_fill_1 FILLER_3_242 ();
 sg13g2_fill_2 FILLER_3_255 ();
 sg13g2_fill_1 FILLER_3_257 ();
 sg13g2_fill_1 FILLER_3_296 ();
 sg13g2_fill_2 FILLER_3_321 ();
 sg13g2_fill_1 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_fill_1 FILLER_4_35 ();
 sg13g2_fill_1 FILLER_4_56 ();
 sg13g2_fill_1 FILLER_4_67 ();
 sg13g2_fill_1 FILLER_4_86 ();
 sg13g2_fill_1 FILLER_4_135 ();
 sg13g2_fill_2 FILLER_4_181 ();
 sg13g2_fill_1 FILLER_4_188 ();
 sg13g2_fill_1 FILLER_4_207 ();
 sg13g2_decap_8 FILLER_4_212 ();
 sg13g2_decap_4 FILLER_4_248 ();
 sg13g2_fill_1 FILLER_4_252 ();
 sg13g2_decap_4 FILLER_4_266 ();
 sg13g2_fill_2 FILLER_4_270 ();
 sg13g2_fill_2 FILLER_4_277 ();
 sg13g2_fill_2 FILLER_4_312 ();
 sg13g2_fill_2 FILLER_4_333 ();
 sg13g2_fill_1 FILLER_4_335 ();
 sg13g2_decap_8 FILLER_4_348 ();
 sg13g2_fill_1 FILLER_4_355 ();
 sg13g2_fill_1 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_4 FILLER_5_35 ();
 sg13g2_fill_1 FILLER_5_39 ();
 sg13g2_fill_2 FILLER_5_45 ();
 sg13g2_fill_2 FILLER_5_76 ();
 sg13g2_fill_2 FILLER_5_83 ();
 sg13g2_fill_1 FILLER_5_85 ();
 sg13g2_fill_2 FILLER_5_104 ();
 sg13g2_fill_1 FILLER_5_106 ();
 sg13g2_fill_1 FILLER_5_121 ();
 sg13g2_fill_2 FILLER_5_145 ();
 sg13g2_fill_1 FILLER_5_164 ();
 sg13g2_fill_2 FILLER_5_182 ();
 sg13g2_fill_1 FILLER_5_184 ();
 sg13g2_decap_8 FILLER_5_195 ();
 sg13g2_decap_8 FILLER_5_202 ();
 sg13g2_decap_8 FILLER_5_209 ();
 sg13g2_fill_1 FILLER_5_216 ();
 sg13g2_fill_2 FILLER_5_231 ();
 sg13g2_fill_2 FILLER_5_237 ();
 sg13g2_fill_1 FILLER_5_249 ();
 sg13g2_fill_1 FILLER_5_257 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_fill_2 FILLER_5_281 ();
 sg13g2_fill_1 FILLER_5_283 ();
 sg13g2_fill_2 FILLER_5_288 ();
 sg13g2_fill_2 FILLER_5_302 ();
 sg13g2_fill_1 FILLER_5_304 ();
 sg13g2_fill_2 FILLER_5_322 ();
 sg13g2_fill_1 FILLER_5_324 ();
 sg13g2_fill_2 FILLER_5_330 ();
 sg13g2_fill_1 FILLER_5_332 ();
 sg13g2_decap_4 FILLER_5_346 ();
 sg13g2_fill_1 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_4 FILLER_6_7 ();
 sg13g2_fill_2 FILLER_6_15 ();
 sg13g2_fill_2 FILLER_6_34 ();
 sg13g2_fill_2 FILLER_6_199 ();
 sg13g2_fill_1 FILLER_6_201 ();
 sg13g2_decap_8 FILLER_6_206 ();
 sg13g2_fill_1 FILLER_6_213 ();
 sg13g2_fill_1 FILLER_6_233 ();
 sg13g2_fill_2 FILLER_6_251 ();
 sg13g2_fill_1 FILLER_6_270 ();
 sg13g2_fill_2 FILLER_6_284 ();
 sg13g2_fill_2 FILLER_6_307 ();
 sg13g2_fill_1 FILLER_6_342 ();
 sg13g2_decap_4 FILLER_6_355 ();
 sg13g2_decap_8 FILLER_6_367 ();
 sg13g2_fill_1 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_20 ();
 sg13g2_fill_2 FILLER_7_59 ();
 sg13g2_fill_2 FILLER_7_102 ();
 sg13g2_fill_2 FILLER_7_113 ();
 sg13g2_decap_8 FILLER_7_214 ();
 sg13g2_fill_1 FILLER_7_221 ();
 sg13g2_fill_1 FILLER_7_244 ();
 sg13g2_fill_1 FILLER_7_267 ();
 sg13g2_fill_2 FILLER_7_289 ();
 sg13g2_fill_1 FILLER_7_291 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_fill_2 FILLER_7_332 ();
 sg13g2_fill_1 FILLER_7_334 ();
 sg13g2_decap_8 FILLER_7_340 ();
 sg13g2_decap_4 FILLER_7_347 ();
 sg13g2_fill_1 FILLER_7_351 ();
 sg13g2_decap_4 FILLER_7_360 ();
 sg13g2_fill_2 FILLER_7_364 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_2 FILLER_8_45 ();
 sg13g2_fill_2 FILLER_8_56 ();
 sg13g2_decap_4 FILLER_8_66 ();
 sg13g2_fill_1 FILLER_8_70 ();
 sg13g2_fill_2 FILLER_8_84 ();
 sg13g2_fill_1 FILLER_8_86 ();
 sg13g2_fill_1 FILLER_8_91 ();
 sg13g2_fill_2 FILLER_8_118 ();
 sg13g2_fill_1 FILLER_8_120 ();
 sg13g2_fill_2 FILLER_8_136 ();
 sg13g2_fill_1 FILLER_8_173 ();
 sg13g2_fill_2 FILLER_8_187 ();
 sg13g2_fill_2 FILLER_8_225 ();
 sg13g2_fill_2 FILLER_8_237 ();
 sg13g2_fill_1 FILLER_8_239 ();
 sg13g2_fill_1 FILLER_8_274 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_fill_2 FILLER_8_315 ();
 sg13g2_fill_1 FILLER_8_317 ();
 sg13g2_decap_8 FILLER_8_327 ();
 sg13g2_decap_4 FILLER_8_334 ();
 sg13g2_fill_2 FILLER_8_338 ();
 sg13g2_fill_1 FILLER_8_345 ();
 sg13g2_fill_1 FILLER_8_353 ();
 sg13g2_fill_2 FILLER_8_375 ();
 sg13g2_fill_1 FILLER_8_377 ();
 sg13g2_fill_1 FILLER_8_391 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_decap_4 FILLER_9_55 ();
 sg13g2_fill_1 FILLER_9_59 ();
 sg13g2_fill_2 FILLER_9_79 ();
 sg13g2_decap_4 FILLER_9_86 ();
 sg13g2_fill_1 FILLER_9_90 ();
 sg13g2_fill_2 FILLER_9_104 ();
 sg13g2_fill_1 FILLER_9_114 ();
 sg13g2_fill_1 FILLER_9_217 ();
 sg13g2_fill_1 FILLER_9_226 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_4 FILLER_9_252 ();
 sg13g2_fill_1 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_267 ();
 sg13g2_decap_8 FILLER_9_274 ();
 sg13g2_decap_4 FILLER_9_281 ();
 sg13g2_fill_1 FILLER_9_285 ();
 sg13g2_fill_1 FILLER_9_291 ();
 sg13g2_fill_2 FILLER_9_296 ();
 sg13g2_fill_1 FILLER_9_321 ();
 sg13g2_fill_1 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_fill_2 FILLER_9_388 ();
 sg13g2_fill_1 FILLER_9_390 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_fill_2 FILLER_10_11 ();
 sg13g2_fill_1 FILLER_10_13 ();
 sg13g2_decap_8 FILLER_10_30 ();
 sg13g2_decap_8 FILLER_10_37 ();
 sg13g2_decap_8 FILLER_10_44 ();
 sg13g2_fill_1 FILLER_10_51 ();
 sg13g2_fill_1 FILLER_10_97 ();
 sg13g2_fill_2 FILLER_10_123 ();
 sg13g2_fill_1 FILLER_10_125 ();
 sg13g2_fill_2 FILLER_10_136 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_fill_2 FILLER_10_203 ();
 sg13g2_fill_1 FILLER_10_205 ();
 sg13g2_decap_8 FILLER_10_215 ();
 sg13g2_fill_2 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_246 ();
 sg13g2_fill_2 FILLER_10_253 ();
 sg13g2_fill_1 FILLER_10_255 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_4 FILLER_10_289 ();
 sg13g2_fill_2 FILLER_10_293 ();
 sg13g2_fill_1 FILLER_10_307 ();
 sg13g2_fill_2 FILLER_10_314 ();
 sg13g2_fill_1 FILLER_10_347 ();
 sg13g2_fill_2 FILLER_10_355 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_14 ();
 sg13g2_fill_1 FILLER_11_29 ();
 sg13g2_fill_2 FILLER_11_38 ();
 sg13g2_fill_1 FILLER_11_40 ();
 sg13g2_fill_2 FILLER_11_45 ();
 sg13g2_fill_1 FILLER_11_47 ();
 sg13g2_fill_2 FILLER_11_80 ();
 sg13g2_decap_4 FILLER_11_86 ();
 sg13g2_fill_2 FILLER_11_90 ();
 sg13g2_fill_1 FILLER_11_118 ();
 sg13g2_fill_2 FILLER_11_148 ();
 sg13g2_decap_8 FILLER_11_155 ();
 sg13g2_fill_1 FILLER_11_162 ();
 sg13g2_fill_2 FILLER_11_193 ();
 sg13g2_fill_1 FILLER_11_200 ();
 sg13g2_fill_2 FILLER_11_206 ();
 sg13g2_fill_1 FILLER_11_208 ();
 sg13g2_fill_1 FILLER_11_218 ();
 sg13g2_fill_2 FILLER_11_232 ();
 sg13g2_fill_1 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_260 ();
 sg13g2_fill_2 FILLER_11_291 ();
 sg13g2_fill_1 FILLER_11_310 ();
 sg13g2_fill_1 FILLER_11_319 ();
 sg13g2_fill_1 FILLER_11_353 ();
 sg13g2_fill_1 FILLER_11_358 ();
 sg13g2_fill_2 FILLER_11_379 ();
 sg13g2_fill_1 FILLER_11_381 ();
 sg13g2_fill_2 FILLER_11_395 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_23 ();
 sg13g2_fill_2 FILLER_12_33 ();
 sg13g2_fill_1 FILLER_12_35 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_fill_1 FILLER_12_62 ();
 sg13g2_fill_1 FILLER_12_68 ();
 sg13g2_decap_4 FILLER_12_74 ();
 sg13g2_fill_1 FILLER_12_86 ();
 sg13g2_decap_8 FILLER_12_153 ();
 sg13g2_decap_8 FILLER_12_160 ();
 sg13g2_fill_1 FILLER_12_170 ();
 sg13g2_fill_1 FILLER_12_197 ();
 sg13g2_decap_4 FILLER_12_224 ();
 sg13g2_fill_2 FILLER_12_250 ();
 sg13g2_fill_1 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_fill_2 FILLER_12_317 ();
 sg13g2_decap_8 FILLER_12_327 ();
 sg13g2_decap_4 FILLER_12_334 ();
 sg13g2_decap_4 FILLER_12_343 ();
 sg13g2_fill_2 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_fill_2 FILLER_12_359 ();
 sg13g2_fill_1 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_fill_2 FILLER_12_373 ();
 sg13g2_fill_1 FILLER_12_380 ();
 sg13g2_decap_4 FILLER_12_385 ();
 sg13g2_fill_1 FILLER_12_389 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_4 ();
 sg13g2_fill_2 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_16 ();
 sg13g2_fill_2 FILLER_13_26 ();
 sg13g2_fill_1 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_38 ();
 sg13g2_decap_8 FILLER_13_45 ();
 sg13g2_decap_4 FILLER_13_52 ();
 sg13g2_fill_1 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_106 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_fill_1 FILLER_13_165 ();
 sg13g2_fill_1 FILLER_13_170 ();
 sg13g2_fill_1 FILLER_13_181 ();
 sg13g2_fill_2 FILLER_13_187 ();
 sg13g2_fill_2 FILLER_13_215 ();
 sg13g2_fill_1 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_268 ();
 sg13g2_fill_1 FILLER_13_275 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_fill_2 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_318 ();
 sg13g2_fill_1 FILLER_13_325 ();
 sg13g2_decap_8 FILLER_13_342 ();
 sg13g2_fill_1 FILLER_13_349 ();
 sg13g2_decap_4 FILLER_13_389 ();
 sg13g2_fill_1 FILLER_13_393 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_19 ();
 sg13g2_fill_1 FILLER_14_33 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_4 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_53 ();
 sg13g2_decap_8 FILLER_14_75 ();
 sg13g2_fill_2 FILLER_14_82 ();
 sg13g2_fill_2 FILLER_14_199 ();
 sg13g2_fill_1 FILLER_14_201 ();
 sg13g2_decap_4 FILLER_14_222 ();
 sg13g2_fill_2 FILLER_14_226 ();
 sg13g2_decap_4 FILLER_14_236 ();
 sg13g2_fill_2 FILLER_14_240 ();
 sg13g2_decap_8 FILLER_14_246 ();
 sg13g2_decap_4 FILLER_14_253 ();
 sg13g2_fill_1 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_274 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_1 FILLER_14_315 ();
 sg13g2_fill_1 FILLER_14_324 ();
 sg13g2_fill_1 FILLER_14_333 ();
 sg13g2_fill_2 FILLER_14_346 ();
 sg13g2_fill_1 FILLER_14_360 ();
 sg13g2_fill_2 FILLER_14_376 ();
 sg13g2_fill_1 FILLER_14_378 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_27 ();
 sg13g2_fill_2 FILLER_15_53 ();
 sg13g2_fill_1 FILLER_15_55 ();
 sg13g2_fill_2 FILLER_15_64 ();
 sg13g2_fill_1 FILLER_15_66 ();
 sg13g2_decap_8 FILLER_15_79 ();
 sg13g2_fill_2 FILLER_15_86 ();
 sg13g2_fill_1 FILLER_15_88 ();
 sg13g2_fill_2 FILLER_15_115 ();
 sg13g2_fill_1 FILLER_15_135 ();
 sg13g2_fill_2 FILLER_15_168 ();
 sg13g2_decap_4 FILLER_15_175 ();
 sg13g2_fill_2 FILLER_15_215 ();
 sg13g2_decap_4 FILLER_15_229 ();
 sg13g2_decap_8 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_250 ();
 sg13g2_fill_1 FILLER_15_260 ();
 sg13g2_decap_4 FILLER_15_282 ();
 sg13g2_fill_2 FILLER_15_345 ();
 sg13g2_fill_2 FILLER_15_365 ();
 sg13g2_decap_4 FILLER_15_380 ();
 sg13g2_fill_1 FILLER_15_384 ();
 sg13g2_fill_2 FILLER_15_390 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_4 ();
 sg13g2_fill_2 FILLER_16_25 ();
 sg13g2_fill_1 FILLER_16_68 ();
 sg13g2_fill_1 FILLER_16_74 ();
 sg13g2_decap_8 FILLER_16_89 ();
 sg13g2_fill_1 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_201 ();
 sg13g2_fill_1 FILLER_16_203 ();
 sg13g2_fill_1 FILLER_16_230 ();
 sg13g2_fill_2 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_251 ();
 sg13g2_fill_1 FILLER_16_286 ();
 sg13g2_fill_2 FILLER_16_296 ();
 sg13g2_fill_1 FILLER_16_298 ();
 sg13g2_fill_2 FILLER_16_311 ();
 sg13g2_fill_2 FILLER_16_343 ();
 sg13g2_fill_1 FILLER_16_372 ();
 sg13g2_fill_2 FILLER_16_390 ();
 sg13g2_fill_1 FILLER_16_392 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_50 ();
 sg13g2_fill_1 FILLER_17_73 ();
 sg13g2_fill_1 FILLER_17_109 ();
 sg13g2_fill_2 FILLER_17_118 ();
 sg13g2_fill_2 FILLER_17_159 ();
 sg13g2_fill_2 FILLER_17_171 ();
 sg13g2_fill_1 FILLER_17_230 ();
 sg13g2_fill_2 FILLER_17_236 ();
 sg13g2_decap_4 FILLER_17_289 ();
 sg13g2_fill_2 FILLER_17_316 ();
 sg13g2_decap_4 FILLER_17_323 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_decap_4 FILLER_17_338 ();
 sg13g2_fill_2 FILLER_17_378 ();
 sg13g2_fill_1 FILLER_17_380 ();
 sg13g2_fill_1 FILLER_17_404 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_11 ();
 sg13g2_fill_2 FILLER_18_23 ();
 sg13g2_fill_2 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_54 ();
 sg13g2_fill_1 FILLER_18_61 ();
 sg13g2_decap_4 FILLER_18_66 ();
 sg13g2_fill_1 FILLER_18_70 ();
 sg13g2_decap_4 FILLER_18_87 ();
 sg13g2_fill_1 FILLER_18_91 ();
 sg13g2_fill_2 FILLER_18_113 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_2 FILLER_18_128 ();
 sg13g2_fill_1 FILLER_18_130 ();
 sg13g2_fill_2 FILLER_18_145 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_fill_2 FILLER_18_185 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_fill_2 FILLER_18_254 ();
 sg13g2_fill_2 FILLER_18_261 ();
 sg13g2_fill_1 FILLER_18_263 ();
 sg13g2_fill_2 FILLER_18_298 ();
 sg13g2_fill_1 FILLER_18_300 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_decap_4 FILLER_18_314 ();
 sg13g2_fill_2 FILLER_18_318 ();
 sg13g2_decap_4 FILLER_18_350 ();
 sg13g2_fill_2 FILLER_18_354 ();
 sg13g2_decap_4 FILLER_18_366 ();
 sg13g2_fill_2 FILLER_18_370 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_4 FILLER_19_58 ();
 sg13g2_fill_2 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_151 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_fill_2 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_fill_2 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_275 ();
 sg13g2_fill_1 FILLER_19_297 ();
 sg13g2_decap_4 FILLER_19_327 ();
 sg13g2_decap_8 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_365 ();
 sg13g2_fill_2 FILLER_20_31 ();
 sg13g2_decap_8 FILLER_20_37 ();
 sg13g2_decap_4 FILLER_20_59 ();
 sg13g2_fill_2 FILLER_20_75 ();
 sg13g2_fill_1 FILLER_20_77 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_fill_2 FILLER_20_188 ();
 sg13g2_fill_1 FILLER_20_212 ();
 sg13g2_fill_1 FILLER_20_222 ();
 sg13g2_decap_4 FILLER_20_246 ();
 sg13g2_fill_1 FILLER_20_254 ();
 sg13g2_fill_2 FILLER_20_265 ();
 sg13g2_fill_1 FILLER_20_267 ();
 sg13g2_fill_2 FILLER_20_289 ();
 sg13g2_decap_4 FILLER_20_334 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_fill_1 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_387 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_13 ();
 sg13g2_fill_1 FILLER_21_15 ();
 sg13g2_fill_1 FILLER_21_23 ();
 sg13g2_fill_2 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_38 ();
 sg13g2_fill_1 FILLER_21_40 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_fill_2 FILLER_21_73 ();
 sg13g2_fill_2 FILLER_21_106 ();
 sg13g2_fill_2 FILLER_21_129 ();
 sg13g2_fill_2 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_161 ();
 sg13g2_fill_2 FILLER_21_181 ();
 sg13g2_fill_2 FILLER_21_192 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_decap_8 FILLER_21_248 ();
 sg13g2_decap_4 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_296 ();
 sg13g2_fill_2 FILLER_21_330 ();
 sg13g2_decap_4 FILLER_21_358 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_fill_2 FILLER_21_371 ();
 sg13g2_fill_1 FILLER_21_373 ();
 sg13g2_fill_2 FILLER_21_391 ();
 sg13g2_fill_1 FILLER_21_393 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_1 FILLER_22_12 ();
 sg13g2_fill_2 FILLER_22_21 ();
 sg13g2_fill_1 FILLER_22_23 ();
 sg13g2_fill_2 FILLER_22_53 ();
 sg13g2_fill_1 FILLER_22_55 ();
 sg13g2_fill_1 FILLER_22_81 ();
 sg13g2_decap_4 FILLER_22_87 ();
 sg13g2_decap_8 FILLER_22_121 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_fill_1 FILLER_22_162 ();
 sg13g2_fill_1 FILLER_22_193 ();
 sg13g2_fill_1 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_366 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_fill_2 FILLER_22_385 ();
 sg13g2_fill_1 FILLER_22_387 ();
 sg13g2_fill_1 FILLER_22_398 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_18 ();
 sg13g2_fill_1 FILLER_23_20 ();
 sg13g2_fill_1 FILLER_23_38 ();
 sg13g2_fill_1 FILLER_23_43 ();
 sg13g2_fill_2 FILLER_23_60 ();
 sg13g2_decap_4 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_74 ();
 sg13g2_fill_1 FILLER_23_81 ();
 sg13g2_decap_4 FILLER_23_86 ();
 sg13g2_fill_1 FILLER_23_90 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_fill_2 FILLER_23_123 ();
 sg13g2_fill_1 FILLER_23_125 ();
 sg13g2_fill_1 FILLER_23_170 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_246 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_4 FILLER_23_277 ();
 sg13g2_fill_2 FILLER_23_289 ();
 sg13g2_fill_1 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_4 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_319 ();
 sg13g2_fill_1 FILLER_23_348 ();
 sg13g2_fill_2 FILLER_23_388 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_19 ();
 sg13g2_fill_1 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_31 ();
 sg13g2_decap_8 FILLER_24_40 ();
 sg13g2_fill_1 FILLER_24_47 ();
 sg13g2_decap_8 FILLER_24_52 ();
 sg13g2_decap_8 FILLER_24_59 ();
 sg13g2_decap_8 FILLER_24_66 ();
 sg13g2_fill_1 FILLER_24_73 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_100 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_decap_4 FILLER_24_139 ();
 sg13g2_fill_2 FILLER_24_143 ();
 sg13g2_decap_8 FILLER_24_149 ();
 sg13g2_decap_4 FILLER_24_156 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_fill_2 FILLER_24_197 ();
 sg13g2_fill_2 FILLER_24_259 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_fill_2 FILLER_24_281 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_fill_2 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_325 ();
 sg13g2_fill_1 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_25 ();
 sg13g2_fill_2 FILLER_25_43 ();
 sg13g2_fill_1 FILLER_25_45 ();
 sg13g2_decap_8 FILLER_25_50 ();
 sg13g2_fill_2 FILLER_25_57 ();
 sg13g2_fill_2 FILLER_25_76 ();
 sg13g2_fill_1 FILLER_25_83 ();
 sg13g2_decap_4 FILLER_25_89 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_fill_1 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_146 ();
 sg13g2_fill_2 FILLER_25_193 ();
 sg13g2_fill_2 FILLER_25_204 ();
 sg13g2_fill_1 FILLER_25_206 ();
 sg13g2_decap_8 FILLER_25_255 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_decap_8 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_289 ();
 sg13g2_decap_4 FILLER_25_296 ();
 sg13g2_fill_1 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_327 ();
 sg13g2_fill_1 FILLER_25_362 ();
 sg13g2_fill_1 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_4 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_26 ();
 sg13g2_fill_1 FILLER_26_64 ();
 sg13g2_fill_2 FILLER_26_81 ();
 sg13g2_fill_1 FILLER_26_126 ();
 sg13g2_fill_2 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_174 ();
 sg13g2_fill_2 FILLER_26_222 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_fill_1 FILLER_26_328 ();
 sg13g2_fill_2 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_390 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_50 ();
 sg13g2_fill_2 FILLER_27_60 ();
 sg13g2_fill_2 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_80 ();
 sg13g2_fill_2 FILLER_27_107 ();
 sg13g2_fill_1 FILLER_27_109 ();
 sg13g2_fill_2 FILLER_27_123 ();
 sg13g2_fill_2 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_310 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_decap_8 FILLER_27_330 ();
 sg13g2_fill_2 FILLER_27_337 ();
 sg13g2_fill_1 FILLER_27_339 ();
 sg13g2_fill_2 FILLER_27_344 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_28_26 ();
 sg13g2_fill_2 FILLER_28_36 ();
 sg13g2_fill_1 FILLER_28_38 ();
 sg13g2_fill_1 FILLER_28_44 ();
 sg13g2_fill_2 FILLER_28_109 ();
 sg13g2_decap_8 FILLER_28_123 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_193 ();
 sg13g2_fill_1 FILLER_28_209 ();
 sg13g2_decap_4 FILLER_28_235 ();
 sg13g2_fill_2 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_fill_1 FILLER_28_340 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_23 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_4 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_67 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_decap_4 FILLER_29_89 ();
 sg13g2_fill_2 FILLER_29_93 ();
 sg13g2_decap_8 FILLER_29_99 ();
 sg13g2_fill_2 FILLER_29_106 ();
 sg13g2_fill_1 FILLER_29_108 ();
 sg13g2_decap_8 FILLER_29_143 ();
 sg13g2_fill_1 FILLER_29_154 ();
 sg13g2_fill_2 FILLER_29_190 ();
 sg13g2_fill_1 FILLER_29_192 ();
 sg13g2_fill_2 FILLER_29_211 ();
 sg13g2_fill_1 FILLER_29_213 ();
 sg13g2_decap_8 FILLER_29_226 ();
 sg13g2_decap_4 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_237 ();
 sg13g2_decap_4 FILLER_29_243 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_fill_2 FILLER_29_262 ();
 sg13g2_decap_4 FILLER_29_268 ();
 sg13g2_fill_1 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_277 ();
 sg13g2_decap_4 FILLER_29_284 ();
 sg13g2_fill_1 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_310 ();
 sg13g2_fill_2 FILLER_29_319 ();
 sg13g2_fill_2 FILLER_29_356 ();
 sg13g2_fill_1 FILLER_29_394 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_2 FILLER_30_31 ();
 sg13g2_fill_1 FILLER_30_71 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_fill_2 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_124 ();
 sg13g2_decap_4 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_156 ();
 sg13g2_fill_1 FILLER_30_175 ();
 sg13g2_fill_2 FILLER_30_198 ();
 sg13g2_decap_4 FILLER_30_222 ();
 sg13g2_fill_1 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_309 ();
 sg13g2_fill_1 FILLER_30_348 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_19 ();
 sg13g2_fill_1 FILLER_31_29 ();
 sg13g2_fill_1 FILLER_31_54 ();
 sg13g2_decap_8 FILLER_31_75 ();
 sg13g2_decap_4 FILLER_31_86 ();
 sg13g2_fill_1 FILLER_31_90 ();
 sg13g2_fill_2 FILLER_31_96 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_130 ();
 sg13g2_fill_2 FILLER_31_137 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_fill_2 FILLER_31_310 ();
 sg13g2_fill_1 FILLER_31_312 ();
 sg13g2_decap_4 FILLER_31_321 ();
 sg13g2_fill_2 FILLER_31_325 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_351 ();
 sg13g2_fill_2 FILLER_31_385 ();
 sg13g2_fill_2 FILLER_31_391 ();
 sg13g2_fill_1 FILLER_31_393 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_101 ();
 sg13g2_fill_2 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_decap_4 FILLER_32_261 ();
 sg13g2_decap_8 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_320 ();
 sg13g2_decap_8 FILLER_32_342 ();
 sg13g2_decap_4 FILLER_32_349 ();
 sg13g2_decap_4 FILLER_32_362 ();
 sg13g2_fill_1 FILLER_32_370 ();
 sg13g2_fill_2 FILLER_32_375 ();
 sg13g2_fill_1 FILLER_32_377 ();
 sg13g2_fill_1 FILLER_32_404 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_41 ();
 sg13g2_decap_8 FILLER_33_48 ();
 sg13g2_decap_8 FILLER_33_55 ();
 sg13g2_fill_2 FILLER_33_62 ();
 sg13g2_decap_4 FILLER_33_71 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_fill_2 FILLER_33_203 ();
 sg13g2_fill_2 FILLER_33_214 ();
 sg13g2_fill_2 FILLER_33_233 ();
 sg13g2_fill_2 FILLER_33_240 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_decap_4 FILLER_33_248 ();
 sg13g2_decap_8 FILLER_33_281 ();
 sg13g2_decap_8 FILLER_33_288 ();
 sg13g2_fill_2 FILLER_33_329 ();
 sg13g2_fill_1 FILLER_33_331 ();
 sg13g2_fill_2 FILLER_33_373 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_26 ();
 sg13g2_decap_4 FILLER_34_33 ();
 sg13g2_fill_2 FILLER_34_37 ();
 sg13g2_fill_1 FILLER_34_43 ();
 sg13g2_decap_8 FILLER_34_52 ();
 sg13g2_fill_2 FILLER_34_59 ();
 sg13g2_fill_1 FILLER_34_82 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_159 ();
 sg13g2_fill_2 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_243 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_280 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_fill_2 FILLER_34_309 ();
 sg13g2_fill_1 FILLER_34_311 ();
 sg13g2_fill_2 FILLER_34_347 ();
 sg13g2_fill_2 FILLER_34_357 ();
 sg13g2_fill_1 FILLER_34_359 ();
 sg13g2_fill_1 FILLER_34_386 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_2 FILLER_35_24 ();
 sg13g2_fill_1 FILLER_35_34 ();
 sg13g2_fill_2 FILLER_35_64 ();
 sg13g2_fill_1 FILLER_35_66 ();
 sg13g2_fill_2 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_132 ();
 sg13g2_fill_2 FILLER_35_171 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_180 ();
 sg13g2_fill_1 FILLER_35_208 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_decap_4 FILLER_35_254 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_fill_1 FILLER_35_282 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_2 FILLER_36_13 ();
 sg13g2_fill_1 FILLER_36_15 ();
 sg13g2_fill_2 FILLER_36_34 ();
 sg13g2_fill_1 FILLER_36_62 ();
 sg13g2_fill_2 FILLER_36_101 ();
 sg13g2_fill_1 FILLER_36_103 ();
 sg13g2_fill_2 FILLER_36_118 ();
 sg13g2_fill_1 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_183 ();
 sg13g2_fill_2 FILLER_36_200 ();
 sg13g2_fill_1 FILLER_36_202 ();
 sg13g2_fill_2 FILLER_36_209 ();
 sg13g2_fill_1 FILLER_36_211 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_250 ();
 sg13g2_fill_1 FILLER_36_252 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_fill_2 FILLER_36_323 ();
 sg13g2_fill_1 FILLER_36_325 ();
 sg13g2_fill_2 FILLER_36_368 ();
 sg13g2_fill_2 FILLER_36_389 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_1 FILLER_37_13 ();
 sg13g2_decap_4 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_46 ();
 sg13g2_fill_1 FILLER_37_52 ();
 sg13g2_fill_1 FILLER_37_104 ();
 sg13g2_fill_1 FILLER_37_123 ();
 sg13g2_fill_2 FILLER_37_150 ();
 sg13g2_decap_4 FILLER_37_178 ();
 sg13g2_fill_2 FILLER_37_186 ();
 sg13g2_fill_1 FILLER_37_188 ();
 sg13g2_fill_1 FILLER_37_204 ();
 sg13g2_fill_2 FILLER_37_261 ();
 sg13g2_fill_1 FILLER_37_271 ();
 sg13g2_fill_2 FILLER_37_305 ();
 sg13g2_fill_1 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_390 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_9 ();
 sg13g2_decap_4 FILLER_38_26 ();
 sg13g2_fill_1 FILLER_38_30 ();
 sg13g2_fill_2 FILLER_38_41 ();
 sg13g2_decap_4 FILLER_38_51 ();
 sg13g2_fill_1 FILLER_38_63 ();
 sg13g2_decap_4 FILLER_38_82 ();
 sg13g2_fill_1 FILLER_38_86 ();
 sg13g2_fill_1 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_decap_4 FILLER_38_244 ();
 sg13g2_decap_8 FILLER_38_261 ();
 sg13g2_decap_8 FILLER_38_268 ();
 sg13g2_decap_8 FILLER_38_275 ();
 sg13g2_decap_8 FILLER_38_282 ();
 sg13g2_fill_2 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_fill_1 FILLER_38_313 ();
 sg13g2_fill_1 FILLER_38_344 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_7 ();
 sg13g2_fill_1 FILLER_39_9 ();
 sg13g2_decap_4 FILLER_39_26 ();
 sg13g2_fill_2 FILLER_39_52 ();
 sg13g2_fill_1 FILLER_39_54 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_4 FILLER_39_84 ();
 sg13g2_fill_1 FILLER_39_88 ();
 sg13g2_fill_2 FILLER_39_93 ();
 sg13g2_decap_8 FILLER_39_134 ();
 sg13g2_fill_2 FILLER_39_141 ();
 sg13g2_fill_1 FILLER_39_143 ();
 sg13g2_fill_1 FILLER_39_158 ();
 sg13g2_fill_1 FILLER_39_167 ();
 sg13g2_decap_8 FILLER_39_180 ();
 sg13g2_fill_2 FILLER_39_187 ();
 sg13g2_fill_1 FILLER_39_189 ();
 sg13g2_decap_4 FILLER_39_194 ();
 sg13g2_decap_4 FILLER_39_235 ();
 sg13g2_fill_1 FILLER_39_249 ();
 sg13g2_decap_8 FILLER_39_254 ();
 sg13g2_decap_8 FILLER_39_261 ();
 sg13g2_fill_2 FILLER_39_268 ();
 sg13g2_fill_2 FILLER_39_278 ();
 sg13g2_fill_1 FILLER_39_289 ();
 sg13g2_fill_2 FILLER_39_307 ();
 sg13g2_fill_2 FILLER_39_388 ();
 sg13g2_fill_1 FILLER_40_0 ();
 sg13g2_decap_4 FILLER_40_28 ();
 sg13g2_fill_1 FILLER_40_40 ();
 sg13g2_fill_1 FILLER_40_54 ();
 sg13g2_fill_1 FILLER_40_60 ();
 sg13g2_decap_8 FILLER_40_82 ();
 sg13g2_fill_2 FILLER_40_89 ();
 sg13g2_decap_4 FILLER_40_96 ();
 sg13g2_fill_2 FILLER_40_100 ();
 sg13g2_decap_4 FILLER_40_126 ();
 sg13g2_fill_2 FILLER_40_164 ();
 sg13g2_decap_8 FILLER_40_170 ();
 sg13g2_fill_2 FILLER_40_177 ();
 sg13g2_fill_1 FILLER_40_179 ();
 sg13g2_decap_8 FILLER_40_184 ();
 sg13g2_decap_4 FILLER_40_198 ();
 sg13g2_decap_8 FILLER_40_206 ();
 sg13g2_decap_4 FILLER_40_213 ();
 sg13g2_fill_1 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_227 ();
 sg13g2_fill_1 FILLER_40_234 ();
 sg13g2_fill_2 FILLER_40_256 ();
 sg13g2_fill_1 FILLER_40_258 ();
 sg13g2_fill_1 FILLER_40_362 ();
 sg13g2_fill_1 FILLER_40_371 ();
 sg13g2_decap_4 FILLER_41_72 ();
 sg13g2_fill_1 FILLER_41_102 ();
 sg13g2_fill_1 FILLER_41_111 ();
 sg13g2_fill_2 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_165 ();
 sg13g2_fill_2 FILLER_41_172 ();
 sg13g2_decap_4 FILLER_41_212 ();
 sg13g2_fill_2 FILLER_41_216 ();
 sg13g2_fill_2 FILLER_41_232 ();
 sg13g2_fill_1 FILLER_41_234 ();
 sg13g2_fill_2 FILLER_41_244 ();
 sg13g2_fill_1 FILLER_41_246 ();
 sg13g2_fill_2 FILLER_41_273 ();
 sg13g2_decap_4 FILLER_41_300 ();
 sg13g2_fill_1 FILLER_41_318 ();
 sg13g2_fill_1 FILLER_41_345 ();
 sg13g2_fill_1 FILLER_41_352 ();
 sg13g2_fill_1 FILLER_41_356 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_fill_1 FILLER_42_9 ();
 sg13g2_decap_4 FILLER_42_14 ();
 sg13g2_fill_2 FILLER_42_18 ();
 sg13g2_decap_4 FILLER_42_28 ();
 sg13g2_fill_2 FILLER_42_37 ();
 sg13g2_decap_4 FILLER_42_50 ();
 sg13g2_fill_2 FILLER_42_54 ();
 sg13g2_decap_8 FILLER_42_61 ();
 sg13g2_decap_8 FILLER_42_68 ();
 sg13g2_decap_4 FILLER_42_75 ();
 sg13g2_fill_1 FILLER_42_118 ();
 sg13g2_fill_2 FILLER_42_129 ();
 sg13g2_fill_1 FILLER_42_131 ();
 sg13g2_decap_8 FILLER_42_141 ();
 sg13g2_fill_2 FILLER_42_148 ();
 sg13g2_fill_1 FILLER_42_150 ();
 sg13g2_fill_2 FILLER_42_193 ();
 sg13g2_fill_1 FILLER_42_224 ();
 sg13g2_fill_2 FILLER_42_233 ();
 sg13g2_decap_4 FILLER_42_243 ();
 sg13g2_fill_2 FILLER_42_252 ();
 sg13g2_fill_2 FILLER_42_269 ();
 sg13g2_fill_1 FILLER_42_330 ();
 sg13g2_fill_2 FILLER_42_343 ();
 sg13g2_fill_2 FILLER_42_393 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_4 ();
 sg13g2_decap_8 FILLER_43_30 ();
 sg13g2_fill_1 FILLER_43_37 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_fill_2 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_75 ();
 sg13g2_decap_8 FILLER_43_82 ();
 sg13g2_fill_1 FILLER_43_104 ();
 sg13g2_fill_2 FILLER_43_123 ();
 sg13g2_fill_2 FILLER_43_147 ();
 sg13g2_fill_1 FILLER_43_149 ();
 sg13g2_fill_1 FILLER_43_183 ();
 sg13g2_decap_8 FILLER_43_233 ();
 sg13g2_decap_4 FILLER_43_240 ();
 sg13g2_fill_2 FILLER_43_244 ();
 sg13g2_fill_1 FILLER_43_272 ();
 sg13g2_fill_2 FILLER_43_286 ();
 sg13g2_fill_2 FILLER_43_362 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_48 ();
 sg13g2_decap_8 FILLER_44_73 ();
 sg13g2_fill_2 FILLER_44_151 ();
 sg13g2_decap_8 FILLER_44_167 ();
 sg13g2_fill_2 FILLER_44_201 ();
 sg13g2_fill_2 FILLER_44_222 ();
 sg13g2_decap_8 FILLER_44_228 ();
 sg13g2_decap_8 FILLER_44_235 ();
 sg13g2_decap_4 FILLER_44_242 ();
 sg13g2_decap_8 FILLER_44_249 ();
 sg13g2_fill_2 FILLER_44_279 ();
 sg13g2_fill_1 FILLER_44_281 ();
 sg13g2_decap_4 FILLER_44_287 ();
 sg13g2_fill_1 FILLER_44_332 ();
 sg13g2_fill_1 FILLER_44_392 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_decap_4 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_65 ();
 sg13g2_fill_1 FILLER_45_146 ();
 sg13g2_fill_2 FILLER_45_187 ();
 sg13g2_fill_2 FILLER_45_194 ();
 sg13g2_fill_1 FILLER_45_217 ();
 sg13g2_fill_1 FILLER_45_258 ();
 sg13g2_fill_2 FILLER_45_303 ();
 sg13g2_fill_1 FILLER_45_342 ();
 sg13g2_fill_1 FILLER_45_364 ();
 sg13g2_decap_4 FILLER_46_28 ();
 sg13g2_fill_1 FILLER_46_32 ();
 sg13g2_fill_2 FILLER_46_67 ();
 sg13g2_fill_1 FILLER_46_120 ();
 sg13g2_fill_1 FILLER_46_133 ();
 sg13g2_fill_2 FILLER_46_139 ();
 sg13g2_fill_1 FILLER_46_141 ();
 sg13g2_fill_2 FILLER_46_156 ();
 sg13g2_fill_1 FILLER_46_162 ();
 sg13g2_fill_1 FILLER_46_198 ();
 sg13g2_decap_4 FILLER_46_212 ();
 sg13g2_decap_8 FILLER_46_220 ();
 sg13g2_fill_2 FILLER_46_227 ();
 sg13g2_fill_1 FILLER_46_378 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_4 ();
 sg13g2_fill_1 FILLER_47_36 ();
 sg13g2_fill_1 FILLER_47_45 ();
 sg13g2_decap_8 FILLER_47_61 ();
 sg13g2_decap_4 FILLER_47_68 ();
 sg13g2_fill_1 FILLER_47_98 ();
 sg13g2_decap_4 FILLER_47_156 ();
 sg13g2_decap_4 FILLER_47_168 ();
 sg13g2_fill_1 FILLER_47_172 ();
 sg13g2_fill_2 FILLER_47_182 ();
 sg13g2_decap_4 FILLER_47_219 ();
 sg13g2_fill_2 FILLER_47_223 ();
 sg13g2_fill_1 FILLER_47_251 ();
 sg13g2_fill_2 FILLER_47_314 ();
 sg13g2_fill_1 FILLER_47_382 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_4 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_11 ();
 sg13g2_decap_8 FILLER_48_16 ();
 sg13g2_decap_8 FILLER_48_53 ();
 sg13g2_fill_2 FILLER_48_60 ();
 sg13g2_decap_8 FILLER_48_66 ();
 sg13g2_fill_1 FILLER_48_73 ();
 sg13g2_fill_2 FILLER_48_95 ();
 sg13g2_fill_1 FILLER_48_97 ();
 sg13g2_fill_2 FILLER_48_131 ();
 sg13g2_fill_1 FILLER_48_137 ();
 sg13g2_decap_8 FILLER_48_146 ();
 sg13g2_decap_8 FILLER_48_153 ();
 sg13g2_fill_1 FILLER_48_160 ();
 sg13g2_fill_2 FILLER_48_166 ();
 sg13g2_fill_1 FILLER_48_209 ();
 sg13g2_fill_1 FILLER_48_221 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_fill_2 FILLER_48_318 ();
 sg13g2_fill_1 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_370 ();
 sg13g2_fill_2 FILLER_48_384 ();
 sg13g2_fill_1 FILLER_49_15 ();
 sg13g2_fill_2 FILLER_49_37 ();
 sg13g2_decap_8 FILLER_49_48 ();
 sg13g2_fill_2 FILLER_49_55 ();
 sg13g2_fill_1 FILLER_49_57 ();
 sg13g2_fill_2 FILLER_49_63 ();
 sg13g2_decap_4 FILLER_49_75 ();
 sg13g2_fill_2 FILLER_49_79 ();
 sg13g2_fill_2 FILLER_49_95 ();
 sg13g2_fill_1 FILLER_49_145 ();
 sg13g2_decap_8 FILLER_49_155 ();
 sg13g2_fill_2 FILLER_49_177 ();
 sg13g2_fill_2 FILLER_49_204 ();
 sg13g2_fill_1 FILLER_49_251 ();
 sg13g2_fill_2 FILLER_49_329 ();
 sg13g2_fill_1 FILLER_49_344 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_32 ();
 sg13g2_decap_8 FILLER_50_38 ();
 sg13g2_fill_1 FILLER_50_45 ();
 sg13g2_fill_1 FILLER_50_101 ();
 sg13g2_fill_1 FILLER_50_111 ();
 sg13g2_fill_2 FILLER_50_130 ();
 sg13g2_fill_2 FILLER_50_145 ();
 sg13g2_decap_4 FILLER_50_201 ();
 sg13g2_fill_1 FILLER_50_205 ();
 sg13g2_fill_1 FILLER_50_215 ();
 sg13g2_fill_1 FILLER_50_229 ();
 sg13g2_fill_1 FILLER_50_291 ();
 sg13g2_fill_2 FILLER_50_319 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_decap_4 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_32 ();
 sg13g2_fill_2 FILLER_51_43 ();
 sg13g2_fill_2 FILLER_51_134 ();
 sg13g2_fill_2 FILLER_51_207 ();
 sg13g2_fill_2 FILLER_51_218 ();
 sg13g2_fill_2 FILLER_51_281 ();
 sg13g2_fill_1 FILLER_51_303 ();
 sg13g2_fill_1 FILLER_51_309 ();
 sg13g2_fill_1 FILLER_51_340 ();
 sg13g2_fill_1 FILLER_51_346 ();
 sg13g2_fill_1 FILLER_51_361 ();
 sg13g2_fill_2 FILLER_52_27 ();
 sg13g2_fill_1 FILLER_52_46 ();
 sg13g2_fill_2 FILLER_52_71 ();
 sg13g2_fill_2 FILLER_52_107 ();
 sg13g2_fill_1 FILLER_52_159 ();
 sg13g2_decap_8 FILLER_52_169 ();
 sg13g2_fill_1 FILLER_52_176 ();
 sg13g2_fill_1 FILLER_52_187 ();
 sg13g2_fill_1 FILLER_52_193 ();
 sg13g2_fill_2 FILLER_52_215 ();
 sg13g2_fill_1 FILLER_52_294 ();
 sg13g2_fill_1 FILLER_52_308 ();
 sg13g2_fill_1 FILLER_52_345 ();
 sg13g2_fill_1 FILLER_52_356 ();
 sg13g2_fill_2 FILLER_52_383 ();
 sg13g2_fill_1 FILLER_52_403 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_28 ();
 sg13g2_fill_1 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_75 ();
 sg13g2_fill_2 FILLER_53_82 ();
 sg13g2_fill_1 FILLER_53_84 ();
 sg13g2_fill_1 FILLER_53_103 ();
 sg13g2_fill_2 FILLER_53_118 ();
 sg13g2_fill_2 FILLER_53_140 ();
 sg13g2_fill_1 FILLER_53_174 ();
 sg13g2_fill_1 FILLER_53_179 ();
 sg13g2_fill_2 FILLER_53_188 ();
 sg13g2_fill_1 FILLER_53_222 ();
 sg13g2_fill_1 FILLER_53_274 ();
 sg13g2_fill_2 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_360 ();
 sg13g2_fill_1 FILLER_53_370 ();
 sg13g2_fill_1 FILLER_53_402 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_fill_2 FILLER_54_6 ();
 sg13g2_fill_1 FILLER_54_21 ();
 sg13g2_fill_2 FILLER_54_52 ();
 sg13g2_decap_8 FILLER_54_68 ();
 sg13g2_decap_8 FILLER_54_75 ();
 sg13g2_decap_8 FILLER_54_82 ();
 sg13g2_fill_2 FILLER_54_89 ();
 sg13g2_fill_1 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_110 ();
 sg13g2_fill_2 FILLER_54_143 ();
 sg13g2_fill_1 FILLER_54_167 ();
 sg13g2_fill_1 FILLER_54_227 ();
 sg13g2_fill_2 FILLER_54_232 ();
 sg13g2_fill_2 FILLER_54_238 ();
 sg13g2_fill_2 FILLER_54_380 ();
 sg13g2_fill_2 FILLER_54_396 ();
 sg13g2_fill_2 FILLER_55_4 ();
 sg13g2_fill_1 FILLER_55_32 ();
 sg13g2_fill_2 FILLER_55_46 ();
 sg13g2_fill_2 FILLER_55_61 ();
 sg13g2_decap_8 FILLER_55_78 ();
 sg13g2_fill_1 FILLER_55_85 ();
 sg13g2_fill_1 FILLER_55_127 ();
 sg13g2_fill_1 FILLER_55_216 ();
 sg13g2_fill_2 FILLER_55_235 ();
 sg13g2_fill_2 FILLER_55_300 ();
 sg13g2_fill_1 FILLER_55_386 ();
 sg13g2_fill_2 FILLER_55_396 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_10 ();
 sg13g2_fill_1 FILLER_56_17 ();
 sg13g2_fill_1 FILLER_56_30 ();
 sg13g2_fill_1 FILLER_56_35 ();
 sg13g2_fill_2 FILLER_56_42 ();
 sg13g2_fill_2 FILLER_56_73 ();
 sg13g2_fill_1 FILLER_56_75 ();
 sg13g2_fill_2 FILLER_56_83 ();
 sg13g2_fill_1 FILLER_56_85 ();
 sg13g2_fill_1 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_188 ();
 sg13g2_fill_2 FILLER_56_291 ();
 sg13g2_fill_1 FILLER_56_320 ();
 sg13g2_fill_1 FILLER_56_336 ();
 sg13g2_fill_1 FILLER_57_4 ();
 sg13g2_fill_1 FILLER_57_30 ();
 sg13g2_fill_1 FILLER_57_80 ();
 sg13g2_fill_2 FILLER_57_243 ();
 sg13g2_fill_1 FILLER_57_284 ();
 sg13g2_fill_1 FILLER_57_319 ();
 sg13g2_fill_1 FILLER_57_341 ();
 sg13g2_fill_2 FILLER_58_40 ();
 sg13g2_fill_2 FILLER_58_48 ();
 sg13g2_fill_2 FILLER_58_62 ();
 sg13g2_fill_1 FILLER_58_145 ();
 sg13g2_fill_2 FILLER_58_159 ();
 sg13g2_fill_1 FILLER_58_308 ();
 sg13g2_fill_1 FILLER_58_326 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_26 ();
 sg13g2_fill_2 FILLER_59_75 ();
 sg13g2_fill_1 FILLER_59_80 ();
 sg13g2_fill_1 FILLER_59_86 ();
 sg13g2_fill_2 FILLER_59_133 ();
 sg13g2_fill_1 FILLER_59_231 ();
 sg13g2_fill_1 FILLER_59_256 ();
 sg13g2_fill_1 FILLER_59_274 ();
 sg13g2_fill_2 FILLER_59_343 ();
 sg13g2_fill_1 FILLER_59_354 ();
 sg13g2_fill_1 FILLER_60_36 ();
 sg13g2_fill_1 FILLER_60_60 ();
 sg13g2_fill_1 FILLER_60_130 ();
 sg13g2_fill_2 FILLER_60_151 ();
 sg13g2_fill_1 FILLER_60_243 ();
 sg13g2_fill_2 FILLER_60_294 ();
 sg13g2_fill_2 FILLER_60_322 ();
 sg13g2_fill_2 FILLER_60_381 ();
 sg13g2_fill_1 FILLER_61_10 ();
 sg13g2_fill_1 FILLER_61_36 ();
 sg13g2_fill_1 FILLER_61_45 ();
 sg13g2_fill_2 FILLER_61_186 ();
 sg13g2_fill_1 FILLER_61_264 ();
 sg13g2_fill_1 FILLER_61_291 ();
 sg13g2_fill_2 FILLER_61_345 ();
 sg13g2_fill_1 FILLER_61_368 ();
 sg13g2_fill_1 FILLER_61_383 ();
 sg13g2_fill_1 FILLER_62_86 ();
 sg13g2_fill_1 FILLER_62_106 ();
 sg13g2_fill_1 FILLER_62_120 ();
 sg13g2_fill_2 FILLER_62_127 ();
 sg13g2_fill_1 FILLER_62_185 ();
 sg13g2_fill_2 FILLER_62_281 ();
 sg13g2_fill_2 FILLER_62_352 ();
 sg13g2_fill_1 FILLER_63_29 ();
 sg13g2_fill_2 FILLER_63_62 ();
 sg13g2_fill_1 FILLER_63_80 ();
 sg13g2_fill_1 FILLER_63_104 ();
 sg13g2_fill_2 FILLER_63_160 ();
 sg13g2_fill_1 FILLER_63_283 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_fill_1 FILLER_64_15 ();
 sg13g2_fill_1 FILLER_64_24 ();
 sg13g2_fill_2 FILLER_64_41 ();
 sg13g2_fill_1 FILLER_64_88 ();
 sg13g2_fill_1 FILLER_64_94 ();
 sg13g2_fill_1 FILLER_64_136 ();
 sg13g2_fill_1 FILLER_64_155 ();
 sg13g2_fill_2 FILLER_64_180 ();
 sg13g2_fill_2 FILLER_64_213 ();
 sg13g2_fill_1 FILLER_64_331 ();
 sg13g2_fill_2 FILLER_64_338 ();
 sg13g2_fill_1 FILLER_65_46 ();
 sg13g2_fill_1 FILLER_65_104 ();
 sg13g2_fill_1 FILLER_65_161 ();
 sg13g2_fill_1 FILLER_65_188 ();
 sg13g2_fill_1 FILLER_65_204 ();
 sg13g2_fill_1 FILLER_65_241 ();
 sg13g2_fill_1 FILLER_65_280 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_34 ();
 sg13g2_fill_1 FILLER_66_61 ();
 sg13g2_fill_1 FILLER_66_96 ();
 sg13g2_fill_2 FILLER_66_154 ();
 sg13g2_fill_1 FILLER_66_182 ();
 sg13g2_fill_1 FILLER_66_189 ();
 sg13g2_fill_1 FILLER_66_308 ();
 sg13g2_fill_1 FILLER_66_337 ();
 sg13g2_fill_1 FILLER_66_382 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_14 ();
 sg13g2_fill_1 FILLER_67_68 ();
 sg13g2_fill_2 FILLER_67_85 ();
 sg13g2_fill_1 FILLER_67_143 ();
 sg13g2_fill_1 FILLER_67_206 ();
 sg13g2_fill_2 FILLER_67_270 ();
 sg13g2_fill_2 FILLER_67_292 ();
 sg13g2_fill_1 FILLER_67_327 ();
 sg13g2_fill_1 FILLER_68_42 ();
 sg13g2_fill_1 FILLER_68_70 ();
 sg13g2_fill_1 FILLER_68_173 ();
 sg13g2_fill_2 FILLER_68_200 ();
 sg13g2_fill_2 FILLER_68_207 ();
 sg13g2_fill_2 FILLER_68_255 ();
 sg13g2_fill_2 FILLER_68_288 ();
 sg13g2_fill_1 FILLER_68_387 ();
 sg13g2_fill_2 FILLER_69_26 ();
 sg13g2_fill_1 FILLER_69_33 ();
 sg13g2_fill_1 FILLER_69_37 ();
 sg13g2_fill_1 FILLER_69_127 ();
 sg13g2_fill_2 FILLER_69_187 ();
 sg13g2_fill_2 FILLER_69_197 ();
 sg13g2_fill_1 FILLER_69_213 ();
 sg13g2_fill_1 FILLER_69_289 ();
 sg13g2_fill_2 FILLER_69_330 ();
 sg13g2_fill_2 FILLER_69_351 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_fill_1 FILLER_70_4 ();
 sg13g2_fill_1 FILLER_70_21 ();
 sg13g2_fill_2 FILLER_70_46 ();
 sg13g2_fill_2 FILLER_70_99 ();
 sg13g2_fill_1 FILLER_70_118 ();
 sg13g2_fill_2 FILLER_70_183 ();
 sg13g2_fill_2 FILLER_70_193 ();
 sg13g2_fill_2 FILLER_70_205 ();
 sg13g2_fill_1 FILLER_70_251 ();
 sg13g2_fill_1 FILLER_70_369 ();
 sg13g2_fill_1 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_127 ();
 sg13g2_fill_2 FILLER_71_167 ();
 sg13g2_fill_1 FILLER_71_188 ();
 sg13g2_fill_1 FILLER_71_385 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_78 ();
 sg13g2_fill_1 FILLER_72_198 ();
 sg13g2_fill_2 FILLER_72_269 ();
 sg13g2_fill_1 FILLER_72_286 ();
 sg13g2_fill_2 FILLER_72_341 ();
 sg13g2_fill_2 FILLER_72_357 ();
 sg13g2_fill_1 FILLER_72_382 ();
 sg13g2_fill_1 FILLER_73_4 ();
 sg13g2_fill_1 FILLER_73_36 ();
 sg13g2_fill_1 FILLER_73_125 ();
 sg13g2_fill_2 FILLER_73_223 ();
 sg13g2_fill_1 FILLER_73_258 ();
 sg13g2_fill_1 FILLER_73_283 ();
 sg13g2_fill_1 FILLER_73_356 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_45 ();
 sg13g2_fill_1 FILLER_74_60 ();
 sg13g2_fill_1 FILLER_74_133 ();
 sg13g2_fill_2 FILLER_74_149 ();
 sg13g2_fill_1 FILLER_74_200 ();
 sg13g2_fill_2 FILLER_74_225 ();
 sg13g2_fill_2 FILLER_74_232 ();
 sg13g2_fill_2 FILLER_74_242 ();
 sg13g2_fill_1 FILLER_74_249 ();
 sg13g2_fill_1 FILLER_74_255 ();
 sg13g2_fill_1 FILLER_74_355 ();
 sg13g2_fill_1 FILLER_74_375 ();
 sg13g2_fill_1 FILLER_74_408 ();
 sg13g2_fill_1 FILLER_75_170 ();
 sg13g2_fill_1 FILLER_75_200 ();
 sg13g2_fill_2 FILLER_75_226 ();
 sg13g2_fill_2 FILLER_75_305 ();
 sg13g2_fill_2 FILLER_75_341 ();
 sg13g2_fill_1 FILLER_76_11 ();
 sg13g2_fill_2 FILLER_76_73 ();
 sg13g2_fill_2 FILLER_76_99 ();
 sg13g2_fill_2 FILLER_76_131 ();
 sg13g2_fill_1 FILLER_76_287 ();
 sg13g2_fill_2 FILLER_76_300 ();
 sg13g2_fill_2 FILLER_76_338 ();
 sg13g2_fill_1 FILLER_76_347 ();
 sg13g2_fill_1 FILLER_76_392 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_fill_1 FILLER_77_62 ();
 sg13g2_fill_1 FILLER_77_173 ();
 sg13g2_fill_2 FILLER_77_253 ();
 sg13g2_fill_1 FILLER_77_272 ();
 sg13g2_fill_1 FILLER_77_287 ();
 sg13g2_fill_1 FILLER_78_11 ();
 sg13g2_fill_1 FILLER_78_144 ();
 sg13g2_fill_1 FILLER_78_154 ();
 sg13g2_fill_1 FILLER_78_190 ();
 sg13g2_fill_1 FILLER_78_196 ();
 sg13g2_fill_2 FILLER_78_260 ();
 sg13g2_fill_2 FILLER_78_306 ();
 sg13g2_fill_1 FILLER_78_339 ();
 sg13g2_fill_1 FILLER_79_38 ();
 sg13g2_fill_2 FILLER_79_164 ();
 sg13g2_fill_2 FILLER_79_227 ();
 sg13g2_fill_1 FILLER_79_315 ();
 sg13g2_fill_1 FILLER_79_360 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_44 ();
 sg13g2_fill_2 FILLER_80_69 ();
 sg13g2_fill_1 FILLER_80_80 ();
 sg13g2_fill_2 FILLER_80_90 ();
 sg13g2_fill_1 FILLER_80_119 ();
 sg13g2_fill_2 FILLER_80_133 ();
 sg13g2_fill_2 FILLER_80_206 ();
 sg13g2_fill_1 FILLER_80_348 ();
 sg13g2_fill_1 FILLER_80_376 ();
 assign uio_oe[0] = net8;
 assign uio_oe[1] = net9;
 assign uio_oe[2] = net10;
 assign uio_oe[3] = net11;
 assign uio_oe[4] = net12;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
 assign uio_out[7] = net23;
 assign uo_out[7] = net24;
endmodule
