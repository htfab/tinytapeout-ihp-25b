module tt_um_tinytapeout_logo_screensaver (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire clknet_0_clk;
 wire \color_index[0] ;
 wire \color_index[1] ;
 wire \color_index[2] ;
 wire dir_x;
 wire dir_y;
 wire \gamepad.decoder.data_reg[0] ;
 wire \gamepad.decoder.data_reg[10] ;
 wire \gamepad.decoder.data_reg[11] ;
 wire \gamepad.decoder.data_reg[1] ;
 wire \gamepad.decoder.data_reg[2] ;
 wire \gamepad.decoder.data_reg[3] ;
 wire \gamepad.decoder.data_reg[4] ;
 wire \gamepad.decoder.data_reg[5] ;
 wire \gamepad.decoder.data_reg[6] ;
 wire \gamepad.decoder.data_reg[7] ;
 wire \gamepad.decoder.data_reg[8] ;
 wire \gamepad.decoder.data_reg[9] ;
 wire \gamepad.driver.pmod_clk_prev ;
 wire \gamepad.driver.pmod_clk_sync[0] ;
 wire \gamepad.driver.pmod_clk_sync[1] ;
 wire \gamepad.driver.pmod_data_sync[0] ;
 wire \gamepad.driver.pmod_data_sync[1] ;
 wire \gamepad.driver.pmod_latch_prev ;
 wire \gamepad.driver.pmod_latch_sync[0] ;
 wire \gamepad.driver.pmod_latch_sync[1] ;
 wire \gamepad.driver.shift_reg[0] ;
 wire \gamepad.driver.shift_reg[10] ;
 wire \gamepad.driver.shift_reg[11] ;
 wire \gamepad.driver.shift_reg[1] ;
 wire \gamepad.driver.shift_reg[2] ;
 wire \gamepad.driver.shift_reg[3] ;
 wire \gamepad.driver.shift_reg[4] ;
 wire \gamepad.driver.shift_reg[5] ;
 wire \gamepad.driver.shift_reg[6] ;
 wire \gamepad.driver.shift_reg[7] ;
 wire \gamepad.driver.shift_reg[8] ;
 wire \gamepad.driver.shift_reg[9] ;
 wire gamepad_start_prev;
 wire hsync;
 wire \logo_left[0] ;
 wire \logo_left[1] ;
 wire \logo_left[2] ;
 wire \logo_left[3] ;
 wire \logo_left[4] ;
 wire \logo_left[5] ;
 wire \logo_left[6] ;
 wire \logo_left[7] ;
 wire \logo_left[8] ;
 wire \logo_left[9] ;
 wire \logo_top[0] ;
 wire \logo_top[1] ;
 wire \logo_top[2] ;
 wire \logo_top[3] ;
 wire \logo_top[4] ;
 wire \logo_top[5] ;
 wire \logo_top[6] ;
 wire \logo_top[7] ;
 wire \logo_top[8] ;
 wire \logo_top[9] ;
 wire manual_mode;
 wire \palette_inst.rrggbb[0] ;
 wire \palette_inst.rrggbb[1] ;
 wire \palette_inst.rrggbb[2] ;
 wire \palette_inst.rrggbb[3] ;
 wire \palette_inst.rrggbb[4] ;
 wire \palette_inst.rrggbb[5] ;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire \prev_y[0] ;
 wire \prev_y[1] ;
 wire \prev_y[2] ;
 wire \prev_y[3] ;
 wire \prev_y[4] ;
 wire \prev_y[5] ;
 wire \prev_y[6] ;
 wire \prev_y[7] ;
 wire \prev_y[8] ;
 wire \prev_y[9] ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire \vga_sync_gen.vsync ;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;

 sg13g2_inv_1 _1685_ (.Y(_0721_),
    .A(net176));
 sg13g2_inv_1 _1686_ (.Y(_0722_),
    .A(net179));
 sg13g2_inv_1 _1687_ (.Y(_0723_),
    .A(net169));
 sg13g2_inv_1 _1688_ (.Y(_0724_),
    .A(net175));
 sg13g2_inv_1 _1689_ (.Y(_0725_),
    .A(net165));
 sg13g2_inv_1 _1690_ (.Y(_0726_),
    .A(net182));
 sg13g2_inv_1 _1691_ (.Y(_0727_),
    .A(net171));
 sg13g2_inv_1 _1692_ (.Y(_0728_),
    .A(net194));
 sg13g2_inv_1 _1693_ (.Y(_0729_),
    .A(net193));
 sg13g2_inv_1 _1694_ (.Y(_0730_),
    .A(net184));
 sg13g2_inv_1 _1695_ (.Y(_0731_),
    .A(\gamepad.driver.shift_reg[0] ));
 sg13g2_inv_1 _1696_ (.Y(_0732_),
    .A(net153));
 sg13g2_inv_1 _1697_ (.Y(_0733_),
    .A(net826));
 sg13g2_inv_2 _1698_ (.Y(_0734_),
    .A(net831));
 sg13g2_inv_2 _1699_ (.Y(_0735_),
    .A(net833));
 sg13g2_inv_1 _1700_ (.Y(_0736_),
    .A(\logo_top[8] ));
 sg13g2_inv_2 _1701_ (.Y(_0737_),
    .A(\logo_top[7] ));
 sg13g2_inv_1 _1702_ (.Y(_0738_),
    .A(\logo_top[4] ));
 sg13g2_inv_1 _1703_ (.Y(_0739_),
    .A(\logo_top[3] ));
 sg13g2_inv_1 _1704_ (.Y(_0740_),
    .A(net132));
 sg13g2_inv_2 _1705_ (.Y(_0741_),
    .A(\logo_left[5] ));
 sg13g2_inv_1 _1706_ (.Y(_0742_),
    .A(\logo_left[4] ));
 sg13g2_inv_1 _1707_ (.Y(_0743_),
    .A(net841));
 sg13g2_inv_1 _1708_ (.Y(_0744_),
    .A(\logo_left[2] ));
 sg13g2_inv_1 _1709_ (.Y(_0745_),
    .A(net136));
 sg13g2_inv_1 _1710_ (.Y(_0746_),
    .A(net149));
 sg13g2_inv_1 _1711_ (.Y(_0747_),
    .A(\pix_y[4] ));
 sg13g2_inv_1 _1712_ (.Y(_0748_),
    .A(net817));
 sg13g2_inv_1 _1713_ (.Y(_0749_),
    .A(net213));
 sg13g2_inv_1 _1714_ (.Y(_0750_),
    .A(net851));
 sg13g2_inv_2 _1715_ (.Y(_0751_),
    .A(net214));
 sg13g2_inv_1 _1716_ (.Y(_0752_),
    .A(net178));
 sg13g2_inv_2 _1717_ (.Y(_0753_),
    .A(net816));
 sg13g2_inv_1 _1718_ (.Y(_0754_),
    .A(\prev_y[0] ));
 sg13g2_inv_1 _1719_ (.Y(_0755_),
    .A(\prev_y[6] ));
 sg13g2_inv_1 _1720_ (.Y(_0756_),
    .A(\prev_y[8] ));
 sg13g2_inv_1 _1721_ (.Y(_0757_),
    .A(\prev_y[9] ));
 sg13g2_inv_1 _1722_ (.Y(_0758_),
    .A(net160));
 sg13g2_inv_1 _1723_ (.Y(_0759_),
    .A(net156));
 sg13g2_inv_1 _1724_ (.Y(_0760_),
    .A(net158));
 sg13g2_inv_1 _1725_ (.Y(_0761_),
    .A(net147));
 sg13g2_inv_1 _1726_ (.Y(_0762_),
    .A(net167));
 sg13g2_inv_1 _1727_ (.Y(_0763_),
    .A(net189));
 sg13g2_inv_1 _1728_ (.Y(_0764_),
    .A(net181));
 sg13g2_inv_1 _1729_ (.Y(_0765_),
    .A(net187));
 sg13g2_inv_1 _1730_ (.Y(_0766_),
    .A(net145));
 sg13g2_inv_1 _1731_ (.Y(_0767_),
    .A(net186));
 sg13g2_inv_1 _1732_ (.Y(_0768_),
    .A(net155));
 sg13g2_inv_1 _1733_ (.Y(_0769_),
    .A(net151));
 sg13g2_inv_1 _1734_ (.Y(_0770_),
    .A(_0010_));
 sg13g2_inv_1 _1735_ (.Y(_0771_),
    .A(_0011_));
 sg13g2_inv_1 _1736_ (.Y(_0772_),
    .A(net2));
 sg13g2_nand2_1 _1737_ (.Y(_0773_),
    .A(net817),
    .B(\pix_y[6] ));
 sg13g2_nor3_2 _1738_ (.A(_0751_),
    .B(_0753_),
    .C(_0773_),
    .Y(_0774_));
 sg13g2_nand4_1 _1739_ (.B(\pix_y[6] ),
    .C(net221),
    .A(net817),
    .Y(_0775_),
    .D(net203));
 sg13g2_nand3b_1 _1740_ (.B(net820),
    .C(net162),
    .Y(_0776_),
    .A_N(\pix_y[2] ));
 sg13g2_nor4_1 _1741_ (.A(net819),
    .B(net815),
    .C(_0775_),
    .D(net163),
    .Y(_0006_));
 sg13g2_and3_1 _1742_ (.X(_0777_),
    .A(\pix_x[4] ),
    .B(\pix_x[5] ),
    .C(net197));
 sg13g2_nor3_1 _1743_ (.A(\pix_x[4] ),
    .B(\pix_x[5] ),
    .C(net197),
    .Y(_0778_));
 sg13g2_nand2_1 _1744_ (.Y(_0779_),
    .A(\pix_x[7] ),
    .B(\pix_x[9] ));
 sg13g2_nor4_1 _1745_ (.A(net199),
    .B(_0777_),
    .C(_0778_),
    .D(_0779_),
    .Y(_0005_));
 sg13g2_nand2b_1 _1746_ (.Y(_0780_),
    .B(\prev_y[1] ),
    .A_N(\pix_y[1] ));
 sg13g2_nand2b_1 _1747_ (.Y(_0781_),
    .B(net816),
    .A_N(\prev_y[7] ));
 sg13g2_nand2b_1 _1748_ (.Y(_0782_),
    .B(net823),
    .A_N(\prev_y[1] ));
 sg13g2_nand2b_1 _1749_ (.Y(_0783_),
    .B(net817),
    .A_N(\prev_y[5] ));
 sg13g2_a22oi_1 _1750_ (.Y(_0784_),
    .B1(\prev_y[8] ),
    .B2(_0751_),
    .A2(\prev_y[4] ),
    .A1(_0747_));
 sg13g2_a22oi_1 _1751_ (.Y(_0785_),
    .B1(_0756_),
    .B2(\pix_y[8] ),
    .A2(\prev_y[7] ),
    .A1(_0753_));
 sg13g2_nand2b_1 _1752_ (.Y(_0786_),
    .B(net819),
    .A_N(\prev_y[4] ));
 sg13g2_xnor2_1 _1753_ (.Y(_0787_),
    .A(net820),
    .B(\prev_y[3] ));
 sg13g2_xnor2_1 _1754_ (.Y(_0788_),
    .A(\pix_y[2] ),
    .B(\prev_y[2] ));
 sg13g2_o21ai_1 _1755_ (.B1(_0782_),
    .Y(_0789_),
    .A1(\pix_y[0] ),
    .A2(_0754_));
 sg13g2_a221oi_1 _1756_ (.B2(\pix_y[6] ),
    .C1(_0789_),
    .B1(_0755_),
    .A1(\pix_y[0] ),
    .Y(_0790_),
    .A2(_0754_));
 sg13g2_a22oi_1 _1757_ (.Y(_0791_),
    .B1(_0757_),
    .B2(net815),
    .A2(\prev_y[6] ),
    .A1(_0749_));
 sg13g2_nand4_1 _1758_ (.B(_0784_),
    .C(_0786_),
    .A(_0783_),
    .Y(_0792_),
    .D(_0791_));
 sg13g2_a221oi_1 _1759_ (.B2(_0752_),
    .C1(_0792_),
    .B1(\prev_y[9] ),
    .A1(_0748_),
    .Y(_0793_),
    .A2(\prev_y[5] ));
 sg13g2_and4_1 _1760_ (.A(_0780_),
    .B(_0781_),
    .C(_0785_),
    .D(_0793_),
    .X(_0794_));
 sg13g2_nand4_1 _1761_ (.B(_0788_),
    .C(_0790_),
    .A(_0787_),
    .Y(_0795_),
    .D(_0794_));
 sg13g2_nor4_1 _1762_ (.A(net819),
    .B(net818),
    .C(\pix_y[6] ),
    .D(net816),
    .Y(_0796_));
 sg13g2_nor2_1 _1763_ (.A(net824),
    .B(net823),
    .Y(_0797_));
 sg13g2_nor4_1 _1764_ (.A(net822),
    .B(net821),
    .C(\pix_y[8] ),
    .D(net815),
    .Y(_0798_));
 sg13g2_nand4_1 _1765_ (.B(_0796_),
    .C(_0797_),
    .A(_0795_),
    .Y(_0799_),
    .D(_0798_));
 sg13g2_inv_1 _1766_ (.Y(_0800_),
    .A(_0799_));
 sg13g2_nor2_2 _1767_ (.A(net828),
    .B(_0799_),
    .Y(_0801_));
 sg13g2_inv_1 _1768_ (.Y(_0802_),
    .A(_0801_));
 sg13g2_nand2_2 _1769_ (.Y(_0803_),
    .A(\logo_top[1] ),
    .B(\logo_top[0] ));
 sg13g2_nand3_1 _1770_ (.B(\logo_top[1] ),
    .C(\logo_top[0] ),
    .A(net836),
    .Y(_0804_));
 sg13g2_and4_1 _1771_ (.A(\logo_top[3] ),
    .B(net836),
    .C(net837),
    .D(net838),
    .X(_0805_));
 sg13g2_nand3_1 _1772_ (.B(\logo_top[4] ),
    .C(_0805_),
    .A(net835),
    .Y(_0806_));
 sg13g2_inv_1 _1773_ (.Y(_0807_),
    .A(_0806_));
 sg13g2_nor2_1 _1774_ (.A(_0013_),
    .B(_0806_),
    .Y(_0808_));
 sg13g2_xor2_1 _1775_ (.B(_0806_),
    .A(_0013_),
    .X(_0809_));
 sg13g2_xnor2_1 _1776_ (.Y(_0810_),
    .A(\logo_top[7] ),
    .B(_0808_));
 sg13g2_inv_1 _1777_ (.Y(_0811_),
    .A(_0810_));
 sg13g2_nor2_1 _1778_ (.A(_0809_),
    .B(_0811_),
    .Y(_0812_));
 sg13g2_and3_1 _1779_ (.X(_0813_),
    .A(\logo_top[7] ),
    .B(\logo_top[6] ),
    .C(_0807_));
 sg13g2_nand2b_1 _1780_ (.Y(_0814_),
    .B(_0014_),
    .A_N(_0813_));
 sg13g2_nand3b_1 _1781_ (.B(_0813_),
    .C(net834),
    .Y(_0815_),
    .A_N(_0014_));
 sg13g2_o21ai_1 _1782_ (.B1(_0815_),
    .Y(_0816_),
    .A1(net834),
    .A2(_0814_));
 sg13g2_nor2_2 _1783_ (.A(net837),
    .B(net838),
    .Y(_0817_));
 sg13g2_nand2_1 _1784_ (.Y(_0818_),
    .A(_0011_),
    .B(_0817_));
 sg13g2_xnor2_1 _1785_ (.Y(_0819_),
    .A(_0739_),
    .B(_0818_));
 sg13g2_nor4_1 _1786_ (.A(net831),
    .B(net835),
    .C(net837),
    .D(_0771_),
    .Y(_0820_));
 sg13g2_and4_1 _1787_ (.A(_0739_),
    .B(net838),
    .C(_0012_),
    .D(_0820_),
    .X(_0821_));
 sg13g2_nand3_1 _1788_ (.B(_0816_),
    .C(_0821_),
    .A(_0812_),
    .Y(_0822_));
 sg13g2_xnor2_1 _1789_ (.Y(_0823_),
    .A(_0014_),
    .B(_0813_));
 sg13g2_nand2b_1 _1790_ (.Y(_0824_),
    .B(_0823_),
    .A_N(net834));
 sg13g2_nand2_1 _1791_ (.Y(_0825_),
    .A(_0737_),
    .B(_0809_));
 sg13g2_inv_1 _1792_ (.Y(_0826_),
    .A(_0825_));
 sg13g2_a21oi_1 _1793_ (.A1(\logo_top[4] ),
    .A2(_0805_),
    .Y(_0827_),
    .B1(net835));
 sg13g2_or2_1 _1794_ (.X(_0828_),
    .B(_0827_),
    .A(_0807_));
 sg13g2_xnor2_1 _1795_ (.Y(_0829_),
    .A(_0012_),
    .B(_0805_));
 sg13g2_nor2_1 _1796_ (.A(_0011_),
    .B(_0803_),
    .Y(_0830_));
 sg13g2_xnor2_1 _1797_ (.Y(_0831_),
    .A(_0739_),
    .B(_0830_));
 sg13g2_or4_1 _1798_ (.A(_0804_),
    .B(_0828_),
    .C(_0829_),
    .D(_0831_),
    .X(_0832_));
 sg13g2_nor3_2 _1799_ (.A(_0824_),
    .B(_0825_),
    .C(_0832_),
    .Y(_0833_));
 sg13g2_nand2_1 _1800_ (.Y(_0834_),
    .A(net831),
    .B(_0833_));
 sg13g2_and2_1 _1801_ (.A(_0822_),
    .B(_0834_),
    .X(_0835_));
 sg13g2_nor2_2 _1802_ (.A(net842),
    .B(net843),
    .Y(_0836_));
 sg13g2_nor4_2 _1803_ (.A(\logo_left[3] ),
    .B(\logo_left[2] ),
    .C(\logo_left[1] ),
    .Y(_0837_),
    .D(net843));
 sg13g2_nand2_1 _1804_ (.Y(_0838_),
    .A(_0008_),
    .B(_0837_));
 sg13g2_xnor2_1 _1805_ (.Y(_0839_),
    .A(_0008_),
    .B(_0837_));
 sg13g2_nand2_1 _1806_ (.Y(_0840_),
    .A(_0007_),
    .B(_0836_));
 sg13g2_xnor2_1 _1807_ (.Y(_0841_),
    .A(net841),
    .B(_0840_));
 sg13g2_nand2_1 _1808_ (.Y(_0842_),
    .A(\logo_left[0] ),
    .B(_0007_));
 sg13g2_or4_1 _1809_ (.A(net833),
    .B(\logo_left[9] ),
    .C(net842),
    .D(_0842_),
    .X(_0843_));
 sg13g2_nor3_1 _1810_ (.A(_0839_),
    .B(_0841_),
    .C(_0843_),
    .Y(_0844_));
 sg13g2_nor2_1 _1811_ (.A(\logo_left[5] ),
    .B(\logo_left[4] ),
    .Y(_0845_));
 sg13g2_nand2_1 _1812_ (.Y(_0846_),
    .A(_0837_),
    .B(_0845_));
 sg13g2_nand3_1 _1813_ (.B(_0837_),
    .C(_0845_),
    .A(_0009_),
    .Y(_0847_));
 sg13g2_xnor2_1 _1814_ (.Y(_0848_),
    .A(_0009_),
    .B(_0846_));
 sg13g2_xnor2_1 _1815_ (.Y(_0849_),
    .A(_0741_),
    .B(_0838_));
 sg13g2_or3_2 _1816_ (.A(net839),
    .B(net840),
    .C(_0846_),
    .X(_0850_));
 sg13g2_nor2_1 _1817_ (.A(_0770_),
    .B(_0850_),
    .Y(_0851_));
 sg13g2_xnor2_1 _1818_ (.Y(_0852_),
    .A(_0770_),
    .B(_0850_));
 sg13g2_xor2_1 _1819_ (.B(_0847_),
    .A(net839),
    .X(_0853_));
 sg13g2_nor2b_1 _1820_ (.A(_0852_),
    .B_N(_0853_),
    .Y(_0854_));
 sg13g2_nand4_1 _1821_ (.B(_0848_),
    .C(_0849_),
    .A(_0844_),
    .Y(_0855_),
    .D(_0854_));
 sg13g2_nand2_2 _1822_ (.Y(_0856_),
    .A(net842),
    .B(net843));
 sg13g2_nand4_1 _1823_ (.B(\logo_left[2] ),
    .C(net842),
    .A(\logo_left[3] ),
    .Y(_0857_),
    .D(net843));
 sg13g2_nand2_1 _1824_ (.Y(_0858_),
    .A(\logo_left[5] ),
    .B(\logo_left[4] ));
 sg13g2_nor2_1 _1825_ (.A(_0857_),
    .B(_0858_),
    .Y(_0859_));
 sg13g2_and3_1 _1826_ (.X(_0860_),
    .A(net839),
    .B(net840),
    .C(_0859_));
 sg13g2_and2_1 _1827_ (.A(_0770_),
    .B(_0860_),
    .X(_0861_));
 sg13g2_xnor2_1 _1828_ (.Y(_0862_),
    .A(\logo_left[9] ),
    .B(_0861_));
 sg13g2_xnor2_1 _1829_ (.Y(_0863_),
    .A(net840),
    .B(_0859_));
 sg13g2_nor2_1 _1830_ (.A(_0008_),
    .B(_0857_),
    .Y(_0864_));
 sg13g2_xnor2_1 _1831_ (.Y(_0865_),
    .A(_0741_),
    .B(_0864_));
 sg13g2_xnor2_1 _1832_ (.Y(_0866_),
    .A(_0742_),
    .B(_0857_));
 sg13g2_nor2_1 _1833_ (.A(_0007_),
    .B(_0856_),
    .Y(_0867_));
 sg13g2_xnor2_1 _1834_ (.Y(_0868_),
    .A(net841),
    .B(_0867_));
 sg13g2_nor3_1 _1835_ (.A(_0735_),
    .B(_0744_),
    .C(_0856_),
    .Y(_0869_));
 sg13g2_nand4_1 _1836_ (.B(_0866_),
    .C(_0868_),
    .A(_0863_),
    .Y(_0870_),
    .D(_0869_));
 sg13g2_or2_1 _1837_ (.X(_0871_),
    .B(_0870_),
    .A(_0865_));
 sg13g2_nor3_1 _1838_ (.A(_0009_),
    .B(_0857_),
    .C(_0858_),
    .Y(_0872_));
 sg13g2_xnor2_1 _1839_ (.Y(_0873_),
    .A(net839),
    .B(_0872_));
 sg13g2_xor2_1 _1840_ (.B(_0860_),
    .A(\logo_left[8] ),
    .X(_0874_));
 sg13g2_nand3_1 _1841_ (.B(\logo_left[8] ),
    .C(_0860_),
    .A(\logo_left[9] ),
    .Y(_0875_));
 sg13g2_nand2_1 _1842_ (.Y(_0876_),
    .A(_0873_),
    .B(_0875_));
 sg13g2_or4_1 _1843_ (.A(_0862_),
    .B(_0871_),
    .C(_0874_),
    .D(_0876_),
    .X(_0877_));
 sg13g2_nand3_1 _1844_ (.B(_0855_),
    .C(_0877_),
    .A(_0835_),
    .Y(_0878_));
 sg13g2_nand2_2 _1845_ (.Y(_0879_),
    .A(_0801_),
    .B(_0878_));
 sg13g2_inv_1 _1846_ (.Y(_0880_),
    .A(_0879_));
 sg13g2_xor2_1 _1847_ (.B(_0879_),
    .A(net134),
    .X(_0881_));
 sg13g2_inv_1 _1848_ (.Y(_0882_),
    .A(_0881_));
 sg13g2_and2_1 _1849_ (.A(net850),
    .B(_0881_),
    .X(_0883_));
 sg13g2_nand2_1 _1850_ (.Y(_0884_),
    .A(net173),
    .B(\color_index[0] ));
 sg13g2_xor2_1 _1851_ (.B(_0884_),
    .A(_0015_),
    .X(_0885_));
 sg13g2_nand3_1 _1852_ (.B(_0878_),
    .C(_0885_),
    .A(_0801_),
    .Y(_0886_));
 sg13g2_o21ai_1 _1853_ (.B1(_0886_),
    .Y(_0887_),
    .A1(net216),
    .A2(_0880_));
 sg13g2_nand2b_1 _1854_ (.Y(_0888_),
    .B(_0879_),
    .A_N(net220));
 sg13g2_nor2_1 _1855_ (.A(\color_index[1] ),
    .B(\color_index[0] ),
    .Y(_0889_));
 sg13g2_nand3_1 _1856_ (.B(_0878_),
    .C(_0884_),
    .A(_0801_),
    .Y(_0890_));
 sg13g2_o21ai_1 _1857_ (.B1(_0888_),
    .Y(_0891_),
    .A1(_0889_),
    .A2(_0890_));
 sg13g2_nand2_1 _1858_ (.Y(_0892_),
    .A(_0887_),
    .B(_0891_));
 sg13g2_nand2_1 _1859_ (.Y(_0000_),
    .A(_0883_),
    .B(net217));
 sg13g2_nand2_1 _1860_ (.Y(_0893_),
    .A(_0883_),
    .B(_0887_));
 sg13g2_nand2_1 _1861_ (.Y(_0894_),
    .A(net850),
    .B(_0891_));
 sg13g2_mux2_1 _1862_ (.A0(_0891_),
    .A1(_0894_),
    .S(_0893_),
    .X(_0001_));
 sg13g2_nor2_1 _1863_ (.A(_0887_),
    .B(_0894_),
    .Y(_0895_));
 sg13g2_mux2_1 _1864_ (.A0(_0883_),
    .A1(_0882_),
    .S(_0895_),
    .X(_0002_));
 sg13g2_a21o_1 _1865_ (.A2(_0887_),
    .A1(net850),
    .B1(_0883_),
    .X(_0115_));
 sg13g2_nand2_1 _1866_ (.Y(_0896_),
    .A(_0893_),
    .B(_0115_));
 sg13g2_or2_1 _1867_ (.X(_0003_),
    .B(_0896_),
    .A(_0895_));
 sg13g2_nand2b_2 _1868_ (.Y(_0897_),
    .B(net843),
    .A_N(\pix_x[0] ));
 sg13g2_nor2b_1 _1869_ (.A(net842),
    .B_N(\pix_x[1] ),
    .Y(_0898_));
 sg13g2_xnor2_1 _1870_ (.Y(_0899_),
    .A(net842),
    .B(\pix_x[1] ));
 sg13g2_xnor2_1 _1871_ (.Y(_0900_),
    .A(_0897_),
    .B(_0899_));
 sg13g2_inv_1 _1872_ (.Y(_0901_),
    .A(_0900_));
 sg13g2_xor2_1 _1873_ (.B(\pix_y[6] ),
    .A(\logo_top[6] ),
    .X(_0902_));
 sg13g2_nor2b_1 _1874_ (.A(net818),
    .B_N(net835),
    .Y(_0903_));
 sg13g2_nor2b_1 _1875_ (.A(\logo_top[3] ),
    .B_N(net821),
    .Y(_0904_));
 sg13g2_xnor2_1 _1876_ (.Y(_0905_),
    .A(\logo_top[3] ),
    .B(net821));
 sg13g2_nand2b_1 _1877_ (.Y(_0906_),
    .B(net822),
    .A_N(\logo_top[2] ));
 sg13g2_nor2b_1 _1878_ (.A(net837),
    .B_N(net823),
    .Y(_0907_));
 sg13g2_nand2b_2 _1879_ (.Y(_0908_),
    .B(net838),
    .A_N(net824));
 sg13g2_xnor2_1 _1880_ (.Y(_0909_),
    .A(net837),
    .B(net823));
 sg13g2_a21oi_2 _1881_ (.B1(_0907_),
    .Y(_0910_),
    .A2(_0909_),
    .A1(_0908_));
 sg13g2_xor2_1 _1882_ (.B(net822),
    .A(net836),
    .X(_0911_));
 sg13g2_inv_1 _1883_ (.Y(_0912_),
    .A(_0911_));
 sg13g2_o21ai_1 _1884_ (.B1(_0906_),
    .Y(_0913_),
    .A1(_0910_),
    .A2(_0911_));
 sg13g2_nand2_2 _1885_ (.Y(_0914_),
    .A(_0905_),
    .B(_0913_));
 sg13g2_a21oi_2 _1886_ (.B1(_0904_),
    .Y(_0915_),
    .A2(_0913_),
    .A1(_0905_));
 sg13g2_xor2_1 _1887_ (.B(net819),
    .A(\logo_top[4] ),
    .X(_0916_));
 sg13g2_nor2_1 _1888_ (.A(_0915_),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_a21oi_2 _1889_ (.B1(_0917_),
    .Y(_0918_),
    .A2(net819),
    .A1(_0738_));
 sg13g2_nand2b_1 _1890_ (.Y(_0919_),
    .B(net818),
    .A_N(net835));
 sg13g2_o21ai_1 _1891_ (.B1(_0919_),
    .Y(_0920_),
    .A1(_0903_),
    .A2(_0918_));
 sg13g2_nand2b_1 _1892_ (.Y(_0921_),
    .B(_0920_),
    .A_N(_0902_));
 sg13g2_xnor2_1 _1893_ (.Y(_0922_),
    .A(_0902_),
    .B(_0920_));
 sg13g2_xor2_1 _1894_ (.B(_0920_),
    .A(_0902_),
    .X(_0923_));
 sg13g2_nor2b_1 _1895_ (.A(_0903_),
    .B_N(_0919_),
    .Y(_0924_));
 sg13g2_xnor2_1 _1896_ (.Y(_0925_),
    .A(_0918_),
    .B(_0924_));
 sg13g2_xor2_1 _1897_ (.B(_0924_),
    .A(_0918_),
    .X(_0926_));
 sg13g2_or2_2 _1898_ (.X(_0927_),
    .B(_0913_),
    .A(_0905_));
 sg13g2_and2_1 _1899_ (.A(_0914_),
    .B(_0927_),
    .X(_0928_));
 sg13g2_nand2_1 _1900_ (.Y(_0929_),
    .A(_0914_),
    .B(_0927_));
 sg13g2_xor2_1 _1901_ (.B(_0909_),
    .A(_0908_),
    .X(_0930_));
 sg13g2_xnor2_1 _1902_ (.Y(_0931_),
    .A(_0908_),
    .B(_0909_));
 sg13g2_xnor2_1 _1903_ (.Y(_0932_),
    .A(net838),
    .B(net824));
 sg13g2_xor2_1 _1904_ (.B(net824),
    .A(net838),
    .X(_0933_));
 sg13g2_nor2_1 _1905_ (.A(net786),
    .B(net801),
    .Y(_0934_));
 sg13g2_nand2_2 _1906_ (.Y(_0935_),
    .A(net792),
    .B(net809));
 sg13g2_a21oi_2 _1907_ (.B1(_0898_),
    .Y(_0936_),
    .A2(_0899_),
    .A1(_0897_));
 sg13g2_a21o_1 _1908_ (.A2(_0899_),
    .A1(_0897_),
    .B1(_0898_),
    .X(_0937_));
 sg13g2_nor2b_1 _1909_ (.A(\logo_left[2] ),
    .B_N(\pix_x[2] ),
    .Y(_0938_));
 sg13g2_xnor2_1 _1910_ (.Y(_0939_),
    .A(\logo_left[2] ),
    .B(\pix_x[2] ));
 sg13g2_nor2b_1 _1911_ (.A(\logo_left[3] ),
    .B_N(\pix_x[3] ),
    .Y(_0940_));
 sg13g2_nand2b_1 _1912_ (.Y(_0941_),
    .B(net841),
    .A_N(\pix_x[3] ));
 sg13g2_xnor2_1 _1913_ (.Y(_0942_),
    .A(net841),
    .B(\pix_x[3] ));
 sg13g2_nand2_1 _1914_ (.Y(_0943_),
    .A(_0939_),
    .B(_0942_));
 sg13g2_a21oi_1 _1915_ (.A1(_0938_),
    .A2(_0941_),
    .Y(_0944_),
    .B1(_0940_));
 sg13g2_o21ai_1 _1916_ (.B1(_0944_),
    .Y(_0945_),
    .A1(_0936_),
    .A2(_0943_));
 sg13g2_nor2b_1 _1917_ (.A(\logo_left[4] ),
    .B_N(\pix_x[4] ),
    .Y(_0946_));
 sg13g2_xnor2_1 _1918_ (.Y(_0947_),
    .A(\logo_left[4] ),
    .B(\pix_x[4] ));
 sg13g2_xor2_1 _1919_ (.B(_0947_),
    .A(_0945_),
    .X(_0948_));
 sg13g2_xnor2_1 _1920_ (.Y(_0949_),
    .A(_0945_),
    .B(_0947_));
 sg13g2_a21o_1 _1921_ (.A2(_0947_),
    .A1(_0945_),
    .B1(_0946_),
    .X(_0950_));
 sg13g2_nor2b_1 _1922_ (.A(\logo_left[5] ),
    .B_N(\pix_x[5] ),
    .Y(_0951_));
 sg13g2_nor2_2 _1923_ (.A(_0741_),
    .B(\pix_x[5] ),
    .Y(_0952_));
 sg13g2_inv_1 _1924_ (.Y(_0953_),
    .A(_0952_));
 sg13g2_nor2_1 _1925_ (.A(_0951_),
    .B(_0952_),
    .Y(_0954_));
 sg13g2_xnor2_1 _1926_ (.Y(_0955_),
    .A(_0950_),
    .B(_0954_));
 sg13g2_xor2_1 _1927_ (.B(_0954_),
    .A(_0950_),
    .X(_0956_));
 sg13g2_nor2_2 _1928_ (.A(net772),
    .B(net733),
    .Y(_0957_));
 sg13g2_nand2_1 _1929_ (.Y(_0958_),
    .A(net776),
    .B(net730));
 sg13g2_nand2b_2 _1930_ (.Y(_0959_),
    .B(\logo_left[6] ),
    .A_N(\pix_x[6] ));
 sg13g2_nand2b_2 _1931_ (.Y(_0960_),
    .B(\pix_x[6] ),
    .A_N(\logo_left[6] ));
 sg13g2_and2_1 _1932_ (.A(_0959_),
    .B(_0960_),
    .X(_0961_));
 sg13g2_nand2_1 _1933_ (.Y(_0962_),
    .A(_0959_),
    .B(_0960_));
 sg13g2_a221oi_1 _1934_ (.B2(_0947_),
    .C1(_0946_),
    .B1(_0945_),
    .A1(_0741_),
    .Y(_0963_),
    .A2(\pix_x[5] ));
 sg13g2_nor3_2 _1935_ (.A(_0952_),
    .B(_0962_),
    .C(_0963_),
    .Y(_0964_));
 sg13g2_or3_1 _1936_ (.A(_0952_),
    .B(_0962_),
    .C(_0963_),
    .X(_0965_));
 sg13g2_a221oi_1 _1937_ (.B2(_0960_),
    .C1(_0951_),
    .B1(_0959_),
    .A1(_0950_),
    .Y(_0966_),
    .A2(_0953_));
 sg13g2_o21ai_1 _1938_ (.B1(_0962_),
    .Y(_0967_),
    .A1(_0952_),
    .A2(_0963_));
 sg13g2_o21ai_1 _1939_ (.B1(_0961_),
    .Y(_0968_),
    .A1(_0952_),
    .A2(_0963_));
 sg13g2_or3_1 _1940_ (.A(_0952_),
    .B(_0961_),
    .C(_0963_),
    .X(_0969_));
 sg13g2_nor2_1 _1941_ (.A(_0964_),
    .B(_0966_),
    .Y(_0970_));
 sg13g2_nand2_2 _1942_ (.Y(_0971_),
    .A(net725),
    .B(net723));
 sg13g2_a21oi_2 _1943_ (.B1(net774),
    .Y(_0972_),
    .A2(net724),
    .A1(net727));
 sg13g2_nor2_2 _1944_ (.A(_0957_),
    .B(_0972_),
    .Y(_0973_));
 sg13g2_a21oi_1 _1945_ (.A1(_0937_),
    .A2(_0939_),
    .Y(_0974_),
    .B1(_0938_));
 sg13g2_xnor2_1 _1946_ (.Y(_0975_),
    .A(_0942_),
    .B(_0974_));
 sg13g2_xor2_1 _1947_ (.B(_0974_),
    .A(_0942_),
    .X(_0976_));
 sg13g2_nor2_2 _1948_ (.A(net773),
    .B(net771),
    .Y(_0977_));
 sg13g2_nand2_1 _1949_ (.Y(_0978_),
    .A(net776),
    .B(_0975_));
 sg13g2_nor2_2 _1950_ (.A(net775),
    .B(_0975_),
    .Y(_0979_));
 sg13g2_nand2_1 _1951_ (.Y(_0980_),
    .A(net773),
    .B(net771));
 sg13g2_xnor2_1 _1952_ (.Y(_0981_),
    .A(net772),
    .B(_0975_));
 sg13g2_xnor2_1 _1953_ (.Y(_0982_),
    .A(net775),
    .B(_0975_));
 sg13g2_nand2_2 _1954_ (.Y(_0983_),
    .A(net690),
    .B(net715));
 sg13g2_a21o_1 _1955_ (.A2(_0983_),
    .A1(_0973_),
    .B1(_0935_),
    .X(_0984_));
 sg13g2_nand2b_2 _1956_ (.Y(_0985_),
    .B(_0911_),
    .A_N(_0910_));
 sg13g2_nand2_2 _1957_ (.Y(_0986_),
    .A(_0910_),
    .B(_0912_));
 sg13g2_nand2_1 _1958_ (.Y(_0987_),
    .A(_0985_),
    .B(_0986_));
 sg13g2_and2_1 _1959_ (.A(_0985_),
    .B(_0986_),
    .X(_0988_));
 sg13g2_nor2_2 _1960_ (.A(net790),
    .B(net800),
    .Y(_0989_));
 sg13g2_nand2_2 _1961_ (.Y(_0990_),
    .A(net786),
    .B(net808));
 sg13g2_nor2_1 _1962_ (.A(net773),
    .B(net732),
    .Y(_0991_));
 sg13g2_a22oi_1 _1963_ (.Y(_0992_),
    .B1(net727),
    .B2(net724),
    .A2(net733),
    .A1(net774));
 sg13g2_nor2_2 _1964_ (.A(net715),
    .B(net685),
    .Y(_0993_));
 sg13g2_o21ai_1 _1965_ (.B1(net780),
    .Y(_0994_),
    .A1(net715),
    .A2(net684));
 sg13g2_and2_1 _1966_ (.A(net764),
    .B(_0994_),
    .X(_0995_));
 sg13g2_nor2_1 _1967_ (.A(net786),
    .B(net807),
    .Y(_0996_));
 sg13g2_nand2_2 _1968_ (.Y(_0997_),
    .A(net790),
    .B(net800));
 sg13g2_a22oi_1 _1969_ (.Y(_0998_),
    .B1(net721),
    .B2(net719),
    .A2(net728),
    .A1(net772));
 sg13g2_nor2_1 _1970_ (.A(net728),
    .B(_0977_),
    .Y(_0999_));
 sg13g2_nand2_1 _1971_ (.Y(_1000_),
    .A(net735),
    .B(net718));
 sg13g2_nand2_2 _1972_ (.Y(_1001_),
    .A(net734),
    .B(_0981_));
 sg13g2_nand2_1 _1973_ (.Y(_1002_),
    .A(net682),
    .B(net681));
 sg13g2_a21oi_1 _1974_ (.A1(net682),
    .A2(net681),
    .Y(_1003_),
    .B1(net684));
 sg13g2_nand2b_1 _1975_ (.Y(_1004_),
    .B(net778),
    .A_N(_1003_));
 sg13g2_nor3_2 _1976_ (.A(_0964_),
    .B(_0966_),
    .C(net770),
    .Y(_1005_));
 sg13g2_nand2_1 _1977_ (.Y(_1006_),
    .A(net693),
    .B(_0975_));
 sg13g2_nor2_2 _1978_ (.A(net774),
    .B(net770),
    .Y(_1007_));
 sg13g2_nand2_1 _1979_ (.Y(_1008_),
    .A(net772),
    .B(_0975_));
 sg13g2_nand2_1 _1980_ (.Y(_1009_),
    .A(net690),
    .B(_1007_));
 sg13g2_nor2_2 _1981_ (.A(net790),
    .B(net807),
    .Y(_1010_));
 sg13g2_nand2_1 _1982_ (.Y(_1011_),
    .A(net734),
    .B(net770));
 sg13g2_nand3_1 _1983_ (.B(net733),
    .C(net770),
    .A(net774),
    .Y(_1012_));
 sg13g2_nand3_1 _1984_ (.B(_1010_),
    .C(_1012_),
    .A(_1009_),
    .Y(_1013_));
 sg13g2_nand4_1 _1985_ (.B(_0995_),
    .C(_1004_),
    .A(_0984_),
    .Y(_1014_),
    .D(_1013_));
 sg13g2_a22oi_1 _1986_ (.Y(_1015_),
    .B1(_0981_),
    .B2(net734),
    .A2(net724),
    .A1(net727));
 sg13g2_nand2_1 _1987_ (.Y(_1016_),
    .A(net689),
    .B(net681));
 sg13g2_o21ai_1 _1988_ (.B1(_0981_),
    .Y(_1017_),
    .A1(net734),
    .A2(net690));
 sg13g2_nor2_1 _1989_ (.A(net766),
    .B(_1017_),
    .Y(_1018_));
 sg13g2_o21ai_1 _1990_ (.B1(_1018_),
    .Y(_1019_),
    .A1(_0993_),
    .A2(net777));
 sg13g2_a21o_2 _1991_ (.A2(_1019_),
    .A1(_1014_),
    .B1(net748),
    .X(_1020_));
 sg13g2_xor2_1 _1992_ (.B(_0916_),
    .A(_0915_),
    .X(_1021_));
 sg13g2_xnor2_1 _1993_ (.Y(_1022_),
    .A(_0915_),
    .B(_0916_));
 sg13g2_nor2_2 _1994_ (.A(net786),
    .B(net757),
    .Y(_1023_));
 sg13g2_nand2_2 _1995_ (.Y(_1024_),
    .A(net791),
    .B(net764));
 sg13g2_nor2_2 _1996_ (.A(net733),
    .B(_0979_),
    .Y(_1025_));
 sg13g2_nand2_2 _1997_ (.Y(_1026_),
    .A(net730),
    .B(net716));
 sg13g2_a21oi_1 _1998_ (.A1(net726),
    .A2(net723),
    .Y(_1027_),
    .B1(net731));
 sg13g2_nand4_1 _1999_ (.B(net721),
    .C(net719),
    .A(net737),
    .Y(_1028_),
    .D(_0978_));
 sg13g2_and2_2 _2000_ (.A(_1026_),
    .B(_1028_),
    .X(_1029_));
 sg13g2_nand2_1 _2001_ (.Y(_1030_),
    .A(_1026_),
    .B(_1028_));
 sg13g2_nor2_1 _2002_ (.A(net728),
    .B(_0983_),
    .Y(_1031_));
 sg13g2_nand4_1 _2003_ (.B(net727),
    .C(net724),
    .A(net735),
    .Y(_1032_),
    .D(_0982_));
 sg13g2_o21ai_1 _2004_ (.B1(net704),
    .Y(_1033_),
    .A1(_1030_),
    .A2(_1031_));
 sg13g2_nor2_2 _2005_ (.A(net790),
    .B(net757),
    .Y(_1034_));
 sg13g2_nand2_2 _2006_ (.Y(_1035_),
    .A(net787),
    .B(net768));
 sg13g2_a21oi_2 _2007_ (.B1(_1007_),
    .Y(_1036_),
    .A2(net770),
    .A1(net734));
 sg13g2_mux2_1 _2008_ (.A0(net718),
    .A1(net716),
    .S(net728),
    .X(_1037_));
 sg13g2_nand3_1 _2009_ (.B(net687),
    .C(net677),
    .A(net801),
    .Y(_1038_));
 sg13g2_nand2_2 _2010_ (.Y(_1039_),
    .A(net728),
    .B(_0979_));
 sg13g2_nor2_1 _2011_ (.A(net775),
    .B(net729),
    .Y(_1040_));
 sg13g2_nand2_1 _2012_ (.Y(_1041_),
    .A(net773),
    .B(net738));
 sg13g2_mux2_2 _2013_ (.A0(net773),
    .A1(net717),
    .S(net730),
    .X(_1042_));
 sg13g2_nand2_2 _2014_ (.Y(_1043_),
    .A(_0971_),
    .B(_1042_));
 sg13g2_nand3_1 _2015_ (.B(_1038_),
    .C(net652),
    .A(_1002_),
    .Y(_1044_));
 sg13g2_o21ai_1 _2016_ (.B1(net749),
    .Y(_1045_),
    .A1(net764),
    .A2(_1003_));
 sg13g2_a21oi_2 _2017_ (.B1(_1045_),
    .Y(_1046_),
    .A2(_1044_),
    .A1(_1034_));
 sg13g2_a21oi_1 _2018_ (.A1(_1033_),
    .A2(_1046_),
    .Y(_1047_),
    .B1(net710));
 sg13g2_nor3_2 _2019_ (.A(net737),
    .B(_0964_),
    .C(_0966_),
    .Y(_1048_));
 sg13g2_nand3_1 _2020_ (.B(net725),
    .C(_0967_),
    .A(net730),
    .Y(_1049_));
 sg13g2_nand2_1 _2021_ (.Y(_1050_),
    .A(net775),
    .B(net693));
 sg13g2_a22oi_1 _2022_ (.Y(_1051_),
    .B1(net722),
    .B2(net720),
    .A2(net737),
    .A1(net773));
 sg13g2_a22oi_1 _2023_ (.Y(_1052_),
    .B1(net725),
    .B2(net723),
    .A2(net731),
    .A1(net776));
 sg13g2_or2_1 _2024_ (.X(_1053_),
    .B(_1052_),
    .A(_1051_));
 sg13g2_nor2_1 _2025_ (.A(net735),
    .B(net718),
    .Y(_1054_));
 sg13g2_a22oi_1 _2026_ (.Y(_1055_),
    .B1(_0977_),
    .B2(net730),
    .A2(net723),
    .A1(net725));
 sg13g2_nor3_2 _2027_ (.A(net803),
    .B(_1051_),
    .C(_1055_),
    .Y(_1056_));
 sg13g2_a21oi_2 _2028_ (.B1(net787),
    .Y(_1057_),
    .A2(_1056_),
    .A1(_1006_));
 sg13g2_o21ai_1 _2029_ (.B1(net768),
    .Y(_1058_),
    .A1(_1053_),
    .A2(_1057_));
 sg13g2_a22oi_1 _2030_ (.Y(_1059_),
    .B1(net718),
    .B2(net737),
    .A2(net720),
    .A1(net722));
 sg13g2_a22oi_1 _2031_ (.Y(_1060_),
    .B1(net716),
    .B2(net730),
    .A2(net723),
    .A1(net725));
 sg13g2_nand2_1 _2032_ (.Y(_1061_),
    .A(net689),
    .B(_1026_));
 sg13g2_or2_1 _2033_ (.X(_1062_),
    .B(net670),
    .A(net673));
 sg13g2_nor2_1 _2034_ (.A(net742),
    .B(_1062_),
    .Y(_1063_));
 sg13g2_nor2_1 _2035_ (.A(_0979_),
    .B(_1049_),
    .Y(_1064_));
 sg13g2_nand4_1 _2036_ (.B(net725),
    .C(net723),
    .A(net728),
    .Y(_1065_),
    .D(net716));
 sg13g2_mux2_2 _2037_ (.A0(net775),
    .A1(net718),
    .S(net735),
    .X(_1066_));
 sg13g2_nand2_1 _2038_ (.Y(_1067_),
    .A(_0971_),
    .B(_1066_));
 sg13g2_mux2_2 _2039_ (.A0(_1025_),
    .A1(_1066_),
    .S(net688),
    .X(_1068_));
 sg13g2_xnor2_1 _2040_ (.Y(_1069_),
    .A(net728),
    .B(_0977_));
 sg13g2_nand4_1 _2041_ (.B(net722),
    .C(net720),
    .A(net730),
    .Y(_1070_),
    .D(_0977_));
 sg13g2_nand2_1 _2042_ (.Y(_1071_),
    .A(_1028_),
    .B(_1070_));
 sg13g2_a221oi_1 _2043_ (.B2(net811),
    .C1(_1071_),
    .B1(_1068_),
    .A1(net716),
    .Y(_1072_),
    .A2(_1048_));
 sg13g2_nor2_1 _2044_ (.A(net790),
    .B(net764),
    .Y(_1073_));
 sg13g2_nand2_2 _2045_ (.Y(_1074_),
    .A(net785),
    .B(net759));
 sg13g2_nand2b_1 _2046_ (.Y(_1075_),
    .B(_1032_),
    .A_N(_1068_));
 sg13g2_nand2_1 _2047_ (.Y(_1076_),
    .A(net700),
    .B(_1075_));
 sg13g2_nor2_1 _2048_ (.A(net678),
    .B(net673),
    .Y(_1077_));
 sg13g2_o21ai_1 _2049_ (.B1(net743),
    .Y(_1078_),
    .A1(net761),
    .A2(_1077_));
 sg13g2_a221oi_1 _2050_ (.B2(_1075_),
    .C1(_1078_),
    .B1(net700),
    .A1(net760),
    .Y(_1079_),
    .A2(_1031_));
 sg13g2_o21ai_1 _2051_ (.B1(_1079_),
    .Y(_1080_),
    .A1(net767),
    .A2(_1072_));
 sg13g2_a21oi_1 _2052_ (.A1(_1058_),
    .A2(_1063_),
    .Y(_1081_),
    .B1(net709));
 sg13g2_a22oi_1 _2053_ (.Y(_1082_),
    .B1(_1080_),
    .B2(_1081_),
    .A2(_1047_),
    .A1(_1020_));
 sg13g2_nor4_2 _2054_ (.A(net772),
    .B(_0964_),
    .C(_0966_),
    .Y(_1083_),
    .D(_0975_));
 sg13g2_nand4_1 _2055_ (.B(net727),
    .C(net724),
    .A(net775),
    .Y(_1084_),
    .D(net770));
 sg13g2_nand2_2 _2056_ (.Y(_1085_),
    .A(net735),
    .B(_1007_));
 sg13g2_nand2_1 _2057_ (.Y(_1086_),
    .A(_1084_),
    .B(_1085_));
 sg13g2_a21oi_2 _2058_ (.B1(net690),
    .Y(_1087_),
    .A2(_1011_),
    .A1(_0981_));
 sg13g2_a22oi_1 _2059_ (.Y(_1088_),
    .B1(net722),
    .B2(net720),
    .A2(net731),
    .A1(net776));
 sg13g2_nand2_2 _2060_ (.Y(_1089_),
    .A(_1001_),
    .B(net669));
 sg13g2_nor2b_2 _2061_ (.A(_1087_),
    .B_N(_1089_),
    .Y(_1090_));
 sg13g2_o21ai_1 _2062_ (.B1(net718),
    .Y(_1091_),
    .A1(net774),
    .A2(net734));
 sg13g2_nor2_1 _2063_ (.A(_0979_),
    .B(_1091_),
    .Y(_1092_));
 sg13g2_o21ai_1 _2064_ (.B1(_0981_),
    .Y(_1093_),
    .A1(net774),
    .A2(net733));
 sg13g2_and2_1 _2065_ (.A(net691),
    .B(_1093_),
    .X(_1094_));
 sg13g2_nor3_1 _2066_ (.A(_0935_),
    .B(_1087_),
    .C(_1094_),
    .Y(_1095_));
 sg13g2_a221oi_1 _2067_ (.B2(net785),
    .C1(_1095_),
    .B1(_1090_),
    .A1(net778),
    .Y(_1096_),
    .A2(_1086_));
 sg13g2_a21o_1 _2068_ (.A2(_1094_),
    .A1(_1010_),
    .B1(net759),
    .X(_1097_));
 sg13g2_nor2_2 _2069_ (.A(net786),
    .B(net766),
    .Y(_1098_));
 sg13g2_nand2_2 _2070_ (.Y(_1099_),
    .A(net790),
    .B(net757));
 sg13g2_a22oi_1 _2071_ (.Y(_1100_),
    .B1(_0981_),
    .B2(net729),
    .A2(net724),
    .A1(net727));
 sg13g2_mux2_1 _2072_ (.A0(net775),
    .A1(net715),
    .S(net732),
    .X(_1101_));
 sg13g2_a22oi_1 _2073_ (.Y(_1102_),
    .B1(net665),
    .B2(net675),
    .A2(net669),
    .A1(_1001_));
 sg13g2_a221oi_1 _2074_ (.B2(net699),
    .C1(net751),
    .B1(_1102_),
    .A1(_1090_),
    .Y(_1103_),
    .A2(net695));
 sg13g2_o21ai_1 _2075_ (.B1(_1103_),
    .Y(_1104_),
    .A1(_1096_),
    .A2(_1097_));
 sg13g2_a21o_2 _2076_ (.A2(_1093_),
    .A1(net691),
    .B1(_1015_),
    .X(_1105_));
 sg13g2_mux2_1 _2077_ (.A0(_1017_),
    .A1(_1105_),
    .S(net809),
    .X(_1106_));
 sg13g2_nand2b_1 _2078_ (.Y(_1107_),
    .B(_1034_),
    .A_N(_1106_));
 sg13g2_o21ai_1 _2079_ (.B1(net750),
    .Y(_1108_),
    .A1(_1017_),
    .A2(_1024_));
 sg13g2_a21oi_1 _2080_ (.A1(net759),
    .A2(_1086_),
    .Y(_1109_),
    .B1(_1108_));
 sg13g2_a21oi_1 _2081_ (.A1(_1107_),
    .A2(_1109_),
    .Y(_1110_),
    .B1(net706));
 sg13g2_nor4_2 _2082_ (.A(net735),
    .B(_0964_),
    .C(_0966_),
    .Y(_1111_),
    .D(net715));
 sg13g2_nor2_2 _2083_ (.A(net731),
    .B(net717),
    .Y(_1112_));
 sg13g2_nand2_1 _2084_ (.Y(_1113_),
    .A(net733),
    .B(_0979_));
 sg13g2_a21o_2 _2085_ (.A2(net663),
    .A1(net672),
    .B1(_1111_),
    .X(_1114_));
 sg13g2_a22oi_1 _2086_ (.Y(_1115_),
    .B1(_0981_),
    .B2(net729),
    .A2(net719),
    .A1(net721));
 sg13g2_o21ai_1 _2087_ (.B1(net693),
    .Y(_1116_),
    .A1(net736),
    .A2(net715));
 sg13g2_a21oi_1 _2088_ (.A1(net686),
    .A2(_1039_),
    .Y(_1117_),
    .B1(_1115_));
 sg13g2_nand2_1 _2089_ (.Y(_1118_),
    .A(net652),
    .B(_1116_));
 sg13g2_a221oi_1 _2090_ (.B2(net652),
    .C1(net751),
    .B1(_1116_),
    .A1(net699),
    .Y(_1119_),
    .A2(_1114_));
 sg13g2_nand2_1 _2091_ (.Y(_1120_),
    .A(net785),
    .B(_1111_));
 sg13g2_nor2_2 _2092_ (.A(net741),
    .B(net765),
    .Y(_1121_));
 sg13g2_nand2_2 _2093_ (.Y(_1122_),
    .A(net750),
    .B(net759));
 sg13g2_a22oi_1 _2094_ (.Y(_1123_),
    .B1(_1007_),
    .B2(net728),
    .A2(net719),
    .A1(net721));
 sg13g2_o21ai_1 _2095_ (.B1(net691),
    .Y(_1124_),
    .A1(net736),
    .A2(_1008_));
 sg13g2_a21oi_1 _2096_ (.A1(net652),
    .A2(_1124_),
    .Y(_1125_),
    .B1(_1122_));
 sg13g2_nor2_1 _2097_ (.A(net745),
    .B(net762),
    .Y(_1126_));
 sg13g2_nand2_2 _2098_ (.Y(_1127_),
    .A(net750),
    .B(net765));
 sg13g2_a221oi_1 _2099_ (.B2(_1102_),
    .C1(_1119_),
    .B1(net662),
    .A1(_1120_),
    .Y(_1128_),
    .A2(_1125_));
 sg13g2_o21ai_1 _2100_ (.B1(net654),
    .Y(_1129_),
    .A1(net711),
    .A2(_1128_));
 sg13g2_a21o_1 _2101_ (.A2(_1110_),
    .A1(_1104_),
    .B1(_1129_),
    .X(_1130_));
 sg13g2_o21ai_1 _2102_ (.B1(_1130_),
    .Y(_1131_),
    .A1(net653),
    .A2(_1082_));
 sg13g2_xnor2_1 _2103_ (.Y(_1132_),
    .A(net843),
    .B(\pix_x[0] ));
 sg13g2_xor2_1 _2104_ (.B(\pix_x[0] ),
    .A(net843),
    .X(_1133_));
 sg13g2_or3_1 _2105_ (.A(net810),
    .B(_1051_),
    .C(_1055_),
    .X(_1134_));
 sg13g2_and2_1 _2106_ (.A(_1005_),
    .B(net700),
    .X(_1135_));
 sg13g2_a21o_1 _2107_ (.A2(_1134_),
    .A1(net700),
    .B1(_1135_),
    .X(_1136_));
 sg13g2_inv_1 _2108_ (.Y(_1137_),
    .A(_1136_));
 sg13g2_a221oi_1 _2109_ (.B2(_1134_),
    .C1(_1135_),
    .B1(net700),
    .A1(net762),
    .Y(_1138_),
    .A2(_1053_));
 sg13g2_nand2_1 _2110_ (.Y(_1139_),
    .A(net777),
    .B(_1062_));
 sg13g2_nand4_1 _2111_ (.B(_1061_),
    .C(_1138_),
    .A(_1049_),
    .Y(_1140_),
    .D(_1139_));
 sg13g2_nor2_1 _2112_ (.A(net678),
    .B(_1048_),
    .Y(_1141_));
 sg13g2_mux2_2 _2113_ (.A0(_1042_),
    .A1(_1066_),
    .S(net688),
    .X(_1142_));
 sg13g2_a22oi_1 _2114_ (.Y(_1143_),
    .B1(net717),
    .B2(net737),
    .A2(net720),
    .A1(net722));
 sg13g2_a221oi_1 _2115_ (.B2(_1039_),
    .C1(_1071_),
    .B1(_1143_),
    .A1(net803),
    .Y(_1144_),
    .A2(_1142_));
 sg13g2_nand2_2 _2116_ (.Y(_1145_),
    .A(net692),
    .B(_0999_));
 sg13g2_nand2_1 _2117_ (.Y(_1146_),
    .A(net692),
    .B(net677));
 sg13g2_and2_1 _2118_ (.A(net692),
    .B(net677),
    .X(_1147_));
 sg13g2_a221oi_1 _2119_ (.B2(net778),
    .C1(_0988_),
    .B1(_1147_),
    .A1(net791),
    .Y(_1148_),
    .A2(_1142_));
 sg13g2_a221oi_1 _2120_ (.B2(_1148_),
    .C1(net743),
    .B1(_1144_),
    .A1(net760),
    .Y(_1149_),
    .A2(_1141_));
 sg13g2_a21o_1 _2121_ (.A2(_1140_),
    .A1(net743),
    .B1(_1149_),
    .X(_1150_));
 sg13g2_or2_1 _2122_ (.X(_1151_),
    .B(net667),
    .A(net671));
 sg13g2_o21ai_1 _2123_ (.B1(_1000_),
    .Y(_1152_),
    .A1(net672),
    .A2(net669));
 sg13g2_nand2_1 _2124_ (.Y(_1153_),
    .A(net808),
    .B(_1152_));
 sg13g2_or2_2 _2125_ (.X(_1154_),
    .B(net683),
    .A(net684));
 sg13g2_nand3_1 _2126_ (.B(_1039_),
    .C(_1154_),
    .A(net801),
    .Y(_1155_));
 sg13g2_a21o_1 _2127_ (.A2(_1155_),
    .A1(_1153_),
    .B1(_1099_),
    .X(_1156_));
 sg13g2_a22oi_1 _2128_ (.Y(_1157_),
    .B1(_1154_),
    .B2(net766),
    .A2(net698),
    .A1(net677));
 sg13g2_nand3_1 _2129_ (.B(_1156_),
    .C(_1157_),
    .A(net739),
    .Y(_1158_));
 sg13g2_and4_2 _2130_ (.A(net772),
    .B(net735),
    .C(net721),
    .D(net719),
    .X(_1159_));
 sg13g2_a21oi_2 _2131_ (.B1(_1159_),
    .Y(_1160_),
    .A2(_1115_),
    .A1(net675));
 sg13g2_nor2_1 _2132_ (.A(net760),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_o21ai_1 _2133_ (.B1(_1161_),
    .Y(_1162_),
    .A1(net780),
    .A2(_1085_));
 sg13g2_o21ai_1 _2134_ (.B1(net808),
    .Y(_1163_),
    .A1(net684),
    .A2(_1123_));
 sg13g2_nand2_1 _2135_ (.Y(_1164_),
    .A(_1160_),
    .B(_1163_));
 sg13g2_nand2_2 _2136_ (.Y(_1165_),
    .A(net754),
    .B(net697));
 sg13g2_a221oi_1 _2137_ (.B2(net695),
    .C1(net740),
    .B1(_1164_),
    .A1(net698),
    .Y(_1166_),
    .A2(_1154_));
 sg13g2_a21oi_1 _2138_ (.A1(_1162_),
    .A2(_1166_),
    .Y(_1167_),
    .B1(net705));
 sg13g2_a221oi_1 _2139_ (.B2(_1167_),
    .C1(net655),
    .B1(_1158_),
    .A1(net705),
    .Y(_1168_),
    .A2(_1150_));
 sg13g2_and4_2 _2140_ (.A(net737),
    .B(net722),
    .C(net720),
    .D(_0979_),
    .X(_1169_));
 sg13g2_nand4_1 _2141_ (.B(net721),
    .C(net719),
    .A(net735),
    .Y(_1170_),
    .D(_0979_));
 sg13g2_nor2_1 _2142_ (.A(_1005_),
    .B(net667),
    .Y(_1171_));
 sg13g2_o21ai_1 _2143_ (.B1(net676),
    .Y(_1172_),
    .A1(_1005_),
    .A2(net667));
 sg13g2_nand2_2 _2144_ (.Y(_1173_),
    .A(_1170_),
    .B(_1172_));
 sg13g2_nand2_1 _2145_ (.Y(_1174_),
    .A(net758),
    .B(net777));
 sg13g2_nor2_2 _2146_ (.A(net764),
    .B(net778),
    .Y(_1175_));
 sg13g2_o21ai_1 _2147_ (.B1(_1175_),
    .Y(_1176_),
    .A1(net788),
    .A2(_1007_));
 sg13g2_nand2_1 _2148_ (.Y(_1177_),
    .A(net789),
    .B(_1085_));
 sg13g2_o21ai_1 _2149_ (.B1(net739),
    .Y(_1178_),
    .A1(_1160_),
    .A2(_1177_));
 sg13g2_a21oi_1 _2150_ (.A1(_1173_),
    .A2(_1176_),
    .Y(_1179_),
    .B1(_1178_));
 sg13g2_a21oi_2 _2151_ (.B1(_1169_),
    .Y(_1180_),
    .A2(net667),
    .A1(net676));
 sg13g2_nor2_2 _2152_ (.A(net761),
    .B(net780),
    .Y(_1181_));
 sg13g2_o21ai_1 _2153_ (.B1(_1181_),
    .Y(_1182_),
    .A1(net668),
    .A2(net666));
 sg13g2_nand3_1 _2154_ (.B(_1180_),
    .C(_1182_),
    .A(net754),
    .Y(_1183_));
 sg13g2_nand3_1 _2155_ (.B(net812),
    .C(net763),
    .A(net754),
    .Y(_1184_));
 sg13g2_a22oi_1 _2156_ (.Y(_1185_),
    .B1(_1183_),
    .B2(_1184_),
    .A2(_1175_),
    .A1(_1173_));
 sg13g2_or3_1 _2157_ (.A(net714),
    .B(_1179_),
    .C(_1185_),
    .X(_1186_));
 sg13g2_a22oi_1 _2158_ (.Y(_1187_),
    .B1(_0977_),
    .B2(net731),
    .A2(net719),
    .A1(net721));
 sg13g2_a21o_1 _2159_ (.A2(net666),
    .A1(net676),
    .B1(net660),
    .X(_1188_));
 sg13g2_a221oi_1 _2160_ (.B2(net702),
    .C1(net744),
    .B1(_1188_),
    .A1(_1043_),
    .Y(_1189_),
    .A2(_1116_));
 sg13g2_a22oi_1 _2161_ (.Y(_1190_),
    .B1(_1181_),
    .B2(_1114_),
    .A2(_1117_),
    .A1(_1034_));
 sg13g2_o21ai_1 _2162_ (.B1(_1190_),
    .Y(_1191_),
    .A1(net661),
    .A2(_1189_));
 sg13g2_a21o_2 _2163_ (.A2(net665),
    .A1(net675),
    .B1(net669),
    .X(_1192_));
 sg13g2_a21oi_1 _2164_ (.A1(net701),
    .A2(net665),
    .Y(_1193_),
    .B1(_1192_));
 sg13g2_a21oi_1 _2165_ (.A1(net704),
    .A2(net660),
    .Y(_1194_),
    .B1(net755));
 sg13g2_a21oi_1 _2166_ (.A1(_1193_),
    .A2(_1194_),
    .Y(_1195_),
    .B1(net707));
 sg13g2_a21oi_1 _2167_ (.A1(_1191_),
    .A2(_1195_),
    .Y(_1196_),
    .B1(net653));
 sg13g2_a21o_1 _2168_ (.A2(_1196_),
    .A1(_1186_),
    .B1(net650),
    .X(_1197_));
 sg13g2_o21ai_1 _2169_ (.B1(_1133_),
    .Y(_1198_),
    .A1(_1168_),
    .A2(_1197_));
 sg13g2_a21o_1 _2170_ (.A2(_1131_),
    .A1(net650),
    .B1(_1198_),
    .X(_1199_));
 sg13g2_o21ai_1 _2171_ (.B1(net787),
    .Y(_1200_),
    .A1(net811),
    .A2(_1142_));
 sg13g2_a22oi_1 _2172_ (.Y(_1201_),
    .B1(net718),
    .B2(net730),
    .A2(net723),
    .A1(net725));
 sg13g2_a221oi_1 _2173_ (.B2(_1039_),
    .C1(_1201_),
    .B1(_1143_),
    .A1(net803),
    .Y(_1202_),
    .A2(_1142_));
 sg13g2_o21ai_1 _2174_ (.B1(_1148_),
    .Y(_1203_),
    .A1(_1200_),
    .A2(_1202_));
 sg13g2_o21ai_1 _2175_ (.B1(_0997_),
    .Y(_1204_),
    .A1(net679),
    .A2(_1048_));
 sg13g2_nor3_2 _2176_ (.A(net767),
    .B(net678),
    .C(_1064_),
    .Y(_1205_));
 sg13g2_nand2_1 _2177_ (.Y(_1206_),
    .A(_1204_),
    .B(_1205_));
 sg13g2_a21oi_1 _2178_ (.A1(_1203_),
    .A2(_1206_),
    .Y(_1207_),
    .B1(net743));
 sg13g2_a21oi_1 _2179_ (.A1(net810),
    .A2(_1062_),
    .Y(_1208_),
    .B1(net752));
 sg13g2_nand2_1 _2180_ (.Y(_1209_),
    .A(_1138_),
    .B(_1208_));
 sg13g2_o21ai_1 _2181_ (.B1(_0989_),
    .Y(_1210_),
    .A1(_1052_),
    .A2(net674));
 sg13g2_o21ai_1 _2182_ (.B1(_1010_),
    .Y(_1211_),
    .A1(net673),
    .A2(net670));
 sg13g2_nand4_1 _2183_ (.B(_1061_),
    .C(_1210_),
    .A(_1049_),
    .Y(_1212_),
    .D(_1211_));
 sg13g2_o21ai_1 _2184_ (.B1(net709),
    .Y(_1213_),
    .A1(_1209_),
    .A2(_1212_));
 sg13g2_a21o_1 _2185_ (.A2(net677),
    .A1(net687),
    .B1(net683),
    .X(_1214_));
 sg13g2_mux2_1 _2186_ (.A0(_1152_),
    .A1(_1214_),
    .S(net802),
    .X(_1215_));
 sg13g2_and2_1 _2187_ (.A(net807),
    .B(_1037_),
    .X(_1216_));
 sg13g2_a21o_1 _2188_ (.A2(_1152_),
    .A1(net800),
    .B1(_1216_),
    .X(_1217_));
 sg13g2_and2_1 _2189_ (.A(_1154_),
    .B(_1181_),
    .X(_1218_));
 sg13g2_a221oi_1 _2190_ (.B2(net687),
    .C1(net683),
    .B1(_1042_),
    .A1(_0990_),
    .Y(_1219_),
    .A2(net684));
 sg13g2_o21ai_1 _2191_ (.B1(net739),
    .Y(_1220_),
    .A1(net758),
    .A2(_1219_));
 sg13g2_a221oi_1 _2192_ (.B2(net698),
    .C1(_1220_),
    .B1(_1217_),
    .A1(net695),
    .Y(_1221_),
    .A2(_1215_));
 sg13g2_or2_1 _2193_ (.X(_1222_),
    .B(_1115_),
    .A(net686));
 sg13g2_o21ai_1 _2194_ (.B1(net808),
    .Y(_1223_),
    .A1(net686),
    .A2(_1115_));
 sg13g2_a21oi_1 _2195_ (.A1(_1160_),
    .A2(_1223_),
    .Y(_1224_),
    .B1(_1099_));
 sg13g2_nor2_1 _2196_ (.A(net740),
    .B(_1224_),
    .Y(_1225_));
 sg13g2_o21ai_1 _2197_ (.B1(net807),
    .Y(_1226_),
    .A1(net684),
    .A2(net682));
 sg13g2_o21ai_1 _2198_ (.B1(net801),
    .Y(_1227_),
    .A1(net684),
    .A2(_1123_));
 sg13g2_a21oi_1 _2199_ (.A1(_1226_),
    .A2(_1227_),
    .Y(_1228_),
    .B1(net696));
 sg13g2_nor2_1 _2200_ (.A(net786),
    .B(_1085_),
    .Y(_1229_));
 sg13g2_nor3_1 _2201_ (.A(net760),
    .B(_1160_),
    .C(_1229_),
    .Y(_1230_));
 sg13g2_nor4_1 _2202_ (.A(net740),
    .B(_1224_),
    .C(_1228_),
    .D(_1230_),
    .Y(_1231_));
 sg13g2_or3_1 _2203_ (.A(net705),
    .B(_1221_),
    .C(_1231_),
    .X(_1232_));
 sg13g2_o21ai_1 _2204_ (.B1(_1232_),
    .Y(_1233_),
    .A1(_1207_),
    .A2(_1213_));
 sg13g2_nor2_2 _2205_ (.A(net767),
    .B(_0990_),
    .Y(_1234_));
 sg13g2_a22oi_1 _2206_ (.Y(_1235_),
    .B1(_1234_),
    .B2(_1007_),
    .A2(_1172_),
    .A1(_1170_));
 sg13g2_o21ai_1 _2207_ (.B1(_1183_),
    .Y(_1236_),
    .A1(net754),
    .A2(_1235_));
 sg13g2_nor3_1 _2208_ (.A(net697),
    .B(net668),
    .C(net665),
    .Y(_1237_));
 sg13g2_a221oi_1 _2209_ (.B2(net666),
    .C1(net659),
    .B1(net675),
    .A1(net788),
    .Y(_1238_),
    .A2(net761));
 sg13g2_o21ai_1 _2210_ (.B1(net745),
    .Y(_1239_),
    .A1(_1237_),
    .A2(_1238_));
 sg13g2_nand3b_1 _2211_ (.B(_1239_),
    .C(net713),
    .Y(_1240_),
    .A_N(_1189_));
 sg13g2_o21ai_1 _2212_ (.B1(_1240_),
    .Y(_1241_),
    .A1(net713),
    .A2(_1236_));
 sg13g2_a21o_1 _2213_ (.A2(_1241_),
    .A1(net657),
    .B1(net650),
    .X(_1242_));
 sg13g2_a21oi_1 _2214_ (.A1(net653),
    .A2(_1233_),
    .Y(_1243_),
    .B1(_1242_));
 sg13g2_a21oi_2 _2215_ (.B1(net685),
    .Y(_1244_),
    .A2(net715),
    .A1(net690));
 sg13g2_or2_1 _2216_ (.X(_1245_),
    .B(_1244_),
    .A(net791));
 sg13g2_nand4_1 _2217_ (.B(_0995_),
    .C(_1004_),
    .A(_0984_),
    .Y(_1246_),
    .D(_1245_));
 sg13g2_a221oi_1 _2218_ (.B2(net792),
    .C1(net715),
    .B1(net685),
    .A1(net729),
    .Y(_1247_),
    .A2(net688));
 sg13g2_nand2_1 _2219_ (.Y(_1248_),
    .A(net759),
    .B(_1247_));
 sg13g2_a21o_1 _2220_ (.A2(_1248_),
    .A1(_1246_),
    .B1(net748),
    .X(_1249_));
 sg13g2_o21ai_1 _2221_ (.B1(net749),
    .Y(_1250_),
    .A1(_1003_),
    .A2(_1174_));
 sg13g2_nor2_2 _2222_ (.A(net763),
    .B(_0997_),
    .Y(_1251_));
 sg13g2_nand2_2 _2223_ (.Y(_1252_),
    .A(net764),
    .B(net778));
 sg13g2_a21oi_1 _2224_ (.A1(_1029_),
    .A2(_1032_),
    .Y(_1253_),
    .B1(_1252_));
 sg13g2_a22oi_1 _2225_ (.Y(_1254_),
    .B1(net677),
    .B2(net687),
    .A2(net681),
    .A1(net682));
 sg13g2_nor3_1 _2226_ (.A(net757),
    .B(net778),
    .C(_1254_),
    .Y(_1255_));
 sg13g2_a21oi_1 _2227_ (.A1(_1002_),
    .A2(net652),
    .Y(_1256_),
    .B1(net764));
 sg13g2_nor4_1 _2228_ (.A(_1250_),
    .B(_1253_),
    .C(_1255_),
    .D(_1256_),
    .Y(_1257_));
 sg13g2_nor2_1 _2229_ (.A(net710),
    .B(_1257_),
    .Y(_1258_));
 sg13g2_o21ai_1 _2230_ (.B1(net779),
    .Y(_1259_),
    .A1(_1052_),
    .A2(net673));
 sg13g2_and2_1 _2231_ (.A(_1063_),
    .B(_1259_),
    .X(_1260_));
 sg13g2_nand3b_1 _2232_ (.B(_1065_),
    .C(_1032_),
    .Y(_1261_),
    .A_N(_1201_));
 sg13g2_nor2_1 _2233_ (.A(net767),
    .B(net777),
    .Y(_1262_));
 sg13g2_nand2_2 _2234_ (.Y(_1263_),
    .A(net757),
    .B(net778));
 sg13g2_nand3_1 _2235_ (.B(_0979_),
    .C(_0989_),
    .A(net743),
    .Y(_1264_));
 sg13g2_o21ai_1 _2236_ (.B1(_1078_),
    .Y(_1265_),
    .A1(net678),
    .A2(_1264_));
 sg13g2_a22oi_1 _2237_ (.Y(_1266_),
    .B1(_1261_),
    .B2(_1262_),
    .A2(_1175_),
    .A1(_1075_));
 sg13g2_a221oi_1 _2238_ (.B2(_1266_),
    .C1(net709),
    .B1(_1265_),
    .A1(_1058_),
    .Y(_1267_),
    .A2(_1260_));
 sg13g2_a21o_1 _2239_ (.A2(_1258_),
    .A1(_1249_),
    .B1(_1267_),
    .X(_1268_));
 sg13g2_nand2_1 _2240_ (.Y(_1269_),
    .A(net695),
    .B(_1105_));
 sg13g2_a22oi_1 _2241_ (.Y(_1270_),
    .B1(_1007_),
    .B2(net734),
    .A2(net724),
    .A1(net727));
 sg13g2_nand2_1 _2242_ (.Y(_1271_),
    .A(_1251_),
    .B(_1270_));
 sg13g2_nand3_1 _2243_ (.B(net729),
    .C(_1034_),
    .A(net772),
    .Y(_1272_));
 sg13g2_nand3_1 _2244_ (.B(_1084_),
    .C(_1085_),
    .A(net699),
    .Y(_1273_));
 sg13g2_nand4_1 _2245_ (.B(_1269_),
    .C(_1272_),
    .A(net750),
    .Y(_1274_),
    .D(_1273_));
 sg13g2_a21oi_1 _2246_ (.A1(net765),
    .A2(_1106_),
    .Y(_1275_),
    .B1(_1274_));
 sg13g2_and3_1 _2247_ (.X(_1276_),
    .A(net741),
    .B(_1090_),
    .C(_1271_));
 sg13g2_o21ai_1 _2248_ (.B1(net711),
    .Y(_1277_),
    .A1(_1275_),
    .A2(_1276_));
 sg13g2_nand2_1 _2249_ (.Y(_1278_),
    .A(_1118_),
    .B(_1127_));
 sg13g2_o21ai_1 _2250_ (.B1(net662),
    .Y(_1279_),
    .A1(_0935_),
    .A2(_1102_));
 sg13g2_a22oi_1 _2251_ (.Y(_1280_),
    .B1(net660),
    .B2(net681),
    .A2(net665),
    .A1(net675));
 sg13g2_or2_1 _2252_ (.X(_1281_),
    .B(_1280_),
    .A(net793));
 sg13g2_o21ai_1 _2253_ (.B1(_1281_),
    .Y(_1282_),
    .A1(net777),
    .A2(_1090_));
 sg13g2_o21ai_1 _2254_ (.B1(_1278_),
    .Y(_1283_),
    .A1(_1279_),
    .A2(_1282_));
 sg13g2_a21oi_1 _2255_ (.A1(net706),
    .A2(_1283_),
    .Y(_1284_),
    .B1(net655));
 sg13g2_a221oi_1 _2256_ (.B2(_1284_),
    .C1(_0923_),
    .B1(_1277_),
    .A1(net655),
    .Y(_1285_),
    .A2(_1268_));
 sg13g2_o21ai_1 _2257_ (.B1(_1132_),
    .Y(_1286_),
    .A1(_1243_),
    .A2(_1285_));
 sg13g2_a21o_1 _2258_ (.A2(_1286_),
    .A1(_1199_),
    .B1(_0900_),
    .X(_1287_));
 sg13g2_xnor2_1 _2259_ (.Y(_1288_),
    .A(_0936_),
    .B(_0939_));
 sg13g2_o21ai_1 _2260_ (.B1(net803),
    .Y(_1289_),
    .A1(net679),
    .A2(_1048_));
 sg13g2_o21ai_1 _2261_ (.B1(net810),
    .Y(_1290_),
    .A1(_1048_),
    .A2(net670));
 sg13g2_a21oi_1 _2262_ (.A1(_1289_),
    .A2(_1290_),
    .Y(_1291_),
    .B1(net794));
 sg13g2_nand2b_1 _2263_ (.Y(_1292_),
    .B(_1205_),
    .A_N(_1291_));
 sg13g2_a21oi_1 _2264_ (.A1(net693),
    .A2(_1042_),
    .Y(_1293_),
    .B1(_1201_));
 sg13g2_nor2_1 _2265_ (.A(net795),
    .B(_1293_),
    .Y(_1294_));
 sg13g2_nand2b_1 _2266_ (.Y(_1295_),
    .B(_1148_),
    .A_N(_1294_));
 sg13g2_nand3_1 _2267_ (.B(_1292_),
    .C(_1295_),
    .A(net752),
    .Y(_1296_));
 sg13g2_nor3_1 _2268_ (.A(net810),
    .B(_1052_),
    .C(net673),
    .Y(_1297_));
 sg13g2_nor3_1 _2269_ (.A(net768),
    .B(_1056_),
    .C(_1297_),
    .Y(_1298_));
 sg13g2_nor2_1 _2270_ (.A(_1212_),
    .B(_1298_),
    .Y(_1299_));
 sg13g2_or3_1 _2271_ (.A(_1136_),
    .B(_1212_),
    .C(_1298_),
    .X(_1300_));
 sg13g2_a21oi_1 _2272_ (.A1(net742),
    .A2(_1300_),
    .Y(_1301_),
    .B1(net712));
 sg13g2_a21o_1 _2273_ (.A2(_1152_),
    .A1(net801),
    .B1(_1066_),
    .X(_1302_));
 sg13g2_a221oi_1 _2274_ (.B2(net698),
    .C1(net749),
    .B1(_1302_),
    .A1(net695),
    .Y(_1303_),
    .A2(_1214_));
 sg13g2_nor2_1 _2275_ (.A(net758),
    .B(_0990_),
    .Y(_1304_));
 sg13g2_a21oi_1 _2276_ (.A1(_1214_),
    .A2(_1304_),
    .Y(_1305_),
    .B1(_1218_));
 sg13g2_o21ai_1 _2277_ (.B1(net801),
    .Y(_1306_),
    .A1(net686),
    .A2(_1115_));
 sg13g2_a21oi_1 _2278_ (.A1(_1163_),
    .A2(_1306_),
    .Y(_1307_),
    .B1(net696));
 sg13g2_nor4_1 _2279_ (.A(net740),
    .B(_1161_),
    .C(_1224_),
    .D(_1307_),
    .Y(_1308_));
 sg13g2_a21o_1 _2280_ (.A2(_1305_),
    .A1(_1303_),
    .B1(_1308_),
    .X(_1309_));
 sg13g2_a221oi_1 _2281_ (.B2(net712),
    .C1(net656),
    .B1(_1309_),
    .A1(_1296_),
    .Y(_1310_),
    .A2(_1301_));
 sg13g2_o21ai_1 _2282_ (.B1(net754),
    .Y(_1311_),
    .A1(net769),
    .A2(_1180_));
 sg13g2_a221oi_1 _2283_ (.B2(_1251_),
    .C1(_1311_),
    .B1(net659),
    .A1(_1151_),
    .Y(_1312_),
    .A2(_1181_));
 sg13g2_nor4_2 _2284_ (.A(net737),
    .B(_0964_),
    .C(_0966_),
    .Y(_1313_),
    .D(net770));
 sg13g2_nand2_1 _2285_ (.Y(_1314_),
    .A(net745),
    .B(_1180_));
 sg13g2_a221oi_1 _2286_ (.B2(net762),
    .C1(_1314_),
    .B1(_1313_),
    .A1(net788),
    .Y(_1315_),
    .A2(_1173_));
 sg13g2_o21ai_1 _2287_ (.B1(net708),
    .Y(_1316_),
    .A1(_1035_),
    .A2(_1180_));
 sg13g2_inv_1 _2288_ (.Y(_1317_),
    .A(_1316_));
 sg13g2_o21ai_1 _2289_ (.B1(_1317_),
    .Y(_1318_),
    .A1(_1312_),
    .A2(_1315_));
 sg13g2_nand2b_1 _2290_ (.Y(_1319_),
    .B(_1042_),
    .A_N(net659));
 sg13g2_a221oi_1 _2291_ (.B2(net701),
    .C1(net744),
    .B1(_1319_),
    .A1(_1043_),
    .Y(_1320_),
    .A2(_1116_));
 sg13g2_a221oi_1 _2292_ (.B2(net723),
    .C1(_1007_),
    .B1(net725),
    .A1(net776),
    .Y(_1321_),
    .A2(net732));
 sg13g2_or2_1 _2293_ (.X(_1322_),
    .B(_1321_),
    .A(net659));
 sg13g2_o21ai_1 _2294_ (.B1(_1098_),
    .Y(_1323_),
    .A1(net659),
    .A2(_1321_));
 sg13g2_o21ai_1 _2295_ (.B1(net701),
    .Y(_1324_),
    .A1(net671),
    .A2(net659));
 sg13g2_nand3_1 _2296_ (.B(_1323_),
    .C(_1324_),
    .A(net744),
    .Y(_1325_));
 sg13g2_a221oi_1 _2297_ (.B2(net777),
    .C1(_1325_),
    .B1(_1322_),
    .A1(net805),
    .Y(_1326_),
    .A2(_1319_));
 sg13g2_o21ai_1 _2298_ (.B1(net713),
    .Y(_1327_),
    .A1(_1320_),
    .A2(_1326_));
 sg13g2_and3_1 _2299_ (.X(_1328_),
    .A(net656),
    .B(_1318_),
    .C(_1327_));
 sg13g2_nor3_1 _2300_ (.A(_0922_),
    .B(_1310_),
    .C(_1328_),
    .Y(_1329_));
 sg13g2_o21ai_1 _2301_ (.B1(net810),
    .Y(_1330_),
    .A1(net679),
    .A2(net674));
 sg13g2_o21ai_1 _2302_ (.B1(net803),
    .Y(_1331_),
    .A1(net674),
    .A2(net670));
 sg13g2_and2_1 _2303_ (.A(_1330_),
    .B(_1331_),
    .X(_1332_));
 sg13g2_a21oi_1 _2304_ (.A1(_1330_),
    .A2(_1331_),
    .Y(_1333_),
    .B1(_1024_));
 sg13g2_a221oi_1 _2305_ (.B2(net811),
    .C1(net679),
    .B1(_1112_),
    .A1(net717),
    .Y(_1334_),
    .A2(net673));
 sg13g2_nor2_2 _2306_ (.A(_1035_),
    .B(_1334_),
    .Y(_1335_));
 sg13g2_a21o_1 _2307_ (.A2(_1261_),
    .A1(net695),
    .B1(net753),
    .X(_1336_));
 sg13g2_nor3_1 _2308_ (.A(_1333_),
    .B(_1335_),
    .C(_1336_),
    .Y(_1337_));
 sg13g2_a21oi_1 _2309_ (.A1(_1076_),
    .A2(_1337_),
    .Y(_1338_),
    .B1(_1260_));
 sg13g2_mux4_1 _2310_ (.S0(net692),
    .A0(_0957_),
    .A1(_0999_),
    .A2(_1054_),
    .A3(_1040_),
    .S1(net802),
    .X(_1339_));
 sg13g2_o21ai_1 _2311_ (.B1(_1339_),
    .Y(_1340_),
    .A1(net787),
    .A2(_1056_));
 sg13g2_nand2b_1 _2312_ (.Y(_1341_),
    .B(_1339_),
    .A_N(_1057_));
 sg13g2_a21oi_1 _2313_ (.A1(net661),
    .A2(_1341_),
    .Y(_1342_),
    .B1(net709));
 sg13g2_nand2b_1 _2314_ (.Y(_1343_),
    .B(_1342_),
    .A_N(_1338_));
 sg13g2_nor2_1 _2315_ (.A(_1099_),
    .B(_1254_),
    .Y(_1344_));
 sg13g2_nor2_1 _2316_ (.A(_1254_),
    .B(_1263_),
    .Y(_1345_));
 sg13g2_a22oi_1 _2317_ (.Y(_1346_),
    .B1(_1066_),
    .B2(net688),
    .A2(_1001_),
    .A1(net683));
 sg13g2_nor2_1 _2318_ (.A(net758),
    .B(_1346_),
    .Y(_1347_));
 sg13g2_nor4_1 _2319_ (.A(_1250_),
    .B(_1255_),
    .C(_1345_),
    .D(_1347_),
    .Y(_1348_));
 sg13g2_a21oi_1 _2320_ (.A1(_0973_),
    .A2(_0983_),
    .Y(_1349_),
    .B1(_1252_));
 sg13g2_nor2_2 _2321_ (.A(net702),
    .B(_1251_),
    .Y(_1350_));
 sg13g2_nor2b_1 _2322_ (.A(_1244_),
    .B_N(_1350_),
    .Y(_1351_));
 sg13g2_o21ai_1 _2323_ (.B1(net739),
    .Y(_1352_),
    .A1(_0993_),
    .A2(_1174_));
 sg13g2_nor3_1 _2324_ (.A(_1349_),
    .B(_1351_),
    .C(_1352_),
    .Y(_1353_));
 sg13g2_o21ai_1 _2325_ (.B1(net706),
    .Y(_1354_),
    .A1(_1348_),
    .A2(_1353_));
 sg13g2_and2_1 _2326_ (.A(net658),
    .B(_1354_),
    .X(_1355_));
 sg13g2_a21oi_1 _2327_ (.A1(net681),
    .A2(net660),
    .Y(_1356_),
    .B1(_1321_));
 sg13g2_nor2_1 _2328_ (.A(net769),
    .B(_1356_),
    .Y(_1357_));
 sg13g2_nor2b_1 _2329_ (.A(_1356_),
    .B_N(_1234_),
    .Y(_1358_));
 sg13g2_a21oi_1 _2330_ (.A1(net681),
    .A2(net669),
    .Y(_1359_),
    .B1(_1321_));
 sg13g2_o21ai_1 _2331_ (.B1(_1271_),
    .Y(_1360_),
    .A1(_1234_),
    .A2(_1359_));
 sg13g2_o21ai_1 _2332_ (.B1(net741),
    .Y(_1361_),
    .A1(_1358_),
    .A2(_1360_));
 sg13g2_a21o_1 _2333_ (.A2(_1089_),
    .A1(_1016_),
    .B1(_1122_),
    .X(_1362_));
 sg13g2_nand3_1 _2334_ (.B(net696),
    .C(_1105_),
    .A(net751),
    .Y(_1363_));
 sg13g2_nand4_1 _2335_ (.B(_1361_),
    .C(_1362_),
    .A(net711),
    .Y(_1364_),
    .D(_1363_));
 sg13g2_nor2_1 _2336_ (.A(net744),
    .B(net780),
    .Y(_1365_));
 sg13g2_o21ai_1 _2337_ (.B1(_1365_),
    .Y(_1366_),
    .A1(_1111_),
    .A2(_1321_));
 sg13g2_nor2_1 _2338_ (.A(_1127_),
    .B(_1356_),
    .Y(_1367_));
 sg13g2_a21oi_1 _2339_ (.A1(net751),
    .A2(net793),
    .Y(_1368_),
    .B1(_1118_));
 sg13g2_nor3_1 _2340_ (.A(net711),
    .B(_1367_),
    .C(_1368_),
    .Y(_1369_));
 sg13g2_a21oi_1 _2341_ (.A1(_1366_),
    .A2(_1369_),
    .Y(_1370_),
    .B1(net658));
 sg13g2_a221oi_1 _2342_ (.B2(_1370_),
    .C1(_0923_),
    .B1(_1364_),
    .A1(_1343_),
    .Y(_1371_),
    .A2(_1355_));
 sg13g2_or3_1 _2343_ (.A(_1132_),
    .B(_1329_),
    .C(_1371_),
    .X(_1372_));
 sg13g2_a21oi_2 _2344_ (.B1(_1321_),
    .Y(_1373_),
    .A2(_1083_),
    .A1(net731));
 sg13g2_nand2_1 _2345_ (.Y(_1374_),
    .A(net755),
    .B(_1373_));
 sg13g2_a22oi_1 _2346_ (.Y(_1375_),
    .B1(_1325_),
    .B2(_1374_),
    .A2(_1322_),
    .A1(_1165_));
 sg13g2_nand2b_2 _2347_ (.Y(_1376_),
    .B(_1172_),
    .A_N(_1159_));
 sg13g2_o21ai_1 _2348_ (.B1(net745),
    .Y(_1377_),
    .A1(net763),
    .A2(_1180_));
 sg13g2_a221oi_1 _2349_ (.B2(net701),
    .C1(_1377_),
    .B1(_1376_),
    .A1(_1098_),
    .Y(_1378_),
    .A2(_1173_));
 sg13g2_o21ai_1 _2350_ (.B1(_1181_),
    .Y(_1379_),
    .A1(net671),
    .A2(net659));
 sg13g2_a21oi_1 _2351_ (.A1(net676),
    .A2(net659),
    .Y(_1380_),
    .B1(_1169_));
 sg13g2_o21ai_1 _2352_ (.B1(_1379_),
    .Y(_1381_),
    .A1(_1035_),
    .A2(_1380_));
 sg13g2_o21ai_1 _2353_ (.B1(net708),
    .Y(_1382_),
    .A1(_1311_),
    .A2(_1381_));
 sg13g2_nor2_1 _2354_ (.A(_1378_),
    .B(_1382_),
    .Y(_1383_));
 sg13g2_o21ai_1 _2355_ (.B1(net656),
    .Y(_1384_),
    .A1(net707),
    .A2(_1375_));
 sg13g2_nor2_1 _2356_ (.A(_1383_),
    .B(_1384_),
    .Y(_1385_));
 sg13g2_a21oi_1 _2357_ (.A1(net700),
    .A2(_1134_),
    .Y(_1386_),
    .B1(net752));
 sg13g2_and4_1 _2358_ (.A(net737),
    .B(net722),
    .C(net720),
    .D(net716),
    .X(_1387_));
 sg13g2_nor2_2 _2359_ (.A(_1313_),
    .B(_1387_),
    .Y(_1388_));
 sg13g2_nor2_1 _2360_ (.A(_0935_),
    .B(_1388_),
    .Y(_1389_));
 sg13g2_o21ai_1 _2361_ (.B1(net768),
    .Y(_1390_),
    .A1(_1294_),
    .A2(_1389_));
 sg13g2_a21oi_1 _2362_ (.A1(net704),
    .A2(_1066_),
    .Y(_1391_),
    .B1(net742));
 sg13g2_a221oi_1 _2363_ (.B2(net804),
    .C1(net679),
    .B1(_1112_),
    .A1(net716),
    .Y(_1392_),
    .A2(_1048_));
 sg13g2_o21ai_1 _2364_ (.B1(_1391_),
    .Y(_1393_),
    .A1(_1099_),
    .A2(_1392_));
 sg13g2_a21oi_1 _2365_ (.A1(net761),
    .A2(_1291_),
    .Y(_1394_),
    .B1(_1393_));
 sg13g2_a221oi_1 _2366_ (.B2(_1394_),
    .C1(net712),
    .B1(_1390_),
    .A1(_1299_),
    .Y(_1395_),
    .A2(_1386_));
 sg13g2_nand2_1 _2367_ (.Y(_1396_),
    .A(_1226_),
    .B(_1306_));
 sg13g2_a22oi_1 _2368_ (.Y(_1397_),
    .B1(_1396_),
    .B2(net703),
    .A2(_1214_),
    .A1(_1034_));
 sg13g2_nor3_1 _2369_ (.A(net760),
    .B(net779),
    .C(_1160_),
    .Y(_1398_));
 sg13g2_a221oi_1 _2370_ (.B2(_1376_),
    .C1(_1398_),
    .B1(_1251_),
    .A1(net699),
    .Y(_1399_),
    .A2(_1222_));
 sg13g2_a221oi_1 _2371_ (.B2(_1225_),
    .C1(net705),
    .B1(_1399_),
    .A1(_1303_),
    .Y(_1400_),
    .A2(_1397_));
 sg13g2_nor3_1 _2372_ (.A(net656),
    .B(_1395_),
    .C(_1400_),
    .Y(_1401_));
 sg13g2_o21ai_1 _2373_ (.B1(_0923_),
    .Y(_1402_),
    .A1(_1385_),
    .A2(_1401_));
 sg13g2_o21ai_1 _2374_ (.B1(net805),
    .Y(_1403_),
    .A1(_1313_),
    .A2(_1387_));
 sg13g2_a21oi_1 _2375_ (.A1(_1346_),
    .A2(_1403_),
    .Y(_1404_),
    .B1(net697));
 sg13g2_nor4_1 _2376_ (.A(_1333_),
    .B(_1335_),
    .C(_1336_),
    .D(_1404_),
    .Y(_1405_));
 sg13g2_a21oi_1 _2377_ (.A1(_1126_),
    .A2(_1340_),
    .Y(_1406_),
    .B1(net709));
 sg13g2_o21ai_1 _2378_ (.B1(_1406_),
    .Y(_1407_),
    .A1(_1260_),
    .A2(_1405_));
 sg13g2_nor2_1 _2379_ (.A(net809),
    .B(net685),
    .Y(_1408_));
 sg13g2_a221oi_1 _2380_ (.B2(_1002_),
    .C1(net696),
    .B1(_1408_),
    .A1(net808),
    .Y(_1409_),
    .A2(_1244_));
 sg13g2_nor4_1 _2381_ (.A(_1255_),
    .B(_1344_),
    .C(_1347_),
    .D(_1409_),
    .Y(_1410_));
 sg13g2_nand2_2 _2382_ (.Y(_1411_),
    .A(net747),
    .B(net699));
 sg13g2_a21oi_1 _2383_ (.A1(net688),
    .A2(_1012_),
    .Y(_1412_),
    .B1(net806));
 sg13g2_a221oi_1 _2384_ (.B2(_1412_),
    .C1(_1411_),
    .B1(_1092_),
    .A1(net806),
    .Y(_1413_),
    .A2(_0993_));
 sg13g2_nor3_1 _2385_ (.A(net748),
    .B(net699),
    .C(_1244_),
    .Y(_1414_));
 sg13g2_nor3_1 _2386_ (.A(net710),
    .B(_1413_),
    .C(_1414_),
    .Y(_1415_));
 sg13g2_o21ai_1 _2387_ (.B1(_1415_),
    .Y(_1416_),
    .A1(net739),
    .A2(_1410_));
 sg13g2_nand3_1 _2388_ (.B(_1407_),
    .C(_1416_),
    .A(net656),
    .Y(_1417_));
 sg13g2_nor2_1 _2389_ (.A(_1035_),
    .B(_1359_),
    .Y(_1418_));
 sg13g2_o21ai_1 _2390_ (.B1(net744),
    .Y(_1419_),
    .A1(_1357_),
    .A2(_1418_));
 sg13g2_o21ai_1 _2391_ (.B1(net703),
    .Y(_1420_),
    .A1(net672),
    .A2(net669));
 sg13g2_nor2_1 _2392_ (.A(net750),
    .B(_1251_),
    .Y(_1421_));
 sg13g2_a22oi_1 _2393_ (.Y(_1422_),
    .B1(_1420_),
    .B2(_1421_),
    .A2(_1089_),
    .A1(_1016_));
 sg13g2_o21ai_1 _2394_ (.B1(net711),
    .Y(_1423_),
    .A1(_1127_),
    .A2(_1247_));
 sg13g2_nor2_1 _2395_ (.A(_1422_),
    .B(_1423_),
    .Y(_1424_));
 sg13g2_nor2_1 _2396_ (.A(net710),
    .B(_1367_),
    .Y(_1425_));
 sg13g2_a221oi_1 _2397_ (.B2(_1373_),
    .C1(net658),
    .B1(_1425_),
    .A1(_1419_),
    .Y(_1426_),
    .A2(_1424_));
 sg13g2_nor2_1 _2398_ (.A(_0923_),
    .B(_1426_),
    .Y(_1427_));
 sg13g2_a21oi_1 _2399_ (.A1(_1417_),
    .A2(_1427_),
    .Y(_1428_),
    .B1(_1133_));
 sg13g2_a21oi_1 _2400_ (.A1(_1402_),
    .A2(_1428_),
    .Y(_1429_),
    .B1(_0901_));
 sg13g2_a21oi_1 _2401_ (.A1(_1372_),
    .A2(_1429_),
    .Y(_1430_),
    .B1(_1288_));
 sg13g2_or3_2 _2402_ (.A(_1005_),
    .B(net667),
    .C(net666),
    .X(_1431_));
 sg13g2_a21o_2 _2403_ (.A2(net667),
    .A1(net675),
    .B1(_1005_),
    .X(_1432_));
 sg13g2_a22oi_1 _2404_ (.Y(_1433_),
    .B1(_1432_),
    .B2(_1024_),
    .A2(_1431_),
    .A1(_1181_));
 sg13g2_o21ai_1 _2405_ (.B1(net707),
    .Y(_1434_),
    .A1(net746),
    .A2(_1433_));
 sg13g2_nand2_1 _2406_ (.Y(_1435_),
    .A(net664),
    .B(_1115_));
 sg13g2_a21oi_2 _2407_ (.B1(_1169_),
    .Y(_1436_),
    .A2(_1115_),
    .A1(net664));
 sg13g2_or2_1 _2408_ (.X(_1437_),
    .B(_1436_),
    .A(net768));
 sg13g2_and3_1 _2409_ (.X(_1438_),
    .A(net788),
    .B(net664),
    .C(_1115_));
 sg13g2_a21o_1 _2410_ (.A2(_1432_),
    .A1(net794),
    .B1(_1438_),
    .X(_1439_));
 sg13g2_a221oi_1 _2411_ (.B2(net794),
    .C1(_1438_),
    .B1(_1432_),
    .A1(net689),
    .Y(_1440_),
    .A2(_1112_));
 sg13g2_o21ai_1 _2412_ (.B1(_1437_),
    .Y(_1441_),
    .A1(net762),
    .A2(_1440_));
 sg13g2_a21oi_1 _2413_ (.A1(net742),
    .A2(_1441_),
    .Y(_1442_),
    .B1(_1434_));
 sg13g2_o21ai_1 _2414_ (.B1(_1170_),
    .Y(_1443_),
    .A1(net668),
    .A2(net666));
 sg13g2_nor2_1 _2415_ (.A(net697),
    .B(_1443_),
    .Y(_1444_));
 sg13g2_nor4_1 _2416_ (.A(net736),
    .B(_0964_),
    .C(_0966_),
    .D(_1008_),
    .Y(_1445_));
 sg13g2_a21o_2 _2417_ (.A2(net664),
    .A1(net672),
    .B1(_1445_),
    .X(_1446_));
 sg13g2_nor3_1 _2418_ (.A(net707),
    .B(_1444_),
    .C(_1446_),
    .Y(_1447_));
 sg13g2_nand2_1 _2419_ (.Y(_1448_),
    .A(net812),
    .B(_1431_));
 sg13g2_o21ai_1 _2420_ (.B1(_1448_),
    .Y(_1449_),
    .A1(_1234_),
    .A2(_1237_));
 sg13g2_a21oi_1 _2421_ (.A1(net696),
    .A2(_1443_),
    .Y(_1450_),
    .B1(net754));
 sg13g2_nand2_1 _2422_ (.Y(_1451_),
    .A(_1449_),
    .B(_1450_));
 sg13g2_a21o_1 _2423_ (.A2(_1451_),
    .A1(_1447_),
    .B1(_1442_),
    .X(_1452_));
 sg13g2_o21ai_1 _2424_ (.B1(_0989_),
    .Y(_1453_),
    .A1(_1051_),
    .A2(net670));
 sg13g2_o21ai_1 _2425_ (.B1(net804),
    .Y(_1454_),
    .A1(net678),
    .A2(net673));
 sg13g2_nand3_1 _2426_ (.B(_1453_),
    .C(_1454_),
    .A(_1211_),
    .Y(_1455_));
 sg13g2_and2_1 _2427_ (.A(_1028_),
    .B(_1049_),
    .X(_1456_));
 sg13g2_nand3_1 _2428_ (.B(_1028_),
    .C(_1049_),
    .A(net761),
    .Y(_1457_));
 sg13g2_nor2b_1 _2429_ (.A(_1457_),
    .B_N(_1204_),
    .Y(_1458_));
 sg13g2_and4_1 _2430_ (.A(net790),
    .B(net800),
    .C(net687),
    .D(net677),
    .X(_1459_));
 sg13g2_a221oi_1 _2431_ (.B2(net790),
    .C1(_1459_),
    .B1(_1142_),
    .A1(_0985_),
    .Y(_1460_),
    .A2(_0986_));
 sg13g2_nand3b_1 _2432_ (.B(_1070_),
    .C(_1028_),
    .Y(_1461_),
    .A_N(_1143_));
 sg13g2_a22oi_1 _2433_ (.Y(_1462_),
    .B1(_1461_),
    .B2(net780),
    .A2(_1142_),
    .A1(_1010_));
 sg13g2_a21o_1 _2434_ (.A2(_1462_),
    .A1(_1460_),
    .B1(_1458_),
    .X(_1463_));
 sg13g2_a21oi_1 _2435_ (.A1(net752),
    .A2(_1463_),
    .Y(_1464_),
    .B1(net712));
 sg13g2_o21ai_1 _2436_ (.B1(_1464_),
    .Y(_1465_),
    .A1(_1209_),
    .A2(_1455_));
 sg13g2_a21oi_1 _2437_ (.A1(net652),
    .A2(_1146_),
    .Y(_1466_),
    .B1(net807));
 sg13g2_o21ai_1 _2438_ (.B1(net698),
    .Y(_1467_),
    .A1(_1216_),
    .A2(_1466_));
 sg13g2_a21oi_1 _2439_ (.A1(_0973_),
    .A2(_1145_),
    .Y(_1468_),
    .B1(net757));
 sg13g2_a21oi_1 _2440_ (.A1(net692),
    .A2(net677),
    .Y(_1469_),
    .B1(net684));
 sg13g2_nor2_1 _2441_ (.A(net800),
    .B(_1039_),
    .Y(_1470_));
 sg13g2_nor3_1 _2442_ (.A(_1099_),
    .B(_1469_),
    .C(_1470_),
    .Y(_1471_));
 sg13g2_nor4_1 _2443_ (.A(net748),
    .B(_1218_),
    .C(_1468_),
    .D(_1471_),
    .Y(_1472_));
 sg13g2_nand2_1 _2444_ (.Y(_1473_),
    .A(net663),
    .B(_1123_));
 sg13g2_a21o_1 _2445_ (.A2(_1473_),
    .A1(_1170_),
    .B1(_1263_),
    .X(_1474_));
 sg13g2_nor2_1 _2446_ (.A(net682),
    .B(net680),
    .Y(_1475_));
 sg13g2_nor3_1 _2447_ (.A(net800),
    .B(net764),
    .C(_1475_),
    .Y(_1476_));
 sg13g2_nand2_1 _2448_ (.Y(_1477_),
    .A(_0934_),
    .B(net758));
 sg13g2_o21ai_1 _2449_ (.B1(net748),
    .Y(_1478_),
    .A1(_1475_),
    .A2(_1477_));
 sg13g2_o21ai_1 _2450_ (.B1(_1436_),
    .Y(_1479_),
    .A1(net791),
    .A2(_1473_));
 sg13g2_a21oi_2 _2451_ (.B1(net682),
    .Y(_1480_),
    .A2(_1012_),
    .A1(net687));
 sg13g2_o21ai_1 _2452_ (.B1(_1226_),
    .Y(_1481_),
    .A1(net807),
    .A2(_1480_));
 sg13g2_a221oi_1 _2453_ (.B2(net698),
    .C1(_1478_),
    .B1(_1481_),
    .A1(net765),
    .Y(_1482_),
    .A2(_1479_));
 sg13g2_a221oi_1 _2454_ (.B2(_1482_),
    .C1(net705),
    .B1(_1474_),
    .A1(_1467_),
    .Y(_1483_),
    .A2(_1472_));
 sg13g2_nor2_1 _2455_ (.A(net655),
    .B(_1483_),
    .Y(_1484_));
 sg13g2_a221oi_1 _2456_ (.B2(_1484_),
    .C1(net650),
    .B1(_1465_),
    .A1(net656),
    .Y(_1485_),
    .A2(_1452_));
 sg13g2_nor3_1 _2457_ (.A(net810),
    .B(_1051_),
    .C(net670),
    .Y(_1486_));
 sg13g2_o21ai_1 _2458_ (.B1(net794),
    .Y(_1487_),
    .A1(net673),
    .A2(net670));
 sg13g2_a21o_1 _2459_ (.A2(_1487_),
    .A1(net777),
    .B1(_1486_),
    .X(_1488_));
 sg13g2_nand4_1 _2460_ (.B(_1058_),
    .C(_1332_),
    .A(net752),
    .Y(_1489_),
    .D(_1488_));
 sg13g2_nor3_1 _2461_ (.A(net787),
    .B(net678),
    .C(_1048_),
    .Y(_1490_));
 sg13g2_nand3_1 _2462_ (.B(_1028_),
    .C(_1049_),
    .A(net787),
    .Y(_1491_));
 sg13g2_nand3b_1 _2463_ (.B(_1491_),
    .C(net767),
    .Y(_1492_),
    .A_N(_1490_));
 sg13g2_and2_1 _2464_ (.A(net760),
    .B(_1010_),
    .X(_1493_));
 sg13g2_a221oi_1 _2465_ (.B2(_1068_),
    .C1(net753),
    .B1(_1493_),
    .A1(_1030_),
    .Y(_1494_),
    .A2(_1234_));
 sg13g2_mux4_1 _2466_ (.S0(net808),
    .A0(net729),
    .A1(_1025_),
    .A2(_1069_),
    .A3(_1066_),
    .S1(net687),
    .X(_0117_));
 sg13g2_nand2_1 _2467_ (.Y(_0118_),
    .A(net695),
    .B(_0117_));
 sg13g2_or2_1 _2468_ (.X(_0119_),
    .B(_1289_),
    .A(net761));
 sg13g2_nand4_1 _2469_ (.B(_1494_),
    .C(_0118_),
    .A(_1492_),
    .Y(_0120_),
    .D(_0119_));
 sg13g2_and2_1 _2470_ (.A(net710),
    .B(_0120_),
    .X(_0121_));
 sg13g2_a221oi_1 _2471_ (.B2(net733),
    .C1(net772),
    .B1(net770),
    .A1(net721),
    .Y(_0122_),
    .A2(net719));
 sg13g2_nand3_1 _2472_ (.B(net690),
    .C(_1011_),
    .A(net774),
    .Y(_0123_));
 sg13g2_a221oi_1 _2473_ (.B2(net809),
    .C1(_0122_),
    .B1(_1036_),
    .A1(net688),
    .Y(_0124_),
    .A2(net681));
 sg13g2_o21ai_1 _2474_ (.B1(_0123_),
    .Y(_0125_),
    .A1(_1408_),
    .A2(_1412_));
 sg13g2_o21ai_1 _2475_ (.B1(net718),
    .Y(_0126_),
    .A1(net733),
    .A2(net716));
 sg13g2_nor2_1 _2476_ (.A(net680),
    .B(_0126_),
    .Y(_0127_));
 sg13g2_nand2_1 _2477_ (.Y(_0128_),
    .A(net792),
    .B(_1036_));
 sg13g2_a21oi_1 _2478_ (.A1(_0127_),
    .A2(_0128_),
    .Y(_0129_),
    .B1(net765));
 sg13g2_a221oi_1 _2479_ (.B2(_0125_),
    .C1(_0129_),
    .B1(net703),
    .A1(_0914_),
    .Y(_0130_),
    .A2(_0927_));
 sg13g2_o21ai_1 _2480_ (.B1(_0130_),
    .Y(_0131_),
    .A1(_1035_),
    .A2(_0124_));
 sg13g2_nor2_1 _2481_ (.A(net685),
    .B(_0122_),
    .Y(_0132_));
 sg13g2_o21ai_1 _2482_ (.B1(_1175_),
    .Y(_0133_),
    .A1(net685),
    .A2(_0122_));
 sg13g2_o21ai_1 _2483_ (.B1(net757),
    .Y(_0134_),
    .A1(_0957_),
    .A2(_0972_));
 sg13g2_nand3_1 _2484_ (.B(_0133_),
    .C(_0134_),
    .A(net748),
    .Y(_0135_));
 sg13g2_nor2_1 _2485_ (.A(net780),
    .B(net778),
    .Y(_0136_));
 sg13g2_o21ai_1 _2486_ (.B1(_0136_),
    .Y(_0137_),
    .A1(_1025_),
    .A2(_1159_));
 sg13g2_o21ai_1 _2487_ (.B1(net780),
    .Y(_0138_),
    .A1(_0972_),
    .A2(_1025_));
 sg13g2_a21oi_1 _2488_ (.A1(_0137_),
    .A2(_0138_),
    .Y(_0139_),
    .B1(net757));
 sg13g2_nor4_1 _2489_ (.A(net786),
    .B(net807),
    .C(net758),
    .D(_1029_),
    .Y(_0140_));
 sg13g2_nor3_1 _2490_ (.A(_0135_),
    .B(_0139_),
    .C(_0140_),
    .Y(_0141_));
 sg13g2_nor2_1 _2491_ (.A(net710),
    .B(_0141_),
    .Y(_0142_));
 sg13g2_a221oi_1 _2492_ (.B2(_0142_),
    .C1(net654),
    .B1(_0131_),
    .A1(_1489_),
    .Y(_0143_),
    .A2(_0121_));
 sg13g2_a221oi_1 _2493_ (.B2(net663),
    .C1(net793),
    .B1(net665),
    .A1(_1000_),
    .Y(_0144_),
    .A2(net669));
 sg13g2_and2_1 _2494_ (.A(net690),
    .B(_1091_),
    .X(_0145_));
 sg13g2_mux2_2 _2495_ (.A0(_1091_),
    .A1(_1101_),
    .S(net688),
    .X(_0146_));
 sg13g2_a221oi_1 _2496_ (.B2(net802),
    .C1(net785),
    .B1(_0146_),
    .A1(_1145_),
    .Y(_0147_),
    .A2(_1192_));
 sg13g2_o21ai_1 _2497_ (.B1(net662),
    .Y(_0148_),
    .A1(_0144_),
    .A2(_0147_));
 sg13g2_nor2_1 _2498_ (.A(net662),
    .B(_1446_),
    .Y(_0149_));
 sg13g2_nor2_1 _2499_ (.A(net711),
    .B(_0149_),
    .Y(_0150_));
 sg13g2_nor2_1 _2500_ (.A(_1270_),
    .B(_0126_),
    .Y(_0151_));
 sg13g2_nand2_1 _2501_ (.Y(_0152_),
    .A(net662),
    .B(_0151_));
 sg13g2_nor2_1 _2502_ (.A(_1091_),
    .B(_1270_),
    .Y(_0153_));
 sg13g2_a22oi_1 _2503_ (.Y(_0154_),
    .B1(_1121_),
    .B2(_0153_),
    .A2(net792),
    .A1(net750));
 sg13g2_o21ai_1 _2504_ (.B1(net809),
    .Y(_0155_),
    .A1(_1270_),
    .A2(_0126_));
 sg13g2_o21ai_1 _2505_ (.B1(net802),
    .Y(_0156_),
    .A1(net680),
    .A2(_0126_));
 sg13g2_nand2_1 _2506_ (.Y(_0157_),
    .A(_0155_),
    .B(_0156_));
 sg13g2_a22oi_1 _2507_ (.Y(_0158_),
    .B1(_0157_),
    .B2(net703),
    .A2(_0154_),
    .A1(_0152_));
 sg13g2_o21ai_1 _2508_ (.B1(_0158_),
    .Y(_0159_),
    .A1(_1099_),
    .A2(_0151_));
 sg13g2_nand3_1 _2509_ (.B(_1084_),
    .C(_1251_),
    .A(net675),
    .Y(_0160_));
 sg13g2_nor2b_1 _2510_ (.A(_0146_),
    .B_N(_0160_),
    .Y(_0161_));
 sg13g2_a21oi_1 _2511_ (.A1(net741),
    .A2(_0161_),
    .Y(_0162_),
    .B1(net706));
 sg13g2_a221oi_1 _2512_ (.B2(_0162_),
    .C1(net655),
    .B1(_0159_),
    .A1(_0148_),
    .Y(_0163_),
    .A2(_0150_));
 sg13g2_nor3_1 _2513_ (.A(_0923_),
    .B(_0143_),
    .C(_0163_),
    .Y(_0164_));
 sg13g2_o21ai_1 _2514_ (.B1(_1133_),
    .Y(_0165_),
    .A1(_1485_),
    .A2(_0164_));
 sg13g2_a21o_1 _2515_ (.A2(_0145_),
    .A1(net809),
    .B1(_1087_),
    .X(_0166_));
 sg13g2_o21ai_1 _2516_ (.B1(net765),
    .Y(_0167_),
    .A1(net777),
    .A2(_0153_));
 sg13g2_a221oi_1 _2517_ (.B2(_0136_),
    .C1(_0167_),
    .B1(_0166_),
    .A1(net785),
    .Y(_0168_),
    .A2(_0146_));
 sg13g2_a221oi_1 _2518_ (.B2(net792),
    .C1(net765),
    .B1(_0145_),
    .A1(_1145_),
    .Y(_0169_),
    .A2(_1192_));
 sg13g2_or2_1 _2519_ (.X(_0170_),
    .B(_0169_),
    .A(net750));
 sg13g2_nand3_1 _2520_ (.B(_0155_),
    .C(_0156_),
    .A(net785),
    .Y(_0171_));
 sg13g2_a21oi_1 _2521_ (.A1(net792),
    .A2(_0127_),
    .Y(_0172_),
    .B1(_1127_));
 sg13g2_nor2_1 _2522_ (.A(_1122_),
    .B(_0153_),
    .Y(_0173_));
 sg13g2_a21oi_1 _2523_ (.A1(_0171_),
    .A2(_0172_),
    .Y(_0174_),
    .B1(_0173_));
 sg13g2_o21ai_1 _2524_ (.B1(_0174_),
    .Y(_0175_),
    .A1(_0168_),
    .A2(_0170_));
 sg13g2_nand4_1 _2525_ (.B(_1058_),
    .C(_1332_),
    .A(net752),
    .Y(_0176_),
    .D(_1487_));
 sg13g2_mux2_1 _2526_ (.A0(_1072_),
    .A1(_1141_),
    .S(net767),
    .X(_0177_));
 sg13g2_a21oi_1 _2527_ (.A1(_1494_),
    .A2(_0177_),
    .Y(_0178_),
    .B1(net653));
 sg13g2_a22oi_1 _2528_ (.Y(_0179_),
    .B1(_0176_),
    .B2(_0178_),
    .A2(_0175_),
    .A1(net653));
 sg13g2_nor2_1 _2529_ (.A(net802),
    .B(net680),
    .Y(_0180_));
 sg13g2_nor2_1 _2530_ (.A(net809),
    .B(_0972_),
    .Y(_0181_));
 sg13g2_nor2_1 _2531_ (.A(net792),
    .B(_1036_),
    .Y(_0182_));
 sg13g2_o21ai_1 _2532_ (.B1(_0182_),
    .Y(_0183_),
    .A1(_0180_),
    .A2(_0181_));
 sg13g2_a21oi_1 _2533_ (.A1(net792),
    .A2(_0132_),
    .Y(_0184_),
    .B1(net759));
 sg13g2_nand2_1 _2534_ (.Y(_0185_),
    .A(net809),
    .B(_0127_));
 sg13g2_a221oi_1 _2535_ (.B2(_0129_),
    .C1(net750),
    .B1(_0185_),
    .A1(_0183_),
    .Y(_0186_),
    .A2(_0184_));
 sg13g2_o21ai_1 _2536_ (.B1(_1010_),
    .Y(_0187_),
    .A1(_1025_),
    .A2(_1159_));
 sg13g2_o21ai_1 _2537_ (.B1(net662),
    .Y(_0188_),
    .A1(_0973_),
    .A2(_0990_));
 sg13g2_o21ai_1 _2538_ (.B1(_0187_),
    .Y(_0189_),
    .A1(net785),
    .A2(_1029_));
 sg13g2_a21oi_1 _2539_ (.A1(_1121_),
    .A2(_0132_),
    .Y(_0190_),
    .B1(net654));
 sg13g2_o21ai_1 _2540_ (.B1(_0190_),
    .Y(_0191_),
    .A1(_0188_),
    .A2(_0189_));
 sg13g2_a221oi_1 _2541_ (.B2(net785),
    .C1(_1122_),
    .B1(_1446_),
    .A1(net652),
    .Y(_0192_),
    .A2(_1124_));
 sg13g2_a221oi_1 _2542_ (.B2(_1114_),
    .C1(_1446_),
    .B1(net699),
    .A1(_0914_),
    .Y(_0193_),
    .A2(_0927_));
 sg13g2_a21oi_1 _2543_ (.A1(_1145_),
    .A2(_1192_),
    .Y(_0194_),
    .B1(_1127_));
 sg13g2_or4_1 _2544_ (.A(net655),
    .B(_0192_),
    .C(_0193_),
    .D(_0194_),
    .X(_0195_));
 sg13g2_o21ai_1 _2545_ (.B1(_0195_),
    .Y(_0196_),
    .A1(_0186_),
    .A2(_0191_));
 sg13g2_a21oi_1 _2546_ (.A1(net706),
    .A2(_0196_),
    .Y(_0197_),
    .B1(_0923_));
 sg13g2_o21ai_1 _2547_ (.B1(_0197_),
    .Y(_0198_),
    .A1(net707),
    .A2(_0179_));
 sg13g2_o21ai_1 _2548_ (.B1(net708),
    .Y(_0199_),
    .A1(net769),
    .A2(_1436_));
 sg13g2_o21ai_1 _2549_ (.B1(net768),
    .Y(_0200_),
    .A1(_1169_),
    .A2(_1432_));
 sg13g2_nand2b_1 _2550_ (.Y(_0201_),
    .B(_0200_),
    .A_N(_0199_));
 sg13g2_nand3_1 _2551_ (.B(net665),
    .C(net663),
    .A(net704),
    .Y(_0202_));
 sg13g2_nand3_1 _2552_ (.B(_1193_),
    .C(_0202_),
    .A(net714),
    .Y(_0203_));
 sg13g2_nand3_1 _2553_ (.B(_0201_),
    .C(_0203_),
    .A(net744),
    .Y(_0204_));
 sg13g2_o21ai_1 _2554_ (.B1(net761),
    .Y(_0205_),
    .A1(net779),
    .A2(_1170_));
 sg13g2_nor2_1 _2555_ (.A(_1432_),
    .B(_0205_),
    .Y(_0206_));
 sg13g2_nor4_1 _2556_ (.A(net795),
    .B(_0964_),
    .C(_0966_),
    .D(net771),
    .Y(_0207_));
 sg13g2_or3_1 _2557_ (.A(net667),
    .B(net666),
    .C(_0207_),
    .X(_0208_));
 sg13g2_and2_1 _2558_ (.A(net787),
    .B(_1432_),
    .X(_0209_));
 sg13g2_a221oi_1 _2559_ (.B2(_0990_),
    .C1(net763),
    .B1(_0208_),
    .A1(net788),
    .Y(_0210_),
    .A2(_1432_));
 sg13g2_o21ai_1 _2560_ (.B1(net707),
    .Y(_0211_),
    .A1(_0206_),
    .A2(_0210_));
 sg13g2_and2_1 _2561_ (.A(_1114_),
    .B(_1251_),
    .X(_0212_));
 sg13g2_nor4_1 _2562_ (.A(net707),
    .B(_1444_),
    .C(_1446_),
    .D(_0212_),
    .Y(_0213_));
 sg13g2_nand3b_1 _2563_ (.B(net754),
    .C(_0211_),
    .Y(_0214_),
    .A_N(_0213_));
 sg13g2_a21oi_1 _2564_ (.A1(_0204_),
    .A2(_0214_),
    .Y(_0215_),
    .B1(net653));
 sg13g2_nand3_1 _2565_ (.B(_1139_),
    .C(_1454_),
    .A(_1138_),
    .Y(_0216_));
 sg13g2_nand2_1 _2566_ (.Y(_0217_),
    .A(net743),
    .B(_0216_));
 sg13g2_a221oi_1 _2567_ (.B2(_1460_),
    .C1(net743),
    .B1(_1144_),
    .A1(net760),
    .Y(_0218_),
    .A2(_1141_));
 sg13g2_nor2_1 _2568_ (.A(net712),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_a21oi_1 _2569_ (.A1(net687),
    .A2(_1012_),
    .Y(_0220_),
    .B1(_1123_));
 sg13g2_nand2_1 _2570_ (.Y(_0221_),
    .A(net786),
    .B(_1154_));
 sg13g2_a21o_1 _2571_ (.A2(_1146_),
    .A1(net652),
    .B1(_1477_),
    .X(_0222_));
 sg13g2_a21o_1 _2572_ (.A2(_1145_),
    .A1(_0973_),
    .B1(_1263_),
    .X(_0223_));
 sg13g2_o21ai_1 _2573_ (.B1(_1436_),
    .Y(_0224_),
    .A1(_0990_),
    .A2(_1473_));
 sg13g2_nand3_1 _2574_ (.B(_0222_),
    .C(_0223_),
    .A(_1157_),
    .Y(_0225_));
 sg13g2_o21ai_1 _2575_ (.B1(_0221_),
    .Y(_0226_),
    .A1(_0935_),
    .A2(_0220_));
 sg13g2_o21ai_1 _2576_ (.B1(net710),
    .Y(_0227_),
    .A1(net739),
    .A2(_1474_));
 sg13g2_a21oi_1 _2577_ (.A1(_1121_),
    .A2(_0226_),
    .Y(_0228_),
    .B1(_0227_));
 sg13g2_a22oi_1 _2578_ (.Y(_0229_),
    .B1(_0225_),
    .B2(net739),
    .A2(_0224_),
    .A1(net662));
 sg13g2_a221oi_1 _2579_ (.B2(_0229_),
    .C1(net655),
    .B1(_0228_),
    .A1(_0217_),
    .Y(_0230_),
    .A2(_0219_));
 sg13g2_nor3_1 _2580_ (.A(net650),
    .B(_0215_),
    .C(_0230_),
    .Y(_0231_));
 sg13g2_nand3b_1 _2581_ (.B(_1132_),
    .C(_0198_),
    .Y(_0232_),
    .A_N(_0231_));
 sg13g2_nand3_1 _2582_ (.B(_0165_),
    .C(_0232_),
    .A(_0900_),
    .Y(_0233_));
 sg13g2_nor3_1 _2583_ (.A(net810),
    .B(_1005_),
    .C(_1053_),
    .Y(_0234_));
 sg13g2_nor3_1 _2584_ (.A(net804),
    .B(_1051_),
    .C(net670),
    .Y(_0235_));
 sg13g2_nand2b_1 _2585_ (.Y(_0236_),
    .B(net661),
    .A_N(_0235_));
 sg13g2_o21ai_1 _2586_ (.B1(net713),
    .Y(_0237_),
    .A1(_0234_),
    .A2(_0236_));
 sg13g2_or3_1 _2587_ (.A(net803),
    .B(_1005_),
    .C(_1053_),
    .X(_0238_));
 sg13g2_nand2_1 _2588_ (.Y(_0239_),
    .A(net704),
    .B(_0238_));
 sg13g2_a21oi_1 _2589_ (.A1(net774),
    .A2(net690),
    .Y(_0240_),
    .B1(net747));
 sg13g2_nor2_1 _2590_ (.A(net787),
    .B(_1039_),
    .Y(_0241_));
 sg13g2_nor4_2 _2591_ (.A(net746),
    .B(net678),
    .C(_1051_),
    .Y(_0242_),
    .D(_0241_));
 sg13g2_o21ai_1 _2592_ (.B1(_0239_),
    .Y(_0243_),
    .A1(net661),
    .A2(_0242_));
 sg13g2_a21oi_1 _2593_ (.A1(net803),
    .A2(_1051_),
    .Y(_0244_),
    .B1(net678));
 sg13g2_nand2_1 _2594_ (.Y(_0245_),
    .A(net803),
    .B(net729));
 sg13g2_nand3_1 _2595_ (.B(_1069_),
    .C(_0245_),
    .A(net689),
    .Y(_0246_));
 sg13g2_a22oi_1 _2596_ (.Y(_0247_),
    .B1(_0246_),
    .B2(_1034_),
    .A2(_0244_),
    .A1(net703));
 sg13g2_nor3_1 _2597_ (.A(_1048_),
    .B(_1083_),
    .C(_0247_),
    .Y(_0248_));
 sg13g2_nand3_1 _2598_ (.B(_1067_),
    .C(_1084_),
    .A(_1049_),
    .Y(_0249_));
 sg13g2_a221oi_1 _2599_ (.B2(net794),
    .C1(net767),
    .B1(_0249_),
    .A1(_1010_),
    .Y(_0250_),
    .A2(_1480_));
 sg13g2_nand3_1 _2600_ (.B(_1065_),
    .C(_1084_),
    .A(_1043_),
    .Y(_0251_));
 sg13g2_a21oi_1 _2601_ (.A1(net700),
    .A2(_0251_),
    .Y(_0252_),
    .B1(net753));
 sg13g2_o21ai_1 _2602_ (.B1(_0252_),
    .Y(_0253_),
    .A1(_0248_),
    .A2(_0250_));
 sg13g2_a21oi_1 _2603_ (.A1(_0243_),
    .A2(_0253_),
    .Y(_0254_),
    .B1(_0237_));
 sg13g2_a21oi_1 _2604_ (.A1(_1008_),
    .A2(net675),
    .Y(_0255_),
    .B1(_1270_));
 sg13g2_a21oi_1 _2605_ (.A1(net802),
    .A2(_0220_),
    .Y(_0256_),
    .B1(_0255_));
 sg13g2_o21ai_1 _2606_ (.B1(_0240_),
    .Y(_0257_),
    .A1(_1408_),
    .A2(_0180_));
 sg13g2_o21ai_1 _2607_ (.B1(_0257_),
    .Y(_0258_),
    .A1(net749),
    .A2(_0256_));
 sg13g2_nand3_1 _2608_ (.B(_1016_),
    .C(_1050_),
    .A(net744),
    .Y(_0259_));
 sg13g2_or4_1 _2609_ (.A(net743),
    .B(net686),
    .C(_1064_),
    .D(_1083_),
    .X(_0260_));
 sg13g2_a21oi_1 _2610_ (.A1(_0259_),
    .A2(_0260_),
    .Y(_0261_),
    .B1(net701));
 sg13g2_a221oi_1 _2611_ (.B2(net701),
    .C1(_0261_),
    .B1(_0258_),
    .A1(net661),
    .Y(_0262_),
    .A2(_0241_));
 sg13g2_o21ai_1 _2612_ (.B1(net656),
    .Y(_0263_),
    .A1(net712),
    .A2(_0262_));
 sg13g2_a21oi_1 _2613_ (.A1(_0971_),
    .A2(_0977_),
    .Y(_0264_),
    .B1(_1387_));
 sg13g2_nand2_1 _2614_ (.Y(_0265_),
    .A(_1172_),
    .B(_0264_));
 sg13g2_nor3_1 _2615_ (.A(net794),
    .B(_0977_),
    .C(_0991_),
    .Y(_0266_));
 sg13g2_o21ai_1 _2616_ (.B1(_1172_),
    .Y(_0267_),
    .A1(net762),
    .A2(_0266_));
 sg13g2_nor3_2 _2617_ (.A(_1005_),
    .B(net667),
    .C(_1201_),
    .Y(_0268_));
 sg13g2_or2_1 _2618_ (.X(_0269_),
    .B(_1111_),
    .A(_1040_));
 sg13g2_a22oi_1 _2619_ (.Y(_0270_),
    .B1(_0269_),
    .B2(net795),
    .A2(_0268_),
    .A1(_0934_));
 sg13g2_a22oi_1 _2620_ (.Y(_0271_),
    .B1(_0267_),
    .B2(_0270_),
    .A2(_0265_),
    .A1(net761));
 sg13g2_nor2_1 _2621_ (.A(_1127_),
    .B(_0255_),
    .Y(_0272_));
 sg13g2_o21ai_1 _2622_ (.B1(net710),
    .Y(_0273_),
    .A1(_1122_),
    .A2(_0269_));
 sg13g2_a21oi_2 _2623_ (.B1(_0273_),
    .Y(_0274_),
    .A2(_0272_),
    .A1(_1120_));
 sg13g2_o21ai_1 _2624_ (.B1(_0274_),
    .Y(_0275_),
    .A1(net754),
    .A2(_0271_));
 sg13g2_o21ai_1 _2625_ (.B1(net707),
    .Y(_0276_),
    .A1(_1126_),
    .A2(_1388_));
 sg13g2_a21oi_1 _2626_ (.A1(net661),
    .A2(_0265_),
    .Y(_0277_),
    .B1(_0276_));
 sg13g2_nor2_1 _2627_ (.A(net657),
    .B(_0277_),
    .Y(_0278_));
 sg13g2_a21oi_1 _2628_ (.A1(_0275_),
    .A2(_0278_),
    .Y(_0279_),
    .B1(_0923_));
 sg13g2_o21ai_1 _2629_ (.B1(_0279_),
    .Y(_0280_),
    .A1(_0254_),
    .A2(_0263_));
 sg13g2_a21o_1 _2630_ (.A2(_1147_),
    .A1(net800),
    .B1(_1042_),
    .X(_0281_));
 sg13g2_o21ai_1 _2631_ (.B1(net739),
    .Y(_0282_),
    .A1(_1099_),
    .A2(_1469_));
 sg13g2_a21oi_1 _2632_ (.A1(net698),
    .A2(_0281_),
    .Y(_0283_),
    .B1(_0282_));
 sg13g2_nor2_1 _2633_ (.A(_1035_),
    .B(_1469_),
    .Y(_0284_));
 sg13g2_o21ai_1 _2634_ (.B1(net801),
    .Y(_0285_),
    .A1(net682),
    .A2(net680));
 sg13g2_a21oi_1 _2635_ (.A1(_1226_),
    .A2(_0285_),
    .Y(_0286_),
    .B1(_1024_));
 sg13g2_nor2_1 _2636_ (.A(_0284_),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_nand3_1 _2637_ (.B(net663),
    .C(_1123_),
    .A(net703),
    .Y(_0288_));
 sg13g2_nand2_1 _2638_ (.Y(_0289_),
    .A(net683),
    .B(net663));
 sg13g2_and4_1 _2639_ (.A(net748),
    .B(_1170_),
    .C(_0288_),
    .D(_0289_),
    .X(_0290_));
 sg13g2_o21ai_1 _2640_ (.B1(_1175_),
    .Y(_0291_),
    .A1(net682),
    .A2(net680));
 sg13g2_a221oi_1 _2641_ (.B2(_0291_),
    .C1(net705),
    .B1(_0290_),
    .A1(_0283_),
    .Y(_0292_),
    .A2(_0287_));
 sg13g2_nor2_1 _2642_ (.A(net804),
    .B(_1456_),
    .Y(_0293_));
 sg13g2_o21ai_1 _2643_ (.B1(net703),
    .Y(_0294_),
    .A1(_1042_),
    .A2(_0293_));
 sg13g2_o21ai_1 _2644_ (.B1(_1456_),
    .Y(_0295_),
    .A1(net810),
    .A2(_1070_));
 sg13g2_nand2_1 _2645_ (.Y(_0296_),
    .A(_1289_),
    .B(_1330_));
 sg13g2_a21oi_1 _2646_ (.A1(net689),
    .A2(_1066_),
    .Y(_0297_),
    .B1(_1143_));
 sg13g2_o21ai_1 _2647_ (.B1(net752),
    .Y(_0298_),
    .A1(_1035_),
    .A2(_0297_));
 sg13g2_a221oi_1 _2648_ (.B2(net701),
    .C1(_0298_),
    .B1(_0296_),
    .A1(net695),
    .Y(_0299_),
    .A2(_0295_));
 sg13g2_nor2_1 _2649_ (.A(net768),
    .B(_1486_),
    .Y(_0300_));
 sg13g2_o21ai_1 _2650_ (.B1(net794),
    .Y(_0301_),
    .A1(net679),
    .A2(net674));
 sg13g2_nand4_1 _2651_ (.B(_1211_),
    .C(_1453_),
    .A(net742),
    .Y(_0302_),
    .D(_0301_));
 sg13g2_a21oi_1 _2652_ (.A1(_0238_),
    .A2(_0300_),
    .Y(_0303_),
    .B1(_0302_));
 sg13g2_nand2b_1 _2653_ (.Y(_0304_),
    .B(net700),
    .A_N(_0234_));
 sg13g2_a221oi_1 _2654_ (.B2(_0304_),
    .C1(net712),
    .B1(_0303_),
    .A1(_0294_),
    .Y(_0305_),
    .A2(_0299_));
 sg13g2_o21ai_1 _2655_ (.B1(net654),
    .Y(_0306_),
    .A1(_0292_),
    .A2(_0305_));
 sg13g2_nor2_1 _2656_ (.A(net780),
    .B(_0268_),
    .Y(_0307_));
 sg13g2_o21ai_1 _2657_ (.B1(net661),
    .Y(_0308_),
    .A1(_0209_),
    .A2(_0307_));
 sg13g2_a21oi_1 _2658_ (.A1(net768),
    .A2(_1435_),
    .Y(_0309_),
    .B1(net752));
 sg13g2_a22oi_1 _2659_ (.Y(_0310_),
    .B1(_1479_),
    .B2(_0309_),
    .A2(_1439_),
    .A1(_1121_));
 sg13g2_nand3_1 _2660_ (.B(_0308_),
    .C(_0310_),
    .A(net708),
    .Y(_0311_));
 sg13g2_a22oi_1 _2661_ (.Y(_0312_),
    .B1(_1121_),
    .B2(net788),
    .A2(net696),
    .A1(net742));
 sg13g2_a21oi_1 _2662_ (.A1(_1171_),
    .A2(_0264_),
    .Y(_0313_),
    .B1(_0312_));
 sg13g2_nor2_1 _2663_ (.A(_1411_),
    .B(_0268_),
    .Y(_0314_));
 sg13g2_o21ai_1 _2664_ (.B1(net713),
    .Y(_0315_),
    .A1(_1165_),
    .A2(_1388_));
 sg13g2_nor3_1 _2665_ (.A(_0313_),
    .B(_0314_),
    .C(_0315_),
    .Y(_0316_));
 sg13g2_nor2_1 _2666_ (.A(net653),
    .B(_0316_),
    .Y(_0317_));
 sg13g2_a21oi_1 _2667_ (.A1(_0311_),
    .A2(_0317_),
    .Y(_0318_),
    .B1(net650));
 sg13g2_a21oi_1 _2668_ (.A1(_0306_),
    .A2(_0318_),
    .Y(_0319_),
    .B1(_1132_));
 sg13g2_a21oi_1 _2669_ (.A1(net807),
    .A2(_0284_),
    .Y(_0320_),
    .B1(_1218_));
 sg13g2_o21ai_1 _2670_ (.B1(_0285_),
    .Y(_0321_),
    .A1(net800),
    .A2(_1480_));
 sg13g2_a221oi_1 _2671_ (.B2(_1473_),
    .C1(net808),
    .B1(_1170_),
    .A1(_0985_),
    .Y(_0322_),
    .A2(_0986_));
 sg13g2_nor2b_1 _2672_ (.A(_0322_),
    .B_N(_0290_),
    .Y(_0323_));
 sg13g2_a21oi_1 _2673_ (.A1(net698),
    .A2(_0321_),
    .Y(_0324_),
    .B1(_1476_));
 sg13g2_a221oi_1 _2674_ (.B2(_0324_),
    .C1(net705),
    .B1(_0323_),
    .A1(_0283_),
    .Y(_0325_),
    .A2(_0320_));
 sg13g2_a21o_1 _2675_ (.A2(_0296_),
    .A1(net788),
    .B1(_1457_),
    .X(_0326_));
 sg13g2_o21ai_1 _2676_ (.B1(_1460_),
    .Y(_0327_),
    .A1(net794),
    .A2(_0297_));
 sg13g2_a21o_1 _2677_ (.A2(_0327_),
    .A1(_0326_),
    .B1(net742),
    .X(_0328_));
 sg13g2_a21oi_1 _2678_ (.A1(_1137_),
    .A2(_0303_),
    .Y(_0329_),
    .B1(net712));
 sg13g2_a21oi_1 _2679_ (.A1(_0328_),
    .A2(_0329_),
    .Y(_0330_),
    .B1(_0325_));
 sg13g2_o21ai_1 _2680_ (.B1(_1435_),
    .Y(_0331_),
    .A1(net704),
    .A2(_1170_));
 sg13g2_a21o_1 _2681_ (.A2(_0331_),
    .A1(net742),
    .B1(_1434_),
    .X(_0332_));
 sg13g2_nor2_1 _2682_ (.A(_1252_),
    .B(_1443_),
    .Y(_0333_));
 sg13g2_and2_1 _2683_ (.A(_1252_),
    .B(_1431_),
    .X(_0334_));
 sg13g2_a21oi_1 _2684_ (.A1(_1169_),
    .A2(_1350_),
    .Y(_0335_),
    .B1(net755));
 sg13g2_o21ai_1 _2685_ (.B1(_0335_),
    .Y(_0336_),
    .A1(_0333_),
    .A2(_0334_));
 sg13g2_a21oi_1 _2686_ (.A1(_1447_),
    .A2(_0336_),
    .Y(_0337_),
    .B1(net653));
 sg13g2_a21oi_1 _2687_ (.A1(_0332_),
    .A2(_0337_),
    .Y(_0338_),
    .B1(net650));
 sg13g2_o21ai_1 _2688_ (.B1(_0338_),
    .Y(_0339_),
    .A1(net656),
    .A2(_0330_));
 sg13g2_o21ai_1 _2689_ (.B1(_1454_),
    .Y(_0340_),
    .A1(net779),
    .A2(_1490_));
 sg13g2_nand3_1 _2690_ (.B(_1491_),
    .C(_0340_),
    .A(net767),
    .Y(_0341_));
 sg13g2_a21oi_2 _2691_ (.B1(_1099_),
    .Y(_0342_),
    .A2(_1456_),
    .A1(_0958_));
 sg13g2_a221oi_1 _2692_ (.B2(_1068_),
    .C1(_0342_),
    .B1(_1493_),
    .A1(_1030_),
    .Y(_0343_),
    .A2(_1234_));
 sg13g2_a21oi_1 _2693_ (.A1(_0341_),
    .A2(_0343_),
    .Y(_0344_),
    .B1(net753));
 sg13g2_a21o_1 _2694_ (.A2(_1488_),
    .A1(_1077_),
    .B1(_1122_),
    .X(_0345_));
 sg13g2_nand2_1 _2695_ (.Y(_0346_),
    .A(_1057_),
    .B(net661));
 sg13g2_nand3b_1 _2696_ (.B(_0345_),
    .C(_0346_),
    .Y(_0347_),
    .A_N(_0237_));
 sg13g2_nand2_1 _2697_ (.Y(_0348_),
    .A(_1035_),
    .B(_1263_));
 sg13g2_o21ai_1 _2698_ (.B1(_0348_),
    .Y(_0349_),
    .A1(_0972_),
    .A2(_1025_));
 sg13g2_o21ai_1 _2699_ (.B1(net703),
    .Y(_0350_),
    .A1(_1025_),
    .A2(_1159_));
 sg13g2_nand4_1 _2700_ (.B(_0133_),
    .C(_0349_),
    .A(net748),
    .Y(_0351_),
    .D(_0350_));
 sg13g2_a21oi_1 _2701_ (.A1(net689),
    .A2(_1012_),
    .Y(_0352_),
    .B1(_0122_));
 sg13g2_nor2_1 _2702_ (.A(_1252_),
    .B(_0352_),
    .Y(_0353_));
 sg13g2_o21ai_1 _2703_ (.B1(_1350_),
    .Y(_0354_),
    .A1(net680),
    .A2(_0122_));
 sg13g2_o21ai_1 _2704_ (.B1(_1175_),
    .Y(_0355_),
    .A1(net680),
    .A2(_1036_));
 sg13g2_nand3_1 _2705_ (.B(_0354_),
    .C(_0355_),
    .A(net741),
    .Y(_0356_));
 sg13g2_o21ai_1 _2706_ (.B1(_0351_),
    .Y(_0357_),
    .A1(_0353_),
    .A2(_0356_));
 sg13g2_a21oi_2 _2707_ (.B1(net654),
    .Y(_0358_),
    .A2(_0357_),
    .A1(net705));
 sg13g2_o21ai_1 _2708_ (.B1(_0358_),
    .Y(_0359_),
    .A1(_0344_),
    .A2(_0347_));
 sg13g2_a22oi_1 _2709_ (.Y(_0360_),
    .B1(net665),
    .B2(net663),
    .A2(_1091_),
    .A1(net691));
 sg13g2_nand2b_1 _2710_ (.Y(_0361_),
    .B(net812),
    .A_N(_0360_));
 sg13g2_a21oi_1 _2711_ (.A1(net802),
    .A2(_0146_),
    .Y(_0362_),
    .B1(net696));
 sg13g2_a221oi_1 _2712_ (.B2(_0362_),
    .C1(net751),
    .B1(_0361_),
    .A1(net696),
    .Y(_0363_),
    .A2(_0161_));
 sg13g2_a21oi_1 _2713_ (.A1(net691),
    .A2(_0981_),
    .Y(_0364_),
    .B1(_1040_));
 sg13g2_a21oi_1 _2714_ (.A1(_1121_),
    .A2(_0364_),
    .Y(_0365_),
    .B1(net706));
 sg13g2_o21ai_1 _2715_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_1165_),
    .A2(_0151_));
 sg13g2_or2_1 _2716_ (.X(_0367_),
    .B(_0366_),
    .A(_0363_));
 sg13g2_a21o_1 _2717_ (.A2(net663),
    .A1(net671),
    .B1(_1313_),
    .X(_0368_));
 sg13g2_a22oi_1 _2718_ (.Y(_0369_),
    .B1(_0368_),
    .B2(_0990_),
    .A2(_1446_),
    .A1(net789));
 sg13g2_nand2b_1 _2719_ (.Y(_0370_),
    .B(_1121_),
    .A_N(_0369_));
 sg13g2_o21ai_1 _2720_ (.B1(net706),
    .Y(_0371_),
    .A1(_1127_),
    .A2(_0360_));
 sg13g2_a21oi_1 _2721_ (.A1(net741),
    .A2(_1446_),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_a21oi_1 _2722_ (.A1(_0370_),
    .A2(_0372_),
    .Y(_0373_),
    .B1(net655));
 sg13g2_a21oi_1 _2723_ (.A1(_0367_),
    .A2(_0373_),
    .Y(_0374_),
    .B1(_0923_));
 sg13g2_a21oi_1 _2724_ (.A1(_0359_),
    .A2(_0374_),
    .Y(_0375_),
    .B1(_1133_));
 sg13g2_a221oi_1 _2725_ (.B2(_0375_),
    .C1(_0900_),
    .B1(_0339_),
    .A1(_0280_),
    .Y(_0376_),
    .A2(_0319_));
 sg13g2_nor2b_1 _2726_ (.A(_0376_),
    .B_N(_1288_),
    .Y(_0377_));
 sg13g2_xor2_1 _2727_ (.B(net815),
    .A(net834),
    .X(_0378_));
 sg13g2_a21oi_1 _2728_ (.A1(_0736_),
    .A2(\pix_y[8] ),
    .Y(_0379_),
    .B1(_0378_));
 sg13g2_o21ai_1 _2729_ (.B1(_0921_),
    .Y(_0380_),
    .A1(\logo_top[6] ),
    .A2(_0749_));
 sg13g2_nor4_1 _2730_ (.A(_0737_),
    .B(net816),
    .C(_0379_),
    .D(_0380_),
    .Y(_0381_));
 sg13g2_a21oi_1 _2731_ (.A1(_0737_),
    .A2(net816),
    .Y(_0382_),
    .B1(_0380_));
 sg13g2_a21oi_1 _2732_ (.A1(\logo_top[7] ),
    .A2(_0753_),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_a21oi_1 _2733_ (.A1(_0379_),
    .A2(_0383_),
    .Y(_0384_),
    .B1(_0381_));
 sg13g2_nand3_1 _2734_ (.B(net816),
    .C(_0380_),
    .A(_0737_),
    .Y(_0385_));
 sg13g2_nor2b_1 _2735_ (.A(\pix_x[7] ),
    .B_N(\logo_left[7] ),
    .Y(_0386_));
 sg13g2_nor2b_1 _2736_ (.A(net839),
    .B_N(\pix_x[7] ),
    .Y(_0387_));
 sg13g2_a21oi_1 _2737_ (.A1(_0960_),
    .A2(net726),
    .Y(_0388_),
    .B1(_0387_));
 sg13g2_nand2b_1 _2738_ (.Y(_0389_),
    .B(_0388_),
    .A_N(_0386_));
 sg13g2_nand2b_1 _2739_ (.Y(_0390_),
    .B(\logo_left[8] ),
    .A_N(\pix_x[8] ));
 sg13g2_xor2_1 _2740_ (.B(\pix_x[8] ),
    .A(\logo_left[8] ),
    .X(_0391_));
 sg13g2_a21o_1 _2741_ (.A2(_0391_),
    .A1(_0386_),
    .B1(_0387_),
    .X(_0392_));
 sg13g2_nand3_1 _2742_ (.B(net726),
    .C(_0392_),
    .A(_0960_),
    .Y(_0393_));
 sg13g2_xnor2_1 _2743_ (.Y(_0394_),
    .A(\logo_left[9] ),
    .B(\pix_x[9] ));
 sg13g2_xnor2_1 _2744_ (.Y(_0395_),
    .A(_0390_),
    .B(_0394_));
 sg13g2_nor2_1 _2745_ (.A(_0736_),
    .B(\pix_y[8] ),
    .Y(_0396_));
 sg13g2_xor2_1 _2746_ (.B(_0396_),
    .A(_0378_),
    .X(_0397_));
 sg13g2_nand2b_1 _2747_ (.Y(_0398_),
    .B(_0389_),
    .A_N(_0387_));
 sg13g2_a221oi_1 _2748_ (.B2(_0391_),
    .C1(_0397_),
    .B1(_0398_),
    .A1(_0389_),
    .Y(_0399_),
    .A2(_0393_));
 sg13g2_nand3_1 _2749_ (.B(_0395_),
    .C(_0399_),
    .A(_0385_),
    .Y(_0400_));
 sg13g2_nor2_1 _2750_ (.A(_0384_),
    .B(_0400_),
    .Y(_0401_));
 sg13g2_and2_1 _2751_ (.A(\pix_x[8] ),
    .B(\pix_x[9] ),
    .X(_0402_));
 sg13g2_nand2_1 _2752_ (.Y(_0403_),
    .A(net849),
    .B(_0779_));
 sg13g2_nor4_2 _2753_ (.A(net815),
    .B(_0774_),
    .C(_0402_),
    .Y(_0404_),
    .D(_0403_));
 sg13g2_o21ai_1 _2754_ (.B1(_0404_),
    .Y(_0405_),
    .A1(net1),
    .A2(_0401_));
 sg13g2_a221oi_1 _2755_ (.B2(_0377_),
    .C1(_0405_),
    .B1(_0233_),
    .A1(_1287_),
    .Y(_0406_),
    .A2(_1430_));
 sg13g2_nand2b_1 _2756_ (.Y(_0407_),
    .B(net713),
    .A_N(_0008_));
 sg13g2_xnor2_1 _2757_ (.Y(_0408_),
    .A(\logo_left[4] ),
    .B(net713));
 sg13g2_o21ai_1 _2758_ (.B1(_0407_),
    .Y(_0409_),
    .A1(net776),
    .A2(_0408_));
 sg13g2_nand2_1 _2759_ (.Y(_0410_),
    .A(\logo_left[5] ),
    .B(net657));
 sg13g2_xnor2_1 _2760_ (.Y(_0411_),
    .A(\logo_left[5] ),
    .B(net657));
 sg13g2_xnor2_1 _2761_ (.Y(_0412_),
    .A(net738),
    .B(_0411_));
 sg13g2_xnor2_1 _2762_ (.Y(_0413_),
    .A(net773),
    .B(_0408_));
 sg13g2_nand2_1 _2763_ (.Y(_0414_),
    .A(net841),
    .B(net755));
 sg13g2_xnor2_1 _2764_ (.Y(_0415_),
    .A(_0743_),
    .B(net744));
 sg13g2_o21ai_1 _2765_ (.B1(_0414_),
    .Y(_0416_),
    .A1(_0975_),
    .A2(_0415_));
 sg13g2_nand2_1 _2766_ (.Y(_0417_),
    .A(_0413_),
    .B(_0416_));
 sg13g2_nand2_1 _2767_ (.Y(_0418_),
    .A(_0007_),
    .B(_1288_));
 sg13g2_xnor2_1 _2768_ (.Y(_0419_),
    .A(net771),
    .B(_0415_));
 sg13g2_and2_1 _2769_ (.A(_0418_),
    .B(_0419_),
    .X(_0420_));
 sg13g2_xnor2_1 _2770_ (.Y(_0421_),
    .A(\pix_x[2] ),
    .B(_0936_));
 sg13g2_nor2_1 _2771_ (.A(net762),
    .B(_0421_),
    .Y(_0422_));
 sg13g2_xnor2_1 _2772_ (.Y(_0423_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_nor3_1 _2773_ (.A(net762),
    .B(_0421_),
    .C(_0423_),
    .Y(_0424_));
 sg13g2_xor2_1 _2774_ (.B(_0416_),
    .A(_0413_),
    .X(_0425_));
 sg13g2_o21ai_1 _2775_ (.B1(_0425_),
    .Y(_0426_),
    .A1(_0420_),
    .A2(_0424_));
 sg13g2_xnor2_1 _2776_ (.Y(_0427_),
    .A(_0409_),
    .B(_0412_));
 sg13g2_a21oi_1 _2777_ (.A1(_0417_),
    .A2(_0426_),
    .Y(_0428_),
    .B1(_0427_));
 sg13g2_a21oi_1 _2778_ (.A1(_0409_),
    .A2(_0412_),
    .Y(_0429_),
    .B1(_0428_));
 sg13g2_o21ai_1 _2779_ (.B1(_0410_),
    .Y(_0430_),
    .A1(net731),
    .A2(_0411_));
 sg13g2_xnor2_1 _2780_ (.Y(_0431_),
    .A(net840),
    .B(net689));
 sg13g2_xnor2_1 _2781_ (.Y(_0432_),
    .A(net650),
    .B(_0431_));
 sg13g2_xnor2_1 _2782_ (.Y(_0433_),
    .A(_0430_),
    .B(_0432_));
 sg13g2_xnor2_1 _2783_ (.Y(_0434_),
    .A(_0429_),
    .B(_0433_));
 sg13g2_nand2_1 _2784_ (.Y(_0435_),
    .A(net2),
    .B(net207));
 sg13g2_o21ai_1 _2785_ (.B1(_0435_),
    .Y(_0436_),
    .A1(net2),
    .A2(_0434_));
 sg13g2_and2_1 _2786_ (.A(_0406_),
    .B(_0436_),
    .X(_0022_));
 sg13g2_nand2b_1 _2787_ (.Y(_0437_),
    .B(net2),
    .A_N(net188));
 sg13g2_and2_1 _2788_ (.A(_0406_),
    .B(_0437_),
    .X(_0023_));
 sg13g2_nor2b_2 _2789_ (.A(\gamepad.driver.pmod_latch_prev ),
    .B_N(\gamepad.driver.pmod_latch_sync[1] ),
    .Y(_0438_));
 sg13g2_nor2_1 _2790_ (.A(net844),
    .B(net799),
    .Y(_0439_));
 sg13g2_a22oi_1 _2791_ (.Y(_0024_),
    .B1(net784),
    .B2(_0759_),
    .A2(net799),
    .A1(_0731_));
 sg13g2_a22oi_1 _2792_ (.Y(_0025_),
    .B1(net784),
    .B2(_0758_),
    .A2(net799),
    .A1(_0730_));
 sg13g2_a22oi_1 _2793_ (.Y(_0026_),
    .B1(net784),
    .B2(_0761_),
    .A2(net799),
    .A1(_0729_));
 sg13g2_a22oi_1 _2794_ (.Y(_0027_),
    .B1(net784),
    .B2(_0760_),
    .A2(net799),
    .A1(_0728_));
 sg13g2_a22oi_1 _2795_ (.Y(_0028_),
    .B1(net783),
    .B2(_0763_),
    .A2(net798),
    .A1(_0727_));
 sg13g2_a22oi_1 _2796_ (.Y(_0029_),
    .B1(net783),
    .B2(_0762_),
    .A2(net798),
    .A1(_0726_));
 sg13g2_a22oi_1 _2797_ (.Y(_0030_),
    .B1(net783),
    .B2(_0765_),
    .A2(net798),
    .A1(_0725_));
 sg13g2_a22oi_1 _2798_ (.Y(_0031_),
    .B1(net783),
    .B2(_0764_),
    .A2(net798),
    .A1(_0724_));
 sg13g2_a22oi_1 _2799_ (.Y(_0032_),
    .B1(net783),
    .B2(_0767_),
    .A2(net798),
    .A1(_0723_));
 sg13g2_a22oi_1 _2800_ (.Y(_0033_),
    .B1(net783),
    .B2(_0766_),
    .A2(net798),
    .A1(_0722_));
 sg13g2_a22oi_1 _2801_ (.Y(_0034_),
    .B1(net783),
    .B2(_0769_),
    .A2(net798),
    .A1(_0721_));
 sg13g2_a22oi_1 _2802_ (.Y(_0035_),
    .B1(net783),
    .B2(_0768_),
    .A2(net798),
    .A1(_0746_));
 sg13g2_nand2_1 _2803_ (.Y(_0440_),
    .A(net143),
    .B(_0799_));
 sg13g2_nand4_1 _2804_ (.B(\gamepad.decoder.data_reg[8] ),
    .C(\gamepad.decoder.data_reg[11] ),
    .A(\gamepad.decoder.data_reg[9] ),
    .Y(_0441_),
    .D(\gamepad.decoder.data_reg[10] ));
 sg13g2_nand4_1 _2805_ (.B(\gamepad.decoder.data_reg[4] ),
    .C(\gamepad.decoder.data_reg[7] ),
    .A(\gamepad.decoder.data_reg[5] ),
    .Y(_0442_),
    .D(\gamepad.decoder.data_reg[6] ));
 sg13g2_nand4_1 _2806_ (.B(\gamepad.decoder.data_reg[0] ),
    .C(\gamepad.decoder.data_reg[3] ),
    .A(\gamepad.decoder.data_reg[1] ),
    .Y(_0443_),
    .D(\gamepad.decoder.data_reg[2] ));
 sg13g2_or3_2 _2807_ (.A(_0441_),
    .B(_0442_),
    .C(_0443_),
    .X(_0444_));
 sg13g2_nand3_1 _2808_ (.B(_0800_),
    .C(_0444_),
    .A(\gamepad.decoder.data_reg[8] ),
    .Y(_0445_));
 sg13g2_a21oi_1 _2809_ (.A1(_0440_),
    .A2(_0445_),
    .Y(_0036_),
    .B1(net845));
 sg13g2_and3_1 _2810_ (.X(_0446_),
    .A(\pix_x[0] ),
    .B(net190),
    .C(net205));
 sg13g2_and2_1 _2811_ (.A(net209),
    .B(_0446_),
    .X(_0447_));
 sg13g2_and2_1 _2812_ (.A(net208),
    .B(_0447_),
    .X(_0448_));
 sg13g2_nor3_1 _2813_ (.A(\pix_x[5] ),
    .B(\pix_x[6] ),
    .C(\pix_x[7] ),
    .Y(_0449_));
 sg13g2_nand3_1 _2814_ (.B(_0448_),
    .C(_0449_),
    .A(_0402_),
    .Y(_0450_));
 sg13g2_nand2_1 _2815_ (.Y(_0451_),
    .A(net849),
    .B(_0450_));
 sg13g2_and3_1 _2816_ (.X(_0037_),
    .A(net849),
    .B(net127),
    .C(_0450_));
 sg13g2_xnor2_1 _2817_ (.Y(_0452_),
    .A(\pix_x[0] ),
    .B(net205));
 sg13g2_nor2_1 _2818_ (.A(net694),
    .B(net206),
    .Y(_0038_));
 sg13g2_a21oi_1 _2819_ (.A1(\pix_x[0] ),
    .A2(\pix_x[1] ),
    .Y(_0453_),
    .B1(net190));
 sg13g2_nor3_1 _2820_ (.A(net845),
    .B(_0446_),
    .C(net191),
    .Y(_0039_));
 sg13g2_o21ai_1 _2821_ (.B1(net849),
    .Y(_0454_),
    .A1(net209),
    .A2(_0446_));
 sg13g2_nor2_1 _2822_ (.A(_0447_),
    .B(_0454_),
    .Y(_0040_));
 sg13g2_o21ai_1 _2823_ (.B1(net849),
    .Y(_0455_),
    .A1(net208),
    .A2(_0447_));
 sg13g2_nor2_1 _2824_ (.A(_0448_),
    .B(_0455_),
    .Y(_0041_));
 sg13g2_and2_1 _2825_ (.A(net210),
    .B(_0448_),
    .X(_0456_));
 sg13g2_nor2_1 _2826_ (.A(net210),
    .B(_0448_),
    .Y(_0457_));
 sg13g2_nor3_1 _2827_ (.A(net694),
    .B(_0456_),
    .C(_0457_),
    .Y(_0042_));
 sg13g2_nor2_1 _2828_ (.A(net197),
    .B(_0456_),
    .Y(_0458_));
 sg13g2_and2_1 _2829_ (.A(_0777_),
    .B(_0447_),
    .X(_0459_));
 sg13g2_nor3_1 _2830_ (.A(net694),
    .B(net198),
    .C(_0459_),
    .Y(_0043_));
 sg13g2_xnor2_1 _2831_ (.Y(_0460_),
    .A(net202),
    .B(_0459_));
 sg13g2_nor2_1 _2832_ (.A(net694),
    .B(_0460_),
    .Y(_0044_));
 sg13g2_a21oi_1 _2833_ (.A1(net202),
    .A2(_0459_),
    .Y(_0461_),
    .B1(net199));
 sg13g2_and3_1 _2834_ (.X(_0462_),
    .A(net202),
    .B(net199),
    .C(_0459_));
 sg13g2_nor3_1 _2835_ (.A(net694),
    .B(_0461_),
    .C(_0462_),
    .Y(_0045_));
 sg13g2_a21oi_1 _2836_ (.A1(net212),
    .A2(_0462_),
    .Y(_0463_),
    .B1(net694));
 sg13g2_o21ai_1 _2837_ (.B1(_0463_),
    .Y(_0464_),
    .A1(net212),
    .A2(_0462_));
 sg13g2_inv_1 _2838_ (.Y(_0046_),
    .A(_0464_));
 sg13g2_and2_1 _2839_ (.A(\gamepad.decoder.data_reg[5] ),
    .B(_0444_),
    .X(_0465_));
 sg13g2_or2_1 _2840_ (.X(_0466_),
    .B(\logo_left[8] ),
    .A(\logo_left[9] ));
 sg13g2_o21ai_1 _2841_ (.B1(_0465_),
    .Y(_0467_),
    .A1(_0850_),
    .A2(_0466_));
 sg13g2_and3_1 _2842_ (.X(_0468_),
    .A(\gamepad.decoder.data_reg[4] ),
    .B(_0862_),
    .C(_0444_));
 sg13g2_and2_2 _2843_ (.A(_0875_),
    .B(_0468_),
    .X(_0469_));
 sg13g2_nand2_1 _2844_ (.Y(_0470_),
    .A(_0875_),
    .B(_0468_));
 sg13g2_nor2_1 _2845_ (.A(net814),
    .B(_0469_),
    .Y(_0471_));
 sg13g2_a21oi_1 _2846_ (.A1(_0467_),
    .A2(_0471_),
    .Y(_0472_),
    .B1(_0799_));
 sg13g2_a21o_2 _2847_ (.A2(_0471_),
    .A1(_0467_),
    .B1(_0799_),
    .X(_0473_));
 sg13g2_o21ai_1 _2848_ (.B1(net847),
    .Y(_0474_),
    .A1(net843),
    .A2(net648));
 sg13g2_a21oi_1 _2849_ (.A1(_0745_),
    .A2(net648),
    .Y(_0047_),
    .B1(_0474_));
 sg13g2_nand2b_1 _2850_ (.Y(_0475_),
    .B(_0856_),
    .A_N(_0836_));
 sg13g2_xnor2_1 _2851_ (.Y(_0476_),
    .A(net651),
    .B(_0475_));
 sg13g2_xor2_1 _2852_ (.B(net842),
    .A(net832),
    .X(_0477_));
 sg13g2_xnor2_1 _2853_ (.Y(_0478_),
    .A(net136),
    .B(_0477_));
 sg13g2_o21ai_1 _2854_ (.B1(net648),
    .Y(_0479_),
    .A1(net827),
    .A2(_0478_));
 sg13g2_a21oi_1 _2855_ (.A1(net827),
    .A2(_0476_),
    .Y(_0480_),
    .B1(_0479_));
 sg13g2_o21ai_1 _2856_ (.B1(net847),
    .Y(_0481_),
    .A1(net842),
    .A2(net648));
 sg13g2_nor2_1 _2857_ (.A(_0480_),
    .B(_0481_),
    .Y(_0048_));
 sg13g2_xor2_1 _2858_ (.B(_0836_),
    .A(_0007_),
    .X(_0482_));
 sg13g2_xnor2_1 _2859_ (.Y(_0483_),
    .A(\logo_left[2] ),
    .B(_0856_));
 sg13g2_o21ai_1 _2860_ (.B1(net827),
    .Y(_0484_),
    .A1(net651),
    .A2(_0483_));
 sg13g2_a21oi_1 _2861_ (.A1(net651),
    .A2(_0482_),
    .Y(_0485_),
    .B1(_0484_));
 sg13g2_xnor2_1 _2862_ (.Y(_0486_),
    .A(net832),
    .B(\logo_left[2] ));
 sg13g2_a21oi_1 _2863_ (.A1(net832),
    .A2(_0856_),
    .Y(_0487_),
    .B1(_0836_));
 sg13g2_nand2_1 _2864_ (.Y(_0488_),
    .A(_0486_),
    .B(_0487_));
 sg13g2_o21ai_1 _2865_ (.B1(net814),
    .Y(_0489_),
    .A1(_0486_),
    .A2(_0487_));
 sg13g2_nor2b_1 _2866_ (.A(_0489_),
    .B_N(_0488_),
    .Y(_0490_));
 sg13g2_nor3_1 _2867_ (.A(_0473_),
    .B(_0485_),
    .C(_0490_),
    .Y(_0491_));
 sg13g2_o21ai_1 _2868_ (.B1(net847),
    .Y(_0492_),
    .A1(net228),
    .A2(net648));
 sg13g2_nor2_1 _2869_ (.A(_0491_),
    .B(_0492_),
    .Y(_0049_));
 sg13g2_nand2_1 _2870_ (.Y(_0493_),
    .A(_0841_),
    .B(net651));
 sg13g2_o21ai_1 _2871_ (.B1(_0493_),
    .Y(_0494_),
    .A1(_0868_),
    .A2(net651));
 sg13g2_xnor2_1 _2872_ (.Y(_0495_),
    .A(net832),
    .B(net841));
 sg13g2_o21ai_1 _2873_ (.B1(_0488_),
    .Y(_0496_),
    .A1(net832),
    .A2(_0744_));
 sg13g2_xnor2_1 _2874_ (.Y(_0497_),
    .A(_0495_),
    .B(_0496_));
 sg13g2_nor2_1 _2875_ (.A(net827),
    .B(_0497_),
    .Y(_0498_));
 sg13g2_a21oi_1 _2876_ (.A1(net827),
    .A2(_0494_),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_a21oi_1 _2877_ (.A1(net841),
    .A2(_0473_),
    .Y(_0500_),
    .B1(net845));
 sg13g2_o21ai_1 _2878_ (.B1(_0500_),
    .Y(_0050_),
    .A1(_0473_),
    .A2(_0499_));
 sg13g2_a21oi_1 _2879_ (.A1(_0866_),
    .A2(_0469_),
    .Y(_0501_),
    .B1(net814));
 sg13g2_o21ai_1 _2880_ (.B1(_0501_),
    .Y(_0502_),
    .A1(_0839_),
    .A2(_0469_));
 sg13g2_xnor2_1 _2881_ (.Y(_0503_),
    .A(net832),
    .B(\logo_left[4] ));
 sg13g2_a21oi_1 _2882_ (.A1(net833),
    .A2(_0743_),
    .Y(_0504_),
    .B1(_0488_));
 sg13g2_a21oi_1 _2883_ (.A1(_0743_),
    .A2(_0744_),
    .Y(_0505_),
    .B1(net833));
 sg13g2_o21ai_1 _2884_ (.B1(_0503_),
    .Y(_0506_),
    .A1(_0504_),
    .A2(_0505_));
 sg13g2_or3_1 _2885_ (.A(_0503_),
    .B(_0504_),
    .C(_0505_),
    .X(_0507_));
 sg13g2_nand3_1 _2886_ (.B(_0506_),
    .C(_0507_),
    .A(net814),
    .Y(_0508_));
 sg13g2_nand3_1 _2887_ (.B(_0502_),
    .C(_0508_),
    .A(net648),
    .Y(_0509_));
 sg13g2_o21ai_1 _2888_ (.B1(_0509_),
    .Y(_0510_),
    .A1(net232),
    .A2(net648));
 sg13g2_nor2_1 _2889_ (.A(net845),
    .B(_0510_),
    .Y(_0051_));
 sg13g2_xor2_1 _2890_ (.B(\logo_left[5] ),
    .A(net832),
    .X(_0511_));
 sg13g2_o21ai_1 _2891_ (.B1(_0506_),
    .Y(_0512_),
    .A1(net832),
    .A2(_0742_));
 sg13g2_o21ai_1 _2892_ (.B1(net827),
    .Y(_0513_),
    .A1(_0865_),
    .A2(net651));
 sg13g2_a21oi_1 _2893_ (.A1(_0849_),
    .A2(net651),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_xor2_1 _2894_ (.B(_0512_),
    .A(_0511_),
    .X(_0515_));
 sg13g2_nor2_1 _2895_ (.A(net827),
    .B(_0515_),
    .Y(_0516_));
 sg13g2_nor3_1 _2896_ (.A(_0473_),
    .B(_0514_),
    .C(_0516_),
    .Y(_0517_));
 sg13g2_o21ai_1 _2897_ (.B1(net847),
    .Y(_0518_),
    .A1(net233),
    .A2(net648));
 sg13g2_nor2_1 _2898_ (.A(_0517_),
    .B(_0518_),
    .Y(_0052_));
 sg13g2_nand2_1 _2899_ (.Y(_0519_),
    .A(_0848_),
    .B(_0470_));
 sg13g2_a21oi_1 _2900_ (.A1(_0863_),
    .A2(_0469_),
    .Y(_0520_),
    .B1(net814));
 sg13g2_xor2_1 _2901_ (.B(net840),
    .A(dir_x),
    .X(_0521_));
 sg13g2_nor2_1 _2902_ (.A(_0506_),
    .B(_0511_),
    .Y(_0522_));
 sg13g2_nor2_1 _2903_ (.A(dir_x),
    .B(_0845_),
    .Y(_0523_));
 sg13g2_nor2_1 _2904_ (.A(_0522_),
    .B(_0523_),
    .Y(_0524_));
 sg13g2_nor2_1 _2905_ (.A(_0521_),
    .B(_0524_),
    .Y(_0525_));
 sg13g2_nand2_1 _2906_ (.Y(_0526_),
    .A(_0521_),
    .B(_0524_));
 sg13g2_nor2_1 _2907_ (.A(net827),
    .B(_0525_),
    .Y(_0527_));
 sg13g2_a22oi_1 _2908_ (.Y(_0528_),
    .B1(_0526_),
    .B2(_0527_),
    .A2(_0520_),
    .A1(_0519_));
 sg13g2_o21ai_1 _2909_ (.B1(net847),
    .Y(_0529_),
    .A1(_0473_),
    .A2(_0528_));
 sg13g2_a21o_1 _2910_ (.A2(_0473_),
    .A1(net840),
    .B1(_0529_),
    .X(_0053_));
 sg13g2_a21oi_1 _2911_ (.A1(net839),
    .A2(_0473_),
    .Y(_0530_),
    .B1(net845));
 sg13g2_xnor2_1 _2912_ (.Y(_0531_),
    .A(net833),
    .B(net839));
 sg13g2_a21oi_1 _2913_ (.A1(_0735_),
    .A2(net840),
    .Y(_0532_),
    .B1(_0525_));
 sg13g2_o21ai_1 _2914_ (.B1(net813),
    .Y(_0533_),
    .A1(_0531_),
    .A2(_0532_));
 sg13g2_a21oi_1 _2915_ (.A1(_0531_),
    .A2(_0532_),
    .Y(_0534_),
    .B1(_0533_));
 sg13g2_nor2_1 _2916_ (.A(_0873_),
    .B(_0470_),
    .Y(_0535_));
 sg13g2_o21ai_1 _2917_ (.B1(net828),
    .Y(_0536_),
    .A1(_0853_),
    .A2(_0469_));
 sg13g2_o21ai_1 _2918_ (.B1(net649),
    .Y(_0537_),
    .A1(_0535_),
    .A2(_0536_));
 sg13g2_o21ai_1 _2919_ (.B1(_0530_),
    .Y(_0054_),
    .A1(_0534_),
    .A2(_0537_));
 sg13g2_nand2_1 _2920_ (.Y(_0538_),
    .A(_0735_),
    .B(\logo_left[8] ));
 sg13g2_xor2_1 _2921_ (.B(\logo_left[8] ),
    .A(net833),
    .X(_0539_));
 sg13g2_nor3_1 _2922_ (.A(_0506_),
    .B(_0511_),
    .C(_0521_),
    .Y(_0540_));
 sg13g2_o21ai_1 _2923_ (.B1(_0735_),
    .Y(_0541_),
    .A1(net839),
    .A2(net840));
 sg13g2_nand2b_1 _2924_ (.Y(_0542_),
    .B(_0541_),
    .A_N(_0523_));
 sg13g2_a21oi_1 _2925_ (.A1(_0531_),
    .A2(_0540_),
    .Y(_0543_),
    .B1(_0542_));
 sg13g2_xor2_1 _2926_ (.B(_0543_),
    .A(_0539_),
    .X(_0544_));
 sg13g2_a22oi_1 _2927_ (.Y(_0545_),
    .B1(net651),
    .B2(_0852_),
    .A2(_0468_),
    .A1(_0874_));
 sg13g2_nand2_1 _2928_ (.Y(_0546_),
    .A(net828),
    .B(_0545_));
 sg13g2_o21ai_1 _2929_ (.B1(_0546_),
    .Y(_0547_),
    .A1(net828),
    .A2(_0544_));
 sg13g2_o21ai_1 _2930_ (.B1(net847),
    .Y(_0548_),
    .A1(net227),
    .A2(net649));
 sg13g2_a21oi_1 _2931_ (.A1(net649),
    .A2(_0547_),
    .Y(_0055_),
    .B1(_0548_));
 sg13g2_o21ai_1 _2932_ (.B1(_0538_),
    .Y(_0549_),
    .A1(_0539_),
    .A2(_0543_));
 sg13g2_xor2_1 _2933_ (.B(\logo_left[9] ),
    .A(net833),
    .X(_0550_));
 sg13g2_xnor2_1 _2934_ (.Y(_0551_),
    .A(_0549_),
    .B(_0550_));
 sg13g2_xor2_1 _2935_ (.B(_0851_),
    .A(\logo_left[9] ),
    .X(_0552_));
 sg13g2_a221oi_1 _2936_ (.B2(_0471_),
    .C1(_0473_),
    .B1(_0552_),
    .A1(net813),
    .Y(_0553_),
    .A2(_0551_));
 sg13g2_o21ai_1 _2937_ (.B1(net848),
    .Y(_0554_),
    .A1(net231),
    .A2(net649));
 sg13g2_nor2_1 _2938_ (.A(_0553_),
    .B(_0554_),
    .Y(_0056_));
 sg13g2_a21oi_1 _2939_ (.A1(_0826_),
    .A2(_0828_),
    .Y(_0555_),
    .B1(_0812_));
 sg13g2_nor2_1 _2940_ (.A(_0824_),
    .B(_0555_),
    .Y(_0556_));
 sg13g2_nand2_1 _2941_ (.Y(_0557_),
    .A(\logo_top[9] ),
    .B(\logo_top[8] ));
 sg13g2_nand3_1 _2942_ (.B(_0444_),
    .C(_0557_),
    .A(\gamepad.decoder.data_reg[6] ),
    .Y(_0558_));
 sg13g2_nor2_1 _2943_ (.A(_0833_),
    .B(_0558_),
    .Y(_0559_));
 sg13g2_o21ai_1 _2944_ (.B1(_0559_),
    .Y(_0560_),
    .A1(_0816_),
    .A2(_0556_));
 sg13g2_nand2_1 _2945_ (.Y(_0561_),
    .A(\gamepad.decoder.data_reg[7] ),
    .B(_0444_));
 sg13g2_nor2_1 _2946_ (.A(\logo_top[3] ),
    .B(net836),
    .Y(_0562_));
 sg13g2_and2_1 _2947_ (.A(_0817_),
    .B(_0562_),
    .X(_0563_));
 sg13g2_nor2_1 _2948_ (.A(net835),
    .B(\logo_top[4] ),
    .Y(_0564_));
 sg13g2_nand2_1 _2949_ (.Y(_0565_),
    .A(_0563_),
    .B(_0564_));
 sg13g2_nor3_2 _2950_ (.A(\logo_top[7] ),
    .B(\logo_top[6] ),
    .C(_0565_),
    .Y(_0566_));
 sg13g2_inv_1 _2951_ (.Y(_0567_),
    .A(_0566_));
 sg13g2_nor3_1 _2952_ (.A(net834),
    .B(\logo_top[8] ),
    .C(_0567_),
    .Y(_0568_));
 sg13g2_o21ai_1 _2953_ (.B1(net826),
    .Y(_0569_),
    .A1(_0561_),
    .A2(_0568_));
 sg13g2_inv_1 _2954_ (.Y(_0570_),
    .A(_0569_));
 sg13g2_a21oi_1 _2955_ (.A1(net646),
    .A2(_0570_),
    .Y(_0571_),
    .B1(_0799_));
 sg13g2_o21ai_1 _2956_ (.B1(net846),
    .Y(_0572_),
    .A1(net838),
    .A2(net642));
 sg13g2_a21oi_1 _2957_ (.A1(_0740_),
    .A2(net642),
    .Y(_0057_),
    .B1(_0572_));
 sg13g2_xnor2_1 _2958_ (.Y(_0573_),
    .A(net837),
    .B(net838));
 sg13g2_xnor2_1 _2959_ (.Y(_0574_),
    .A(net647),
    .B(_0573_));
 sg13g2_xor2_1 _2960_ (.B(net837),
    .A(net830),
    .X(_0575_));
 sg13g2_xnor2_1 _2961_ (.Y(_0576_),
    .A(net132),
    .B(_0575_));
 sg13g2_o21ai_1 _2962_ (.B1(net642),
    .Y(_0577_),
    .A1(net825),
    .A2(_0576_));
 sg13g2_a21oi_1 _2963_ (.A1(net825),
    .A2(_0574_),
    .Y(_0578_),
    .B1(_0577_));
 sg13g2_o21ai_1 _2964_ (.B1(net846),
    .Y(_0579_),
    .A1(net837),
    .A2(net642));
 sg13g2_nor2_1 _2965_ (.A(_0578_),
    .B(_0579_),
    .Y(_0058_));
 sg13g2_xnor2_1 _2966_ (.Y(_0580_),
    .A(net836),
    .B(_0803_));
 sg13g2_xnor2_1 _2967_ (.Y(_0581_),
    .A(_0771_),
    .B(_0817_));
 sg13g2_o21ai_1 _2968_ (.B1(net825),
    .Y(_0582_),
    .A1(net647),
    .A2(_0580_));
 sg13g2_a21oi_1 _2969_ (.A1(net647),
    .A2(_0581_),
    .Y(_0583_),
    .B1(_0582_));
 sg13g2_xnor2_1 _2970_ (.Y(_0584_),
    .A(net830),
    .B(net836));
 sg13g2_a21oi_1 _2971_ (.A1(net830),
    .A2(_0803_),
    .Y(_0585_),
    .B1(_0817_));
 sg13g2_and2_1 _2972_ (.A(_0584_),
    .B(_0585_),
    .X(_0586_));
 sg13g2_o21ai_1 _2973_ (.B1(net813),
    .Y(_0587_),
    .A1(_0584_),
    .A2(_0585_));
 sg13g2_o21ai_1 _2974_ (.B1(net644),
    .Y(_0588_),
    .A1(_0586_),
    .A2(_0587_));
 sg13g2_nor2_1 _2975_ (.A(net836),
    .B(net642),
    .Y(_0589_));
 sg13g2_o21ai_1 _2976_ (.B1(net846),
    .Y(_0590_),
    .A1(_0583_),
    .A2(_0588_));
 sg13g2_nor2_1 _2977_ (.A(_0589_),
    .B(_0590_),
    .Y(_0059_));
 sg13g2_nor2_1 _2978_ (.A(_0831_),
    .B(net647),
    .Y(_0591_));
 sg13g2_a21oi_1 _2979_ (.A1(_0819_),
    .A2(net647),
    .Y(_0592_),
    .B1(_0591_));
 sg13g2_xor2_1 _2980_ (.B(\logo_top[3] ),
    .A(net830),
    .X(_0593_));
 sg13g2_a21oi_1 _2981_ (.A1(_0734_),
    .A2(net836),
    .Y(_0594_),
    .B1(_0586_));
 sg13g2_xnor2_1 _2982_ (.Y(_0595_),
    .A(_0593_),
    .B(_0594_));
 sg13g2_nor2_1 _2983_ (.A(net230),
    .B(net642),
    .Y(_0596_));
 sg13g2_o21ai_1 _2984_ (.B1(net642),
    .Y(_0597_),
    .A1(net825),
    .A2(_0595_));
 sg13g2_a21oi_1 _2985_ (.A1(net825),
    .A2(_0592_),
    .Y(_0598_),
    .B1(_0597_));
 sg13g2_o21ai_1 _2986_ (.B1(net846),
    .Y(_0060_),
    .A1(_0596_),
    .A2(_0598_));
 sg13g2_nand2_1 _2987_ (.Y(_0599_),
    .A(_0012_),
    .B(_0563_));
 sg13g2_xor2_1 _2988_ (.B(_0563_),
    .A(_0012_),
    .X(_0600_));
 sg13g2_nor2_1 _2989_ (.A(_0829_),
    .B(net645),
    .Y(_0601_));
 sg13g2_a21oi_1 _2990_ (.A1(net645),
    .A2(_0600_),
    .Y(_0602_),
    .B1(_0601_));
 sg13g2_xnor2_1 _2991_ (.Y(_0603_),
    .A(net830),
    .B(\logo_top[4] ));
 sg13g2_o21ai_1 _2992_ (.B1(_0586_),
    .Y(_0604_),
    .A1(_0734_),
    .A2(\logo_top[3] ));
 sg13g2_o21ai_1 _2993_ (.B1(_0604_),
    .Y(_0605_),
    .A1(net830),
    .A2(_0562_));
 sg13g2_nand2_1 _2994_ (.Y(_0606_),
    .A(_0603_),
    .B(_0605_));
 sg13g2_xnor2_1 _2995_ (.Y(_0607_),
    .A(_0603_),
    .B(_0605_));
 sg13g2_o21ai_1 _2996_ (.B1(net643),
    .Y(_0608_),
    .A1(net825),
    .A2(_0607_));
 sg13g2_a21oi_1 _2997_ (.A1(net825),
    .A2(_0602_),
    .Y(_0609_),
    .B1(_0608_));
 sg13g2_o21ai_1 _2998_ (.B1(net846),
    .Y(_0610_),
    .A1(net223),
    .A2(net644));
 sg13g2_nor2_1 _2999_ (.A(_0609_),
    .B(_0610_),
    .Y(_0061_));
 sg13g2_xor2_1 _3000_ (.B(_0599_),
    .A(net835),
    .X(_0611_));
 sg13g2_o21ai_1 _3001_ (.B1(_0606_),
    .Y(_0612_),
    .A1(net830),
    .A2(_0738_));
 sg13g2_xnor2_1 _3002_ (.Y(_0613_),
    .A(net830),
    .B(\logo_top[5] ));
 sg13g2_xnor2_1 _3003_ (.Y(_0614_),
    .A(_0612_),
    .B(_0613_));
 sg13g2_o21ai_1 _3004_ (.B1(net643),
    .Y(_0615_),
    .A1(net825),
    .A2(_0614_));
 sg13g2_nand2b_1 _3005_ (.Y(_0616_),
    .B(_0828_),
    .A_N(net645));
 sg13g2_a21oi_1 _3006_ (.A1(net645),
    .A2(_0611_),
    .Y(_0617_),
    .B1(net813));
 sg13g2_a21oi_1 _3007_ (.A1(_0616_),
    .A2(_0617_),
    .Y(_0618_),
    .B1(_0615_));
 sg13g2_o21ai_1 _3008_ (.B1(net846),
    .Y(_0619_),
    .A1(net835),
    .A2(net642));
 sg13g2_nor2_1 _3009_ (.A(_0618_),
    .B(_0619_),
    .Y(_0062_));
 sg13g2_nand3_1 _3010_ (.B(_0563_),
    .C(_0564_),
    .A(_0013_),
    .Y(_0620_));
 sg13g2_xnor2_1 _3011_ (.Y(_0621_),
    .A(_0013_),
    .B(_0565_));
 sg13g2_nor2_1 _3012_ (.A(_0809_),
    .B(net645),
    .Y(_0622_));
 sg13g2_a21oi_1 _3013_ (.A1(net646),
    .A2(_0621_),
    .Y(_0623_),
    .B1(_0622_));
 sg13g2_xor2_1 _3014_ (.B(\logo_top[6] ),
    .A(net831),
    .X(_0624_));
 sg13g2_or2_1 _3015_ (.X(_0625_),
    .B(_0564_),
    .A(net831));
 sg13g2_nand3_1 _3016_ (.B(_0605_),
    .C(_0613_),
    .A(_0603_),
    .Y(_0626_));
 sg13g2_nand3_1 _3017_ (.B(_0625_),
    .C(_0626_),
    .A(_0624_),
    .Y(_0627_));
 sg13g2_a21oi_1 _3018_ (.A1(_0625_),
    .A2(_0626_),
    .Y(_0628_),
    .B1(_0624_));
 sg13g2_nand2_1 _3019_ (.Y(_0629_),
    .A(net813),
    .B(_0627_));
 sg13g2_o21ai_1 _3020_ (.B1(net643),
    .Y(_0630_),
    .A1(_0628_),
    .A2(_0629_));
 sg13g2_a21oi_1 _3021_ (.A1(net826),
    .A2(_0623_),
    .Y(_0631_),
    .B1(_0630_));
 sg13g2_nor2_1 _3022_ (.A(\logo_top[6] ),
    .B(net643),
    .Y(_0632_));
 sg13g2_o21ai_1 _3023_ (.B1(net848),
    .Y(_0063_),
    .A1(_0631_),
    .A2(_0632_));
 sg13g2_xnor2_1 _3024_ (.Y(_0633_),
    .A(_0737_),
    .B(_0620_));
 sg13g2_o21ai_1 _3025_ (.B1(net826),
    .Y(_0634_),
    .A1(_0811_),
    .A2(net645));
 sg13g2_a21oi_1 _3026_ (.A1(net645),
    .A2(_0633_),
    .Y(_0635_),
    .B1(_0634_));
 sg13g2_xor2_1 _3027_ (.B(\logo_top[7] ),
    .A(net831),
    .X(_0636_));
 sg13g2_a21o_1 _3028_ (.A2(\logo_top[6] ),
    .A1(_0734_),
    .B1(_0628_),
    .X(_0637_));
 sg13g2_xor2_1 _3029_ (.B(_0637_),
    .A(_0636_),
    .X(_0638_));
 sg13g2_o21ai_1 _3030_ (.B1(net644),
    .Y(_0639_),
    .A1(net826),
    .A2(_0638_));
 sg13g2_nor2_1 _3031_ (.A(_0635_),
    .B(_0639_),
    .Y(_0640_));
 sg13g2_nor2_1 _3032_ (.A(\logo_top[7] ),
    .B(net644),
    .Y(_0641_));
 sg13g2_o21ai_1 _3033_ (.B1(net848),
    .Y(_0064_),
    .A1(_0640_),
    .A2(_0641_));
 sg13g2_nand2_1 _3034_ (.Y(_0642_),
    .A(_0014_),
    .B(_0566_));
 sg13g2_xnor2_1 _3035_ (.Y(_0643_),
    .A(_0014_),
    .B(_0566_));
 sg13g2_mux2_1 _3036_ (.A0(_0823_),
    .A1(_0643_),
    .S(net645),
    .X(_0644_));
 sg13g2_nand2_1 _3037_ (.Y(_0645_),
    .A(_0734_),
    .B(\logo_top[8] ));
 sg13g2_xnor2_1 _3038_ (.Y(_0646_),
    .A(dir_y),
    .B(\logo_top[8] ));
 sg13g2_nor3_1 _3039_ (.A(_0624_),
    .B(_0626_),
    .C(_0636_),
    .Y(_0647_));
 sg13g2_o21ai_1 _3040_ (.B1(_0734_),
    .Y(_0648_),
    .A1(\logo_top[7] ),
    .A2(\logo_top[6] ));
 sg13g2_nand2_1 _3041_ (.Y(_0649_),
    .A(_0625_),
    .B(_0648_));
 sg13g2_o21ai_1 _3042_ (.B1(_0646_),
    .Y(_0650_),
    .A1(_0647_),
    .A2(_0649_));
 sg13g2_or3_1 _3043_ (.A(_0646_),
    .B(_0647_),
    .C(_0649_),
    .X(_0651_));
 sg13g2_nand3_1 _3044_ (.B(_0650_),
    .C(_0651_),
    .A(net813),
    .Y(_0652_));
 sg13g2_nand2_1 _3045_ (.Y(_0653_),
    .A(net643),
    .B(_0652_));
 sg13g2_a21oi_1 _3046_ (.A1(net826),
    .A2(_0644_),
    .Y(_0654_),
    .B1(_0653_));
 sg13g2_o21ai_1 _3047_ (.B1(net846),
    .Y(_0655_),
    .A1(net224),
    .A2(net643));
 sg13g2_nor2_1 _3048_ (.A(_0654_),
    .B(_0655_),
    .Y(_0065_));
 sg13g2_xor2_1 _3049_ (.B(net834),
    .A(dir_y),
    .X(_0656_));
 sg13g2_nand3_1 _3050_ (.B(_0650_),
    .C(_0656_),
    .A(_0645_),
    .Y(_0657_));
 sg13g2_a21o_1 _3051_ (.A2(_0650_),
    .A1(_0645_),
    .B1(_0656_),
    .X(_0658_));
 sg13g2_nand3_1 _3052_ (.B(_0657_),
    .C(_0658_),
    .A(net813),
    .Y(_0659_));
 sg13g2_xnor2_1 _3053_ (.Y(_0660_),
    .A(net834),
    .B(_0642_));
 sg13g2_nand3_1 _3054_ (.B(net646),
    .C(_0660_),
    .A(net826),
    .Y(_0661_));
 sg13g2_nand3_1 _3055_ (.B(_0659_),
    .C(_0661_),
    .A(net643),
    .Y(_0662_));
 sg13g2_o21ai_1 _3056_ (.B1(net848),
    .Y(_0663_),
    .A1(net834),
    .A2(net643));
 sg13g2_nor2b_1 _3057_ (.A(_0663_),
    .B_N(_0662_),
    .Y(_0066_));
 sg13g2_o21ai_1 _3058_ (.B1(_0444_),
    .Y(_0664_),
    .A1(\gamepad.decoder.data_reg[5] ),
    .A2(\gamepad.decoder.data_reg[4] ));
 sg13g2_nand3_1 _3059_ (.B(_0877_),
    .C(_0664_),
    .A(_0855_),
    .Y(_0665_));
 sg13g2_a21o_1 _3060_ (.A2(_0665_),
    .A1(_0801_),
    .B1(_0735_),
    .X(_0666_));
 sg13g2_nand2_1 _3061_ (.Y(_0667_),
    .A(_0855_),
    .B(_0465_));
 sg13g2_nand4_1 _3062_ (.B(_0877_),
    .C(_0665_),
    .A(_0801_),
    .Y(_0668_),
    .D(_0667_));
 sg13g2_nand3_1 _3063_ (.B(_0666_),
    .C(_0668_),
    .A(net847),
    .Y(_0067_));
 sg13g2_o21ai_1 _3064_ (.B1(_0444_),
    .Y(_0669_),
    .A1(\gamepad.decoder.data_reg[7] ),
    .A2(\gamepad.decoder.data_reg[6] ));
 sg13g2_a21oi_1 _3065_ (.A1(_0835_),
    .A2(_0669_),
    .Y(_0670_),
    .B1(_0802_));
 sg13g2_nand2b_1 _3066_ (.Y(_0671_),
    .B(_0822_),
    .A_N(_0561_));
 sg13g2_nand2_1 _3067_ (.Y(_0672_),
    .A(_0834_),
    .B(_0671_));
 sg13g2_o21ai_1 _3068_ (.B1(net846),
    .Y(_0673_),
    .A1(net831),
    .A2(_0670_));
 sg13g2_a21oi_1 _3069_ (.A1(_0670_),
    .A2(_0672_),
    .Y(_0068_),
    .B1(_0673_));
 sg13g2_or2_1 _3070_ (.X(_0674_),
    .B(_0445_),
    .A(gamepad_start_prev));
 sg13g2_o21ai_1 _3071_ (.B1(net847),
    .Y(_0675_),
    .A1(net138),
    .A2(_0674_));
 sg13g2_a21oi_1 _3072_ (.A1(net813),
    .A2(_0674_),
    .Y(_0069_),
    .B1(net139));
 sg13g2_nand2_1 _3073_ (.Y(_0676_),
    .A(\color_index[0] ),
    .B(_0879_));
 sg13g2_nand2_1 _3074_ (.Y(_0677_),
    .A(net134),
    .B(_0880_));
 sg13g2_a21oi_1 _3075_ (.A1(_0676_),
    .A2(_0677_),
    .Y(_0070_),
    .B1(net844));
 sg13g2_nand2_1 _3076_ (.Y(_0678_),
    .A(net173),
    .B(_0879_));
 sg13g2_o21ai_1 _3077_ (.B1(net850),
    .Y(_0679_),
    .A1(net173),
    .A2(\color_index[0] ));
 sg13g2_a21oi_1 _3078_ (.A1(_0890_),
    .A2(_0678_),
    .Y(_0071_),
    .B1(_0679_));
 sg13g2_nand2_1 _3079_ (.Y(_0680_),
    .A(net141),
    .B(_0879_));
 sg13g2_a21oi_1 _3080_ (.A1(_0886_),
    .A2(_0680_),
    .Y(_0072_),
    .B1(net844));
 sg13g2_and2_1 _3081_ (.A(net824),
    .B(net849),
    .X(_0073_));
 sg13g2_and2_1 _3082_ (.A(net823),
    .B(net849),
    .X(_0074_));
 sg13g2_and2_1 _3083_ (.A(net822),
    .B(net852),
    .X(_0075_));
 sg13g2_and2_1 _3084_ (.A(net820),
    .B(net852),
    .X(_0076_));
 sg13g2_and2_1 _3085_ (.A(net819),
    .B(net851),
    .X(_0077_));
 sg13g2_nor2_1 _3086_ (.A(_0748_),
    .B(net844),
    .Y(_0078_));
 sg13g2_nor2_1 _3087_ (.A(_0749_),
    .B(net845),
    .Y(_0079_));
 sg13g2_nor2_1 _3088_ (.A(net844),
    .B(_0753_),
    .Y(_0080_));
 sg13g2_nor2_1 _3089_ (.A(net844),
    .B(_0751_),
    .Y(_0081_));
 sg13g2_nor2_1 _3090_ (.A(net844),
    .B(_0752_),
    .Y(_0082_));
 sg13g2_xnor2_1 _3091_ (.Y(_0681_),
    .A(net762),
    .B(_0421_));
 sg13g2_nand2_1 _3092_ (.Y(_0682_),
    .A(net201),
    .B(net2));
 sg13g2_o21ai_1 _3093_ (.B1(_0682_),
    .Y(_0683_),
    .A1(net2),
    .A2(_0681_));
 sg13g2_and2_1 _3094_ (.A(_0406_),
    .B(_0683_),
    .X(_0083_));
 sg13g2_xnor2_1 _3095_ (.Y(_0684_),
    .A(_0422_),
    .B(_0423_));
 sg13g2_mux2_1 _3096_ (.A0(net204),
    .A1(_0684_),
    .S(_0772_),
    .X(_0685_));
 sg13g2_and2_1 _3097_ (.A(_0406_),
    .B(_0685_),
    .X(_0084_));
 sg13g2_nor3_1 _3098_ (.A(_0420_),
    .B(_0424_),
    .C(_0425_),
    .Y(_0686_));
 sg13g2_nand2_1 _3099_ (.Y(_0687_),
    .A(_0772_),
    .B(_0426_));
 sg13g2_nand2_1 _3100_ (.Y(_0688_),
    .A(net2),
    .B(net195));
 sg13g2_o21ai_1 _3101_ (.B1(_0688_),
    .Y(_0689_),
    .A1(_0686_),
    .A2(_0687_));
 sg13g2_and2_1 _3102_ (.A(_0406_),
    .B(_0689_),
    .X(_0085_));
 sg13g2_nand2b_1 _3103_ (.Y(_0690_),
    .B(net2),
    .A_N(net196));
 sg13g2_and3_1 _3104_ (.X(_0691_),
    .A(_0417_),
    .B(_0426_),
    .C(_0427_));
 sg13g2_o21ai_1 _3105_ (.B1(_0772_),
    .Y(_0692_),
    .A1(_0428_),
    .A2(_0691_));
 sg13g2_and3_1 _3106_ (.X(_0086_),
    .A(_0406_),
    .B(_0690_),
    .C(_0692_));
 sg13g2_nor2b_2 _3107_ (.A(\gamepad.driver.pmod_clk_prev ),
    .B_N(\gamepad.driver.pmod_clk_sync[1] ),
    .Y(_0693_));
 sg13g2_nor2_1 _3108_ (.A(net844),
    .B(net797),
    .Y(_0694_));
 sg13g2_a22oi_1 _3109_ (.Y(_0087_),
    .B1(net782),
    .B2(_0731_),
    .A2(net797),
    .A1(_0732_));
 sg13g2_a22oi_1 _3110_ (.Y(_0088_),
    .B1(net782),
    .B2(_0730_),
    .A2(net797),
    .A1(_0731_));
 sg13g2_a22oi_1 _3111_ (.Y(_0089_),
    .B1(net782),
    .B2(_0729_),
    .A2(net797),
    .A1(_0730_));
 sg13g2_a22oi_1 _3112_ (.Y(_0090_),
    .B1(net782),
    .B2(_0728_),
    .A2(net797),
    .A1(_0729_));
 sg13g2_a22oi_1 _3113_ (.Y(_0091_),
    .B1(net781),
    .B2(_0727_),
    .A2(net796),
    .A1(_0728_));
 sg13g2_a22oi_1 _3114_ (.Y(_0092_),
    .B1(net781),
    .B2(_0726_),
    .A2(net796),
    .A1(_0727_));
 sg13g2_a22oi_1 _3115_ (.Y(_0093_),
    .B1(net781),
    .B2(_0725_),
    .A2(net796),
    .A1(_0726_));
 sg13g2_a22oi_1 _3116_ (.Y(_0094_),
    .B1(net781),
    .B2(_0724_),
    .A2(net796),
    .A1(_0725_));
 sg13g2_a22oi_1 _3117_ (.Y(_0095_),
    .B1(net781),
    .B2(_0723_),
    .A2(net796),
    .A1(_0724_));
 sg13g2_a22oi_1 _3118_ (.Y(_0096_),
    .B1(net781),
    .B2(_0722_),
    .A2(net796),
    .A1(_0723_));
 sg13g2_a22oi_1 _3119_ (.Y(_0097_),
    .B1(net781),
    .B2(_0721_),
    .A2(net796),
    .A1(_0722_));
 sg13g2_a22oi_1 _3120_ (.Y(_0098_),
    .B1(net781),
    .B2(_0746_),
    .A2(net796),
    .A1(_0721_));
 sg13g2_and2_1 _3121_ (.A(net851),
    .B(net5),
    .X(_0099_));
 sg13g2_and2_1 _3122_ (.A(net851),
    .B(net129),
    .X(_0100_));
 sg13g2_and2_1 _3123_ (.A(net851),
    .B(net4),
    .X(_0101_));
 sg13g2_and2_1 _3124_ (.A(net850),
    .B(net131),
    .X(_0102_));
 sg13g2_and2_1 _3125_ (.A(net850),
    .B(net3),
    .X(_0103_));
 sg13g2_and2_1 _3126_ (.A(net850),
    .B(net130),
    .X(_0104_));
 sg13g2_nand3_1 _3127_ (.B(_0751_),
    .C(_0797_),
    .A(net822),
    .Y(_0695_));
 sg13g2_nand3_1 _3128_ (.B(net815),
    .C(_0796_),
    .A(net820),
    .Y(_0696_));
 sg13g2_o21ai_1 _3129_ (.B1(net849),
    .Y(_0697_),
    .A1(_0695_),
    .A2(_0696_));
 sg13g2_nor2_1 _3130_ (.A(_0450_),
    .B(_0697_),
    .Y(_0698_));
 sg13g2_a22oi_1 _3131_ (.Y(_0699_),
    .B1(_0698_),
    .B2(net128),
    .A2(_0073_),
    .A1(_0450_));
 sg13g2_inv_1 _3132_ (.Y(_0105_),
    .A(_0699_));
 sg13g2_and3_1 _3133_ (.X(_0700_),
    .A(net824),
    .B(net823),
    .C(_0451_));
 sg13g2_a21oi_1 _3134_ (.A1(net824),
    .A2(_0451_),
    .Y(_0701_),
    .B1(net823));
 sg13g2_and2_2 _3135_ (.A(net694),
    .B(_0697_),
    .X(_0702_));
 sg13g2_nand2_1 _3136_ (.Y(_0703_),
    .A(net694),
    .B(_0697_));
 sg13g2_nor3_1 _3137_ (.A(_0700_),
    .B(_0701_),
    .C(_0702_),
    .Y(_0106_));
 sg13g2_nand2_1 _3138_ (.Y(_0704_),
    .A(net822),
    .B(_0700_));
 sg13g2_inv_1 _3139_ (.Y(_0705_),
    .A(_0704_));
 sg13g2_nor2_1 _3140_ (.A(_0702_),
    .B(_0705_),
    .Y(_0706_));
 sg13g2_o21ai_1 _3141_ (.B1(_0706_),
    .Y(_0707_),
    .A1(net822),
    .A2(_0700_));
 sg13g2_inv_1 _3142_ (.Y(_0107_),
    .A(_0707_));
 sg13g2_nand2_1 _3143_ (.Y(_0708_),
    .A(net820),
    .B(_0706_));
 sg13g2_nand4_1 _3144_ (.B(net823),
    .C(net822),
    .A(net824),
    .Y(_0709_),
    .D(_0698_));
 sg13g2_o21ai_1 _3145_ (.B1(_0708_),
    .Y(_0108_),
    .A1(net820),
    .A2(_0709_));
 sg13g2_and3_2 _3146_ (.X(_0710_),
    .A(net820),
    .B(net819),
    .C(_0705_));
 sg13g2_a21oi_1 _3147_ (.A1(net820),
    .A2(_0705_),
    .Y(_0711_),
    .B1(net819));
 sg13g2_nor3_1 _3148_ (.A(_0702_),
    .B(_0710_),
    .C(_0711_),
    .Y(_0109_));
 sg13g2_nand3b_1 _3149_ (.B(net817),
    .C(_0703_),
    .Y(_0712_),
    .A_N(_0710_));
 sg13g2_nand2b_1 _3150_ (.Y(_0713_),
    .B(_0710_),
    .A_N(_0697_));
 sg13g2_o21ai_1 _3151_ (.B1(_0712_),
    .Y(_0110_),
    .A1(net817),
    .A2(_0713_));
 sg13g2_nor2b_1 _3152_ (.A(_0773_),
    .B_N(_0710_),
    .Y(_0714_));
 sg13g2_a21oi_1 _3153_ (.A1(net817),
    .A2(_0710_),
    .Y(_0715_),
    .B1(net213));
 sg13g2_nor3_1 _3154_ (.A(_0702_),
    .B(_0714_),
    .C(_0715_),
    .Y(_0111_));
 sg13g2_nor3_1 _3155_ (.A(net203),
    .B(_0773_),
    .C(_0713_),
    .Y(_0716_));
 sg13g2_nand3b_1 _3156_ (.B(net816),
    .C(_0703_),
    .Y(_0717_),
    .A_N(_0714_));
 sg13g2_nand2b_1 _3157_ (.Y(_0112_),
    .B(_0717_),
    .A_N(_0716_));
 sg13g2_a21oi_1 _3158_ (.A1(_0774_),
    .A2(_0710_),
    .Y(_0718_),
    .B1(_0702_));
 sg13g2_nand4_1 _3159_ (.B(net213),
    .C(net816),
    .A(net817),
    .Y(_0719_),
    .D(_0710_));
 sg13g2_a221oi_1 _3160_ (.B2(_0751_),
    .C1(_0702_),
    .B1(_0719_),
    .A1(_0774_),
    .Y(_0113_),
    .A2(_0710_));
 sg13g2_nor3_1 _3161_ (.A(net815),
    .B(_0775_),
    .C(_0713_),
    .Y(_0720_));
 sg13g2_a21o_1 _3162_ (.A2(_0718_),
    .A1(net815),
    .B1(_0720_),
    .X(_0114_));
 sg13g2_a21o_1 _3163_ (.A2(_0891_),
    .A1(net850),
    .B1(_0115_),
    .X(_0116_));
 sg13g2_dfrbp_1 _3164_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net87),
    .D(_0022_),
    .Q_N(_1573_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _3165_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net40),
    .D(_0023_),
    .Q_N(_1572_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _3166_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net39),
    .D(net157),
    .Q_N(_1571_),
    .Q(\gamepad.decoder.data_reg[0] ));
 sg13g2_dfrbp_1 _3167_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net37),
    .D(net161),
    .Q_N(_1570_),
    .Q(\gamepad.decoder.data_reg[1] ));
 sg13g2_dfrbp_1 _3168_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net35),
    .D(net148),
    .Q_N(_1569_),
    .Q(\gamepad.decoder.data_reg[2] ));
 sg13g2_dfrbp_1 _3169_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net33),
    .D(net159),
    .Q_N(_1568_),
    .Q(\gamepad.decoder.data_reg[3] ));
 sg13g2_dfrbp_1 _3170_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net31),
    .D(_0028_),
    .Q_N(_1567_),
    .Q(\gamepad.decoder.data_reg[4] ));
 sg13g2_dfrbp_1 _3171_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net29),
    .D(net168),
    .Q_N(_1566_),
    .Q(\gamepad.decoder.data_reg[5] ));
 sg13g2_dfrbp_1 _3172_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net27),
    .D(_0030_),
    .Q_N(_1565_),
    .Q(\gamepad.decoder.data_reg[6] ));
 sg13g2_dfrbp_1 _3173_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net25),
    .D(_0031_),
    .Q_N(_1564_),
    .Q(\gamepad.decoder.data_reg[7] ));
 sg13g2_dfrbp_1 _3174_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net23),
    .D(_0032_),
    .Q_N(_1563_),
    .Q(\gamepad.decoder.data_reg[8] ));
 sg13g2_dfrbp_1 _3175_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net124),
    .D(net146),
    .Q_N(_1562_),
    .Q(\gamepad.decoder.data_reg[9] ));
 sg13g2_dfrbp_1 _3176_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net117),
    .D(net152),
    .Q_N(_1561_),
    .Q(\gamepad.decoder.data_reg[10] ));
 sg13g2_dfrbp_1 _3177_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net115),
    .D(_0035_),
    .Q_N(_1560_),
    .Q(\gamepad.decoder.data_reg[11] ));
 sg13g2_dfrbp_1 _3178_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net113),
    .D(net144),
    .Q_N(_1559_),
    .Q(gamepad_start_prev));
 sg13g2_dfrbp_1 _3179_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net111),
    .D(_0037_),
    .Q_N(_0021_),
    .Q(\pix_x[0] ));
 sg13g2_dfrbp_1 _3180_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net110),
    .D(_0038_),
    .Q_N(_1558_),
    .Q(\pix_x[1] ));
 sg13g2_dfrbp_1 _3181_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net109),
    .D(net192),
    .Q_N(_1557_),
    .Q(\pix_x[2] ));
 sg13g2_dfrbp_1 _3182_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net108),
    .D(_0040_),
    .Q_N(_1556_),
    .Q(\pix_x[3] ));
 sg13g2_dfrbp_1 _3183_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net106),
    .D(_0041_),
    .Q_N(_1555_),
    .Q(\pix_x[4] ));
 sg13g2_dfrbp_1 _3184_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net105),
    .D(_0042_),
    .Q_N(_1554_),
    .Q(\pix_x[5] ));
 sg13g2_dfrbp_1 _3185_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net104),
    .D(_0043_),
    .Q_N(_1553_),
    .Q(\pix_x[6] ));
 sg13g2_dfrbp_1 _3186_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net103),
    .D(_0044_),
    .Q_N(_1552_),
    .Q(\pix_x[7] ));
 sg13g2_dfrbp_1 _3187_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net102),
    .D(_0045_),
    .Q_N(_1551_),
    .Q(\pix_x[8] ));
 sg13g2_dfrbp_1 _3188_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net101),
    .D(_0046_),
    .Q_N(_1550_),
    .Q(\pix_x[9] ));
 sg13g2_dfrbp_1 _3189_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net100),
    .D(net137),
    .Q_N(_0020_),
    .Q(\logo_left[0] ));
 sg13g2_dfrbp_1 _3190_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net98),
    .D(_0048_),
    .Q_N(_1549_),
    .Q(\logo_left[1] ));
 sg13g2_dfrbp_1 _3191_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net96),
    .D(_0049_),
    .Q_N(_0007_),
    .Q(\logo_left[2] ));
 sg13g2_dfrbp_1 _3192_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net94),
    .D(_0050_),
    .Q_N(_1548_),
    .Q(\logo_left[3] ));
 sg13g2_dfrbp_1 _3193_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net92),
    .D(_0051_),
    .Q_N(_0008_),
    .Q(\logo_left[4] ));
 sg13g2_dfrbp_1 _3194_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net90),
    .D(_0052_),
    .Q_N(_1547_),
    .Q(\logo_left[5] ));
 sg13g2_dfrbp_1 _3195_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net86),
    .D(_0053_),
    .Q_N(_0009_),
    .Q(\logo_left[6] ));
 sg13g2_dfrbp_1 _3196_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net84),
    .D(_0054_),
    .Q_N(_1546_),
    .Q(\logo_left[7] ));
 sg13g2_dfrbp_1 _3197_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net82),
    .D(_0055_),
    .Q_N(_0010_),
    .Q(\logo_left[8] ));
 sg13g2_dfrbp_1 _3198_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net80),
    .D(_0056_),
    .Q_N(_1545_),
    .Q(\logo_left[9] ));
 sg13g2_dfrbp_1 _3199_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net78),
    .D(net133),
    .Q_N(_0019_),
    .Q(\logo_top[0] ));
 sg13g2_dfrbp_1 _3200_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net76),
    .D(_0058_),
    .Q_N(_1544_),
    .Q(\logo_top[1] ));
 sg13g2_dfrbp_1 _3201_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net74),
    .D(_0059_),
    .Q_N(_0011_),
    .Q(\logo_top[2] ));
 sg13g2_dfrbp_1 _3202_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net72),
    .D(_0060_),
    .Q_N(_1543_),
    .Q(\logo_top[3] ));
 sg13g2_dfrbp_1 _3203_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net70),
    .D(_0061_),
    .Q_N(_0012_),
    .Q(\logo_top[4] ));
 sg13g2_dfrbp_1 _3204_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net68),
    .D(_0062_),
    .Q_N(_1542_),
    .Q(\logo_top[5] ));
 sg13g2_dfrbp_1 _3205_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net66),
    .D(_0063_),
    .Q_N(_0013_),
    .Q(\logo_top[6] ));
 sg13g2_dfrbp_1 _3206_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net64),
    .D(_0064_),
    .Q_N(_1541_),
    .Q(\logo_top[7] ));
 sg13g2_dfrbp_1 _3207_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net62),
    .D(_0065_),
    .Q_N(_0014_),
    .Q(\logo_top[8] ));
 sg13g2_dfrbp_1 _3208_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net60),
    .D(_0066_),
    .Q_N(_1540_),
    .Q(\logo_top[9] ));
 sg13g2_dfrbp_1 _3209_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net58),
    .D(_0067_),
    .Q_N(_1539_),
    .Q(dir_x));
 sg13g2_dfrbp_1 _3210_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net56),
    .D(_0068_),
    .Q_N(_1538_),
    .Q(dir_y));
 sg13g2_dfrbp_1 _3211_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net54),
    .D(net140),
    .Q_N(_0004_),
    .Q(manual_mode));
 sg13g2_dfrbp_1 _3212_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net52),
    .D(net135),
    .Q_N(_0018_),
    .Q(\color_index[0] ));
 sg13g2_dfrbp_1 _3213_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net50),
    .D(net174),
    .Q_N(_0016_),
    .Q(\color_index[1] ));
 sg13g2_dfrbp_1 _3214_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net48),
    .D(net142),
    .Q_N(_0015_),
    .Q(\color_index[2] ));
 sg13g2_dfrbp_1 _3215_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net46),
    .D(_0073_),
    .Q_N(_1537_),
    .Q(\prev_y[0] ));
 sg13g2_dfrbp_1 _3216_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net45),
    .D(_0074_),
    .Q_N(_1536_),
    .Q(\prev_y[1] ));
 sg13g2_dfrbp_1 _3217_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net44),
    .D(_0075_),
    .Q_N(_1535_),
    .Q(\prev_y[2] ));
 sg13g2_dfrbp_1 _3218_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net43),
    .D(_0076_),
    .Q_N(_1534_),
    .Q(\prev_y[3] ));
 sg13g2_dfrbp_1 _3219_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net42),
    .D(_0077_),
    .Q_N(_1533_),
    .Q(\prev_y[4] ));
 sg13g2_dfrbp_1 _3220_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net41),
    .D(_0078_),
    .Q_N(_1532_),
    .Q(\prev_y[5] ));
 sg13g2_dfrbp_1 _3221_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net38),
    .D(_0079_),
    .Q_N(_1531_),
    .Q(\prev_y[6] ));
 sg13g2_dfrbp_1 _3222_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net36),
    .D(_0080_),
    .Q_N(_1530_),
    .Q(\prev_y[7] ));
 sg13g2_dfrbp_1 _3223_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net34),
    .D(_0081_),
    .Q_N(_1529_),
    .Q(\prev_y[8] ));
 sg13g2_dfrbp_1 _3224_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net32),
    .D(_0082_),
    .Q_N(_1528_),
    .Q(\prev_y[9] ));
 sg13g2_dfrbp_1 _3225_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net30),
    .D(_0083_),
    .Q_N(_1527_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _3226_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net28),
    .D(_0084_),
    .Q_N(_1526_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _3227_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net26),
    .D(_0085_),
    .Q_N(_1525_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _3228_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net88),
    .D(_0086_),
    .Q_N(_1574_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _3229_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net107),
    .D(net125),
    .Q_N(_1575_),
    .Q(\gamepad.driver.pmod_clk_prev ));
 sg13g2_dfrbp_1 _3230_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net24),
    .D(net126),
    .Q_N(_1524_),
    .Q(\gamepad.driver.pmod_latch_prev ));
 sg13g2_dfrbp_1 _3231_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net22),
    .D(net154),
    .Q_N(_1523_),
    .Q(\gamepad.driver.shift_reg[0] ));
 sg13g2_dfrbp_1 _3232_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net116),
    .D(net185),
    .Q_N(_1522_),
    .Q(\gamepad.driver.shift_reg[1] ));
 sg13g2_dfrbp_1 _3233_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net112),
    .D(_0089_),
    .Q_N(_1521_),
    .Q(\gamepad.driver.shift_reg[2] ));
 sg13g2_dfrbp_1 _3234_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net97),
    .D(_0090_),
    .Q_N(_1520_),
    .Q(\gamepad.driver.shift_reg[3] ));
 sg13g2_dfrbp_1 _3235_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net93),
    .D(net172),
    .Q_N(_1519_),
    .Q(\gamepad.driver.shift_reg[4] ));
 sg13g2_dfrbp_1 _3236_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net89),
    .D(net183),
    .Q_N(_1518_),
    .Q(\gamepad.driver.shift_reg[5] ));
 sg13g2_dfrbp_1 _3237_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net83),
    .D(net166),
    .Q_N(_1517_),
    .Q(\gamepad.driver.shift_reg[6] ));
 sg13g2_dfrbp_1 _3238_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net79),
    .D(_0094_),
    .Q_N(_1516_),
    .Q(\gamepad.driver.shift_reg[7] ));
 sg13g2_dfrbp_1 _3239_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net75),
    .D(net170),
    .Q_N(_1515_),
    .Q(\gamepad.driver.shift_reg[8] ));
 sg13g2_dfrbp_1 _3240_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net71),
    .D(net180),
    .Q_N(_1514_),
    .Q(\gamepad.driver.shift_reg[9] ));
 sg13g2_dfrbp_1 _3241_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net67),
    .D(net177),
    .Q_N(_1513_),
    .Q(\gamepad.driver.shift_reg[10] ));
 sg13g2_dfrbp_1 _3242_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net63),
    .D(net150),
    .Q_N(_1512_),
    .Q(\gamepad.driver.shift_reg[11] ));
 sg13g2_dfrbp_1 _3243_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net59),
    .D(_0099_),
    .Q_N(_1511_),
    .Q(\gamepad.driver.pmod_data_sync[0] ));
 sg13g2_dfrbp_1 _3244_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net57),
    .D(_0100_),
    .Q_N(_1510_),
    .Q(\gamepad.driver.pmod_data_sync[1] ));
 sg13g2_dfrbp_1 _3245_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net55),
    .D(_0101_),
    .Q_N(_1509_),
    .Q(\gamepad.driver.pmod_clk_sync[0] ));
 sg13g2_dfrbp_1 _3246_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net53),
    .D(_0102_),
    .Q_N(_1508_),
    .Q(\gamepad.driver.pmod_clk_sync[1] ));
 sg13g2_dfrbp_1 _3247_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net51),
    .D(_0103_),
    .Q_N(_1507_),
    .Q(\gamepad.driver.pmod_latch_sync[0] ));
 sg13g2_dfrbp_1 _3248_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net118),
    .D(_0104_),
    .Q_N(_1576_),
    .Q(\gamepad.driver.pmod_latch_sync[1] ));
 sg13g2_dfrbp_1 _3249_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net49),
    .D(net200),
    .Q_N(_1506_),
    .Q(hsync));
 sg13g2_dfrbp_1 _3250_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net47),
    .D(_0105_),
    .Q_N(_0017_),
    .Q(\pix_y[0] ));
 sg13g2_dfrbp_1 _3251_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net114),
    .D(_0106_),
    .Q_N(_1505_),
    .Q(\pix_y[1] ));
 sg13g2_dfrbp_1 _3252_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net95),
    .D(_0107_),
    .Q_N(_1504_),
    .Q(\pix_y[2] ));
 sg13g2_dfrbp_1 _3253_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net85),
    .D(_0108_),
    .Q_N(_1503_),
    .Q(\pix_y[3] ));
 sg13g2_dfrbp_1 _3254_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net77),
    .D(_0109_),
    .Q_N(_1502_),
    .Q(\pix_y[4] ));
 sg13g2_dfrbp_1 _3255_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net69),
    .D(_0110_),
    .Q_N(_1501_),
    .Q(\pix_y[5] ));
 sg13g2_dfrbp_1 _3256_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net61),
    .D(_0111_),
    .Q_N(_1500_),
    .Q(\pix_y[6] ));
 sg13g2_dfrbp_1 _3257_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net99),
    .D(_0112_),
    .Q_N(_1499_),
    .Q(\pix_y[7] ));
 sg13g2_dfrbp_1 _3258_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net81),
    .D(_0113_),
    .Q_N(_1498_),
    .Q(\pix_y[8] ));
 sg13g2_dfrbp_1 _3259_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net119),
    .D(_0114_),
    .Q_N(_1577_),
    .Q(\pix_y[9] ));
 sg13g2_dfrbp_1 _3260_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net120),
    .D(net164),
    .Q_N(_1578_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_dfrbp_1 _3261_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net121),
    .D(_0000_),
    .Q_N(_1579_),
    .Q(\palette_inst.rrggbb[0] ));
 sg13g2_dfrbp_1 _3262_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net122),
    .D(_0001_),
    .Q_N(_1580_),
    .Q(\palette_inst.rrggbb[1] ));
 sg13g2_dfrbp_1 _3263_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net123),
    .D(_0002_),
    .Q_N(_1581_),
    .Q(\palette_inst.rrggbb[2] ));
 sg13g2_dfrbp_1 _3264_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net65),
    .D(_0003_),
    .Q_N(_1497_),
    .Q(\palette_inst.rrggbb[3] ));
 sg13g2_dfrbp_1 _3265_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net91),
    .D(_0115_),
    .Q_N(_1496_),
    .Q(\palette_inst.rrggbb[4] ));
 sg13g2_dfrbp_1 _3266_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net73),
    .D(_0116_),
    .Q_N(_1495_),
    .Q(\palette_inst.rrggbb[5] ));
 sg13g2_tiehi _3174__23 (.L_HI(net23));
 sg13g2_tiehi _3230__24 (.L_HI(net24));
 sg13g2_tiehi _3173__25 (.L_HI(net25));
 sg13g2_tiehi _3227__26 (.L_HI(net26));
 sg13g2_tiehi _3172__27 (.L_HI(net27));
 sg13g2_tiehi _3226__28 (.L_HI(net28));
 sg13g2_tiehi _3171__29 (.L_HI(net29));
 sg13g2_tiehi _3225__30 (.L_HI(net30));
 sg13g2_tiehi _3170__31 (.L_HI(net31));
 sg13g2_tiehi _3224__32 (.L_HI(net32));
 sg13g2_tiehi _3169__33 (.L_HI(net33));
 sg13g2_tiehi _3223__34 (.L_HI(net34));
 sg13g2_tiehi _3168__35 (.L_HI(net35));
 sg13g2_tiehi _3222__36 (.L_HI(net36));
 sg13g2_tiehi _3167__37 (.L_HI(net37));
 sg13g2_tiehi _3221__38 (.L_HI(net38));
 sg13g2_tiehi _3166__39 (.L_HI(net39));
 sg13g2_tiehi _3165__40 (.L_HI(net40));
 sg13g2_tiehi _3220__41 (.L_HI(net41));
 sg13g2_tiehi _3219__42 (.L_HI(net42));
 sg13g2_tiehi _3218__43 (.L_HI(net43));
 sg13g2_tiehi _3217__44 (.L_HI(net44));
 sg13g2_tiehi _3216__45 (.L_HI(net45));
 sg13g2_tiehi _3215__46 (.L_HI(net46));
 sg13g2_tiehi _3250__47 (.L_HI(net47));
 sg13g2_tiehi _3214__48 (.L_HI(net48));
 sg13g2_tiehi _3249__49 (.L_HI(net49));
 sg13g2_tiehi _3213__50 (.L_HI(net50));
 sg13g2_tiehi _3247__51 (.L_HI(net51));
 sg13g2_tiehi _3212__52 (.L_HI(net52));
 sg13g2_tiehi _3246__53 (.L_HI(net53));
 sg13g2_tiehi _3211__54 (.L_HI(net54));
 sg13g2_tiehi _3245__55 (.L_HI(net55));
 sg13g2_tiehi _3210__56 (.L_HI(net56));
 sg13g2_tiehi _3244__57 (.L_HI(net57));
 sg13g2_tiehi _3209__58 (.L_HI(net58));
 sg13g2_tiehi _3243__59 (.L_HI(net59));
 sg13g2_tiehi _3208__60 (.L_HI(net60));
 sg13g2_tiehi _3256__61 (.L_HI(net61));
 sg13g2_tiehi _3207__62 (.L_HI(net62));
 sg13g2_tiehi _3242__63 (.L_HI(net63));
 sg13g2_tiehi _3206__64 (.L_HI(net64));
 sg13g2_tiehi _3264__65 (.L_HI(net65));
 sg13g2_tiehi _3205__66 (.L_HI(net66));
 sg13g2_tiehi _3241__67 (.L_HI(net67));
 sg13g2_tiehi _3204__68 (.L_HI(net68));
 sg13g2_tiehi _3255__69 (.L_HI(net69));
 sg13g2_tiehi _3203__70 (.L_HI(net70));
 sg13g2_tiehi _3240__71 (.L_HI(net71));
 sg13g2_tiehi _3202__72 (.L_HI(net72));
 sg13g2_tiehi _3266__73 (.L_HI(net73));
 sg13g2_tiehi _3201__74 (.L_HI(net74));
 sg13g2_tiehi _3239__75 (.L_HI(net75));
 sg13g2_tiehi _3200__76 (.L_HI(net76));
 sg13g2_tiehi _3254__77 (.L_HI(net77));
 sg13g2_tiehi _3199__78 (.L_HI(net78));
 sg13g2_tiehi _3238__79 (.L_HI(net79));
 sg13g2_tiehi _3198__80 (.L_HI(net80));
 sg13g2_tiehi _3258__81 (.L_HI(net81));
 sg13g2_tiehi _3197__82 (.L_HI(net82));
 sg13g2_tiehi _3237__83 (.L_HI(net83));
 sg13g2_tiehi _3196__84 (.L_HI(net84));
 sg13g2_tiehi _3253__85 (.L_HI(net85));
 sg13g2_tiehi _3195__86 (.L_HI(net86));
 sg13g2_tiehi _3164__87 (.L_HI(net87));
 sg13g2_tiehi _3228__88 (.L_HI(net88));
 sg13g2_tiehi _3236__89 (.L_HI(net89));
 sg13g2_tiehi _3194__90 (.L_HI(net90));
 sg13g2_tiehi _3265__91 (.L_HI(net91));
 sg13g2_tiehi _3193__92 (.L_HI(net92));
 sg13g2_tiehi _3235__93 (.L_HI(net93));
 sg13g2_tiehi _3192__94 (.L_HI(net94));
 sg13g2_tiehi _3252__95 (.L_HI(net95));
 sg13g2_tiehi _3191__96 (.L_HI(net96));
 sg13g2_tiehi _3234__97 (.L_HI(net97));
 sg13g2_tiehi _3190__98 (.L_HI(net98));
 sg13g2_tiehi _3257__99 (.L_HI(net99));
 sg13g2_tiehi _3189__100 (.L_HI(net100));
 sg13g2_tiehi _3188__101 (.L_HI(net101));
 sg13g2_tiehi _3187__102 (.L_HI(net102));
 sg13g2_tiehi _3186__103 (.L_HI(net103));
 sg13g2_tiehi _3185__104 (.L_HI(net104));
 sg13g2_tiehi _3184__105 (.L_HI(net105));
 sg13g2_tiehi _3183__106 (.L_HI(net106));
 sg13g2_tiehi _3229__107 (.L_HI(net107));
 sg13g2_tiehi _3182__108 (.L_HI(net108));
 sg13g2_tiehi _3181__109 (.L_HI(net109));
 sg13g2_tiehi _3180__110 (.L_HI(net110));
 sg13g2_tiehi _3179__111 (.L_HI(net111));
 sg13g2_tiehi _3233__112 (.L_HI(net112));
 sg13g2_tiehi _3178__113 (.L_HI(net113));
 sg13g2_tiehi _3251__114 (.L_HI(net114));
 sg13g2_tiehi _3177__115 (.L_HI(net115));
 sg13g2_tiehi _3232__116 (.L_HI(net116));
 sg13g2_tiehi _3176__117 (.L_HI(net117));
 sg13g2_tiehi _3248__118 (.L_HI(net118));
 sg13g2_tiehi _3259__119 (.L_HI(net119));
 sg13g2_tiehi _3260__120 (.L_HI(net120));
 sg13g2_tiehi _3261__121 (.L_HI(net121));
 sg13g2_tiehi _3262__122 (.L_HI(net122));
 sg13g2_tiehi _3263__123 (.L_HI(net123));
 sg13g2_tiehi _3175__124 (.L_HI(net124));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_7 (.L_LO(net7));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_8 (.L_LO(net8));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_9 (.L_LO(net9));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_10 (.L_LO(net10));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_11 (.L_LO(net11));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_12 (.L_LO(net12));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_13 (.L_LO(net13));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_14 (.L_LO(net14));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_15 (.L_LO(net15));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_16 (.L_LO(net16));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_17 (.L_LO(net17));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_18 (.L_LO(net18));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_19 (.L_LO(net19));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_20 (.L_LO(net20));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_21 (.L_LO(net21));
 sg13g2_tiehi _3231__22 (.L_HI(net22));
 sg13g2_buf_2 _3386_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_2 _3387_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout642 (.A(net644),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_0571_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(net646),
    .X(net645));
 sg13g2_buf_1 fanout646 (.A(net647),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_0560_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_0472_),
    .X(net648));
 sg13g2_buf_1 fanout649 (.A(_0472_),
    .X(net649));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(_0922_));
 sg13g2_buf_2 fanout651 (.A(_0470_),
    .X(net651));
 sg13g2_buf_4 fanout652 (.X(net652),
    .A(_1043_));
 sg13g2_buf_4 fanout653 (.X(net653),
    .A(net654));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(_0926_));
 sg13g2_buf_2 fanout655 (.A(net658),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(net658),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_0925_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(net660),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_1187_),
    .X(net660));
 sg13g2_buf_4 fanout661 (.X(net661),
    .A(net662));
 sg13g2_buf_4 fanout662 (.X(net662),
    .A(_1126_));
 sg13g2_buf_4 fanout663 (.X(net663),
    .A(_1113_));
 sg13g2_buf_2 fanout664 (.A(_1113_),
    .X(net664));
 sg13g2_buf_4 fanout665 (.X(net665),
    .A(_1100_));
 sg13g2_buf_2 fanout666 (.A(_1100_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(net669),
    .X(net668));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(_1088_));
 sg13g2_buf_2 fanout670 (.A(net672),
    .X(net670));
 sg13g2_buf_1 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_4 fanout672 (.X(net672),
    .A(_1060_));
 sg13g2_buf_2 fanout673 (.A(_1059_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_1059_),
    .X(net674));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(_1041_));
 sg13g2_buf_1 fanout676 (.A(_1041_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_1037_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(net679),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(_1027_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_1015_),
    .X(net680));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(_1001_));
 sg13g2_buf_2 fanout682 (.A(_0998_),
    .X(net682));
 sg13g2_buf_1 fanout683 (.A(_0998_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(net686),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(net686),
    .X(net685));
 sg13g2_buf_4 fanout686 (.X(net686),
    .A(_0992_));
 sg13g2_buf_4 fanout687 (.X(net687),
    .A(net688));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(net689));
 sg13g2_buf_4 fanout689 (.X(net689),
    .A(_0971_));
 sg13g2_buf_2 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(net693),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_0970_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_0451_),
    .X(net694));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(_1098_));
 sg13g2_buf_4 fanout696 (.X(net696),
    .A(_1074_));
 sg13g2_buf_1 fanout697 (.A(_1074_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(net702),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(net702),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(net702));
 sg13g2_buf_4 fanout702 (.X(net702),
    .A(_1073_));
 sg13g2_buf_4 fanout703 (.X(net703),
    .A(_1023_));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(_1023_));
 sg13g2_buf_2 fanout705 (.A(_1022_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_1022_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(net709),
    .X(net707));
 sg13g2_buf_1 fanout708 (.A(net709),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_1022_),
    .X(net709));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(net714));
 sg13g2_buf_2 fanout711 (.A(net714),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(net713),
    .X(net712));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(net714));
 sg13g2_buf_2 fanout714 (.A(_1021_),
    .X(net714));
 sg13g2_buf_4 fanout715 (.X(net715),
    .A(_0982_));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(_0980_));
 sg13g2_buf_1 fanout717 (.A(_0980_),
    .X(net717));
 sg13g2_buf_4 fanout718 (.X(net718),
    .A(_0978_));
 sg13g2_buf_4 fanout719 (.X(net719),
    .A(_0969_));
 sg13g2_buf_2 fanout720 (.A(_0969_),
    .X(net720));
 sg13g2_buf_4 fanout721 (.X(net721),
    .A(_0968_));
 sg13g2_buf_2 fanout722 (.A(_0968_),
    .X(net722));
 sg13g2_buf_4 fanout723 (.X(net723),
    .A(net724));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(_0967_));
 sg13g2_buf_4 fanout725 (.X(net725),
    .A(net726));
 sg13g2_buf_2 fanout726 (.A(net727),
    .X(net726));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(_0965_));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(net729));
 sg13g2_buf_4 fanout729 (.X(net729),
    .A(net732));
 sg13g2_buf_2 fanout730 (.A(net731),
    .X(net730));
 sg13g2_buf_4 fanout731 (.X(net731),
    .A(net732));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(_0956_));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(net736));
 sg13g2_buf_2 fanout734 (.A(net736),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(net736),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(net738),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(net738),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_0955_),
    .X(net738));
 sg13g2_buf_4 fanout739 (.X(net739),
    .A(net741));
 sg13g2_buf_1 fanout740 (.A(net741),
    .X(net740));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(net747));
 sg13g2_buf_2 fanout742 (.A(net746),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(net746),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(net746),
    .X(net744));
 sg13g2_buf_1 fanout745 (.A(net746),
    .X(net745));
 sg13g2_buf_4 fanout746 (.X(net746),
    .A(net747));
 sg13g2_buf_2 fanout747 (.A(_0929_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(net749),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(net756),
    .X(net749));
 sg13g2_buf_4 fanout750 (.X(net750),
    .A(net756));
 sg13g2_buf_1 fanout751 (.A(net756),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(net753),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(net756),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(net755),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(net756),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_0928_),
    .X(net756));
 sg13g2_buf_4 fanout757 (.X(net757),
    .A(net758));
 sg13g2_buf_2 fanout758 (.A(net759),
    .X(net758));
 sg13g2_buf_4 fanout759 (.X(net759),
    .A(net760));
 sg13g2_buf_4 fanout760 (.X(net760),
    .A(_0988_));
 sg13g2_buf_4 fanout761 (.X(net761),
    .A(net763));
 sg13g2_buf_4 fanout762 (.X(net762),
    .A(net763));
 sg13g2_buf_4 fanout763 (.X(net763),
    .A(_0988_));
 sg13g2_buf_2 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_4 fanout765 (.X(net765),
    .A(net766));
 sg13g2_buf_4 fanout766 (.X(net766),
    .A(_0987_));
 sg13g2_buf_2 fanout767 (.A(net769),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(net769),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_0987_),
    .X(net769));
 sg13g2_buf_4 fanout770 (.X(net770),
    .A(_0976_));
 sg13g2_buf_2 fanout771 (.A(_0976_),
    .X(net771));
 sg13g2_buf_4 fanout772 (.X(net772),
    .A(_0949_));
 sg13g2_buf_2 fanout773 (.A(_0949_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_4 fanout775 (.X(net775),
    .A(net776));
 sg13g2_buf_4 fanout776 (.X(net776),
    .A(_0948_));
 sg13g2_buf_4 fanout777 (.X(net777),
    .A(_0997_));
 sg13g2_buf_4 fanout778 (.X(net778),
    .A(_0996_));
 sg13g2_buf_2 fanout779 (.A(_0996_),
    .X(net779));
 sg13g2_buf_4 fanout780 (.X(net780),
    .A(_0989_));
 sg13g2_buf_4 fanout781 (.X(net781),
    .A(_0694_));
 sg13g2_buf_2 fanout782 (.A(_0694_),
    .X(net782));
 sg13g2_buf_4 fanout783 (.X(net783),
    .A(_0439_));
 sg13g2_buf_1 fanout784 (.A(_0439_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(net789),
    .X(net785));
 sg13g2_buf_4 fanout786 (.X(net786),
    .A(net789));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(net788));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(net789));
 sg13g2_buf_2 fanout789 (.A(_0931_),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(net791));
 sg13g2_buf_2 fanout791 (.A(net793),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(net793),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_0930_),
    .X(net793));
 sg13g2_buf_4 fanout794 (.X(net794),
    .A(net795));
 sg13g2_buf_4 fanout795 (.X(net795),
    .A(_0930_));
 sg13g2_buf_4 fanout796 (.X(net796),
    .A(_0693_));
 sg13g2_buf_1 fanout797 (.A(_0693_),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(_0438_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_0438_),
    .X(net799));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(net801));
 sg13g2_buf_2 fanout801 (.A(net802),
    .X(net801));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(net806));
 sg13g2_buf_4 fanout803 (.X(net803),
    .A(net805));
 sg13g2_buf_1 fanout804 (.A(net805),
    .X(net804));
 sg13g2_buf_4 fanout805 (.X(net805),
    .A(net806));
 sg13g2_buf_2 fanout806 (.A(_0933_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(net808),
    .X(net807));
 sg13g2_buf_4 fanout808 (.X(net808),
    .A(net812));
 sg13g2_buf_2 fanout809 (.A(net812),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(net811),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(net812),
    .X(net811));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(_0932_));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(_0733_));
 sg13g2_buf_2 fanout814 (.A(_0733_),
    .X(net814));
 sg13g2_buf_4 fanout815 (.X(net815),
    .A(net178));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(net203));
 sg13g2_buf_2 fanout817 (.A(net818),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(\pix_y[5] ),
    .X(net818));
 sg13g2_buf_4 fanout819 (.X(net819),
    .A(net211));
 sg13g2_buf_2 fanout820 (.A(net821),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(\pix_y[3] ),
    .X(net821));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(net222));
 sg13g2_buf_4 fanout823 (.X(net823),
    .A(net162));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(net219));
 sg13g2_buf_2 fanout825 (.A(net829),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(net829),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(net829),
    .X(net827));
 sg13g2_buf_1 fanout828 (.A(net829),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(manual_mode),
    .X(net829));
 sg13g2_buf_4 fanout830 (.X(net830),
    .A(net831));
 sg13g2_buf_4 fanout831 (.X(net831),
    .A(net234));
 sg13g2_buf_4 fanout832 (.X(net832),
    .A(net833));
 sg13g2_buf_4 fanout833 (.X(net833),
    .A(dir_x));
 sg13g2_buf_4 fanout834 (.X(net834),
    .A(net226));
 sg13g2_buf_2 fanout835 (.A(\logo_top[5] ),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(net229),
    .X(net836));
 sg13g2_buf_4 fanout837 (.X(net837),
    .A(net218));
 sg13g2_buf_4 fanout838 (.X(net838),
    .A(\logo_top[0] ));
 sg13g2_buf_2 fanout839 (.A(\logo_left[7] ),
    .X(net839));
 sg13g2_buf_4 fanout840 (.X(net840),
    .A(net225));
 sg13g2_buf_4 fanout841 (.X(net841),
    .A(\logo_left[3] ));
 sg13g2_buf_4 fanout842 (.X(net842),
    .A(net215));
 sg13g2_buf_4 fanout843 (.X(net843),
    .A(\logo_left[0] ));
 sg13g2_buf_4 fanout844 (.X(net844),
    .A(net845));
 sg13g2_buf_4 fanout845 (.X(net845),
    .A(_0750_));
 sg13g2_buf_4 fanout846 (.X(net846),
    .A(net848));
 sg13g2_buf_4 fanout847 (.X(net847),
    .A(net848));
 sg13g2_buf_2 fanout848 (.A(rst_n),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(net852),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(net852),
    .X(net850));
 sg13g2_buf_1 fanout851 (.A(net852),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(rst_n),
    .X(net852));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_tielo tt_um_tinytapeout_logo_screensaver_6 (.L_LO(net6));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\gamepad.driver.pmod_clk_sync[1] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold2 (.A(\gamepad.driver.pmod_latch_sync[1] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0021_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0017_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold5 (.A(\gamepad.driver.pmod_data_sync[0] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold6 (.A(\gamepad.driver.pmod_latch_sync[0] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold7 (.A(\gamepad.driver.pmod_clk_sync[0] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0019_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0057_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0018_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0070_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0020_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0047_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0004_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0675_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0069_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold17 (.A(\color_index[2] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0072_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold19 (.A(gamepad_start_prev),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0036_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold21 (.A(\gamepad.decoder.data_reg[9] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0033_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold23 (.A(\gamepad.decoder.data_reg[2] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0026_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold25 (.A(\gamepad.driver.shift_reg[11] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0098_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold27 (.A(\gamepad.decoder.data_reg[10] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0034_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold29 (.A(\gamepad.driver.pmod_data_sync[1] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0087_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold31 (.A(\gamepad.decoder.data_reg[11] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold32 (.A(\gamepad.decoder.data_reg[0] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0024_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold34 (.A(\gamepad.decoder.data_reg[3] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0027_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold36 (.A(\gamepad.decoder.data_reg[1] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0025_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold38 (.A(\pix_y[1] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0776_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0006_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold41 (.A(\gamepad.driver.shift_reg[6] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0093_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold43 (.A(\gamepad.decoder.data_reg[5] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0029_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold45 (.A(\gamepad.driver.shift_reg[8] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0095_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold47 (.A(\gamepad.driver.shift_reg[4] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold48 (.A(_0091_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold49 (.A(\color_index[1] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0071_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold51 (.A(\gamepad.driver.shift_reg[7] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold52 (.A(\gamepad.driver.shift_reg[10] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0097_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold54 (.A(\pix_y[9] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold55 (.A(\gamepad.driver.shift_reg[9] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0096_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold57 (.A(\gamepad.decoder.data_reg[7] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold58 (.A(\gamepad.driver.shift_reg[5] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0092_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold60 (.A(\gamepad.driver.shift_reg[1] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0088_),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold62 (.A(\gamepad.decoder.data_reg[8] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold63 (.A(\gamepad.decoder.data_reg[6] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold64 (.A(\palette_inst.rrggbb[5] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold65 (.A(\gamepad.decoder.data_reg[4] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold66 (.A(\pix_x[2] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0453_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0039_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold69 (.A(\gamepad.driver.shift_reg[2] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold70 (.A(\gamepad.driver.shift_reg[3] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold71 (.A(\palette_inst.rrggbb[2] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold72 (.A(\palette_inst.rrggbb[3] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold73 (.A(\pix_x[6] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0458_),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold75 (.A(\pix_x[8] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0005_),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold77 (.A(\palette_inst.rrggbb[0] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold78 (.A(\pix_x[7] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold79 (.A(\pix_y[7] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold80 (.A(\palette_inst.rrggbb[1] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold81 (.A(\pix_x[1] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0452_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold83 (.A(\palette_inst.rrggbb[4] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold84 (.A(\pix_x[4] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold85 (.A(\pix_x[3] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold86 (.A(\pix_x[5] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold87 (.A(\pix_y[4] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold88 (.A(\pix_x[9] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold89 (.A(\pix_y[6] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold90 (.A(\pix_y[8] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold91 (.A(\logo_left[1] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0015_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0892_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold94 (.A(\logo_top[1] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold95 (.A(\pix_y[0] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0016_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold97 (.A(\pix_y[8] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold98 (.A(\pix_y[2] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold99 (.A(\logo_top[4] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold100 (.A(\logo_top[8] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold101 (.A(\logo_left[6] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold102 (.A(\logo_top[9] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold103 (.A(\logo_left[8] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold104 (.A(\logo_left[2] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold105 (.A(\logo_top[2] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold106 (.A(\logo_top[3] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold107 (.A(\logo_left[9] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold108 (.A(\logo_left[4] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold109 (.A(\logo_left[5] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold110 (.A(dir_y),
    .X(net234));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_fill_2 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_150 ();
 sg13g2_decap_8 FILLER_15_157 ();
 sg13g2_decap_8 FILLER_15_164 ();
 sg13g2_decap_8 FILLER_15_171 ();
 sg13g2_decap_8 FILLER_15_178 ();
 sg13g2_decap_8 FILLER_15_185 ();
 sg13g2_decap_8 FILLER_15_192 ();
 sg13g2_decap_8 FILLER_15_199 ();
 sg13g2_decap_8 FILLER_15_206 ();
 sg13g2_decap_8 FILLER_15_213 ();
 sg13g2_decap_8 FILLER_15_220 ();
 sg13g2_decap_8 FILLER_15_227 ();
 sg13g2_decap_8 FILLER_15_234 ();
 sg13g2_decap_8 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_decap_8 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_262 ();
 sg13g2_decap_8 FILLER_15_269 ();
 sg13g2_decap_8 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_283 ();
 sg13g2_decap_8 FILLER_15_290 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_346 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_15_388 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_fill_2 FILLER_16_119 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_decap_8 FILLER_16_162 ();
 sg13g2_decap_8 FILLER_16_169 ();
 sg13g2_decap_8 FILLER_16_176 ();
 sg13g2_decap_8 FILLER_16_183 ();
 sg13g2_decap_8 FILLER_16_190 ();
 sg13g2_decap_8 FILLER_16_197 ();
 sg13g2_decap_8 FILLER_16_204 ();
 sg13g2_decap_8 FILLER_16_211 ();
 sg13g2_decap_8 FILLER_16_218 ();
 sg13g2_decap_8 FILLER_16_225 ();
 sg13g2_decap_8 FILLER_16_232 ();
 sg13g2_decap_8 FILLER_16_239 ();
 sg13g2_decap_8 FILLER_16_246 ();
 sg13g2_decap_8 FILLER_16_253 ();
 sg13g2_decap_8 FILLER_16_260 ();
 sg13g2_decap_8 FILLER_16_267 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_decap_8 FILLER_16_295 ();
 sg13g2_decap_8 FILLER_16_302 ();
 sg13g2_decap_8 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_decap_8 FILLER_16_323 ();
 sg13g2_decap_8 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_fill_2 FILLER_17_98 ();
 sg13g2_fill_1 FILLER_17_105 ();
 sg13g2_fill_2 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_125 ();
 sg13g2_fill_2 FILLER_17_134 ();
 sg13g2_fill_1 FILLER_17_136 ();
 sg13g2_decap_8 FILLER_17_166 ();
 sg13g2_decap_8 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_180 ();
 sg13g2_decap_8 FILLER_17_187 ();
 sg13g2_decap_8 FILLER_17_194 ();
 sg13g2_decap_8 FILLER_17_201 ();
 sg13g2_decap_8 FILLER_17_208 ();
 sg13g2_decap_8 FILLER_17_215 ();
 sg13g2_decap_8 FILLER_17_222 ();
 sg13g2_decap_8 FILLER_17_229 ();
 sg13g2_decap_8 FILLER_17_236 ();
 sg13g2_decap_8 FILLER_17_243 ();
 sg13g2_decap_8 FILLER_17_250 ();
 sg13g2_decap_8 FILLER_17_257 ();
 sg13g2_decap_8 FILLER_17_264 ();
 sg13g2_decap_8 FILLER_17_271 ();
 sg13g2_decap_8 FILLER_17_278 ();
 sg13g2_decap_8 FILLER_17_285 ();
 sg13g2_decap_8 FILLER_17_292 ();
 sg13g2_decap_8 FILLER_17_299 ();
 sg13g2_decap_8 FILLER_17_306 ();
 sg13g2_decap_8 FILLER_17_313 ();
 sg13g2_decap_8 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_17_327 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_fill_1 FILLER_18_84 ();
 sg13g2_fill_2 FILLER_18_90 ();
 sg13g2_decap_4 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_134 ();
 sg13g2_fill_1 FILLER_18_140 ();
 sg13g2_fill_1 FILLER_18_158 ();
 sg13g2_decap_8 FILLER_18_174 ();
 sg13g2_decap_8 FILLER_18_181 ();
 sg13g2_decap_8 FILLER_18_188 ();
 sg13g2_decap_8 FILLER_18_195 ();
 sg13g2_decap_8 FILLER_18_202 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_decap_8 FILLER_18_223 ();
 sg13g2_decap_8 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_237 ();
 sg13g2_decap_8 FILLER_18_244 ();
 sg13g2_decap_8 FILLER_18_251 ();
 sg13g2_decap_8 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_272 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_decap_8 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_293 ();
 sg13g2_decap_8 FILLER_18_300 ();
 sg13g2_decap_8 FILLER_18_307 ();
 sg13g2_decap_8 FILLER_18_314 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_decap_8 FILLER_18_356 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_4 FILLER_19_70 ();
 sg13g2_decap_4 FILLER_19_114 ();
 sg13g2_fill_2 FILLER_19_118 ();
 sg13g2_decap_4 FILLER_19_125 ();
 sg13g2_fill_2 FILLER_19_129 ();
 sg13g2_fill_1 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_146 ();
 sg13g2_decap_8 FILLER_19_153 ();
 sg13g2_decap_4 FILLER_19_160 ();
 sg13g2_decap_4 FILLER_19_177 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_decap_8 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_249 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_84 ();
 sg13g2_fill_1 FILLER_20_96 ();
 sg13g2_fill_1 FILLER_20_108 ();
 sg13g2_decap_8 FILLER_20_124 ();
 sg13g2_fill_1 FILLER_20_131 ();
 sg13g2_fill_2 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_142 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_fill_1 FILLER_20_154 ();
 sg13g2_fill_2 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_192 ();
 sg13g2_decap_8 FILLER_20_199 ();
 sg13g2_decap_8 FILLER_20_206 ();
 sg13g2_decap_8 FILLER_20_213 ();
 sg13g2_decap_8 FILLER_20_220 ();
 sg13g2_decap_8 FILLER_20_227 ();
 sg13g2_decap_8 FILLER_20_234 ();
 sg13g2_decap_8 FILLER_20_241 ();
 sg13g2_decap_8 FILLER_20_248 ();
 sg13g2_decap_8 FILLER_20_255 ();
 sg13g2_decap_8 FILLER_20_262 ();
 sg13g2_decap_8 FILLER_20_269 ();
 sg13g2_decap_8 FILLER_20_276 ();
 sg13g2_decap_8 FILLER_20_283 ();
 sg13g2_decap_8 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_297 ();
 sg13g2_decap_8 FILLER_20_304 ();
 sg13g2_decap_8 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_fill_2 FILLER_21_70 ();
 sg13g2_fill_1 FILLER_21_72 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_4 FILLER_21_105 ();
 sg13g2_fill_2 FILLER_21_113 ();
 sg13g2_fill_1 FILLER_21_115 ();
 sg13g2_decap_4 FILLER_21_126 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_146 ();
 sg13g2_fill_1 FILLER_21_148 ();
 sg13g2_fill_2 FILLER_21_166 ();
 sg13g2_fill_1 FILLER_21_168 ();
 sg13g2_fill_2 FILLER_21_180 ();
 sg13g2_fill_1 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_211 ();
 sg13g2_decap_8 FILLER_21_218 ();
 sg13g2_decap_8 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_232 ();
 sg13g2_decap_8 FILLER_21_239 ();
 sg13g2_decap_8 FILLER_21_246 ();
 sg13g2_decap_8 FILLER_21_253 ();
 sg13g2_decap_8 FILLER_21_260 ();
 sg13g2_decap_8 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_274 ();
 sg13g2_decap_8 FILLER_21_281 ();
 sg13g2_decap_8 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_295 ();
 sg13g2_decap_8 FILLER_21_302 ();
 sg13g2_decap_8 FILLER_21_309 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_fill_2 FILLER_22_72 ();
 sg13g2_decap_4 FILLER_22_79 ();
 sg13g2_fill_2 FILLER_22_83 ();
 sg13g2_fill_1 FILLER_22_94 ();
 sg13g2_decap_8 FILLER_22_99 ();
 sg13g2_decap_8 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_113 ();
 sg13g2_fill_2 FILLER_22_120 ();
 sg13g2_fill_1 FILLER_22_122 ();
 sg13g2_fill_2 FILLER_22_133 ();
 sg13g2_fill_2 FILLER_22_139 ();
 sg13g2_fill_2 FILLER_22_172 ();
 sg13g2_fill_1 FILLER_22_174 ();
 sg13g2_decap_8 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_201 ();
 sg13g2_decap_8 FILLER_22_208 ();
 sg13g2_decap_8 FILLER_22_215 ();
 sg13g2_decap_8 FILLER_22_222 ();
 sg13g2_fill_2 FILLER_22_229 ();
 sg13g2_decap_8 FILLER_22_257 ();
 sg13g2_decap_8 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_271 ();
 sg13g2_decap_8 FILLER_22_278 ();
 sg13g2_decap_8 FILLER_22_285 ();
 sg13g2_decap_8 FILLER_22_292 ();
 sg13g2_decap_8 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_4 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_54 ();
 sg13g2_fill_2 FILLER_23_68 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_89 ();
 sg13g2_fill_1 FILLER_23_91 ();
 sg13g2_decap_4 FILLER_23_109 ();
 sg13g2_decap_4 FILLER_23_123 ();
 sg13g2_fill_1 FILLER_23_127 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_decap_4 FILLER_23_167 ();
 sg13g2_fill_1 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_decap_8 FILLER_23_205 ();
 sg13g2_decap_8 FILLER_23_212 ();
 sg13g2_decap_4 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_223 ();
 sg13g2_decap_8 FILLER_23_251 ();
 sg13g2_decap_8 FILLER_23_258 ();
 sg13g2_decap_8 FILLER_23_265 ();
 sg13g2_decap_8 FILLER_23_272 ();
 sg13g2_decap_8 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_286 ();
 sg13g2_decap_8 FILLER_23_293 ();
 sg13g2_decap_8 FILLER_23_300 ();
 sg13g2_decap_8 FILLER_23_307 ();
 sg13g2_decap_8 FILLER_23_314 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_35 ();
 sg13g2_fill_1 FILLER_24_37 ();
 sg13g2_fill_1 FILLER_24_60 ();
 sg13g2_fill_1 FILLER_24_77 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_fill_1 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_145 ();
 sg13g2_decap_8 FILLER_24_152 ();
 sg13g2_decap_8 FILLER_24_159 ();
 sg13g2_decap_8 FILLER_24_166 ();
 sg13g2_decap_4 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_177 ();
 sg13g2_decap_8 FILLER_24_183 ();
 sg13g2_decap_8 FILLER_24_190 ();
 sg13g2_decap_8 FILLER_24_197 ();
 sg13g2_decap_8 FILLER_24_204 ();
 sg13g2_decap_8 FILLER_24_211 ();
 sg13g2_decap_4 FILLER_24_218 ();
 sg13g2_fill_2 FILLER_24_222 ();
 sg13g2_fill_2 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_246 ();
 sg13g2_decap_4 FILLER_24_257 ();
 sg13g2_fill_2 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_267 ();
 sg13g2_decap_8 FILLER_24_274 ();
 sg13g2_decap_8 FILLER_24_281 ();
 sg13g2_decap_8 FILLER_24_288 ();
 sg13g2_decap_8 FILLER_24_295 ();
 sg13g2_decap_8 FILLER_24_302 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_decap_8 FILLER_24_316 ();
 sg13g2_decap_8 FILLER_24_323 ();
 sg13g2_decap_8 FILLER_24_330 ();
 sg13g2_decap_8 FILLER_24_337 ();
 sg13g2_decap_8 FILLER_24_344 ();
 sg13g2_decap_8 FILLER_24_351 ();
 sg13g2_decap_8 FILLER_24_358 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_decap_8 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_379 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_fill_1 FILLER_25_53 ();
 sg13g2_fill_1 FILLER_25_64 ();
 sg13g2_fill_2 FILLER_25_75 ();
 sg13g2_fill_1 FILLER_25_101 ();
 sg13g2_fill_2 FILLER_25_106 ();
 sg13g2_fill_1 FILLER_25_108 ();
 sg13g2_fill_2 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_fill_1 FILLER_25_135 ();
 sg13g2_fill_1 FILLER_25_141 ();
 sg13g2_fill_2 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_149 ();
 sg13g2_decap_8 FILLER_25_186 ();
 sg13g2_decap_4 FILLER_25_193 ();
 sg13g2_decap_4 FILLER_25_210 ();
 sg13g2_fill_1 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_278 ();
 sg13g2_decap_8 FILLER_25_285 ();
 sg13g2_decap_8 FILLER_25_296 ();
 sg13g2_decap_8 FILLER_25_303 ();
 sg13g2_decap_8 FILLER_25_310 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_42 ();
 sg13g2_fill_2 FILLER_26_46 ();
 sg13g2_fill_2 FILLER_26_59 ();
 sg13g2_fill_1 FILLER_26_61 ();
 sg13g2_decap_4 FILLER_26_67 ();
 sg13g2_fill_1 FILLER_26_71 ();
 sg13g2_decap_8 FILLER_26_82 ();
 sg13g2_decap_4 FILLER_26_89 ();
 sg13g2_decap_8 FILLER_26_97 ();
 sg13g2_fill_2 FILLER_26_104 ();
 sg13g2_fill_2 FILLER_26_121 ();
 sg13g2_decap_4 FILLER_26_129 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_163 ();
 sg13g2_fill_1 FILLER_26_179 ();
 sg13g2_fill_2 FILLER_26_185 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_decap_8 FILLER_26_321 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_4 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_61 ();
 sg13g2_decap_8 FILLER_27_68 ();
 sg13g2_decap_8 FILLER_27_75 ();
 sg13g2_decap_8 FILLER_27_87 ();
 sg13g2_fill_2 FILLER_27_107 ();
 sg13g2_fill_1 FILLER_27_124 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_decap_8 FILLER_27_144 ();
 sg13g2_decap_8 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_158 ();
 sg13g2_fill_2 FILLER_27_179 ();
 sg13g2_fill_1 FILLER_27_181 ();
 sg13g2_fill_1 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_201 ();
 sg13g2_decap_8 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_215 ();
 sg13g2_fill_1 FILLER_27_217 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_decap_8 FILLER_27_253 ();
 sg13g2_decap_8 FILLER_27_260 ();
 sg13g2_decap_4 FILLER_27_267 ();
 sg13g2_fill_2 FILLER_27_271 ();
 sg13g2_decap_8 FILLER_27_299 ();
 sg13g2_decap_8 FILLER_27_306 ();
 sg13g2_decap_8 FILLER_27_313 ();
 sg13g2_decap_8 FILLER_27_320 ();
 sg13g2_decap_8 FILLER_27_327 ();
 sg13g2_decap_8 FILLER_27_334 ();
 sg13g2_decap_8 FILLER_27_341 ();
 sg13g2_decap_8 FILLER_27_348 ();
 sg13g2_decap_8 FILLER_27_355 ();
 sg13g2_decap_8 FILLER_27_362 ();
 sg13g2_decap_8 FILLER_27_369 ();
 sg13g2_decap_8 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_decap_8 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_59 ();
 sg13g2_fill_1 FILLER_28_85 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_4 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_142 ();
 sg13g2_decap_4 FILLER_28_153 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_fill_2 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_186 ();
 sg13g2_decap_8 FILLER_28_193 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_4 FILLER_28_214 ();
 sg13g2_decap_4 FILLER_28_234 ();
 sg13g2_fill_2 FILLER_28_243 ();
 sg13g2_decap_8 FILLER_28_295 ();
 sg13g2_decap_8 FILLER_28_302 ();
 sg13g2_decap_8 FILLER_28_309 ();
 sg13g2_decap_8 FILLER_28_316 ();
 sg13g2_decap_8 FILLER_28_323 ();
 sg13g2_decap_8 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_337 ();
 sg13g2_decap_8 FILLER_28_344 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_decap_8 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_365 ();
 sg13g2_decap_8 FILLER_28_372 ();
 sg13g2_decap_8 FILLER_28_379 ();
 sg13g2_decap_8 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_393 ();
 sg13g2_decap_8 FILLER_28_400 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_59 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_fill_1 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_88 ();
 sg13g2_fill_1 FILLER_29_90 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_109 ();
 sg13g2_decap_4 FILLER_29_118 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_fill_2 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_fill_2 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_194 ();
 sg13g2_decap_8 FILLER_29_201 ();
 sg13g2_decap_8 FILLER_29_208 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_decap_8 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_229 ();
 sg13g2_fill_1 FILLER_29_282 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_307 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_334 ();
 sg13g2_decap_8 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_348 ();
 sg13g2_decap_8 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_29_362 ();
 sg13g2_decap_8 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_51 ();
 sg13g2_fill_1 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_89 ();
 sg13g2_fill_2 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_111 ();
 sg13g2_fill_2 FILLER_30_118 ();
 sg13g2_fill_1 FILLER_30_120 ();
 sg13g2_decap_8 FILLER_30_127 ();
 sg13g2_decap_4 FILLER_30_134 ();
 sg13g2_decap_8 FILLER_30_143 ();
 sg13g2_decap_8 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_215 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_4 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_fill_2 FILLER_30_276 ();
 sg13g2_decap_4 FILLER_30_283 ();
 sg13g2_fill_2 FILLER_30_287 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_decap_8 FILLER_30_349 ();
 sg13g2_decap_8 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_30_363 ();
 sg13g2_decap_8 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_decap_8 FILLER_30_391 ();
 sg13g2_decap_8 FILLER_30_398 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_4 FILLER_31_70 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_fill_1 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_89 ();
 sg13g2_decap_8 FILLER_31_95 ();
 sg13g2_decap_4 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_106 ();
 sg13g2_decap_4 FILLER_31_115 ();
 sg13g2_fill_2 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_127 ();
 sg13g2_fill_1 FILLER_31_134 ();
 sg13g2_decap_4 FILLER_31_139 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_decap_8 FILLER_31_149 ();
 sg13g2_decap_4 FILLER_31_156 ();
 sg13g2_decap_4 FILLER_31_165 ();
 sg13g2_fill_1 FILLER_31_169 ();
 sg13g2_fill_1 FILLER_31_178 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_4 FILLER_31_231 ();
 sg13g2_fill_1 FILLER_31_235 ();
 sg13g2_decap_8 FILLER_31_241 ();
 sg13g2_fill_1 FILLER_31_248 ();
 sg13g2_decap_8 FILLER_31_255 ();
 sg13g2_decap_8 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_269 ();
 sg13g2_decap_8 FILLER_31_279 ();
 sg13g2_fill_2 FILLER_31_286 ();
 sg13g2_fill_1 FILLER_31_288 ();
 sg13g2_fill_2 FILLER_31_293 ();
 sg13g2_fill_1 FILLER_31_295 ();
 sg13g2_fill_2 FILLER_31_300 ();
 sg13g2_fill_1 FILLER_31_302 ();
 sg13g2_decap_8 FILLER_31_325 ();
 sg13g2_decap_8 FILLER_31_332 ();
 sg13g2_decap_8 FILLER_31_339 ();
 sg13g2_decap_8 FILLER_31_346 ();
 sg13g2_decap_8 FILLER_31_353 ();
 sg13g2_decap_8 FILLER_31_360 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_4 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_46 ();
 sg13g2_fill_2 FILLER_32_59 ();
 sg13g2_fill_1 FILLER_32_61 ();
 sg13g2_decap_4 FILLER_32_76 ();
 sg13g2_fill_1 FILLER_32_80 ();
 sg13g2_decap_4 FILLER_32_92 ();
 sg13g2_fill_2 FILLER_32_111 ();
 sg13g2_decap_8 FILLER_32_138 ();
 sg13g2_decap_8 FILLER_32_145 ();
 sg13g2_decap_4 FILLER_32_152 ();
 sg13g2_decap_4 FILLER_32_170 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_decap_8 FILLER_32_204 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_fill_1 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_251 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_fill_2 FILLER_32_283 ();
 sg13g2_fill_1 FILLER_32_285 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_decap_8 FILLER_32_312 ();
 sg13g2_decap_8 FILLER_32_319 ();
 sg13g2_decap_8 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_347 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_4 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_4 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_32 ();
 sg13g2_decap_4 FILLER_33_58 ();
 sg13g2_fill_1 FILLER_33_95 ();
 sg13g2_fill_2 FILLER_33_120 ();
 sg13g2_fill_1 FILLER_33_122 ();
 sg13g2_decap_4 FILLER_33_127 ();
 sg13g2_decap_4 FILLER_33_140 ();
 sg13g2_fill_1 FILLER_33_144 ();
 sg13g2_fill_2 FILLER_33_171 ();
 sg13g2_fill_1 FILLER_33_173 ();
 sg13g2_decap_8 FILLER_33_179 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_4 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_233 ();
 sg13g2_fill_1 FILLER_33_239 ();
 sg13g2_fill_1 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_255 ();
 sg13g2_fill_1 FILLER_33_277 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_fill_2 FILLER_34_59 ();
 sg13g2_fill_1 FILLER_34_61 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_fill_2 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_fill_1 FILLER_34_100 ();
 sg13g2_fill_1 FILLER_34_110 ();
 sg13g2_fill_1 FILLER_34_123 ();
 sg13g2_fill_2 FILLER_34_148 ();
 sg13g2_fill_2 FILLER_34_158 ();
 sg13g2_fill_2 FILLER_34_177 ();
 sg13g2_decap_8 FILLER_34_184 ();
 sg13g2_decap_8 FILLER_34_191 ();
 sg13g2_decap_8 FILLER_34_198 ();
 sg13g2_fill_2 FILLER_34_211 ();
 sg13g2_fill_1 FILLER_34_218 ();
 sg13g2_fill_2 FILLER_34_228 ();
 sg13g2_fill_2 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_241 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_1 FILLER_34_293 ();
 sg13g2_decap_4 FILLER_34_303 ();
 sg13g2_decap_8 FILLER_34_311 ();
 sg13g2_decap_8 FILLER_34_318 ();
 sg13g2_decap_8 FILLER_34_325 ();
 sg13g2_decap_8 FILLER_34_332 ();
 sg13g2_decap_8 FILLER_34_339 ();
 sg13g2_decap_8 FILLER_34_346 ();
 sg13g2_decap_8 FILLER_34_353 ();
 sg13g2_decap_8 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_4 FILLER_35_28 ();
 sg13g2_fill_1 FILLER_35_32 ();
 sg13g2_decap_8 FILLER_35_52 ();
 sg13g2_decap_4 FILLER_35_59 ();
 sg13g2_decap_8 FILLER_35_74 ();
 sg13g2_fill_2 FILLER_35_81 ();
 sg13g2_fill_1 FILLER_35_93 ();
 sg13g2_fill_1 FILLER_35_109 ();
 sg13g2_decap_8 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_181 ();
 sg13g2_decap_4 FILLER_35_193 ();
 sg13g2_fill_1 FILLER_35_197 ();
 sg13g2_decap_4 FILLER_35_202 ();
 sg13g2_fill_1 FILLER_35_217 ();
 sg13g2_fill_1 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_fill_2 FILLER_35_273 ();
 sg13g2_fill_1 FILLER_35_275 ();
 sg13g2_fill_2 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_decap_8 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_338 ();
 sg13g2_decap_8 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_352 ();
 sg13g2_decap_8 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_44 ();
 sg13g2_decap_8 FILLER_36_50 ();
 sg13g2_fill_2 FILLER_36_57 ();
 sg13g2_fill_2 FILLER_36_72 ();
 sg13g2_decap_8 FILLER_36_89 ();
 sg13g2_decap_8 FILLER_36_96 ();
 sg13g2_decap_8 FILLER_36_103 ();
 sg13g2_decap_8 FILLER_36_110 ();
 sg13g2_fill_1 FILLER_36_117 ();
 sg13g2_decap_4 FILLER_36_124 ();
 sg13g2_decap_8 FILLER_36_142 ();
 sg13g2_fill_2 FILLER_36_149 ();
 sg13g2_fill_2 FILLER_36_166 ();
 sg13g2_fill_1 FILLER_36_168 ();
 sg13g2_fill_2 FILLER_36_179 ();
 sg13g2_fill_1 FILLER_36_181 ();
 sg13g2_fill_2 FILLER_36_195 ();
 sg13g2_fill_1 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_decap_4 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_230 ();
 sg13g2_fill_1 FILLER_36_240 ();
 sg13g2_decap_8 FILLER_36_250 ();
 sg13g2_decap_4 FILLER_36_257 ();
 sg13g2_fill_1 FILLER_36_261 ();
 sg13g2_decap_8 FILLER_36_267 ();
 sg13g2_decap_8 FILLER_36_274 ();
 sg13g2_decap_8 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_288 ();
 sg13g2_decap_4 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_320 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_36_346 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_decap_8 FILLER_36_360 ();
 sg13g2_decap_8 FILLER_36_367 ();
 sg13g2_decap_8 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_fill_2 FILLER_37_35 ();
 sg13g2_decap_4 FILLER_37_58 ();
 sg13g2_fill_1 FILLER_37_62 ();
 sg13g2_fill_1 FILLER_37_79 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_decap_8 FILLER_37_111 ();
 sg13g2_decap_8 FILLER_37_118 ();
 sg13g2_fill_2 FILLER_37_125 ();
 sg13g2_fill_1 FILLER_37_127 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_fill_2 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_decap_4 FILLER_37_174 ();
 sg13g2_fill_2 FILLER_37_178 ();
 sg13g2_decap_8 FILLER_37_201 ();
 sg13g2_decap_8 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_215 ();
 sg13g2_fill_1 FILLER_37_240 ();
 sg13g2_decap_4 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_fill_1 FILLER_37_274 ();
 sg13g2_fill_1 FILLER_37_306 ();
 sg13g2_decap_8 FILLER_37_317 ();
 sg13g2_decap_8 FILLER_37_324 ();
 sg13g2_decap_8 FILLER_37_331 ();
 sg13g2_decap_8 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_345 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_decap_8 FILLER_37_359 ();
 sg13g2_decap_8 FILLER_37_366 ();
 sg13g2_decap_8 FILLER_37_373 ();
 sg13g2_decap_8 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_387 ();
 sg13g2_decap_8 FILLER_37_394 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_35 ();
 sg13g2_fill_1 FILLER_38_37 ();
 sg13g2_fill_1 FILLER_38_60 ();
 sg13g2_fill_2 FILLER_38_89 ();
 sg13g2_fill_1 FILLER_38_91 ();
 sg13g2_fill_1 FILLER_38_107 ();
 sg13g2_decap_4 FILLER_38_121 ();
 sg13g2_fill_2 FILLER_38_125 ();
 sg13g2_decap_4 FILLER_38_144 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_4 FILLER_38_161 ();
 sg13g2_fill_2 FILLER_38_165 ();
 sg13g2_decap_8 FILLER_38_171 ();
 sg13g2_decap_4 FILLER_38_178 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_decap_8 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_297 ();
 sg13g2_fill_2 FILLER_38_302 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_324 ();
 sg13g2_decap_8 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_352 ();
 sg13g2_decap_8 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_366 ();
 sg13g2_decap_8 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_4 FILLER_39_50 ();
 sg13g2_fill_2 FILLER_39_62 ();
 sg13g2_fill_1 FILLER_39_64 ();
 sg13g2_fill_2 FILLER_39_72 ();
 sg13g2_fill_1 FILLER_39_80 ();
 sg13g2_decap_8 FILLER_39_99 ();
 sg13g2_fill_1 FILLER_39_106 ();
 sg13g2_decap_4 FILLER_39_132 ();
 sg13g2_fill_1 FILLER_39_136 ();
 sg13g2_decap_8 FILLER_39_145 ();
 sg13g2_decap_8 FILLER_39_152 ();
 sg13g2_fill_2 FILLER_39_159 ();
 sg13g2_fill_1 FILLER_39_166 ();
 sg13g2_decap_4 FILLER_39_173 ();
 sg13g2_fill_2 FILLER_39_177 ();
 sg13g2_decap_4 FILLER_39_188 ();
 sg13g2_fill_1 FILLER_39_192 ();
 sg13g2_decap_8 FILLER_39_198 ();
 sg13g2_decap_4 FILLER_39_205 ();
 sg13g2_fill_1 FILLER_39_209 ();
 sg13g2_decap_8 FILLER_39_230 ();
 sg13g2_fill_1 FILLER_39_266 ();
 sg13g2_fill_2 FILLER_39_298 ();
 sg13g2_fill_1 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_324 ();
 sg13g2_decap_8 FILLER_39_331 ();
 sg13g2_decap_8 FILLER_39_338 ();
 sg13g2_decap_8 FILLER_39_345 ();
 sg13g2_decap_8 FILLER_39_352 ();
 sg13g2_decap_8 FILLER_39_359 ();
 sg13g2_decap_8 FILLER_39_366 ();
 sg13g2_decap_8 FILLER_39_373 ();
 sg13g2_decap_8 FILLER_39_380 ();
 sg13g2_decap_8 FILLER_39_387 ();
 sg13g2_decap_8 FILLER_39_394 ();
 sg13g2_decap_8 FILLER_39_401 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_4 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_60 ();
 sg13g2_decap_8 FILLER_40_67 ();
 sg13g2_fill_1 FILLER_40_82 ();
 sg13g2_fill_1 FILLER_40_87 ();
 sg13g2_decap_8 FILLER_40_96 ();
 sg13g2_decap_8 FILLER_40_103 ();
 sg13g2_fill_2 FILLER_40_110 ();
 sg13g2_fill_2 FILLER_40_134 ();
 sg13g2_fill_2 FILLER_40_158 ();
 sg13g2_fill_1 FILLER_40_160 ();
 sg13g2_fill_1 FILLER_40_174 ();
 sg13g2_decap_8 FILLER_40_186 ();
 sg13g2_decap_8 FILLER_40_198 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_fill_1 FILLER_40_231 ();
 sg13g2_fill_1 FILLER_40_248 ();
 sg13g2_fill_2 FILLER_40_253 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_fill_2 FILLER_40_273 ();
 sg13g2_fill_1 FILLER_40_275 ();
 sg13g2_fill_2 FILLER_40_310 ();
 sg13g2_fill_1 FILLER_40_312 ();
 sg13g2_decap_8 FILLER_40_348 ();
 sg13g2_decap_8 FILLER_40_355 ();
 sg13g2_decap_8 FILLER_40_362 ();
 sg13g2_decap_8 FILLER_40_369 ();
 sg13g2_decap_8 FILLER_40_376 ();
 sg13g2_decap_8 FILLER_40_383 ();
 sg13g2_decap_8 FILLER_40_390 ();
 sg13g2_decap_8 FILLER_40_397 ();
 sg13g2_decap_4 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_fill_2 FILLER_41_49 ();
 sg13g2_fill_1 FILLER_41_51 ();
 sg13g2_decap_8 FILLER_41_60 ();
 sg13g2_decap_8 FILLER_41_67 ();
 sg13g2_decap_8 FILLER_41_74 ();
 sg13g2_decap_8 FILLER_41_81 ();
 sg13g2_decap_8 FILLER_41_88 ();
 sg13g2_decap_8 FILLER_41_95 ();
 sg13g2_decap_8 FILLER_41_106 ();
 sg13g2_fill_2 FILLER_41_113 ();
 sg13g2_fill_2 FILLER_41_126 ();
 sg13g2_fill_1 FILLER_41_128 ();
 sg13g2_fill_1 FILLER_41_148 ();
 sg13g2_fill_2 FILLER_41_157 ();
 sg13g2_fill_1 FILLER_41_159 ();
 sg13g2_fill_1 FILLER_41_180 ();
 sg13g2_fill_1 FILLER_41_190 ();
 sg13g2_fill_2 FILLER_41_204 ();
 sg13g2_decap_8 FILLER_41_240 ();
 sg13g2_decap_8 FILLER_41_247 ();
 sg13g2_decap_8 FILLER_41_254 ();
 sg13g2_decap_8 FILLER_41_261 ();
 sg13g2_decap_8 FILLER_41_268 ();
 sg13g2_decap_8 FILLER_41_275 ();
 sg13g2_fill_2 FILLER_41_282 ();
 sg13g2_fill_2 FILLER_41_314 ();
 sg13g2_decap_4 FILLER_41_320 ();
 sg13g2_fill_1 FILLER_41_324 ();
 sg13g2_fill_2 FILLER_41_340 ();
 sg13g2_fill_1 FILLER_41_342 ();
 sg13g2_fill_2 FILLER_41_349 ();
 sg13g2_fill_2 FILLER_41_364 ();
 sg13g2_fill_1 FILLER_41_369 ();
 sg13g2_decap_8 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_4 FILLER_42_42 ();
 sg13g2_fill_1 FILLER_42_46 ();
 sg13g2_decap_4 FILLER_42_60 ();
 sg13g2_fill_2 FILLER_42_64 ();
 sg13g2_decap_8 FILLER_42_74 ();
 sg13g2_decap_4 FILLER_42_81 ();
 sg13g2_fill_2 FILLER_42_90 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_4 FILLER_42_126 ();
 sg13g2_fill_1 FILLER_42_130 ();
 sg13g2_fill_2 FILLER_42_143 ();
 sg13g2_fill_2 FILLER_42_155 ();
 sg13g2_fill_1 FILLER_42_157 ();
 sg13g2_fill_2 FILLER_42_171 ();
 sg13g2_fill_2 FILLER_42_187 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_4 FILLER_42_217 ();
 sg13g2_fill_1 FILLER_42_221 ();
 sg13g2_decap_8 FILLER_42_226 ();
 sg13g2_fill_1 FILLER_42_233 ();
 sg13g2_fill_2 FILLER_42_239 ();
 sg13g2_fill_1 FILLER_42_251 ();
 sg13g2_fill_2 FILLER_42_257 ();
 sg13g2_fill_1 FILLER_42_267 ();
 sg13g2_decap_8 FILLER_42_271 ();
 sg13g2_fill_2 FILLER_42_278 ();
 sg13g2_decap_8 FILLER_42_285 ();
 sg13g2_fill_2 FILLER_42_292 ();
 sg13g2_fill_1 FILLER_42_294 ();
 sg13g2_fill_1 FILLER_42_300 ();
 sg13g2_decap_4 FILLER_42_311 ();
 sg13g2_fill_1 FILLER_42_315 ();
 sg13g2_fill_2 FILLER_42_328 ();
 sg13g2_fill_1 FILLER_42_339 ();
 sg13g2_decap_8 FILLER_42_401 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_fill_2 FILLER_43_35 ();
 sg13g2_fill_2 FILLER_43_71 ();
 sg13g2_fill_1 FILLER_43_79 ();
 sg13g2_decap_4 FILLER_43_91 ();
 sg13g2_fill_2 FILLER_43_95 ();
 sg13g2_fill_2 FILLER_43_107 ();
 sg13g2_fill_1 FILLER_43_117 ();
 sg13g2_decap_8 FILLER_43_124 ();
 sg13g2_fill_2 FILLER_43_131 ();
 sg13g2_fill_1 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_143 ();
 sg13g2_decap_4 FILLER_43_150 ();
 sg13g2_fill_1 FILLER_43_154 ();
 sg13g2_fill_2 FILLER_43_159 ();
 sg13g2_decap_8 FILLER_43_169 ();
 sg13g2_fill_2 FILLER_43_176 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_fill_2 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_283 ();
 sg13g2_decap_8 FILLER_43_290 ();
 sg13g2_decap_8 FILLER_43_297 ();
 sg13g2_decap_4 FILLER_43_304 ();
 sg13g2_decap_8 FILLER_43_400 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_fill_2 FILLER_44_42 ();
 sg13g2_fill_1 FILLER_44_73 ();
 sg13g2_decap_8 FILLER_44_97 ();
 sg13g2_decap_8 FILLER_44_104 ();
 sg13g2_decap_4 FILLER_44_111 ();
 sg13g2_fill_2 FILLER_44_115 ();
 sg13g2_fill_2 FILLER_44_125 ();
 sg13g2_fill_1 FILLER_44_127 ();
 sg13g2_decap_8 FILLER_44_153 ();
 sg13g2_decap_8 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_167 ();
 sg13g2_fill_1 FILLER_44_169 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_4 FILLER_44_195 ();
 sg13g2_fill_2 FILLER_44_199 ();
 sg13g2_fill_2 FILLER_44_227 ();
 sg13g2_fill_1 FILLER_44_229 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_4 FILLER_44_245 ();
 sg13g2_fill_1 FILLER_44_249 ();
 sg13g2_decap_4 FILLER_44_258 ();
 sg13g2_fill_1 FILLER_44_262 ();
 sg13g2_fill_1 FILLER_44_267 ();
 sg13g2_fill_2 FILLER_44_272 ();
 sg13g2_decap_4 FILLER_44_279 ();
 sg13g2_fill_1 FILLER_44_283 ();
 sg13g2_decap_8 FILLER_44_288 ();
 sg13g2_decap_8 FILLER_44_295 ();
 sg13g2_decap_8 FILLER_44_302 ();
 sg13g2_decap_8 FILLER_44_309 ();
 sg13g2_decap_4 FILLER_44_316 ();
 sg13g2_fill_1 FILLER_44_320 ();
 sg13g2_decap_8 FILLER_44_330 ();
 sg13g2_fill_1 FILLER_44_366 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_fill_1 FILLER_45_49 ();
 sg13g2_fill_1 FILLER_45_55 ();
 sg13g2_decap_4 FILLER_45_69 ();
 sg13g2_fill_1 FILLER_45_73 ();
 sg13g2_decap_8 FILLER_45_79 ();
 sg13g2_fill_1 FILLER_45_86 ();
 sg13g2_fill_2 FILLER_45_97 ();
 sg13g2_fill_1 FILLER_45_99 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_fill_1 FILLER_45_112 ();
 sg13g2_decap_4 FILLER_45_127 ();
 sg13g2_decap_4 FILLER_45_151 ();
 sg13g2_fill_1 FILLER_45_155 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_fill_2 FILLER_45_182 ();
 sg13g2_fill_2 FILLER_45_230 ();
 sg13g2_fill_2 FILLER_45_266 ();
 sg13g2_fill_1 FILLER_45_268 ();
 sg13g2_decap_4 FILLER_45_274 ();
 sg13g2_fill_1 FILLER_45_292 ();
 sg13g2_decap_8 FILLER_45_327 ();
 sg13g2_decap_8 FILLER_45_334 ();
 sg13g2_fill_1 FILLER_45_341 ();
 sg13g2_fill_2 FILLER_45_348 ();
 sg13g2_fill_1 FILLER_45_391 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_fill_2 FILLER_46_35 ();
 sg13g2_fill_2 FILLER_46_53 ();
 sg13g2_fill_1 FILLER_46_55 ();
 sg13g2_decap_4 FILLER_46_70 ();
 sg13g2_fill_2 FILLER_46_82 ();
 sg13g2_fill_2 FILLER_46_92 ();
 sg13g2_decap_8 FILLER_46_122 ();
 sg13g2_fill_2 FILLER_46_129 ();
 sg13g2_fill_1 FILLER_46_131 ();
 sg13g2_fill_2 FILLER_46_157 ();
 sg13g2_fill_2 FILLER_46_174 ();
 sg13g2_fill_1 FILLER_46_176 ();
 sg13g2_decap_8 FILLER_46_187 ();
 sg13g2_decap_8 FILLER_46_194 ();
 sg13g2_fill_2 FILLER_46_201 ();
 sg13g2_fill_1 FILLER_46_246 ();
 sg13g2_fill_2 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_337 ();
 sg13g2_decap_4 FILLER_46_344 ();
 sg13g2_fill_1 FILLER_46_369 ();
 sg13g2_fill_2 FILLER_46_398 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_fill_2 FILLER_47_28 ();
 sg13g2_fill_1 FILLER_47_30 ();
 sg13g2_fill_2 FILLER_47_57 ();
 sg13g2_fill_1 FILLER_47_59 ();
 sg13g2_fill_2 FILLER_47_70 ();
 sg13g2_fill_1 FILLER_47_72 ();
 sg13g2_fill_2 FILLER_47_78 ();
 sg13g2_decap_8 FILLER_47_131 ();
 sg13g2_decap_4 FILLER_47_138 ();
 sg13g2_fill_1 FILLER_47_147 ();
 sg13g2_decap_4 FILLER_47_153 ();
 sg13g2_fill_1 FILLER_47_179 ();
 sg13g2_decap_8 FILLER_47_192 ();
 sg13g2_decap_8 FILLER_47_199 ();
 sg13g2_fill_2 FILLER_47_206 ();
 sg13g2_fill_1 FILLER_47_213 ();
 sg13g2_decap_8 FILLER_47_219 ();
 sg13g2_decap_4 FILLER_47_230 ();
 sg13g2_fill_1 FILLER_47_234 ();
 sg13g2_decap_4 FILLER_47_239 ();
 sg13g2_fill_1 FILLER_47_243 ();
 sg13g2_decap_8 FILLER_47_249 ();
 sg13g2_decap_4 FILLER_47_276 ();
 sg13g2_fill_1 FILLER_47_316 ();
 sg13g2_fill_2 FILLER_47_381 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_60 ();
 sg13g2_decap_8 FILLER_48_67 ();
 sg13g2_decap_4 FILLER_48_74 ();
 sg13g2_fill_2 FILLER_48_100 ();
 sg13g2_decap_8 FILLER_48_106 ();
 sg13g2_decap_4 FILLER_48_120 ();
 sg13g2_fill_2 FILLER_48_124 ();
 sg13g2_fill_2 FILLER_48_131 ();
 sg13g2_fill_2 FILLER_48_143 ();
 sg13g2_fill_1 FILLER_48_145 ();
 sg13g2_fill_1 FILLER_48_152 ();
 sg13g2_decap_8 FILLER_48_158 ();
 sg13g2_decap_8 FILLER_48_165 ();
 sg13g2_decap_8 FILLER_48_172 ();
 sg13g2_decap_4 FILLER_48_179 ();
 sg13g2_fill_1 FILLER_48_183 ();
 sg13g2_decap_8 FILLER_48_192 ();
 sg13g2_decap_8 FILLER_48_199 ();
 sg13g2_fill_1 FILLER_48_206 ();
 sg13g2_decap_8 FILLER_48_233 ();
 sg13g2_decap_8 FILLER_48_240 ();
 sg13g2_decap_4 FILLER_48_247 ();
 sg13g2_fill_1 FILLER_48_251 ();
 sg13g2_decap_4 FILLER_48_256 ();
 sg13g2_fill_2 FILLER_48_264 ();
 sg13g2_fill_1 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_297 ();
 sg13g2_fill_2 FILLER_48_304 ();
 sg13g2_fill_1 FILLER_48_306 ();
 sg13g2_fill_2 FILLER_48_312 ();
 sg13g2_fill_1 FILLER_48_346 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_54 ();
 sg13g2_decap_4 FILLER_49_61 ();
 sg13g2_fill_1 FILLER_49_65 ();
 sg13g2_fill_2 FILLER_49_71 ();
 sg13g2_fill_1 FILLER_49_73 ();
 sg13g2_decap_8 FILLER_49_79 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_fill_1 FILLER_49_119 ();
 sg13g2_fill_1 FILLER_49_129 ();
 sg13g2_fill_2 FILLER_49_135 ();
 sg13g2_fill_1 FILLER_49_142 ();
 sg13g2_fill_2 FILLER_49_148 ();
 sg13g2_decap_8 FILLER_49_156 ();
 sg13g2_fill_2 FILLER_49_163 ();
 sg13g2_decap_4 FILLER_49_175 ();
 sg13g2_fill_2 FILLER_49_184 ();
 sg13g2_decap_8 FILLER_49_194 ();
 sg13g2_decap_8 FILLER_49_227 ();
 sg13g2_decap_8 FILLER_49_234 ();
 sg13g2_decap_4 FILLER_49_241 ();
 sg13g2_fill_2 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_265 ();
 sg13g2_decap_8 FILLER_49_272 ();
 sg13g2_decap_8 FILLER_49_279 ();
 sg13g2_decap_8 FILLER_49_286 ();
 sg13g2_fill_1 FILLER_49_293 ();
 sg13g2_fill_1 FILLER_49_298 ();
 sg13g2_fill_1 FILLER_49_309 ();
 sg13g2_fill_1 FILLER_49_320 ();
 sg13g2_fill_2 FILLER_49_329 ();
 sg13g2_fill_1 FILLER_49_339 ();
 sg13g2_fill_2 FILLER_49_398 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_fill_1 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_53 ();
 sg13g2_fill_1 FILLER_50_60 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_4 FILLER_50_84 ();
 sg13g2_fill_1 FILLER_50_88 ();
 sg13g2_decap_8 FILLER_50_96 ();
 sg13g2_decap_8 FILLER_50_103 ();
 sg13g2_decap_4 FILLER_50_120 ();
 sg13g2_fill_1 FILLER_50_129 ();
 sg13g2_fill_1 FILLER_50_176 ();
 sg13g2_decap_4 FILLER_50_199 ();
 sg13g2_fill_2 FILLER_50_203 ();
 sg13g2_decap_8 FILLER_50_218 ();
 sg13g2_fill_2 FILLER_50_225 ();
 sg13g2_decap_4 FILLER_50_232 ();
 sg13g2_fill_2 FILLER_50_236 ();
 sg13g2_fill_2 FILLER_50_268 ();
 sg13g2_decap_8 FILLER_50_275 ();
 sg13g2_decap_8 FILLER_50_282 ();
 sg13g2_decap_8 FILLER_50_326 ();
 sg13g2_decap_8 FILLER_50_333 ();
 sg13g2_fill_2 FILLER_50_340 ();
 sg13g2_fill_2 FILLER_50_354 ();
 sg13g2_fill_1 FILLER_50_369 ();
 sg13g2_fill_1 FILLER_50_386 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_35 ();
 sg13g2_fill_1 FILLER_51_65 ();
 sg13g2_decap_4 FILLER_51_80 ();
 sg13g2_fill_1 FILLER_51_84 ();
 sg13g2_fill_2 FILLER_51_90 ();
 sg13g2_fill_1 FILLER_51_103 ();
 sg13g2_fill_1 FILLER_51_122 ();
 sg13g2_decap_4 FILLER_51_130 ();
 sg13g2_fill_2 FILLER_51_161 ();
 sg13g2_fill_1 FILLER_51_175 ();
 sg13g2_fill_2 FILLER_51_181 ();
 sg13g2_fill_1 FILLER_51_183 ();
 sg13g2_decap_4 FILLER_51_196 ();
 sg13g2_fill_1 FILLER_51_200 ();
 sg13g2_decap_4 FILLER_51_209 ();
 sg13g2_fill_1 FILLER_51_213 ();
 sg13g2_fill_1 FILLER_51_219 ();
 sg13g2_fill_2 FILLER_51_242 ();
 sg13g2_fill_1 FILLER_51_249 ();
 sg13g2_fill_2 FILLER_51_268 ();
 sg13g2_fill_1 FILLER_51_313 ();
 sg13g2_decap_8 FILLER_51_345 ();
 sg13g2_decap_8 FILLER_51_352 ();
 sg13g2_decap_8 FILLER_51_359 ();
 sg13g2_fill_2 FILLER_51_366 ();
 sg13g2_fill_1 FILLER_51_368 ();
 sg13g2_fill_1 FILLER_51_375 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_4 FILLER_52_35 ();
 sg13g2_fill_2 FILLER_52_39 ();
 sg13g2_fill_1 FILLER_52_50 ();
 sg13g2_fill_1 FILLER_52_65 ();
 sg13g2_fill_2 FILLER_52_76 ();
 sg13g2_decap_8 FILLER_52_99 ();
 sg13g2_decap_4 FILLER_52_106 ();
 sg13g2_decap_4 FILLER_52_131 ();
 sg13g2_fill_2 FILLER_52_135 ();
 sg13g2_fill_2 FILLER_52_142 ();
 sg13g2_fill_1 FILLER_52_144 ();
 sg13g2_decap_8 FILLER_52_150 ();
 sg13g2_decap_8 FILLER_52_157 ();
 sg13g2_decap_8 FILLER_52_164 ();
 sg13g2_decap_8 FILLER_52_171 ();
 sg13g2_decap_8 FILLER_52_178 ();
 sg13g2_decap_8 FILLER_52_185 ();
 sg13g2_fill_2 FILLER_52_220 ();
 sg13g2_fill_1 FILLER_52_222 ();
 sg13g2_fill_2 FILLER_52_231 ();
 sg13g2_fill_1 FILLER_52_269 ();
 sg13g2_decap_8 FILLER_52_302 ();
 sg13g2_fill_1 FILLER_52_309 ();
 sg13g2_decap_8 FILLER_52_314 ();
 sg13g2_fill_1 FILLER_52_321 ();
 sg13g2_decap_4 FILLER_52_348 ();
 sg13g2_fill_1 FILLER_52_381 ();
 sg13g2_fill_1 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_4 FILLER_53_28 ();
 sg13g2_decap_4 FILLER_53_87 ();
 sg13g2_fill_2 FILLER_53_109 ();
 sg13g2_fill_2 FILLER_53_123 ();
 sg13g2_fill_2 FILLER_53_131 ();
 sg13g2_fill_1 FILLER_53_133 ();
 sg13g2_fill_1 FILLER_53_142 ();
 sg13g2_decap_8 FILLER_53_151 ();
 sg13g2_fill_1 FILLER_53_158 ();
 sg13g2_fill_1 FILLER_53_167 ();
 sg13g2_decap_8 FILLER_53_177 ();
 sg13g2_decap_8 FILLER_53_192 ();
 sg13g2_decap_4 FILLER_53_199 ();
 sg13g2_fill_1 FILLER_53_203 ();
 sg13g2_decap_4 FILLER_53_217 ();
 sg13g2_fill_2 FILLER_53_261 ();
 sg13g2_fill_1 FILLER_53_263 ();
 sg13g2_fill_1 FILLER_53_270 ();
 sg13g2_decap_8 FILLER_53_294 ();
 sg13g2_decap_8 FILLER_53_301 ();
 sg13g2_decap_8 FILLER_53_308 ();
 sg13g2_decap_4 FILLER_53_315 ();
 sg13g2_decap_8 FILLER_53_323 ();
 sg13g2_decap_4 FILLER_53_338 ();
 sg13g2_fill_1 FILLER_53_342 ();
 sg13g2_fill_2 FILLER_53_375 ();
 sg13g2_fill_1 FILLER_53_382 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_4 FILLER_54_35 ();
 sg13g2_fill_1 FILLER_54_39 ();
 sg13g2_fill_1 FILLER_54_50 ();
 sg13g2_fill_2 FILLER_54_67 ();
 sg13g2_fill_1 FILLER_54_69 ();
 sg13g2_fill_1 FILLER_54_75 ();
 sg13g2_decap_4 FILLER_54_80 ();
 sg13g2_fill_2 FILLER_54_84 ();
 sg13g2_fill_2 FILLER_54_98 ();
 sg13g2_decap_4 FILLER_54_118 ();
 sg13g2_fill_2 FILLER_54_122 ();
 sg13g2_decap_4 FILLER_54_133 ();
 sg13g2_fill_1 FILLER_54_137 ();
 sg13g2_decap_4 FILLER_54_155 ();
 sg13g2_decap_8 FILLER_54_183 ();
 sg13g2_decap_8 FILLER_54_198 ();
 sg13g2_decap_8 FILLER_54_205 ();
 sg13g2_fill_2 FILLER_54_212 ();
 sg13g2_fill_1 FILLER_54_214 ();
 sg13g2_decap_8 FILLER_54_222 ();
 sg13g2_fill_2 FILLER_54_229 ();
 sg13g2_decap_4 FILLER_54_244 ();
 sg13g2_fill_2 FILLER_54_248 ();
 sg13g2_fill_2 FILLER_54_262 ();
 sg13g2_decap_4 FILLER_54_268 ();
 sg13g2_fill_2 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_292 ();
 sg13g2_decap_8 FILLER_54_297 ();
 sg13g2_decap_4 FILLER_54_307 ();
 sg13g2_fill_1 FILLER_54_311 ();
 sg13g2_fill_2 FILLER_54_317 ();
 sg13g2_fill_1 FILLER_54_324 ();
 sg13g2_fill_1 FILLER_54_351 ();
 sg13g2_fill_2 FILLER_54_361 ();
 sg13g2_fill_1 FILLER_54_399 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_4 FILLER_55_42 ();
 sg13g2_fill_1 FILLER_55_46 ();
 sg13g2_decap_4 FILLER_55_52 ();
 sg13g2_decap_8 FILLER_55_66 ();
 sg13g2_decap_8 FILLER_55_73 ();
 sg13g2_fill_1 FILLER_55_85 ();
 sg13g2_fill_2 FILLER_55_91 ();
 sg13g2_decap_4 FILLER_55_104 ();
 sg13g2_decap_8 FILLER_55_113 ();
 sg13g2_fill_1 FILLER_55_129 ();
 sg13g2_decap_8 FILLER_55_134 ();
 sg13g2_decap_8 FILLER_55_141 ();
 sg13g2_decap_8 FILLER_55_148 ();
 sg13g2_fill_2 FILLER_55_155 ();
 sg13g2_fill_2 FILLER_55_162 ();
 sg13g2_decap_8 FILLER_55_174 ();
 sg13g2_fill_2 FILLER_55_181 ();
 sg13g2_decap_4 FILLER_55_207 ();
 sg13g2_decap_8 FILLER_55_229 ();
 sg13g2_decap_8 FILLER_55_236 ();
 sg13g2_decap_8 FILLER_55_243 ();
 sg13g2_fill_2 FILLER_55_250 ();
 sg13g2_fill_1 FILLER_55_252 ();
 sg13g2_fill_1 FILLER_55_261 ();
 sg13g2_decap_8 FILLER_55_269 ();
 sg13g2_decap_8 FILLER_55_276 ();
 sg13g2_decap_4 FILLER_55_283 ();
 sg13g2_decap_4 FILLER_55_322 ();
 sg13g2_fill_1 FILLER_55_326 ();
 sg13g2_decap_4 FILLER_55_331 ();
 sg13g2_fill_1 FILLER_55_335 ();
 sg13g2_decap_8 FILLER_55_340 ();
 sg13g2_fill_1 FILLER_55_347 ();
 sg13g2_fill_2 FILLER_55_376 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_4 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_60 ();
 sg13g2_decap_8 FILLER_56_67 ();
 sg13g2_fill_1 FILLER_56_74 ();
 sg13g2_fill_2 FILLER_56_80 ();
 sg13g2_fill_2 FILLER_56_97 ();
 sg13g2_fill_1 FILLER_56_99 ();
 sg13g2_fill_2 FILLER_56_118 ();
 sg13g2_fill_1 FILLER_56_120 ();
 sg13g2_fill_2 FILLER_56_131 ();
 sg13g2_fill_1 FILLER_56_133 ();
 sg13g2_fill_2 FILLER_56_144 ();
 sg13g2_fill_1 FILLER_56_146 ();
 sg13g2_decap_8 FILLER_56_156 ();
 sg13g2_decap_4 FILLER_56_163 ();
 sg13g2_fill_2 FILLER_56_172 ();
 sg13g2_decap_8 FILLER_56_192 ();
 sg13g2_decap_8 FILLER_56_199 ();
 sg13g2_fill_1 FILLER_56_206 ();
 sg13g2_fill_1 FILLER_56_226 ();
 sg13g2_decap_8 FILLER_56_239 ();
 sg13g2_decap_4 FILLER_56_246 ();
 sg13g2_fill_2 FILLER_56_250 ();
 sg13g2_decap_4 FILLER_56_260 ();
 sg13g2_decap_8 FILLER_56_272 ();
 sg13g2_decap_8 FILLER_56_279 ();
 sg13g2_decap_8 FILLER_56_286 ();
 sg13g2_fill_1 FILLER_56_315 ();
 sg13g2_decap_8 FILLER_56_345 ();
 sg13g2_decap_4 FILLER_56_352 ();
 sg13g2_fill_1 FILLER_56_356 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_fill_1 FILLER_57_35 ();
 sg13g2_fill_1 FILLER_57_50 ();
 sg13g2_fill_2 FILLER_57_64 ();
 sg13g2_decap_4 FILLER_57_76 ();
 sg13g2_fill_2 FILLER_57_80 ();
 sg13g2_decap_8 FILLER_57_90 ();
 sg13g2_decap_8 FILLER_57_97 ();
 sg13g2_fill_2 FILLER_57_109 ();
 sg13g2_fill_1 FILLER_57_111 ();
 sg13g2_fill_1 FILLER_57_136 ();
 sg13g2_fill_2 FILLER_57_160 ();
 sg13g2_fill_1 FILLER_57_162 ();
 sg13g2_fill_1 FILLER_57_171 ();
 sg13g2_decap_8 FILLER_57_200 ();
 sg13g2_decap_8 FILLER_57_225 ();
 sg13g2_decap_8 FILLER_57_275 ();
 sg13g2_decap_4 FILLER_57_287 ();
 sg13g2_fill_2 FILLER_57_291 ();
 sg13g2_decap_4 FILLER_57_313 ();
 sg13g2_decap_8 FILLER_57_327 ();
 sg13g2_fill_1 FILLER_57_334 ();
 sg13g2_decap_8 FILLER_57_356 ();
 sg13g2_decap_4 FILLER_57_363 ();
 sg13g2_fill_1 FILLER_57_367 ();
 sg13g2_fill_2 FILLER_57_372 ();
 sg13g2_fill_1 FILLER_57_374 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_fill_1 FILLER_58_42 ();
 sg13g2_fill_2 FILLER_58_68 ();
 sg13g2_fill_1 FILLER_58_70 ();
 sg13g2_decap_4 FILLER_58_84 ();
 sg13g2_decap_4 FILLER_58_98 ();
 sg13g2_decap_4 FILLER_58_115 ();
 sg13g2_fill_2 FILLER_58_119 ();
 sg13g2_decap_4 FILLER_58_125 ();
 sg13g2_fill_2 FILLER_58_139 ();
 sg13g2_decap_4 FILLER_58_166 ();
 sg13g2_fill_1 FILLER_58_181 ();
 sg13g2_decap_8 FILLER_58_200 ();
 sg13g2_fill_1 FILLER_58_207 ();
 sg13g2_decap_4 FILLER_58_219 ();
 sg13g2_fill_1 FILLER_58_223 ();
 sg13g2_fill_1 FILLER_58_230 ();
 sg13g2_fill_2 FILLER_58_261 ();
 sg13g2_fill_1 FILLER_58_263 ();
 sg13g2_fill_2 FILLER_58_272 ();
 sg13g2_decap_8 FILLER_58_300 ();
 sg13g2_decap_8 FILLER_58_307 ();
 sg13g2_fill_2 FILLER_58_314 ();
 sg13g2_fill_1 FILLER_58_316 ();
 sg13g2_fill_2 FILLER_58_335 ();
 sg13g2_fill_2 FILLER_58_342 ();
 sg13g2_fill_2 FILLER_58_370 ();
 sg13g2_fill_1 FILLER_58_372 ();
 sg13g2_fill_1 FILLER_58_385 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_fill_2 FILLER_59_79 ();
 sg13g2_decap_4 FILLER_59_86 ();
 sg13g2_fill_2 FILLER_59_109 ();
 sg13g2_fill_1 FILLER_59_111 ();
 sg13g2_fill_1 FILLER_59_117 ();
 sg13g2_fill_1 FILLER_59_137 ();
 sg13g2_fill_2 FILLER_59_143 ();
 sg13g2_fill_2 FILLER_59_149 ();
 sg13g2_fill_1 FILLER_59_169 ();
 sg13g2_decap_8 FILLER_59_175 ();
 sg13g2_decap_8 FILLER_59_182 ();
 sg13g2_decap_4 FILLER_59_189 ();
 sg13g2_fill_2 FILLER_59_193 ();
 sg13g2_decap_8 FILLER_59_203 ();
 sg13g2_fill_2 FILLER_59_210 ();
 sg13g2_decap_8 FILLER_59_221 ();
 sg13g2_decap_4 FILLER_59_228 ();
 sg13g2_fill_1 FILLER_59_236 ();
 sg13g2_decap_8 FILLER_59_253 ();
 sg13g2_decap_8 FILLER_59_260 ();
 sg13g2_decap_8 FILLER_59_267 ();
 sg13g2_fill_1 FILLER_59_274 ();
 sg13g2_fill_2 FILLER_59_283 ();
 sg13g2_decap_8 FILLER_59_289 ();
 sg13g2_decap_8 FILLER_59_296 ();
 sg13g2_decap_4 FILLER_59_303 ();
 sg13g2_decap_4 FILLER_59_319 ();
 sg13g2_decap_8 FILLER_59_363 ();
 sg13g2_decap_4 FILLER_59_370 ();
 sg13g2_fill_1 FILLER_59_374 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_fill_2 FILLER_60_42 ();
 sg13g2_fill_2 FILLER_60_49 ();
 sg13g2_fill_1 FILLER_60_51 ();
 sg13g2_fill_1 FILLER_60_62 ();
 sg13g2_fill_2 FILLER_60_82 ();
 sg13g2_fill_1 FILLER_60_84 ();
 sg13g2_fill_2 FILLER_60_95 ();
 sg13g2_fill_1 FILLER_60_97 ();
 sg13g2_decap_4 FILLER_60_103 ();
 sg13g2_fill_1 FILLER_60_107 ();
 sg13g2_fill_1 FILLER_60_117 ();
 sg13g2_decap_8 FILLER_60_128 ();
 sg13g2_decap_8 FILLER_60_135 ();
 sg13g2_decap_8 FILLER_60_142 ();
 sg13g2_fill_1 FILLER_60_149 ();
 sg13g2_decap_8 FILLER_60_165 ();
 sg13g2_decap_8 FILLER_60_172 ();
 sg13g2_decap_8 FILLER_60_179 ();
 sg13g2_decap_4 FILLER_60_186 ();
 sg13g2_fill_1 FILLER_60_190 ();
 sg13g2_fill_2 FILLER_60_199 ();
 sg13g2_fill_1 FILLER_60_201 ();
 sg13g2_fill_2 FILLER_60_207 ();
 sg13g2_fill_1 FILLER_60_209 ();
 sg13g2_decap_4 FILLER_60_223 ();
 sg13g2_fill_2 FILLER_60_227 ();
 sg13g2_fill_1 FILLER_60_234 ();
 sg13g2_decap_4 FILLER_60_244 ();
 sg13g2_fill_2 FILLER_60_248 ();
 sg13g2_decap_4 FILLER_60_262 ();
 sg13g2_fill_2 FILLER_60_266 ();
 sg13g2_decap_4 FILLER_60_273 ();
 sg13g2_fill_1 FILLER_60_277 ();
 sg13g2_decap_8 FILLER_60_286 ();
 sg13g2_fill_2 FILLER_60_293 ();
 sg13g2_fill_2 FILLER_60_339 ();
 sg13g2_decap_8 FILLER_60_344 ();
 sg13g2_decap_4 FILLER_60_351 ();
 sg13g2_fill_2 FILLER_60_381 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_50 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_fill_1 FILLER_61_69 ();
 sg13g2_decap_8 FILLER_61_95 ();
 sg13g2_decap_8 FILLER_61_102 ();
 sg13g2_fill_1 FILLER_61_109 ();
 sg13g2_decap_4 FILLER_61_123 ();
 sg13g2_fill_2 FILLER_61_127 ();
 sg13g2_decap_8 FILLER_61_141 ();
 sg13g2_decap_4 FILLER_61_148 ();
 sg13g2_fill_2 FILLER_61_152 ();
 sg13g2_decap_8 FILLER_61_163 ();
 sg13g2_fill_2 FILLER_61_170 ();
 sg13g2_fill_2 FILLER_61_188 ();
 sg13g2_decap_8 FILLER_61_232 ();
 sg13g2_fill_1 FILLER_61_239 ();
 sg13g2_fill_2 FILLER_61_292 ();
 sg13g2_fill_1 FILLER_61_294 ();
 sg13g2_fill_2 FILLER_61_301 ();
 sg13g2_fill_1 FILLER_61_335 ();
 sg13g2_fill_1 FILLER_61_364 ();
 sg13g2_decap_8 FILLER_61_369 ();
 sg13g2_fill_1 FILLER_61_376 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_4 FILLER_62_42 ();
 sg13g2_decap_4 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_64 ();
 sg13g2_fill_2 FILLER_62_71 ();
 sg13g2_fill_1 FILLER_62_73 ();
 sg13g2_decap_8 FILLER_62_94 ();
 sg13g2_fill_1 FILLER_62_101 ();
 sg13g2_decap_4 FILLER_62_127 ();
 sg13g2_fill_1 FILLER_62_139 ();
 sg13g2_fill_1 FILLER_62_160 ();
 sg13g2_decap_8 FILLER_62_166 ();
 sg13g2_decap_8 FILLER_62_173 ();
 sg13g2_decap_4 FILLER_62_180 ();
 sg13g2_fill_1 FILLER_62_184 ();
 sg13g2_decap_8 FILLER_62_204 ();
 sg13g2_decap_8 FILLER_62_211 ();
 sg13g2_decap_8 FILLER_62_218 ();
 sg13g2_decap_8 FILLER_62_229 ();
 sg13g2_decap_4 FILLER_62_236 ();
 sg13g2_decap_8 FILLER_62_249 ();
 sg13g2_fill_2 FILLER_62_282 ();
 sg13g2_fill_1 FILLER_62_284 ();
 sg13g2_decap_8 FILLER_62_337 ();
 sg13g2_decap_8 FILLER_62_344 ();
 sg13g2_decap_4 FILLER_62_351 ();
 sg13g2_fill_1 FILLER_62_355 ();
 sg13g2_decap_8 FILLER_62_361 ();
 sg13g2_decap_8 FILLER_62_368 ();
 sg13g2_decap_8 FILLER_62_375 ();
 sg13g2_fill_1 FILLER_62_382 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_4 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_fill_1 FILLER_63_77 ();
 sg13g2_decap_4 FILLER_63_83 ();
 sg13g2_decap_8 FILLER_63_93 ();
 sg13g2_decap_8 FILLER_63_100 ();
 sg13g2_fill_2 FILLER_63_107 ();
 sg13g2_fill_1 FILLER_63_117 ();
 sg13g2_fill_2 FILLER_63_132 ();
 sg13g2_fill_1 FILLER_63_134 ();
 sg13g2_decap_8 FILLER_63_152 ();
 sg13g2_decap_8 FILLER_63_159 ();
 sg13g2_decap_8 FILLER_63_166 ();
 sg13g2_fill_2 FILLER_63_173 ();
 sg13g2_fill_1 FILLER_63_175 ();
 sg13g2_fill_1 FILLER_63_193 ();
 sg13g2_fill_2 FILLER_63_199 ();
 sg13g2_fill_1 FILLER_63_201 ();
 sg13g2_decap_4 FILLER_63_207 ();
 sg13g2_fill_2 FILLER_63_219 ();
 sg13g2_fill_1 FILLER_63_221 ();
 sg13g2_decap_8 FILLER_63_257 ();
 sg13g2_fill_2 FILLER_63_264 ();
 sg13g2_decap_4 FILLER_63_293 ();
 sg13g2_fill_1 FILLER_63_297 ();
 sg13g2_fill_2 FILLER_63_312 ();
 sg13g2_fill_1 FILLER_63_319 ();
 sg13g2_decap_8 FILLER_63_324 ();
 sg13g2_decap_4 FILLER_63_331 ();
 sg13g2_fill_2 FILLER_63_335 ();
 sg13g2_fill_1 FILLER_63_385 ();
 sg13g2_fill_1 FILLER_63_399 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_fill_1 FILLER_64_49 ();
 sg13g2_fill_2 FILLER_64_55 ();
 sg13g2_fill_1 FILLER_64_57 ();
 sg13g2_fill_2 FILLER_64_74 ();
 sg13g2_fill_1 FILLER_64_76 ();
 sg13g2_fill_2 FILLER_64_84 ();
 sg13g2_fill_1 FILLER_64_86 ();
 sg13g2_decap_8 FILLER_64_93 ();
 sg13g2_decap_8 FILLER_64_100 ();
 sg13g2_decap_8 FILLER_64_107 ();
 sg13g2_decap_4 FILLER_64_114 ();
 sg13g2_fill_2 FILLER_64_118 ();
 sg13g2_decap_4 FILLER_64_125 ();
 sg13g2_fill_1 FILLER_64_129 ();
 sg13g2_fill_1 FILLER_64_150 ();
 sg13g2_fill_2 FILLER_64_189 ();
 sg13g2_fill_1 FILLER_64_229 ();
 sg13g2_decap_8 FILLER_64_260 ();
 sg13g2_decap_8 FILLER_64_267 ();
 sg13g2_decap_8 FILLER_64_274 ();
 sg13g2_decap_8 FILLER_64_281 ();
 sg13g2_decap_8 FILLER_64_288 ();
 sg13g2_decap_8 FILLER_64_295 ();
 sg13g2_decap_4 FILLER_64_302 ();
 sg13g2_fill_1 FILLER_64_306 ();
 sg13g2_fill_1 FILLER_64_311 ();
 sg13g2_decap_4 FILLER_64_317 ();
 sg13g2_fill_1 FILLER_64_321 ();
 sg13g2_decap_8 FILLER_64_337 ();
 sg13g2_decap_4 FILLER_64_344 ();
 sg13g2_fill_1 FILLER_64_352 ();
 sg13g2_decap_8 FILLER_64_363 ();
 sg13g2_decap_8 FILLER_64_374 ();
 sg13g2_decap_4 FILLER_64_381 ();
 sg13g2_decap_4 FILLER_64_391 ();
 sg13g2_fill_1 FILLER_64_395 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_fill_1 FILLER_65_49 ();
 sg13g2_decap_4 FILLER_65_73 ();
 sg13g2_fill_1 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_99 ();
 sg13g2_decap_4 FILLER_65_118 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_4 FILLER_65_133 ();
 sg13g2_fill_1 FILLER_65_137 ();
 sg13g2_decap_8 FILLER_65_159 ();
 sg13g2_fill_1 FILLER_65_166 ();
 sg13g2_fill_2 FILLER_65_175 ();
 sg13g2_fill_1 FILLER_65_177 ();
 sg13g2_fill_2 FILLER_65_186 ();
 sg13g2_fill_1 FILLER_65_188 ();
 sg13g2_fill_2 FILLER_65_198 ();
 sg13g2_fill_1 FILLER_65_200 ();
 sg13g2_fill_1 FILLER_65_206 ();
 sg13g2_fill_2 FILLER_65_212 ();
 sg13g2_fill_1 FILLER_65_214 ();
 sg13g2_decap_8 FILLER_65_249 ();
 sg13g2_fill_1 FILLER_65_256 ();
 sg13g2_decap_8 FILLER_65_273 ();
 sg13g2_decap_8 FILLER_65_283 ();
 sg13g2_decap_4 FILLER_65_290 ();
 sg13g2_fill_1 FILLER_65_294 ();
 sg13g2_fill_1 FILLER_65_316 ();
 sg13g2_fill_1 FILLER_65_350 ();
 sg13g2_decap_4 FILLER_65_370 ();
 sg13g2_fill_1 FILLER_65_374 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_4 FILLER_66_49 ();
 sg13g2_fill_2 FILLER_66_53 ();
 sg13g2_fill_1 FILLER_66_73 ();
 sg13g2_fill_1 FILLER_66_120 ();
 sg13g2_decap_8 FILLER_66_136 ();
 sg13g2_decap_8 FILLER_66_143 ();
 sg13g2_decap_8 FILLER_66_150 ();
 sg13g2_fill_1 FILLER_66_157 ();
 sg13g2_fill_2 FILLER_66_163 ();
 sg13g2_fill_1 FILLER_66_165 ();
 sg13g2_decap_8 FILLER_66_179 ();
 sg13g2_decap_8 FILLER_66_186 ();
 sg13g2_decap_8 FILLER_66_193 ();
 sg13g2_decap_8 FILLER_66_200 ();
 sg13g2_fill_1 FILLER_66_207 ();
 sg13g2_fill_1 FILLER_66_224 ();
 sg13g2_fill_2 FILLER_66_243 ();
 sg13g2_fill_1 FILLER_66_271 ();
 sg13g2_fill_2 FILLER_66_307 ();
 sg13g2_fill_2 FILLER_66_339 ();
 sg13g2_fill_2 FILLER_66_381 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_fill_1 FILLER_67_63 ();
 sg13g2_fill_2 FILLER_67_70 ();
 sg13g2_fill_2 FILLER_67_76 ();
 sg13g2_fill_1 FILLER_67_78 ();
 sg13g2_fill_1 FILLER_67_97 ();
 sg13g2_decap_4 FILLER_67_104 ();
 sg13g2_fill_1 FILLER_67_108 ();
 sg13g2_fill_1 FILLER_67_115 ();
 sg13g2_decap_8 FILLER_67_130 ();
 sg13g2_decap_4 FILLER_67_137 ();
 sg13g2_fill_1 FILLER_67_141 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_fill_1 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_180 ();
 sg13g2_fill_1 FILLER_67_187 ();
 sg13g2_decap_8 FILLER_67_249 ();
 sg13g2_fill_2 FILLER_67_260 ();
 sg13g2_decap_4 FILLER_67_299 ();
 sg13g2_fill_2 FILLER_67_329 ();
 sg13g2_decap_4 FILLER_67_368 ();
 sg13g2_fill_2 FILLER_67_372 ();
 sg13g2_fill_1 FILLER_67_399 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_fill_2 FILLER_68_63 ();
 sg13g2_fill_1 FILLER_68_65 ();
 sg13g2_decap_8 FILLER_68_71 ();
 sg13g2_decap_4 FILLER_68_78 ();
 sg13g2_fill_2 FILLER_68_82 ();
 sg13g2_decap_4 FILLER_68_105 ();
 sg13g2_fill_2 FILLER_68_117 ();
 sg13g2_fill_1 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_125 ();
 sg13g2_decap_8 FILLER_68_132 ();
 sg13g2_fill_2 FILLER_68_139 ();
 sg13g2_decap_8 FILLER_68_150 ();
 sg13g2_fill_2 FILLER_68_173 ();
 sg13g2_decap_8 FILLER_68_200 ();
 sg13g2_fill_2 FILLER_68_207 ();
 sg13g2_fill_2 FILLER_68_214 ();
 sg13g2_decap_8 FILLER_68_299 ();
 sg13g2_decap_8 FILLER_68_306 ();
 sg13g2_fill_1 FILLER_68_313 ();
 sg13g2_fill_2 FILLER_68_318 ();
 sg13g2_decap_8 FILLER_68_378 ();
 sg13g2_decap_8 FILLER_68_385 ();
 sg13g2_decap_4 FILLER_68_392 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_89 ();
 sg13g2_fill_1 FILLER_69_96 ();
 sg13g2_decap_4 FILLER_69_102 ();
 sg13g2_fill_1 FILLER_69_106 ();
 sg13g2_fill_1 FILLER_69_131 ();
 sg13g2_decap_4 FILLER_69_154 ();
 sg13g2_fill_1 FILLER_69_158 ();
 sg13g2_fill_2 FILLER_69_173 ();
 sg13g2_fill_1 FILLER_69_175 ();
 sg13g2_decap_8 FILLER_69_197 ();
 sg13g2_decap_4 FILLER_69_204 ();
 sg13g2_fill_2 FILLER_69_208 ();
 sg13g2_fill_1 FILLER_69_236 ();
 sg13g2_fill_1 FILLER_69_247 ();
 sg13g2_fill_2 FILLER_69_264 ();
 sg13g2_fill_2 FILLER_69_289 ();
 sg13g2_fill_1 FILLER_69_291 ();
 sg13g2_decap_8 FILLER_69_305 ();
 sg13g2_decap_4 FILLER_69_312 ();
 sg13g2_fill_1 FILLER_69_325 ();
 sg13g2_decap_8 FILLER_69_384 ();
 sg13g2_decap_8 FILLER_69_391 ();
 sg13g2_decap_4 FILLER_69_398 ();
 sg13g2_fill_1 FILLER_69_402 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_4 FILLER_70_112 ();
 sg13g2_fill_1 FILLER_70_116 ();
 sg13g2_fill_2 FILLER_70_127 ();
 sg13g2_fill_1 FILLER_70_129 ();
 sg13g2_fill_1 FILLER_70_144 ();
 sg13g2_fill_2 FILLER_70_163 ();
 sg13g2_fill_1 FILLER_70_165 ();
 sg13g2_decap_8 FILLER_70_170 ();
 sg13g2_decap_4 FILLER_70_177 ();
 sg13g2_decap_8 FILLER_70_191 ();
 sg13g2_decap_8 FILLER_70_198 ();
 sg13g2_decap_4 FILLER_70_205 ();
 sg13g2_fill_2 FILLER_70_235 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_decap_8 FILLER_70_300 ();
 sg13g2_fill_1 FILLER_70_307 ();
 sg13g2_decap_4 FILLER_70_331 ();
 sg13g2_fill_1 FILLER_70_373 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_4 FILLER_71_138 ();
 sg13g2_fill_2 FILLER_71_171 ();
 sg13g2_fill_1 FILLER_71_173 ();
 sg13g2_decap_8 FILLER_71_181 ();
 sg13g2_decap_4 FILLER_71_188 ();
 sg13g2_decap_8 FILLER_71_197 ();
 sg13g2_fill_2 FILLER_71_204 ();
 sg13g2_decap_8 FILLER_71_210 ();
 sg13g2_fill_2 FILLER_71_217 ();
 sg13g2_decap_4 FILLER_71_223 ();
 sg13g2_fill_1 FILLER_71_236 ();
 sg13g2_fill_1 FILLER_71_242 ();
 sg13g2_fill_1 FILLER_71_304 ();
 sg13g2_fill_1 FILLER_71_338 ();
 sg13g2_fill_2 FILLER_71_365 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_4 FILLER_72_119 ();
 sg13g2_fill_1 FILLER_72_123 ();
 sg13g2_decap_4 FILLER_72_132 ();
 sg13g2_fill_2 FILLER_72_136 ();
 sg13g2_fill_1 FILLER_72_167 ();
 sg13g2_fill_1 FILLER_72_184 ();
 sg13g2_decap_8 FILLER_72_221 ();
 sg13g2_fill_2 FILLER_72_254 ();
 sg13g2_fill_1 FILLER_72_256 ();
 sg13g2_fill_1 FILLER_72_262 ();
 sg13g2_fill_1 FILLER_72_271 ();
 sg13g2_fill_2 FILLER_72_303 ();
 sg13g2_decap_4 FILLER_72_321 ();
 sg13g2_fill_1 FILLER_72_340 ();
 sg13g2_fill_2 FILLER_72_345 ();
 sg13g2_fill_1 FILLER_72_354 ();
 sg13g2_fill_1 FILLER_72_381 ();
 sg13g2_fill_2 FILLER_72_398 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_fill_2 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_4 FILLER_73_161 ();
 sg13g2_fill_1 FILLER_73_165 ();
 sg13g2_fill_2 FILLER_73_184 ();
 sg13g2_decap_8 FILLER_73_222 ();
 sg13g2_decap_8 FILLER_73_229 ();
 sg13g2_fill_1 FILLER_73_236 ();
 sg13g2_decap_4 FILLER_73_250 ();
 sg13g2_fill_1 FILLER_73_258 ();
 sg13g2_decap_4 FILLER_73_289 ();
 sg13g2_fill_2 FILLER_73_293 ();
 sg13g2_fill_2 FILLER_73_341 ();
 sg13g2_decap_4 FILLER_73_360 ();
 sg13g2_fill_2 FILLER_73_364 ();
 sg13g2_decap_4 FILLER_73_370 ();
 sg13g2_fill_2 FILLER_73_374 ();
 sg13g2_fill_1 FILLER_73_380 ();
 sg13g2_fill_2 FILLER_73_386 ();
 sg13g2_fill_1 FILLER_73_388 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_fill_2 FILLER_74_175 ();
 sg13g2_fill_1 FILLER_74_177 ();
 sg13g2_decap_4 FILLER_74_190 ();
 sg13g2_fill_2 FILLER_74_194 ();
 sg13g2_fill_2 FILLER_74_201 ();
 sg13g2_fill_1 FILLER_74_203 ();
 sg13g2_fill_1 FILLER_74_239 ();
 sg13g2_decap_8 FILLER_74_244 ();
 sg13g2_decap_8 FILLER_74_251 ();
 sg13g2_decap_8 FILLER_74_258 ();
 sg13g2_decap_8 FILLER_74_265 ();
 sg13g2_fill_2 FILLER_74_272 ();
 sg13g2_decap_8 FILLER_74_278 ();
 sg13g2_decap_8 FILLER_74_285 ();
 sg13g2_decap_8 FILLER_74_292 ();
 sg13g2_decap_4 FILLER_74_299 ();
 sg13g2_fill_2 FILLER_74_303 ();
 sg13g2_decap_8 FILLER_74_309 ();
 sg13g2_decap_4 FILLER_74_326 ();
 sg13g2_decap_8 FILLER_74_356 ();
 sg13g2_fill_2 FILLER_74_363 ();
 sg13g2_decap_8 FILLER_74_391 ();
 sg13g2_decap_8 FILLER_74_398 ();
 sg13g2_decap_4 FILLER_74_405 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_4 FILLER_75_175 ();
 sg13g2_fill_2 FILLER_75_179 ();
 sg13g2_decap_8 FILLER_75_186 ();
 sg13g2_decap_4 FILLER_75_193 ();
 sg13g2_fill_1 FILLER_75_201 ();
 sg13g2_fill_1 FILLER_75_206 ();
 sg13g2_decap_8 FILLER_75_211 ();
 sg13g2_fill_1 FILLER_75_231 ();
 sg13g2_fill_2 FILLER_75_236 ();
 sg13g2_fill_1 FILLER_75_238 ();
 sg13g2_fill_2 FILLER_75_243 ();
 sg13g2_decap_8 FILLER_75_271 ();
 sg13g2_fill_2 FILLER_75_278 ();
 sg13g2_fill_1 FILLER_75_280 ();
 sg13g2_decap_4 FILLER_75_289 ();
 sg13g2_decap_8 FILLER_75_298 ();
 sg13g2_decap_8 FILLER_75_305 ();
 sg13g2_decap_8 FILLER_75_347 ();
 sg13g2_decap_4 FILLER_75_354 ();
 sg13g2_fill_1 FILLER_75_358 ();
 sg13g2_fill_1 FILLER_75_368 ();
 sg13g2_decap_8 FILLER_75_378 ();
 sg13g2_fill_2 FILLER_75_385 ();
 sg13g2_fill_1 FILLER_75_387 ();
 sg13g2_decap_8 FILLER_75_395 ();
 sg13g2_decap_8 FILLER_75_402 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_4 FILLER_76_168 ();
 sg13g2_fill_2 FILLER_76_172 ();
 sg13g2_fill_1 FILLER_76_195 ();
 sg13g2_decap_8 FILLER_76_201 ();
 sg13g2_fill_2 FILLER_76_208 ();
 sg13g2_fill_1 FILLER_76_210 ();
 sg13g2_decap_4 FILLER_76_215 ();
 sg13g2_fill_2 FILLER_76_232 ();
 sg13g2_fill_1 FILLER_76_234 ();
 sg13g2_decap_4 FILLER_76_270 ();
 sg13g2_fill_2 FILLER_76_274 ();
 sg13g2_fill_1 FILLER_76_297 ();
 sg13g2_fill_1 FILLER_76_308 ();
 sg13g2_fill_2 FILLER_76_318 ();
 sg13g2_decap_4 FILLER_76_339 ();
 sg13g2_decap_4 FILLER_76_374 ();
 sg13g2_fill_2 FILLER_76_378 ();
 sg13g2_fill_2 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_4 FILLER_77_161 ();
 sg13g2_fill_2 FILLER_77_165 ();
 sg13g2_fill_2 FILLER_77_197 ();
 sg13g2_fill_1 FILLER_77_199 ();
 sg13g2_fill_1 FILLER_77_267 ();
 sg13g2_decap_8 FILLER_77_324 ();
 sg13g2_decap_8 FILLER_77_331 ();
 sg13g2_decap_8 FILLER_77_338 ();
 sg13g2_fill_2 FILLER_77_345 ();
 sg13g2_fill_2 FILLER_77_352 ();
 sg13g2_fill_1 FILLER_77_354 ();
 sg13g2_decap_8 FILLER_77_401 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_fill_1 FILLER_78_161 ();
 sg13g2_fill_2 FILLER_78_233 ();
 sg13g2_fill_1 FILLER_78_235 ();
 sg13g2_decap_8 FILLER_78_253 ();
 sg13g2_fill_1 FILLER_78_260 ();
 sg13g2_fill_2 FILLER_78_287 ();
 sg13g2_fill_2 FILLER_78_312 ();
 sg13g2_fill_1 FILLER_78_323 ();
 sg13g2_fill_1 FILLER_78_350 ();
 sg13g2_decap_4 FILLER_78_403 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_fill_1 FILLER_79_228 ();
 sg13g2_fill_2 FILLER_79_234 ();
 sg13g2_fill_1 FILLER_79_236 ();
 sg13g2_fill_2 FILLER_79_263 ();
 sg13g2_fill_2 FILLER_79_291 ();
 sg13g2_fill_1 FILLER_79_293 ();
 sg13g2_decap_8 FILLER_79_390 ();
 sg13g2_decap_8 FILLER_79_397 ();
 sg13g2_decap_4 FILLER_79_404 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_fill_1 FILLER_80_187 ();
 sg13g2_fill_1 FILLER_80_193 ();
 sg13g2_decap_8 FILLER_80_202 ();
 sg13g2_fill_2 FILLER_80_213 ();
 sg13g2_fill_1 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_225 ();
 sg13g2_decap_8 FILLER_80_232 ();
 sg13g2_decap_8 FILLER_80_239 ();
 sg13g2_fill_2 FILLER_80_246 ();
 sg13g2_decap_8 FILLER_80_252 ();
 sg13g2_decap_8 FILLER_80_259 ();
 sg13g2_decap_4 FILLER_80_266 ();
 sg13g2_fill_2 FILLER_80_287 ();
 sg13g2_fill_2 FILLER_80_293 ();
 sg13g2_fill_1 FILLER_80_304 ();
 sg13g2_decap_4 FILLER_80_309 ();
 sg13g2_fill_1 FILLER_80_313 ();
 sg13g2_fill_1 FILLER_80_335 ();
 sg13g2_fill_2 FILLER_80_348 ();
 sg13g2_fill_1 FILLER_80_350 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_fill_2 FILLER_80_365 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net11;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net13;
 assign uio_out[0] = net14;
 assign uio_out[1] = net15;
 assign uio_out[2] = net16;
 assign uio_out[3] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
endmodule
