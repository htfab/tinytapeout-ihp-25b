module tt_um_gamepad_pmod_demo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire clknet_0_clk;
 wire \driver.decoder.data_reg[0] ;
 wire \driver.decoder.data_reg[10] ;
 wire \driver.decoder.data_reg[11] ;
 wire \driver.decoder.data_reg[1] ;
 wire \driver.decoder.data_reg[2] ;
 wire \driver.decoder.data_reg[3] ;
 wire \driver.decoder.data_reg[4] ;
 wire \driver.decoder.data_reg[5] ;
 wire \driver.decoder.data_reg[6] ;
 wire \driver.decoder.data_reg[7] ;
 wire \driver.decoder.data_reg[8] ;
 wire \driver.decoder.data_reg[9] ;
 wire \driver.driver.pmod_clk_prev ;
 wire \driver.driver.pmod_clk_sync[0] ;
 wire \driver.driver.pmod_clk_sync[1] ;
 wire \driver.driver.pmod_data_sync[0] ;
 wire \driver.driver.pmod_data_sync[1] ;
 wire \driver.driver.pmod_latch_prev ;
 wire \driver.driver.pmod_latch_sync[0] ;
 wire \driver.driver.pmod_latch_sync[1] ;
 wire \driver.driver.shift_reg[0] ;
 wire \driver.driver.shift_reg[10] ;
 wire \driver.driver.shift_reg[11] ;
 wire \driver.driver.shift_reg[1] ;
 wire \driver.driver.shift_reg[2] ;
 wire \driver.driver.shift_reg[3] ;
 wire \driver.driver.shift_reg[4] ;
 wire \driver.driver.shift_reg[5] ;
 wire \driver.driver.shift_reg[6] ;
 wire \driver.driver.shift_reg[7] ;
 wire \driver.driver.shift_reg[8] ;
 wire \driver.driver.shift_reg[9] ;
 wire hsync;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire \vga_sync_gen.vsync ;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;

 sg13g2_inv_1 _0643_ (.Y(_0071_),
    .A(net132));
 sg13g2_inv_1 _0644_ (.Y(_0072_),
    .A(net126));
 sg13g2_inv_1 _0645_ (.Y(_0073_),
    .A(net130));
 sg13g2_inv_1 _0646_ (.Y(_0074_),
    .A(net110));
 sg13g2_inv_1 _0647_ (.Y(_0075_),
    .A(net112));
 sg13g2_inv_1 _0648_ (.Y(_0076_),
    .A(net138));
 sg13g2_inv_1 _0649_ (.Y(_0077_),
    .A(net124));
 sg13g2_inv_1 _0650_ (.Y(_0078_),
    .A(net128));
 sg13g2_inv_1 _0651_ (.Y(_0079_),
    .A(net140));
 sg13g2_inv_1 _0652_ (.Y(_0080_),
    .A(net114));
 sg13g2_inv_1 _0653_ (.Y(_0081_),
    .A(\driver.driver.shift_reg[0] ));
 sg13g2_inv_1 _0654_ (.Y(_0082_),
    .A(net93));
 sg13g2_inv_1 _0655_ (.Y(_0083_),
    .A(net84));
 sg13g2_inv_1 _0656_ (.Y(_0084_),
    .A(net91));
 sg13g2_inv_1 _0657_ (.Y(_0085_),
    .A(net190));
 sg13g2_inv_1 _0658_ (.Y(_0086_),
    .A(net195));
 sg13g2_inv_2 _0659_ (.Y(_0087_),
    .A(net197));
 sg13g2_inv_1 _0660_ (.Y(_0088_),
    .A(net201));
 sg13g2_inv_1 _0661_ (.Y(_0089_),
    .A(net211));
 sg13g2_inv_2 _0662_ (.Y(_0090_),
    .A(\pix_x[2] ));
 sg13g2_inv_1 _0663_ (.Y(_0091_),
    .A(\pix_x[3] ));
 sg13g2_inv_1 _0664_ (.Y(_0092_),
    .A(_0011_));
 sg13g2_inv_1 _0665_ (.Y(_0093_),
    .A(net116));
 sg13g2_inv_1 _0666_ (.Y(_0094_),
    .A(net104));
 sg13g2_inv_1 _0667_ (.Y(_0095_),
    .A(net106));
 sg13g2_inv_1 _0668_ (.Y(_0096_),
    .A(net118));
 sg13g2_inv_1 _0669_ (.Y(_0097_),
    .A(net98));
 sg13g2_inv_1 _0670_ (.Y(_0098_),
    .A(net108));
 sg13g2_inv_1 _0671_ (.Y(_0099_),
    .A(net100));
 sg13g2_inv_1 _0672_ (.Y(_0100_),
    .A(net89));
 sg13g2_inv_1 _0673_ (.Y(_0101_),
    .A(net120));
 sg13g2_inv_1 _0674_ (.Y(_0102_),
    .A(net102));
 sg13g2_inv_1 _0675_ (.Y(_0103_),
    .A(net122));
 sg13g2_inv_1 _0676_ (.Y(_0104_),
    .A(net136));
 sg13g2_nand3_1 _0677_ (.B(net194),
    .C(net195),
    .A(\pix_y[7] ),
    .Y(_0105_));
 sg13g2_nor2b_1 _0678_ (.A(\pix_y[9] ),
    .B_N(net190),
    .Y(_0106_));
 sg13g2_nand2b_2 _0679_ (.Y(_0107_),
    .B(net190),
    .A_N(net188));
 sg13g2_nand4_1 _0680_ (.B(_0088_),
    .C(net199),
    .A(_0087_),
    .Y(_0108_),
    .D(net134));
 sg13g2_nor3_1 _0681_ (.A(_0105_),
    .B(_0107_),
    .C(net143),
    .Y(_0001_));
 sg13g2_and2_1 _0682_ (.A(\pix_x[8] ),
    .B(\pix_x[9] ),
    .X(_0109_));
 sg13g2_nand2_1 _0683_ (.Y(_0110_),
    .A(\pix_x[8] ),
    .B(\pix_x[9] ));
 sg13g2_nor2_1 _0684_ (.A(net205),
    .B(net207),
    .Y(_0111_));
 sg13g2_or2_1 _0685_ (.X(_0112_),
    .B(net206),
    .A(net204));
 sg13g2_and2_1 _0686_ (.A(net203),
    .B(\pix_x[9] ),
    .X(_0113_));
 sg13g2_o21ai_1 _0687_ (.B1(_0113_),
    .Y(_0114_),
    .A1(net209),
    .A2(_0112_));
 sg13g2_nor2b_2 _0688_ (.A(\pix_x[8] ),
    .B_N(\pix_x[9] ),
    .Y(_0115_));
 sg13g2_nand2_1 _0689_ (.Y(_0116_),
    .A(net206),
    .B(net209));
 sg13g2_and2_1 _0690_ (.A(net202),
    .B(net204),
    .X(_0117_));
 sg13g2_nand2b_1 _0691_ (.Y(_0118_),
    .B(_0117_),
    .A_N(_0116_));
 sg13g2_a21oi_1 _0692_ (.A1(_0115_),
    .A2(_0118_),
    .Y(_0119_),
    .B1(net80));
 sg13g2_a21oi_1 _0693_ (.A1(_0110_),
    .A2(_0114_),
    .Y(_0000_),
    .B1(_0119_));
 sg13g2_nand4_1 _0694_ (.B(net102),
    .C(net122),
    .A(net120),
    .Y(_0120_),
    .D(net136));
 sg13g2_nand4_1 _0695_ (.B(net108),
    .C(net100),
    .A(net98),
    .Y(_0121_),
    .D(net89));
 sg13g2_nand4_1 _0696_ (.B(net104),
    .C(net106),
    .A(net116),
    .Y(_0122_),
    .D(net118));
 sg13g2_nor3_2 _0697_ (.A(_0120_),
    .B(_0121_),
    .C(_0122_),
    .Y(_0123_));
 sg13g2_inv_1 _0698_ (.Y(_0124_),
    .A(_0123_));
 sg13g2_nand2_2 _0699_ (.Y(_0125_),
    .A(net197),
    .B(net198));
 sg13g2_nor2b_1 _0700_ (.A(net193),
    .B_N(net195),
    .Y(_0126_));
 sg13g2_nand2b_1 _0701_ (.Y(_0127_),
    .B(net195),
    .A_N(net194));
 sg13g2_mux2_1 _0702_ (.A0(_0126_),
    .A1(net193),
    .S(_0125_),
    .X(_0128_));
 sg13g2_nor2_1 _0703_ (.A(net202),
    .B(net204),
    .Y(_0129_));
 sg13g2_nor3_2 _0704_ (.A(net203),
    .B(net204),
    .C(net206),
    .Y(_0130_));
 sg13g2_nor2_2 _0705_ (.A(net189),
    .B(net188),
    .Y(_0131_));
 sg13g2_inv_1 _0706_ (.Y(_0132_),
    .A(_0131_));
 sg13g2_nand2_1 _0707_ (.Y(_0133_),
    .A(\pix_y[7] ),
    .B(_0131_));
 sg13g2_and4_1 _0708_ (.A(net191),
    .B(_0115_),
    .C(_0130_),
    .D(_0131_),
    .X(_0134_));
 sg13g2_and3_2 _0709_ (.X(_0135_),
    .A(_0105_),
    .B(_0128_),
    .C(_0134_));
 sg13g2_nand3_1 _0710_ (.B(_0128_),
    .C(_0134_),
    .A(_0105_),
    .Y(_0136_));
 sg13g2_nand2_2 _0711_ (.Y(_0137_),
    .A(net200),
    .B(net198));
 sg13g2_nand2_2 _0712_ (.Y(_0138_),
    .A(net196),
    .B(net197));
 sg13g2_nand3_1 _0713_ (.B(net196),
    .C(net197),
    .A(net194),
    .Y(_0139_));
 sg13g2_or2_1 _0714_ (.X(_0140_),
    .B(_0139_),
    .A(_0137_));
 sg13g2_nand2b_1 _0715_ (.Y(_0141_),
    .B(\pix_y[4] ),
    .A_N(net195));
 sg13g2_nand2b_1 _0716_ (.Y(_0142_),
    .B(_0137_),
    .A_N(_0141_));
 sg13g2_nor2_1 _0717_ (.A(net195),
    .B(\pix_y[4] ),
    .Y(_0143_));
 sg13g2_or2_2 _0718_ (.X(_0144_),
    .B(\pix_y[4] ),
    .A(net196));
 sg13g2_nor2b_2 _0719_ (.A(net191),
    .B_N(net193),
    .Y(_0145_));
 sg13g2_nand2b_1 _0720_ (.Y(_0146_),
    .B(net194),
    .A_N(net191));
 sg13g2_nor4_2 _0721_ (.A(net189),
    .B(net188),
    .C(_0143_),
    .Y(_0147_),
    .D(_0146_));
 sg13g2_nor2_1 _0722_ (.A(net191),
    .B(net193),
    .Y(_0148_));
 sg13g2_or2_1 _0723_ (.X(_0149_),
    .B(net194),
    .A(net191));
 sg13g2_nand2_1 _0724_ (.Y(_0150_),
    .A(net193),
    .B(_0086_));
 sg13g2_a21oi_1 _0725_ (.A1(net193),
    .A2(_0144_),
    .Y(_0151_),
    .B1(net191));
 sg13g2_and3_1 _0726_ (.X(_0152_),
    .A(_0140_),
    .B(_0142_),
    .C(_0147_));
 sg13g2_nand3_1 _0727_ (.B(_0142_),
    .C(_0147_),
    .A(_0140_),
    .Y(_0153_));
 sg13g2_nor2_1 _0728_ (.A(\pix_x[8] ),
    .B(\pix_x[9] ),
    .Y(_0154_));
 sg13g2_or2_1 _0729_ (.X(_0155_),
    .B(\pix_x[9] ),
    .A(\pix_x[8] ));
 sg13g2_and3_1 _0730_ (.X(_0156_),
    .A(net206),
    .B(_0129_),
    .C(_0154_));
 sg13g2_nand3_1 _0731_ (.B(_0129_),
    .C(_0154_),
    .A(net206),
    .Y(_0157_));
 sg13g2_and4_2 _0732_ (.A(_0140_),
    .B(_0142_),
    .C(_0147_),
    .D(_0156_),
    .X(_0158_));
 sg13g2_nand4_1 _0733_ (.B(_0142_),
    .C(_0147_),
    .A(_0140_),
    .Y(_0159_),
    .D(_0156_));
 sg13g2_nand2_2 _0734_ (.Y(_0160_),
    .A(_0005_),
    .B(_0115_));
 sg13g2_nand2b_1 _0735_ (.Y(_0161_),
    .B(net207),
    .A_N(\pix_x[4] ));
 sg13g2_xor2_1 _0736_ (.B(net208),
    .A(net207),
    .X(_0162_));
 sg13g2_nand2b_1 _0737_ (.Y(_0163_),
    .B(net204),
    .A_N(net202));
 sg13g2_o21ai_1 _0738_ (.B1(net204),
    .Y(_0164_),
    .A1(net207),
    .A2(net208));
 sg13g2_nand2_2 _0739_ (.Y(_0165_),
    .A(net205),
    .B(_0162_));
 sg13g2_nor3_2 _0740_ (.A(net203),
    .B(_0160_),
    .C(_0165_),
    .Y(_0166_));
 sg13g2_or3_1 _0741_ (.A(net202),
    .B(_0160_),
    .C(_0165_),
    .X(_0167_));
 sg13g2_nor2_2 _0742_ (.A(_0153_),
    .B(_0167_),
    .Y(_0168_));
 sg13g2_nand2_1 _0743_ (.Y(_0169_),
    .A(_0152_),
    .B(_0166_));
 sg13g2_a21oi_2 _0744_ (.B1(_0158_),
    .Y(_0170_),
    .A2(_0166_),
    .A1(_0152_));
 sg13g2_a221oi_1 _0745_ (.B2(_0167_),
    .C1(_0153_),
    .B1(_0157_),
    .A1(net201),
    .Y(_0171_),
    .A2(net199));
 sg13g2_xor2_1 _0746_ (.B(_0171_),
    .A(_0015_),
    .X(_0172_));
 sg13g2_or2_1 _0747_ (.X(_0173_),
    .B(net198),
    .A(net197));
 sg13g2_nand2_1 _0748_ (.Y(_0174_),
    .A(_0125_),
    .B(_0173_));
 sg13g2_and2_1 _0749_ (.A(_0106_),
    .B(_0115_),
    .X(_0175_));
 sg13g2_nand2_1 _0750_ (.Y(_0176_),
    .A(net197),
    .B(_0131_));
 sg13g2_nand4_1 _0751_ (.B(_0141_),
    .C(_0175_),
    .A(_0130_),
    .Y(_0177_),
    .D(_0176_));
 sg13g2_a21oi_1 _0752_ (.A1(_0148_),
    .A2(_0173_),
    .Y(_0178_),
    .B1(_0086_));
 sg13g2_nor2_1 _0753_ (.A(\pix_y[1] ),
    .B(\pix_y[0] ),
    .Y(_0179_));
 sg13g2_or2_1 _0754_ (.X(_0180_),
    .B(\pix_y[0] ),
    .A(net134));
 sg13g2_nand2b_1 _0755_ (.Y(_0181_),
    .B(\pix_y[5] ),
    .A_N(net200));
 sg13g2_o21ai_1 _0756_ (.B1(_0131_),
    .Y(_0182_),
    .A1(_0180_),
    .A2(_0181_));
 sg13g2_o21ai_1 _0757_ (.B1(_0086_),
    .Y(_0183_),
    .A1(net198),
    .A2(_0146_));
 sg13g2_nand3b_1 _0758_ (.B(_0182_),
    .C(_0183_),
    .Y(_0184_),
    .A_N(_0178_));
 sg13g2_nor2_2 _0759_ (.A(_0177_),
    .B(_0184_),
    .Y(_0185_));
 sg13g2_a21oi_1 _0760_ (.A1(_0135_),
    .A2(_0174_),
    .Y(_0186_),
    .B1(_0185_));
 sg13g2_nor2b_1 _0761_ (.A(net200),
    .B_N(net198),
    .Y(_0187_));
 sg13g2_o21ai_1 _0762_ (.B1(net199),
    .Y(_0188_),
    .A1(net200),
    .A2(_0180_));
 sg13g2_nor2_1 _0763_ (.A(_0107_),
    .B(_0149_),
    .Y(_0189_));
 sg13g2_and3_1 _0764_ (.X(_0190_),
    .A(_0106_),
    .B(_0138_),
    .C(_0148_));
 sg13g2_o21ai_1 _0765_ (.B1(_0190_),
    .Y(_0191_),
    .A1(_0086_),
    .A2(_0188_));
 sg13g2_nand4_1 _0766_ (.B(_0087_),
    .C(_0179_),
    .A(net195),
    .Y(_0192_),
    .D(_0187_));
 sg13g2_nor3_1 _0767_ (.A(_0107_),
    .B(_0149_),
    .C(_0192_),
    .Y(_0193_));
 sg13g2_a21oi_1 _0768_ (.A1(_0132_),
    .A2(_0191_),
    .Y(_0194_),
    .B1(_0193_));
 sg13g2_a21o_1 _0769_ (.A2(_0191_),
    .A1(_0132_),
    .B1(_0193_),
    .X(_0195_));
 sg13g2_nand4_1 _0770_ (.B(_0145_),
    .C(_0179_),
    .A(_0143_),
    .Y(_0196_),
    .D(_0187_));
 sg13g2_nand4_1 _0771_ (.B(_0130_),
    .C(_0151_),
    .A(_0115_),
    .Y(_0197_),
    .D(_0196_));
 sg13g2_a21oi_1 _0772_ (.A1(_0106_),
    .A2(_0188_),
    .Y(_0198_),
    .B1(_0189_));
 sg13g2_nor2_1 _0773_ (.A(_0197_),
    .B(_0198_),
    .Y(_0199_));
 sg13g2_nor3_2 _0774_ (.A(_0194_),
    .B(_0197_),
    .C(_0198_),
    .Y(_0200_));
 sg13g2_o21ai_1 _0775_ (.B1(net179),
    .Y(_0201_),
    .A1(_0177_),
    .A2(_0184_));
 sg13g2_o21ai_1 _0776_ (.B1(_0186_),
    .Y(_0202_),
    .A1(_0135_),
    .A2(_0172_));
 sg13g2_nor2_1 _0777_ (.A(net202),
    .B(_0155_),
    .Y(_0203_));
 sg13g2_nor2b_1 _0778_ (.A(_0007_),
    .B_N(net205),
    .Y(_0204_));
 sg13g2_or2_1 _0779_ (.X(_0205_),
    .B(net149),
    .A(\pix_x[1] ));
 sg13g2_or3_2 _0780_ (.A(\pix_x[2] ),
    .B(\pix_x[1] ),
    .C(\pix_x[0] ),
    .X(_0206_));
 sg13g2_nor4_1 _0781_ (.A(net210),
    .B(_0161_),
    .C(_0163_),
    .D(_0206_),
    .Y(_0207_));
 sg13g2_o21ai_1 _0782_ (.B1(_0203_),
    .Y(_0208_),
    .A1(_0204_),
    .A2(_0207_));
 sg13g2_nor3_2 _0783_ (.A(_0133_),
    .B(_0150_),
    .C(_0208_),
    .Y(_0209_));
 sg13g2_nand2b_1 _0784_ (.Y(_0210_),
    .B(net189),
    .A_N(net192));
 sg13g2_o21ai_1 _0785_ (.B1(_0189_),
    .Y(_0211_),
    .A1(net193),
    .A2(net195));
 sg13g2_nor2_1 _0786_ (.A(_0208_),
    .B(_0211_),
    .Y(_0212_));
 sg13g2_or2_2 _0787_ (.X(_0213_),
    .B(net176),
    .A(_0209_));
 sg13g2_a21oi_1 _0788_ (.A1(_0174_),
    .A2(_0200_),
    .Y(_0214_),
    .B1(_0213_));
 sg13g2_a22oi_1 _0789_ (.Y(_0215_),
    .B1(_0214_),
    .B2(_0202_),
    .A2(_0213_),
    .A1(_0087_));
 sg13g2_inv_2 _0790_ (.Y(_0216_),
    .A(net166));
 sg13g2_or2_1 _0791_ (.X(_0217_),
    .B(net199),
    .A(net201));
 sg13g2_a221oi_1 _0792_ (.B2(_0217_),
    .C1(_0201_),
    .B1(_0171_),
    .A1(net199),
    .Y(_0218_),
    .A2(net178));
 sg13g2_nor2b_1 _0793_ (.A(_0014_),
    .B_N(_0201_),
    .Y(_0219_));
 sg13g2_or2_1 _0794_ (.X(_0220_),
    .B(_0219_),
    .A(_0218_));
 sg13g2_nor2_1 _0795_ (.A(_0218_),
    .B(_0219_),
    .Y(_0221_));
 sg13g2_nor2b_2 _0796_ (.A(_0008_),
    .B_N(_0209_),
    .Y(_0222_));
 sg13g2_o21ai_1 _0797_ (.B1(_0012_),
    .Y(_0223_),
    .A1(_0137_),
    .A2(_0141_));
 sg13g2_nand2_1 _0798_ (.Y(_0224_),
    .A(_0145_),
    .B(_0223_));
 sg13g2_a21oi_1 _0799_ (.A1(_0145_),
    .A2(_0223_),
    .Y(_0225_),
    .B1(_0092_));
 sg13g2_xor2_1 _0800_ (.B(_0225_),
    .A(_0009_),
    .X(_0226_));
 sg13g2_xor2_1 _0801_ (.B(_0125_),
    .A(_0012_),
    .X(_0227_));
 sg13g2_nor2_1 _0802_ (.A(net200),
    .B(_0012_),
    .Y(_0228_));
 sg13g2_a21oi_1 _0803_ (.A1(net200),
    .A2(_0227_),
    .Y(_0229_),
    .B1(_0228_));
 sg13g2_nor2_1 _0804_ (.A(net189),
    .B(_0009_),
    .Y(_0230_));
 sg13g2_nor2b_1 _0805_ (.A(net193),
    .B_N(net191),
    .Y(_0231_));
 sg13g2_nand2b_1 _0806_ (.Y(_0232_),
    .B(_0231_),
    .A_N(_0223_));
 sg13g2_a221oi_1 _0807_ (.B2(_0224_),
    .C1(_0229_),
    .B1(_0232_),
    .A1(_0008_),
    .Y(_0233_),
    .A2(_0230_));
 sg13g2_a21oi_1 _0808_ (.A1(_0226_),
    .A2(_0233_),
    .Y(_0234_),
    .B1(net178));
 sg13g2_o21ai_1 _0809_ (.B1(net179),
    .Y(_0235_),
    .A1(_0008_),
    .A2(_0230_));
 sg13g2_nand2b_1 _0810_ (.Y(_0236_),
    .B(_0010_),
    .A_N(net192));
 sg13g2_nand2b_1 _0811_ (.Y(_0237_),
    .B(net192),
    .A_N(_0010_));
 sg13g2_a22oi_1 _0812_ (.Y(_0238_),
    .B1(_0237_),
    .B2(_0144_),
    .A2(_0236_),
    .A1(_0138_));
 sg13g2_nand4_1 _0813_ (.B(net194),
    .C(net196),
    .A(net192),
    .Y(_0239_),
    .D(net197));
 sg13g2_xor2_1 _0814_ (.B(_0239_),
    .A(_0009_),
    .X(_0240_));
 sg13g2_nand3_1 _0815_ (.B(_0238_),
    .C(_0240_),
    .A(_0008_),
    .Y(_0241_));
 sg13g2_a21o_1 _0816_ (.A2(_0241_),
    .A1(net178),
    .B1(_0235_),
    .X(_0242_));
 sg13g2_o21ai_1 _0817_ (.B1(_0010_),
    .Y(_0243_),
    .A1(_0125_),
    .A2(_0127_));
 sg13g2_nand2_1 _0818_ (.Y(_0244_),
    .A(net189),
    .B(_0008_));
 sg13g2_o21ai_1 _0819_ (.B1(_0009_),
    .Y(_0245_),
    .A1(net189),
    .A2(_0008_));
 sg13g2_nand3_1 _0820_ (.B(_0243_),
    .C(_0244_),
    .A(net191),
    .Y(_0246_));
 sg13g2_nand3b_1 _0821_ (.B(_0008_),
    .C(_0010_),
    .Y(_0247_),
    .A_N(net192));
 sg13g2_nor2_1 _0822_ (.A(_0009_),
    .B(_0247_),
    .Y(_0248_));
 sg13g2_o21ai_1 _0823_ (.B1(_0248_),
    .Y(_0249_),
    .A1(_0125_),
    .A2(_0127_));
 sg13g2_o21ai_1 _0824_ (.B1(_0249_),
    .Y(_0250_),
    .A1(_0245_),
    .A2(_0246_));
 sg13g2_nor2_1 _0825_ (.A(net179),
    .B(_0227_),
    .Y(_0251_));
 sg13g2_a22oi_1 _0826_ (.Y(_0252_),
    .B1(_0250_),
    .B2(_0251_),
    .A2(_0199_),
    .A1(_0195_));
 sg13g2_o21ai_1 _0827_ (.B1(_0252_),
    .Y(_0253_),
    .A1(_0234_),
    .A2(_0242_));
 sg13g2_a21oi_1 _0828_ (.A1(_0010_),
    .A2(_0011_),
    .Y(_0254_),
    .B1(_0150_));
 sg13g2_a21oi_1 _0829_ (.A1(_0247_),
    .A2(_0254_),
    .Y(_0255_),
    .B1(_0173_));
 sg13g2_a21oi_1 _0830_ (.A1(_0010_),
    .A2(_0210_),
    .Y(_0256_),
    .B1(_0011_));
 sg13g2_nor3_1 _0831_ (.A(_0092_),
    .B(_0127_),
    .C(_0244_),
    .Y(_0257_));
 sg13g2_a21oi_1 _0832_ (.A1(_0236_),
    .A2(_0244_),
    .Y(_0258_),
    .B1(_0173_));
 sg13g2_nor2_1 _0833_ (.A(_0257_),
    .B(_0258_),
    .Y(_0259_));
 sg13g2_or3_1 _0834_ (.A(_0255_),
    .B(_0256_),
    .C(_0259_),
    .X(_0260_));
 sg13g2_a21oi_1 _0835_ (.A1(_0200_),
    .A2(_0260_),
    .Y(_0261_),
    .B1(net176));
 sg13g2_a221oi_1 _0836_ (.B2(_0253_),
    .C1(_0209_),
    .B1(_0261_),
    .A1(net176),
    .Y(_0262_),
    .A2(_0257_));
 sg13g2_nor2_2 _0837_ (.A(_0222_),
    .B(_0262_),
    .Y(_0263_));
 sg13g2_o21ai_1 _0838_ (.B1(_0088_),
    .Y(_0264_),
    .A1(_0153_),
    .A2(_0167_));
 sg13g2_nand3_1 _0839_ (.B(_0152_),
    .C(_0166_),
    .A(net201),
    .Y(_0265_));
 sg13g2_a21oi_2 _0840_ (.B1(_0158_),
    .Y(_0266_),
    .A2(_0265_),
    .A1(_0264_));
 sg13g2_nor2_2 _0841_ (.A(_0013_),
    .B(_0159_),
    .Y(_0267_));
 sg13g2_nor2_2 _0842_ (.A(_0266_),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_or2_1 _0843_ (.X(_0269_),
    .B(_0267_),
    .A(_0266_));
 sg13g2_nor3_1 _0844_ (.A(_0222_),
    .B(_0262_),
    .C(net167),
    .Y(_0270_));
 sg13g2_nor3_2 _0845_ (.A(_0107_),
    .B(_0144_),
    .C(_0149_),
    .Y(_0271_));
 sg13g2_nor3_2 _0846_ (.A(net189),
    .B(net188),
    .C(_0239_),
    .Y(_0272_));
 sg13g2_nor2_2 _0847_ (.A(_0271_),
    .B(_0272_),
    .Y(_0273_));
 sg13g2_or2_1 _0848_ (.X(_0274_),
    .B(_0272_),
    .A(_0271_));
 sg13g2_nor2b_1 _0849_ (.A(\pix_x[9] ),
    .B_N(\pix_x[8] ),
    .Y(_0275_));
 sg13g2_o21ai_1 _0850_ (.B1(_0275_),
    .Y(_0276_),
    .A1(_0271_),
    .A2(_0272_));
 sg13g2_nand4_1 _0851_ (.B(_0162_),
    .C(_0274_),
    .A(_0117_),
    .Y(_0277_),
    .D(_0275_));
 sg13g2_nand2_2 _0852_ (.Y(_0278_),
    .A(_0136_),
    .B(_0277_));
 sg13g2_a21o_1 _0853_ (.A2(net208),
    .A1(net207),
    .B1(net204),
    .X(_0279_));
 sg13g2_and2_2 _0854_ (.A(_0164_),
    .B(_0279_),
    .X(_0280_));
 sg13g2_and3_2 _0855_ (.X(_0281_),
    .A(_0203_),
    .B(_0274_),
    .C(_0280_));
 sg13g2_nand3_1 _0856_ (.B(_0274_),
    .C(_0280_),
    .A(_0203_),
    .Y(_0282_));
 sg13g2_nor2_1 _0857_ (.A(_0209_),
    .B(_0281_),
    .Y(_0283_));
 sg13g2_or2_1 _0858_ (.X(_0284_),
    .B(_0281_),
    .A(_0209_));
 sg13g2_nor2_1 _0859_ (.A(net202),
    .B(_0280_),
    .Y(_0285_));
 sg13g2_nor2_1 _0860_ (.A(_0160_),
    .B(_0273_),
    .Y(_0286_));
 sg13g2_nor3_2 _0861_ (.A(_0160_),
    .B(_0273_),
    .C(_0285_),
    .Y(_0287_));
 sg13g2_nor2_2 _0862_ (.A(_0185_),
    .B(_0287_),
    .Y(_0288_));
 sg13g2_or2_2 _0863_ (.X(_0289_),
    .B(_0287_),
    .A(_0185_));
 sg13g2_nand2_1 _0864_ (.Y(_0290_),
    .A(_0169_),
    .B(_0288_));
 sg13g2_nor2_1 _0865_ (.A(net208),
    .B(net210),
    .Y(_0291_));
 sg13g2_o21ai_1 _0866_ (.B1(net206),
    .Y(_0292_),
    .A1(net209),
    .A2(net210));
 sg13g2_nor3_1 _0867_ (.A(net206),
    .B(net208),
    .C(net210),
    .Y(_0293_));
 sg13g2_nand3b_1 _0868_ (.B(_0129_),
    .C(_0292_),
    .Y(_0294_),
    .A_N(_0293_));
 sg13g2_or2_2 _0869_ (.X(_0295_),
    .B(_0294_),
    .A(_0276_));
 sg13g2_o21ai_1 _0870_ (.B1(_0159_),
    .Y(_0296_),
    .A1(_0276_),
    .A2(_0294_));
 sg13g2_or2_1 _0871_ (.X(_0297_),
    .B(_0296_),
    .A(_0289_));
 sg13g2_nor4_2 _0872_ (.A(_0168_),
    .B(_0185_),
    .C(_0287_),
    .Y(_0298_),
    .D(_0296_));
 sg13g2_nor2b_1 _0873_ (.A(_0281_),
    .B_N(_0298_),
    .Y(_0299_));
 sg13g2_nand2_2 _0874_ (.Y(_0300_),
    .A(_0283_),
    .B(_0298_));
 sg13g2_o21ai_1 _0875_ (.B1(_0116_),
    .Y(_0301_),
    .A1(net209),
    .A2(_0112_));
 sg13g2_a21oi_1 _0876_ (.A1(net202),
    .A2(_0301_),
    .Y(_0302_),
    .B1(_0005_));
 sg13g2_nand3_1 _0877_ (.B(net209),
    .C(_0091_),
    .A(net202),
    .Y(_0303_));
 sg13g2_nor3_1 _0878_ (.A(_0112_),
    .B(_0206_),
    .C(_0303_),
    .Y(_0304_));
 sg13g2_nor2_1 _0879_ (.A(_0302_),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_nor4_2 _0880_ (.A(_0117_),
    .B(_0155_),
    .C(_0273_),
    .Y(_0306_),
    .D(_0305_));
 sg13g2_or4_2 _0881_ (.A(_0117_),
    .B(_0155_),
    .C(_0273_),
    .D(_0305_),
    .X(_0307_));
 sg13g2_nor2_2 _0882_ (.A(net177),
    .B(_0306_),
    .Y(_0308_));
 sg13g2_nand2b_1 _0883_ (.Y(_0309_),
    .B(_0307_),
    .A_N(net176));
 sg13g2_nor3_2 _0884_ (.A(_0278_),
    .B(_0300_),
    .C(_0309_),
    .Y(_0310_));
 sg13g2_nor3_2 _0885_ (.A(_0222_),
    .B(_0262_),
    .C(net169),
    .Y(_0311_));
 sg13g2_nand2_1 _0886_ (.Y(_0312_),
    .A(_0136_),
    .B(_0298_));
 sg13g2_a221oi_1 _0887_ (.B2(_0312_),
    .C1(net173),
    .B1(_0311_),
    .A1(net164),
    .Y(_0313_),
    .A2(_0310_));
 sg13g2_nand2_1 _0888_ (.Y(_0314_),
    .A(_0288_),
    .B(_0308_));
 sg13g2_and2_1 _0889_ (.A(_0170_),
    .B(_0288_),
    .X(_0315_));
 sg13g2_nand2_1 _0890_ (.Y(_0316_),
    .A(net179),
    .B(_0315_));
 sg13g2_nand3_1 _0891_ (.B(_0308_),
    .C(_0315_),
    .A(net179),
    .Y(_0317_));
 sg13g2_a221oi_1 _0892_ (.B2(net164),
    .C1(net171),
    .B1(_0317_),
    .A1(_0311_),
    .Y(_0318_),
    .A2(_0314_));
 sg13g2_o21ai_1 _0893_ (.B1(_0215_),
    .Y(_0319_),
    .A1(_0313_),
    .A2(_0318_));
 sg13g2_nand3_1 _0894_ (.B(_0144_),
    .C(net178),
    .A(_0138_),
    .Y(_0320_));
 sg13g2_nand2b_1 _0895_ (.Y(_0321_),
    .B(_0229_),
    .A_N(net178));
 sg13g2_nand3_1 _0896_ (.B(_0320_),
    .C(_0321_),
    .A(net179),
    .Y(_0322_));
 sg13g2_nor3_1 _0897_ (.A(_0200_),
    .B(net176),
    .C(_0251_),
    .Y(_0323_));
 sg13g2_a22oi_1 _0898_ (.Y(_0324_),
    .B1(_0322_),
    .B2(_0323_),
    .A2(net176),
    .A1(_0012_));
 sg13g2_or2_1 _0899_ (.X(_0325_),
    .B(_0324_),
    .A(_0209_));
 sg13g2_nand2_2 _0900_ (.Y(_0326_),
    .A(\pix_x[2] ),
    .B(_0325_));
 sg13g2_inv_1 _0901_ (.Y(_0327_),
    .A(_0326_));
 sg13g2_nor2_1 _0902_ (.A(net171),
    .B(net169),
    .Y(_0328_));
 sg13g2_nand2_2 _0903_ (.Y(_0329_),
    .A(net173),
    .B(net167));
 sg13g2_nor2_1 _0904_ (.A(_0290_),
    .B(_0329_),
    .Y(_0330_));
 sg13g2_nor2_1 _0905_ (.A(net171),
    .B(net168),
    .Y(_0331_));
 sg13g2_nand2_1 _0906_ (.Y(_0332_),
    .A(net173),
    .B(net169));
 sg13g2_and4_1 _0907_ (.A(_0169_),
    .B(_0288_),
    .C(_0295_),
    .D(_0307_),
    .X(_0333_));
 sg13g2_nor2_1 _0908_ (.A(_0278_),
    .B(_0332_),
    .Y(_0334_));
 sg13g2_a21oi_1 _0909_ (.A1(_0333_),
    .A2(_0334_),
    .Y(_0335_),
    .B1(_0330_));
 sg13g2_nand2b_2 _0910_ (.Y(_0336_),
    .B(_0307_),
    .A_N(_0209_));
 sg13g2_nand2_1 _0911_ (.Y(_0337_),
    .A(_0268_),
    .B(_0282_));
 sg13g2_nor3_1 _0912_ (.A(_0290_),
    .B(_0336_),
    .C(_0337_),
    .Y(_0338_));
 sg13g2_or3_1 _0913_ (.A(_0201_),
    .B(_0287_),
    .C(_0336_),
    .X(_0339_));
 sg13g2_nand2_1 _0914_ (.Y(_0340_),
    .A(_0169_),
    .B(_0277_));
 sg13g2_nor3_1 _0915_ (.A(net169),
    .B(_0339_),
    .C(_0340_),
    .Y(_0341_));
 sg13g2_o21ai_1 _0916_ (.B1(net170),
    .Y(_0342_),
    .A1(_0338_),
    .A2(_0341_));
 sg13g2_nand3_1 _0917_ (.B(_0335_),
    .C(_0342_),
    .A(_0263_),
    .Y(_0343_));
 sg13g2_a21oi_1 _0918_ (.A1(_0216_),
    .A2(_0343_),
    .Y(_0344_),
    .B1(_0326_));
 sg13g2_nor2b_1 _0919_ (.A(net177),
    .B_N(_0298_),
    .Y(_0345_));
 sg13g2_nand2_1 _0920_ (.Y(_0346_),
    .A(net179),
    .B(_0345_));
 sg13g2_nand2_1 _0921_ (.Y(_0347_),
    .A(_0277_),
    .B(_0282_));
 sg13g2_nor2_1 _0922_ (.A(_0346_),
    .B(_0347_),
    .Y(_0348_));
 sg13g2_o21ai_1 _0923_ (.B1(_0331_),
    .Y(_0349_),
    .A1(_0336_),
    .A2(_0348_));
 sg13g2_and4_1 _0924_ (.A(_0159_),
    .B(_0264_),
    .C(_0265_),
    .D(_0295_),
    .X(_0350_));
 sg13g2_a21oi_1 _0925_ (.A1(net167),
    .A2(_0299_),
    .Y(_0351_),
    .B1(_0350_));
 sg13g2_nor3_1 _0926_ (.A(net176),
    .B(net173),
    .C(_0351_),
    .Y(_0352_));
 sg13g2_nor3_1 _0927_ (.A(_0158_),
    .B(_0213_),
    .C(_0347_),
    .Y(_0353_));
 sg13g2_nor2_1 _0928_ (.A(_0135_),
    .B(_0329_),
    .Y(_0354_));
 sg13g2_a221oi_1 _0929_ (.B2(_0354_),
    .C1(net166),
    .B1(_0353_),
    .A1(net168),
    .Y(_0355_),
    .A2(_0306_));
 sg13g2_nor2b_1 _0930_ (.A(_0352_),
    .B_N(_0355_),
    .Y(_0356_));
 sg13g2_and2_1 _0931_ (.A(_0090_),
    .B(_0325_),
    .X(_0357_));
 sg13g2_nand2_1 _0932_ (.Y(_0358_),
    .A(_0090_),
    .B(_0325_));
 sg13g2_nand2_1 _0933_ (.Y(_0359_),
    .A(_0263_),
    .B(_0357_));
 sg13g2_o21ai_1 _0934_ (.B1(_0307_),
    .Y(_0360_),
    .A1(_0266_),
    .A2(_0267_));
 sg13g2_nor2_1 _0935_ (.A(_0284_),
    .B(_0297_),
    .Y(_0361_));
 sg13g2_nor2_1 _0936_ (.A(_0158_),
    .B(_0340_),
    .Y(_0362_));
 sg13g2_nand3_1 _0937_ (.B(_0170_),
    .C(_0277_),
    .A(net179),
    .Y(_0363_));
 sg13g2_nor3_1 _0938_ (.A(_0306_),
    .B(_0329_),
    .C(_0361_),
    .Y(_0364_));
 sg13g2_nor3_1 _0939_ (.A(_0309_),
    .B(_0332_),
    .C(_0363_),
    .Y(_0365_));
 sg13g2_a21o_1 _0940_ (.A2(net167),
    .A1(_0200_),
    .B1(net172),
    .X(_0366_));
 sg13g2_nor3_1 _0941_ (.A(net168),
    .B(_0284_),
    .C(_0317_),
    .Y(_0367_));
 sg13g2_a21oi_1 _0942_ (.A1(_0308_),
    .A2(_0362_),
    .Y(_0368_),
    .B1(_0268_));
 sg13g2_nor3_1 _0943_ (.A(_0366_),
    .B(_0367_),
    .C(_0368_),
    .Y(_0369_));
 sg13g2_or3_1 _0944_ (.A(_0364_),
    .B(_0365_),
    .C(_0369_),
    .X(_0370_));
 sg13g2_a221oi_1 _0945_ (.B2(net166),
    .C1(_0359_),
    .B1(_0370_),
    .A1(_0349_),
    .Y(_0371_),
    .A2(_0356_));
 sg13g2_a21o_1 _0946_ (.A2(_0344_),
    .A1(_0319_),
    .B1(_0371_),
    .X(_0372_));
 sg13g2_a221oi_1 _0947_ (.B2(_0314_),
    .C1(net170),
    .B1(_0311_),
    .A1(net164),
    .Y(_0373_),
    .A2(_0297_));
 sg13g2_a21oi_1 _0948_ (.A1(_0135_),
    .A2(net164),
    .Y(_0374_),
    .B1(net172));
 sg13g2_nand3_1 _0949_ (.B(_0295_),
    .C(_0308_),
    .A(_0283_),
    .Y(_0375_));
 sg13g2_nor4_1 _0950_ (.A(_0222_),
    .B(_0262_),
    .C(net169),
    .D(_0375_),
    .Y(_0376_));
 sg13g2_a221oi_1 _0951_ (.B2(_0376_),
    .C1(net172),
    .B1(_0277_),
    .A1(_0135_),
    .Y(_0377_),
    .A2(net164));
 sg13g2_nor4_1 _0952_ (.A(_0177_),
    .B(_0184_),
    .C(net172),
    .D(net169),
    .Y(_0378_));
 sg13g2_or4_1 _0953_ (.A(_0358_),
    .B(_0373_),
    .C(_0377_),
    .D(_0378_),
    .X(_0379_));
 sg13g2_a21oi_1 _0954_ (.A1(net164),
    .A2(_0310_),
    .Y(_0380_),
    .B1(net170));
 sg13g2_nor3_1 _0955_ (.A(_0284_),
    .B(_0289_),
    .C(_0363_),
    .Y(_0381_));
 sg13g2_nand4_1 _0956_ (.B(_0308_),
    .C(_0311_),
    .A(net173),
    .Y(_0382_),
    .D(_0381_));
 sg13g2_o21ai_1 _0957_ (.B1(_0382_),
    .Y(_0383_),
    .A1(_0374_),
    .A2(_0380_));
 sg13g2_a21oi_1 _0958_ (.A1(_0327_),
    .A2(_0383_),
    .Y(_0384_),
    .B1(_0216_));
 sg13g2_nor3_1 _0959_ (.A(_0213_),
    .B(_0289_),
    .C(_0363_),
    .Y(_0385_));
 sg13g2_a221oi_1 _0960_ (.B2(net164),
    .C1(net172),
    .B1(_0385_),
    .A1(_0310_),
    .Y(_0386_),
    .A2(_0311_));
 sg13g2_a21oi_2 _0961_ (.B1(net170),
    .Y(_0387_),
    .A2(_0311_),
    .A1(_0278_));
 sg13g2_nor4_2 _0962_ (.A(_0222_),
    .B(_0262_),
    .C(net167),
    .Y(_0388_),
    .D(_0375_));
 sg13g2_nand2_1 _0963_ (.Y(_0389_),
    .A(_0159_),
    .B(_0388_));
 sg13g2_nor4_1 _0964_ (.A(net168),
    .B(_0281_),
    .C(_0287_),
    .D(_0336_),
    .Y(_0390_));
 sg13g2_a21oi_1 _0965_ (.A1(net168),
    .A2(_0333_),
    .Y(_0391_),
    .B1(_0390_));
 sg13g2_nand2_1 _0966_ (.Y(_0392_),
    .A(net165),
    .B(_0391_));
 sg13g2_a221oi_1 _0967_ (.B2(net170),
    .C1(_0358_),
    .B1(_0392_),
    .A1(_0387_),
    .Y(_0393_),
    .A2(_0389_));
 sg13g2_nor3_1 _0968_ (.A(_0326_),
    .B(_0386_),
    .C(_0387_),
    .Y(_0394_));
 sg13g2_nor2_1 _0969_ (.A(_0393_),
    .B(_0394_),
    .Y(_0395_));
 sg13g2_a22oi_1 _0970_ (.Y(_0396_),
    .B1(_0395_),
    .B2(_0216_),
    .A2(_0384_),
    .A1(_0379_));
 sg13g2_nor2_1 _0971_ (.A(_0278_),
    .B(_0289_),
    .Y(_0397_));
 sg13g2_nor4_1 _0972_ (.A(net176),
    .B(_0222_),
    .C(_0262_),
    .D(net167),
    .Y(_0398_));
 sg13g2_o21ai_1 _0973_ (.B1(_0397_),
    .Y(_0399_),
    .A1(_0376_),
    .A2(_0398_));
 sg13g2_nand2b_1 _0974_ (.Y(_0400_),
    .B(net165),
    .A_N(net178));
 sg13g2_a22oi_1 _0975_ (.Y(_0401_),
    .B1(_0400_),
    .B2(_0387_),
    .A2(_0399_),
    .A1(net170));
 sg13g2_nor2_1 _0976_ (.A(net166),
    .B(_0401_),
    .Y(_0402_));
 sg13g2_nor2_1 _0977_ (.A(_0339_),
    .B(_0347_),
    .Y(_0403_));
 sg13g2_a221oi_1 _0978_ (.B2(_0311_),
    .C1(net170),
    .B1(_0403_),
    .A1(_0388_),
    .Y(_0404_),
    .A2(_0397_));
 sg13g2_nand3b_1 _0979_ (.B(net165),
    .C(net167),
    .Y(_0405_),
    .A_N(net178));
 sg13g2_a21oi_1 _0980_ (.A1(_0374_),
    .A2(_0405_),
    .Y(_0406_),
    .B1(_0404_));
 sg13g2_o21ai_1 _0981_ (.B1(_0357_),
    .Y(_0407_),
    .A1(_0216_),
    .A2(_0406_));
 sg13g2_nor3_1 _0982_ (.A(_0222_),
    .B(_0262_),
    .C(_0345_),
    .Y(_0408_));
 sg13g2_nor2_1 _0983_ (.A(_0332_),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_nand3_1 _0984_ (.B(_0282_),
    .C(_0288_),
    .A(net178),
    .Y(_0410_));
 sg13g2_nor2_1 _0985_ (.A(net177),
    .B(_0410_),
    .Y(_0411_));
 sg13g2_nor2_1 _0986_ (.A(_0306_),
    .B(_0411_),
    .Y(_0412_));
 sg13g2_a21oi_1 _0987_ (.A1(net165),
    .A2(_0412_),
    .Y(_0413_),
    .B1(_0329_));
 sg13g2_nor3_1 _0988_ (.A(_0377_),
    .B(_0409_),
    .C(_0413_),
    .Y(_0414_));
 sg13g2_nor2_1 _0989_ (.A(_0200_),
    .B(_0363_),
    .Y(_0415_));
 sg13g2_nor4_1 _0990_ (.A(_0222_),
    .B(_0262_),
    .C(net169),
    .D(_0415_),
    .Y(_0416_));
 sg13g2_o21ai_1 _0991_ (.B1(net172),
    .Y(_0417_),
    .A1(_0388_),
    .A2(_0416_));
 sg13g2_o21ai_1 _0992_ (.B1(net169),
    .Y(_0418_),
    .A1(_0336_),
    .A2(_0410_));
 sg13g2_nand2b_1 _0993_ (.Y(_0419_),
    .B(_0300_),
    .A_N(_0360_));
 sg13g2_a21oi_1 _0994_ (.A1(_0418_),
    .A2(_0419_),
    .Y(_0420_),
    .B1(net173));
 sg13g2_a21oi_1 _0995_ (.A1(net165),
    .A2(_0420_),
    .Y(_0421_),
    .B1(net166));
 sg13g2_a21oi_1 _0996_ (.A1(_0417_),
    .A2(_0421_),
    .Y(_0422_),
    .B1(_0326_));
 sg13g2_o21ai_1 _0997_ (.B1(_0422_),
    .Y(_0423_),
    .A1(_0216_),
    .A2(_0414_));
 sg13g2_o21ai_1 _0998_ (.B1(_0423_),
    .Y(_0424_),
    .A1(_0402_),
    .A2(_0407_));
 sg13g2_a221oi_1 _0999_ (.B2(_0346_),
    .C1(net173),
    .B1(_0311_),
    .A1(net164),
    .Y(_0425_),
    .A2(_0310_));
 sg13g2_a221oi_1 _1000_ (.B2(net165),
    .C1(net171),
    .B1(_0412_),
    .A1(_0135_),
    .Y(_0426_),
    .A2(_0270_));
 sg13g2_o21ai_1 _1001_ (.B1(_0215_),
    .Y(_0427_),
    .A1(_0425_),
    .A2(_0426_));
 sg13g2_or2_1 _1002_ (.X(_0428_),
    .B(_0381_),
    .A(_0360_));
 sg13g2_and2_1 _1003_ (.A(net171),
    .B(_0418_),
    .X(_0429_));
 sg13g2_o21ai_1 _1004_ (.B1(_0307_),
    .Y(_0430_),
    .A1(_0278_),
    .A2(_0300_));
 sg13g2_and2_1 _1005_ (.A(_0331_),
    .B(_0430_),
    .X(_0431_));
 sg13g2_a221oi_1 _1006_ (.B2(_0429_),
    .C1(_0431_),
    .B1(_0428_),
    .A1(_0315_),
    .Y(_0432_),
    .A2(_0328_));
 sg13g2_a21o_1 _1007_ (.A2(_0432_),
    .A1(net165),
    .B1(net166),
    .X(_0433_));
 sg13g2_nand3_1 _1008_ (.B(_0427_),
    .C(_0433_),
    .A(_0357_),
    .Y(_0434_));
 sg13g2_or2_1 _1009_ (.X(_0435_),
    .B(_0353_),
    .A(_0268_));
 sg13g2_o21ai_1 _1010_ (.B1(_0435_),
    .Y(_0436_),
    .A1(_0316_),
    .A2(_0337_));
 sg13g2_nor4_1 _1011_ (.A(_0213_),
    .B(net167),
    .C(_0281_),
    .D(_0363_),
    .Y(_0437_));
 sg13g2_a221oi_1 _1012_ (.B2(net173),
    .C1(_0306_),
    .B1(_0437_),
    .A1(_0297_),
    .Y(_0438_),
    .A2(_0328_));
 sg13g2_o21ai_1 _1013_ (.B1(_0438_),
    .Y(_0439_),
    .A1(_0366_),
    .A2(_0436_));
 sg13g2_nand2_1 _1014_ (.Y(_0440_),
    .A(net166),
    .B(_0439_));
 sg13g2_a21oi_1 _1015_ (.A1(net172),
    .A2(_0266_),
    .Y(_0441_),
    .B1(_0298_));
 sg13g2_a21oi_1 _1016_ (.A1(net172),
    .A2(_0278_),
    .Y(_0442_),
    .B1(_0441_));
 sg13g2_a221oi_1 _1017_ (.B2(_0307_),
    .C1(net166),
    .B1(_0442_),
    .A1(net170),
    .Y(_0443_),
    .A2(_0350_));
 sg13g2_nand3_1 _1018_ (.B(_0327_),
    .C(_0440_),
    .A(net165),
    .Y(_0444_));
 sg13g2_o21ai_1 _1019_ (.B1(_0434_),
    .Y(_0445_),
    .A1(_0443_),
    .A2(_0444_));
 sg13g2_mux4_1 _1020_ (.S0(net210),
    .A0(_0424_),
    .A1(_0445_),
    .A2(_0372_),
    .A3(_0396_),
    .S1(net208),
    .X(_0446_));
 sg13g2_nand4_1 _1021_ (.B(_0111_),
    .C(_0135_),
    .A(\driver.decoder.data_reg[2] ),
    .Y(_0447_),
    .D(_0446_));
 sg13g2_mux4_1 _1022_ (.S0(net210),
    .A0(_0372_),
    .A1(_0396_),
    .A2(_0424_),
    .A3(_0445_),
    .S1(net208),
    .X(_0448_));
 sg13g2_nand2_1 _1023_ (.Y(_0449_),
    .A(_0281_),
    .B(_0448_));
 sg13g2_nand3_1 _1024_ (.B(_0281_),
    .C(_0448_),
    .A(net213),
    .Y(_0450_));
 sg13g2_nand4_1 _1025_ (.B(_0111_),
    .C(_0185_),
    .A(\driver.decoder.data_reg[11] ),
    .Y(_0451_),
    .D(_0446_));
 sg13g2_and3_1 _1026_ (.X(_0452_),
    .A(_0447_),
    .B(_0450_),
    .C(_0451_));
 sg13g2_nor2b_1 _1027_ (.A(_0165_),
    .B_N(_0448_),
    .Y(_0453_));
 sg13g2_nand2_1 _1028_ (.Y(_0454_),
    .A(\driver.decoder.data_reg[0] ),
    .B(_0168_));
 sg13g2_o21ai_1 _1029_ (.B1(_0454_),
    .Y(_0455_),
    .A1(_0104_),
    .A2(_0277_));
 sg13g2_mux4_1 _1030_ (.S0(net210),
    .A0(_0396_),
    .A1(_0424_),
    .A2(_0445_),
    .A3(_0372_),
    .S1(net208),
    .X(_0456_));
 sg13g2_o21ai_1 _1031_ (.B1(net210),
    .Y(_0457_),
    .A1(_0206_),
    .A2(_0275_));
 sg13g2_and2_1 _1032_ (.A(_0164_),
    .B(_0457_),
    .X(_0458_));
 sg13g2_xnor2_1 _1033_ (.Y(_0459_),
    .A(_0007_),
    .B(_0291_));
 sg13g2_or2_1 _1034_ (.X(_0460_),
    .B(_0459_),
    .A(_0163_));
 sg13g2_nor3_1 _1035_ (.A(_0091_),
    .B(_0161_),
    .C(_0206_),
    .Y(_0461_));
 sg13g2_nor4_2 _1036_ (.A(_0276_),
    .B(_0458_),
    .C(_0460_),
    .Y(_0462_),
    .D(_0461_));
 sg13g2_and3_1 _1037_ (.X(_0463_),
    .A(net102),
    .B(_0456_),
    .C(_0462_));
 sg13g2_xnor2_1 _1038_ (.Y(_0464_),
    .A(_0002_),
    .B(_0293_));
 sg13g2_nor3_1 _1039_ (.A(_0295_),
    .B(_0459_),
    .C(_0464_),
    .Y(_0465_));
 sg13g2_and2_1 _1040_ (.A(_0456_),
    .B(_0465_),
    .X(_0466_));
 sg13g2_a221oi_1 _1041_ (.B2(net120),
    .C1(_0463_),
    .B1(_0466_),
    .A1(_0453_),
    .Y(_0467_),
    .A2(_0455_));
 sg13g2_and2_1 _1042_ (.A(_0204_),
    .B(_0446_),
    .X(_0468_));
 sg13g2_a22oi_1 _1043_ (.Y(_0469_),
    .B1(net177),
    .B2(\driver.decoder.data_reg[6] ),
    .A2(_0209_),
    .A1(\driver.decoder.data_reg[7] ));
 sg13g2_inv_1 _1044_ (.Y(_0470_),
    .A(_0469_));
 sg13g2_and4_1 _1045_ (.A(_0002_),
    .B(_0162_),
    .C(_0306_),
    .D(_0448_),
    .X(_0471_));
 sg13g2_a22oi_1 _1046_ (.Y(_0472_),
    .B1(_0471_),
    .B2(net108),
    .A2(_0470_),
    .A1(_0468_));
 sg13g2_nor2_1 _1047_ (.A(net205),
    .B(_0007_),
    .Y(_0473_));
 sg13g2_nand3_1 _1048_ (.B(_0446_),
    .C(_0473_),
    .A(_0158_),
    .Y(_0474_));
 sg13g2_nand4_1 _1049_ (.B(_0158_),
    .C(_0446_),
    .A(\driver.decoder.data_reg[1] ),
    .Y(_0475_),
    .D(_0473_));
 sg13g2_nand3_1 _1050_ (.B(_0286_),
    .C(_0448_),
    .A(_0280_),
    .Y(_0476_));
 sg13g2_nand4_1 _1051_ (.B(_0280_),
    .C(_0286_),
    .A(\driver.decoder.data_reg[3] ),
    .Y(_0477_),
    .D(_0448_));
 sg13g2_and2_1 _1052_ (.A(_0475_),
    .B(_0477_),
    .X(_0478_));
 sg13g2_nand4_1 _1053_ (.B(_0467_),
    .C(_0472_),
    .A(_0452_),
    .Y(_0479_),
    .D(_0478_));
 sg13g2_and3_1 _1054_ (.X(_0480_),
    .A(_0449_),
    .B(_0474_),
    .C(_0476_));
 sg13g2_nand3_1 _1055_ (.B(_0474_),
    .C(_0476_),
    .A(_0449_),
    .Y(_0481_));
 sg13g2_nand3_1 _1056_ (.B(_0201_),
    .C(_0446_),
    .A(_0111_),
    .Y(_0482_));
 sg13g2_o21ai_1 _1057_ (.B1(_0456_),
    .Y(_0483_),
    .A1(_0462_),
    .A2(_0465_));
 sg13g2_nand3b_1 _1058_ (.B(_0482_),
    .C(_0483_),
    .Y(_0484_),
    .A_N(_0471_));
 sg13g2_and3_1 _1059_ (.X(_0485_),
    .A(_0204_),
    .B(_0213_),
    .C(_0446_));
 sg13g2_a21o_1 _1060_ (.A2(_0453_),
    .A1(_0340_),
    .B1(_0485_),
    .X(_0486_));
 sg13g2_nor2_1 _1061_ (.A(_0484_),
    .B(_0486_),
    .Y(_0487_));
 sg13g2_nor3_1 _1062_ (.A(_0481_),
    .B(_0484_),
    .C(_0486_),
    .Y(_0488_));
 sg13g2_nor4_1 _1063_ (.A(net188),
    .B(_0089_),
    .C(_0109_),
    .D(_0113_),
    .Y(_0489_));
 sg13g2_o21ai_1 _1064_ (.B1(_0489_),
    .Y(_0490_),
    .A1(_0085_),
    .A2(_0105_));
 sg13g2_a221oi_1 _1065_ (.B2(_0487_),
    .C1(_0490_),
    .B1(_0480_),
    .A1(_0124_),
    .Y(_0018_),
    .A2(_0479_));
 sg13g2_nor2b_1 _1066_ (.A(\driver.driver.pmod_latch_prev ),
    .B_N(net77),
    .Y(_0491_));
 sg13g2_nor2b_1 _1067_ (.A(net187),
    .B_N(net212),
    .Y(_0492_));
 sg13g2_a22oi_1 _1068_ (.Y(_0019_),
    .B1(net183),
    .B2(_0094_),
    .A2(net187),
    .A1(_0081_));
 sg13g2_a22oi_1 _1069_ (.Y(_0020_),
    .B1(net183),
    .B2(_0093_),
    .A2(net187),
    .A1(_0080_));
 sg13g2_a22oi_1 _1070_ (.Y(_0021_),
    .B1(net182),
    .B2(_0096_),
    .A2(net186),
    .A1(_0079_));
 sg13g2_a22oi_1 _1071_ (.Y(_0022_),
    .B1(net182),
    .B2(_0095_),
    .A2(net186),
    .A1(_0078_));
 sg13g2_a22oi_1 _1072_ (.Y(_0023_),
    .B1(net182),
    .B2(_0098_),
    .A2(net186),
    .A1(_0077_));
 sg13g2_a22oi_1 _1073_ (.Y(_0024_),
    .B1(net182),
    .B2(_0097_),
    .A2(net186),
    .A1(_0076_));
 sg13g2_a22oi_1 _1074_ (.Y(_0025_),
    .B1(net182),
    .B2(_0100_),
    .A2(net186),
    .A1(_0075_));
 sg13g2_a22oi_1 _1075_ (.Y(_0026_),
    .B1(net182),
    .B2(_0099_),
    .A2(net186),
    .A1(_0074_));
 sg13g2_a22oi_1 _1076_ (.Y(_0027_),
    .B1(net182),
    .B2(_0102_),
    .A2(net186),
    .A1(_0073_));
 sg13g2_a22oi_1 _1077_ (.Y(_0028_),
    .B1(net182),
    .B2(_0101_),
    .A2(net186),
    .A1(_0072_));
 sg13g2_a22oi_1 _1078_ (.Y(_0029_),
    .B1(net183),
    .B2(_0104_),
    .A2(net187),
    .A1(_0071_));
 sg13g2_a22oi_1 _1079_ (.Y(_0030_),
    .B1(net183),
    .B2(_0103_),
    .A2(net187),
    .A1(_0084_));
 sg13g2_nand2_2 _1080_ (.Y(_0493_),
    .A(net157),
    .B(net149));
 sg13g2_nor3_2 _1081_ (.A(_0090_),
    .B(_0091_),
    .C(_0493_),
    .Y(_0494_));
 sg13g2_nand4_1 _1082_ (.B(_0109_),
    .C(_0130_),
    .A(net209),
    .Y(_0495_),
    .D(_0494_));
 sg13g2_and2_1 _1083_ (.A(net211),
    .B(_0495_),
    .X(_0496_));
 sg13g2_nand2_2 _1084_ (.Y(_0497_),
    .A(net211),
    .B(_0495_));
 sg13g2_and2_1 _1085_ (.A(net79),
    .B(net175),
    .X(_0031_));
 sg13g2_and3_1 _1086_ (.X(_0032_),
    .A(net150),
    .B(_0493_),
    .C(net175));
 sg13g2_xnor2_1 _1087_ (.Y(_0498_),
    .A(_0090_),
    .B(_0493_));
 sg13g2_nor2_1 _1088_ (.A(_0497_),
    .B(net158),
    .Y(_0033_));
 sg13g2_nor2_1 _1089_ (.A(net95),
    .B(_0493_),
    .Y(_0499_));
 sg13g2_xnor2_1 _1090_ (.Y(_0500_),
    .A(\pix_x[3] ),
    .B(net96));
 sg13g2_nor2_1 _1091_ (.A(_0497_),
    .B(net97),
    .Y(_0034_));
 sg13g2_xor2_1 _1092_ (.B(_0494_),
    .A(net87),
    .X(_0501_));
 sg13g2_nor2_1 _1093_ (.A(_0497_),
    .B(net88),
    .Y(_0035_));
 sg13g2_nand2b_1 _1094_ (.Y(_0502_),
    .B(_0494_),
    .A_N(_0116_));
 sg13g2_inv_1 _1095_ (.Y(_0503_),
    .A(_0502_));
 sg13g2_a21oi_1 _1096_ (.A1(net209),
    .A2(_0494_),
    .Y(_0504_),
    .B1(net206));
 sg13g2_nor3_1 _1097_ (.A(_0497_),
    .B(_0503_),
    .C(net216),
    .Y(_0036_));
 sg13g2_xor2_1 _1098_ (.B(_0502_),
    .A(net204),
    .X(_0505_));
 sg13g2_nor2_1 _1099_ (.A(_0497_),
    .B(_0505_),
    .Y(_0037_));
 sg13g2_nor2_1 _1100_ (.A(_0002_),
    .B(_0502_),
    .Y(_0506_));
 sg13g2_o21ai_1 _1101_ (.B1(net175),
    .Y(_0507_),
    .A1(net203),
    .A2(_0506_));
 sg13g2_a21oi_1 _1102_ (.A1(net203),
    .A2(_0506_),
    .Y(_0038_),
    .B1(_0507_));
 sg13g2_nor2b_1 _1103_ (.A(_0118_),
    .B_N(_0494_),
    .Y(_0508_));
 sg13g2_xnor2_1 _1104_ (.Y(_0509_),
    .A(net163),
    .B(_0508_));
 sg13g2_nor2_1 _1105_ (.A(_0497_),
    .B(_0509_),
    .Y(_0039_));
 sg13g2_a21oi_1 _1106_ (.A1(\pix_x[8] ),
    .A2(_0508_),
    .Y(_0510_),
    .B1(net145));
 sg13g2_a21oi_1 _1107_ (.A1(_0109_),
    .A2(_0508_),
    .Y(_0511_),
    .B1(_0497_));
 sg13g2_nor2b_1 _1108_ (.A(net146),
    .B_N(_0511_),
    .Y(_0040_));
 sg13g2_nor3_1 _1109_ (.A(_0123_),
    .B(_0488_),
    .C(_0490_),
    .Y(_0042_));
 sg13g2_nor4_1 _1110_ (.A(_0123_),
    .B(net214),
    .C(_0488_),
    .D(_0490_),
    .Y(_0041_));
 sg13g2_and2_1 _1111_ (.A(net212),
    .B(net1),
    .X(_0043_));
 sg13g2_and2_1 _1112_ (.A(net212),
    .B(net86),
    .X(_0044_));
 sg13g2_nand2_1 _1113_ (.Y(_0512_),
    .A(\pix_y[0] ),
    .B(net175));
 sg13g2_nand3b_1 _1114_ (.B(net188),
    .C(_0179_),
    .Y(_0513_),
    .A_N(net190));
 sg13g2_nand4_1 _1115_ (.B(net198),
    .C(_0143_),
    .A(net200),
    .Y(_0514_),
    .D(_0148_));
 sg13g2_o21ai_1 _1116_ (.B1(net211),
    .Y(_0515_),
    .A1(_0513_),
    .A2(_0514_));
 sg13g2_or2_2 _1117_ (.X(_0516_),
    .B(_0515_),
    .A(_0495_));
 sg13g2_o21ai_1 _1118_ (.B1(_0512_),
    .Y(_0045_),
    .A1(_0083_),
    .A2(_0516_));
 sg13g2_nand2_1 _1119_ (.Y(_0517_),
    .A(net134),
    .B(net174));
 sg13g2_nand2_1 _1120_ (.Y(_0518_),
    .A(net134),
    .B(\pix_y[0] ));
 sg13g2_nand2_1 _1121_ (.Y(_0519_),
    .A(_0180_),
    .B(_0518_));
 sg13g2_o21ai_1 _1122_ (.B1(_0517_),
    .Y(_0046_),
    .A1(_0516_),
    .A2(_0519_));
 sg13g2_nor2_1 _1123_ (.A(net174),
    .B(_0518_),
    .Y(_0520_));
 sg13g2_and2_2 _1124_ (.A(_0497_),
    .B(_0515_),
    .X(_0521_));
 sg13g2_xnor2_1 _1125_ (.Y(_0522_),
    .A(net200),
    .B(_0520_));
 sg13g2_nor2_1 _1126_ (.A(_0521_),
    .B(net221),
    .Y(_0047_));
 sg13g2_nand2_1 _1127_ (.Y(_0523_),
    .A(net198),
    .B(net175));
 sg13g2_nor2_1 _1128_ (.A(net152),
    .B(_0518_),
    .Y(_0524_));
 sg13g2_xnor2_1 _1129_ (.Y(_0525_),
    .A(net198),
    .B(net153));
 sg13g2_o21ai_1 _1130_ (.B1(_0523_),
    .Y(_0048_),
    .A1(_0516_),
    .A2(_0525_));
 sg13g2_or2_2 _1131_ (.X(_0526_),
    .B(_0518_),
    .A(_0137_));
 sg13g2_nor2_1 _1132_ (.A(net174),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_nor2_1 _1133_ (.A(net197),
    .B(_0527_),
    .Y(_0528_));
 sg13g2_nor3_1 _1134_ (.A(_0087_),
    .B(net174),
    .C(_0526_),
    .Y(_0529_));
 sg13g2_nor3_1 _1135_ (.A(_0521_),
    .B(_0528_),
    .C(_0529_),
    .Y(_0049_));
 sg13g2_nand2_1 _1136_ (.Y(_0530_),
    .A(net196),
    .B(net174));
 sg13g2_nor2_1 _1137_ (.A(net154),
    .B(_0526_),
    .Y(_0531_));
 sg13g2_xnor2_1 _1138_ (.Y(_0532_),
    .A(net196),
    .B(_0531_));
 sg13g2_o21ai_1 _1139_ (.B1(_0530_),
    .Y(_0050_),
    .A1(_0516_),
    .A2(net155));
 sg13g2_nor3_1 _1140_ (.A(_0139_),
    .B(net174),
    .C(_0526_),
    .Y(_0533_));
 sg13g2_a21oi_1 _1141_ (.A1(net196),
    .A2(_0529_),
    .Y(_0534_),
    .B1(net194));
 sg13g2_nor3_1 _1142_ (.A(_0521_),
    .B(_0533_),
    .C(net160),
    .Y(_0051_));
 sg13g2_nand2_1 _1143_ (.Y(_0535_),
    .A(net192),
    .B(net174));
 sg13g2_nor3_1 _1144_ (.A(_0010_),
    .B(_0138_),
    .C(_0526_),
    .Y(_0536_));
 sg13g2_xnor2_1 _1145_ (.Y(_0537_),
    .A(net192),
    .B(_0536_));
 sg13g2_o21ai_1 _1146_ (.B1(_0535_),
    .Y(_0052_),
    .A1(_0516_),
    .A2(_0537_));
 sg13g2_nand2_1 _1147_ (.Y(_0538_),
    .A(net192),
    .B(_0533_));
 sg13g2_xor2_1 _1148_ (.B(_0538_),
    .A(net189),
    .X(_0539_));
 sg13g2_nor2_1 _1149_ (.A(_0521_),
    .B(_0539_),
    .Y(_0053_));
 sg13g2_nand2_1 _1150_ (.Y(_0540_),
    .A(net188),
    .B(net174));
 sg13g2_nor3_1 _1151_ (.A(_0009_),
    .B(_0239_),
    .C(_0526_),
    .Y(_0541_));
 sg13g2_xnor2_1 _1152_ (.Y(_0542_),
    .A(net188),
    .B(_0541_));
 sg13g2_o21ai_1 _1153_ (.B1(_0540_),
    .Y(_0054_),
    .A1(_0516_),
    .A2(_0542_));
 sg13g2_nor2b_1 _1154_ (.A(\driver.driver.pmod_clk_prev ),
    .B_N(net78),
    .Y(_0543_));
 sg13g2_nor2b_1 _1155_ (.A(net185),
    .B_N(net212),
    .Y(_0544_));
 sg13g2_a22oi_1 _1156_ (.Y(_0055_),
    .B1(net181),
    .B2(_0081_),
    .A2(net185),
    .A1(_0082_));
 sg13g2_a22oi_1 _1157_ (.Y(_0056_),
    .B1(net181),
    .B2(_0080_),
    .A2(net185),
    .A1(_0081_));
 sg13g2_a22oi_1 _1158_ (.Y(_0057_),
    .B1(net181),
    .B2(_0079_),
    .A2(net185),
    .A1(_0080_));
 sg13g2_a22oi_1 _1159_ (.Y(_0058_),
    .B1(net180),
    .B2(_0078_),
    .A2(net184),
    .A1(_0079_));
 sg13g2_a22oi_1 _1160_ (.Y(_0059_),
    .B1(net180),
    .B2(_0077_),
    .A2(net184),
    .A1(_0078_));
 sg13g2_a22oi_1 _1161_ (.Y(_0060_),
    .B1(net180),
    .B2(_0076_),
    .A2(net184),
    .A1(_0077_));
 sg13g2_a22oi_1 _1162_ (.Y(_0061_),
    .B1(net180),
    .B2(_0075_),
    .A2(net184),
    .A1(_0076_));
 sg13g2_a22oi_1 _1163_ (.Y(_0062_),
    .B1(net180),
    .B2(_0074_),
    .A2(net184),
    .A1(_0075_));
 sg13g2_a22oi_1 _1164_ (.Y(_0063_),
    .B1(net180),
    .B2(_0073_),
    .A2(net184),
    .A1(_0074_));
 sg13g2_a22oi_1 _1165_ (.Y(_0064_),
    .B1(net180),
    .B2(_0072_),
    .A2(net184),
    .A1(_0073_));
 sg13g2_a22oi_1 _1166_ (.Y(_0065_),
    .B1(net180),
    .B2(_0071_),
    .A2(net184),
    .A1(_0072_));
 sg13g2_a22oi_1 _1167_ (.Y(_0066_),
    .B1(net181),
    .B2(_0084_),
    .A2(net185),
    .A1(_0071_));
 sg13g2_and2_1 _1168_ (.A(net211),
    .B(net3),
    .X(_0067_));
 sg13g2_and2_1 _1169_ (.A(net211),
    .B(net82),
    .X(_0068_));
 sg13g2_and2_1 _1170_ (.A(net211),
    .B(net2),
    .X(_0069_));
 sg13g2_and2_1 _1171_ (.A(net211),
    .B(net83),
    .X(_0070_));
 sg13g2_dfrbp_1 _1172_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net47),
    .D(_0018_),
    .Q_N(_0582_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _1173_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net63),
    .D(net105),
    .Q_N(_0581_),
    .Q(\driver.decoder.data_reg[0] ));
 sg13g2_dfrbp_1 _1174_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net61),
    .D(net117),
    .Q_N(_0580_),
    .Q(\driver.decoder.data_reg[1] ));
 sg13g2_dfrbp_1 _1175_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net56),
    .D(net119),
    .Q_N(_0579_),
    .Q(\driver.decoder.data_reg[2] ));
 sg13g2_dfrbp_1 _1176_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net54),
    .D(net107),
    .Q_N(_0578_),
    .Q(\driver.decoder.data_reg[3] ));
 sg13g2_dfrbp_1 _1177_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net52),
    .D(net109),
    .Q_N(_0577_),
    .Q(\driver.decoder.data_reg[4] ));
 sg13g2_dfrbp_1 _1178_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net50),
    .D(net99),
    .Q_N(_0576_),
    .Q(\driver.decoder.data_reg[5] ));
 sg13g2_dfrbp_1 _1179_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net48),
    .D(net90),
    .Q_N(_0575_),
    .Q(\driver.decoder.data_reg[6] ));
 sg13g2_dfrbp_1 _1180_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net45),
    .D(net101),
    .Q_N(_0574_),
    .Q(\driver.decoder.data_reg[7] ));
 sg13g2_dfrbp_1 _1181_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net43),
    .D(net103),
    .Q_N(_0573_),
    .Q(\driver.decoder.data_reg[8] ));
 sg13g2_dfrbp_1 _1182_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net41),
    .D(net121),
    .Q_N(_0572_),
    .Q(\driver.decoder.data_reg[9] ));
 sg13g2_dfrbp_1 _1183_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net39),
    .D(net137),
    .Q_N(_0571_),
    .Q(\driver.decoder.data_reg[10] ));
 sg13g2_dfrbp_1 _1184_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net37),
    .D(net123),
    .Q_N(_0570_),
    .Q(\driver.decoder.data_reg[11] ));
 sg13g2_dfrbp_1 _1185_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net35),
    .D(_0031_),
    .Q_N(_0017_),
    .Q(\pix_x[0] ));
 sg13g2_dfrbp_1 _1186_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net34),
    .D(net151),
    .Q_N(_0569_),
    .Q(\pix_x[1] ));
 sg13g2_dfrbp_1 _1187_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net33),
    .D(_0033_),
    .Q_N(_0004_),
    .Q(\pix_x[2] ));
 sg13g2_dfrbp_1 _1188_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net32),
    .D(_0034_),
    .Q_N(_0568_),
    .Q(\pix_x[3] ));
 sg13g2_dfrbp_1 _1189_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net31),
    .D(_0035_),
    .Q_N(_0003_),
    .Q(\pix_x[4] ));
 sg13g2_dfrbp_1 _1190_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net30),
    .D(_0036_),
    .Q_N(_0007_),
    .Q(\pix_x[5] ));
 sg13g2_dfrbp_1 _1191_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net29),
    .D(_0037_),
    .Q_N(_0002_),
    .Q(\pix_x[6] ));
 sg13g2_dfrbp_1 _1192_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net28),
    .D(net148),
    .Q_N(_0005_),
    .Q(\pix_x[7] ));
 sg13g2_dfrbp_1 _1193_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net27),
    .D(_0039_),
    .Q_N(_0567_),
    .Q(\pix_x[8] ));
 sg13g2_dfrbp_1 _1194_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net26),
    .D(_0040_),
    .Q_N(_0006_),
    .Q(\pix_x[9] ));
 sg13g2_dfrbp_1 _1195_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net25),
    .D(_0041_),
    .Q_N(_0566_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _1196_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net24),
    .D(_0042_),
    .Q_N(_0565_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _1197_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net23),
    .D(_0043_),
    .Q_N(_0564_),
    .Q(\driver.driver.pmod_latch_sync[0] ));
 sg13g2_dfrbp_1 _1198_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net58),
    .D(_0044_),
    .Q_N(_0583_),
    .Q(\driver.driver.pmod_latch_sync[1] ));
 sg13g2_dfrbp_1 _1199_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net22),
    .D(net81),
    .Q_N(_0563_),
    .Q(hsync));
 sg13g2_dfrbp_1 _1200_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net21),
    .D(net85),
    .Q_N(_0016_),
    .Q(\pix_y[0] ));
 sg13g2_dfrbp_1 _1201_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net76),
    .D(net135),
    .Q_N(_0562_),
    .Q(\pix_y[1] ));
 sg13g2_dfrbp_1 _1202_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net74),
    .D(_0047_),
    .Q_N(_0013_),
    .Q(\pix_y[2] ));
 sg13g2_dfrbp_1 _1203_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net72),
    .D(_0048_),
    .Q_N(_0014_),
    .Q(\pix_y[3] ));
 sg13g2_dfrbp_1 _1204_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net70),
    .D(_0049_),
    .Q_N(_0015_),
    .Q(\pix_y[4] ));
 sg13g2_dfrbp_1 _1205_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net68),
    .D(net156),
    .Q_N(_0012_),
    .Q(\pix_y[5] ));
 sg13g2_dfrbp_1 _1206_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net66),
    .D(_0051_),
    .Q_N(_0010_),
    .Q(\pix_y[6] ));
 sg13g2_dfrbp_1 _1207_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net64),
    .D(net219),
    .Q_N(_0011_),
    .Q(\pix_y[7] ));
 sg13g2_dfrbp_1 _1208_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net57),
    .D(_0053_),
    .Q_N(_0009_),
    .Q(\pix_y[8] ));
 sg13g2_dfrbp_1 _1209_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net59),
    .D(net162),
    .Q_N(_0008_),
    .Q(\pix_y[9] ));
 sg13g2_dfrbp_1 _1210_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net60),
    .D(net144),
    .Q_N(_0584_),
    .Q(\vga_sync_gen.vsync ));
 sg13g2_dfrbp_1 _1211_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net65),
    .D(net78),
    .Q_N(_0585_),
    .Q(\driver.driver.pmod_clk_prev ));
 sg13g2_dfrbp_1 _1212_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net53),
    .D(net77),
    .Q_N(_0561_),
    .Q(\driver.driver.pmod_latch_prev ));
 sg13g2_dfrbp_1 _1213_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net49),
    .D(net94),
    .Q_N(_0560_),
    .Q(\driver.driver.shift_reg[0] ));
 sg13g2_dfrbp_1 _1214_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net44),
    .D(net115),
    .Q_N(_0559_),
    .Q(\driver.driver.shift_reg[1] ));
 sg13g2_dfrbp_1 _1215_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net40),
    .D(net141),
    .Q_N(_0558_),
    .Q(\driver.driver.shift_reg[2] ));
 sg13g2_dfrbp_1 _1216_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net36),
    .D(net129),
    .Q_N(_0557_),
    .Q(\driver.driver.shift_reg[3] ));
 sg13g2_dfrbp_1 _1217_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net75),
    .D(net125),
    .Q_N(_0556_),
    .Q(\driver.driver.shift_reg[4] ));
 sg13g2_dfrbp_1 _1218_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net71),
    .D(net139),
    .Q_N(_0555_),
    .Q(\driver.driver.shift_reg[5] ));
 sg13g2_dfrbp_1 _1219_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net67),
    .D(net113),
    .Q_N(_0554_),
    .Q(\driver.driver.shift_reg[6] ));
 sg13g2_dfrbp_1 _1220_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net62),
    .D(net111),
    .Q_N(_0553_),
    .Q(\driver.driver.shift_reg[7] ));
 sg13g2_dfrbp_1 _1221_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net51),
    .D(net131),
    .Q_N(_0552_),
    .Q(\driver.driver.shift_reg[8] ));
 sg13g2_dfrbp_1 _1222_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net42),
    .D(net127),
    .Q_N(_0551_),
    .Q(\driver.driver.shift_reg[9] ));
 sg13g2_dfrbp_1 _1223_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net20),
    .D(net133),
    .Q_N(_0550_),
    .Q(\driver.driver.shift_reg[10] ));
 sg13g2_dfrbp_1 _1224_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net69),
    .D(net92),
    .Q_N(_0549_),
    .Q(\driver.driver.shift_reg[11] ));
 sg13g2_dfrbp_1 _1225_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net55),
    .D(_0067_),
    .Q_N(_0548_),
    .Q(\driver.driver.pmod_data_sync[0] ));
 sg13g2_dfrbp_1 _1226_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net46),
    .D(_0068_),
    .Q_N(_0547_),
    .Q(\driver.driver.pmod_data_sync[1] ));
 sg13g2_dfrbp_1 _1227_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net38),
    .D(_0069_),
    .Q_N(_0546_),
    .Q(\driver.driver.pmod_clk_sync[0] ));
 sg13g2_dfrbp_1 _1228_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net73),
    .D(_0070_),
    .Q_N(_0545_),
    .Q(\driver.driver.pmod_clk_sync[1] ));
 sg13g2_tiehi _1200__21 (.L_HI(net21));
 sg13g2_tiehi _1199__22 (.L_HI(net22));
 sg13g2_tiehi _1197__23 (.L_HI(net23));
 sg13g2_tiehi _1196__24 (.L_HI(net24));
 sg13g2_tiehi _1195__25 (.L_HI(net25));
 sg13g2_tiehi _1194__26 (.L_HI(net26));
 sg13g2_tiehi _1193__27 (.L_HI(net27));
 sg13g2_tiehi _1192__28 (.L_HI(net28));
 sg13g2_tiehi _1191__29 (.L_HI(net29));
 sg13g2_tiehi _1190__30 (.L_HI(net30));
 sg13g2_tiehi _1189__31 (.L_HI(net31));
 sg13g2_tiehi _1188__32 (.L_HI(net32));
 sg13g2_tiehi _1187__33 (.L_HI(net33));
 sg13g2_tiehi _1186__34 (.L_HI(net34));
 sg13g2_tiehi _1185__35 (.L_HI(net35));
 sg13g2_tiehi _1216__36 (.L_HI(net36));
 sg13g2_tiehi _1184__37 (.L_HI(net37));
 sg13g2_tiehi _1227__38 (.L_HI(net38));
 sg13g2_tiehi _1183__39 (.L_HI(net39));
 sg13g2_tiehi _1215__40 (.L_HI(net40));
 sg13g2_tiehi _1182__41 (.L_HI(net41));
 sg13g2_tiehi _1222__42 (.L_HI(net42));
 sg13g2_tiehi _1181__43 (.L_HI(net43));
 sg13g2_tiehi _1214__44 (.L_HI(net44));
 sg13g2_tiehi _1180__45 (.L_HI(net45));
 sg13g2_tiehi _1226__46 (.L_HI(net46));
 sg13g2_tiehi _1172__47 (.L_HI(net47));
 sg13g2_tiehi _1179__48 (.L_HI(net48));
 sg13g2_tiehi _1213__49 (.L_HI(net49));
 sg13g2_tiehi _1178__50 (.L_HI(net50));
 sg13g2_tiehi _1221__51 (.L_HI(net51));
 sg13g2_tiehi _1177__52 (.L_HI(net52));
 sg13g2_tiehi _1212__53 (.L_HI(net53));
 sg13g2_tiehi _1176__54 (.L_HI(net54));
 sg13g2_tiehi _1225__55 (.L_HI(net55));
 sg13g2_tiehi _1175__56 (.L_HI(net56));
 sg13g2_tiehi _1208__57 (.L_HI(net57));
 sg13g2_tiehi _1198__58 (.L_HI(net58));
 sg13g2_tiehi _1209__59 (.L_HI(net59));
 sg13g2_tiehi _1210__60 (.L_HI(net60));
 sg13g2_tiehi _1174__61 (.L_HI(net61));
 sg13g2_tiehi _1220__62 (.L_HI(net62));
 sg13g2_tiehi _1173__63 (.L_HI(net63));
 sg13g2_tiehi _1207__64 (.L_HI(net64));
 sg13g2_tiehi _1211__65 (.L_HI(net65));
 sg13g2_tiehi _1206__66 (.L_HI(net66));
 sg13g2_tiehi _1219__67 (.L_HI(net67));
 sg13g2_tiehi _1205__68 (.L_HI(net68));
 sg13g2_tiehi _1224__69 (.L_HI(net69));
 sg13g2_tiehi _1204__70 (.L_HI(net70));
 sg13g2_tiehi _1218__71 (.L_HI(net71));
 sg13g2_tiehi _1203__72 (.L_HI(net72));
 sg13g2_tiehi _1228__73 (.L_HI(net73));
 sg13g2_tiehi _1202__74 (.L_HI(net74));
 sg13g2_tiehi _1217__75 (.L_HI(net75));
 sg13g2_tiehi _1201__76 (.L_HI(net76));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_gamepad_pmod_demo_5 (.L_LO(net5));
 sg13g2_tielo tt_um_gamepad_pmod_demo_6 (.L_LO(net6));
 sg13g2_tielo tt_um_gamepad_pmod_demo_7 (.L_LO(net7));
 sg13g2_tielo tt_um_gamepad_pmod_demo_8 (.L_LO(net8));
 sg13g2_tielo tt_um_gamepad_pmod_demo_9 (.L_LO(net9));
 sg13g2_tielo tt_um_gamepad_pmod_demo_10 (.L_LO(net10));
 sg13g2_tielo tt_um_gamepad_pmod_demo_11 (.L_LO(net11));
 sg13g2_tielo tt_um_gamepad_pmod_demo_12 (.L_LO(net12));
 sg13g2_tielo tt_um_gamepad_pmod_demo_13 (.L_LO(net13));
 sg13g2_tielo tt_um_gamepad_pmod_demo_14 (.L_LO(net14));
 sg13g2_tielo tt_um_gamepad_pmod_demo_15 (.L_LO(net15));
 sg13g2_tielo tt_um_gamepad_pmod_demo_16 (.L_LO(net16));
 sg13g2_tielo tt_um_gamepad_pmod_demo_17 (.L_LO(net17));
 sg13g2_tielo tt_um_gamepad_pmod_demo_18 (.L_LO(net18));
 sg13g2_tielo tt_um_gamepad_pmod_demo_19 (.L_LO(net19));
 sg13g2_tiehi _1223__20 (.L_HI(net20));
 sg13g2_buf_1 _1302_ (.A(uo_out[6]),
    .X(uo_out[0]));
 sg13g2_buf_1 _1303_ (.A(uo_out[5]),
    .X(uo_out[1]));
 sg13g2_buf_1 _1304_ (.A(uo_out[6]),
    .X(uo_out[2]));
 sg13g2_buf_1 _1305_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1306_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout164 (.A(_0270_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_0263_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_0215_),
    .X(net166));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(_0269_));
 sg13g2_buf_1 fanout168 (.A(_0269_),
    .X(net168));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(_0268_));
 sg13g2_buf_2 fanout170 (.A(_0221_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_0221_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_0220_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_0220_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_0496_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_0212_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_0212_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_0170_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_0136_),
    .X(net179));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(_0544_));
 sg13g2_buf_2 fanout181 (.A(_0544_),
    .X(net181));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(_0492_));
 sg13g2_buf_2 fanout183 (.A(_0492_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_0543_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_0543_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_0491_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_0491_),
    .X(net187));
 sg13g2_buf_4 fanout188 (.X(net188),
    .A(net161));
 sg13g2_buf_4 fanout189 (.X(net189),
    .A(net217));
 sg13g2_buf_2 fanout190 (.A(\pix_y[8] ),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(\pix_y[7] ),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(net218),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(net194),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(net159),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(\pix_y[5] ),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(net223),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(net199),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(net142),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(net220),
    .X(net200));
 sg13g2_buf_1 fanout201 (.A(\pix_y[2] ),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(net203),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(net147),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(net222),
    .X(net204));
 sg13g2_buf_1 fanout205 (.A(\pix_x[6] ),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(net215),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(\pix_x[5] ),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(net209),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(\pix_x[4] ),
    .X(net209));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(\pix_x[3] ));
 sg13g2_buf_4 fanout211 (.X(net211),
    .A(rst_n));
 sg13g2_buf_1 fanout212 (.A(rst_n),
    .X(net212));
 sg13g2_buf_1 input1 (.A(ui_in[4]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[5]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[6]),
    .X(net3));
 sg13g2_tielo tt_um_gamepad_pmod_demo_4 (.L_LO(net4));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\driver.driver.pmod_latch_sync[1] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold2 (.A(\driver.driver.pmod_clk_sync[1] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0017_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0006_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0000_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold6 (.A(\driver.driver.pmod_data_sync[0] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold7 (.A(\driver.driver.pmod_clk_sync[0] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0016_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0045_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold10 (.A(\driver.driver.pmod_latch_sync[0] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0003_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0501_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold13 (.A(\driver.decoder.data_reg[6] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0025_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold15 (.A(\driver.driver.shift_reg[11] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0066_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold17 (.A(\driver.driver.pmod_data_sync[1] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0055_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0004_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0499_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0500_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold22 (.A(\driver.decoder.data_reg[5] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0024_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold24 (.A(\driver.decoder.data_reg[7] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0026_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold26 (.A(\driver.decoder.data_reg[8] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0027_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold28 (.A(\driver.decoder.data_reg[0] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0019_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold30 (.A(\driver.decoder.data_reg[3] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0022_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold32 (.A(\driver.decoder.data_reg[4] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0023_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold34 (.A(\driver.driver.shift_reg[7] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0062_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold36 (.A(\driver.driver.shift_reg[6] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0061_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold38 (.A(\driver.driver.shift_reg[1] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0056_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold40 (.A(\driver.decoder.data_reg[1] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0020_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold42 (.A(\driver.decoder.data_reg[2] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0021_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold44 (.A(\driver.decoder.data_reg[9] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0028_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold46 (.A(\driver.decoder.data_reg[11] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0030_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold48 (.A(\driver.driver.shift_reg[4] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0059_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold50 (.A(\driver.driver.shift_reg[9] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0064_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold52 (.A(\driver.driver.shift_reg[3] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0058_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold54 (.A(\driver.driver.shift_reg[8] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0063_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold56 (.A(\driver.driver.shift_reg[10] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0065_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold58 (.A(\pix_y[1] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0046_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold60 (.A(\driver.decoder.data_reg[10] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0029_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold62 (.A(\driver.driver.shift_reg[5] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0060_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold64 (.A(\driver.driver.shift_reg[2] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0057_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold66 (.A(\pix_y[3] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0108_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0001_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold69 (.A(\pix_x[9] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0510_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold71 (.A(\pix_x[7] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0038_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold73 (.A(\pix_x[0] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0205_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0032_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0013_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0524_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0015_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0532_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0050_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold81 (.A(\pix_x[1] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0498_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold83 (.A(\pix_y[6] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0534_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold85 (.A(\pix_y[9] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0054_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold87 (.A(\pix_x[8] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold88 (.A(\driver.decoder.data_reg[5] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0479_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold90 (.A(\pix_x[5] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0504_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold92 (.A(\pix_y[8] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold93 (.A(\pix_y[7] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0052_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold95 (.A(\pix_y[2] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0522_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold97 (.A(\pix_x[6] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold98 (.A(\pix_y[4] ),
    .X(net223));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_fill_2 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_4 FILLER_14_168 ();
 sg13g2_fill_2 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_185 ();
 sg13g2_decap_8 FILLER_14_192 ();
 sg13g2_decap_8 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_decap_4 FILLER_14_213 ();
 sg13g2_fill_1 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_222 ();
 sg13g2_decap_8 FILLER_14_229 ();
 sg13g2_decap_8 FILLER_14_240 ();
 sg13g2_decap_8 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_254 ();
 sg13g2_decap_8 FILLER_14_261 ();
 sg13g2_decap_8 FILLER_14_268 ();
 sg13g2_decap_8 FILLER_14_275 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_decap_8 FILLER_14_289 ();
 sg13g2_decap_8 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_310 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_decap_8 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_decap_8 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_366 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_387 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_134 ();
 sg13g2_decap_8 FILLER_15_141 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_fill_2 FILLER_15_155 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_fill_1 FILLER_15_196 ();
 sg13g2_fill_2 FILLER_15_210 ();
 sg13g2_fill_1 FILLER_15_244 ();
 sg13g2_decap_4 FILLER_15_250 ();
 sg13g2_fill_1 FILLER_15_254 ();
 sg13g2_decap_8 FILLER_15_265 ();
 sg13g2_decap_8 FILLER_15_272 ();
 sg13g2_decap_8 FILLER_15_279 ();
 sg13g2_decap_8 FILLER_15_286 ();
 sg13g2_decap_8 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_300 ();
 sg13g2_decap_8 FILLER_15_307 ();
 sg13g2_decap_8 FILLER_15_314 ();
 sg13g2_decap_8 FILLER_15_321 ();
 sg13g2_decap_8 FILLER_15_328 ();
 sg13g2_decap_8 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_4 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_66 ();
 sg13g2_fill_1 FILLER_16_73 ();
 sg13g2_fill_1 FILLER_16_85 ();
 sg13g2_fill_2 FILLER_16_115 ();
 sg13g2_decap_4 FILLER_16_124 ();
 sg13g2_decap_4 FILLER_16_148 ();
 sg13g2_fill_1 FILLER_16_152 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_decap_4 FILLER_16_165 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_decap_4 FILLER_16_184 ();
 sg13g2_decap_8 FILLER_16_206 ();
 sg13g2_decap_4 FILLER_16_213 ();
 sg13g2_decap_8 FILLER_16_222 ();
 sg13g2_decap_4 FILLER_16_229 ();
 sg13g2_decap_4 FILLER_16_251 ();
 sg13g2_fill_2 FILLER_16_269 ();
 sg13g2_fill_1 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_4 FILLER_17_35 ();
 sg13g2_decap_4 FILLER_17_67 ();
 sg13g2_fill_1 FILLER_17_81 ();
 sg13g2_decap_8 FILLER_17_94 ();
 sg13g2_fill_2 FILLER_17_101 ();
 sg13g2_decap_8 FILLER_17_108 ();
 sg13g2_decap_4 FILLER_17_115 ();
 sg13g2_fill_2 FILLER_17_124 ();
 sg13g2_decap_8 FILLER_17_136 ();
 sg13g2_decap_8 FILLER_17_143 ();
 sg13g2_decap_8 FILLER_17_150 ();
 sg13g2_decap_8 FILLER_17_157 ();
 sg13g2_fill_1 FILLER_17_164 ();
 sg13g2_decap_8 FILLER_17_202 ();
 sg13g2_fill_2 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_fill_2 FILLER_17_233 ();
 sg13g2_decap_4 FILLER_17_248 ();
 sg13g2_fill_2 FILLER_17_275 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_decap_8 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_decap_8 FILLER_17_311 ();
 sg13g2_decap_8 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_325 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_34 ();
 sg13g2_fill_1 FILLER_18_36 ();
 sg13g2_decap_8 FILLER_18_41 ();
 sg13g2_decap_4 FILLER_18_48 ();
 sg13g2_fill_1 FILLER_18_52 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_4 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_88 ();
 sg13g2_fill_2 FILLER_18_100 ();
 sg13g2_fill_2 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_137 ();
 sg13g2_fill_1 FILLER_18_139 ();
 sg13g2_fill_1 FILLER_18_145 ();
 sg13g2_fill_1 FILLER_18_161 ();
 sg13g2_fill_1 FILLER_18_174 ();
 sg13g2_decap_4 FILLER_18_183 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_4 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_222 ();
 sg13g2_fill_2 FILLER_18_239 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_fill_2 FILLER_18_255 ();
 sg13g2_fill_1 FILLER_18_257 ();
 sg13g2_fill_2 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_decap_4 FILLER_18_270 ();
 sg13g2_fill_2 FILLER_18_274 ();
 sg13g2_decap_8 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_310 ();
 sg13g2_decap_8 FILLER_18_317 ();
 sg13g2_decap_8 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_331 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_4 FILLER_19_52 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_fill_1 FILLER_19_81 ();
 sg13g2_decap_4 FILLER_19_92 ();
 sg13g2_fill_2 FILLER_19_96 ();
 sg13g2_decap_8 FILLER_19_107 ();
 sg13g2_decap_4 FILLER_19_114 ();
 sg13g2_fill_2 FILLER_19_118 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_4 FILLER_19_147 ();
 sg13g2_fill_1 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_172 ();
 sg13g2_decap_4 FILLER_19_180 ();
 sg13g2_fill_1 FILLER_19_184 ();
 sg13g2_decap_4 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_fill_1 FILLER_19_240 ();
 sg13g2_decap_4 FILLER_19_250 ();
 sg13g2_fill_2 FILLER_19_254 ();
 sg13g2_fill_2 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_275 ();
 sg13g2_fill_2 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_32 ();
 sg13g2_fill_2 FILLER_20_39 ();
 sg13g2_fill_1 FILLER_20_41 ();
 sg13g2_fill_1 FILLER_20_86 ();
 sg13g2_fill_2 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_109 ();
 sg13g2_fill_1 FILLER_20_130 ();
 sg13g2_fill_1 FILLER_20_135 ();
 sg13g2_decap_4 FILLER_20_150 ();
 sg13g2_fill_1 FILLER_20_154 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_fill_1 FILLER_20_172 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_decap_4 FILLER_20_189 ();
 sg13g2_fill_2 FILLER_20_197 ();
 sg13g2_decap_8 FILLER_20_204 ();
 sg13g2_decap_8 FILLER_20_211 ();
 sg13g2_decap_4 FILLER_20_222 ();
 sg13g2_fill_2 FILLER_20_226 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_decap_4 FILLER_20_238 ();
 sg13g2_fill_1 FILLER_20_251 ();
 sg13g2_fill_2 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_259 ();
 sg13g2_fill_1 FILLER_20_265 ();
 sg13g2_fill_2 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_297 ();
 sg13g2_decap_8 FILLER_20_304 ();
 sg13g2_decap_8 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_325 ();
 sg13g2_fill_2 FILLER_20_332 ();
 sg13g2_fill_1 FILLER_20_334 ();
 sg13g2_decap_4 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_352 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_8 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_66 ();
 sg13g2_fill_1 FILLER_21_95 ();
 sg13g2_fill_2 FILLER_21_100 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_107 ();
 sg13g2_decap_8 FILLER_21_114 ();
 sg13g2_fill_1 FILLER_21_121 ();
 sg13g2_decap_8 FILLER_21_134 ();
 sg13g2_decap_4 FILLER_21_148 ();
 sg13g2_fill_2 FILLER_21_156 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_decap_8 FILLER_21_164 ();
 sg13g2_fill_2 FILLER_21_171 ();
 sg13g2_fill_1 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_181 ();
 sg13g2_fill_2 FILLER_21_187 ();
 sg13g2_fill_2 FILLER_21_194 ();
 sg13g2_fill_2 FILLER_21_209 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_fill_2 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_fill_1 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_297 ();
 sg13g2_decap_4 FILLER_21_304 ();
 sg13g2_fill_2 FILLER_21_308 ();
 sg13g2_fill_1 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_4 ();
 sg13g2_fill_1 FILLER_22_18 ();
 sg13g2_fill_2 FILLER_22_71 ();
 sg13g2_decap_4 FILLER_22_85 ();
 sg13g2_fill_1 FILLER_22_89 ();
 sg13g2_decap_8 FILLER_22_135 ();
 sg13g2_decap_8 FILLER_22_142 ();
 sg13g2_decap_4 FILLER_22_160 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_decap_4 FILLER_22_191 ();
 sg13g2_fill_2 FILLER_22_195 ();
 sg13g2_decap_8 FILLER_22_202 ();
 sg13g2_decap_4 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_218 ();
 sg13g2_decap_4 FILLER_22_225 ();
 sg13g2_fill_2 FILLER_22_241 ();
 sg13g2_fill_1 FILLER_22_243 ();
 sg13g2_decap_8 FILLER_22_260 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_269 ();
 sg13g2_fill_1 FILLER_22_274 ();
 sg13g2_decap_8 FILLER_22_292 ();
 sg13g2_decap_8 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_306 ();
 sg13g2_decap_4 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_337 ();
 sg13g2_decap_4 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_4 FILLER_22_386 ();
 sg13g2_decap_4 FILLER_22_393 ();
 sg13g2_fill_1 FILLER_22_397 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_19 ();
 sg13g2_decap_8 FILLER_23_40 ();
 sg13g2_fill_2 FILLER_23_47 ();
 sg13g2_fill_1 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_83 ();
 sg13g2_decap_4 FILLER_23_90 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_127 ();
 sg13g2_fill_1 FILLER_23_129 ();
 sg13g2_fill_2 FILLER_23_144 ();
 sg13g2_fill_1 FILLER_23_146 ();
 sg13g2_decap_4 FILLER_23_163 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_decap_8 FILLER_23_173 ();
 sg13g2_decap_4 FILLER_23_180 ();
 sg13g2_fill_2 FILLER_23_184 ();
 sg13g2_decap_4 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_195 ();
 sg13g2_fill_2 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_226 ();
 sg13g2_decap_8 FILLER_23_233 ();
 sg13g2_decap_8 FILLER_23_240 ();
 sg13g2_fill_2 FILLER_23_247 ();
 sg13g2_fill_2 FILLER_23_256 ();
 sg13g2_fill_2 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_291 ();
 sg13g2_fill_1 FILLER_23_346 ();
 sg13g2_fill_2 FILLER_23_362 ();
 sg13g2_fill_1 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_16 ();
 sg13g2_fill_2 FILLER_24_53 ();
 sg13g2_fill_1 FILLER_24_66 ();
 sg13g2_decap_8 FILLER_24_72 ();
 sg13g2_decap_8 FILLER_24_79 ();
 sg13g2_decap_4 FILLER_24_86 ();
 sg13g2_fill_2 FILLER_24_90 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_fill_2 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_fill_1 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_136 ();
 sg13g2_decap_8 FILLER_24_143 ();
 sg13g2_decap_8 FILLER_24_155 ();
 sg13g2_fill_1 FILLER_24_162 ();
 sg13g2_fill_2 FILLER_24_176 ();
 sg13g2_decap_4 FILLER_24_195 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_212 ();
 sg13g2_decap_8 FILLER_24_219 ();
 sg13g2_fill_2 FILLER_24_226 ();
 sg13g2_fill_1 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_275 ();
 sg13g2_decap_4 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_325 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_fill_1 FILLER_25_31 ();
 sg13g2_fill_1 FILLER_25_50 ();
 sg13g2_fill_2 FILLER_25_72 ();
 sg13g2_fill_1 FILLER_25_74 ();
 sg13g2_decap_4 FILLER_25_81 ();
 sg13g2_fill_1 FILLER_25_85 ();
 sg13g2_fill_2 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_115 ();
 sg13g2_fill_1 FILLER_25_134 ();
 sg13g2_decap_4 FILLER_25_140 ();
 sg13g2_fill_1 FILLER_25_144 ();
 sg13g2_fill_2 FILLER_25_153 ();
 sg13g2_fill_1 FILLER_25_155 ();
 sg13g2_decap_4 FILLER_25_178 ();
 sg13g2_fill_2 FILLER_25_182 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_191 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_fill_1 FILLER_25_206 ();
 sg13g2_decap_4 FILLER_25_219 ();
 sg13g2_decap_8 FILLER_25_244 ();
 sg13g2_decap_8 FILLER_25_251 ();
 sg13g2_fill_1 FILLER_25_258 ();
 sg13g2_decap_4 FILLER_25_264 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_fill_1 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_15 ();
 sg13g2_fill_1 FILLER_26_17 ();
 sg13g2_decap_8 FILLER_26_57 ();
 sg13g2_fill_2 FILLER_26_64 ();
 sg13g2_fill_1 FILLER_26_66 ();
 sg13g2_decap_8 FILLER_26_71 ();
 sg13g2_decap_4 FILLER_26_78 ();
 sg13g2_fill_1 FILLER_26_82 ();
 sg13g2_decap_8 FILLER_26_87 ();
 sg13g2_decap_8 FILLER_26_94 ();
 sg13g2_fill_1 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_116 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_132 ();
 sg13g2_decap_8 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_149 ();
 sg13g2_decap_4 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_decap_8 FILLER_26_194 ();
 sg13g2_decap_4 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_decap_8 FILLER_26_223 ();
 sg13g2_fill_2 FILLER_26_230 ();
 sg13g2_fill_1 FILLER_26_232 ();
 sg13g2_decap_8 FILLER_26_254 ();
 sg13g2_decap_8 FILLER_26_272 ();
 sg13g2_decap_8 FILLER_26_279 ();
 sg13g2_decap_8 FILLER_26_297 ();
 sg13g2_decap_8 FILLER_26_304 ();
 sg13g2_decap_4 FILLER_26_311 ();
 sg13g2_fill_2 FILLER_26_315 ();
 sg13g2_fill_2 FILLER_26_321 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_fill_1 FILLER_26_384 ();
 sg13g2_fill_2 FILLER_26_398 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_25 ();
 sg13g2_decap_4 FILLER_27_47 ();
 sg13g2_fill_2 FILLER_27_107 ();
 sg13g2_fill_1 FILLER_27_109 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_121 ();
 sg13g2_decap_8 FILLER_27_142 ();
 sg13g2_decap_8 FILLER_27_149 ();
 sg13g2_decap_8 FILLER_27_172 ();
 sg13g2_decap_4 FILLER_27_179 ();
 sg13g2_fill_1 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_fill_2 FILLER_27_236 ();
 sg13g2_fill_1 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_260 ();
 sg13g2_fill_2 FILLER_27_271 ();
 sg13g2_decap_4 FILLER_27_278 ();
 sg13g2_fill_2 FILLER_27_288 ();
 sg13g2_decap_4 FILLER_27_314 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_21 ();
 sg13g2_fill_2 FILLER_28_46 ();
 sg13g2_decap_4 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_fill_2 FILLER_28_155 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_176 ();
 sg13g2_decap_8 FILLER_28_183 ();
 sg13g2_decap_4 FILLER_28_190 ();
 sg13g2_fill_2 FILLER_28_194 ();
 sg13g2_decap_4 FILLER_28_201 ();
 sg13g2_decap_8 FILLER_28_209 ();
 sg13g2_decap_8 FILLER_28_216 ();
 sg13g2_fill_2 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_225 ();
 sg13g2_decap_8 FILLER_28_239 ();
 sg13g2_fill_2 FILLER_28_246 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_274 ();
 sg13g2_fill_2 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_289 ();
 sg13g2_decap_8 FILLER_28_296 ();
 sg13g2_decap_4 FILLER_28_303 ();
 sg13g2_fill_1 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_338 ();
 sg13g2_fill_2 FILLER_28_398 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_14 ();
 sg13g2_fill_2 FILLER_29_48 ();
 sg13g2_fill_1 FILLER_29_50 ();
 sg13g2_decap_4 FILLER_29_78 ();
 sg13g2_fill_2 FILLER_29_82 ();
 sg13g2_fill_2 FILLER_29_96 ();
 sg13g2_fill_1 FILLER_29_98 ();
 sg13g2_decap_4 FILLER_29_122 ();
 sg13g2_fill_2 FILLER_29_126 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_fill_1 FILLER_29_151 ();
 sg13g2_decap_4 FILLER_29_171 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_187 ();
 sg13g2_decap_4 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_236 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_257 ();
 sg13g2_decap_4 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_fill_2 FILLER_29_315 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_47 ();
 sg13g2_decap_8 FILLER_30_80 ();
 sg13g2_fill_2 FILLER_30_87 ();
 sg13g2_fill_1 FILLER_30_89 ();
 sg13g2_fill_2 FILLER_30_102 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_152 ();
 sg13g2_fill_2 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_fill_1 FILLER_30_190 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_226 ();
 sg13g2_decap_4 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_250 ();
 sg13g2_decap_8 FILLER_30_257 ();
 sg13g2_fill_1 FILLER_30_264 ();
 sg13g2_decap_8 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_381 ();
 sg13g2_fill_2 FILLER_30_391 ();
 sg13g2_fill_1 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_fill_2 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_65 ();
 sg13g2_decap_8 FILLER_31_79 ();
 sg13g2_decap_4 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_120 ();
 sg13g2_decap_4 FILLER_31_127 ();
 sg13g2_fill_2 FILLER_31_131 ();
 sg13g2_decap_8 FILLER_31_146 ();
 sg13g2_decap_4 FILLER_31_153 ();
 sg13g2_fill_2 FILLER_31_157 ();
 sg13g2_fill_2 FILLER_31_169 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_decap_8 FILLER_31_177 ();
 sg13g2_decap_8 FILLER_31_184 ();
 sg13g2_fill_1 FILLER_31_191 ();
 sg13g2_decap_4 FILLER_31_204 ();
 sg13g2_decap_8 FILLER_31_213 ();
 sg13g2_fill_2 FILLER_31_220 ();
 sg13g2_decap_4 FILLER_31_257 ();
 sg13g2_decap_8 FILLER_31_291 ();
 sg13g2_fill_2 FILLER_31_298 ();
 sg13g2_fill_2 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_51 ();
 sg13g2_fill_1 FILLER_32_83 ();
 sg13g2_fill_1 FILLER_32_89 ();
 sg13g2_fill_2 FILLER_32_99 ();
 sg13g2_fill_1 FILLER_32_115 ();
 sg13g2_fill_2 FILLER_32_125 ();
 sg13g2_decap_8 FILLER_32_146 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_decap_4 FILLER_32_158 ();
 sg13g2_fill_1 FILLER_32_162 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_fill_1 FILLER_32_175 ();
 sg13g2_fill_2 FILLER_32_193 ();
 sg13g2_fill_1 FILLER_32_195 ();
 sg13g2_decap_4 FILLER_32_229 ();
 sg13g2_decap_8 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_244 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_fill_1 FILLER_32_266 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_276 ();
 sg13g2_decap_8 FILLER_32_283 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_336 ();
 sg13g2_fill_2 FILLER_32_389 ();
 sg13g2_fill_1 FILLER_32_391 ();
 sg13g2_fill_1 FILLER_32_396 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_4 FILLER_33_70 ();
 sg13g2_fill_1 FILLER_33_74 ();
 sg13g2_fill_2 FILLER_33_101 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_fill_2 FILLER_33_187 ();
 sg13g2_fill_1 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_207 ();
 sg13g2_fill_1 FILLER_33_222 ();
 sg13g2_fill_2 FILLER_33_254 ();
 sg13g2_fill_1 FILLER_33_311 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_351 ();
 sg13g2_fill_1 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_89 ();
 sg13g2_fill_1 FILLER_34_100 ();
 sg13g2_fill_1 FILLER_34_126 ();
 sg13g2_decap_4 FILLER_34_131 ();
 sg13g2_fill_1 FILLER_34_135 ();
 sg13g2_fill_2 FILLER_34_153 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_fill_2 FILLER_34_191 ();
 sg13g2_fill_1 FILLER_34_233 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_4 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_258 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_decap_8 FILLER_34_265 ();
 sg13g2_decap_4 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_276 ();
 sg13g2_decap_4 FILLER_34_289 ();
 sg13g2_fill_2 FILLER_34_336 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_fill_1 FILLER_34_357 ();
 sg13g2_fill_2 FILLER_34_367 ();
 sg13g2_fill_2 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_4 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_fill_1 FILLER_35_206 ();
 sg13g2_decap_4 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_237 ();
 sg13g2_fill_1 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_276 ();
 sg13g2_fill_1 FILLER_35_303 ();
 sg13g2_fill_2 FILLER_35_310 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_fill_2 FILLER_36_145 ();
 sg13g2_decap_8 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_194 ();
 sg13g2_decap_8 FILLER_36_201 ();
 sg13g2_decap_8 FILLER_36_208 ();
 sg13g2_fill_2 FILLER_36_215 ();
 sg13g2_decap_8 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_fill_2 FILLER_36_285 ();
 sg13g2_fill_2 FILLER_36_291 ();
 sg13g2_decap_8 FILLER_36_302 ();
 sg13g2_decap_8 FILLER_36_327 ();
 sg13g2_decap_4 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_decap_4 FILLER_36_354 ();
 sg13g2_fill_1 FILLER_36_358 ();
 sg13g2_decap_8 FILLER_36_376 ();
 sg13g2_decap_8 FILLER_36_383 ();
 sg13g2_decap_8 FILLER_36_390 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_decap_4 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_156 ();
 sg13g2_decap_4 FILLER_37_163 ();
 sg13g2_decap_8 FILLER_37_197 ();
 sg13g2_decap_8 FILLER_37_204 ();
 sg13g2_decap_8 FILLER_37_211 ();
 sg13g2_decap_8 FILLER_37_218 ();
 sg13g2_decap_4 FILLER_37_225 ();
 sg13g2_fill_1 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_268 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_fill_2 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_249 ();
 sg13g2_decap_4 FILLER_38_256 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_277 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_decap_8 FILLER_38_284 ();
 sg13g2_decap_4 FILLER_38_291 ();
 sg13g2_fill_1 FILLER_38_308 ();
 sg13g2_fill_1 FILLER_38_314 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_decap_4 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_353 ();
 sg13g2_decap_8 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_366 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
endmodule
