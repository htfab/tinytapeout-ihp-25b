module tt_um_bleeptrack_prism (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \dist_x[0] ;
 wire \dist_y[0] ;
 wire hsync;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net1;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 sg13g2_inv_1 _438_ (.Y(_390_),
    .A(\hvsync_gen.vpos[3] ));
 sg13g2_inv_1 _439_ (.Y(_391_),
    .A(net46));
 sg13g2_inv_1 _440_ (.Y(_392_),
    .A(\hvsync_gen.hpos[7] ));
 sg13g2_inv_1 _441_ (.Y(_393_),
    .A(net96));
 sg13g2_inv_1 _442_ (.Y(_394_),
    .A(net89));
 sg13g2_inv_1 _443_ (.Y(_395_),
    .A(_006_));
 sg13g2_inv_1 _444_ (.Y(_396_),
    .A(_011_));
 sg13g2_inv_1 _445_ (.Y(_055_),
    .A(net74));
 sg13g2_inv_1 _446_ (.Y(_056_),
    .A(\counter[4] ));
 sg13g2_inv_1 _447_ (.Y(_057_),
    .A(_019_));
 sg13g2_inv_1 _448_ (.Y(_058_),
    .A(\counter[6] ));
 sg13g2_inv_1 _449_ (.Y(_059_),
    .A(\counter[7] ));
 sg13g2_inv_1 _450_ (.Y(_060_),
    .A(\counter[9] ));
 sg13g2_and4_1 _451_ (.A(\hvsync_gen.vpos[7] ),
    .B(\hvsync_gen.vpos[6] ),
    .C(net45),
    .D(\hvsync_gen.vpos[8] ),
    .X(_061_));
 sg13g2_nor3_1 _452_ (.A(\hvsync_gen.vpos[2] ),
    .B(\hvsync_gen.vpos[4] ),
    .C(net76),
    .Y(_062_));
 sg13g2_and4_1 _453_ (.A(\hvsync_gen.vpos[1] ),
    .B(\hvsync_gen.vpos[3] ),
    .C(_061_),
    .D(net77),
    .X(_001_));
 sg13g2_nand2_1 _454_ (.Y(_063_),
    .A(net48),
    .B(\hvsync_gen.hpos[8] ));
 sg13g2_nor2_1 _455_ (.A(net50),
    .B(\hvsync_gen.hpos[4] ),
    .Y(_064_));
 sg13g2_nand2_1 _456_ (.Y(_065_),
    .A(\hvsync_gen.hpos[7] ),
    .B(net48));
 sg13g2_a21o_1 _457_ (.A2(_064_),
    .A1(_393_),
    .B1(_065_),
    .X(_066_));
 sg13g2_nor2_1 _458_ (.A(_392_),
    .B(_393_),
    .Y(_067_));
 sg13g2_nand3_1 _459_ (.B(\hvsync_gen.hpos[4] ),
    .C(_067_),
    .A(net50),
    .Y(_068_));
 sg13g2_nor2b_1 _460_ (.A(\hvsync_gen.hpos[8] ),
    .B_N(net48),
    .Y(_069_));
 sg13g2_a21oi_1 _461_ (.A1(_068_),
    .A2(_069_),
    .Y(_070_),
    .B1(net65));
 sg13g2_a21oi_1 _462_ (.A1(_063_),
    .A2(_066_),
    .Y(_000_),
    .B1(net66));
 sg13g2_a21oi_2 _463_ (.B1(_002_),
    .Y(_071_),
    .A2(_394_),
    .A1(_392_));
 sg13g2_nor3_2 _464_ (.A(net44),
    .B(_061_),
    .C(_071_),
    .Y(_072_));
 sg13g2_and2_1 _465_ (.A(net45),
    .B(net46),
    .X(_073_));
 sg13g2_nand2_1 _466_ (.Y(_074_),
    .A(\hvsync_gen.vpos[5] ),
    .B(\hvsync_gen.vpos[4] ));
 sg13g2_nor2_2 _467_ (.A(\hvsync_gen.vpos[8] ),
    .B(net44),
    .Y(_075_));
 sg13g2_or2_1 _468_ (.X(_076_),
    .B(net44),
    .A(\hvsync_gen.vpos[8] ));
 sg13g2_nand4_1 _469_ (.B(\hvsync_gen.vpos[6] ),
    .C(net45),
    .A(\hvsync_gen.vpos[7] ),
    .Y(_077_),
    .D(net46));
 sg13g2_nand2_1 _470_ (.Y(_078_),
    .A(_075_),
    .B(_077_));
 sg13g2_nor2_1 _471_ (.A(\hvsync_gen.vpos[1] ),
    .B(net47),
    .Y(_079_));
 sg13g2_nor3_1 _472_ (.A(\hvsync_gen.vpos[1] ),
    .B(net47),
    .C(\hvsync_gen.vpos[2] ),
    .Y(_080_));
 sg13g2_nor4_2 _473_ (.A(\hvsync_gen.vpos[1] ),
    .B(net47),
    .C(\hvsync_gen.vpos[3] ),
    .Y(_081_),
    .D(\hvsync_gen.vpos[2] ));
 sg13g2_a21oi_2 _474_ (.B1(_081_),
    .Y(_082_),
    .A2(_077_),
    .A1(_075_));
 sg13g2_a221oi_1 _475_ (.B2(_390_),
    .C1(_074_),
    .B1(_080_),
    .A1(_075_),
    .Y(_083_),
    .A2(_077_));
 sg13g2_o21ai_1 _476_ (.B1(_075_),
    .Y(_084_),
    .A1(_077_),
    .A2(_081_));
 sg13g2_a21o_1 _477_ (.A2(_075_),
    .A1(_074_),
    .B1(_083_),
    .X(_085_));
 sg13g2_xor2_1 _478_ (.B(_085_),
    .A(\hvsync_gen.vpos[6] ),
    .X(_086_));
 sg13g2_nor2_1 _479_ (.A(\hvsync_gen.hpos[7] ),
    .B(\hvsync_gen.hpos[6] ),
    .Y(_087_));
 sg13g2_nor2_1 _480_ (.A(net95),
    .B(\hvsync_gen.hpos[1] ),
    .Y(_088_));
 sg13g2_or2_1 _481_ (.X(_089_),
    .B(\hvsync_gen.hpos[1] ),
    .A(net51));
 sg13g2_nor4_2 _482_ (.A(net51),
    .B(\hvsync_gen.hpos[3] ),
    .C(\hvsync_gen.hpos[2] ),
    .Y(_090_),
    .D(\hvsync_gen.hpos[1] ));
 sg13g2_nor3_1 _483_ (.A(net50),
    .B(\hvsync_gen.hpos[4] ),
    .C(\hvsync_gen.hpos[7] ),
    .Y(_091_));
 sg13g2_a21o_1 _484_ (.A2(_091_),
    .A1(_090_),
    .B1(_087_),
    .X(_092_));
 sg13g2_a221oi_1 _485_ (.B2(_091_),
    .C1(_394_),
    .B1(_090_),
    .A1(_392_),
    .Y(_093_),
    .A2(_393_));
 sg13g2_nor2_1 _486_ (.A(net48),
    .B(_093_),
    .Y(_094_));
 sg13g2_or2_2 _487_ (.X(_095_),
    .B(_093_),
    .A(net49));
 sg13g2_nor2b_1 _488_ (.A(\hvsync_gen.hpos[4] ),
    .B_N(_090_),
    .Y(_096_));
 sg13g2_nand2_1 _489_ (.Y(_097_),
    .A(_064_),
    .B(_090_));
 sg13g2_xnor2_1 _490_ (.Y(_098_),
    .A(_012_),
    .B(_097_));
 sg13g2_mux2_2 _491_ (.A0(\hvsync_gen.hpos[6] ),
    .A1(_098_),
    .S(_095_),
    .X(_099_));
 sg13g2_a22oi_1 _492_ (.Y(_100_),
    .B1(_082_),
    .B2(_055_),
    .A2(_075_),
    .A1(_391_));
 sg13g2_xnor2_1 _493_ (.Y(_101_),
    .A(net45),
    .B(_100_));
 sg13g2_nor2_1 _494_ (.A(_013_),
    .B(_095_),
    .Y(_102_));
 sg13g2_xnor2_1 _495_ (.Y(_103_),
    .A(\hvsync_gen.hpos[5] ),
    .B(_096_));
 sg13g2_a21oi_2 _496_ (.B1(_102_),
    .Y(_104_),
    .A2(_103_),
    .A1(_095_));
 sg13g2_and2_1 _497_ (.A(_101_),
    .B(_104_),
    .X(_105_));
 sg13g2_xnor2_1 _498_ (.Y(_106_),
    .A(net46),
    .B(_082_));
 sg13g2_nand2_1 _499_ (.Y(_107_),
    .A(_015_),
    .B(_094_));
 sg13g2_xnor2_1 _500_ (.Y(_108_),
    .A(\hvsync_gen.hpos[4] ),
    .B(_090_));
 sg13g2_o21ai_1 _501_ (.B1(_107_),
    .Y(_109_),
    .A1(_094_),
    .A2(_108_));
 sg13g2_nor2b_1 _502_ (.A(_109_),
    .B_N(_106_),
    .Y(_110_));
 sg13g2_xor2_1 _503_ (.B(_109_),
    .A(_106_),
    .X(_111_));
 sg13g2_and2_1 _504_ (.A(net51),
    .B(\hvsync_gen.hpos[1] ),
    .X(_112_));
 sg13g2_nor2_1 _505_ (.A(_088_),
    .B(_112_),
    .Y(_113_));
 sg13g2_or3_1 _506_ (.A(net49),
    .B(_007_),
    .C(_093_),
    .X(_114_));
 sg13g2_o21ai_1 _507_ (.B1(_113_),
    .Y(_115_),
    .A1(net49),
    .A2(_093_));
 sg13g2_nand2_1 _508_ (.Y(_116_),
    .A(_114_),
    .B(_115_));
 sg13g2_nand2_2 _509_ (.Y(_117_),
    .A(net82),
    .B(net47));
 sg13g2_nand2b_1 _510_ (.Y(_118_),
    .B(_117_),
    .A_N(_079_));
 sg13g2_mux2_1 _511_ (.A0(_008_),
    .A1(_118_),
    .S(_084_),
    .X(_119_));
 sg13g2_a21oi_1 _512_ (.A1(_114_),
    .A2(_115_),
    .Y(_120_),
    .B1(_119_));
 sg13g2_nand3_1 _513_ (.B(_115_),
    .C(_119_),
    .A(_114_),
    .Y(_121_));
 sg13g2_nand2b_1 _514_ (.Y(_122_),
    .B(_121_),
    .A_N(_120_));
 sg13g2_and2_1 _515_ (.A(net51),
    .B(\dist_y[0] ),
    .X(_123_));
 sg13g2_a21oi_1 _516_ (.A1(_121_),
    .A2(_123_),
    .Y(_124_),
    .B1(_120_));
 sg13g2_o21ai_1 _517_ (.B1(_089_),
    .Y(_125_),
    .A1(net49),
    .A2(_093_));
 sg13g2_xnor2_1 _518_ (.Y(_126_),
    .A(_004_),
    .B(_125_));
 sg13g2_nor2_1 _519_ (.A(_005_),
    .B(_084_),
    .Y(_127_));
 sg13g2_xnor2_1 _520_ (.Y(_128_),
    .A(\hvsync_gen.vpos[2] ),
    .B(_079_));
 sg13g2_a21oi_2 _521_ (.B1(_127_),
    .Y(_129_),
    .A2(_128_),
    .A1(_084_));
 sg13g2_nor2_1 _522_ (.A(_126_),
    .B(_129_),
    .Y(_130_));
 sg13g2_and2_1 _523_ (.A(_126_),
    .B(_129_),
    .X(_131_));
 sg13g2_nand2b_1 _524_ (.Y(_132_),
    .B(\hvsync_gen.vpos[3] ),
    .A_N(_080_));
 sg13g2_nor2_1 _525_ (.A(_017_),
    .B(_084_),
    .Y(_133_));
 sg13g2_a21oi_2 _526_ (.B1(_133_),
    .Y(_134_),
    .A2(_132_),
    .A1(_082_));
 sg13g2_inv_1 _527_ (.Y(_135_),
    .A(_134_));
 sg13g2_nand2_1 _528_ (.Y(_136_),
    .A(_004_),
    .B(_088_));
 sg13g2_xnor2_1 _529_ (.Y(_137_),
    .A(\hvsync_gen.hpos[3] ),
    .B(_136_));
 sg13g2_mux2_2 _530_ (.A0(_016_),
    .A1(_137_),
    .S(_095_),
    .X(_138_));
 sg13g2_nor2_1 _531_ (.A(_134_),
    .B(_138_),
    .Y(_139_));
 sg13g2_nand2_1 _532_ (.Y(_140_),
    .A(_134_),
    .B(_138_));
 sg13g2_xnor2_1 _533_ (.Y(_141_),
    .A(_134_),
    .B(_138_));
 sg13g2_or4_1 _534_ (.A(_124_),
    .B(_130_),
    .C(_131_),
    .D(_141_),
    .X(_142_));
 sg13g2_a21oi_1 _535_ (.A1(_130_),
    .A2(_140_),
    .Y(_143_),
    .B1(_139_));
 sg13g2_a21o_1 _536_ (.A2(_143_),
    .A1(_142_),
    .B1(_111_),
    .X(_144_));
 sg13g2_nor2_1 _537_ (.A(_101_),
    .B(_104_),
    .Y(_145_));
 sg13g2_nor2_1 _538_ (.A(_110_),
    .B(_145_),
    .Y(_146_));
 sg13g2_a21o_1 _539_ (.A2(_146_),
    .A1(_144_),
    .B1(_105_),
    .X(_147_));
 sg13g2_a21o_1 _540_ (.A2(_097_),
    .A1(_067_),
    .B1(_092_),
    .X(_148_));
 sg13g2_nor2_1 _541_ (.A(_087_),
    .B(_095_),
    .Y(_149_));
 sg13g2_nor4_1 _542_ (.A(net48),
    .B(_067_),
    .C(_087_),
    .D(_093_),
    .Y(_150_));
 sg13g2_a21oi_2 _543_ (.B1(_150_),
    .Y(_151_),
    .A2(_148_),
    .A1(_095_));
 sg13g2_a21oi_1 _544_ (.A1(\hvsync_gen.vpos[6] ),
    .A2(_073_),
    .Y(_152_),
    .B1(_076_));
 sg13g2_a21oi_1 _545_ (.A1(_396_),
    .A2(_083_),
    .Y(_153_),
    .B1(_152_));
 sg13g2_xnor2_1 _546_ (.Y(_154_),
    .A(\hvsync_gen.vpos[7] ),
    .B(_153_));
 sg13g2_inv_1 _547_ (.Y(_155_),
    .A(_154_));
 sg13g2_nor2_1 _548_ (.A(_151_),
    .B(_155_),
    .Y(_156_));
 sg13g2_nand2_1 _549_ (.Y(_157_),
    .A(_151_),
    .B(_155_));
 sg13g2_xnor2_1 _550_ (.Y(_158_),
    .A(_151_),
    .B(_154_));
 sg13g2_a22oi_1 _551_ (.Y(_159_),
    .B1(_147_),
    .B2(_158_),
    .A2(_099_),
    .A1(_086_));
 sg13g2_or2_1 _552_ (.X(_160_),
    .B(_099_),
    .A(_086_));
 sg13g2_nand2_1 _553_ (.Y(_161_),
    .A(_158_),
    .B(_160_));
 sg13g2_a21o_1 _554_ (.A2(_161_),
    .A1(_147_),
    .B1(_159_),
    .X(_162_));
 sg13g2_nand3_1 _555_ (.B(_142_),
    .C(_143_),
    .A(_111_),
    .Y(_163_));
 sg13g2_nor2_1 _556_ (.A(net51),
    .B(\dist_y[0] ),
    .Y(_164_));
 sg13g2_mux2_1 _557_ (.A0(_123_),
    .A1(_164_),
    .S(_122_),
    .X(_165_));
 sg13g2_mux2_1 _558_ (.A0(_130_),
    .A1(_131_),
    .S(_141_),
    .X(_166_));
 sg13g2_nand2_1 _559_ (.Y(_167_),
    .A(_124_),
    .B(_166_));
 sg13g2_a22oi_1 _560_ (.Y(_168_),
    .B1(_167_),
    .B2(_142_),
    .A2(_163_),
    .A1(_144_));
 sg13g2_nand2_1 _561_ (.Y(_169_),
    .A(_165_),
    .B(_168_));
 sg13g2_nor2_1 _562_ (.A(_105_),
    .B(_145_),
    .Y(_170_));
 sg13g2_nor2b_1 _563_ (.A(_110_),
    .B_N(_144_),
    .Y(_171_));
 sg13g2_xnor2_1 _564_ (.Y(_172_),
    .A(_170_),
    .B(_171_));
 sg13g2_a22oi_1 _565_ (.Y(_173_),
    .B1(_169_),
    .B2(_172_),
    .A2(_161_),
    .A1(_159_));
 sg13g2_nor3_1 _566_ (.A(_010_),
    .B(_077_),
    .C(_081_),
    .Y(_174_));
 sg13g2_o21ai_1 _567_ (.B1(_010_),
    .Y(_175_),
    .A1(_077_),
    .A2(_081_));
 sg13g2_nand2_1 _568_ (.Y(_176_),
    .A(_084_),
    .B(_175_));
 sg13g2_o21ai_1 _569_ (.B1(_078_),
    .Y(_177_),
    .A1(_174_),
    .A2(_176_));
 sg13g2_a21oi_1 _570_ (.A1(net48),
    .A2(_092_),
    .Y(_178_),
    .B1(_149_));
 sg13g2_xnor2_1 _571_ (.Y(_179_),
    .A(\hvsync_gen.hpos[8] ),
    .B(_178_));
 sg13g2_nand2_1 _572_ (.Y(_180_),
    .A(_177_),
    .B(_179_));
 sg13g2_a21o_1 _573_ (.A2(_099_),
    .A1(_086_),
    .B1(_161_),
    .X(_181_));
 sg13g2_a221oi_1 _574_ (.B2(_146_),
    .C1(_181_),
    .B1(_144_),
    .A1(_101_),
    .Y(_182_),
    .A2(_104_));
 sg13g2_o21ai_1 _575_ (.B1(_157_),
    .Y(_183_),
    .A1(_156_),
    .A2(_160_));
 sg13g2_or2_1 _576_ (.X(_184_),
    .B(_183_),
    .A(_182_));
 sg13g2_nand2_1 _577_ (.Y(_185_),
    .A(\hvsync_gen.hpos[8] ),
    .B(_149_));
 sg13g2_nor2_1 _578_ (.A(_009_),
    .B(_092_),
    .Y(_186_));
 sg13g2_xnor2_1 _579_ (.Y(_187_),
    .A(_002_),
    .B(_186_));
 sg13g2_o21ai_1 _580_ (.B1(_185_),
    .Y(_188_),
    .A1(_094_),
    .A2(_187_));
 sg13g2_a21oi_1 _581_ (.A1(_075_),
    .A2(_077_),
    .Y(_189_),
    .B1(net44));
 sg13g2_or2_1 _582_ (.X(_190_),
    .B(_189_),
    .A(_175_));
 sg13g2_o21ai_1 _583_ (.B1(_190_),
    .Y(_191_),
    .A1(net44),
    .A2(_176_));
 sg13g2_xnor2_1 _584_ (.Y(_192_),
    .A(_188_),
    .B(_191_));
 sg13g2_o21ai_1 _585_ (.B1(_192_),
    .Y(_193_),
    .A1(_182_),
    .A2(_183_));
 sg13g2_and2_1 _586_ (.A(_180_),
    .B(_193_),
    .X(_194_));
 sg13g2_o21ai_1 _587_ (.B1(_192_),
    .Y(_195_),
    .A1(_177_),
    .A2(_179_));
 sg13g2_a22oi_1 _588_ (.Y(_196_),
    .B1(_195_),
    .B2(_184_),
    .A2(_193_),
    .A1(_180_));
 sg13g2_a21o_1 _589_ (.A2(_173_),
    .A1(_162_),
    .B1(_196_),
    .X(_197_));
 sg13g2_a221oi_1 _590_ (.B2(_195_),
    .C1(_196_),
    .B1(_194_),
    .A1(_162_),
    .Y(_198_),
    .A2(_173_));
 sg13g2_xnor2_1 _591_ (.Y(_199_),
    .A(\hvsync_gen.hpos[1] ),
    .B(net50));
 sg13g2_xnor2_1 _592_ (.Y(_200_),
    .A(net45),
    .B(_199_));
 sg13g2_nand2b_1 _593_ (.Y(_201_),
    .B(_200_),
    .A_N(_020_));
 sg13g2_xnor2_1 _594_ (.Y(_202_),
    .A(net46),
    .B(\hvsync_gen.hpos[4] ));
 sg13g2_xnor2_1 _595_ (.Y(_203_),
    .A(net51),
    .B(_202_));
 sg13g2_nand2_1 _596_ (.Y(_204_),
    .A(net51),
    .B(\counter[0] ));
 sg13g2_xnor2_1 _597_ (.Y(_205_),
    .A(\hvsync_gen.hpos[1] ),
    .B(_006_));
 sg13g2_nand2b_1 _598_ (.Y(_206_),
    .B(_205_),
    .A_N(_204_));
 sg13g2_nand2_1 _599_ (.Y(_207_),
    .A(\hvsync_gen.hpos[1] ),
    .B(\counter[1] ));
 sg13g2_xnor2_1 _600_ (.Y(_208_),
    .A(\hvsync_gen.hpos[2] ),
    .B(\counter[2] ));
 sg13g2_a21oi_1 _601_ (.A1(_206_),
    .A2(_207_),
    .Y(_209_),
    .B1(_208_));
 sg13g2_nor2b_1 _602_ (.A(_003_),
    .B_N(\hvsync_gen.hpos[2] ),
    .Y(_210_));
 sg13g2_xor2_1 _603_ (.B(\counter[3] ),
    .A(\hvsync_gen.hpos[3] ),
    .X(_211_));
 sg13g2_o21ai_1 _604_ (.B1(_211_),
    .Y(_212_),
    .A1(_209_),
    .A2(_210_));
 sg13g2_nand2b_1 _605_ (.Y(_213_),
    .B(\hvsync_gen.hpos[3] ),
    .A_N(_018_));
 sg13g2_xnor2_1 _606_ (.Y(_214_),
    .A(\counter[4] ),
    .B(_203_));
 sg13g2_a21oi_1 _607_ (.A1(_212_),
    .A2(_213_),
    .Y(_215_),
    .B1(_214_));
 sg13g2_a21oi_1 _608_ (.A1(_057_),
    .A2(_203_),
    .Y(_216_),
    .B1(_215_));
 sg13g2_xnor2_1 _609_ (.Y(_217_),
    .A(\counter[5] ),
    .B(_200_));
 sg13g2_o21ai_1 _610_ (.B1(_201_),
    .Y(_218_),
    .A1(_216_),
    .A2(_217_));
 sg13g2_xor2_1 _611_ (.B(\counter[6] ),
    .A(\hvsync_gen.hpos[6] ),
    .X(_219_));
 sg13g2_xor2_1 _612_ (.B(\hvsync_gen.hpos[2] ),
    .A(\hvsync_gen.vpos[6] ),
    .X(_220_));
 sg13g2_xnor2_1 _613_ (.Y(_221_),
    .A(_219_),
    .B(_220_));
 sg13g2_and2_1 _614_ (.A(_218_),
    .B(_221_),
    .X(_222_));
 sg13g2_xor2_1 _615_ (.B(_217_),
    .A(_216_),
    .X(_223_));
 sg13g2_and3_1 _616_ (.X(_224_),
    .A(_212_),
    .B(_213_),
    .C(_214_));
 sg13g2_o21ai_1 _617_ (.B1(_221_),
    .Y(_225_),
    .A1(_058_),
    .A2(_021_));
 sg13g2_xor2_1 _618_ (.B(\counter[7] ),
    .A(\hvsync_gen.hpos[7] ),
    .X(_226_));
 sg13g2_xor2_1 _619_ (.B(\hvsync_gen.hpos[3] ),
    .A(\hvsync_gen.vpos[7] ),
    .X(_227_));
 sg13g2_xnor2_1 _620_ (.Y(_228_),
    .A(_226_),
    .B(_227_));
 sg13g2_xnor2_1 _621_ (.Y(_229_),
    .A(_225_),
    .B(_228_));
 sg13g2_or3_1 _622_ (.A(_209_),
    .B(_210_),
    .C(_211_),
    .X(_230_));
 sg13g2_nand2_1 _623_ (.Y(_231_),
    .A(_212_),
    .B(_230_));
 sg13g2_o21ai_1 _624_ (.B1(_231_),
    .Y(_232_),
    .A1(_215_),
    .A2(_224_));
 sg13g2_nor4_1 _625_ (.A(_222_),
    .B(_223_),
    .C(_229_),
    .D(_232_),
    .Y(_233_));
 sg13g2_o21ai_1 _626_ (.B1(_233_),
    .Y(_234_),
    .A1(_218_),
    .A2(_221_));
 sg13g2_xor2_1 _627_ (.B(_205_),
    .A(_204_),
    .X(_235_));
 sg13g2_nor2_1 _628_ (.A(_234_),
    .B(_235_),
    .Y(_236_));
 sg13g2_o21ai_1 _629_ (.B1(_072_),
    .Y(_237_),
    .A1(_198_),
    .A2(_236_));
 sg13g2_nand3_1 _630_ (.B(_114_),
    .C(_115_),
    .A(\counter[1] ),
    .Y(_238_));
 sg13g2_a21o_1 _631_ (.A2(_115_),
    .A1(_114_),
    .B1(\counter[1] ),
    .X(_239_));
 sg13g2_a21oi_1 _632_ (.A1(_238_),
    .A2(_239_),
    .Y(_240_),
    .B1(_119_));
 sg13g2_a21oi_1 _633_ (.A1(_395_),
    .A2(_116_),
    .Y(_241_),
    .B1(_240_));
 sg13g2_xor2_1 _634_ (.B(_126_),
    .A(_003_),
    .X(_242_));
 sg13g2_nand2b_1 _635_ (.Y(_243_),
    .B(_242_),
    .A_N(_129_));
 sg13g2_xor2_1 _636_ (.B(_242_),
    .A(_129_),
    .X(_244_));
 sg13g2_nor2_1 _637_ (.A(_241_),
    .B(_244_),
    .Y(_245_));
 sg13g2_xor2_1 _638_ (.B(_244_),
    .A(_241_),
    .X(_246_));
 sg13g2_nand3_1 _639_ (.B(_238_),
    .C(_239_),
    .A(_119_),
    .Y(_247_));
 sg13g2_xor2_1 _640_ (.B(\counter[0] ),
    .A(net51),
    .X(_248_));
 sg13g2_nand2_1 _641_ (.Y(_249_),
    .A(net47),
    .B(_248_));
 sg13g2_nand2_1 _642_ (.Y(_250_),
    .A(_204_),
    .B(_249_));
 sg13g2_nand2_1 _643_ (.Y(_251_),
    .A(_247_),
    .B(_250_));
 sg13g2_nor2_1 _644_ (.A(_240_),
    .B(_251_),
    .Y(_252_));
 sg13g2_xnor2_1 _645_ (.Y(_253_),
    .A(_246_),
    .B(_252_));
 sg13g2_a21oi_2 _646_ (.B1(_237_),
    .Y(uo_out[4]),
    .A2(_253_),
    .A1(_198_));
 sg13g2_nand3_1 _647_ (.B(_207_),
    .C(_208_),
    .A(_206_),
    .Y(_254_));
 sg13g2_nand2b_1 _648_ (.Y(_255_),
    .B(_254_),
    .A_N(_209_));
 sg13g2_nor2_1 _649_ (.A(_234_),
    .B(_255_),
    .Y(_256_));
 sg13g2_o21ai_1 _650_ (.B1(_072_),
    .Y(_257_),
    .A1(_198_),
    .A2(_256_));
 sg13g2_xnor2_1 _651_ (.Y(_258_),
    .A(net47),
    .B(_248_));
 sg13g2_a21oi_2 _652_ (.B1(_257_),
    .Y(uo_out[0]),
    .A2(_258_),
    .A1(_198_));
 sg13g2_xnor2_1 _653_ (.Y(_259_),
    .A(\counter[6] ),
    .B(_099_));
 sg13g2_nor2b_1 _654_ (.A(_086_),
    .B_N(_259_),
    .Y(_260_));
 sg13g2_xor2_1 _655_ (.B(_259_),
    .A(_086_),
    .X(_261_));
 sg13g2_xnor2_1 _656_ (.Y(_262_),
    .A(\counter[5] ),
    .B(_104_));
 sg13g2_nand2b_1 _657_ (.Y(_263_),
    .B(_262_),
    .A_N(_101_));
 sg13g2_or2_1 _658_ (.X(_264_),
    .B(_104_),
    .A(_020_));
 sg13g2_a21oi_2 _659_ (.B1(_261_),
    .Y(_265_),
    .A2(_264_),
    .A1(_263_));
 sg13g2_xnor2_1 _660_ (.Y(_266_),
    .A(_056_),
    .B(_109_));
 sg13g2_inv_1 _661_ (.Y(_267_),
    .A(_266_));
 sg13g2_xor2_1 _662_ (.B(_266_),
    .A(_106_),
    .X(_268_));
 sg13g2_nor2_1 _663_ (.A(_018_),
    .B(_138_),
    .Y(_269_));
 sg13g2_xnor2_1 _664_ (.Y(_270_),
    .A(\counter[3] ),
    .B(_138_));
 sg13g2_a21oi_1 _665_ (.A1(_135_),
    .A2(_270_),
    .Y(_271_),
    .B1(_269_));
 sg13g2_nor2_1 _666_ (.A(_268_),
    .B(_271_),
    .Y(_272_));
 sg13g2_xnor2_1 _667_ (.Y(_273_),
    .A(_268_),
    .B(_271_));
 sg13g2_xnor2_1 _668_ (.Y(_274_),
    .A(_135_),
    .B(_270_));
 sg13g2_inv_1 _669_ (.Y(_275_),
    .A(_274_));
 sg13g2_o21ai_1 _670_ (.B1(_243_),
    .Y(_276_),
    .A1(_003_),
    .A2(_126_));
 sg13g2_a221oi_1 _671_ (.B2(_276_),
    .C1(_245_),
    .B1(_275_),
    .A1(_246_),
    .Y(_277_),
    .A2(_252_));
 sg13g2_nor2_1 _672_ (.A(_275_),
    .B(_276_),
    .Y(_278_));
 sg13g2_or3_1 _673_ (.A(_273_),
    .B(_277_),
    .C(_278_),
    .X(_279_));
 sg13g2_xor2_1 _674_ (.B(_262_),
    .A(_101_),
    .X(_280_));
 sg13g2_inv_1 _675_ (.Y(_281_),
    .A(_280_));
 sg13g2_nor2_1 _676_ (.A(_019_),
    .B(_109_),
    .Y(_282_));
 sg13g2_a21oi_1 _677_ (.A1(_106_),
    .A2(_267_),
    .Y(_283_),
    .B1(_282_));
 sg13g2_a21o_1 _678_ (.A2(_267_),
    .A1(_106_),
    .B1(_282_),
    .X(_284_));
 sg13g2_a21oi_1 _679_ (.A1(_281_),
    .A2(_284_),
    .Y(_285_),
    .B1(_272_));
 sg13g2_nor2_1 _680_ (.A(_281_),
    .B(_284_),
    .Y(_286_));
 sg13g2_a21o_1 _681_ (.A2(_285_),
    .A1(_279_),
    .B1(_286_),
    .X(_287_));
 sg13g2_nand3_1 _682_ (.B(_263_),
    .C(_264_),
    .A(_261_),
    .Y(_288_));
 sg13g2_nand2b_1 _683_ (.Y(_289_),
    .B(_288_),
    .A_N(_265_));
 sg13g2_a221oi_1 _684_ (.B2(_279_),
    .C1(_289_),
    .B1(_285_),
    .A1(_280_),
    .Y(_290_),
    .A2(_283_));
 sg13g2_nor2_1 _685_ (.A(_021_),
    .B(_099_),
    .Y(_291_));
 sg13g2_nor2_1 _686_ (.A(_260_),
    .B(_291_),
    .Y(_292_));
 sg13g2_nand2_1 _687_ (.Y(_293_),
    .A(\counter[7] ),
    .B(_151_));
 sg13g2_xnor2_1 _688_ (.Y(_294_),
    .A(\counter[7] ),
    .B(_151_));
 sg13g2_xnor2_1 _689_ (.Y(_295_),
    .A(_155_),
    .B(_294_));
 sg13g2_nor2b_1 _690_ (.A(_292_),
    .B_N(_295_),
    .Y(_296_));
 sg13g2_xnor2_1 _691_ (.Y(_297_),
    .A(_292_),
    .B(_295_));
 sg13g2_inv_1 _692_ (.Y(_298_),
    .A(_297_));
 sg13g2_o21ai_1 _693_ (.B1(_298_),
    .Y(_299_),
    .A1(_265_),
    .A2(_290_));
 sg13g2_nor3_1 _694_ (.A(_265_),
    .B(_290_),
    .C(_298_),
    .Y(_300_));
 sg13g2_nor2b_1 _695_ (.A(_300_),
    .B_N(_198_),
    .Y(_301_));
 sg13g2_a21oi_2 _696_ (.B1(_237_),
    .Y(uo_out[5]),
    .A2(_301_),
    .A1(_299_));
 sg13g2_o21ai_1 _697_ (.B1(_273_),
    .Y(_302_),
    .A1(_277_),
    .A2(_278_));
 sg13g2_nand2_1 _698_ (.Y(_303_),
    .A(_279_),
    .B(_302_));
 sg13g2_a21oi_2 _699_ (.B1(_257_),
    .Y(uo_out[1]),
    .A2(_303_),
    .A1(_198_));
 sg13g2_o21ai_1 _700_ (.B1(_293_),
    .Y(_304_),
    .A1(_154_),
    .A2(_294_));
 sg13g2_and2_1 _701_ (.A(\counter[8] ),
    .B(_179_),
    .X(_305_));
 sg13g2_xor2_1 _702_ (.B(_179_),
    .A(\counter[8] ),
    .X(_306_));
 sg13g2_xor2_1 _703_ (.B(_306_),
    .A(_177_),
    .X(_307_));
 sg13g2_a21oi_1 _704_ (.A1(_304_),
    .A2(_307_),
    .Y(_308_),
    .B1(_296_));
 sg13g2_a221oi_1 _705_ (.B2(_307_),
    .C1(_296_),
    .B1(_304_),
    .A1(_265_),
    .Y(_309_),
    .A2(_297_));
 sg13g2_nor2_1 _706_ (.A(_304_),
    .B(_307_),
    .Y(_310_));
 sg13g2_nand2_1 _707_ (.Y(_311_),
    .A(_288_),
    .B(_297_));
 sg13g2_a221oi_1 _708_ (.B2(_308_),
    .C1(_310_),
    .B1(_311_),
    .A1(_287_),
    .Y(_312_),
    .A2(_309_));
 sg13g2_a21oi_1 _709_ (.A1(_177_),
    .A2(_306_),
    .Y(_313_),
    .B1(_305_));
 sg13g2_xnor2_1 _710_ (.Y(_314_),
    .A(\counter[9] ),
    .B(_192_));
 sg13g2_xnor2_1 _711_ (.Y(_315_),
    .A(_313_),
    .B(_314_));
 sg13g2_or2_1 _712_ (.X(_316_),
    .B(_315_),
    .A(_312_));
 sg13g2_a221oi_1 _713_ (.B2(_315_),
    .C1(_197_),
    .B1(_312_),
    .A1(_194_),
    .Y(_317_),
    .A2(_195_));
 sg13g2_a21oi_2 _714_ (.B1(_237_),
    .Y(uo_out[6]),
    .A2(_317_),
    .A1(_316_));
 sg13g2_xnor2_1 _715_ (.Y(_318_),
    .A(_287_),
    .B(_289_));
 sg13g2_a21oi_2 _716_ (.B1(_257_),
    .Y(uo_out[2]),
    .A2(_318_),
    .A1(_198_));
 sg13g2_and3_2 _717_ (.X(_319_),
    .A(\hvsync_gen.hpos[3] ),
    .B(\hvsync_gen.hpos[2] ),
    .C(_112_));
 sg13g2_and2_1 _718_ (.A(net94),
    .B(_319_),
    .X(_320_));
 sg13g2_nor4_1 _719_ (.A(net50),
    .B(\hvsync_gen.hpos[7] ),
    .C(\hvsync_gen.hpos[6] ),
    .D(_063_),
    .Y(_321_));
 sg13g2_and2_1 _720_ (.A(_320_),
    .B(_321_),
    .X(_322_));
 sg13g2_nor2b_1 _721_ (.A(_322_),
    .B_N(net52),
    .Y(_323_));
 sg13g2_nand2b_1 _722_ (.Y(_324_),
    .B(net52),
    .A_N(_322_));
 sg13g2_and2_1 _723_ (.A(net62),
    .B(net41),
    .X(_025_));
 sg13g2_and2_1 _724_ (.A(_113_),
    .B(net42),
    .X(_026_));
 sg13g2_o21ai_1 _725_ (.B1(net53),
    .Y(_325_),
    .A1(net88),
    .A2(_112_));
 sg13g2_a21oi_1 _726_ (.A1(net88),
    .A2(_112_),
    .Y(_027_),
    .B1(_325_));
 sg13g2_nand2b_1 _727_ (.Y(_326_),
    .B(_112_),
    .A_N(net92));
 sg13g2_xor2_1 _728_ (.B(_326_),
    .A(\hvsync_gen.hpos[3] ),
    .X(_327_));
 sg13g2_nor2_1 _729_ (.A(_324_),
    .B(net93),
    .Y(_028_));
 sg13g2_o21ai_1 _730_ (.B1(net52),
    .Y(_328_),
    .A1(net94),
    .A2(_319_));
 sg13g2_nor2_1 _731_ (.A(_320_),
    .B(_328_),
    .Y(_029_));
 sg13g2_nor2b_1 _732_ (.A(net68),
    .B_N(_319_),
    .Y(_329_));
 sg13g2_o21ai_1 _733_ (.B1(net41),
    .Y(_330_),
    .A1(net50),
    .A2(_329_));
 sg13g2_a21oi_1 _734_ (.A1(net50),
    .A2(_329_),
    .Y(_030_),
    .B1(_330_));
 sg13g2_nand2_1 _735_ (.Y(_331_),
    .A(net50),
    .B(_320_));
 sg13g2_xnor2_1 _736_ (.Y(_332_),
    .A(_393_),
    .B(_331_));
 sg13g2_nor2_1 _737_ (.A(_324_),
    .B(_332_),
    .Y(_031_));
 sg13g2_nor2_1 _738_ (.A(net83),
    .B(_331_),
    .Y(_333_));
 sg13g2_o21ai_1 _739_ (.B1(net41),
    .Y(_334_),
    .A1(\hvsync_gen.hpos[7] ),
    .A2(_333_));
 sg13g2_a21oi_1 _740_ (.A1(\hvsync_gen.hpos[7] ),
    .A2(_333_),
    .Y(_032_),
    .B1(_334_));
 sg13g2_nand2b_1 _741_ (.Y(_335_),
    .B(_319_),
    .A_N(_068_));
 sg13g2_o21ai_1 _742_ (.B1(net41),
    .Y(_336_),
    .A1(_394_),
    .A2(_335_));
 sg13g2_a21oi_1 _743_ (.A1(_394_),
    .A2(_335_),
    .Y(_033_),
    .B1(_336_));
 sg13g2_nor2_1 _744_ (.A(net73),
    .B(_335_),
    .Y(_337_));
 sg13g2_o21ai_1 _745_ (.B1(net41),
    .Y(_338_),
    .A1(net48),
    .A2(_337_));
 sg13g2_a21oi_1 _746_ (.A1(net48),
    .A2(_337_),
    .Y(_034_),
    .B1(_338_));
 sg13g2_and2_1 _747_ (.A(net53),
    .B(_023_),
    .X(_035_));
 sg13g2_nand2_1 _748_ (.Y(_339_),
    .A(\counter[1] ),
    .B(\counter[0] ));
 sg13g2_o21ai_1 _749_ (.B1(net53),
    .Y(_340_),
    .A1(\counter[1] ),
    .A2(\counter[0] ));
 sg13g2_nor2b_1 _750_ (.A(_340_),
    .B_N(_339_),
    .Y(_036_));
 sg13g2_xnor2_1 _751_ (.Y(_341_),
    .A(\counter[2] ),
    .B(_339_));
 sg13g2_and2_1 _752_ (.A(net53),
    .B(_341_),
    .X(_037_));
 sg13g2_nor2_1 _753_ (.A(_003_),
    .B(_339_),
    .Y(_342_));
 sg13g2_o21ai_1 _754_ (.B1(net53),
    .Y(_343_),
    .A1(\counter[3] ),
    .A2(_342_));
 sg13g2_a21oi_1 _755_ (.A1(\counter[3] ),
    .A2(_342_),
    .Y(_038_),
    .B1(_343_));
 sg13g2_nand4_1 _756_ (.B(\counter[1] ),
    .C(\counter[0] ),
    .A(\counter[2] ),
    .Y(_344_),
    .D(\counter[3] ));
 sg13g2_nor2_1 _757_ (.A(_056_),
    .B(_344_),
    .Y(_345_));
 sg13g2_o21ai_1 _758_ (.B1(net53),
    .Y(_346_),
    .A1(_056_),
    .A2(_344_));
 sg13g2_a21oi_1 _759_ (.A1(_056_),
    .A2(_344_),
    .Y(_039_),
    .B1(_346_));
 sg13g2_nor2_1 _760_ (.A(_019_),
    .B(_344_),
    .Y(_347_));
 sg13g2_o21ai_1 _761_ (.B1(net53),
    .Y(_348_),
    .A1(\counter[5] ),
    .A2(_347_));
 sg13g2_a21oi_1 _762_ (.A1(\counter[5] ),
    .A2(_347_),
    .Y(_040_),
    .B1(_348_));
 sg13g2_nand2_2 _763_ (.Y(_349_),
    .A(\counter[5] ),
    .B(_345_));
 sg13g2_o21ai_1 _764_ (.B1(net52),
    .Y(_350_),
    .A1(_058_),
    .A2(_349_));
 sg13g2_a21oi_1 _765_ (.A1(_058_),
    .A2(_349_),
    .Y(_041_),
    .B1(_350_));
 sg13g2_nor2_1 _766_ (.A(_021_),
    .B(_349_),
    .Y(_351_));
 sg13g2_o21ai_1 _767_ (.B1(net52),
    .Y(_352_),
    .A1(\counter[7] ),
    .A2(_351_));
 sg13g2_a21oi_1 _768_ (.A1(\counter[7] ),
    .A2(_351_),
    .Y(_042_),
    .B1(_352_));
 sg13g2_nor3_1 _769_ (.A(_058_),
    .B(_059_),
    .C(_349_),
    .Y(_353_));
 sg13g2_or2_1 _770_ (.X(_354_),
    .B(_353_),
    .A(\counter[8] ));
 sg13g2_nand2_1 _771_ (.Y(_355_),
    .A(\counter[8] ),
    .B(_353_));
 sg13g2_and3_1 _772_ (.X(_043_),
    .A(net52),
    .B(_354_),
    .C(_355_));
 sg13g2_o21ai_1 _773_ (.B1(net52),
    .Y(_356_),
    .A1(_060_),
    .A2(_355_));
 sg13g2_a21oi_1 _774_ (.A1(_060_),
    .A2(_355_),
    .Y(_044_),
    .B1(_356_));
 sg13g2_nor3_1 _775_ (.A(net45),
    .B(net46),
    .C(\hvsync_gen.vpos[8] ),
    .Y(_357_));
 sg13g2_nand2_1 _776_ (.Y(_358_),
    .A(\hvsync_gen.vpos[3] ),
    .B(\hvsync_gen.vpos[2] ));
 sg13g2_nor4_1 _777_ (.A(\hvsync_gen.vpos[1] ),
    .B(net47),
    .C(\hvsync_gen.vpos[6] ),
    .D(_358_),
    .Y(_359_));
 sg13g2_nand3_1 _778_ (.B(_357_),
    .C(_359_),
    .A(net44),
    .Y(_360_));
 sg13g2_o21ai_1 _779_ (.B1(net52),
    .Y(_361_),
    .A1(\hvsync_gen.vpos[7] ),
    .A2(_360_));
 sg13g2_inv_1 _780_ (.Y(_362_),
    .A(_361_));
 sg13g2_nand2_2 _781_ (.Y(_363_),
    .A(_322_),
    .B(_362_));
 sg13g2_inv_1 _782_ (.Y(_364_),
    .A(_363_));
 sg13g2_a22oi_1 _783_ (.Y(_365_),
    .B1(_364_),
    .B2(net63),
    .A2(net42),
    .A1(net47));
 sg13g2_inv_1 _784_ (.Y(_045_),
    .A(net64));
 sg13g2_nand2_1 _785_ (.Y(_366_),
    .A(net82),
    .B(net42));
 sg13g2_o21ai_1 _786_ (.B1(_366_),
    .Y(_046_),
    .A1(_118_),
    .A2(_363_));
 sg13g2_nor2_1 _787_ (.A(_117_),
    .B(net42),
    .Y(_367_));
 sg13g2_nor2_2 _788_ (.A(net41),
    .B(_362_),
    .Y(_368_));
 sg13g2_xnor2_1 _789_ (.Y(_369_),
    .A(net87),
    .B(_367_));
 sg13g2_nor2_1 _790_ (.A(_368_),
    .B(_369_),
    .Y(_047_));
 sg13g2_nand2_1 _791_ (.Y(_370_),
    .A(\hvsync_gen.vpos[3] ),
    .B(net42));
 sg13g2_nor2_1 _792_ (.A(net79),
    .B(_117_),
    .Y(_371_));
 sg13g2_xnor2_1 _793_ (.Y(_372_),
    .A(\hvsync_gen.vpos[3] ),
    .B(_371_));
 sg13g2_o21ai_1 _794_ (.B1(_370_),
    .Y(_048_),
    .A1(_363_),
    .A2(net80));
 sg13g2_nand2_1 _795_ (.Y(_373_),
    .A(net46),
    .B(net42));
 sg13g2_nor2_2 _796_ (.A(_117_),
    .B(_358_),
    .Y(_374_));
 sg13g2_xnor2_1 _797_ (.Y(_375_),
    .A(_055_),
    .B(_374_));
 sg13g2_o21ai_1 _798_ (.B1(_373_),
    .Y(_049_),
    .A1(_363_),
    .A2(_375_));
 sg13g2_nand2_1 _799_ (.Y(_376_),
    .A(net45),
    .B(net42));
 sg13g2_a21oi_1 _800_ (.A1(net46),
    .A2(_374_),
    .Y(_377_),
    .B1(net45));
 sg13g2_nand2_1 _801_ (.Y(_378_),
    .A(_073_),
    .B(_374_));
 sg13g2_nand2b_1 _802_ (.Y(_379_),
    .B(_378_),
    .A_N(_377_));
 sg13g2_o21ai_1 _803_ (.B1(_376_),
    .Y(_050_),
    .A1(_363_),
    .A2(_379_));
 sg13g2_nor2_1 _804_ (.A(net41),
    .B(_378_),
    .Y(_380_));
 sg13g2_xnor2_1 _805_ (.Y(_381_),
    .A(net91),
    .B(_380_));
 sg13g2_nor2_1 _806_ (.A(_368_),
    .B(_381_),
    .Y(_051_));
 sg13g2_nand2_1 _807_ (.Y(_382_),
    .A(\hvsync_gen.vpos[7] ),
    .B(net41));
 sg13g2_nor2_1 _808_ (.A(net70),
    .B(_378_),
    .Y(_383_));
 sg13g2_xnor2_1 _809_ (.Y(_384_),
    .A(\hvsync_gen.vpos[7] ),
    .B(_383_));
 sg13g2_o21ai_1 _810_ (.B1(_382_),
    .Y(_052_),
    .A1(_363_),
    .A2(net71));
 sg13g2_nand3_1 _811_ (.B(net97),
    .C(_380_),
    .A(\hvsync_gen.vpos[7] ),
    .Y(_385_));
 sg13g2_xor2_1 _812_ (.B(net98),
    .A(net85),
    .X(_386_));
 sg13g2_nor2_1 _813_ (.A(_368_),
    .B(_386_),
    .Y(_053_));
 sg13g2_nand2_1 _814_ (.Y(_387_),
    .A(net44),
    .B(net42));
 sg13g2_nor4_1 _815_ (.A(net86),
    .B(_077_),
    .C(_117_),
    .D(_358_),
    .Y(_388_));
 sg13g2_xnor2_1 _816_ (.Y(_389_),
    .A(net44),
    .B(_388_));
 sg13g2_o21ai_1 _817_ (.B1(_387_),
    .Y(_054_),
    .A1(_363_),
    .A2(_389_));
 sg13g2_dfrbp_1 _818_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net37),
    .D(_025_),
    .Q_N(_024_),
    .Q(\dist_x[0] ));
 sg13g2_dfrbp_1 _819_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net36),
    .D(_026_),
    .Q_N(_007_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _820_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net35),
    .D(_027_),
    .Q_N(_004_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _821_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net34),
    .D(_028_),
    .Q_N(_016_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _822_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net33),
    .D(_029_),
    .Q_N(_015_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _823_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net32),
    .D(net69),
    .Q_N(_013_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _824_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net31),
    .D(_031_),
    .Q_N(_012_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _825_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net30),
    .D(net84),
    .Q_N(_403_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _826_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net29),
    .D(_033_),
    .Q_N(_009_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _827_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net28),
    .D(_034_),
    .Q_N(_002_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _828_ (.CLK(net43),
    .RESET_B(net27),
    .D(_035_),
    .Q_N(_023_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _829_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net26),
    .D(_036_),
    .Q_N(_006_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _830_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net25),
    .D(_037_),
    .Q_N(_003_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _831_ (.CLK(net43),
    .RESET_B(net24),
    .D(_038_),
    .Q_N(_018_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _832_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net23),
    .D(_039_),
    .Q_N(_019_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _833_ (.CLK(net43),
    .RESET_B(net22),
    .D(_040_),
    .Q_N(_020_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _834_ (.CLK(net43),
    .RESET_B(net21),
    .D(_041_),
    .Q_N(_021_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _835_ (.CLK(net43),
    .RESET_B(net20),
    .D(_042_),
    .Q_N(_402_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _836_ (.CLK(net43),
    .RESET_B(net19),
    .D(_043_),
    .Q_N(_401_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _837_ (.CLK(net43),
    .RESET_B(net61),
    .D(_044_),
    .Q_N(_404_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _838_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net18),
    .D(net67),
    .Q_N(_400_),
    .Q(hsync));
 sg13g2_dfrbp_1 _839_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net17),
    .D(_045_),
    .Q_N(_022_),
    .Q(\dist_y[0] ));
 sg13g2_dfrbp_1 _840_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net59),
    .D(_046_),
    .Q_N(_008_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _841_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net57),
    .D(_047_),
    .Q_N(_005_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _842_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net55),
    .D(net81),
    .Q_N(_017_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _843_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net40),
    .D(net75),
    .Q_N(_014_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _844_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net38),
    .D(_050_),
    .Q_N(_399_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _845_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net58),
    .D(_051_),
    .Q_N(_011_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _846_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net54),
    .D(net72),
    .Q_N(_398_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _847_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net60),
    .D(_053_),
    .Q_N(_010_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _848_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net56),
    .D(_054_),
    .Q_N(_405_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _849_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net39),
    .D(net78),
    .Q_N(_397_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_tiehi _838__18 (.L_HI(net18));
 sg13g2_tiehi _836__19 (.L_HI(net19));
 sg13g2_tiehi _835__20 (.L_HI(net20));
 sg13g2_tiehi _834__21 (.L_HI(net21));
 sg13g2_tiehi _833__22 (.L_HI(net22));
 sg13g2_tiehi _832__23 (.L_HI(net23));
 sg13g2_tiehi _831__24 (.L_HI(net24));
 sg13g2_tiehi _830__25 (.L_HI(net25));
 sg13g2_tiehi _829__26 (.L_HI(net26));
 sg13g2_tiehi _828__27 (.L_HI(net27));
 sg13g2_tiehi _827__28 (.L_HI(net28));
 sg13g2_tiehi _826__29 (.L_HI(net29));
 sg13g2_tiehi _825__30 (.L_HI(net30));
 sg13g2_tiehi _824__31 (.L_HI(net31));
 sg13g2_tiehi _823__32 (.L_HI(net32));
 sg13g2_tiehi _822__33 (.L_HI(net33));
 sg13g2_tiehi _821__34 (.L_HI(net34));
 sg13g2_tiehi _820__35 (.L_HI(net35));
 sg13g2_tiehi _819__36 (.L_HI(net36));
 sg13g2_tiehi _818__37 (.L_HI(net37));
 sg13g2_tiehi _844__38 (.L_HI(net38));
 sg13g2_tiehi _849__39 (.L_HI(net39));
 sg13g2_tiehi _843__40 (.L_HI(net40));
 sg13g2_tiehi _846__41 (.L_HI(net54));
 sg13g2_tiehi _842__42 (.L_HI(net55));
 sg13g2_tiehi _848__43 (.L_HI(net56));
 sg13g2_tiehi _841__44 (.L_HI(net57));
 sg13g2_tiehi _845__45 (.L_HI(net58));
 sg13g2_tiehi _840__46 (.L_HI(net59));
 sg13g2_tiehi _847__47 (.L_HI(net60));
 sg13g2_tiehi _837__48 (.L_HI(net61));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_bleeptrack_prism_2 (.L_LO(net2));
 sg13g2_tielo tt_um_bleeptrack_prism_3 (.L_LO(net3));
 sg13g2_tielo tt_um_bleeptrack_prism_4 (.L_LO(net4));
 sg13g2_tielo tt_um_bleeptrack_prism_5 (.L_LO(net5));
 sg13g2_tielo tt_um_bleeptrack_prism_6 (.L_LO(net6));
 sg13g2_tielo tt_um_bleeptrack_prism_7 (.L_LO(net7));
 sg13g2_tielo tt_um_bleeptrack_prism_8 (.L_LO(net8));
 sg13g2_tielo tt_um_bleeptrack_prism_9 (.L_LO(net9));
 sg13g2_tielo tt_um_bleeptrack_prism_10 (.L_LO(net10));
 sg13g2_tielo tt_um_bleeptrack_prism_11 (.L_LO(net11));
 sg13g2_tielo tt_um_bleeptrack_prism_12 (.L_LO(net12));
 sg13g2_tielo tt_um_bleeptrack_prism_13 (.L_LO(net13));
 sg13g2_tielo tt_um_bleeptrack_prism_14 (.L_LO(net14));
 sg13g2_tielo tt_um_bleeptrack_prism_15 (.L_LO(net15));
 sg13g2_tielo tt_um_bleeptrack_prism_16 (.L_LO(net16));
 sg13g2_tiehi _839__17 (.L_HI(net17));
 sg13g2_buf_1 _898_ (.A(net43),
    .X(uo_out[3]));
 sg13g2_buf_2 _899_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout41 (.A(_323_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_323_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(\hvsync_gen.vsync ),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(net76),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(net90),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(\hvsync_gen.vpos[4] ),
    .X(net46));
 sg13g2_buf_4 fanout47 (.X(net47),
    .A(\dist_y[0] ));
 sg13g2_buf_2 fanout48 (.A(net49),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(\hvsync_gen.hpos[9] ),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(\hvsync_gen.hpos[5] ),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(\dist_x[0] ),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(rst_n),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(rst_n),
    .X(net53));
 sg13g2_tielo tt_um_bleeptrack_prism_1 (.L_LO(net1));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_024_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold2 (.A(_022_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold3 (.A(_365_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold4 (.A(_002_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold5 (.A(_070_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold6 (.A(_000_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold7 (.A(_015_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold8 (.A(_030_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold9 (.A(_011_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold10 (.A(_384_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold11 (.A(_052_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold12 (.A(_009_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold13 (.A(_014_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold14 (.A(_049_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold15 (.A(\hvsync_gen.vpos[9] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold16 (.A(_062_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold17 (.A(_001_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold18 (.A(_005_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold19 (.A(_372_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold20 (.A(_048_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold21 (.A(\hvsync_gen.vpos[1] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold22 (.A(_012_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold23 (.A(_032_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold24 (.A(\hvsync_gen.vpos[8] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold25 (.A(_010_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold26 (.A(\hvsync_gen.vpos[2] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold27 (.A(\hvsync_gen.hpos[2] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold28 (.A(\hvsync_gen.hpos[8] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold29 (.A(\hvsync_gen.vpos[5] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold30 (.A(\hvsync_gen.vpos[6] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold31 (.A(_004_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold32 (.A(_327_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold33 (.A(\hvsync_gen.hpos[4] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold34 (.A(\dist_x[0] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold35 (.A(\hvsync_gen.hpos[6] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold36 (.A(\hvsync_gen.vpos[6] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold37 (.A(_385_),
    .X(net98));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_4 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_225 ();
 sg13g2_decap_8 FILLER_16_232 ();
 sg13g2_fill_1 FILLER_16_239 ();
 sg13g2_decap_8 FILLER_16_244 ();
 sg13g2_decap_8 FILLER_16_251 ();
 sg13g2_decap_8 FILLER_16_262 ();
 sg13g2_decap_8 FILLER_16_269 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_299 ();
 sg13g2_decap_8 FILLER_17_306 ();
 sg13g2_decap_8 FILLER_17_313 ();
 sg13g2_decap_8 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_17_327 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_decap_8 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_348 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_362 ();
 sg13g2_decap_8 FILLER_17_369 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_decap_8 FILLER_17_383 ();
 sg13g2_decap_8 FILLER_17_390 ();
 sg13g2_decap_8 FILLER_17_397 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_4 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_198 ();
 sg13g2_fill_1 FILLER_18_220 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_4 FILLER_18_232 ();
 sg13g2_fill_1 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_246 ();
 sg13g2_decap_4 FILLER_18_316 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_156 ();
 sg13g2_decap_4 FILLER_19_161 ();
 sg13g2_fill_2 FILLER_19_170 ();
 sg13g2_fill_1 FILLER_19_172 ();
 sg13g2_fill_2 FILLER_19_177 ();
 sg13g2_fill_1 FILLER_19_179 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_225 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_decap_4 FILLER_19_277 ();
 sg13g2_fill_2 FILLER_19_302 ();
 sg13g2_fill_2 FILLER_19_313 ();
 sg13g2_fill_1 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_4 FILLER_19_403 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_4 FILLER_20_140 ();
 sg13g2_fill_2 FILLER_20_144 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_208 ();
 sg13g2_decap_8 FILLER_20_248 ();
 sg13g2_fill_2 FILLER_20_255 ();
 sg13g2_fill_1 FILLER_20_283 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_fill_2 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_126 ();
 sg13g2_decap_4 FILLER_21_141 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_decap_8 FILLER_21_163 ();
 sg13g2_fill_2 FILLER_21_170 ();
 sg13g2_decap_4 FILLER_21_210 ();
 sg13g2_fill_2 FILLER_21_214 ();
 sg13g2_fill_2 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_decap_8 FILLER_21_255 ();
 sg13g2_decap_4 FILLER_21_262 ();
 sg13g2_fill_2 FILLER_21_266 ();
 sg13g2_decap_4 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_281 ();
 sg13g2_fill_2 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_fill_2 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_97 ();
 sg13g2_fill_2 FILLER_22_104 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_fill_2 FILLER_22_183 ();
 sg13g2_fill_1 FILLER_22_185 ();
 sg13g2_fill_1 FILLER_22_205 ();
 sg13g2_fill_2 FILLER_22_211 ();
 sg13g2_fill_1 FILLER_22_213 ();
 sg13g2_decap_4 FILLER_22_222 ();
 sg13g2_decap_4 FILLER_22_240 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_fill_2 FILLER_22_279 ();
 sg13g2_decap_4 FILLER_22_289 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_fill_2 FILLER_22_307 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_fill_2 FILLER_22_322 ();
 sg13g2_fill_1 FILLER_22_324 ();
 sg13g2_fill_2 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_4 FILLER_23_77 ();
 sg13g2_fill_1 FILLER_23_81 ();
 sg13g2_fill_2 FILLER_23_113 ();
 sg13g2_fill_1 FILLER_23_115 ();
 sg13g2_fill_1 FILLER_23_135 ();
 sg13g2_decap_4 FILLER_23_172 ();
 sg13g2_decap_8 FILLER_23_181 ();
 sg13g2_decap_8 FILLER_23_188 ();
 sg13g2_decap_4 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_decap_4 FILLER_23_208 ();
 sg13g2_decap_8 FILLER_23_234 ();
 sg13g2_decap_4 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_259 ();
 sg13g2_decap_4 FILLER_23_274 ();
 sg13g2_fill_2 FILLER_23_278 ();
 sg13g2_decap_8 FILLER_23_297 ();
 sg13g2_decap_4 FILLER_23_304 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_330 ();
 sg13g2_fill_2 FILLER_23_340 ();
 sg13g2_fill_1 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_96 ();
 sg13g2_decap_4 FILLER_24_103 ();
 sg13g2_decap_4 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_139 ();
 sg13g2_fill_2 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_156 ();
 sg13g2_fill_2 FILLER_24_163 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_196 ();
 sg13g2_decap_4 FILLER_24_229 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_4 FILLER_24_257 ();
 sg13g2_fill_2 FILLER_24_261 ();
 sg13g2_decap_4 FILLER_24_301 ();
 sg13g2_fill_2 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_4 FILLER_25_77 ();
 sg13g2_fill_1 FILLER_25_107 ();
 sg13g2_fill_1 FILLER_25_135 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_fill_1 FILLER_25_165 ();
 sg13g2_decap_4 FILLER_25_176 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_decap_4 FILLER_25_208 ();
 sg13g2_fill_2 FILLER_25_212 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_decap_4 FILLER_25_232 ();
 sg13g2_decap_4 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_4 FILLER_25_272 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_decap_8 FILLER_25_282 ();
 sg13g2_fill_2 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_296 ();
 sg13g2_fill_2 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_310 ();
 sg13g2_fill_1 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_102 ();
 sg13g2_fill_1 FILLER_26_113 ();
 sg13g2_decap_8 FILLER_26_136 ();
 sg13g2_fill_1 FILLER_26_143 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_184 ();
 sg13g2_fill_2 FILLER_26_204 ();
 sg13g2_fill_1 FILLER_26_206 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_decap_4 FILLER_26_231 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_decap_4 FILLER_26_244 ();
 sg13g2_fill_2 FILLER_26_248 ();
 sg13g2_decap_4 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_267 ();
 sg13g2_decap_4 FILLER_26_273 ();
 sg13g2_fill_2 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_323 ();
 sg13g2_fill_2 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_fill_2 FILLER_27_156 ();
 sg13g2_fill_2 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_168 ();
 sg13g2_fill_2 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_177 ();
 sg13g2_fill_1 FILLER_27_195 ();
 sg13g2_fill_2 FILLER_27_222 ();
 sg13g2_decap_8 FILLER_27_240 ();
 sg13g2_fill_2 FILLER_27_255 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_decap_8 FILLER_27_270 ();
 sg13g2_fill_2 FILLER_27_277 ();
 sg13g2_decap_8 FILLER_27_290 ();
 sg13g2_decap_4 FILLER_27_297 ();
 sg13g2_fill_1 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_306 ();
 sg13g2_decap_8 FILLER_27_313 ();
 sg13g2_decap_4 FILLER_27_320 ();
 sg13g2_fill_2 FILLER_27_324 ();
 sg13g2_decap_8 FILLER_27_341 ();
 sg13g2_decap_8 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_108 ();
 sg13g2_decap_8 FILLER_28_115 ();
 sg13g2_fill_2 FILLER_28_122 ();
 sg13g2_fill_1 FILLER_28_124 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_decap_4 FILLER_28_171 ();
 sg13g2_decap_8 FILLER_28_179 ();
 sg13g2_fill_1 FILLER_28_190 ();
 sg13g2_decap_8 FILLER_28_199 ();
 sg13g2_decap_8 FILLER_28_206 ();
 sg13g2_fill_2 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_decap_4 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_230 ();
 sg13g2_fill_2 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_248 ();
 sg13g2_decap_4 FILLER_28_255 ();
 sg13g2_decap_4 FILLER_28_267 ();
 sg13g2_fill_2 FILLER_28_271 ();
 sg13g2_decap_8 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_286 ();
 sg13g2_fill_2 FILLER_28_318 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_decap_4 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_4 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_decap_8 FILLER_29_132 ();
 sg13g2_decap_4 FILLER_29_139 ();
 sg13g2_fill_2 FILLER_29_143 ();
 sg13g2_decap_8 FILLER_29_149 ();
 sg13g2_decap_8 FILLER_29_156 ();
 sg13g2_decap_8 FILLER_29_163 ();
 sg13g2_fill_1 FILLER_29_170 ();
 sg13g2_fill_1 FILLER_29_193 ();
 sg13g2_decap_4 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_228 ();
 sg13g2_decap_4 FILLER_29_261 ();
 sg13g2_fill_2 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_287 ();
 sg13g2_decap_4 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_fill_2 FILLER_29_342 ();
 sg13g2_fill_1 FILLER_29_344 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_156 ();
 sg13g2_fill_2 FILLER_30_163 ();
 sg13g2_decap_8 FILLER_30_180 ();
 sg13g2_decap_4 FILLER_30_187 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_fill_1 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_223 ();
 sg13g2_decap_8 FILLER_30_230 ();
 sg13g2_decap_4 FILLER_30_237 ();
 sg13g2_fill_2 FILLER_30_241 ();
 sg13g2_decap_4 FILLER_30_247 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_decap_4 FILLER_30_257 ();
 sg13g2_decap_4 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_278 ();
 sg13g2_decap_8 FILLER_30_285 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_296 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_305 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_decap_4 FILLER_30_339 ();
 sg13g2_decap_4 FILLER_30_347 ();
 sg13g2_fill_2 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_373 ();
 sg13g2_decap_8 FILLER_30_380 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_4 FILLER_31_140 ();
 sg13g2_fill_1 FILLER_31_144 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_4 FILLER_31_168 ();
 sg13g2_fill_2 FILLER_31_172 ();
 sg13g2_decap_4 FILLER_31_187 ();
 sg13g2_fill_2 FILLER_31_191 ();
 sg13g2_decap_4 FILLER_31_198 ();
 sg13g2_fill_2 FILLER_31_202 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_decap_8 FILLER_31_219 ();
 sg13g2_decap_8 FILLER_31_226 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_fill_2 FILLER_31_251 ();
 sg13g2_fill_2 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_fill_2 FILLER_31_316 ();
 sg13g2_fill_1 FILLER_31_318 ();
 sg13g2_decap_8 FILLER_31_331 ();
 sg13g2_decap_4 FILLER_31_353 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_4 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_151 ();
 sg13g2_fill_2 FILLER_32_165 ();
 sg13g2_fill_2 FILLER_32_171 ();
 sg13g2_fill_1 FILLER_32_173 ();
 sg13g2_decap_4 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_188 ();
 sg13g2_decap_8 FILLER_32_195 ();
 sg13g2_fill_2 FILLER_32_202 ();
 sg13g2_fill_1 FILLER_32_204 ();
 sg13g2_decap_4 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_253 ();
 sg13g2_decap_8 FILLER_32_260 ();
 sg13g2_fill_1 FILLER_32_267 ();
 sg13g2_fill_2 FILLER_32_288 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_decap_8 FILLER_32_299 ();
 sg13g2_decap_4 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_310 ();
 sg13g2_decap_4 FILLER_32_328 ();
 sg13g2_fill_2 FILLER_32_332 ();
 sg13g2_decap_8 FILLER_32_342 ();
 sg13g2_decap_8 FILLER_32_349 ();
 sg13g2_fill_2 FILLER_32_356 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_363 ();
 sg13g2_decap_8 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_32_377 ();
 sg13g2_decap_8 FILLER_32_384 ();
 sg13g2_decap_8 FILLER_32_391 ();
 sg13g2_decap_8 FILLER_32_398 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_4 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_156 ();
 sg13g2_fill_2 FILLER_33_160 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_fill_2 FILLER_33_171 ();
 sg13g2_decap_4 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_fill_1 FILLER_33_216 ();
 sg13g2_decap_8 FILLER_33_227 ();
 sg13g2_decap_4 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_decap_4 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_decap_8 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_fill_2 FILLER_33_284 ();
 sg13g2_decap_4 FILLER_33_290 ();
 sg13g2_fill_2 FILLER_33_294 ();
 sg13g2_fill_2 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_326 ();
 sg13g2_fill_1 FILLER_33_333 ();
 sg13g2_decap_4 FILLER_33_344 ();
 sg13g2_decap_8 FILLER_33_374 ();
 sg13g2_decap_8 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_388 ();
 sg13g2_decap_8 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_fill_1 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_145 ();
 sg13g2_decap_4 FILLER_34_152 ();
 sg13g2_fill_2 FILLER_34_156 ();
 sg13g2_decap_8 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_174 ();
 sg13g2_decap_8 FILLER_34_180 ();
 sg13g2_decap_8 FILLER_34_187 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_decap_4 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_230 ();
 sg13g2_fill_2 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_269 ();
 sg13g2_decap_8 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_decap_8 FILLER_34_305 ();
 sg13g2_fill_2 FILLER_34_312 ();
 sg13g2_decap_8 FILLER_34_318 ();
 sg13g2_fill_2 FILLER_34_325 ();
 sg13g2_decap_4 FILLER_34_336 ();
 sg13g2_fill_1 FILLER_34_340 ();
 sg13g2_decap_4 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_367 ();
 sg13g2_decap_8 FILLER_34_374 ();
 sg13g2_decap_8 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_34_388 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_fill_1 FILLER_35_154 ();
 sg13g2_fill_1 FILLER_35_188 ();
 sg13g2_decap_8 FILLER_35_202 ();
 sg13g2_decap_8 FILLER_35_209 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_decap_4 FILLER_35_230 ();
 sg13g2_decap_4 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_279 ();
 sg13g2_fill_2 FILLER_35_288 ();
 sg13g2_fill_1 FILLER_35_290 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_326 ();
 sg13g2_fill_1 FILLER_35_328 ();
 sg13g2_fill_2 FILLER_35_335 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_141 ();
 sg13g2_decap_8 FILLER_36_148 ();
 sg13g2_decap_8 FILLER_36_155 ();
 sg13g2_fill_1 FILLER_36_162 ();
 sg13g2_decap_4 FILLER_36_171 ();
 sg13g2_fill_2 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_196 ();
 sg13g2_decap_4 FILLER_36_214 ();
 sg13g2_fill_1 FILLER_36_218 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_fill_1 FILLER_36_233 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_276 ();
 sg13g2_decap_4 FILLER_36_283 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_299 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_4 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_138 ();
 sg13g2_fill_1 FILLER_37_145 ();
 sg13g2_fill_1 FILLER_37_179 ();
 sg13g2_decap_8 FILLER_37_206 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_219 ();
 sg13g2_fill_1 FILLER_37_221 ();
 sg13g2_decap_8 FILLER_37_328 ();
 sg13g2_decap_8 FILLER_37_335 ();
 sg13g2_decap_8 FILLER_37_342 ();
 sg13g2_decap_8 FILLER_37_349 ();
 sg13g2_decap_8 FILLER_37_356 ();
 sg13g2_decap_8 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_370 ();
 sg13g2_decap_8 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_37_384 ();
 sg13g2_decap_8 FILLER_37_391 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_168 ();
 sg13g2_fill_1 FILLER_38_177 ();
 sg13g2_decap_4 FILLER_38_187 ();
 sg13g2_fill_1 FILLER_38_195 ();
 sg13g2_decap_8 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_decap_4 FILLER_38_227 ();
 sg13g2_fill_2 FILLER_38_231 ();
 sg13g2_decap_4 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_decap_8 FILLER_38_248 ();
 sg13g2_decap_8 FILLER_38_255 ();
 sg13g2_decap_4 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_4 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_286 ();
 sg13g2_decap_8 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_300 ();
 sg13g2_decap_4 FILLER_38_307 ();
 sg13g2_fill_2 FILLER_38_311 ();
 sg13g2_decap_8 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_324 ();
 sg13g2_decap_8 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_352 ();
 sg13g2_decap_8 FILLER_38_359 ();
 sg13g2_decap_8 FILLER_38_366 ();
 sg13g2_decap_8 FILLER_38_373 ();
 sg13g2_decap_8 FILLER_38_380 ();
 sg13g2_decap_8 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_394 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
endmodule
