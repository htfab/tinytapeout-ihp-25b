module tt_um_dumbrv_yliu_hashed (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire clk_regs;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire \core.e2m_addr[0] ;
 wire \core.e2m_addr[10] ;
 wire \core.e2m_addr[11] ;
 wire \core.e2m_addr[12] ;
 wire \core.e2m_addr[13] ;
 wire \core.e2m_addr[14] ;
 wire \core.e2m_addr[15] ;
 wire \core.e2m_addr[16] ;
 wire \core.e2m_addr[17] ;
 wire \core.e2m_addr[18] ;
 wire \core.e2m_addr[19] ;
 wire \core.e2m_addr[1] ;
 wire \core.e2m_addr[20] ;
 wire \core.e2m_addr[21] ;
 wire \core.e2m_addr[22] ;
 wire \core.e2m_addr[23] ;
 wire \core.e2m_addr[24] ;
 wire \core.e2m_addr[25] ;
 wire \core.e2m_addr[26] ;
 wire \core.e2m_addr[27] ;
 wire \core.e2m_addr[28] ;
 wire \core.e2m_addr[29] ;
 wire \core.e2m_addr[2] ;
 wire \core.e2m_addr[30] ;
 wire \core.e2m_addr[31] ;
 wire \core.e2m_addr[3] ;
 wire \core.e2m_addr[4] ;
 wire \core.e2m_addr[5] ;
 wire \core.e2m_addr[6] ;
 wire \core.e2m_addr[7] ;
 wire \core.e2m_addr[8] ;
 wire \core.e2m_addr[9] ;
 wire \core.e2m_data[0] ;
 wire \core.e2m_data[10] ;
 wire \core.e2m_data[11] ;
 wire \core.e2m_data[12] ;
 wire \core.e2m_data[13] ;
 wire \core.e2m_data[14] ;
 wire \core.e2m_data[15] ;
 wire \core.e2m_data[16] ;
 wire \core.e2m_data[17] ;
 wire \core.e2m_data[18] ;
 wire \core.e2m_data[19] ;
 wire \core.e2m_data[1] ;
 wire \core.e2m_data[20] ;
 wire \core.e2m_data[21] ;
 wire \core.e2m_data[22] ;
 wire \core.e2m_data[23] ;
 wire \core.e2m_data[24] ;
 wire \core.e2m_data[25] ;
 wire \core.e2m_data[26] ;
 wire \core.e2m_data[27] ;
 wire \core.e2m_data[28] ;
 wire \core.e2m_data[29] ;
 wire \core.e2m_data[2] ;
 wire \core.e2m_data[30] ;
 wire \core.e2m_data[31] ;
 wire \core.e2m_data[3] ;
 wire \core.e2m_data[4] ;
 wire \core.e2m_data[5] ;
 wire \core.e2m_data[6] ;
 wire \core.e2m_data[7] ;
 wire \core.e2m_data[8] ;
 wire \core.e2m_data[9] ;
 wire \core.f2e_addr[10] ;
 wire \core.f2e_addr[11] ;
 wire \core.f2e_addr[12] ;
 wire \core.f2e_addr[13] ;
 wire \core.f2e_addr[14] ;
 wire \core.f2e_addr[15] ;
 wire \core.f2e_addr[1] ;
 wire \core.f2e_addr[2] ;
 wire \core.f2e_addr[3] ;
 wire \core.f2e_addr[4] ;
 wire \core.f2e_addr[5] ;
 wire \core.f2e_addr[6] ;
 wire \core.f2e_addr[7] ;
 wire \core.f2e_addr[8] ;
 wire \core.f2e_addr[9] ;
 wire \core.f2e_inst[0] ;
 wire \core.f2e_inst[10] ;
 wire \core.f2e_inst[11] ;
 wire \core.f2e_inst[12] ;
 wire \core.f2e_inst[13] ;
 wire \core.f2e_inst[14] ;
 wire \core.f2e_inst[15] ;
 wire \core.f2e_inst[16] ;
 wire \core.f2e_inst[17] ;
 wire \core.f2e_inst[18] ;
 wire \core.f2e_inst[19] ;
 wire \core.f2e_inst[1] ;
 wire \core.f2e_inst[20] ;
 wire \core.f2e_inst[21] ;
 wire \core.f2e_inst[22] ;
 wire \core.f2e_inst[23] ;
 wire \core.f2e_inst[24] ;
 wire \core.f2e_inst[25] ;
 wire \core.f2e_inst[26] ;
 wire \core.f2e_inst[27] ;
 wire \core.f2e_inst[28] ;
 wire \core.f2e_inst[29] ;
 wire \core.f2e_inst[2] ;
 wire \core.f2e_inst[30] ;
 wire \core.f2e_inst[31] ;
 wire \core.f2e_inst[3] ;
 wire \core.f2e_inst[4] ;
 wire \core.f2e_inst[5] ;
 wire \core.f2e_inst[6] ;
 wire \core.f2e_inst[7] ;
 wire \core.f2e_inst[8] ;
 wire \core.f2e_inst[9] ;
 wire \core.fetch.cmd_data[0] ;
 wire \core.fetch.cmd_data[1] ;
 wire \core.fetch.cmd_data[2] ;
 wire \core.fetch.cmd_data[3] ;
 wire \core.fetch.cmd_data[4] ;
 wire \core.fetch.cmd_data[5] ;
 wire \core.fetch.cmd_data[6] ;
 wire \core.fetch.cmd_data[7] ;
 wire \core.fetch.cmd_valid ;
 wire \core.fetch.data[0] ;
 wire \core.fetch.data[10] ;
 wire \core.fetch.data[11] ;
 wire \core.fetch.data[12] ;
 wire \core.fetch.data[13] ;
 wire \core.fetch.data[14] ;
 wire \core.fetch.data[15] ;
 wire \core.fetch.data[16] ;
 wire \core.fetch.data[17] ;
 wire \core.fetch.data[18] ;
 wire \core.fetch.data[19] ;
 wire \core.fetch.data[1] ;
 wire \core.fetch.data[20] ;
 wire \core.fetch.data[21] ;
 wire \core.fetch.data[22] ;
 wire \core.fetch.data[23] ;
 wire \core.fetch.data[24] ;
 wire \core.fetch.data[25] ;
 wire \core.fetch.data[26] ;
 wire \core.fetch.data[27] ;
 wire \core.fetch.data[28] ;
 wire \core.fetch.data[29] ;
 wire \core.fetch.data[2] ;
 wire \core.fetch.data[30] ;
 wire \core.fetch.data[31] ;
 wire \core.fetch.data[3] ;
 wire \core.fetch.data[4] ;
 wire \core.fetch.data[5] ;
 wire \core.fetch.data[6] ;
 wire \core.fetch.data[7] ;
 wire \core.fetch.data[8] ;
 wire \core.fetch.data[9] ;
 wire \core.fetch.data_size[0] ;
 wire \core.fetch.data_size[1] ;
 wire \core.fetch.data_size[2] ;
 wire \core.fetch.inst[32] ;
 wire \core.fetch.inst[33] ;
 wire \core.fetch.inst[34] ;
 wire \core.fetch.inst[35] ;
 wire \core.fetch.inst[36] ;
 wire \core.fetch.inst[37] ;
 wire \core.fetch.inst[38] ;
 wire \core.fetch.inst[39] ;
 wire \core.fetch.inst[40] ;
 wire \core.fetch.inst[41] ;
 wire \core.fetch.inst[42] ;
 wire \core.fetch.inst[43] ;
 wire \core.fetch.inst[44] ;
 wire \core.fetch.inst[45] ;
 wire \core.fetch.inst[46] ;
 wire \core.fetch.inst[47] ;
 wire \core.fetch.inst_size[0] ;
 wire \core.fetch.inst_size[1] ;
 wire \core.fetch.inst_size[2] ;
 wire \core.fetch.rd_addr_i[0] ;
 wire \core.fetch.rd_addr_i[10] ;
 wire \core.fetch.rd_addr_i[11] ;
 wire \core.fetch.rd_addr_i[12] ;
 wire \core.fetch.rd_addr_i[13] ;
 wire \core.fetch.rd_addr_i[14] ;
 wire \core.fetch.rd_addr_i[15] ;
 wire \core.fetch.rd_addr_i[1] ;
 wire \core.fetch.rd_addr_i[2] ;
 wire \core.fetch.rd_addr_i[3] ;
 wire \core.fetch.rd_addr_i[4] ;
 wire \core.fetch.rd_addr_i[5] ;
 wire \core.fetch.rd_addr_i[6] ;
 wire \core.fetch.rd_addr_i[7] ;
 wire \core.fetch.rd_addr_i[8] ;
 wire \core.fetch.rd_addr_i[9] ;
 wire \core.fetch.spi_reader.addr[0] ;
 wire \core.fetch.spi_reader.addr[10] ;
 wire \core.fetch.spi_reader.addr[11] ;
 wire \core.fetch.spi_reader.addr[12] ;
 wire \core.fetch.spi_reader.addr[13] ;
 wire \core.fetch.spi_reader.addr[14] ;
 wire \core.fetch.spi_reader.addr[15] ;
 wire \core.fetch.spi_reader.addr[1] ;
 wire \core.fetch.spi_reader.addr[2] ;
 wire \core.fetch.spi_reader.addr[3] ;
 wire \core.fetch.spi_reader.addr[4] ;
 wire \core.fetch.spi_reader.addr[5] ;
 wire \core.fetch.spi_reader.addr[6] ;
 wire \core.fetch.spi_reader.addr[7] ;
 wire \core.fetch.spi_reader.addr[8] ;
 wire \core.fetch.spi_reader.addr[9] ;
 wire \core.fetch.spi_reader.cache_bit ;
 wire \core.fetch.spi_reader.counter[0] ;
 wire \core.fetch.spi_reader.counter[1] ;
 wire \core.fetch.spi_reader.counter[2] ;
 wire \core.fetch.spi_reader.counter[3] ;
 wire \core.fetch.spi_reader.counter[4] ;
 wire \core.fetch.spi_reader.counter[5] ;
 wire \core.fetch.spi_reader.cs ;
 wire \core.fetch.spi_reader.dirty ;
 wire \core.fetch.spi_reader.sck ;
 wire \core.fetch.spi_reader.state[0] ;
 wire \core.fetch.spi_reader.state[1] ;
 wire \core.fetch.spi_reader.state[2] ;
 wire \core.fetch.state[0] ;
 wire \core.fetch.state[1] ;
 wire \core.gpio.stray_data_i[0] ;
 wire \core.gpio.stray_data_i[10] ;
 wire \core.gpio.stray_data_i[11] ;
 wire \core.gpio.stray_data_i[12] ;
 wire \core.gpio.stray_data_i[13] ;
 wire \core.gpio.stray_data_i[14] ;
 wire \core.gpio.stray_data_i[15] ;
 wire \core.gpio.stray_data_i[16] ;
 wire \core.gpio.stray_data_i[17] ;
 wire \core.gpio.stray_data_i[18] ;
 wire \core.gpio.stray_data_i[19] ;
 wire \core.gpio.stray_data_i[1] ;
 wire \core.gpio.stray_data_i[20] ;
 wire \core.gpio.stray_data_i[21] ;
 wire \core.gpio.stray_data_i[22] ;
 wire \core.gpio.stray_data_i[23] ;
 wire \core.gpio.stray_data_i[24] ;
 wire \core.gpio.stray_data_i[25] ;
 wire \core.gpio.stray_data_i[26] ;
 wire \core.gpio.stray_data_i[27] ;
 wire \core.gpio.stray_data_i[28] ;
 wire \core.gpio.stray_data_i[29] ;
 wire \core.gpio.stray_data_i[2] ;
 wire \core.gpio.stray_data_i[30] ;
 wire \core.gpio.stray_data_i[31] ;
 wire \core.gpio.stray_data_i[3] ;
 wire \core.gpio.stray_data_i[4] ;
 wire \core.gpio.stray_data_i[5] ;
 wire \core.gpio.stray_data_i[6] ;
 wire \core.gpio.stray_data_i[7] ;
 wire \core.gpio.stray_data_i[8] ;
 wire \core.gpio.stray_data_i[9] ;
 wire \core.gpio.stray_wr_i ;
 wire \core.lsu.accept ;
 wire \core.lsu.dreg[0] ;
 wire \core.lsu.dreg[1] ;
 wire \core.lsu.dreg[2] ;
 wire \core.lsu.dreg[3] ;
 wire \core.lsu.is_byte ;
 wire \core.lsu.is_half ;
 wire \core.lsu.is_signed ;
 wire \core.lsu.spi.addr[0] ;
 wire \core.lsu.spi.addr[10] ;
 wire \core.lsu.spi.addr[11] ;
 wire \core.lsu.spi.addr[12] ;
 wire \core.lsu.spi.addr[13] ;
 wire \core.lsu.spi.addr[14] ;
 wire \core.lsu.spi.addr[15] ;
 wire \core.lsu.spi.addr[1] ;
 wire \core.lsu.spi.addr[2] ;
 wire \core.lsu.spi.addr[3] ;
 wire \core.lsu.spi.addr[4] ;
 wire \core.lsu.spi.addr[5] ;
 wire \core.lsu.spi.addr[6] ;
 wire \core.lsu.spi.addr[7] ;
 wire \core.lsu.spi.addr[8] ;
 wire \core.lsu.spi.addr[9] ;
 wire \core.lsu.spi.buffer[0] ;
 wire \core.lsu.spi.buffer[1] ;
 wire \core.lsu.spi.buffer[2] ;
 wire \core.lsu.spi.buffer[3] ;
 wire \core.lsu.spi.buffer[4] ;
 wire \core.lsu.spi.buffer[5] ;
 wire \core.lsu.spi.buffer[6] ;
 wire \core.lsu.spi.buffer[7] ;
 wire \core.lsu.spi.cache_bit ;
 wire \core.lsu.spi.counter[0] ;
 wire \core.lsu.spi.counter[1] ;
 wire \core.lsu.spi.counter[2] ;
 wire \core.lsu.spi.counter[3] ;
 wire \core.lsu.spi.counter[4] ;
 wire \core.lsu.spi.counter[5] ;
 wire \core.lsu.spi.cs ;
 wire \core.lsu.spi.dirty ;
 wire \core.lsu.spi.iswr ;
 wire \core.lsu.spi.sck ;
 wire \core.lsu.spi.state[0] ;
 wire \core.lsu.spi.state[1] ;
 wire \core.lsu.spi.state[2] ;
 wire \core.lsu.spi_valid ;
 wire \core.lsu.state[0] ;
 wire \core.lsu.state[1] ;
 wire \core.lsu.state[2] ;
 wire \core.lsu.write_index[0] ;
 wire \core.lsu.write_index[1] ;
 wire \core.lsu.write_index[2] ;
 wire \core.work.alu.is_mem ;
 wire \core.work.alu.is_sign ;
 wire \core.work.alu.is_wr ;
 wire \core.work.alu.ls_size_b ;
 wire \core.work.alu.ls_size_h ;
 wire \core.work.alu.sval2[0] ;
 wire \core.work.alu.sval2[10] ;
 wire \core.work.alu.sval2[11] ;
 wire \core.work.alu.sval2[12] ;
 wire \core.work.alu.sval2[13] ;
 wire \core.work.alu.sval2[14] ;
 wire \core.work.alu.sval2[15] ;
 wire \core.work.alu.sval2[16] ;
 wire \core.work.alu.sval2[17] ;
 wire \core.work.alu.sval2[18] ;
 wire \core.work.alu.sval2[19] ;
 wire \core.work.alu.sval2[1] ;
 wire \core.work.alu.sval2[20] ;
 wire \core.work.alu.sval2[21] ;
 wire \core.work.alu.sval2[22] ;
 wire \core.work.alu.sval2[23] ;
 wire \core.work.alu.sval2[24] ;
 wire \core.work.alu.sval2[25] ;
 wire \core.work.alu.sval2[26] ;
 wire \core.work.alu.sval2[27] ;
 wire \core.work.alu.sval2[28] ;
 wire \core.work.alu.sval2[29] ;
 wire \core.work.alu.sval2[2] ;
 wire \core.work.alu.sval2[30] ;
 wire \core.work.alu.sval2[31] ;
 wire \core.work.alu.sval2[3] ;
 wire \core.work.alu.sval2[4] ;
 wire \core.work.alu.sval2[5] ;
 wire \core.work.alu.sval2[6] ;
 wire \core.work.alu.sval2[7] ;
 wire \core.work.alu.sval2[8] ;
 wire \core.work.alu.sval2[9] ;
 wire \core.work.dreg[0] ;
 wire \core.work.dreg[1] ;
 wire \core.work.dreg[2] ;
 wire \core.work.dreg[3] ;
 wire \core.work.inst_was_short ;
 wire \core.work.op[4] ;
 wire \core.work.registers.genblk1[10].latch[0] ;
 wire \core.work.registers.genblk1[10].latch[10] ;
 wire \core.work.registers.genblk1[10].latch[11] ;
 wire \core.work.registers.genblk1[10].latch[12] ;
 wire \core.work.registers.genblk1[10].latch[13] ;
 wire \core.work.registers.genblk1[10].latch[14] ;
 wire \core.work.registers.genblk1[10].latch[15] ;
 wire \core.work.registers.genblk1[10].latch[16] ;
 wire \core.work.registers.genblk1[10].latch[17] ;
 wire \core.work.registers.genblk1[10].latch[18] ;
 wire \core.work.registers.genblk1[10].latch[19] ;
 wire \core.work.registers.genblk1[10].latch[1] ;
 wire \core.work.registers.genblk1[10].latch[20] ;
 wire \core.work.registers.genblk1[10].latch[21] ;
 wire \core.work.registers.genblk1[10].latch[22] ;
 wire \core.work.registers.genblk1[10].latch[23] ;
 wire \core.work.registers.genblk1[10].latch[24] ;
 wire \core.work.registers.genblk1[10].latch[25] ;
 wire \core.work.registers.genblk1[10].latch[26] ;
 wire \core.work.registers.genblk1[10].latch[27] ;
 wire \core.work.registers.genblk1[10].latch[28] ;
 wire \core.work.registers.genblk1[10].latch[29] ;
 wire \core.work.registers.genblk1[10].latch[2] ;
 wire \core.work.registers.genblk1[10].latch[30] ;
 wire \core.work.registers.genblk1[10].latch[31] ;
 wire \core.work.registers.genblk1[10].latch[3] ;
 wire \core.work.registers.genblk1[10].latch[4] ;
 wire \core.work.registers.genblk1[10].latch[5] ;
 wire \core.work.registers.genblk1[10].latch[6] ;
 wire \core.work.registers.genblk1[10].latch[7] ;
 wire \core.work.registers.genblk1[10].latch[8] ;
 wire \core.work.registers.genblk1[10].latch[9] ;
 wire \core.work.registers.genblk1[10].we ;
 wire \core.work.registers.genblk1[11].latch[0] ;
 wire \core.work.registers.genblk1[11].latch[10] ;
 wire \core.work.registers.genblk1[11].latch[11] ;
 wire \core.work.registers.genblk1[11].latch[12] ;
 wire \core.work.registers.genblk1[11].latch[13] ;
 wire \core.work.registers.genblk1[11].latch[14] ;
 wire \core.work.registers.genblk1[11].latch[15] ;
 wire \core.work.registers.genblk1[11].latch[16] ;
 wire \core.work.registers.genblk1[11].latch[17] ;
 wire \core.work.registers.genblk1[11].latch[18] ;
 wire \core.work.registers.genblk1[11].latch[19] ;
 wire \core.work.registers.genblk1[11].latch[1] ;
 wire \core.work.registers.genblk1[11].latch[20] ;
 wire \core.work.registers.genblk1[11].latch[21] ;
 wire \core.work.registers.genblk1[11].latch[22] ;
 wire \core.work.registers.genblk1[11].latch[23] ;
 wire \core.work.registers.genblk1[11].latch[24] ;
 wire \core.work.registers.genblk1[11].latch[25] ;
 wire \core.work.registers.genblk1[11].latch[26] ;
 wire \core.work.registers.genblk1[11].latch[27] ;
 wire \core.work.registers.genblk1[11].latch[28] ;
 wire \core.work.registers.genblk1[11].latch[29] ;
 wire \core.work.registers.genblk1[11].latch[2] ;
 wire \core.work.registers.genblk1[11].latch[30] ;
 wire \core.work.registers.genblk1[11].latch[31] ;
 wire \core.work.registers.genblk1[11].latch[3] ;
 wire \core.work.registers.genblk1[11].latch[4] ;
 wire \core.work.registers.genblk1[11].latch[5] ;
 wire \core.work.registers.genblk1[11].latch[6] ;
 wire \core.work.registers.genblk1[11].latch[7] ;
 wire \core.work.registers.genblk1[11].latch[8] ;
 wire \core.work.registers.genblk1[11].latch[9] ;
 wire \core.work.registers.genblk1[11].we ;
 wire \core.work.registers.genblk1[12].latch[0] ;
 wire \core.work.registers.genblk1[12].latch[10] ;
 wire \core.work.registers.genblk1[12].latch[11] ;
 wire \core.work.registers.genblk1[12].latch[12] ;
 wire \core.work.registers.genblk1[12].latch[13] ;
 wire \core.work.registers.genblk1[12].latch[14] ;
 wire \core.work.registers.genblk1[12].latch[15] ;
 wire \core.work.registers.genblk1[12].latch[16] ;
 wire \core.work.registers.genblk1[12].latch[17] ;
 wire \core.work.registers.genblk1[12].latch[18] ;
 wire \core.work.registers.genblk1[12].latch[19] ;
 wire \core.work.registers.genblk1[12].latch[1] ;
 wire \core.work.registers.genblk1[12].latch[20] ;
 wire \core.work.registers.genblk1[12].latch[21] ;
 wire \core.work.registers.genblk1[12].latch[22] ;
 wire \core.work.registers.genblk1[12].latch[23] ;
 wire \core.work.registers.genblk1[12].latch[24] ;
 wire \core.work.registers.genblk1[12].latch[25] ;
 wire \core.work.registers.genblk1[12].latch[26] ;
 wire \core.work.registers.genblk1[12].latch[27] ;
 wire \core.work.registers.genblk1[12].latch[28] ;
 wire \core.work.registers.genblk1[12].latch[29] ;
 wire \core.work.registers.genblk1[12].latch[2] ;
 wire \core.work.registers.genblk1[12].latch[30] ;
 wire \core.work.registers.genblk1[12].latch[31] ;
 wire \core.work.registers.genblk1[12].latch[3] ;
 wire \core.work.registers.genblk1[12].latch[4] ;
 wire \core.work.registers.genblk1[12].latch[5] ;
 wire \core.work.registers.genblk1[12].latch[6] ;
 wire \core.work.registers.genblk1[12].latch[7] ;
 wire \core.work.registers.genblk1[12].latch[8] ;
 wire \core.work.registers.genblk1[12].latch[9] ;
 wire \core.work.registers.genblk1[12].we ;
 wire \core.work.registers.genblk1[13].latch[0] ;
 wire \core.work.registers.genblk1[13].latch[10] ;
 wire \core.work.registers.genblk1[13].latch[11] ;
 wire \core.work.registers.genblk1[13].latch[12] ;
 wire \core.work.registers.genblk1[13].latch[13] ;
 wire \core.work.registers.genblk1[13].latch[14] ;
 wire \core.work.registers.genblk1[13].latch[15] ;
 wire \core.work.registers.genblk1[13].latch[16] ;
 wire \core.work.registers.genblk1[13].latch[17] ;
 wire \core.work.registers.genblk1[13].latch[18] ;
 wire \core.work.registers.genblk1[13].latch[19] ;
 wire \core.work.registers.genblk1[13].latch[1] ;
 wire \core.work.registers.genblk1[13].latch[20] ;
 wire \core.work.registers.genblk1[13].latch[21] ;
 wire \core.work.registers.genblk1[13].latch[22] ;
 wire \core.work.registers.genblk1[13].latch[23] ;
 wire \core.work.registers.genblk1[13].latch[24] ;
 wire \core.work.registers.genblk1[13].latch[25] ;
 wire \core.work.registers.genblk1[13].latch[26] ;
 wire \core.work.registers.genblk1[13].latch[27] ;
 wire \core.work.registers.genblk1[13].latch[28] ;
 wire \core.work.registers.genblk1[13].latch[29] ;
 wire \core.work.registers.genblk1[13].latch[2] ;
 wire \core.work.registers.genblk1[13].latch[30] ;
 wire \core.work.registers.genblk1[13].latch[31] ;
 wire \core.work.registers.genblk1[13].latch[3] ;
 wire \core.work.registers.genblk1[13].latch[4] ;
 wire \core.work.registers.genblk1[13].latch[5] ;
 wire \core.work.registers.genblk1[13].latch[6] ;
 wire \core.work.registers.genblk1[13].latch[7] ;
 wire \core.work.registers.genblk1[13].latch[8] ;
 wire \core.work.registers.genblk1[13].latch[9] ;
 wire \core.work.registers.genblk1[13].we ;
 wire \core.work.registers.genblk1[14].latch[0] ;
 wire \core.work.registers.genblk1[14].latch[10] ;
 wire \core.work.registers.genblk1[14].latch[11] ;
 wire \core.work.registers.genblk1[14].latch[12] ;
 wire \core.work.registers.genblk1[14].latch[13] ;
 wire \core.work.registers.genblk1[14].latch[14] ;
 wire \core.work.registers.genblk1[14].latch[15] ;
 wire \core.work.registers.genblk1[14].latch[16] ;
 wire \core.work.registers.genblk1[14].latch[17] ;
 wire \core.work.registers.genblk1[14].latch[18] ;
 wire \core.work.registers.genblk1[14].latch[19] ;
 wire \core.work.registers.genblk1[14].latch[1] ;
 wire \core.work.registers.genblk1[14].latch[20] ;
 wire \core.work.registers.genblk1[14].latch[21] ;
 wire \core.work.registers.genblk1[14].latch[22] ;
 wire \core.work.registers.genblk1[14].latch[23] ;
 wire \core.work.registers.genblk1[14].latch[24] ;
 wire \core.work.registers.genblk1[14].latch[25] ;
 wire \core.work.registers.genblk1[14].latch[26] ;
 wire \core.work.registers.genblk1[14].latch[27] ;
 wire \core.work.registers.genblk1[14].latch[28] ;
 wire \core.work.registers.genblk1[14].latch[29] ;
 wire \core.work.registers.genblk1[14].latch[2] ;
 wire \core.work.registers.genblk1[14].latch[30] ;
 wire \core.work.registers.genblk1[14].latch[31] ;
 wire \core.work.registers.genblk1[14].latch[3] ;
 wire \core.work.registers.genblk1[14].latch[4] ;
 wire \core.work.registers.genblk1[14].latch[5] ;
 wire \core.work.registers.genblk1[14].latch[6] ;
 wire \core.work.registers.genblk1[14].latch[7] ;
 wire \core.work.registers.genblk1[14].latch[8] ;
 wire \core.work.registers.genblk1[14].latch[9] ;
 wire \core.work.registers.genblk1[14].we ;
 wire \core.work.registers.genblk1[15].latch[0] ;
 wire \core.work.registers.genblk1[15].latch[10] ;
 wire \core.work.registers.genblk1[15].latch[11] ;
 wire \core.work.registers.genblk1[15].latch[12] ;
 wire \core.work.registers.genblk1[15].latch[13] ;
 wire \core.work.registers.genblk1[15].latch[14] ;
 wire \core.work.registers.genblk1[15].latch[15] ;
 wire \core.work.registers.genblk1[15].latch[16] ;
 wire \core.work.registers.genblk1[15].latch[17] ;
 wire \core.work.registers.genblk1[15].latch[18] ;
 wire \core.work.registers.genblk1[15].latch[19] ;
 wire \core.work.registers.genblk1[15].latch[1] ;
 wire \core.work.registers.genblk1[15].latch[20] ;
 wire \core.work.registers.genblk1[15].latch[21] ;
 wire \core.work.registers.genblk1[15].latch[22] ;
 wire \core.work.registers.genblk1[15].latch[23] ;
 wire \core.work.registers.genblk1[15].latch[24] ;
 wire \core.work.registers.genblk1[15].latch[25] ;
 wire \core.work.registers.genblk1[15].latch[26] ;
 wire \core.work.registers.genblk1[15].latch[27] ;
 wire \core.work.registers.genblk1[15].latch[28] ;
 wire \core.work.registers.genblk1[15].latch[29] ;
 wire \core.work.registers.genblk1[15].latch[2] ;
 wire \core.work.registers.genblk1[15].latch[30] ;
 wire \core.work.registers.genblk1[15].latch[31] ;
 wire \core.work.registers.genblk1[15].latch[3] ;
 wire \core.work.registers.genblk1[15].latch[4] ;
 wire \core.work.registers.genblk1[15].latch[5] ;
 wire \core.work.registers.genblk1[15].latch[6] ;
 wire \core.work.registers.genblk1[15].latch[7] ;
 wire \core.work.registers.genblk1[15].latch[8] ;
 wire \core.work.registers.genblk1[15].latch[9] ;
 wire \core.work.registers.genblk1[15].we ;
 wire \core.work.registers.genblk1[1].latch[0] ;
 wire \core.work.registers.genblk1[1].latch[10] ;
 wire \core.work.registers.genblk1[1].latch[11] ;
 wire \core.work.registers.genblk1[1].latch[12] ;
 wire \core.work.registers.genblk1[1].latch[13] ;
 wire \core.work.registers.genblk1[1].latch[14] ;
 wire \core.work.registers.genblk1[1].latch[15] ;
 wire \core.work.registers.genblk1[1].latch[16] ;
 wire \core.work.registers.genblk1[1].latch[17] ;
 wire \core.work.registers.genblk1[1].latch[18] ;
 wire \core.work.registers.genblk1[1].latch[19] ;
 wire \core.work.registers.genblk1[1].latch[1] ;
 wire \core.work.registers.genblk1[1].latch[20] ;
 wire \core.work.registers.genblk1[1].latch[21] ;
 wire \core.work.registers.genblk1[1].latch[22] ;
 wire \core.work.registers.genblk1[1].latch[23] ;
 wire \core.work.registers.genblk1[1].latch[24] ;
 wire \core.work.registers.genblk1[1].latch[25] ;
 wire \core.work.registers.genblk1[1].latch[26] ;
 wire \core.work.registers.genblk1[1].latch[27] ;
 wire \core.work.registers.genblk1[1].latch[28] ;
 wire \core.work.registers.genblk1[1].latch[29] ;
 wire \core.work.registers.genblk1[1].latch[2] ;
 wire \core.work.registers.genblk1[1].latch[30] ;
 wire \core.work.registers.genblk1[1].latch[31] ;
 wire \core.work.registers.genblk1[1].latch[3] ;
 wire \core.work.registers.genblk1[1].latch[4] ;
 wire \core.work.registers.genblk1[1].latch[5] ;
 wire \core.work.registers.genblk1[1].latch[6] ;
 wire \core.work.registers.genblk1[1].latch[7] ;
 wire \core.work.registers.genblk1[1].latch[8] ;
 wire \core.work.registers.genblk1[1].latch[9] ;
 wire \core.work.registers.genblk1[1].we ;
 wire \core.work.registers.genblk1[2].latch[0] ;
 wire \core.work.registers.genblk1[2].latch[10] ;
 wire \core.work.registers.genblk1[2].latch[11] ;
 wire \core.work.registers.genblk1[2].latch[12] ;
 wire \core.work.registers.genblk1[2].latch[13] ;
 wire \core.work.registers.genblk1[2].latch[14] ;
 wire \core.work.registers.genblk1[2].latch[15] ;
 wire \core.work.registers.genblk1[2].latch[16] ;
 wire \core.work.registers.genblk1[2].latch[17] ;
 wire \core.work.registers.genblk1[2].latch[18] ;
 wire \core.work.registers.genblk1[2].latch[19] ;
 wire \core.work.registers.genblk1[2].latch[1] ;
 wire \core.work.registers.genblk1[2].latch[20] ;
 wire \core.work.registers.genblk1[2].latch[21] ;
 wire \core.work.registers.genblk1[2].latch[22] ;
 wire \core.work.registers.genblk1[2].latch[23] ;
 wire \core.work.registers.genblk1[2].latch[24] ;
 wire \core.work.registers.genblk1[2].latch[25] ;
 wire \core.work.registers.genblk1[2].latch[26] ;
 wire \core.work.registers.genblk1[2].latch[27] ;
 wire \core.work.registers.genblk1[2].latch[28] ;
 wire \core.work.registers.genblk1[2].latch[29] ;
 wire \core.work.registers.genblk1[2].latch[2] ;
 wire \core.work.registers.genblk1[2].latch[30] ;
 wire \core.work.registers.genblk1[2].latch[31] ;
 wire \core.work.registers.genblk1[2].latch[3] ;
 wire \core.work.registers.genblk1[2].latch[4] ;
 wire \core.work.registers.genblk1[2].latch[5] ;
 wire \core.work.registers.genblk1[2].latch[6] ;
 wire \core.work.registers.genblk1[2].latch[7] ;
 wire \core.work.registers.genblk1[2].latch[8] ;
 wire \core.work.registers.genblk1[2].latch[9] ;
 wire \core.work.registers.genblk1[2].we ;
 wire \core.work.registers.genblk1[3].latch[0] ;
 wire \core.work.registers.genblk1[3].latch[10] ;
 wire \core.work.registers.genblk1[3].latch[11] ;
 wire \core.work.registers.genblk1[3].latch[12] ;
 wire \core.work.registers.genblk1[3].latch[13] ;
 wire \core.work.registers.genblk1[3].latch[14] ;
 wire \core.work.registers.genblk1[3].latch[15] ;
 wire \core.work.registers.genblk1[3].latch[16] ;
 wire \core.work.registers.genblk1[3].latch[17] ;
 wire \core.work.registers.genblk1[3].latch[18] ;
 wire \core.work.registers.genblk1[3].latch[19] ;
 wire \core.work.registers.genblk1[3].latch[1] ;
 wire \core.work.registers.genblk1[3].latch[20] ;
 wire \core.work.registers.genblk1[3].latch[21] ;
 wire \core.work.registers.genblk1[3].latch[22] ;
 wire \core.work.registers.genblk1[3].latch[23] ;
 wire \core.work.registers.genblk1[3].latch[24] ;
 wire \core.work.registers.genblk1[3].latch[25] ;
 wire \core.work.registers.genblk1[3].latch[26] ;
 wire \core.work.registers.genblk1[3].latch[27] ;
 wire \core.work.registers.genblk1[3].latch[28] ;
 wire \core.work.registers.genblk1[3].latch[29] ;
 wire \core.work.registers.genblk1[3].latch[2] ;
 wire \core.work.registers.genblk1[3].latch[30] ;
 wire \core.work.registers.genblk1[3].latch[31] ;
 wire \core.work.registers.genblk1[3].latch[3] ;
 wire \core.work.registers.genblk1[3].latch[4] ;
 wire \core.work.registers.genblk1[3].latch[5] ;
 wire \core.work.registers.genblk1[3].latch[6] ;
 wire \core.work.registers.genblk1[3].latch[7] ;
 wire \core.work.registers.genblk1[3].latch[8] ;
 wire \core.work.registers.genblk1[3].latch[9] ;
 wire \core.work.registers.genblk1[3].we ;
 wire \core.work.registers.genblk1[4].latch[0] ;
 wire \core.work.registers.genblk1[4].latch[10] ;
 wire \core.work.registers.genblk1[4].latch[11] ;
 wire \core.work.registers.genblk1[4].latch[12] ;
 wire \core.work.registers.genblk1[4].latch[13] ;
 wire \core.work.registers.genblk1[4].latch[14] ;
 wire \core.work.registers.genblk1[4].latch[15] ;
 wire \core.work.registers.genblk1[4].latch[16] ;
 wire \core.work.registers.genblk1[4].latch[17] ;
 wire \core.work.registers.genblk1[4].latch[18] ;
 wire \core.work.registers.genblk1[4].latch[19] ;
 wire \core.work.registers.genblk1[4].latch[1] ;
 wire \core.work.registers.genblk1[4].latch[20] ;
 wire \core.work.registers.genblk1[4].latch[21] ;
 wire \core.work.registers.genblk1[4].latch[22] ;
 wire \core.work.registers.genblk1[4].latch[23] ;
 wire \core.work.registers.genblk1[4].latch[24] ;
 wire \core.work.registers.genblk1[4].latch[25] ;
 wire \core.work.registers.genblk1[4].latch[26] ;
 wire \core.work.registers.genblk1[4].latch[27] ;
 wire \core.work.registers.genblk1[4].latch[28] ;
 wire \core.work.registers.genblk1[4].latch[29] ;
 wire \core.work.registers.genblk1[4].latch[2] ;
 wire \core.work.registers.genblk1[4].latch[30] ;
 wire \core.work.registers.genblk1[4].latch[31] ;
 wire \core.work.registers.genblk1[4].latch[3] ;
 wire \core.work.registers.genblk1[4].latch[4] ;
 wire \core.work.registers.genblk1[4].latch[5] ;
 wire \core.work.registers.genblk1[4].latch[6] ;
 wire \core.work.registers.genblk1[4].latch[7] ;
 wire \core.work.registers.genblk1[4].latch[8] ;
 wire \core.work.registers.genblk1[4].latch[9] ;
 wire \core.work.registers.genblk1[4].we ;
 wire \core.work.registers.genblk1[5].latch[0] ;
 wire \core.work.registers.genblk1[5].latch[10] ;
 wire \core.work.registers.genblk1[5].latch[11] ;
 wire \core.work.registers.genblk1[5].latch[12] ;
 wire \core.work.registers.genblk1[5].latch[13] ;
 wire \core.work.registers.genblk1[5].latch[14] ;
 wire \core.work.registers.genblk1[5].latch[15] ;
 wire \core.work.registers.genblk1[5].latch[16] ;
 wire \core.work.registers.genblk1[5].latch[17] ;
 wire \core.work.registers.genblk1[5].latch[18] ;
 wire \core.work.registers.genblk1[5].latch[19] ;
 wire \core.work.registers.genblk1[5].latch[1] ;
 wire \core.work.registers.genblk1[5].latch[20] ;
 wire \core.work.registers.genblk1[5].latch[21] ;
 wire \core.work.registers.genblk1[5].latch[22] ;
 wire \core.work.registers.genblk1[5].latch[23] ;
 wire \core.work.registers.genblk1[5].latch[24] ;
 wire \core.work.registers.genblk1[5].latch[25] ;
 wire \core.work.registers.genblk1[5].latch[26] ;
 wire \core.work.registers.genblk1[5].latch[27] ;
 wire \core.work.registers.genblk1[5].latch[28] ;
 wire \core.work.registers.genblk1[5].latch[29] ;
 wire \core.work.registers.genblk1[5].latch[2] ;
 wire \core.work.registers.genblk1[5].latch[30] ;
 wire \core.work.registers.genblk1[5].latch[31] ;
 wire \core.work.registers.genblk1[5].latch[3] ;
 wire \core.work.registers.genblk1[5].latch[4] ;
 wire \core.work.registers.genblk1[5].latch[5] ;
 wire \core.work.registers.genblk1[5].latch[6] ;
 wire \core.work.registers.genblk1[5].latch[7] ;
 wire \core.work.registers.genblk1[5].latch[8] ;
 wire \core.work.registers.genblk1[5].latch[9] ;
 wire \core.work.registers.genblk1[5].we ;
 wire \core.work.registers.genblk1[6].latch[0] ;
 wire \core.work.registers.genblk1[6].latch[10] ;
 wire \core.work.registers.genblk1[6].latch[11] ;
 wire \core.work.registers.genblk1[6].latch[12] ;
 wire \core.work.registers.genblk1[6].latch[13] ;
 wire \core.work.registers.genblk1[6].latch[14] ;
 wire \core.work.registers.genblk1[6].latch[15] ;
 wire \core.work.registers.genblk1[6].latch[16] ;
 wire \core.work.registers.genblk1[6].latch[17] ;
 wire \core.work.registers.genblk1[6].latch[18] ;
 wire \core.work.registers.genblk1[6].latch[19] ;
 wire \core.work.registers.genblk1[6].latch[1] ;
 wire \core.work.registers.genblk1[6].latch[20] ;
 wire \core.work.registers.genblk1[6].latch[21] ;
 wire \core.work.registers.genblk1[6].latch[22] ;
 wire \core.work.registers.genblk1[6].latch[23] ;
 wire \core.work.registers.genblk1[6].latch[24] ;
 wire \core.work.registers.genblk1[6].latch[25] ;
 wire \core.work.registers.genblk1[6].latch[26] ;
 wire \core.work.registers.genblk1[6].latch[27] ;
 wire \core.work.registers.genblk1[6].latch[28] ;
 wire \core.work.registers.genblk1[6].latch[29] ;
 wire \core.work.registers.genblk1[6].latch[2] ;
 wire \core.work.registers.genblk1[6].latch[30] ;
 wire \core.work.registers.genblk1[6].latch[31] ;
 wire \core.work.registers.genblk1[6].latch[3] ;
 wire \core.work.registers.genblk1[6].latch[4] ;
 wire \core.work.registers.genblk1[6].latch[5] ;
 wire \core.work.registers.genblk1[6].latch[6] ;
 wire \core.work.registers.genblk1[6].latch[7] ;
 wire \core.work.registers.genblk1[6].latch[8] ;
 wire \core.work.registers.genblk1[6].latch[9] ;
 wire \core.work.registers.genblk1[6].we ;
 wire \core.work.registers.genblk1[7].latch[0] ;
 wire \core.work.registers.genblk1[7].latch[10] ;
 wire \core.work.registers.genblk1[7].latch[11] ;
 wire \core.work.registers.genblk1[7].latch[12] ;
 wire \core.work.registers.genblk1[7].latch[13] ;
 wire \core.work.registers.genblk1[7].latch[14] ;
 wire \core.work.registers.genblk1[7].latch[15] ;
 wire \core.work.registers.genblk1[7].latch[16] ;
 wire \core.work.registers.genblk1[7].latch[17] ;
 wire \core.work.registers.genblk1[7].latch[18] ;
 wire \core.work.registers.genblk1[7].latch[19] ;
 wire \core.work.registers.genblk1[7].latch[1] ;
 wire \core.work.registers.genblk1[7].latch[20] ;
 wire \core.work.registers.genblk1[7].latch[21] ;
 wire \core.work.registers.genblk1[7].latch[22] ;
 wire \core.work.registers.genblk1[7].latch[23] ;
 wire \core.work.registers.genblk1[7].latch[24] ;
 wire \core.work.registers.genblk1[7].latch[25] ;
 wire \core.work.registers.genblk1[7].latch[26] ;
 wire \core.work.registers.genblk1[7].latch[27] ;
 wire \core.work.registers.genblk1[7].latch[28] ;
 wire \core.work.registers.genblk1[7].latch[29] ;
 wire \core.work.registers.genblk1[7].latch[2] ;
 wire \core.work.registers.genblk1[7].latch[30] ;
 wire \core.work.registers.genblk1[7].latch[31] ;
 wire \core.work.registers.genblk1[7].latch[3] ;
 wire \core.work.registers.genblk1[7].latch[4] ;
 wire \core.work.registers.genblk1[7].latch[5] ;
 wire \core.work.registers.genblk1[7].latch[6] ;
 wire \core.work.registers.genblk1[7].latch[7] ;
 wire \core.work.registers.genblk1[7].latch[8] ;
 wire \core.work.registers.genblk1[7].latch[9] ;
 wire \core.work.registers.genblk1[7].we ;
 wire \core.work.registers.genblk1[8].latch[0] ;
 wire \core.work.registers.genblk1[8].latch[10] ;
 wire \core.work.registers.genblk1[8].latch[11] ;
 wire \core.work.registers.genblk1[8].latch[12] ;
 wire \core.work.registers.genblk1[8].latch[13] ;
 wire \core.work.registers.genblk1[8].latch[14] ;
 wire \core.work.registers.genblk1[8].latch[15] ;
 wire \core.work.registers.genblk1[8].latch[16] ;
 wire \core.work.registers.genblk1[8].latch[17] ;
 wire \core.work.registers.genblk1[8].latch[18] ;
 wire \core.work.registers.genblk1[8].latch[19] ;
 wire \core.work.registers.genblk1[8].latch[1] ;
 wire \core.work.registers.genblk1[8].latch[20] ;
 wire \core.work.registers.genblk1[8].latch[21] ;
 wire \core.work.registers.genblk1[8].latch[22] ;
 wire \core.work.registers.genblk1[8].latch[23] ;
 wire \core.work.registers.genblk1[8].latch[24] ;
 wire \core.work.registers.genblk1[8].latch[25] ;
 wire \core.work.registers.genblk1[8].latch[26] ;
 wire \core.work.registers.genblk1[8].latch[27] ;
 wire \core.work.registers.genblk1[8].latch[28] ;
 wire \core.work.registers.genblk1[8].latch[29] ;
 wire \core.work.registers.genblk1[8].latch[2] ;
 wire \core.work.registers.genblk1[8].latch[30] ;
 wire \core.work.registers.genblk1[8].latch[31] ;
 wire \core.work.registers.genblk1[8].latch[3] ;
 wire \core.work.registers.genblk1[8].latch[4] ;
 wire \core.work.registers.genblk1[8].latch[5] ;
 wire \core.work.registers.genblk1[8].latch[6] ;
 wire \core.work.registers.genblk1[8].latch[7] ;
 wire \core.work.registers.genblk1[8].latch[8] ;
 wire \core.work.registers.genblk1[8].latch[9] ;
 wire \core.work.registers.genblk1[8].we ;
 wire \core.work.registers.genblk1[9].latch[0] ;
 wire \core.work.registers.genblk1[9].latch[10] ;
 wire \core.work.registers.genblk1[9].latch[11] ;
 wire \core.work.registers.genblk1[9].latch[12] ;
 wire \core.work.registers.genblk1[9].latch[13] ;
 wire \core.work.registers.genblk1[9].latch[14] ;
 wire \core.work.registers.genblk1[9].latch[15] ;
 wire \core.work.registers.genblk1[9].latch[16] ;
 wire \core.work.registers.genblk1[9].latch[17] ;
 wire \core.work.registers.genblk1[9].latch[18] ;
 wire \core.work.registers.genblk1[9].latch[19] ;
 wire \core.work.registers.genblk1[9].latch[1] ;
 wire \core.work.registers.genblk1[9].latch[20] ;
 wire \core.work.registers.genblk1[9].latch[21] ;
 wire \core.work.registers.genblk1[9].latch[22] ;
 wire \core.work.registers.genblk1[9].latch[23] ;
 wire \core.work.registers.genblk1[9].latch[24] ;
 wire \core.work.registers.genblk1[9].latch[25] ;
 wire \core.work.registers.genblk1[9].latch[26] ;
 wire \core.work.registers.genblk1[9].latch[27] ;
 wire \core.work.registers.genblk1[9].latch[28] ;
 wire \core.work.registers.genblk1[9].latch[29] ;
 wire \core.work.registers.genblk1[9].latch[2] ;
 wire \core.work.registers.genblk1[9].latch[30] ;
 wire \core.work.registers.genblk1[9].latch[31] ;
 wire \core.work.registers.genblk1[9].latch[3] ;
 wire \core.work.registers.genblk1[9].latch[4] ;
 wire \core.work.registers.genblk1[9].latch[5] ;
 wire \core.work.registers.genblk1[9].latch[6] ;
 wire \core.work.registers.genblk1[9].latch[7] ;
 wire \core.work.registers.genblk1[9].latch[8] ;
 wire \core.work.registers.genblk1[9].latch[9] ;
 wire \core.work.registers.genblk1[9].we ;
 wire \core.work.registers.state[0] ;
 wire \core.work.registers.state[1] ;
 wire \core.work.registers.state[2] ;
 wire \core.work.registers.tmp[0] ;
 wire \core.work.registers.tmp[10] ;
 wire \core.work.registers.tmp[11] ;
 wire \core.work.registers.tmp[12] ;
 wire \core.work.registers.tmp[13] ;
 wire \core.work.registers.tmp[14] ;
 wire \core.work.registers.tmp[15] ;
 wire \core.work.registers.tmp[16] ;
 wire \core.work.registers.tmp[17] ;
 wire \core.work.registers.tmp[18] ;
 wire \core.work.registers.tmp[19] ;
 wire \core.work.registers.tmp[1] ;
 wire \core.work.registers.tmp[20] ;
 wire \core.work.registers.tmp[21] ;
 wire \core.work.registers.tmp[22] ;
 wire \core.work.registers.tmp[23] ;
 wire \core.work.registers.tmp[24] ;
 wire \core.work.registers.tmp[25] ;
 wire \core.work.registers.tmp[26] ;
 wire \core.work.registers.tmp[27] ;
 wire \core.work.registers.tmp[28] ;
 wire \core.work.registers.tmp[29] ;
 wire \core.work.registers.tmp[2] ;
 wire \core.work.registers.tmp[30] ;
 wire \core.work.registers.tmp[31] ;
 wire \core.work.registers.tmp[3] ;
 wire \core.work.registers.tmp[4] ;
 wire \core.work.registers.tmp[5] ;
 wire \core.work.registers.tmp[6] ;
 wire \core.work.registers.tmp[7] ;
 wire \core.work.registers.tmp[8] ;
 wire \core.work.registers.tmp[9] ;
 wire \core.work.registers.wr_reg[0] ;
 wire \core.work.registers.wr_reg[1] ;
 wire \core.work.registers.wr_reg[2] ;
 wire \core.work.registers.wr_reg[3] ;
 wire \core.work.state[0] ;
 wire \core.work.state[1] ;
 wire net336;
 wire net337;
 wire net12;
 wire net338;
 wire net339;
 wire net340;
 wire net13;
 wire net341;
 wire net14;
 wire net15;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_47_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_leaf_53_clk_regs;
 wire clknet_leaf_54_clk_regs;
 wire clknet_leaf_55_clk_regs;
 wire clknet_leaf_56_clk_regs;
 wire clknet_leaf_57_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire delaynet_0_clk;
 wire delaynet_1_clk;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;

 sg13g2_inv_1 _06014_ (.Y(_00579_),
    .A(net579));
 sg13g2_inv_1 _06015_ (.Y(_00580_),
    .A(net3527));
 sg13g2_inv_1 _06016_ (.Y(_00581_),
    .A(\core.fetch.inst_size[1] ));
 sg13g2_inv_1 _06017_ (.Y(_00582_),
    .A(\core.f2e_inst[1] ));
 sg13g2_inv_1 _06018_ (.Y(_00583_),
    .A(net717));
 sg13g2_inv_1 _06019_ (.Y(_00584_),
    .A(net836));
 sg13g2_inv_2 _06020_ (.Y(_00585_),
    .A(net746));
 sg13g2_inv_1 _06021_ (.Y(_00586_),
    .A(net445));
 sg13g2_inv_1 _06022_ (.Y(_00587_),
    .A(_00018_));
 sg13g2_inv_1 _06023_ (.Y(_00588_),
    .A(\core.fetch.state[0] ));
 sg13g2_inv_1 _06024_ (.Y(_00589_),
    .A(net3500));
 sg13g2_inv_4 _06025_ (.A(net3561),
    .Y(_00590_));
 sg13g2_inv_1 _06026_ (.Y(_00591_),
    .A(net3499));
 sg13g2_inv_1 _06027_ (.Y(_00592_),
    .A(net3553));
 sg13g2_inv_1 _06028_ (.Y(_00593_),
    .A(\core.e2m_addr[7] ));
 sg13g2_inv_2 _06029_ (.Y(_00594_),
    .A(\core.e2m_addr[6] ));
 sg13g2_inv_4 _06030_ (.A(net3493),
    .Y(_00595_));
 sg13g2_inv_2 _06031_ (.Y(_00596_),
    .A(net3549));
 sg13g2_inv_1 _06032_ (.Y(_00597_),
    .A(net704));
 sg13g2_inv_1 _06033_ (.Y(_00598_),
    .A(\core.work.alu.sval2[15] ));
 sg13g2_inv_2 _06034_ (.Y(_00599_),
    .A(net3478));
 sg13g2_inv_4 _06035_ (.A(net3480),
    .Y(_00600_));
 sg13g2_inv_4 _06036_ (.A(net3484),
    .Y(_00601_));
 sg13g2_inv_1 _06037_ (.Y(_00602_),
    .A(\core.work.alu.sval2[10] ));
 sg13g2_inv_1 _06038_ (.Y(_00603_),
    .A(net892));
 sg13g2_inv_1 _06039_ (.Y(_00604_),
    .A(\core.work.alu.sval2[31] ));
 sg13g2_inv_4 _06040_ (.A(net3443),
    .Y(_00605_));
 sg13g2_inv_1 _06041_ (.Y(_00606_),
    .A(\core.work.alu.sval2[30] ));
 sg13g2_inv_1 _06042_ (.Y(_00607_),
    .A(net3444));
 sg13g2_inv_1 _06043_ (.Y(_00608_),
    .A(net3540));
 sg13g2_inv_1 _06044_ (.Y(_00609_),
    .A(net3445));
 sg13g2_inv_1 _06045_ (.Y(_00610_),
    .A(net832));
 sg13g2_inv_4 _06046_ (.A(net3448),
    .Y(_00611_));
 sg13g2_inv_1 _06047_ (.Y(_00612_),
    .A(net791));
 sg13g2_inv_4 _06048_ (.A(\core.e2m_addr[26] ),
    .Y(_00613_));
 sg13g2_inv_1 _06049_ (.Y(_00614_),
    .A(net3533));
 sg13g2_inv_1 _06050_ (.Y(_00615_),
    .A(\core.e2m_addr[24] ));
 sg13g2_inv_1 _06051_ (.Y(_00616_),
    .A(net3534));
 sg13g2_inv_1 _06052_ (.Y(_00617_),
    .A(net3453));
 sg13g2_inv_1 _06053_ (.Y(_00618_),
    .A(\core.work.alu.sval2[22] ));
 sg13g2_inv_1 _06054_ (.Y(_00619_),
    .A(\core.work.alu.sval2[21] ));
 sg13g2_inv_1 _06055_ (.Y(_00620_),
    .A(net3458));
 sg13g2_inv_1 _06056_ (.Y(_00621_),
    .A(net459));
 sg13g2_inv_2 _06057_ (.Y(_00622_),
    .A(net3465));
 sg13g2_inv_1 _06058_ (.Y(_00623_),
    .A(\core.e2m_addr[19] ));
 sg13g2_inv_1 _06059_ (.Y(_00624_),
    .A(net3531));
 sg13g2_inv_1 _06060_ (.Y(_00625_),
    .A(\core.work.alu.sval2[18] ));
 sg13g2_inv_1 _06061_ (.Y(_00626_),
    .A(net708));
 sg13g2_inv_1 _06062_ (.Y(_00627_),
    .A(net3532));
 sg13g2_inv_1 _06063_ (.Y(_00628_),
    .A(net3470));
 sg13g2_inv_2 _06064_ (.Y(_00629_),
    .A(net865));
 sg13g2_inv_1 _06065_ (.Y(_00630_),
    .A(net666));
 sg13g2_inv_1 _06066_ (.Y(_00631_),
    .A(net3566));
 sg13g2_inv_1 _06067_ (.Y(_00632_),
    .A(net781));
 sg13g2_inv_1 _06068_ (.Y(_00633_),
    .A(net829));
 sg13g2_inv_1 _06069_ (.Y(_00634_),
    .A(_00021_));
 sg13g2_inv_1 _06070_ (.Y(_00635_),
    .A(net798));
 sg13g2_inv_1 _06071_ (.Y(_00636_),
    .A(net3442));
 sg13g2_inv_1 _06072_ (.Y(_00637_),
    .A(_00027_));
 sg13g2_inv_1 _06073_ (.Y(_00638_),
    .A(_00028_));
 sg13g2_inv_1 _06074_ (.Y(_00639_),
    .A(_00030_));
 sg13g2_inv_2 _06075_ (.Y(_00640_),
    .A(_00033_));
 sg13g2_inv_1 _06076_ (.Y(_00641_),
    .A(_00035_));
 sg13g2_inv_2 _06077_ (.Y(_00642_),
    .A(_00036_));
 sg13g2_inv_1 _06078_ (.Y(_00643_),
    .A(_00037_));
 sg13g2_inv_1 _06079_ (.Y(_00644_),
    .A(_00043_));
 sg13g2_inv_2 _06080_ (.Y(_00645_),
    .A(_00046_));
 sg13g2_inv_1 _06081_ (.Y(_00646_),
    .A(_00048_));
 sg13g2_inv_1 _06082_ (.Y(_00647_),
    .A(_00049_));
 sg13g2_inv_2 _06083_ (.Y(_00648_),
    .A(_00052_));
 sg13g2_inv_1 _06084_ (.Y(_00649_),
    .A(net3577));
 sg13g2_inv_1 _06085_ (.Y(_00650_),
    .A(\core.fetch.data_size[1] ));
 sg13g2_inv_1 _06086_ (.Y(_00651_),
    .A(net762));
 sg13g2_inv_2 _06087_ (.Y(_00652_),
    .A(\core.fetch.rd_addr_i[0] ));
 sg13g2_inv_2 _06088_ (.Y(_00653_),
    .A(net834));
 sg13g2_inv_1 _06089_ (.Y(_00654_),
    .A(net841));
 sg13g2_inv_2 _06090_ (.Y(_00655_),
    .A(net809));
 sg13g2_inv_2 _06091_ (.Y(_00656_),
    .A(_00062_));
 sg13g2_inv_1 _06092_ (.Y(_00657_),
    .A(net3503));
 sg13g2_inv_1 _06093_ (.Y(_00658_),
    .A(\core.fetch.spi_reader.addr[3] ));
 sg13g2_inv_1 _06094_ (.Y(_00659_),
    .A(\core.fetch.spi_reader.addr[2] ));
 sg13g2_inv_1 _06095_ (.Y(_00660_),
    .A(net613));
 sg13g2_inv_1 _06096_ (.Y(_00661_),
    .A(\core.fetch.spi_reader.addr[7] ));
 sg13g2_inv_1 _06097_ (.Y(_00662_),
    .A(_00070_));
 sg13g2_inv_1 _06098_ (.Y(_00663_),
    .A(net759));
 sg13g2_inv_1 _06099_ (.Y(_00664_),
    .A(net777));
 sg13g2_inv_1 _06100_ (.Y(_00665_),
    .A(_00080_));
 sg13g2_inv_2 _06101_ (.Y(_00666_),
    .A(\core.lsu.spi.cs ));
 sg13g2_inv_1 _06102_ (.Y(_00667_),
    .A(net550));
 sg13g2_inv_1 _06103_ (.Y(_00668_),
    .A(_00088_));
 sg13g2_inv_1 _06104_ (.Y(_00669_),
    .A(net372));
 sg13g2_inv_1 _06105_ (.Y(_00670_),
    .A(_00090_));
 sg13g2_inv_1 _06106_ (.Y(_00671_),
    .A(net549));
 sg13g2_inv_1 _06107_ (.Y(_00672_),
    .A(net819));
 sg13g2_inv_1 _06108_ (.Y(_00673_),
    .A(net609));
 sg13g2_inv_1 _06109_ (.Y(_00674_),
    .A(_00093_));
 sg13g2_inv_1 _06110_ (.Y(_00675_),
    .A(net578));
 sg13g2_inv_1 _06111_ (.Y(_00676_),
    .A(net472));
 sg13g2_inv_1 _06112_ (.Y(_00677_),
    .A(net506));
 sg13g2_inv_1 _06113_ (.Y(_00678_),
    .A(\core.f2e_inst[18] ));
 sg13g2_inv_1 _06114_ (.Y(_00679_),
    .A(net585));
 sg13g2_inv_1 _06115_ (.Y(_00680_),
    .A(\core.f2e_inst[2] ));
 sg13g2_inv_2 _06116_ (.Y(_00681_),
    .A(net884));
 sg13g2_inv_1 _06117_ (.Y(_00682_),
    .A(net531));
 sg13g2_inv_1 _06118_ (.Y(_00683_),
    .A(\core.f2e_inst[3] ));
 sg13g2_inv_2 _06119_ (.Y(_00684_),
    .A(net571));
 sg13g2_inv_1 _06120_ (.Y(_00685_),
    .A(net520));
 sg13g2_inv_4 _06121_ (.A(\core.fetch.cmd_data[4] ),
    .Y(_00686_));
 sg13g2_inv_1 _06122_ (.Y(_00687_),
    .A(\core.f2e_inst[21] ));
 sg13g2_inv_1 _06123_ (.Y(_00688_),
    .A(net581));
 sg13g2_inv_4 _06124_ (.A(\core.fetch.cmd_data[5] ),
    .Y(_00689_));
 sg13g2_inv_1 _06125_ (.Y(_00690_),
    .A(net536));
 sg13g2_inv_4 _06126_ (.A(net565),
    .Y(_00691_));
 sg13g2_inv_1 _06127_ (.Y(_00692_),
    .A(net539));
 sg13g2_inv_2 _06128_ (.Y(_00693_),
    .A(\core.fetch.cmd_data[7] ));
 sg13g2_inv_1 _06129_ (.Y(_00694_),
    .A(net528));
 sg13g2_inv_1 _06130_ (.Y(_00695_),
    .A(\core.f2e_inst[8] ));
 sg13g2_inv_1 _06131_ (.Y(_00696_),
    .A(net524));
 sg13g2_inv_1 _06132_ (.Y(_00697_),
    .A(net553));
 sg13g2_inv_1 _06133_ (.Y(_00698_),
    .A(net564));
 sg13g2_inv_2 _06134_ (.Y(_00699_),
    .A(\core.f2e_inst[11] ));
 sg13g2_inv_1 _06135_ (.Y(_00700_),
    .A(net563));
 sg13g2_inv_2 _06136_ (.Y(_00701_),
    .A(net3507));
 sg13g2_inv_1 _06137_ (.Y(_00702_),
    .A(net530));
 sg13g2_inv_1 _06138_ (.Y(_00703_),
    .A(\core.f2e_inst[30] ));
 sg13g2_inv_1 _06139_ (.Y(_00704_),
    .A(net574));
 sg13g2_inv_2 _06140_ (.Y(_00705_),
    .A(\core.f2e_inst[14] ));
 sg13g2_inv_1 _06141_ (.Y(_00706_),
    .A(\core.f2e_inst[31] ));
 sg13g2_inv_1 _06142_ (.Y(_00707_),
    .A(net534));
 sg13g2_inv_2 _06143_ (.Y(_00708_),
    .A(\core.f2e_inst[15] ));
 sg13g2_inv_1 _06144_ (.Y(_00709_),
    .A(net374));
 sg13g2_inv_1 _06145_ (.Y(_00710_),
    .A(net457));
 sg13g2_inv_1 _06146_ (.Y(_00711_),
    .A(net463));
 sg13g2_inv_1 _06147_ (.Y(_00712_),
    .A(net546));
 sg13g2_inv_2 _06148_ (.Y(_00713_),
    .A(net454));
 sg13g2_inv_1 _06149_ (.Y(_00714_),
    .A(_00110_));
 sg13g2_inv_1 _06150_ (.Y(_00715_),
    .A(_00111_));
 sg13g2_inv_1 _06151_ (.Y(_00716_),
    .A(_00112_));
 sg13g2_inv_1 _06152_ (.Y(_00717_),
    .A(_00113_));
 sg13g2_inv_1 _06153_ (.Y(_00718_),
    .A(_00114_));
 sg13g2_inv_1 _06154_ (.Y(_00719_),
    .A(_00115_));
 sg13g2_inv_1 _06155_ (.Y(_00720_),
    .A(_00116_));
 sg13g2_inv_1 _06156_ (.Y(_00721_),
    .A(_00118_));
 sg13g2_inv_1 _06157_ (.Y(_00722_),
    .A(_00119_));
 sg13g2_inv_1 _06158_ (.Y(_00723_),
    .A(_00123_));
 sg13g2_inv_1 _06159_ (.Y(_00724_),
    .A(net634));
 sg13g2_inv_1 _06160_ (.Y(_00725_),
    .A(net738));
 sg13g2_inv_1 _06161_ (.Y(_00726_),
    .A(net646));
 sg13g2_inv_1 _06162_ (.Y(_00727_),
    .A(net807));
 sg13g2_inv_1 _06163_ (.Y(_00728_),
    .A(net750));
 sg13g2_inv_1 _06164_ (.Y(_00729_),
    .A(net650));
 sg13g2_inv_1 _06165_ (.Y(_00730_),
    .A(_00141_));
 sg13g2_inv_1 _06166_ (.Y(_00731_),
    .A(_00145_));
 sg13g2_inv_1 _06167_ (.Y(_00732_),
    .A(_00146_));
 sg13g2_inv_1 _06168_ (.Y(_00733_),
    .A(_00153_));
 sg13g2_inv_1 _11282__2 (.Y(net342),
    .A(clknet_2_1__leaf_clk));
 sg13g2_nand3_1 _06170_ (.B(_00651_),
    .C(_00058_),
    .A(\core.work.registers.state[1] ),
    .Y(_00734_));
 sg13g2_or2_1 _06171_ (.X(_00735_),
    .B(\core.work.registers.state[0] ),
    .A(\core.work.registers.state[1] ));
 sg13g2_nand3b_1 _06172_ (.B(_00651_),
    .C(net544),
    .Y(_00736_),
    .A_N(\core.work.registers.state[1] ));
 sg13g2_and2_1 _06173_ (.A(_00734_),
    .B(_00736_),
    .X(_00737_));
 sg13g2_nand2_1 _06174_ (.Y(_00738_),
    .A(_00734_),
    .B(_00736_));
 sg13g2_nand3_1 _06175_ (.B(\core.work.registers.wr_reg[1] ),
    .C(_00738_),
    .A(\core.work.registers.wr_reg[0] ),
    .Y(_00739_));
 sg13g2_nand2_2 _06176_ (.Y(_00740_),
    .A(\core.work.registers.wr_reg[2] ),
    .B(\core.work.registers.wr_reg[3] ));
 sg13g2_nor2_1 _06177_ (.A(_00739_),
    .B(_00740_),
    .Y(_00008_));
 sg13g2_nor2_2 _06178_ (.A(\core.work.registers.wr_reg[0] ),
    .B(_00737_),
    .Y(_00741_));
 sg13g2_nand2_2 _06179_ (.Y(_00742_),
    .A(\core.work.registers.wr_reg[1] ),
    .B(_00741_));
 sg13g2_nor2_1 _06180_ (.A(_00740_),
    .B(_00742_),
    .Y(_00007_));
 sg13g2_nand3b_1 _06181_ (.B(_00738_),
    .C(\core.work.registers.wr_reg[0] ),
    .Y(_00743_),
    .A_N(\core.work.registers.wr_reg[1] ));
 sg13g2_nor2_1 _06182_ (.A(_00740_),
    .B(_00743_),
    .Y(_00006_));
 sg13g2_nand2b_2 _06183_ (.Y(_00744_),
    .B(_00741_),
    .A_N(\core.work.registers.wr_reg[1] ));
 sg13g2_nor2_1 _06184_ (.A(_00740_),
    .B(_00744_),
    .Y(_00005_));
 sg13g2_nand2b_2 _06185_ (.Y(_00745_),
    .B(\core.work.registers.wr_reg[3] ),
    .A_N(\core.work.registers.wr_reg[2] ));
 sg13g2_nor2_1 _06186_ (.A(_00739_),
    .B(_00745_),
    .Y(_00004_));
 sg13g2_nor2_1 _06187_ (.A(_00742_),
    .B(_00745_),
    .Y(_00003_));
 sg13g2_nor2_1 _06188_ (.A(_00743_),
    .B(_00745_),
    .Y(_00017_));
 sg13g2_nor2_1 _06189_ (.A(_00744_),
    .B(_00745_),
    .Y(_00016_));
 sg13g2_nand2b_2 _06190_ (.Y(_00746_),
    .B(\core.work.registers.wr_reg[2] ),
    .A_N(\core.work.registers.wr_reg[3] ));
 sg13g2_nor2_1 _06191_ (.A(_00739_),
    .B(_00746_),
    .Y(_00015_));
 sg13g2_nor2_1 _06192_ (.A(_00742_),
    .B(_00746_),
    .Y(_00014_));
 sg13g2_nor2_1 _06193_ (.A(_00743_),
    .B(_00746_),
    .Y(_00013_));
 sg13g2_nor2_1 _06194_ (.A(_00744_),
    .B(_00746_),
    .Y(_00012_));
 sg13g2_nor3_1 _06195_ (.A(\core.work.registers.wr_reg[2] ),
    .B(\core.work.registers.wr_reg[3] ),
    .C(_00739_),
    .Y(_00011_));
 sg13g2_nor3_1 _06196_ (.A(\core.work.registers.wr_reg[2] ),
    .B(\core.work.registers.wr_reg[3] ),
    .C(_00742_),
    .Y(_00010_));
 sg13g2_nor3_1 _06197_ (.A(\core.work.registers.wr_reg[2] ),
    .B(\core.work.registers.wr_reg[3] ),
    .C(_00743_),
    .Y(_00009_));
 sg13g2_nor2b_2 _06198_ (.A(\core.fetch.spi_reader.state[0] ),
    .B_N(_00060_),
    .Y(_00747_));
 sg13g2_nor2b_2 _06199_ (.A(net3567),
    .B_N(_00747_),
    .Y(_00748_));
 sg13g2_nand2b_2 _06200_ (.Y(_00749_),
    .B(_00747_),
    .A_N(net3567));
 sg13g2_and4_1 _06201_ (.A(\core.fetch.rd_addr_i[9] ),
    .B(\core.fetch.rd_addr_i[8] ),
    .C(\core.fetch.rd_addr_i[11] ),
    .D(\core.fetch.rd_addr_i[10] ),
    .X(_00750_));
 sg13g2_nand4_1 _06202_ (.B(\core.fetch.rd_addr_i[8] ),
    .C(\core.fetch.rd_addr_i[11] ),
    .A(\core.fetch.rd_addr_i[9] ),
    .Y(_00751_),
    .D(\core.fetch.rd_addr_i[10] ));
 sg13g2_nand2_2 _06203_ (.Y(_00752_),
    .A(\core.fetch.rd_addr_i[5] ),
    .B(\core.fetch.rd_addr_i[4] ));
 sg13g2_nand4_1 _06204_ (.B(\core.fetch.rd_addr_i[4] ),
    .C(\core.fetch.rd_addr_i[7] ),
    .A(\core.fetch.rd_addr_i[5] ),
    .Y(_00753_),
    .D(\core.fetch.rd_addr_i[6] ));
 sg13g2_and2_1 _06205_ (.A(\core.fetch.data_size[2] ),
    .B(\core.fetch.rd_addr_i[2] ),
    .X(_00754_));
 sg13g2_nand2b_2 _06206_ (.Y(_00755_),
    .B(_00754_),
    .A_N(_00066_));
 sg13g2_nand2_1 _06207_ (.Y(_00756_),
    .A(net3576),
    .B(net3526));
 sg13g2_nand2_2 _06208_ (.Y(_00757_),
    .A(net3577),
    .B(\core.fetch.rd_addr_i[0] ));
 sg13g2_nor2_1 _06209_ (.A(net3576),
    .B(net3526),
    .Y(_00758_));
 sg13g2_xor2_1 _06210_ (.B(net3526),
    .A(net3576),
    .X(_00759_));
 sg13g2_o21ai_1 _06211_ (.B1(_00756_),
    .Y(_00760_),
    .A1(_00757_),
    .A2(_00758_));
 sg13g2_xor2_1 _06212_ (.B(\core.fetch.rd_addr_i[2] ),
    .A(\core.fetch.data_size[2] ),
    .X(_00761_));
 sg13g2_nand3_1 _06213_ (.B(_00760_),
    .C(_00761_),
    .A(\core.fetch.rd_addr_i[3] ),
    .Y(_00762_));
 sg13g2_a21oi_2 _06214_ (.B1(_00753_),
    .Y(_00763_),
    .A2(_00762_),
    .A1(_00755_));
 sg13g2_nand3_1 _06215_ (.B(_00750_),
    .C(_00763_),
    .A(net3525),
    .Y(_00764_));
 sg13g2_and2_1 _06216_ (.A(\core.fetch.state[1] ),
    .B(\core.fetch.state[0] ),
    .X(_00765_));
 sg13g2_nand2_1 _06217_ (.Y(_00766_),
    .A(\core.fetch.state[1] ),
    .B(\core.fetch.state[0] ));
 sg13g2_nand4_1 _06218_ (.B(net3525),
    .C(_00750_),
    .A(\core.fetch.rd_addr_i[13] ),
    .Y(_00767_),
    .D(_00763_));
 sg13g2_nor2_1 _06219_ (.A(_00073_),
    .B(_00767_),
    .Y(_00768_));
 sg13g2_or2_1 _06220_ (.X(_00769_),
    .B(_00768_),
    .A(_00072_));
 sg13g2_a21oi_1 _06221_ (.A1(_00072_),
    .A2(_00768_),
    .Y(_00770_),
    .B1(net3353));
 sg13g2_nand2_1 _06222_ (.Y(_00771_),
    .A(\core.fetch.inst_size[2] ),
    .B(\core.f2e_addr[2] ));
 sg13g2_nand2_2 _06223_ (.Y(_00772_),
    .A(net3528),
    .B(net3503));
 sg13g2_xnor2_1 _06224_ (.Y(_00773_),
    .A(\core.fetch.inst_size[2] ),
    .B(\core.f2e_addr[2] ));
 sg13g2_o21ai_1 _06225_ (.B1(_00771_),
    .Y(_00774_),
    .A1(_00772_),
    .A2(_00773_));
 sg13g2_and3_1 _06226_ (.X(_00775_),
    .A(\core.f2e_addr[3] ),
    .B(net3564),
    .C(_00774_));
 sg13g2_nand2_1 _06227_ (.Y(_00776_),
    .A(\core.f2e_addr[6] ),
    .B(\core.f2e_addr[5] ));
 sg13g2_inv_1 _06228_ (.Y(_00777_),
    .A(_00776_));
 sg13g2_and4_2 _06229_ (.A(\core.f2e_addr[3] ),
    .B(net3564),
    .C(_00774_),
    .D(_00777_),
    .X(_00778_));
 sg13g2_nand3_1 _06230_ (.B(\core.f2e_addr[8] ),
    .C(_00778_),
    .A(net3563),
    .Y(_00779_));
 sg13g2_nand4_1 _06231_ (.B(\core.f2e_addr[9] ),
    .C(\core.f2e_addr[8] ),
    .A(net3563),
    .Y(_00780_),
    .D(_00778_));
 sg13g2_and2_1 _06232_ (.A(\core.f2e_addr[10] ),
    .B(\core.f2e_addr[9] ),
    .X(_00781_));
 sg13g2_or2_1 _06233_ (.X(_00782_),
    .B(_00780_),
    .A(_00663_));
 sg13g2_nand2_1 _06234_ (.Y(_00783_),
    .A(\core.f2e_addr[14] ),
    .B(\core.f2e_addr[13] ));
 sg13g2_and3_1 _06235_ (.X(_00784_),
    .A(\core.f2e_addr[12] ),
    .B(\core.f2e_addr[11] ),
    .C(_00781_));
 sg13g2_nand3_1 _06236_ (.B(\core.f2e_addr[11] ),
    .C(_00781_),
    .A(\core.f2e_addr[12] ),
    .Y(_00785_));
 sg13g2_nor3_1 _06237_ (.A(_00779_),
    .B(_00783_),
    .C(_00785_),
    .Y(_00786_));
 sg13g2_xnor2_1 _06238_ (.Y(_00787_),
    .A(\core.f2e_addr[15] ),
    .B(_00786_));
 sg13g2_a22oi_1 _06239_ (.Y(_00788_),
    .B1(_00787_),
    .B2(net3353),
    .A2(_00770_),
    .A1(_00769_));
 sg13g2_inv_1 _06240_ (.Y(_00789_),
    .A(_00788_));
 sg13g2_nor2_1 _06241_ (.A(\core.fetch.spi_reader.addr[15] ),
    .B(_00789_),
    .Y(_00790_));
 sg13g2_xor2_1 _06242_ (.B(_00788_),
    .A(_00071_),
    .X(_00791_));
 sg13g2_nand2_1 _06243_ (.Y(_00792_),
    .A(\core.fetch.rd_addr_i[8] ),
    .B(_00763_));
 sg13g2_xnor2_1 _06244_ (.Y(_00793_),
    .A(_00082_),
    .B(_00792_));
 sg13g2_nand2b_1 _06245_ (.Y(_00794_),
    .B(_00779_),
    .A_N(\core.f2e_addr[9] ));
 sg13g2_a21oi_1 _06246_ (.A1(_00780_),
    .A2(_00794_),
    .Y(_00795_),
    .B1(net3356));
 sg13g2_a21oi_2 _06247_ (.B1(_00795_),
    .Y(_00796_),
    .A2(_00793_),
    .A1(net3356));
 sg13g2_nor2b_1 _06248_ (.A(\core.fetch.spi_reader.addr[9] ),
    .B_N(_00796_),
    .Y(_00797_));
 sg13g2_nand2b_1 _06249_ (.Y(_00798_),
    .B(\core.fetch.spi_reader.addr[9] ),
    .A_N(_00796_));
 sg13g2_nor2b_1 _06250_ (.A(_00797_),
    .B_N(_00798_),
    .Y(_00799_));
 sg13g2_xnor2_1 _06251_ (.Y(_00800_),
    .A(_00655_),
    .B(_00763_));
 sg13g2_a21oi_1 _06252_ (.A1(\core.f2e_addr[7] ),
    .A2(_00778_),
    .Y(_00801_),
    .B1(\core.f2e_addr[8] ));
 sg13g2_nor2_1 _06253_ (.A(net3357),
    .B(_00801_),
    .Y(_00802_));
 sg13g2_a22oi_1 _06254_ (.Y(_00803_),
    .B1(_00802_),
    .B2(_00779_),
    .A2(_00800_),
    .A1(net3356));
 sg13g2_xnor2_1 _06255_ (.Y(_00804_),
    .A(_00083_),
    .B(_00803_));
 sg13g2_nand2_1 _06256_ (.Y(_00805_),
    .A(_00799_),
    .B(_00804_));
 sg13g2_xor2_1 _06257_ (.B(_00778_),
    .A(\core.f2e_addr[7] ),
    .X(_00806_));
 sg13g2_a21oi_2 _06258_ (.B1(_00654_),
    .Y(_00807_),
    .A2(_00762_),
    .A1(_00755_));
 sg13g2_a21o_1 _06259_ (.A2(_00762_),
    .A1(_00755_),
    .B1(_00752_),
    .X(_00808_));
 sg13g2_or2_1 _06260_ (.X(_00809_),
    .B(_00808_),
    .A(_00065_));
 sg13g2_xor2_1 _06261_ (.B(_00809_),
    .A(_00064_),
    .X(_00810_));
 sg13g2_mux2_2 _06262_ (.A0(_00806_),
    .A1(_00810_),
    .S(net3357),
    .X(_00811_));
 sg13g2_and2_1 _06263_ (.A(_00661_),
    .B(_00811_),
    .X(_00812_));
 sg13g2_nand2b_2 _06264_ (.Y(_00813_),
    .B(\core.fetch.spi_reader.addr[7] ),
    .A_N(_00811_));
 sg13g2_xnor2_1 _06265_ (.Y(_00814_),
    .A(\core.f2e_addr[5] ),
    .B(_00775_));
 sg13g2_nand2_1 _06266_ (.Y(_00815_),
    .A(net3352),
    .B(_00814_));
 sg13g2_xnor2_1 _06267_ (.Y(_00816_),
    .A(_00069_),
    .B(_00807_));
 sg13g2_o21ai_1 _06268_ (.B1(_00815_),
    .Y(_00817_),
    .A1(net3352),
    .A2(_00816_));
 sg13g2_xnor2_1 _06269_ (.Y(_00818_),
    .A(_00068_),
    .B(_00817_));
 sg13g2_xor2_1 _06270_ (.B(_00774_),
    .A(\core.f2e_addr[3] ),
    .X(_00819_));
 sg13g2_nor2_1 _06271_ (.A(net3357),
    .B(_00819_),
    .Y(_00820_));
 sg13g2_a21oi_1 _06272_ (.A1(_00760_),
    .A2(_00761_),
    .Y(_00821_),
    .B1(_00754_));
 sg13g2_xnor2_1 _06273_ (.Y(_00822_),
    .A(_00653_),
    .B(_00821_));
 sg13g2_a21oi_2 _06274_ (.B1(_00820_),
    .Y(_00823_),
    .A2(_00822_),
    .A1(net3357));
 sg13g2_nor2_1 _06275_ (.A(_00658_),
    .B(_00823_),
    .Y(_00824_));
 sg13g2_nand2_1 _06276_ (.Y(_00825_),
    .A(_00658_),
    .B(_00823_));
 sg13g2_xnor2_1 _06277_ (.Y(_00826_),
    .A(_00757_),
    .B(_00759_));
 sg13g2_a21oi_1 _06278_ (.A1(_00581_),
    .A2(_00657_),
    .Y(_00827_),
    .B1(net3355));
 sg13g2_a22oi_1 _06279_ (.Y(_00828_),
    .B1(_00827_),
    .B2(_00772_),
    .A2(_00826_),
    .A1(net3355));
 sg13g2_or2_1 _06280_ (.X(_00829_),
    .B(_00828_),
    .A(\core.fetch.spi_reader.addr[1] ));
 sg13g2_nand2_1 _06281_ (.Y(_00830_),
    .A(_00649_),
    .B(_00652_));
 sg13g2_and2_1 _06282_ (.A(_00757_),
    .B(net3355),
    .X(_00831_));
 sg13g2_a22oi_1 _06283_ (.Y(_00832_),
    .B1(_00830_),
    .B2(_00831_),
    .A2(net3354),
    .A1(_00656_));
 sg13g2_nor2b_2 _06284_ (.A(_00061_),
    .B_N(_00832_),
    .Y(_00833_));
 sg13g2_xnor2_1 _06285_ (.Y(_00834_),
    .A(\core.fetch.spi_reader.addr[1] ),
    .B(_00828_));
 sg13g2_nor2_1 _06286_ (.A(_00833_),
    .B(_00834_),
    .Y(_00835_));
 sg13g2_or2_1 _06287_ (.X(_00836_),
    .B(_00834_),
    .A(_00833_));
 sg13g2_o21ai_1 _06288_ (.B1(_00829_),
    .Y(_00837_),
    .A1(_00833_),
    .A2(_00834_));
 sg13g2_xor2_1 _06289_ (.B(_00761_),
    .A(_00760_),
    .X(_00838_));
 sg13g2_o21ai_1 _06290_ (.B1(net3354),
    .Y(_00839_),
    .A1(_00772_),
    .A2(_00773_));
 sg13g2_a21oi_1 _06291_ (.A1(_00772_),
    .A2(_00773_),
    .Y(_00840_),
    .B1(_00839_));
 sg13g2_a21oi_2 _06292_ (.B1(_00840_),
    .Y(_00841_),
    .A2(_00838_),
    .A1(net3355));
 sg13g2_xnor2_1 _06293_ (.Y(_00842_),
    .A(_00063_),
    .B(_00841_));
 sg13g2_nor2_1 _06294_ (.A(\core.fetch.spi_reader.addr[2] ),
    .B(_00841_),
    .Y(_00843_));
 sg13g2_a221oi_1 _06295_ (.B2(_00842_),
    .C1(_00843_),
    .B1(_00837_),
    .A1(_00658_),
    .Y(_00844_),
    .A2(_00823_));
 sg13g2_or2_1 _06296_ (.X(_00845_),
    .B(_00844_),
    .A(_00824_));
 sg13g2_and3_1 _06297_ (.X(_00846_),
    .A(_00654_),
    .B(_00755_),
    .C(_00762_));
 sg13g2_nor3_2 _06298_ (.A(net3353),
    .B(_00807_),
    .C(_00846_),
    .Y(_00847_));
 sg13g2_or3_2 _06299_ (.A(net3353),
    .B(_00807_),
    .C(_00846_),
    .X(_00848_));
 sg13g2_a21oi_1 _06300_ (.A1(\core.f2e_addr[3] ),
    .A2(_00774_),
    .Y(_00849_),
    .B1(net3564));
 sg13g2_nor3_2 _06301_ (.A(net3356),
    .B(_00775_),
    .C(_00849_),
    .Y(_00850_));
 sg13g2_inv_1 _06302_ (.Y(_00851_),
    .A(_00850_));
 sg13g2_nor2_1 _06303_ (.A(_00847_),
    .B(_00850_),
    .Y(_00852_));
 sg13g2_nor3_1 _06304_ (.A(_00070_),
    .B(_00847_),
    .C(_00850_),
    .Y(_00853_));
 sg13g2_a21oi_1 _06305_ (.A1(_00848_),
    .A2(_00851_),
    .Y(_00854_),
    .B1(_00662_));
 sg13g2_nor2_1 _06306_ (.A(_00853_),
    .B(_00854_),
    .Y(_00855_));
 sg13g2_nor4_1 _06307_ (.A(_00824_),
    .B(_00844_),
    .C(_00853_),
    .D(_00854_),
    .Y(_00856_));
 sg13g2_nand2_1 _06308_ (.Y(_00857_),
    .A(_00818_),
    .B(_00855_));
 sg13g2_nand2_1 _06309_ (.Y(_00858_),
    .A(\core.fetch.spi_reader.addr[5] ),
    .B(_00817_));
 sg13g2_nor2_1 _06310_ (.A(\core.fetch.spi_reader.addr[4] ),
    .B(_00852_),
    .Y(_00859_));
 sg13g2_nor2_1 _06311_ (.A(\core.fetch.spi_reader.addr[5] ),
    .B(_00817_),
    .Y(_00860_));
 sg13g2_a221oi_1 _06312_ (.B2(_00859_),
    .C1(_00860_),
    .B1(_00858_),
    .A1(_00818_),
    .Y(_00861_),
    .A2(_00856_));
 sg13g2_a21oi_1 _06313_ (.A1(_00065_),
    .A2(_00808_),
    .Y(_00862_),
    .B1(net3352));
 sg13g2_a21oi_1 _06314_ (.A1(\core.f2e_addr[5] ),
    .A2(_00775_),
    .Y(_00863_),
    .B1(\core.f2e_addr[6] ));
 sg13g2_nor3_1 _06315_ (.A(net3356),
    .B(_00778_),
    .C(_00863_),
    .Y(_00864_));
 sg13g2_a21oi_2 _06316_ (.B1(_00864_),
    .Y(_00865_),
    .A2(_00862_),
    .A1(_00809_));
 sg13g2_xor2_1 _06317_ (.B(_00865_),
    .A(_00067_),
    .X(_00866_));
 sg13g2_nor2_1 _06318_ (.A(\core.fetch.spi_reader.addr[6] ),
    .B(_00865_),
    .Y(_00867_));
 sg13g2_a21oi_1 _06319_ (.A1(_00661_),
    .A2(_00811_),
    .Y(_00868_),
    .B1(_00867_));
 sg13g2_o21ai_1 _06320_ (.B1(_00868_),
    .Y(_00869_),
    .A1(_00861_),
    .A2(_00866_));
 sg13g2_and4_1 _06321_ (.A(_00799_),
    .B(_00804_),
    .C(_00813_),
    .D(_00869_),
    .X(_00870_));
 sg13g2_nor2_1 _06322_ (.A(\core.fetch.spi_reader.addr[8] ),
    .B(_00803_),
    .Y(_00871_));
 sg13g2_a21oi_1 _06323_ (.A1(_00798_),
    .A2(_00871_),
    .Y(_00872_),
    .B1(_00797_));
 sg13g2_nor2b_1 _06324_ (.A(_00870_),
    .B_N(_00872_),
    .Y(_00873_));
 sg13g2_nand3_1 _06325_ (.B(\core.fetch.rd_addr_i[8] ),
    .C(_00763_),
    .A(\core.fetch.rd_addr_i[9] ),
    .Y(_00874_));
 sg13g2_nor2_1 _06326_ (.A(_00080_),
    .B(_00874_),
    .Y(_00875_));
 sg13g2_and2_1 _06327_ (.A(_00078_),
    .B(_00782_),
    .X(_00876_));
 sg13g2_nor2_1 _06328_ (.A(_00078_),
    .B(_00782_),
    .Y(_00877_));
 sg13g2_o21ai_1 _06329_ (.B1(net3352),
    .Y(_00878_),
    .A1(_00876_),
    .A2(_00877_));
 sg13g2_xnor2_1 _06330_ (.Y(_00879_),
    .A(_00079_),
    .B(_00875_));
 sg13g2_o21ai_1 _06331_ (.B1(_00878_),
    .Y(_00880_),
    .A1(net3352),
    .A2(_00879_));
 sg13g2_nand2_1 _06332_ (.Y(_00881_),
    .A(net3568),
    .B(_00880_));
 sg13g2_nor2_1 _06333_ (.A(net3568),
    .B(_00880_),
    .Y(_00882_));
 sg13g2_xor2_1 _06334_ (.B(_00880_),
    .A(net3568),
    .X(_00883_));
 sg13g2_xnor2_1 _06335_ (.Y(_00884_),
    .A(_00665_),
    .B(_00874_));
 sg13g2_a21oi_1 _06336_ (.A1(_00663_),
    .A2(_00780_),
    .Y(_00885_),
    .B1(net3356));
 sg13g2_a22oi_1 _06337_ (.Y(_00886_),
    .B1(_00885_),
    .B2(_00782_),
    .A2(_00884_),
    .A1(net3356));
 sg13g2_xnor2_1 _06338_ (.Y(_00887_),
    .A(_00081_),
    .B(_00886_));
 sg13g2_nand2_1 _06339_ (.Y(_00888_),
    .A(_00883_),
    .B(_00887_));
 sg13g2_nor2_1 _06340_ (.A(\core.fetch.spi_reader.addr[10] ),
    .B(_00886_),
    .Y(_00889_));
 sg13g2_o21ai_1 _06341_ (.B1(_00881_),
    .Y(_00890_),
    .A1(_00882_),
    .A2(_00889_));
 sg13g2_o21ai_1 _06342_ (.B1(_00890_),
    .Y(_00891_),
    .A1(_00873_),
    .A2(_00888_));
 sg13g2_nor3_1 _06343_ (.A(_00075_),
    .B(_00779_),
    .C(_00785_),
    .Y(_00892_));
 sg13g2_xnor2_1 _06344_ (.Y(_00893_),
    .A(_00073_),
    .B(_00767_));
 sg13g2_xnor2_1 _06345_ (.Y(_00894_),
    .A(\core.f2e_addr[14] ),
    .B(_00892_));
 sg13g2_mux2_2 _06346_ (.A0(_00893_),
    .A1(_00894_),
    .S(net3352),
    .X(_00895_));
 sg13g2_nor2b_1 _06347_ (.A(_00074_),
    .B_N(_00895_),
    .Y(_00896_));
 sg13g2_xnor2_1 _06348_ (.Y(_00897_),
    .A(_00074_),
    .B(_00895_));
 sg13g2_inv_1 _06349_ (.Y(_00898_),
    .A(_00897_));
 sg13g2_or2_1 _06350_ (.X(_00899_),
    .B(_00895_),
    .A(\core.fetch.spi_reader.addr[14] ));
 sg13g2_nand2_1 _06351_ (.Y(_00900_),
    .A(_00898_),
    .B(_00899_));
 sg13g2_xor2_1 _06352_ (.B(_00764_),
    .A(_00076_),
    .X(_00901_));
 sg13g2_o21ai_1 _06353_ (.B1(_00075_),
    .Y(_00902_),
    .A1(_00779_),
    .A2(_00785_));
 sg13g2_nor2b_1 _06354_ (.A(_00892_),
    .B_N(_00902_),
    .Y(_00903_));
 sg13g2_mux2_2 _06355_ (.A0(_00901_),
    .A1(_00903_),
    .S(net3352),
    .X(_00904_));
 sg13g2_nand2b_1 _06356_ (.Y(_00905_),
    .B(_00904_),
    .A_N(\core.fetch.spi_reader.addr[13] ));
 sg13g2_nand2b_1 _06357_ (.Y(_00906_),
    .B(\core.fetch.spi_reader.addr[13] ),
    .A_N(_00904_));
 sg13g2_and2_1 _06358_ (.A(_00905_),
    .B(_00906_),
    .X(_00907_));
 sg13g2_a21o_1 _06359_ (.A2(_00763_),
    .A1(_00750_),
    .B1(net3525),
    .X(_00908_));
 sg13g2_a21o_1 _06360_ (.A2(_00908_),
    .A1(_00764_),
    .B1(net3352),
    .X(_00909_));
 sg13g2_xor2_1 _06361_ (.B(_00877_),
    .A(\core.f2e_addr[12] ),
    .X(_00910_));
 sg13g2_o21ai_1 _06362_ (.B1(_00909_),
    .Y(_00911_),
    .A1(net3356),
    .A2(_00910_));
 sg13g2_nor2_1 _06363_ (.A(\core.fetch.spi_reader.addr[12] ),
    .B(_00911_),
    .Y(_00912_));
 sg13g2_nand2_1 _06364_ (.Y(_00913_),
    .A(_00907_),
    .B(_00912_));
 sg13g2_and2_1 _06365_ (.A(_00905_),
    .B(_00913_),
    .X(_00914_));
 sg13g2_inv_1 _06366_ (.Y(_00915_),
    .A(_00914_));
 sg13g2_o21ai_1 _06367_ (.B1(_00899_),
    .Y(_00916_),
    .A1(_00898_),
    .A2(_00914_));
 sg13g2_xnor2_1 _06368_ (.Y(_00917_),
    .A(_00077_),
    .B(_00911_));
 sg13g2_or2_1 _06369_ (.X(_00918_),
    .B(_00912_),
    .A(_00907_));
 sg13g2_xor2_1 _06370_ (.B(_00887_),
    .A(_00873_),
    .X(_00919_));
 sg13g2_xnor2_1 _06371_ (.Y(_00920_),
    .A(_00799_),
    .B(_00871_));
 sg13g2_a21oi_1 _06372_ (.A1(_00813_),
    .A2(_00869_),
    .Y(_00921_),
    .B1(_00804_));
 sg13g2_a21o_1 _06373_ (.A2(_00921_),
    .A1(_00920_),
    .B1(_00870_),
    .X(_00922_));
 sg13g2_nor2_1 _06374_ (.A(_00887_),
    .B(_00889_),
    .Y(_00923_));
 sg13g2_xor2_1 _06375_ (.B(_00923_),
    .A(_00883_),
    .X(_00924_));
 sg13g2_xor2_1 _06376_ (.B(_00866_),
    .A(_00861_),
    .X(_00925_));
 sg13g2_nand2b_2 _06377_ (.Y(_00926_),
    .B(_00813_),
    .A_N(_00812_));
 sg13g2_o21ai_1 _06378_ (.B1(_00866_),
    .Y(_00927_),
    .A1(\core.fetch.spi_reader.addr[6] ),
    .A2(_00865_));
 sg13g2_xnor2_1 _06379_ (.Y(_00928_),
    .A(_00926_),
    .B(_00927_));
 sg13g2_xor2_1 _06380_ (.B(_00855_),
    .A(_00845_),
    .X(_00929_));
 sg13g2_nor2_1 _06381_ (.A(_00855_),
    .B(_00859_),
    .Y(_00930_));
 sg13g2_nor2b_1 _06382_ (.A(_00824_),
    .B_N(_00825_),
    .Y(_00931_));
 sg13g2_nor2_1 _06383_ (.A(_00842_),
    .B(_00843_),
    .Y(_00932_));
 sg13g2_xnor2_1 _06384_ (.Y(_00933_),
    .A(_00837_),
    .B(_00842_));
 sg13g2_and2_1 _06385_ (.A(\core.fetch.spi_reader.dirty ),
    .B(_00933_),
    .X(_00934_));
 sg13g2_o21ai_1 _06386_ (.B1(_00934_),
    .Y(_00935_),
    .A1(_00931_),
    .A2(_00932_));
 sg13g2_a21oi_1 _06387_ (.A1(_00931_),
    .A2(_00932_),
    .Y(_00936_),
    .B1(_00935_));
 sg13g2_xor2_1 _06388_ (.B(_00930_),
    .A(_00818_),
    .X(_00937_));
 sg13g2_nand3_1 _06389_ (.B(_00936_),
    .C(_00937_),
    .A(_00929_),
    .Y(_00938_));
 sg13g2_nand2_1 _06390_ (.Y(_00939_),
    .A(_00907_),
    .B(_00917_));
 sg13g2_inv_1 _06391_ (.Y(_00940_),
    .A(_00939_));
 sg13g2_and2_1 _06392_ (.A(_00842_),
    .B(_00931_),
    .X(_00941_));
 sg13g2_nor2b_1 _06393_ (.A(_00832_),
    .B_N(_00061_),
    .Y(_00942_));
 sg13g2_nor2_1 _06394_ (.A(_00836_),
    .B(_00942_),
    .Y(_00943_));
 sg13g2_o21ai_1 _06395_ (.B1(_00837_),
    .Y(_00944_),
    .A1(_00836_),
    .A2(_00942_));
 sg13g2_a21o_1 _06396_ (.A2(_00841_),
    .A1(\core.fetch.spi_reader.addr[2] ),
    .B1(_00824_),
    .X(_00945_));
 sg13g2_a22oi_1 _06397_ (.Y(_00946_),
    .B1(_00945_),
    .B2(_00825_),
    .A2(_00944_),
    .A1(_00941_));
 sg13g2_nor4_1 _06398_ (.A(_00857_),
    .B(_00866_),
    .C(_00926_),
    .D(_00946_),
    .Y(_00947_));
 sg13g2_nand2_1 _06399_ (.Y(_00948_),
    .A(\core.fetch.spi_reader.addr[6] ),
    .B(_00865_));
 sg13g2_a21oi_1 _06400_ (.A1(_00813_),
    .A2(_00948_),
    .Y(_00949_),
    .B1(_00812_));
 sg13g2_a22oi_1 _06401_ (.Y(_00950_),
    .B1(_00852_),
    .B2(\core.fetch.spi_reader.addr[4] ),
    .A2(_00817_),
    .A1(\core.fetch.spi_reader.addr[5] ));
 sg13g2_nor4_1 _06402_ (.A(_00860_),
    .B(_00866_),
    .C(_00926_),
    .D(_00950_),
    .Y(_00951_));
 sg13g2_or3_1 _06403_ (.A(_00947_),
    .B(_00949_),
    .C(_00951_),
    .X(_00952_));
 sg13g2_nand2_1 _06404_ (.Y(_00953_),
    .A(_00791_),
    .B(_00897_));
 sg13g2_nand4_1 _06405_ (.B(_00897_),
    .C(_00907_),
    .A(_00791_),
    .Y(_00954_),
    .D(_00917_));
 sg13g2_inv_1 _06406_ (.Y(_00955_),
    .A(_00954_));
 sg13g2_nand3_1 _06407_ (.B(_00905_),
    .C(_00911_),
    .A(\core.fetch.spi_reader.addr[12] ),
    .Y(_00956_));
 sg13g2_a21oi_1 _06408_ (.A1(_00906_),
    .A2(_00956_),
    .Y(_00957_),
    .B1(_00953_));
 sg13g2_a221oi_1 _06409_ (.B2(_00896_),
    .C1(_00957_),
    .B1(_00791_),
    .A1(\core.fetch.spi_reader.addr[15] ),
    .Y(_00958_),
    .A2(_00789_));
 sg13g2_nand2_1 _06410_ (.Y(_00959_),
    .A(\core.fetch.spi_reader.addr[8] ),
    .B(_00803_));
 sg13g2_a21o_1 _06411_ (.A2(_00959_),
    .A1(_00798_),
    .B1(_00797_),
    .X(_00960_));
 sg13g2_a22oi_1 _06412_ (.Y(_00961_),
    .B1(_00886_),
    .B2(\core.fetch.spi_reader.addr[10] ),
    .A2(_00880_),
    .A1(net3568));
 sg13g2_or2_1 _06413_ (.X(_00962_),
    .B(_00961_),
    .A(_00882_));
 sg13g2_o21ai_1 _06414_ (.B1(_00962_),
    .Y(_00963_),
    .A1(_00888_),
    .A2(_00960_));
 sg13g2_nor3_2 _06415_ (.A(_00805_),
    .B(_00888_),
    .C(_00954_),
    .Y(_00964_));
 sg13g2_a22oi_1 _06416_ (.Y(_00965_),
    .B1(_00964_),
    .B2(_00952_),
    .A2(_00963_),
    .A1(_00955_));
 sg13g2_nand2_1 _06417_ (.Y(_00966_),
    .A(_00941_),
    .B(_00943_));
 sg13g2_nor4_2 _06418_ (.A(_00857_),
    .B(_00866_),
    .C(_00926_),
    .Y(_00967_),
    .D(_00966_));
 sg13g2_a22oi_1 _06419_ (.Y(_00968_),
    .B1(_00967_),
    .B2(_00964_),
    .A2(_00965_),
    .A1(_00958_));
 sg13g2_a21oi_1 _06420_ (.A1(_00891_),
    .A2(_00940_),
    .Y(_00969_),
    .B1(_00915_));
 sg13g2_xnor2_1 _06421_ (.Y(_00970_),
    .A(_00897_),
    .B(_00969_));
 sg13g2_a221oi_1 _06422_ (.B2(_00891_),
    .C1(_00790_),
    .B1(_00955_),
    .A1(_00791_),
    .Y(_00971_),
    .A2(_00916_));
 sg13g2_a21o_1 _06423_ (.A2(_00918_),
    .A1(_00913_),
    .B1(_00917_),
    .X(_00972_));
 sg13g2_mux2_1 _06424_ (.A0(_00972_),
    .A1(_00939_),
    .S(_00891_),
    .X(_00973_));
 sg13g2_xor2_1 _06425_ (.B(_00900_),
    .A(_00791_),
    .X(_00974_));
 sg13g2_nor4_1 _06426_ (.A(_00925_),
    .B(_00928_),
    .C(_00938_),
    .D(_00974_),
    .Y(_00975_));
 sg13g2_nand4_1 _06427_ (.B(_00922_),
    .C(_00924_),
    .A(_00919_),
    .Y(_00976_),
    .D(_00975_));
 sg13g2_or4_1 _06428_ (.A(_00968_),
    .B(_00971_),
    .C(_00973_),
    .D(_00976_),
    .X(_00977_));
 sg13g2_nor2_1 _06429_ (.A(_00970_),
    .B(_00977_),
    .Y(_00978_));
 sg13g2_o21ai_1 _06430_ (.B1(net3565),
    .Y(_00979_),
    .A1(_00970_),
    .A2(_00977_));
 sg13g2_nor3_2 _06431_ (.A(\core.fetch.spi_reader.state[0] ),
    .B(net3567),
    .C(_00633_),
    .Y(_00980_));
 sg13g2_or3_1 _06432_ (.A(\core.fetch.spi_reader.state[0] ),
    .B(net3567),
    .C(_00633_),
    .X(_00981_));
 sg13g2_or3_1 _06433_ (.A(\core.fetch.spi_reader.counter[3] ),
    .B(\core.fetch.spi_reader.counter[2] ),
    .C(\core.fetch.spi_reader.counter[4] ),
    .X(_00982_));
 sg13g2_nor2_1 _06434_ (.A(\core.fetch.spi_reader.counter[1] ),
    .B(\core.fetch.spi_reader.counter[0] ),
    .Y(_00983_));
 sg13g2_nor4_2 _06435_ (.A(\core.fetch.spi_reader.counter[1] ),
    .B(\core.fetch.spi_reader.counter[0] ),
    .C(\core.fetch.spi_reader.counter[5] ),
    .Y(_00984_),
    .D(_00982_));
 sg13g2_and2_2 _06436_ (.A(net3210),
    .B(_00984_),
    .X(_00985_));
 sg13g2_nand2_2 _06437_ (.Y(_00986_),
    .A(net3208),
    .B(_00984_));
 sg13g2_nor2_1 _06438_ (.A(_00019_),
    .B(net3206),
    .Y(_00987_));
 sg13g2_nand2_2 _06439_ (.Y(_00988_),
    .A(\core.fetch.spi_reader.state[1] ),
    .B(\core.fetch.spi_reader.state[2] ));
 sg13g2_nor2_2 _06440_ (.A(_00985_),
    .B(_00987_),
    .Y(_00989_));
 sg13g2_inv_1 _06441_ (.Y(_00990_),
    .A(_00989_));
 sg13g2_nand2_1 _06442_ (.Y(_00991_),
    .A(_00988_),
    .B(_00989_));
 sg13g2_and2_2 _06443_ (.A(net3567),
    .B(_00747_),
    .X(_00992_));
 sg13g2_nand2_2 _06444_ (.Y(_00993_),
    .A(net3567),
    .B(_00747_));
 sg13g2_nand2_1 _06445_ (.Y(_00994_),
    .A(\core.fetch.spi_reader.state[0] ),
    .B(_00988_));
 sg13g2_a21oi_1 _06446_ (.A1(_00993_),
    .A2(_00994_),
    .Y(_00995_),
    .B1(net3362));
 sg13g2_or3_1 _06447_ (.A(net867),
    .B(_00991_),
    .C(_00995_),
    .X(_00996_));
 sg13g2_nor2_1 _06448_ (.A(uio_out[0]),
    .B(_00987_),
    .Y(_00997_));
 sg13g2_a21o_1 _06449_ (.A2(_00979_),
    .A1(_00748_),
    .B1(_00996_),
    .X(_00000_));
 sg13g2_nor2_2 _06450_ (.A(\core.lsu.spi.state[1] ),
    .B(\core.lsu.spi.state[0] ),
    .Y(_00998_));
 sg13g2_inv_1 _06451_ (.Y(_00999_),
    .A(_00998_));
 sg13g2_nand2_2 _06452_ (.Y(_01000_),
    .A(_00084_),
    .B(_00998_));
 sg13g2_nor2_1 _06453_ (.A(_00018_),
    .B(_01000_),
    .Y(_01001_));
 sg13g2_nor3_1 _06454_ (.A(net615),
    .B(uio_out[4]),
    .C(_01000_),
    .Y(_01002_));
 sg13g2_nand2_1 _06455_ (.Y(_01003_),
    .A(\core.lsu.write_index[2] ),
    .B(\core.fetch.rd_addr_i[2] ));
 sg13g2_nor2_1 _06456_ (.A(_00066_),
    .B(_01003_),
    .Y(_01004_));
 sg13g2_and2_1 _06457_ (.A(\core.lsu.write_index[1] ),
    .B(net3526),
    .X(_01005_));
 sg13g2_and2_1 _06458_ (.A(\core.lsu.write_index[0] ),
    .B(\core.fetch.rd_addr_i[0] ),
    .X(_01006_));
 sg13g2_xor2_1 _06459_ (.B(net3526),
    .A(\core.lsu.write_index[1] ),
    .X(_01007_));
 sg13g2_a21oi_2 _06460_ (.B1(_01005_),
    .Y(_01008_),
    .A2(_01007_),
    .A1(_01006_));
 sg13g2_xnor2_1 _06461_ (.Y(_01009_),
    .A(\core.lsu.write_index[2] ),
    .B(\core.fetch.rd_addr_i[2] ));
 sg13g2_nor3_1 _06462_ (.A(_00653_),
    .B(_01008_),
    .C(_01009_),
    .Y(_01010_));
 sg13g2_nor2_2 _06463_ (.A(_01004_),
    .B(_01010_),
    .Y(_01011_));
 sg13g2_nor3_2 _06464_ (.A(_00751_),
    .B(_00753_),
    .C(_01011_),
    .Y(_01012_));
 sg13g2_nand2_1 _06465_ (.Y(_01013_),
    .A(\core.fetch.rd_addr_i[12] ),
    .B(_01012_));
 sg13g2_nand3_1 _06466_ (.B(net3525),
    .C(_01012_),
    .A(\core.fetch.rd_addr_i[13] ),
    .Y(_01014_));
 sg13g2_nor2_1 _06467_ (.A(_00073_),
    .B(_01014_),
    .Y(_01015_));
 sg13g2_xor2_1 _06468_ (.B(_01014_),
    .A(_00073_),
    .X(_01016_));
 sg13g2_xor2_1 _06469_ (.B(_01016_),
    .A(_00091_),
    .X(_01017_));
 sg13g2_xor2_1 _06470_ (.B(_01013_),
    .A(_00076_),
    .X(_01018_));
 sg13g2_xnor2_1 _06471_ (.Y(_01019_),
    .A(_00672_),
    .B(_01018_));
 sg13g2_xnor2_1 _06472_ (.Y(_01020_),
    .A(net3525),
    .B(_01012_));
 sg13g2_xor2_1 _06473_ (.B(_01020_),
    .A(_00092_),
    .X(_01021_));
 sg13g2_nor2_1 _06474_ (.A(_01019_),
    .B(_01021_),
    .Y(_01022_));
 sg13g2_nor3_2 _06475_ (.A(_00655_),
    .B(_00753_),
    .C(_01011_),
    .Y(_01023_));
 sg13g2_nand3_1 _06476_ (.B(_00665_),
    .C(_01023_),
    .A(\core.fetch.rd_addr_i[9] ),
    .Y(_01024_));
 sg13g2_xor2_1 _06477_ (.B(_01024_),
    .A(_00079_),
    .X(_01025_));
 sg13g2_nand2b_1 _06478_ (.Y(_01026_),
    .B(\core.lsu.spi.addr[11] ),
    .A_N(_01025_));
 sg13g2_nor2b_1 _06479_ (.A(\core.lsu.spi.addr[11] ),
    .B_N(_01025_),
    .Y(_01027_));
 sg13g2_xnor2_1 _06480_ (.Y(_01028_),
    .A(\core.lsu.spi.addr[11] ),
    .B(_01025_));
 sg13g2_a21o_1 _06481_ (.A2(_01023_),
    .A1(\core.fetch.rd_addr_i[9] ),
    .B1(_00665_),
    .X(_01029_));
 sg13g2_and2_1 _06482_ (.A(_01024_),
    .B(_01029_),
    .X(_01030_));
 sg13g2_xnor2_1 _06483_ (.Y(_01031_),
    .A(_00674_),
    .B(_01030_));
 sg13g2_nand2_1 _06484_ (.Y(_01032_),
    .A(_01028_),
    .B(_01031_));
 sg13g2_xnor2_1 _06485_ (.Y(_01033_),
    .A(_00082_),
    .B(_01023_));
 sg13g2_xor2_1 _06486_ (.B(_01033_),
    .A(_00094_),
    .X(_01034_));
 sg13g2_o21ai_1 _06487_ (.B1(_00655_),
    .Y(_01035_),
    .A1(_00753_),
    .A2(_01011_));
 sg13g2_nand2b_2 _06488_ (.Y(_01036_),
    .B(_01035_),
    .A_N(_01023_));
 sg13g2_xor2_1 _06489_ (.B(_01036_),
    .A(_00095_),
    .X(_01037_));
 sg13g2_nand2b_1 _06490_ (.Y(_01038_),
    .B(_01034_),
    .A_N(_01037_));
 sg13g2_o21ai_1 _06491_ (.B1(\core.fetch.rd_addr_i[4] ),
    .Y(_01039_),
    .A1(_01004_),
    .A2(_01010_));
 sg13g2_nor3_2 _06492_ (.A(_00065_),
    .B(_00752_),
    .C(_01011_),
    .Y(_01040_));
 sg13g2_xor2_1 _06493_ (.B(_01040_),
    .A(_00064_),
    .X(_01041_));
 sg13g2_nor2_1 _06494_ (.A(\core.lsu.spi.addr[7] ),
    .B(_01041_),
    .Y(_01042_));
 sg13g2_and2_1 _06495_ (.A(net3520),
    .B(_01041_),
    .X(_01043_));
 sg13g2_xor2_1 _06496_ (.B(_01039_),
    .A(_00069_),
    .X(_01044_));
 sg13g2_xnor2_1 _06497_ (.Y(_01045_),
    .A(_00088_),
    .B(_01044_));
 sg13g2_xnor2_1 _06498_ (.Y(_01046_),
    .A(\core.fetch.rd_addr_i[4] ),
    .B(_01011_));
 sg13g2_xnor2_1 _06499_ (.Y(_01047_),
    .A(_00089_),
    .B(_01046_));
 sg13g2_or2_1 _06500_ (.X(_01048_),
    .B(_01047_),
    .A(_01045_));
 sg13g2_o21ai_1 _06501_ (.B1(_01003_),
    .Y(_01049_),
    .A1(_01008_),
    .A2(_01009_));
 sg13g2_xnor2_1 _06502_ (.Y(_01050_),
    .A(_00653_),
    .B(_01049_));
 sg13g2_nor2b_1 _06503_ (.A(\core.lsu.spi.addr[3] ),
    .B_N(_01050_),
    .Y(_01051_));
 sg13g2_nand2b_1 _06504_ (.Y(_01052_),
    .B(\core.lsu.spi.addr[3] ),
    .A_N(_01050_));
 sg13g2_xor2_1 _06505_ (.B(_01007_),
    .A(_01006_),
    .X(_01053_));
 sg13g2_nor2b_1 _06506_ (.A(\core.lsu.spi.addr[1] ),
    .B_N(_01053_),
    .Y(_01054_));
 sg13g2_xor2_1 _06507_ (.B(\core.fetch.rd_addr_i[0] ),
    .A(\core.lsu.write_index[0] ),
    .X(_01055_));
 sg13g2_or2_1 _06508_ (.X(_01056_),
    .B(_01055_),
    .A(_00085_));
 sg13g2_xnor2_1 _06509_ (.Y(_01057_),
    .A(\core.lsu.spi.addr[1] ),
    .B(_01053_));
 sg13g2_a21oi_1 _06510_ (.A1(_01056_),
    .A2(_01057_),
    .Y(_01058_),
    .B1(_01054_));
 sg13g2_xnor2_1 _06511_ (.Y(_01059_),
    .A(_01008_),
    .B(_01009_));
 sg13g2_xor2_1 _06512_ (.B(_01059_),
    .A(_00086_),
    .X(_01060_));
 sg13g2_or2_1 _06513_ (.X(_01061_),
    .B(_01059_),
    .A(\core.lsu.spi.addr[2] ));
 sg13g2_o21ai_1 _06514_ (.B1(_01061_),
    .Y(_01062_),
    .A1(_01058_),
    .A2(_01060_));
 sg13g2_a21oi_1 _06515_ (.A1(_01052_),
    .A2(_01062_),
    .Y(_01063_),
    .B1(_01051_));
 sg13g2_nor3_1 _06516_ (.A(_01045_),
    .B(_01047_),
    .C(_01063_),
    .Y(_01064_));
 sg13g2_or2_1 _06517_ (.X(_01065_),
    .B(_01063_),
    .A(_01048_));
 sg13g2_nand2b_1 _06518_ (.Y(_01066_),
    .B(_01044_),
    .A_N(\core.lsu.spi.addr[5] ));
 sg13g2_nand2b_1 _06519_ (.Y(_01067_),
    .B(_01046_),
    .A_N(\core.lsu.spi.addr[4] ));
 sg13g2_o21ai_1 _06520_ (.B1(_01066_),
    .Y(_01068_),
    .A1(_01045_),
    .A2(_01067_));
 sg13g2_nor2_1 _06521_ (.A(_01064_),
    .B(_01068_),
    .Y(_01069_));
 sg13g2_o21ai_1 _06522_ (.B1(_00065_),
    .Y(_01070_),
    .A1(_00752_),
    .A2(_01011_));
 sg13g2_nor2b_2 _06523_ (.A(_01040_),
    .B_N(_01070_),
    .Y(_01071_));
 sg13g2_xor2_1 _06524_ (.B(_01071_),
    .A(_00087_),
    .X(_01072_));
 sg13g2_o21ai_1 _06525_ (.B1(_01072_),
    .Y(_01073_),
    .A1(_01064_),
    .A2(_01068_));
 sg13g2_and2_1 _06526_ (.A(_00667_),
    .B(_01071_),
    .X(_01074_));
 sg13g2_nor2_1 _06527_ (.A(_01042_),
    .B(_01074_),
    .Y(_01075_));
 sg13g2_a21o_1 _06528_ (.A2(_01075_),
    .A1(_01073_),
    .B1(_01043_),
    .X(_01076_));
 sg13g2_a221oi_1 _06529_ (.B2(_01075_),
    .C1(_01038_),
    .B1(_01073_),
    .A1(net3520),
    .Y(_01077_),
    .A2(_01041_));
 sg13g2_nor2_1 _06530_ (.A(\core.lsu.spi.addr[8] ),
    .B(_01036_),
    .Y(_01078_));
 sg13g2_a22oi_1 _06531_ (.Y(_01079_),
    .B1(_01034_),
    .B2(_01078_),
    .A2(_01033_),
    .A1(_00675_));
 sg13g2_nor2b_1 _06532_ (.A(_01077_),
    .B_N(_01079_),
    .Y(_01080_));
 sg13g2_and2_1 _06533_ (.A(_00673_),
    .B(_01030_),
    .X(_01081_));
 sg13g2_o21ai_1 _06534_ (.B1(_01026_),
    .Y(_01082_),
    .A1(_01027_),
    .A2(_01081_));
 sg13g2_o21ai_1 _06535_ (.B1(_01082_),
    .Y(_01083_),
    .A1(_01032_),
    .A2(_01080_));
 sg13g2_nand2_1 _06536_ (.Y(_01084_),
    .A(_01022_),
    .B(_01083_));
 sg13g2_nor2_1 _06537_ (.A(\core.lsu.spi.addr[12] ),
    .B(_01020_),
    .Y(_01085_));
 sg13g2_nor2b_1 _06538_ (.A(_01019_),
    .B_N(_01085_),
    .Y(_01086_));
 sg13g2_a21oi_1 _06539_ (.A1(_00672_),
    .A2(_01018_),
    .Y(_01087_),
    .B1(_01086_));
 sg13g2_a21o_1 _06540_ (.A2(_01087_),
    .A1(_01084_),
    .B1(_01017_),
    .X(_01088_));
 sg13g2_nand2_1 _06541_ (.Y(_01089_),
    .A(_01017_),
    .B(_01087_));
 sg13g2_xor2_1 _06542_ (.B(_01085_),
    .A(_01019_),
    .X(_01090_));
 sg13g2_nand3_1 _06543_ (.B(_01089_),
    .C(_01090_),
    .A(_01021_),
    .Y(_01091_));
 sg13g2_o21ai_1 _06544_ (.B1(_01084_),
    .Y(_01092_),
    .A1(_01083_),
    .A2(_01091_));
 sg13g2_nand2_1 _06545_ (.Y(_01093_),
    .A(_01031_),
    .B(_01079_));
 sg13g2_xnor2_1 _06546_ (.Y(_01094_),
    .A(_01034_),
    .B(_01078_));
 sg13g2_nor2_1 _06547_ (.A(_01031_),
    .B(_01081_),
    .Y(_01095_));
 sg13g2_nor2_1 _06548_ (.A(_01028_),
    .B(_01095_),
    .Y(_01096_));
 sg13g2_xnor2_1 _06549_ (.Y(_01097_),
    .A(_01045_),
    .B(_01067_));
 sg13g2_nand3_1 _06550_ (.B(_01063_),
    .C(_01097_),
    .A(_01047_),
    .Y(_01098_));
 sg13g2_a221oi_1 _06551_ (.B2(_01065_),
    .C1(_01096_),
    .B1(_01098_),
    .A1(_01028_),
    .Y(_01099_),
    .A2(_01095_));
 sg13g2_xnor2_1 _06552_ (.Y(_01100_),
    .A(_00072_),
    .B(_01015_));
 sg13g2_xnor2_1 _06553_ (.Y(_01101_),
    .A(_00090_),
    .B(_01100_));
 sg13g2_a21oi_1 _06554_ (.A1(_00671_),
    .A2(_01016_),
    .Y(_01102_),
    .B1(_01017_));
 sg13g2_xor2_1 _06555_ (.B(_01041_),
    .A(net3520),
    .X(_01103_));
 sg13g2_inv_1 _06556_ (.Y(_01104_),
    .A(_01103_));
 sg13g2_nor3_1 _06557_ (.A(_01072_),
    .B(_01074_),
    .C(_01104_),
    .Y(_01105_));
 sg13g2_nand2b_1 _06558_ (.Y(_01106_),
    .B(_01052_),
    .A_N(_01051_));
 sg13g2_nand2_1 _06559_ (.Y(_01107_),
    .A(_01060_),
    .B(_01061_));
 sg13g2_nand2b_1 _06560_ (.Y(_01108_),
    .B(\core.gpio.stray_wr_i ),
    .A_N(\core.lsu.spi.iswr ));
 sg13g2_nand2b_1 _06561_ (.Y(_01109_),
    .B(\core.lsu.spi.iswr ),
    .A_N(\core.gpio.stray_wr_i ));
 sg13g2_and2_1 _06562_ (.A(\core.lsu.spi.dirty ),
    .B(_01109_),
    .X(_01110_));
 sg13g2_xnor2_1 _06563_ (.Y(_01111_),
    .A(_01058_),
    .B(_01060_));
 sg13g2_nand3_1 _06564_ (.B(_01110_),
    .C(_01111_),
    .A(_01108_),
    .Y(_01112_));
 sg13g2_xnor2_1 _06565_ (.Y(_01113_),
    .A(_01106_),
    .B(_01107_));
 sg13g2_o21ai_1 _06566_ (.B1(_01104_),
    .Y(_01114_),
    .A1(_01072_),
    .A2(_01074_));
 sg13g2_o21ai_1 _06567_ (.B1(_01114_),
    .Y(_01115_),
    .A1(_00090_),
    .A2(_01100_));
 sg13g2_nor4_1 _06568_ (.A(_01105_),
    .B(_01112_),
    .C(_01113_),
    .D(_01115_),
    .Y(_01116_));
 sg13g2_xor2_1 _06569_ (.B(_01072_),
    .A(_01069_),
    .X(_01117_));
 sg13g2_nand4_1 _06570_ (.B(_01076_),
    .C(_01093_),
    .A(_01037_),
    .Y(_01118_),
    .D(_01094_));
 sg13g2_nand2b_1 _06571_ (.Y(_01119_),
    .B(_01118_),
    .A_N(_01077_));
 sg13g2_a21oi_1 _06572_ (.A1(_01076_),
    .A2(_01079_),
    .Y(_01120_),
    .B1(_01031_));
 sg13g2_xor2_1 _06573_ (.B(_01102_),
    .A(_01101_),
    .X(_01121_));
 sg13g2_nand3_1 _06574_ (.B(_01116_),
    .C(_01117_),
    .A(_01099_),
    .Y(_01122_));
 sg13g2_nor3_1 _06575_ (.A(_01120_),
    .B(_01121_),
    .C(_01122_),
    .Y(_01123_));
 sg13g2_nand4_1 _06576_ (.B(_01092_),
    .C(_01119_),
    .A(_01088_),
    .Y(_01124_),
    .D(_01123_));
 sg13g2_nand2_1 _06577_ (.Y(_00002_),
    .A(net616),
    .B(_01124_));
 sg13g2_nor2_2 _06578_ (.A(\core.lsu.state[0] ),
    .B(\core.lsu.state[1] ),
    .Y(_01125_));
 sg13g2_nand2_2 _06579_ (.Y(_01126_),
    .A(_00021_),
    .B(_01125_));
 sg13g2_nand2_1 _06580_ (.Y(_01127_),
    .A(net3501),
    .B(net3502));
 sg13g2_nor3_2 _06581_ (.A(net730),
    .B(\core.lsu.accept ),
    .C(_01127_),
    .Y(_01128_));
 sg13g2_nor2b_2 _06582_ (.A(_01126_),
    .B_N(net731),
    .Y(_00001_));
 sg13g2_nand2_1 _06583_ (.Y(_01129_),
    .A(_00631_),
    .B(net3355));
 sg13g2_nor2_1 _06584_ (.A(\core.fetch.data_size[0] ),
    .B(net3576),
    .Y(_01130_));
 sg13g2_nor2b_1 _06585_ (.A(net3524),
    .B_N(\core.lsu.is_half ),
    .Y(_01131_));
 sg13g2_nor2_1 _06586_ (.A(net3524),
    .B(\core.lsu.is_half ),
    .Y(_01132_));
 sg13g2_xnor2_1 _06587_ (.Y(_01133_),
    .A(_00650_),
    .B(_01131_));
 sg13g2_xor2_1 _06588_ (.B(_01130_),
    .A(\core.fetch.data_size[2] ),
    .X(_01134_));
 sg13g2_xor2_1 _06589_ (.B(net3524),
    .A(net3577),
    .X(_01135_));
 sg13g2_nor3_2 _06590_ (.A(_01133_),
    .B(_01134_),
    .C(_01135_),
    .Y(_01136_));
 sg13g2_nor2_1 _06591_ (.A(_01129_),
    .B(_01136_),
    .Y(_01137_));
 sg13g2_nor2_2 _06592_ (.A(net3578),
    .B(_00588_),
    .Y(_01138_));
 sg13g2_nor2_1 _06593_ (.A(_00019_),
    .B(net3354),
    .Y(_01139_));
 sg13g2_nand2b_2 _06594_ (.Y(_01140_),
    .B(\core.lsu.state[1] ),
    .A_N(\core.lsu.state[2] ));
 sg13g2_inv_1 _06595_ (.Y(_01141_),
    .A(_01140_));
 sg13g2_nor2_1 _06596_ (.A(\core.lsu.state[0] ),
    .B(_01140_),
    .Y(_01142_));
 sg13g2_or2_2 _06597_ (.X(_01143_),
    .B(_01140_),
    .A(\core.lsu.state[0] ));
 sg13g2_a21oi_1 _06598_ (.A1(_01136_),
    .A2(_01143_),
    .Y(_01144_),
    .B1(_01129_));
 sg13g2_nor3_1 _06599_ (.A(_01138_),
    .B(_01139_),
    .C(_01144_),
    .Y(_01145_));
 sg13g2_nand2_1 _06600_ (.Y(_01146_),
    .A(net3527),
    .B(net806));
 sg13g2_nor2_1 _06601_ (.A(_01143_),
    .B(_01146_),
    .Y(_01147_));
 sg13g2_nand2_1 _06602_ (.Y(_01148_),
    .A(\core.work.alu.sval2[31] ),
    .B(_00605_));
 sg13g2_xor2_1 _06603_ (.B(net3453),
    .A(\core.work.alu.sval2[23] ),
    .X(_01149_));
 sg13g2_and2_1 _06604_ (.A(\core.work.alu.sval2[22] ),
    .B(net3455),
    .X(_01150_));
 sg13g2_xor2_1 _06605_ (.B(net3455),
    .A(\core.work.alu.sval2[22] ),
    .X(_01151_));
 sg13g2_or2_1 _06606_ (.X(_01152_),
    .B(_01151_),
    .A(_01149_));
 sg13g2_xnor2_1 _06607_ (.Y(_01153_),
    .A(net3530),
    .B(net3465));
 sg13g2_xnor2_1 _06608_ (.Y(_01154_),
    .A(\core.work.alu.sval2[21] ),
    .B(net3458));
 sg13g2_nand2_1 _06609_ (.Y(_01155_),
    .A(_01153_),
    .B(_01154_));
 sg13g2_nor2_1 _06610_ (.A(_01152_),
    .B(_01155_),
    .Y(_01156_));
 sg13g2_xor2_1 _06611_ (.B(net3531),
    .A(\core.e2m_addr[19] ),
    .X(_01157_));
 sg13g2_nor2_1 _06612_ (.A(_00625_),
    .B(_00626_),
    .Y(_01158_));
 sg13g2_xor2_1 _06613_ (.B(\core.e2m_addr[18] ),
    .A(\core.work.alu.sval2[18] ),
    .X(_01159_));
 sg13g2_nor2_1 _06614_ (.A(_01157_),
    .B(_01159_),
    .Y(_01160_));
 sg13g2_inv_1 _06615_ (.Y(_01161_),
    .A(_01160_));
 sg13g2_nand2_1 _06616_ (.Y(_01162_),
    .A(net3535),
    .B(net3472));
 sg13g2_xor2_1 _06617_ (.B(net3472),
    .A(net3535),
    .X(_01163_));
 sg13g2_xor2_1 _06618_ (.B(net3470),
    .A(net3532),
    .X(_01164_));
 sg13g2_nor2_1 _06619_ (.A(_01163_),
    .B(_01164_),
    .Y(_01165_));
 sg13g2_nand2_1 _06620_ (.Y(_01166_),
    .A(net3487),
    .B(\core.work.alu.sval2[10] ));
 sg13g2_xor2_1 _06621_ (.B(\core.work.alu.sval2[10] ),
    .A(net3487),
    .X(_01167_));
 sg13g2_xnor2_1 _06622_ (.Y(_01168_),
    .A(net3486),
    .B(\core.work.alu.sval2[10] ));
 sg13g2_nor2_1 _06623_ (.A(\core.e2m_addr[11] ),
    .B(\core.work.alu.sval2[11] ),
    .Y(_01169_));
 sg13g2_nand2_1 _06624_ (.Y(_01170_),
    .A(\core.e2m_addr[11] ),
    .B(\core.work.alu.sval2[11] ));
 sg13g2_xnor2_1 _06625_ (.Y(_01171_),
    .A(\core.e2m_addr[11] ),
    .B(\core.work.alu.sval2[11] ));
 sg13g2_nor2_1 _06626_ (.A(\core.e2m_addr[9] ),
    .B(net3542),
    .Y(_01172_));
 sg13g2_nand2_1 _06627_ (.Y(_01173_),
    .A(net3488),
    .B(net3542));
 sg13g2_xnor2_1 _06628_ (.Y(_01174_),
    .A(net3488),
    .B(net3542));
 sg13g2_nand2_1 _06629_ (.Y(_01175_),
    .A(\core.e2m_addr[8] ),
    .B(\core.work.alu.sval2[8] ));
 sg13g2_xnor2_1 _06630_ (.Y(_01176_),
    .A(\core.e2m_addr[8] ),
    .B(\core.work.alu.sval2[8] ));
 sg13g2_and4_2 _06631_ (.A(_01168_),
    .B(_01171_),
    .C(_01174_),
    .D(_01176_),
    .X(_01177_));
 sg13g2_xnor2_1 _06632_ (.Y(_01178_),
    .A(\core.work.alu.sval2[15] ),
    .B(net3478));
 sg13g2_nand2b_1 _06633_ (.Y(_01179_),
    .B(net3481),
    .A_N(\core.work.alu.sval2[14] ));
 sg13g2_xor2_1 _06634_ (.B(net3481),
    .A(\core.work.alu.sval2[14] ),
    .X(_01180_));
 sg13g2_nor2b_1 _06635_ (.A(_01180_),
    .B_N(_01178_),
    .Y(_01181_));
 sg13g2_nor2_1 _06636_ (.A(\core.work.alu.sval2[13] ),
    .B(net3483),
    .Y(_01182_));
 sg13g2_nand2_1 _06637_ (.Y(_01183_),
    .A(\core.work.alu.sval2[13] ),
    .B(net3483));
 sg13g2_nor2b_1 _06638_ (.A(_01182_),
    .B_N(_01183_),
    .Y(_01184_));
 sg13g2_nand2b_1 _06639_ (.Y(_01185_),
    .B(_01183_),
    .A_N(_01182_));
 sg13g2_nand2_1 _06640_ (.Y(_01186_),
    .A(net3541),
    .B(net3485));
 sg13g2_xnor2_1 _06641_ (.Y(_01187_),
    .A(net3541),
    .B(net3485));
 sg13g2_nand4_1 _06642_ (.B(_01181_),
    .C(_01185_),
    .A(_01177_),
    .Y(_01188_),
    .D(_01187_));
 sg13g2_nor2_1 _06643_ (.A(_00593_),
    .B(\core.work.alu.sval2[7] ),
    .Y(_01189_));
 sg13g2_xnor2_1 _06644_ (.Y(_01190_),
    .A(\core.e2m_addr[7] ),
    .B(\core.work.alu.sval2[7] ));
 sg13g2_nor2_1 _06645_ (.A(\core.work.alu.sval2[6] ),
    .B(_00594_),
    .Y(_01191_));
 sg13g2_nor2_1 _06646_ (.A(net3543),
    .B(_00595_),
    .Y(_01192_));
 sg13g2_nor2_1 _06647_ (.A(net3543),
    .B(net3494),
    .Y(_01193_));
 sg13g2_xor2_1 _06648_ (.B(net3494),
    .A(\core.work.alu.sval2[5] ),
    .X(_01194_));
 sg13g2_xnor2_1 _06649_ (.Y(_01195_),
    .A(net3543),
    .B(net3493));
 sg13g2_nor2_1 _06650_ (.A(_00596_),
    .B(_00597_),
    .Y(_01196_));
 sg13g2_xor2_1 _06651_ (.B(\core.e2m_addr[4] ),
    .A(net3549),
    .X(_01197_));
 sg13g2_nand2_1 _06652_ (.Y(_01198_),
    .A(net3553),
    .B(\core.e2m_addr[3] ));
 sg13g2_xnor2_1 _06653_ (.Y(_01199_),
    .A(net3553),
    .B(\core.e2m_addr[3] ));
 sg13g2_nor2b_1 _06654_ (.A(net3557),
    .B_N(net3498),
    .Y(_01200_));
 sg13g2_nand2b_1 _06655_ (.Y(_01201_),
    .B(\core.e2m_addr[1] ),
    .A_N(net3560));
 sg13g2_nand2_1 _06656_ (.Y(_01202_),
    .A(net3560),
    .B(net3499));
 sg13g2_nor2_1 _06657_ (.A(net3560),
    .B(net3499),
    .Y(_01203_));
 sg13g2_xor2_1 _06658_ (.B(net3499),
    .A(net3560),
    .X(_01204_));
 sg13g2_nor2b_1 _06659_ (.A(net3500),
    .B_N(net3539),
    .Y(_01205_));
 sg13g2_o21ai_1 _06660_ (.B1(_01201_),
    .Y(_01206_),
    .A1(_01204_),
    .A2(_01205_));
 sg13g2_and2_1 _06661_ (.A(net3557),
    .B(net3498),
    .X(_01207_));
 sg13g2_or2_1 _06662_ (.X(_01208_),
    .B(net3497),
    .A(net3558));
 sg13g2_xnor2_1 _06663_ (.Y(_01209_),
    .A(net3557),
    .B(net3498));
 sg13g2_a21oi_1 _06664_ (.A1(_01206_),
    .A2(_01209_),
    .Y(_01210_),
    .B1(_01200_));
 sg13g2_and2_1 _06665_ (.A(_01199_),
    .B(_01209_),
    .X(_01211_));
 sg13g2_and2_1 _06666_ (.A(_01199_),
    .B(_01200_),
    .X(_01212_));
 sg13g2_a221oi_1 _06667_ (.B2(_01211_),
    .C1(_01212_),
    .B1(_01206_),
    .A1(_00592_),
    .Y(_01213_),
    .A2(net3496));
 sg13g2_nand2_1 _06668_ (.Y(_01214_),
    .A(_00596_),
    .B(net3495));
 sg13g2_o21ai_1 _06669_ (.B1(_01214_),
    .Y(_01215_),
    .A1(_01197_),
    .A2(_01213_));
 sg13g2_a21o_1 _06670_ (.A2(_01215_),
    .A1(_01195_),
    .B1(_01192_),
    .X(_01216_));
 sg13g2_xor2_1 _06671_ (.B(\core.e2m_addr[6] ),
    .A(\core.work.alu.sval2[6] ),
    .X(_01217_));
 sg13g2_xnor2_1 _06672_ (.Y(_01218_),
    .A(\core.work.alu.sval2[6] ),
    .B(\core.e2m_addr[6] ));
 sg13g2_and2_1 _06673_ (.A(_01216_),
    .B(_01218_),
    .X(_01219_));
 sg13g2_and2_1 _06674_ (.A(_01190_),
    .B(_01218_),
    .X(_01220_));
 sg13g2_o21ai_1 _06675_ (.B1(_01190_),
    .Y(_01221_),
    .A1(_01191_),
    .A2(_01219_));
 sg13g2_a221oi_1 _06676_ (.B2(_01220_),
    .C1(_01189_),
    .B1(_01216_),
    .A1(_01190_),
    .Y(_01222_),
    .A2(_01191_));
 sg13g2_nand2b_1 _06677_ (.Y(_01223_),
    .B(_01221_),
    .A_N(_01189_));
 sg13g2_nor2_1 _06678_ (.A(_01188_),
    .B(_01222_),
    .Y(_01224_));
 sg13g2_a21oi_1 _06679_ (.A1(\core.work.alu.sval2[15] ),
    .A2(_00599_),
    .Y(_01225_),
    .B1(_01179_));
 sg13g2_nand2b_1 _06680_ (.Y(_01226_),
    .B(net3483),
    .A_N(\core.work.alu.sval2[13] ));
 sg13g2_nand2b_1 _06681_ (.Y(_01227_),
    .B(net3485),
    .A_N(net3541));
 sg13g2_nand2b_1 _06682_ (.Y(_01228_),
    .B(\core.e2m_addr[11] ),
    .A_N(\core.work.alu.sval2[11] ));
 sg13g2_nor2b_1 _06683_ (.A(\core.work.alu.sval2[8] ),
    .B_N(\core.e2m_addr[8] ),
    .Y(_01229_));
 sg13g2_nand2_1 _06684_ (.Y(_01230_),
    .A(net3486),
    .B(_00602_));
 sg13g2_nor2b_1 _06685_ (.A(net3542),
    .B_N(net3488),
    .Y(_01231_));
 sg13g2_a221oi_1 _06686_ (.B2(_01229_),
    .C1(_01231_),
    .B1(_01174_),
    .A1(net3486),
    .Y(_01232_),
    .A2(_00602_));
 sg13g2_o21ai_1 _06687_ (.B1(_01171_),
    .Y(_01233_),
    .A1(net3486),
    .A2(_00602_));
 sg13g2_o21ai_1 _06688_ (.B1(_01228_),
    .Y(_01234_),
    .A1(_01232_),
    .A2(_01233_));
 sg13g2_nor2b_1 _06689_ (.A(_01234_),
    .B_N(_01227_),
    .Y(_01235_));
 sg13g2_a21o_1 _06690_ (.A2(_00601_),
    .A1(net3541),
    .B1(_01184_),
    .X(_01236_));
 sg13g2_o21ai_1 _06691_ (.B1(_01226_),
    .Y(_01237_),
    .A1(_01235_),
    .A2(_01236_));
 sg13g2_a221oi_1 _06692_ (.B2(_01237_),
    .C1(_01225_),
    .B1(_01181_),
    .A1(_00598_),
    .Y(_01238_),
    .A2(net3478));
 sg13g2_nor2b_1 _06693_ (.A(_01224_),
    .B_N(_01238_),
    .Y(_01239_));
 sg13g2_o21ai_1 _06694_ (.B1(_01238_),
    .Y(_01240_),
    .A1(_01188_),
    .A2(_01222_));
 sg13g2_nand2b_1 _06695_ (.Y(_01241_),
    .B(net3471),
    .A_N(net3535));
 sg13g2_a21oi_1 _06696_ (.A1(net3532),
    .A2(_00628_),
    .Y(_01242_),
    .B1(_01241_));
 sg13g2_a221oi_1 _06697_ (.B2(_01240_),
    .C1(_01242_),
    .B1(_01165_),
    .A1(_00627_),
    .Y(_01243_),
    .A2(net3469));
 sg13g2_nand2_1 _06698_ (.Y(_01244_),
    .A(_00625_),
    .B(\core.e2m_addr[18] ));
 sg13g2_a21oi_1 _06699_ (.A1(_00623_),
    .A2(net3531),
    .Y(_01245_),
    .B1(_01244_));
 sg13g2_a21oi_1 _06700_ (.A1(\core.e2m_addr[19] ),
    .A2(_00624_),
    .Y(_01246_),
    .B1(_01245_));
 sg13g2_o21ai_1 _06701_ (.B1(_01246_),
    .Y(_01247_),
    .A1(_01161_),
    .A2(_01243_));
 sg13g2_nor2_1 _06702_ (.A(net3530),
    .B(_00622_),
    .Y(_01248_));
 sg13g2_a21oi_1 _06703_ (.A1(_00619_),
    .A2(net3457),
    .Y(_01249_),
    .B1(_01248_));
 sg13g2_nor2_1 _06704_ (.A(_00619_),
    .B(net3457),
    .Y(_01250_));
 sg13g2_nor3_1 _06705_ (.A(_01152_),
    .B(_01249_),
    .C(_01250_),
    .Y(_01251_));
 sg13g2_nand2_1 _06706_ (.Y(_01252_),
    .A(_00618_),
    .B(net3455));
 sg13g2_o21ai_1 _06707_ (.B1(_00617_),
    .Y(_01253_),
    .A1(net3534),
    .A2(_01252_));
 sg13g2_nand2_1 _06708_ (.Y(_01254_),
    .A(net3534),
    .B(_01252_));
 sg13g2_a221oi_1 _06709_ (.B2(_01254_),
    .C1(_01251_),
    .B1(_01253_),
    .A1(_01156_),
    .Y(_01255_),
    .A2(_01247_));
 sg13g2_nor2_1 _06710_ (.A(net3537),
    .B(_00611_),
    .Y(_01256_));
 sg13g2_nand2_1 _06711_ (.Y(_01257_),
    .A(net3537),
    .B(_00611_));
 sg13g2_nand2b_2 _06712_ (.Y(_01258_),
    .B(_01257_),
    .A_N(_01256_));
 sg13g2_nor2_1 _06713_ (.A(\core.work.alu.sval2[26] ),
    .B(_00613_),
    .Y(_01259_));
 sg13g2_xor2_1 _06714_ (.B(\core.e2m_addr[26] ),
    .A(\core.work.alu.sval2[26] ),
    .X(_01260_));
 sg13g2_nor2_1 _06715_ (.A(_01258_),
    .B(_01260_),
    .Y(_01261_));
 sg13g2_nor2_1 _06716_ (.A(net3533),
    .B(_00615_),
    .Y(_01262_));
 sg13g2_xor2_1 _06717_ (.B(net3451),
    .A(net3533),
    .X(_01263_));
 sg13g2_nand2b_1 _06718_ (.Y(_01264_),
    .B(net3536),
    .A_N(net3450));
 sg13g2_nand2b_2 _06719_ (.Y(_01265_),
    .B(net3450),
    .A_N(net3536));
 sg13g2_nand2_2 _06720_ (.Y(_01266_),
    .A(_01264_),
    .B(_01265_));
 sg13g2_nor4_2 _06721_ (.A(_01258_),
    .B(_01260_),
    .C(_01263_),
    .Y(_01267_),
    .D(_01266_));
 sg13g2_inv_1 _06722_ (.Y(_01268_),
    .A(_01267_));
 sg13g2_nand2_1 _06723_ (.Y(_01269_),
    .A(_01262_),
    .B(_01264_));
 sg13g2_nand2_1 _06724_ (.Y(_01270_),
    .A(_01265_),
    .B(_01269_));
 sg13g2_a221oi_1 _06725_ (.B2(_01270_),
    .C1(_01256_),
    .B1(_01261_),
    .A1(_01257_),
    .Y(_01271_),
    .A2(_01259_));
 sg13g2_o21ai_1 _06726_ (.B1(_01271_),
    .Y(_01272_),
    .A1(_01255_),
    .A2(_01268_));
 sg13g2_xor2_1 _06727_ (.B(\core.e2m_addr[31] ),
    .A(\core.work.alu.sval2[31] ),
    .X(_01273_));
 sg13g2_nand2_1 _06728_ (.Y(_01274_),
    .A(_00606_),
    .B(\core.e2m_addr[30] ));
 sg13g2_xnor2_1 _06729_ (.Y(_01275_),
    .A(\core.work.alu.sval2[30] ),
    .B(\core.e2m_addr[30] ));
 sg13g2_xor2_1 _06730_ (.B(net3444),
    .A(\core.work.alu.sval2[30] ),
    .X(_01276_));
 sg13g2_nor2_1 _06731_ (.A(_01273_),
    .B(_01276_),
    .Y(_01277_));
 sg13g2_nand2_1 _06732_ (.Y(_01278_),
    .A(_00608_),
    .B(net3446));
 sg13g2_nor2_1 _06733_ (.A(_00608_),
    .B(net3446),
    .Y(_01279_));
 sg13g2_xnor2_1 _06734_ (.Y(_01280_),
    .A(net3540),
    .B(net3445));
 sg13g2_xor2_1 _06735_ (.B(net3445),
    .A(net3540),
    .X(_01281_));
 sg13g2_nand2_1 _06736_ (.Y(_01282_),
    .A(\core.work.alu.sval2[28] ),
    .B(net3447));
 sg13g2_xor2_1 _06737_ (.B(\core.e2m_addr[28] ),
    .A(\core.work.alu.sval2[28] ),
    .X(_01283_));
 sg13g2_inv_1 _06738_ (.Y(_01284_),
    .A(_01283_));
 sg13g2_nor4_2 _06739_ (.A(_01273_),
    .B(_01276_),
    .C(_01281_),
    .Y(_01285_),
    .D(_01283_));
 sg13g2_nand2_1 _06740_ (.Y(_01286_),
    .A(_00610_),
    .B(net3447));
 sg13g2_o21ai_1 _06741_ (.B1(_01278_),
    .Y(_01287_),
    .A1(_01279_),
    .A2(_01286_));
 sg13g2_nand2b_1 _06742_ (.Y(_01288_),
    .B(_01148_),
    .A_N(_01274_));
 sg13g2_o21ai_1 _06743_ (.B1(_01288_),
    .Y(_01289_),
    .A1(\core.work.alu.sval2[31] ),
    .A2(_00605_));
 sg13g2_a221oi_1 _06744_ (.B2(_01277_),
    .C1(_01289_),
    .B1(_01287_),
    .A1(_01272_),
    .Y(_01290_),
    .A2(_01285_));
 sg13g2_nand2_1 _06745_ (.Y(_01291_),
    .A(_01272_),
    .B(_01284_));
 sg13g2_nand3_1 _06746_ (.B(_01280_),
    .C(_01284_),
    .A(_01272_),
    .Y(_01292_));
 sg13g2_nor2b_1 _06747_ (.A(_01287_),
    .B_N(_01292_),
    .Y(_01293_));
 sg13g2_o21ai_1 _06748_ (.B1(_01274_),
    .Y(_01294_),
    .A1(_01276_),
    .A2(_01293_));
 sg13g2_o21ai_1 _06749_ (.B1(_01148_),
    .Y(_01295_),
    .A1(_01273_),
    .A2(_01290_));
 sg13g2_and2_2 _06750_ (.A(\core.work.alu.is_sign ),
    .B(\core.work.alu.is_wr ),
    .X(_01296_));
 sg13g2_nand2_2 _06751_ (.Y(_01297_),
    .A(\core.work.alu.is_sign ),
    .B(\core.work.alu.is_wr ));
 sg13g2_nor2b_1 _06752_ (.A(net3441),
    .B_N(\core.work.alu.ls_size_b ),
    .Y(_01298_));
 sg13g2_nand2_1 _06753_ (.Y(_01299_),
    .A(_01296_),
    .B(_01298_));
 sg13g2_nand3_1 _06754_ (.B(\core.work.alu.ls_size_b ),
    .C(_01296_),
    .A(net3441),
    .Y(_01300_));
 sg13g2_nand2b_1 _06755_ (.Y(_01301_),
    .B(net3441),
    .A_N(\core.work.alu.ls_size_b ));
 sg13g2_nor2_1 _06756_ (.A(_01297_),
    .B(_01301_),
    .Y(_01302_));
 sg13g2_xor2_1 _06757_ (.B(net3500),
    .A(net3538),
    .X(_01303_));
 sg13g2_nor4_2 _06758_ (.A(_01194_),
    .B(_01197_),
    .C(_01204_),
    .Y(_01304_),
    .D(_01303_));
 sg13g2_nand4_1 _06759_ (.B(_01267_),
    .C(_01285_),
    .A(_01156_),
    .Y(_01305_),
    .D(_01304_));
 sg13g2_nand4_1 _06760_ (.B(_01165_),
    .C(_01211_),
    .A(_01160_),
    .Y(_01306_),
    .D(_01220_));
 sg13g2_nor3_2 _06761_ (.A(_01188_),
    .B(_01305_),
    .C(_01306_),
    .Y(_01307_));
 sg13g2_nor2b_2 _06762_ (.A(\core.work.alu.is_sign ),
    .B_N(\core.work.alu.is_wr ),
    .Y(_01308_));
 sg13g2_nand2_2 _06763_ (.Y(_01309_),
    .A(_00629_),
    .B(net3440));
 sg13g2_nand2_1 _06764_ (.Y(_01310_),
    .A(_01298_),
    .B(_01308_));
 sg13g2_nor2_1 _06765_ (.A(_01307_),
    .B(_01310_),
    .Y(_01311_));
 sg13g2_nor2_2 _06766_ (.A(net3441),
    .B(\core.work.alu.ls_size_b ),
    .Y(_01312_));
 sg13g2_and2_1 _06767_ (.A(_01308_),
    .B(_01312_),
    .X(_01313_));
 sg13g2_nor2_2 _06768_ (.A(\core.work.alu.is_sign ),
    .B(net3440),
    .Y(_01314_));
 sg13g2_a221oi_1 _06769_ (.B2(_01312_),
    .C1(_01311_),
    .B1(_01314_),
    .A1(_01307_),
    .Y(_01315_),
    .A2(_01313_));
 sg13g2_o21ai_1 _06770_ (.B1(_01315_),
    .Y(_01316_),
    .A1(_01290_),
    .A2(_01300_));
 sg13g2_a21oi_2 _06771_ (.B1(_01316_),
    .Y(_01317_),
    .A2(_01302_),
    .A1(_01290_));
 sg13g2_nand2_1 _06772_ (.Y(_01318_),
    .A(_01296_),
    .B(_01312_));
 sg13g2_mux2_1 _06773_ (.A0(_01318_),
    .A1(_01299_),
    .S(_01295_),
    .X(_01319_));
 sg13g2_nand2_2 _06774_ (.Y(_01320_),
    .A(\core.work.op[4] ),
    .B(_00630_));
 sg13g2_a21oi_2 _06775_ (.B1(_01320_),
    .Y(_01321_),
    .A2(_01319_),
    .A1(_01317_));
 sg13g2_a21o_2 _06776_ (.A2(_01319_),
    .A1(_01317_),
    .B1(_01320_),
    .X(_01322_));
 sg13g2_nor2_2 _06777_ (.A(net3501),
    .B(net3502),
    .Y(_01323_));
 sg13g2_and2_2 _06778_ (.A(net3513),
    .B(net3512),
    .X(_01324_));
 sg13g2_nand2_2 _06779_ (.Y(_01325_),
    .A(net3513),
    .B(net3512));
 sg13g2_a21oi_2 _06780_ (.B1(\core.fetch.inst_size[2] ),
    .Y(_01326_),
    .A2(net3338),
    .A1(net3528));
 sg13g2_nor3_2 _06781_ (.A(net3501),
    .B(net3502),
    .C(_01326_),
    .Y(_01327_));
 sg13g2_or3_1 _06782_ (.A(net3501),
    .B(net3502),
    .C(_01326_),
    .X(_01328_));
 sg13g2_nor2b_1 _06783_ (.A(\core.fetch.state[0] ),
    .B_N(net3578),
    .Y(_01329_));
 sg13g2_and2_1 _06784_ (.A(net3044),
    .B(_01329_),
    .X(_01330_));
 sg13g2_nand2_1 _06785_ (.Y(_01331_),
    .A(_00019_),
    .B(_01330_));
 sg13g2_nor2_1 _06786_ (.A(net3578),
    .B(\core.fetch.state[0] ),
    .Y(_01332_));
 sg13g2_nand4_1 _06787_ (.B(net3528),
    .C(_01143_),
    .A(net3527),
    .Y(_01333_),
    .D(_01332_));
 sg13g2_o21ai_1 _06788_ (.B1(_01333_),
    .Y(_01334_),
    .A1(\core.fetch.state[0] ),
    .A2(net3044));
 sg13g2_nand2_1 _06789_ (.Y(_01335_),
    .A(net3566),
    .B(_01330_));
 sg13g2_o21ai_1 _06790_ (.B1(_01335_),
    .Y(_01336_),
    .A1(_00062_),
    .A2(_01331_));
 sg13g2_nor2_1 _06791_ (.A(_01334_),
    .B(_01336_),
    .Y(_01337_));
 sg13g2_o21ai_1 _06792_ (.B1(_01145_),
    .Y(_01338_),
    .A1(net2737),
    .A2(_01337_));
 sg13g2_nor3_1 _06793_ (.A(net3578),
    .B(_01321_),
    .C(_01338_),
    .Y(_01339_));
 sg13g2_nand2_1 _06794_ (.Y(_01340_),
    .A(_01147_),
    .B(_01339_));
 sg13g2_nand2_1 _06795_ (.Y(_00183_),
    .A(_01145_),
    .B(_01340_));
 sg13g2_a21o_1 _06796_ (.A2(_01338_),
    .A1(net3578),
    .B1(_01339_),
    .X(_00184_));
 sg13g2_nor2b_1 _06797_ (.A(\core.fetch.data_size[2] ),
    .B_N(net3585),
    .Y(_01341_));
 sg13g2_nand4_1 _06798_ (.B(net3355),
    .C(_00985_),
    .A(net3566),
    .Y(_01342_),
    .D(_01341_));
 sg13g2_nor3_1 _06799_ (.A(net3577),
    .B(net3576),
    .C(_01342_),
    .Y(_01343_));
 sg13g2_mux2_1 _06800_ (.A0(net492),
    .A1(net3570),
    .S(net2849),
    .X(_00185_));
 sg13g2_mux2_1 _06801_ (.A0(net610),
    .A1(net587),
    .S(net2849),
    .X(_00186_));
 sg13g2_nor2_1 _06802_ (.A(net569),
    .B(net2849),
    .Y(_01344_));
 sg13g2_a21oi_1 _06803_ (.A1(_00681_),
    .A2(net2849),
    .Y(_00187_),
    .B1(_01344_));
 sg13g2_nor2_1 _06804_ (.A(net465),
    .B(net2850),
    .Y(_01345_));
 sg13g2_a21oi_1 _06805_ (.A1(_00684_),
    .A2(net2850),
    .Y(_00188_),
    .B1(_01345_));
 sg13g2_nor2_1 _06806_ (.A(net593),
    .B(net2849),
    .Y(_01346_));
 sg13g2_a21oi_1 _06807_ (.A1(_00686_),
    .A2(net2849),
    .Y(_00189_),
    .B1(_01346_));
 sg13g2_nor2_1 _06808_ (.A(net401),
    .B(net2850),
    .Y(_01347_));
 sg13g2_a21oi_1 _06809_ (.A1(_00689_),
    .A2(net2850),
    .Y(_00190_),
    .B1(_01347_));
 sg13g2_nor2_1 _06810_ (.A(net442),
    .B(net2849),
    .Y(_01348_));
 sg13g2_a21oi_1 _06811_ (.A1(_00691_),
    .A2(net2850),
    .Y(_00191_),
    .B1(_01348_));
 sg13g2_nor2_1 _06812_ (.A(net455),
    .B(net2849),
    .Y(_01349_));
 sg13g2_a21oi_1 _06813_ (.A1(_00693_),
    .A2(net2850),
    .Y(_00192_),
    .B1(_01349_));
 sg13g2_nor3_2 _06814_ (.A(_00649_),
    .B(net3576),
    .C(_01342_),
    .Y(_01350_));
 sg13g2_mux2_1 _06815_ (.A0(net490),
    .A1(net3570),
    .S(_01350_),
    .X(_00193_));
 sg13g2_mux2_1 _06816_ (.A0(net479),
    .A1(net3569),
    .S(_01350_),
    .X(_00194_));
 sg13g2_mux2_1 _06817_ (.A0(net504),
    .A1(\core.fetch.cmd_data[2] ),
    .S(_01350_),
    .X(_00195_));
 sg13g2_mux2_1 _06818_ (.A0(net640),
    .A1(net571),
    .S(_01350_),
    .X(_00196_));
 sg13g2_mux2_1 _06819_ (.A0(net642),
    .A1(\core.fetch.cmd_data[4] ),
    .S(_01350_),
    .X(_00197_));
 sg13g2_mux2_1 _06820_ (.A0(net397),
    .A1(\core.fetch.cmd_data[5] ),
    .S(_01350_),
    .X(_00198_));
 sg13g2_mux2_1 _06821_ (.A0(net390),
    .A1(\core.fetch.cmd_data[6] ),
    .S(_01350_),
    .X(_00199_));
 sg13g2_mux2_1 _06822_ (.A0(net522),
    .A1(\core.fetch.cmd_data[7] ),
    .S(_01350_),
    .X(_00200_));
 sg13g2_nor3_1 _06823_ (.A(net3577),
    .B(_00650_),
    .C(_01342_),
    .Y(_01351_));
 sg13g2_nor2_1 _06824_ (.A(\core.fetch.data[16] ),
    .B(net2848),
    .Y(_01352_));
 sg13g2_a21oi_1 _06825_ (.A1(net477),
    .A2(net2848),
    .Y(_00201_),
    .B1(_01352_));
 sg13g2_nor2_1 _06826_ (.A(\core.fetch.data[17] ),
    .B(net2848),
    .Y(_01353_));
 sg13g2_a21oi_1 _06827_ (.A1(net515),
    .A2(net2848),
    .Y(_00202_),
    .B1(_01353_));
 sg13g2_nor2_1 _06828_ (.A(\core.fetch.data[18] ),
    .B(net2847),
    .Y(_01354_));
 sg13g2_a21oi_1 _06829_ (.A1(net601),
    .A2(net2847),
    .Y(_00203_),
    .B1(_01354_));
 sg13g2_nor2_1 _06830_ (.A(\core.fetch.data[19] ),
    .B(net2847),
    .Y(_01355_));
 sg13g2_a21oi_1 _06831_ (.A1(net452),
    .A2(net2848),
    .Y(_00204_),
    .B1(_01355_));
 sg13g2_nor2_1 _06832_ (.A(\core.fetch.data[20] ),
    .B(net2847),
    .Y(_01356_));
 sg13g2_a21oi_1 _06833_ (.A1(net500),
    .A2(net2847),
    .Y(_00205_),
    .B1(_01356_));
 sg13g2_nor2_1 _06834_ (.A(\core.fetch.data[21] ),
    .B(net2848),
    .Y(_01357_));
 sg13g2_a21oi_1 _06835_ (.A1(net421),
    .A2(_01351_),
    .Y(_00206_),
    .B1(_01357_));
 sg13g2_nor2_1 _06836_ (.A(\core.fetch.data[22] ),
    .B(net2847),
    .Y(_01358_));
 sg13g2_a21oi_1 _06837_ (.A1(net429),
    .A2(net2847),
    .Y(_00207_),
    .B1(_01358_));
 sg13g2_nor2_1 _06838_ (.A(\core.fetch.data[23] ),
    .B(net2847),
    .Y(_01359_));
 sg13g2_a21oi_1 _06839_ (.A1(net411),
    .A2(net2848),
    .Y(_00208_),
    .B1(_01359_));
 sg13g2_nand2_1 _06840_ (.Y(_01360_),
    .A(net3577),
    .B(net3576));
 sg13g2_nor2_1 _06841_ (.A(_01342_),
    .B(_01360_),
    .Y(_01361_));
 sg13g2_mux2_1 _06842_ (.A0(net464),
    .A1(net3570),
    .S(net2845),
    .X(_00209_));
 sg13g2_mux2_1 _06843_ (.A0(net370),
    .A1(net3569),
    .S(net2845),
    .X(_00210_));
 sg13g2_nor2_1 _06844_ (.A(net404),
    .B(net2845),
    .Y(_01362_));
 sg13g2_a21oi_1 _06845_ (.A1(_00681_),
    .A2(net2845),
    .Y(_00211_),
    .B1(_01362_));
 sg13g2_nor2_1 _06846_ (.A(net383),
    .B(net2846),
    .Y(_01363_));
 sg13g2_a21oi_1 _06847_ (.A1(_00684_),
    .A2(net2845),
    .Y(_00212_),
    .B1(_01363_));
 sg13g2_nor2_1 _06848_ (.A(net367),
    .B(net2846),
    .Y(_01364_));
 sg13g2_a21oi_1 _06849_ (.A1(_00686_),
    .A2(net2846),
    .Y(_00213_),
    .B1(_01364_));
 sg13g2_nor2_1 _06850_ (.A(net388),
    .B(net2845),
    .Y(_01365_));
 sg13g2_a21oi_1 _06851_ (.A1(_00689_),
    .A2(net2845),
    .Y(_00214_),
    .B1(_01365_));
 sg13g2_nor2_1 _06852_ (.A(net423),
    .B(net2846),
    .Y(_01366_));
 sg13g2_a21oi_1 _06853_ (.A1(_00691_),
    .A2(net2846),
    .Y(_00215_),
    .B1(_01366_));
 sg13g2_nor2_1 _06854_ (.A(net416),
    .B(net2846),
    .Y(_01367_));
 sg13g2_a21oi_1 _06855_ (.A1(_00693_),
    .A2(net2845),
    .Y(_00216_),
    .B1(_01367_));
 sg13g2_nor2_1 _06856_ (.A(net2737),
    .B(_01327_),
    .Y(_01368_));
 sg13g2_nor2b_1 _06857_ (.A(_01147_),
    .B_N(_01332_),
    .Y(_01369_));
 sg13g2_nand2_1 _06858_ (.Y(_01370_),
    .A(_00986_),
    .B(_01139_));
 sg13g2_or2_2 _06859_ (.X(_01371_),
    .B(_01332_),
    .A(net3355));
 sg13g2_inv_1 _06860_ (.Y(_01372_),
    .A(_01371_));
 sg13g2_nand3_1 _06861_ (.B(_01370_),
    .C(_01371_),
    .A(_01129_),
    .Y(_01373_));
 sg13g2_a21oi_1 _06862_ (.A1(net2736),
    .A2(net3044),
    .Y(_01374_),
    .B1(net3578));
 sg13g2_a221oi_1 _06863_ (.B2(_00588_),
    .C1(_01373_),
    .B1(_01374_),
    .A1(_01368_),
    .Y(_01375_),
    .A2(_01369_));
 sg13g2_nand4_1 _06864_ (.B(\core.fetch.state[0] ),
    .C(net3566),
    .A(net3578),
    .Y(_01376_),
    .D(_01370_));
 sg13g2_and2_1 _06865_ (.A(_00649_),
    .B(_01376_),
    .X(_01377_));
 sg13g2_a21oi_1 _06866_ (.A1(net3577),
    .A2(_01375_),
    .Y(_00217_),
    .B1(_01377_));
 sg13g2_nand2_1 _06867_ (.Y(_01378_),
    .A(net3355),
    .B(_01360_));
 sg13g2_and2_1 _06868_ (.A(_01375_),
    .B(_01378_),
    .X(_01379_));
 sg13g2_a21oi_1 _06869_ (.A1(net3577),
    .A2(_01375_),
    .Y(_01380_),
    .B1(net3576));
 sg13g2_nor2_1 _06870_ (.A(_01379_),
    .B(_01380_),
    .Y(_00218_));
 sg13g2_nor2_1 _06871_ (.A(_01360_),
    .B(_01376_),
    .Y(_01381_));
 sg13g2_nor2_1 _06872_ (.A(net796),
    .B(_01381_),
    .Y(_01382_));
 sg13g2_a21oi_1 _06873_ (.A1(net796),
    .A2(_01379_),
    .Y(_00219_),
    .B1(_01382_));
 sg13g2_nand2_1 _06874_ (.Y(_01383_),
    .A(net3575),
    .B(net356));
 sg13g2_nand2b_1 _06875_ (.Y(_01384_),
    .B(net3572),
    .A_N(net3574));
 sg13g2_o21ai_1 _06876_ (.B1(_01384_),
    .Y(_00220_),
    .A1(_00984_),
    .A2(net357));
 sg13g2_nand2_1 _06877_ (.Y(_01385_),
    .A(net3584),
    .B(net3575));
 sg13g2_nand2_1 _06878_ (.Y(_01386_),
    .A(net418),
    .B(net3333));
 sg13g2_nand2b_1 _06879_ (.Y(_01387_),
    .B(net3572),
    .A_N(\core.fetch.spi_reader.cache_bit ));
 sg13g2_o21ai_1 _06880_ (.B1(_01387_),
    .Y(_01388_),
    .A1(net3573),
    .A2(\core.fetch.cmd_data[0] ));
 sg13g2_a21oi_1 _06881_ (.A1(_00979_),
    .A2(_01388_),
    .Y(_01389_),
    .B1(_00749_));
 sg13g2_nor3_2 _06882_ (.A(_00632_),
    .B(net3567),
    .C(\core.fetch.spi_reader.state[2] ),
    .Y(_01390_));
 sg13g2_nand3b_1 _06883_ (.B(_00633_),
    .C(\core.fetch.spi_reader.state[0] ),
    .Y(_01391_),
    .A_N(net3567));
 sg13g2_nor2_1 _06884_ (.A(_00747_),
    .B(_01390_),
    .Y(_01392_));
 sg13g2_nor2b_1 _06885_ (.A(net3572),
    .B_N(\core.fetch.spi_reader.counter[0] ),
    .Y(_01393_));
 sg13g2_nor4_1 _06886_ (.A(\core.fetch.spi_reader.counter[1] ),
    .B(\core.fetch.spi_reader.counter[5] ),
    .C(_00982_),
    .D(_01393_),
    .Y(_01394_));
 sg13g2_inv_1 _06887_ (.Y(_01395_),
    .A(_01394_));
 sg13g2_nand2b_1 _06888_ (.Y(_01396_),
    .B(_00992_),
    .A_N(_00061_));
 sg13g2_nand2b_1 _06889_ (.Y(_01397_),
    .B(_01390_),
    .A_N(_00083_));
 sg13g2_a22oi_1 _06890_ (.Y(_01398_),
    .B1(_01396_),
    .B2(_01397_),
    .A2(_01388_),
    .A1(net3362));
 sg13g2_a21oi_1 _06891_ (.A1(net3200),
    .A2(_01398_),
    .Y(_01399_),
    .B1(_01392_));
 sg13g2_nand2_1 _06892_ (.Y(_01400_),
    .A(net3565),
    .B(net3200));
 sg13g2_o21ai_1 _06893_ (.B1(_01400_),
    .Y(_01401_),
    .A1(_00992_),
    .A2(_01390_));
 sg13g2_o21ai_1 _06894_ (.B1(_01399_),
    .Y(_01402_),
    .A1(_01388_),
    .A2(_01401_));
 sg13g2_a21oi_1 _06895_ (.A1(_01388_),
    .A2(_01392_),
    .Y(_01403_),
    .B1(net3333));
 sg13g2_o21ai_1 _06896_ (.B1(_01403_),
    .Y(_01404_),
    .A1(_01389_),
    .A2(_01402_));
 sg13g2_nand2_1 _06897_ (.Y(_00221_),
    .A(_01386_),
    .B(_01404_));
 sg13g2_mux2_1 _06898_ (.A0(_00097_),
    .A1(net870),
    .S(net3571),
    .X(_01405_));
 sg13g2_a21o_1 _06899_ (.A2(_01405_),
    .A1(_00979_),
    .B1(_00749_),
    .X(_01406_));
 sg13g2_a22oi_1 _06900_ (.Y(_01407_),
    .B1(_01390_),
    .B2(\core.fetch.spi_reader.addr[9] ),
    .A2(_00992_),
    .A1(\core.fetch.spi_reader.addr[1] ));
 sg13g2_nor2_1 _06901_ (.A(_01400_),
    .B(_01407_),
    .Y(_01408_));
 sg13g2_nor2_1 _06902_ (.A(_01401_),
    .B(_01405_),
    .Y(_01409_));
 sg13g2_nor3_1 _06903_ (.A(net3039),
    .B(_01408_),
    .C(_01409_),
    .Y(_01410_));
 sg13g2_a221oi_1 _06904_ (.B2(_01410_),
    .C1(net3333),
    .B1(_01406_),
    .A1(net3039),
    .Y(_01411_),
    .A2(_01405_));
 sg13g2_a21o_1 _06905_ (.A2(net3333),
    .A1(net3569),
    .B1(_01411_),
    .X(_00222_));
 sg13g2_a21oi_2 _06906_ (.B1(net3039),
    .Y(_01412_),
    .A2(_00979_),
    .A1(_00748_));
 sg13g2_mux2_1 _06907_ (.A0(net871),
    .A1(_00097_),
    .S(net3571),
    .X(_01413_));
 sg13g2_or2_1 _06908_ (.X(_01414_),
    .B(_01413_),
    .A(_01412_));
 sg13g2_nor2_1 _06909_ (.A(_00063_),
    .B(_00993_),
    .Y(_01415_));
 sg13g2_nor2_1 _06910_ (.A(_00081_),
    .B(_01391_),
    .Y(_01416_));
 sg13g2_o21ai_1 _06911_ (.B1(net3200),
    .Y(_01417_),
    .A1(_01415_),
    .A2(_01416_));
 sg13g2_o21ai_1 _06912_ (.B1(_01417_),
    .Y(_01418_),
    .A1(_01401_),
    .A2(_01413_));
 sg13g2_a21oi_1 _06913_ (.A1(net3362),
    .A2(_01413_),
    .Y(_01419_),
    .B1(net3039));
 sg13g2_a21oi_1 _06914_ (.A1(_01418_),
    .A2(_01419_),
    .Y(_01420_),
    .B1(net3333));
 sg13g2_a22oi_1 _06915_ (.Y(_00223_),
    .B1(_01414_),
    .B2(_01420_),
    .A2(net3333),
    .A1(_00681_));
 sg13g2_nor2b_1 _06916_ (.A(net3571),
    .B_N(_00099_),
    .Y(_01421_));
 sg13g2_a221oi_1 _06917_ (.B2(_01412_),
    .C1(_01421_),
    .B1(_01401_),
    .A1(net3571),
    .Y(_01422_),
    .A2(net871));
 sg13g2_a22oi_1 _06918_ (.Y(_01423_),
    .B1(_01390_),
    .B2(net3568),
    .A2(_00992_),
    .A1(net494));
 sg13g2_nor2_1 _06919_ (.A(_01400_),
    .B(_01423_),
    .Y(_01424_));
 sg13g2_nor3_1 _06920_ (.A(net3334),
    .B(net872),
    .C(_01424_),
    .Y(_01425_));
 sg13g2_a21oi_1 _06921_ (.A1(_00684_),
    .A2(net3334),
    .Y(_00224_),
    .B1(_01425_));
 sg13g2_mux2_1 _06922_ (.A0(_00100_),
    .A1(net877),
    .S(net3571),
    .X(_01426_));
 sg13g2_or2_1 _06923_ (.X(_01427_),
    .B(net878),
    .A(_01412_));
 sg13g2_nor2_1 _06924_ (.A(_00070_),
    .B(_00993_),
    .Y(_01428_));
 sg13g2_nor2_1 _06925_ (.A(_00077_),
    .B(_01391_),
    .Y(_01429_));
 sg13g2_o21ai_1 _06926_ (.B1(net3200),
    .Y(_01430_),
    .A1(_01428_),
    .A2(_01429_));
 sg13g2_o21ai_1 _06927_ (.B1(_01430_),
    .Y(_01431_),
    .A1(_01401_),
    .A2(_01426_));
 sg13g2_a21oi_1 _06928_ (.A1(net3362),
    .A2(_01426_),
    .Y(_01432_),
    .B1(net3039));
 sg13g2_a21oi_1 _06929_ (.A1(_01431_),
    .A2(_01432_),
    .Y(_01433_),
    .B1(net3334));
 sg13g2_a22oi_1 _06930_ (.Y(_00225_),
    .B1(_01427_),
    .B2(_01433_),
    .A2(net3334),
    .A1(_00686_));
 sg13g2_mux2_1 _06931_ (.A0(net888),
    .A1(net890),
    .S(net3571),
    .X(_01434_));
 sg13g2_or2_1 _06932_ (.X(_01435_),
    .B(_01434_),
    .A(_01412_));
 sg13g2_nand2_1 _06933_ (.Y(_01436_),
    .A(\core.fetch.spi_reader.addr[13] ),
    .B(_01390_));
 sg13g2_o21ai_1 _06934_ (.B1(_01436_),
    .Y(_01437_),
    .A1(_00068_),
    .A2(_00993_));
 sg13g2_nand2_1 _06935_ (.Y(_01438_),
    .A(net3200),
    .B(_01437_));
 sg13g2_o21ai_1 _06936_ (.B1(_01438_),
    .Y(_01439_),
    .A1(_01401_),
    .A2(_01434_));
 sg13g2_a21oi_1 _06937_ (.A1(net3362),
    .A2(_01434_),
    .Y(_01440_),
    .B1(net3039));
 sg13g2_a21oi_1 _06938_ (.A1(_01439_),
    .A2(_01440_),
    .Y(_01441_),
    .B1(net3334));
 sg13g2_a22oi_1 _06939_ (.Y(_00226_),
    .B1(_01435_),
    .B2(_01441_),
    .A2(net3334),
    .A1(_00689_));
 sg13g2_mux2_1 _06940_ (.A0(_00102_),
    .A1(net888),
    .S(net3571),
    .X(_01442_));
 sg13g2_or2_1 _06941_ (.X(_01443_),
    .B(net889),
    .A(_01412_));
 sg13g2_nor2_1 _06942_ (.A(_00074_),
    .B(_01391_),
    .Y(_01444_));
 sg13g2_nor2_1 _06943_ (.A(_00067_),
    .B(_00993_),
    .Y(_01445_));
 sg13g2_o21ai_1 _06944_ (.B1(net3200),
    .Y(_01446_),
    .A1(_01444_),
    .A2(_01445_));
 sg13g2_o21ai_1 _06945_ (.B1(_01446_),
    .Y(_01447_),
    .A1(_01401_),
    .A2(_01442_));
 sg13g2_a21oi_1 _06946_ (.A1(net3362),
    .A2(_01442_),
    .Y(_01448_),
    .B1(net3039));
 sg13g2_a21oi_1 _06947_ (.A1(_01447_),
    .A2(_01448_),
    .Y(_01449_),
    .B1(net3334));
 sg13g2_a22oi_1 _06948_ (.Y(_00227_),
    .B1(_01443_),
    .B2(_01449_),
    .A2(net3334),
    .A1(_00691_));
 sg13g2_mux2_1 _06949_ (.A0(net893),
    .A1(_00102_),
    .S(net3571),
    .X(_01450_));
 sg13g2_or2_1 _06950_ (.X(_01451_),
    .B(net894),
    .A(_01412_));
 sg13g2_nand2_1 _06951_ (.Y(_01452_),
    .A(\core.fetch.spi_reader.addr[7] ),
    .B(_00992_));
 sg13g2_o21ai_1 _06952_ (.B1(_01452_),
    .Y(_01453_),
    .A1(_00071_),
    .A2(_01391_));
 sg13g2_nand2_1 _06953_ (.Y(_01454_),
    .A(net3200),
    .B(_01453_));
 sg13g2_o21ai_1 _06954_ (.B1(_01454_),
    .Y(_01455_),
    .A1(_01401_),
    .A2(_01450_));
 sg13g2_a21oi_1 _06955_ (.A1(net3362),
    .A2(_01450_),
    .Y(_01456_),
    .B1(net3039));
 sg13g2_a21oi_1 _06956_ (.A1(_01455_),
    .A2(_01456_),
    .Y(_01457_),
    .B1(net3333));
 sg13g2_a22oi_1 _06957_ (.Y(_00228_),
    .B1(_01451_),
    .B2(_01457_),
    .A2(net3333),
    .A1(_00693_));
 sg13g2_nand2b_1 _06958_ (.Y(_01458_),
    .B(net3584),
    .A_N(uio_out[0]));
 sg13g2_nor3_1 _06959_ (.A(net3572),
    .B(_00984_),
    .C(_01458_),
    .Y(_01459_));
 sg13g2_mux2_1 _06960_ (.A0(net387),
    .A1(net9),
    .S(_01459_),
    .X(_00229_));
 sg13g2_nor2_1 _06961_ (.A(net3565),
    .B(_00749_),
    .Y(_01460_));
 sg13g2_o21ai_1 _06962_ (.B1(_00989_),
    .Y(_01461_),
    .A1(\core.fetch.spi_reader.state[2] ),
    .A2(_00749_));
 sg13g2_nand3_1 _06963_ (.B(_00964_),
    .C(_00967_),
    .A(\core.fetch.spi_reader.dirty ),
    .Y(_01462_));
 sg13g2_o21ai_1 _06964_ (.B1(_01461_),
    .Y(_01463_),
    .A1(_00749_),
    .A2(_01462_));
 sg13g2_nor4_1 _06965_ (.A(_00987_),
    .B(_01458_),
    .C(_01460_),
    .D(_01463_),
    .Y(_01464_));
 sg13g2_nor2_1 _06966_ (.A(net496),
    .B(net2752),
    .Y(_01465_));
 sg13g2_nand2_1 _06967_ (.Y(_01466_),
    .A(_00832_),
    .B(net3206));
 sg13g2_o21ai_1 _06968_ (.B1(_01466_),
    .Y(_01467_),
    .A1(_00061_),
    .A2(net3206));
 sg13g2_a21oi_1 _06969_ (.A1(net2752),
    .A2(_01467_),
    .Y(_00230_),
    .B1(_01465_));
 sg13g2_nand2_2 _06970_ (.Y(_01468_),
    .A(\core.fetch.spi_reader.addr[0] ),
    .B(\core.fetch.spi_reader.addr[1] ));
 sg13g2_or2_1 _06971_ (.X(_01469_),
    .B(\core.fetch.spi_reader.addr[1] ),
    .A(\core.fetch.spi_reader.addr[0] ));
 sg13g2_nand3_1 _06972_ (.B(_01468_),
    .C(_01469_),
    .A(net3210),
    .Y(_01470_));
 sg13g2_o21ai_1 _06973_ (.B1(_01470_),
    .Y(_01471_),
    .A1(_00828_),
    .A2(net3210));
 sg13g2_mux2_1 _06974_ (.A0(net739),
    .A1(_01471_),
    .S(net2752),
    .X(_00231_));
 sg13g2_o21ai_1 _06975_ (.B1(net3210),
    .Y(_01472_),
    .A1(\core.fetch.spi_reader.addr[2] ),
    .A2(_01468_));
 sg13g2_a21oi_1 _06976_ (.A1(net628),
    .A2(_01468_),
    .Y(_01473_),
    .B1(_01472_));
 sg13g2_a21oi_1 _06977_ (.A1(_00841_),
    .A2(net3207),
    .Y(_01474_),
    .B1(_01473_));
 sg13g2_mux2_1 _06978_ (.A0(net628),
    .A1(_01474_),
    .S(net2752),
    .X(_00232_));
 sg13g2_nor2_1 _06979_ (.A(net494),
    .B(net2752),
    .Y(_01475_));
 sg13g2_nor2_1 _06980_ (.A(_00063_),
    .B(_01468_),
    .Y(_01476_));
 sg13g2_xnor2_1 _06981_ (.Y(_01477_),
    .A(net494),
    .B(_01476_));
 sg13g2_nand2_1 _06982_ (.Y(_01478_),
    .A(net3210),
    .B(_01477_));
 sg13g2_o21ai_1 _06983_ (.B1(_01478_),
    .Y(_01479_),
    .A1(_00823_),
    .A2(net3210));
 sg13g2_a21oi_1 _06984_ (.A1(net2752),
    .A2(_01479_),
    .Y(_00233_),
    .B1(_01475_));
 sg13g2_nor2_1 _06985_ (.A(net588),
    .B(net2754),
    .Y(_01480_));
 sg13g2_nor3_2 _06986_ (.A(_00658_),
    .B(_00659_),
    .C(_01468_),
    .Y(_01481_));
 sg13g2_xor2_1 _06987_ (.B(_01481_),
    .A(net588),
    .X(_01482_));
 sg13g2_nor2_1 _06988_ (.A(_00852_),
    .B(net3208),
    .Y(_01483_));
 sg13g2_a21oi_1 _06989_ (.A1(net3208),
    .A2(_01482_),
    .Y(_01484_),
    .B1(_01483_));
 sg13g2_a21oi_1 _06990_ (.A1(net2754),
    .A2(_01484_),
    .Y(_00234_),
    .B1(_01480_));
 sg13g2_a21o_1 _06991_ (.A2(_01481_),
    .A1(_00662_),
    .B1(\core.fetch.spi_reader.addr[5] ),
    .X(_01485_));
 sg13g2_nand3_1 _06992_ (.B(_00662_),
    .C(_01481_),
    .A(\core.fetch.spi_reader.addr[5] ),
    .Y(_01486_));
 sg13g2_nand3_1 _06993_ (.B(_01485_),
    .C(_01486_),
    .A(net3208),
    .Y(_01487_));
 sg13g2_o21ai_1 _06994_ (.B1(_01487_),
    .Y(_01488_),
    .A1(_00817_),
    .A2(net3208));
 sg13g2_mux2_1 _06995_ (.A0(net645),
    .A1(_01488_),
    .S(net2754),
    .X(_00235_));
 sg13g2_nor2_1 _06996_ (.A(net674),
    .B(net2754),
    .Y(_01489_));
 sg13g2_and3_1 _06997_ (.X(_01490_),
    .A(\core.fetch.spi_reader.addr[5] ),
    .B(\core.fetch.spi_reader.addr[4] ),
    .C(_01481_));
 sg13g2_xor2_1 _06998_ (.B(_01490_),
    .A(\core.fetch.spi_reader.addr[6] ),
    .X(_01491_));
 sg13g2_nand2_1 _06999_ (.Y(_01492_),
    .A(_00865_),
    .B(net3207));
 sg13g2_o21ai_1 _07000_ (.B1(_01492_),
    .Y(_01493_),
    .A1(net3207),
    .A2(_01491_));
 sg13g2_a21oi_1 _07001_ (.A1(net2754),
    .A2(_01493_),
    .Y(_00236_),
    .B1(_01489_));
 sg13g2_nor2_1 _07002_ (.A(net695),
    .B(net2754),
    .Y(_01494_));
 sg13g2_nor2b_1 _07003_ (.A(_00067_),
    .B_N(_01490_),
    .Y(_01495_));
 sg13g2_xnor2_1 _07004_ (.Y(_01496_),
    .A(\core.fetch.spi_reader.addr[7] ),
    .B(_01495_));
 sg13g2_nand2_1 _07005_ (.Y(_01497_),
    .A(net3208),
    .B(_01496_));
 sg13g2_o21ai_1 _07006_ (.B1(_01497_),
    .Y(_01498_),
    .A1(_00811_),
    .A2(net3208));
 sg13g2_a21oi_1 _07007_ (.A1(net2754),
    .A2(_01498_),
    .Y(_00237_),
    .B1(_01494_));
 sg13g2_nor2_1 _07008_ (.A(net676),
    .B(net2755),
    .Y(_01499_));
 sg13g2_and3_2 _07009_ (.X(_01500_),
    .A(\core.fetch.spi_reader.addr[7] ),
    .B(\core.fetch.spi_reader.addr[6] ),
    .C(_01490_));
 sg13g2_xor2_1 _07010_ (.B(_01500_),
    .A(\core.fetch.spi_reader.addr[8] ),
    .X(_01501_));
 sg13g2_nand2_1 _07011_ (.Y(_01502_),
    .A(_00803_),
    .B(net3207));
 sg13g2_o21ai_1 _07012_ (.B1(_01502_),
    .Y(_01503_),
    .A1(net3207),
    .A2(_01501_));
 sg13g2_a21oi_1 _07013_ (.A1(net2754),
    .A2(_01503_),
    .Y(_00238_),
    .B1(_01499_));
 sg13g2_nor2_1 _07014_ (.A(net801),
    .B(net2755),
    .Y(_01504_));
 sg13g2_nand2b_1 _07015_ (.Y(_01505_),
    .B(_01500_),
    .A_N(_00083_));
 sg13g2_a21oi_1 _07016_ (.A1(\core.fetch.spi_reader.addr[9] ),
    .A2(_01505_),
    .Y(_01506_),
    .B1(net3207));
 sg13g2_o21ai_1 _07017_ (.B1(_01506_),
    .Y(_01507_),
    .A1(\core.fetch.spi_reader.addr[9] ),
    .A2(_01505_));
 sg13g2_o21ai_1 _07018_ (.B1(_01507_),
    .Y(_01508_),
    .A1(_00796_),
    .A2(net3209));
 sg13g2_a21oi_1 _07019_ (.A1(net2755),
    .A2(_01508_),
    .Y(_00239_),
    .B1(_01504_));
 sg13g2_nor2_1 _07020_ (.A(net655),
    .B(net2755),
    .Y(_01509_));
 sg13g2_and4_1 _07021_ (.A(\core.fetch.spi_reader.addr[10] ),
    .B(\core.fetch.spi_reader.addr[9] ),
    .C(\core.fetch.spi_reader.addr[8] ),
    .D(_01500_),
    .X(_01510_));
 sg13g2_and2_1 _07022_ (.A(\core.fetch.spi_reader.addr[9] ),
    .B(_01500_),
    .X(_01511_));
 sg13g2_nand2_1 _07023_ (.Y(_01512_),
    .A(\core.fetch.spi_reader.addr[8] ),
    .B(_01511_));
 sg13g2_xnor2_1 _07024_ (.Y(_01513_),
    .A(\core.fetch.spi_reader.addr[10] ),
    .B(_01512_));
 sg13g2_nor2_1 _07025_ (.A(_00886_),
    .B(net3209),
    .Y(_01514_));
 sg13g2_a21oi_1 _07026_ (.A1(net3209),
    .A2(_01513_),
    .Y(_01515_),
    .B1(_01514_));
 sg13g2_a21oi_1 _07027_ (.A1(net2755),
    .A2(_01515_),
    .Y(_00240_),
    .B1(_01509_));
 sg13g2_nor2_1 _07028_ (.A(net3568),
    .B(net2755),
    .Y(_01516_));
 sg13g2_nor2_1 _07029_ (.A(_00880_),
    .B(net3209),
    .Y(_01517_));
 sg13g2_nor2_1 _07030_ (.A(_00081_),
    .B(_01512_),
    .Y(_01518_));
 sg13g2_xor2_1 _07031_ (.B(_01518_),
    .A(net3568),
    .X(_01519_));
 sg13g2_a21oi_1 _07032_ (.A1(net3208),
    .A2(_01519_),
    .Y(_01520_),
    .B1(_01517_));
 sg13g2_a21oi_1 _07033_ (.A1(net2755),
    .A2(_01520_),
    .Y(_00241_),
    .B1(_01516_));
 sg13g2_nor2_1 _07034_ (.A(net596),
    .B(net2752),
    .Y(_01521_));
 sg13g2_nand2_1 _07035_ (.Y(_01522_),
    .A(_00911_),
    .B(net3207));
 sg13g2_nand4_1 _07036_ (.B(\core.fetch.spi_reader.addr[10] ),
    .C(\core.fetch.spi_reader.addr[8] ),
    .A(net3568),
    .Y(_01523_),
    .D(_01511_));
 sg13g2_xnor2_1 _07037_ (.Y(_01524_),
    .A(net596),
    .B(_01523_));
 sg13g2_o21ai_1 _07038_ (.B1(_01522_),
    .Y(_01525_),
    .A1(net3207),
    .A2(_01524_));
 sg13g2_a21oi_1 _07039_ (.A1(net2752),
    .A2(_01525_),
    .Y(_00242_),
    .B1(_01521_));
 sg13g2_nor2_1 _07040_ (.A(net705),
    .B(net2753),
    .Y(_01526_));
 sg13g2_nor2_1 _07041_ (.A(_00077_),
    .B(_01523_),
    .Y(_01527_));
 sg13g2_xnor2_1 _07042_ (.Y(_01528_),
    .A(\core.fetch.spi_reader.addr[13] ),
    .B(_01527_));
 sg13g2_nor2_1 _07043_ (.A(net3206),
    .B(_01528_),
    .Y(_01529_));
 sg13g2_a21oi_1 _07044_ (.A1(_00904_),
    .A2(net3206),
    .Y(_01530_),
    .B1(_01529_));
 sg13g2_a21oi_1 _07045_ (.A1(net2753),
    .A2(_01530_),
    .Y(_00243_),
    .B1(_01526_));
 sg13g2_nor2_1 _07046_ (.A(net469),
    .B(net2753),
    .Y(_01531_));
 sg13g2_and4_1 _07047_ (.A(\core.fetch.spi_reader.addr[13] ),
    .B(\core.fetch.spi_reader.addr[12] ),
    .C(\core.fetch.spi_reader.addr[11] ),
    .D(_01510_),
    .X(_01532_));
 sg13g2_xor2_1 _07048_ (.B(_01532_),
    .A(net469),
    .X(_01533_));
 sg13g2_nor2_1 _07049_ (.A(_00895_),
    .B(net3210),
    .Y(_01534_));
 sg13g2_a21oi_1 _07050_ (.A1(net3210),
    .A2(_01533_),
    .Y(_01535_),
    .B1(_01534_));
 sg13g2_a21oi_1 _07051_ (.A1(net2753),
    .A2(_01535_),
    .Y(_00244_),
    .B1(_01531_));
 sg13g2_nor2_1 _07052_ (.A(net547),
    .B(net2753),
    .Y(_01536_));
 sg13g2_nor2b_1 _07053_ (.A(_00074_),
    .B_N(_01532_),
    .Y(_01537_));
 sg13g2_xnor2_1 _07054_ (.Y(_01538_),
    .A(net547),
    .B(_01537_));
 sg13g2_nor2_1 _07055_ (.A(net3206),
    .B(_01538_),
    .Y(_01539_));
 sg13g2_a21oi_1 _07056_ (.A1(_00788_),
    .A2(net3206),
    .Y(_01540_),
    .B1(_01539_));
 sg13g2_a21oi_1 _07057_ (.A1(net2753),
    .A2(_01540_),
    .Y(_00245_),
    .B1(_01536_));
 sg13g2_nor2_1 _07058_ (.A(_00019_),
    .B(_00994_),
    .Y(_01541_));
 sg13g2_a21oi_1 _07059_ (.A1(_00993_),
    .A2(_01391_),
    .Y(_01542_),
    .B1(_00019_));
 sg13g2_or2_1 _07060_ (.X(_01543_),
    .B(_01542_),
    .A(_01541_));
 sg13g2_a21oi_1 _07061_ (.A1(_01395_),
    .A2(_01543_),
    .Y(_01544_),
    .B1(_01460_));
 sg13g2_and3_1 _07062_ (.X(_01545_),
    .A(_00988_),
    .B(_00997_),
    .C(_01544_));
 sg13g2_inv_1 _07063_ (.Y(_01546_),
    .A(_01545_));
 sg13g2_and3_1 _07064_ (.X(_01547_),
    .A(net3206),
    .B(_00993_),
    .C(_00994_));
 sg13g2_inv_1 _07065_ (.Y(_01548_),
    .A(_01547_));
 sg13g2_o21ai_1 _07066_ (.B1(_01545_),
    .Y(_01549_),
    .A1(_00019_),
    .A2(_00993_));
 sg13g2_a21oi_1 _07067_ (.A1(_01462_),
    .A2(_01547_),
    .Y(_01550_),
    .B1(_01549_));
 sg13g2_a21oi_1 _07068_ (.A1(_00632_),
    .A2(_01546_),
    .Y(_00246_),
    .B1(_01550_));
 sg13g2_mux2_1 _07069_ (.A0(net470),
    .A1(_01542_),
    .S(_01545_),
    .X(_00247_));
 sg13g2_a221oi_1 _07070_ (.B2(_00978_),
    .C1(_01546_),
    .B1(_01547_),
    .A1(_01391_),
    .Y(_01551_),
    .A2(_01541_));
 sg13g2_a21oi_1 _07071_ (.A1(_00633_),
    .A2(_01546_),
    .Y(_00248_),
    .B1(_01551_));
 sg13g2_nand2_1 _07072_ (.Y(_01552_),
    .A(_01327_),
    .B(_01329_));
 sg13g2_a21oi_1 _07073_ (.A1(_01333_),
    .A2(_01552_),
    .Y(_01553_),
    .B1(net2737));
 sg13g2_nor3_1 _07074_ (.A(_01138_),
    .B(_01374_),
    .C(_01553_),
    .Y(_01554_));
 sg13g2_o21ai_1 _07075_ (.B1(_01329_),
    .Y(_01555_),
    .A1(net3566),
    .A2(_00656_));
 sg13g2_a21oi_1 _07076_ (.A1(net3565),
    .A2(_00985_),
    .Y(_01556_),
    .B1(_01555_));
 sg13g2_and2_1 _07077_ (.A(net2736),
    .B(_01556_),
    .X(_01557_));
 sg13g2_nand3_1 _07078_ (.B(net3565),
    .C(_00986_),
    .A(\core.fetch.state[0] ),
    .Y(_01558_));
 sg13g2_nand3b_1 _07079_ (.B(_01558_),
    .C(net3578),
    .Y(_01559_),
    .A_N(_01137_));
 sg13g2_o21ai_1 _07080_ (.B1(_01554_),
    .Y(_01560_),
    .A1(_01557_),
    .A2(_01559_));
 sg13g2_o21ai_1 _07081_ (.B1(_01560_),
    .Y(_00249_),
    .A1(_00631_),
    .A2(_01554_));
 sg13g2_nor2b_1 _07082_ (.A(_01460_),
    .B_N(net3575),
    .Y(_01561_));
 sg13g2_nand3_1 _07083_ (.B(_00989_),
    .C(_01561_),
    .A(_00988_),
    .Y(_01562_));
 sg13g2_o21ai_1 _07084_ (.B1(net436),
    .Y(_01563_),
    .A1(_00995_),
    .A2(_01562_));
 sg13g2_o21ai_1 _07085_ (.B1(_01563_),
    .Y(_00250_),
    .A1(_01548_),
    .A2(_01562_));
 sg13g2_nor2_2 _07086_ (.A(_01138_),
    .B(_01368_),
    .Y(_01564_));
 sg13g2_a21oi_1 _07087_ (.A1(net3503),
    .A2(\core.f2e_addr[2] ),
    .Y(_01565_),
    .B1(_01324_));
 sg13g2_o21ai_1 _07088_ (.B1(_01565_),
    .Y(_01566_),
    .A1(net3503),
    .A2(\core.f2e_addr[2] ));
 sg13g2_nand2_1 _07089_ (.Y(_01567_),
    .A(net636),
    .B(_01324_));
 sg13g2_a21oi_1 _07090_ (.A1(_01566_),
    .A2(_01567_),
    .Y(_01568_),
    .B1(net2739));
 sg13g2_a21oi_1 _07091_ (.A1(net629),
    .A2(net2739),
    .Y(_01569_),
    .B1(_01568_));
 sg13g2_nor2_1 _07092_ (.A(\core.f2e_addr[2] ),
    .B(net2733),
    .Y(_01570_));
 sg13g2_a21oi_1 _07093_ (.A1(net2733),
    .A2(_01569_),
    .Y(_00251_),
    .B1(_01570_));
 sg13g2_nor2_2 _07094_ (.A(net3503),
    .B(net3349),
    .Y(_01571_));
 sg13g2_nor2b_1 _07095_ (.A(_01571_),
    .B_N(\core.f2e_addr[2] ),
    .Y(_01572_));
 sg13g2_nand2_1 _07096_ (.Y(_01573_),
    .A(\core.f2e_addr[2] ),
    .B(\core.f2e_addr[3] ));
 sg13g2_nor2_1 _07097_ (.A(_01571_),
    .B(_01573_),
    .Y(_01574_));
 sg13g2_nor2_1 _07098_ (.A(\core.f2e_addr[3] ),
    .B(_01572_),
    .Y(_01575_));
 sg13g2_nor3_1 _07099_ (.A(net2740),
    .B(_01574_),
    .C(_01575_),
    .Y(_01576_));
 sg13g2_a21oi_1 _07100_ (.A1(net457),
    .A2(net2740),
    .Y(_01577_),
    .B1(_01576_));
 sg13g2_nor2_1 _07101_ (.A(net622),
    .B(net2734),
    .Y(_01578_));
 sg13g2_a21oi_1 _07102_ (.A1(net2733),
    .A2(_01577_),
    .Y(_00252_),
    .B1(_01578_));
 sg13g2_nor2_1 _07103_ (.A(net427),
    .B(net2734),
    .Y(_01579_));
 sg13g2_and2_2 _07104_ (.A(net3564),
    .B(_01574_),
    .X(_01580_));
 sg13g2_nor2_1 _07105_ (.A(net3564),
    .B(_01574_),
    .Y(_01581_));
 sg13g2_nor3_1 _07106_ (.A(net2740),
    .B(_01580_),
    .C(_01581_),
    .Y(_01582_));
 sg13g2_a21oi_1 _07107_ (.A1(\core.e2m_data[4] ),
    .A2(net2740),
    .Y(_01583_),
    .B1(_01582_));
 sg13g2_a21oi_1 _07108_ (.A1(net2734),
    .A2(_01583_),
    .Y(_00253_),
    .B1(_01579_));
 sg13g2_xnor2_1 _07109_ (.Y(_01584_),
    .A(\core.f2e_addr[5] ),
    .B(_01580_));
 sg13g2_nor2_1 _07110_ (.A(net2740),
    .B(_01584_),
    .Y(_01585_));
 sg13g2_a21oi_1 _07111_ (.A1(net546),
    .A2(net2739),
    .Y(_01586_),
    .B1(_01585_));
 sg13g2_nor2_1 _07112_ (.A(net698),
    .B(net2734),
    .Y(_01587_));
 sg13g2_a21oi_1 _07113_ (.A1(net2734),
    .A2(_01586_),
    .Y(_00254_),
    .B1(_01587_));
 sg13g2_a21oi_1 _07114_ (.A1(\core.f2e_addr[5] ),
    .A2(_01580_),
    .Y(_01588_),
    .B1(\core.f2e_addr[6] ));
 sg13g2_a21oi_1 _07115_ (.A1(_00777_),
    .A2(_01580_),
    .Y(_01589_),
    .B1(_01588_));
 sg13g2_mux2_1 _07116_ (.A0(net517),
    .A1(_01589_),
    .S(_01322_),
    .X(_01590_));
 sg13g2_nand2_1 _07117_ (.Y(_01591_),
    .A(net2733),
    .B(_01590_));
 sg13g2_o21ai_1 _07118_ (.B1(_01591_),
    .Y(_00255_),
    .A1(_00660_),
    .A2(net2733));
 sg13g2_nand3_1 _07119_ (.B(_00777_),
    .C(_01580_),
    .A(net3563),
    .Y(_01592_));
 sg13g2_a21o_1 _07120_ (.A2(_01580_),
    .A1(_00777_),
    .B1(net3563),
    .X(_01593_));
 sg13g2_a21oi_1 _07121_ (.A1(_01592_),
    .A2(_01593_),
    .Y(_01594_),
    .B1(net2739));
 sg13g2_a21oi_1 _07122_ (.A1(_00713_),
    .A2(net2739),
    .Y(_01595_),
    .B1(_01594_));
 sg13g2_mux2_1 _07123_ (.A0(net3563),
    .A1(_01595_),
    .S(net2733),
    .X(_00256_));
 sg13g2_nor2_1 _07124_ (.A(_00776_),
    .B(_01573_),
    .Y(_01596_));
 sg13g2_and4_1 _07125_ (.A(net3564),
    .B(net3563),
    .C(\core.f2e_addr[8] ),
    .D(_01596_),
    .X(_01597_));
 sg13g2_nand4_1 _07126_ (.B(net3563),
    .C(\core.f2e_addr[8] ),
    .A(net3564),
    .Y(_01598_),
    .D(_01596_));
 sg13g2_nor2_2 _07127_ (.A(_01571_),
    .B(_01598_),
    .Y(_01599_));
 sg13g2_a21oi_1 _07128_ (.A1(_00664_),
    .A2(_01592_),
    .Y(_01600_),
    .B1(_01599_));
 sg13g2_mux2_1 _07129_ (.A0(net560),
    .A1(_01600_),
    .S(net2736),
    .X(_01601_));
 sg13g2_nand2_1 _07130_ (.Y(_01602_),
    .A(net2733),
    .B(_01601_));
 sg13g2_o21ai_1 _07131_ (.B1(_01602_),
    .Y(_00257_),
    .A1(_00664_),
    .A2(net2733));
 sg13g2_xnor2_1 _07132_ (.Y(_01603_),
    .A(\core.f2e_addr[9] ),
    .B(_01599_));
 sg13g2_nor2_1 _07133_ (.A(net2739),
    .B(_01603_),
    .Y(_01604_));
 sg13g2_a21oi_1 _07134_ (.A1(net635),
    .A2(net2739),
    .Y(_01605_),
    .B1(_01604_));
 sg13g2_nor2_1 _07135_ (.A(net670),
    .B(net2732),
    .Y(_01606_));
 sg13g2_a21oi_1 _07136_ (.A1(net2732),
    .A2(_01605_),
    .Y(_00258_),
    .B1(_01606_));
 sg13g2_a21oi_1 _07137_ (.A1(\core.f2e_addr[9] ),
    .A2(_01599_),
    .Y(_01607_),
    .B1(\core.f2e_addr[10] ));
 sg13g2_nand2_1 _07138_ (.Y(_01608_),
    .A(_00781_),
    .B(_01599_));
 sg13g2_nor2b_1 _07139_ (.A(_01607_),
    .B_N(_01608_),
    .Y(_01609_));
 sg13g2_mux2_1 _07140_ (.A0(net542),
    .A1(_01609_),
    .S(net2736),
    .X(_01610_));
 sg13g2_nand2_1 _07141_ (.Y(_01611_),
    .A(net2732),
    .B(_01610_));
 sg13g2_o21ai_1 _07142_ (.B1(_01611_),
    .Y(_00259_),
    .A1(_00663_),
    .A2(net2732));
 sg13g2_nor2_1 _07143_ (.A(net685),
    .B(net2732),
    .Y(_01612_));
 sg13g2_xor2_1 _07144_ (.B(_01608_),
    .A(\core.f2e_addr[11] ),
    .X(_01613_));
 sg13g2_nor2_1 _07145_ (.A(net2739),
    .B(_01613_),
    .Y(_01614_));
 sg13g2_a21oi_1 _07146_ (.A1(net619),
    .A2(net2741),
    .Y(_01615_),
    .B1(_01614_));
 sg13g2_a21oi_1 _07147_ (.A1(net2732),
    .A2(_01615_),
    .Y(_00260_),
    .B1(_01612_));
 sg13g2_nor2_1 _07148_ (.A(net612),
    .B(net2731),
    .Y(_01616_));
 sg13g2_nand2_1 _07149_ (.Y(_01617_),
    .A(\core.f2e_addr[11] ),
    .B(net3349));
 sg13g2_o21ai_1 _07150_ (.B1(_01617_),
    .Y(_01618_),
    .A1(_00078_),
    .A2(net3349));
 sg13g2_nand3_1 _07151_ (.B(_01599_),
    .C(_01618_),
    .A(_00781_),
    .Y(_01619_));
 sg13g2_xor2_1 _07152_ (.B(_01619_),
    .A(\core.f2e_addr[12] ),
    .X(_01620_));
 sg13g2_nor2_1 _07153_ (.A(net2738),
    .B(_01620_),
    .Y(_01621_));
 sg13g2_a21oi_1 _07154_ (.A1(net521),
    .A2(net2738),
    .Y(_01622_),
    .B1(_01621_));
 sg13g2_a21oi_1 _07155_ (.A1(net2731),
    .A2(_01622_),
    .Y(_00261_),
    .B1(_01616_));
 sg13g2_nor2_1 _07156_ (.A(\core.f2e_addr[13] ),
    .B(net2731),
    .Y(_01623_));
 sg13g2_nand2_1 _07157_ (.Y(_01624_),
    .A(_00784_),
    .B(_01599_));
 sg13g2_xor2_1 _07158_ (.B(_01624_),
    .A(\core.f2e_addr[13] ),
    .X(_01625_));
 sg13g2_nor2_1 _07159_ (.A(net2738),
    .B(_01625_),
    .Y(_01626_));
 sg13g2_a21oi_1 _07160_ (.A1(net597),
    .A2(net2738),
    .Y(_01627_),
    .B1(_01626_));
 sg13g2_a21oi_1 _07161_ (.A1(net2731),
    .A2(_01627_),
    .Y(_00262_),
    .B1(_01623_));
 sg13g2_nor2_1 _07162_ (.A(net669),
    .B(net2731),
    .Y(_01628_));
 sg13g2_nand3_1 _07163_ (.B(net3349),
    .C(_01597_),
    .A(_00784_),
    .Y(_01629_));
 sg13g2_nor2_1 _07164_ (.A(_00075_),
    .B(net3349),
    .Y(_01630_));
 sg13g2_nand3_1 _07165_ (.B(_00784_),
    .C(net3349),
    .A(\core.f2e_addr[13] ),
    .Y(_01631_));
 sg13g2_nand4_1 _07166_ (.B(_00784_),
    .C(_01597_),
    .A(net3503),
    .Y(_01632_),
    .D(_01630_));
 sg13g2_o21ai_1 _07167_ (.B1(_01632_),
    .Y(_01633_),
    .A1(_01598_),
    .A2(_01631_));
 sg13g2_xnor2_1 _07168_ (.Y(_01634_),
    .A(\core.f2e_addr[14] ),
    .B(_01633_));
 sg13g2_nor2_1 _07169_ (.A(net2738),
    .B(_01634_),
    .Y(_01635_));
 sg13g2_a21oi_1 _07170_ (.A1(net644),
    .A2(net2738),
    .Y(_01636_),
    .B1(_01635_));
 sg13g2_a21oi_1 _07171_ (.A1(net2731),
    .A2(_01636_),
    .Y(_00263_),
    .B1(_01628_));
 sg13g2_nor2_1 _07172_ (.A(\core.f2e_addr[15] ),
    .B(net2731),
    .Y(_01637_));
 sg13g2_nand4_1 _07173_ (.B(_00784_),
    .C(_01325_),
    .A(net3503),
    .Y(_01638_),
    .D(_01597_));
 sg13g2_a21oi_1 _07174_ (.A1(_01629_),
    .A2(_01638_),
    .Y(_01639_),
    .B1(_00783_));
 sg13g2_xnor2_1 _07175_ (.Y(_01640_),
    .A(\core.f2e_addr[15] ),
    .B(_01639_));
 sg13g2_nor2_1 _07176_ (.A(net2738),
    .B(_01640_),
    .Y(_01641_));
 sg13g2_a21oi_1 _07177_ (.A1(net617),
    .A2(net2738),
    .Y(_01642_),
    .B1(_01641_));
 sg13g2_a21oi_1 _07178_ (.A1(net2731),
    .A2(_01642_),
    .Y(_00264_),
    .B1(_01637_));
 sg13g2_nand2_1 _07179_ (.Y(_01643_),
    .A(_01323_),
    .B(_01326_));
 sg13g2_and3_1 _07180_ (.X(_01644_),
    .A(net3595),
    .B(_01127_),
    .C(_01643_));
 sg13g2_nor2b_2 _07181_ (.A(net3501),
    .B_N(net3502),
    .Y(_01645_));
 sg13g2_nand2b_2 _07182_ (.Y(_01646_),
    .B(net859),
    .A_N(\core.work.state[1] ));
 sg13g2_a21oi_2 _07183_ (.B1(\core.gpio.stray_wr_i ),
    .Y(_01647_),
    .A2(_01125_),
    .A1(_00021_));
 sg13g2_nand2_2 _07184_ (.Y(_01648_),
    .A(\core.lsu.dreg[1] ),
    .B(_01647_));
 sg13g2_xnor2_1 _07185_ (.Y(_01649_),
    .A(net3472),
    .B(_01648_));
 sg13g2_nand2_2 _07186_ (.Y(_01650_),
    .A(\core.lsu.dreg[0] ),
    .B(_01647_));
 sg13g2_nand2_2 _07187_ (.Y(_01651_),
    .A(\core.lsu.dreg[2] ),
    .B(_01647_));
 sg13g2_xnor2_1 _07188_ (.Y(_01652_),
    .A(net3470),
    .B(_01651_));
 sg13g2_nand2_2 _07189_ (.Y(_01653_),
    .A(\core.lsu.dreg[3] ),
    .B(_01647_));
 sg13g2_xnor2_1 _07190_ (.Y(_01654_),
    .A(net3468),
    .B(_01653_));
 sg13g2_nor2_1 _07191_ (.A(net3468),
    .B(net3469),
    .Y(_01655_));
 sg13g2_nor3_2 _07192_ (.A(net3468),
    .B(net3470),
    .C(net3472),
    .Y(_01656_));
 sg13g2_nand2b_1 _07193_ (.Y(_01657_),
    .B(_01655_),
    .A_N(net3471));
 sg13g2_o21ai_1 _07194_ (.B1(_01650_),
    .Y(_01658_),
    .A1(net3475),
    .A2(net3323));
 sg13g2_o21ai_1 _07195_ (.B1(_01658_),
    .Y(_01659_),
    .A1(net3475),
    .A2(_01650_));
 sg13g2_or4_1 _07196_ (.A(_01649_),
    .B(_01652_),
    .C(_01654_),
    .D(_01659_),
    .X(_01660_));
 sg13g2_nand3b_1 _07197_ (.B(net3499),
    .C(net3500),
    .Y(_01661_),
    .A_N(net3496));
 sg13g2_nor2_1 _07198_ (.A(net3497),
    .B(_01661_),
    .Y(_01662_));
 sg13g2_nor3_2 _07199_ (.A(net3497),
    .B(\core.e2m_addr[6] ),
    .C(_01661_),
    .Y(_01663_));
 sg13g2_nor2b_1 _07200_ (.A(net3495),
    .B_N(net3493),
    .Y(_01664_));
 sg13g2_and2_2 _07201_ (.A(_01663_),
    .B(_01664_),
    .X(_01665_));
 sg13g2_nor2b_2 _07202_ (.A(_00020_),
    .B_N(_01664_),
    .Y(_01666_));
 sg13g2_and2_1 _07203_ (.A(_01662_),
    .B(_01666_),
    .X(_01667_));
 sg13g2_nand2_2 _07204_ (.Y(_01668_),
    .A(_01662_),
    .B(_01666_));
 sg13g2_and2_1 _07205_ (.A(net3495),
    .B(_01663_),
    .X(_01669_));
 sg13g2_nand2_2 _07206_ (.Y(_01670_),
    .A(net3495),
    .B(_01663_));
 sg13g2_nor2_2 _07207_ (.A(_00595_),
    .B(_01670_),
    .Y(_01671_));
 sg13g2_nand2_2 _07208_ (.Y(_01672_),
    .A(net3493),
    .B(_01669_));
 sg13g2_nand2_2 _07209_ (.Y(_01673_),
    .A(net3035),
    .B(_01672_));
 sg13g2_xnor2_1 _07210_ (.Y(_01674_),
    .A(net3456),
    .B(_01651_));
 sg13g2_nor3_1 _07211_ (.A(net3454),
    .B(net3456),
    .C(net3459),
    .Y(_01675_));
 sg13g2_o21ai_1 _07212_ (.B1(_01650_),
    .Y(_01676_),
    .A1(net3462),
    .A2(net3314));
 sg13g2_o21ai_1 _07213_ (.B1(_01676_),
    .Y(_01677_),
    .A1(net3462),
    .A2(_01650_));
 sg13g2_xnor2_1 _07214_ (.Y(_01678_),
    .A(net3454),
    .B(_01653_));
 sg13g2_xnor2_1 _07215_ (.Y(_01679_),
    .A(net3459),
    .B(_01648_));
 sg13g2_nor4_2 _07216_ (.A(_01674_),
    .B(_01677_),
    .C(_01678_),
    .Y(_01680_),
    .D(_01679_));
 sg13g2_o21ai_1 _07217_ (.B1(_01680_),
    .Y(_01681_),
    .A1(_01665_),
    .A2(_01673_));
 sg13g2_nand2_1 _07218_ (.Y(_01682_),
    .A(_00595_),
    .B(_01663_));
 sg13g2_nor2_1 _07219_ (.A(net3492),
    .B(_01670_),
    .Y(_01683_));
 sg13g2_nor3_1 _07220_ (.A(_01665_),
    .B(net3038),
    .C(net3031),
    .Y(_01684_));
 sg13g2_and4_2 _07221_ (.A(net3500),
    .B(net3499),
    .C(net3497),
    .D(_01666_),
    .X(_01685_));
 sg13g2_nand4_1 _07222_ (.B(net3499),
    .C(net3497),
    .A(net3500),
    .Y(_01686_),
    .D(_01666_));
 sg13g2_nor2_1 _07223_ (.A(net3496),
    .B(_01686_),
    .Y(_01687_));
 sg13g2_nand2b_1 _07224_ (.Y(_01688_),
    .B(_01685_),
    .A_N(\core.e2m_addr[3] ));
 sg13g2_nor2_1 _07225_ (.A(_01663_),
    .B(net3038),
    .Y(_01689_));
 sg13g2_a22oi_1 _07226_ (.Y(_01690_),
    .B1(net2912),
    .B2(_01689_),
    .A2(_01681_),
    .A1(_01660_));
 sg13g2_nor3_1 _07227_ (.A(\core.e2m_addr[6] ),
    .B(_00597_),
    .C(_01661_),
    .Y(_01691_));
 sg13g2_nand3b_1 _07228_ (.B(_00594_),
    .C(net3495),
    .Y(_01692_),
    .A_N(_01661_));
 sg13g2_nand3_1 _07229_ (.B(_01686_),
    .C(net3195),
    .A(_01682_),
    .Y(_01693_));
 sg13g2_nand2_1 _07230_ (.Y(_01694_),
    .A(net3488),
    .B(_01693_));
 sg13g2_xnor2_1 _07231_ (.Y(_01695_),
    .A(_01651_),
    .B(_01694_));
 sg13g2_nand2_1 _07232_ (.Y(_01696_),
    .A(net3486),
    .B(_01693_));
 sg13g2_a21oi_1 _07233_ (.A1(net3486),
    .A2(_01693_),
    .Y(_01697_),
    .B1(_01653_));
 sg13g2_nand2_1 _07234_ (.Y(_01698_),
    .A(\core.e2m_addr[8] ),
    .B(_01693_));
 sg13g2_xor2_1 _07235_ (.B(_01698_),
    .A(_01648_),
    .X(_01699_));
 sg13g2_nand3_1 _07236_ (.B(_01650_),
    .C(_01651_),
    .A(_01648_),
    .Y(_01700_));
 sg13g2_a22oi_1 _07237_ (.Y(_01701_),
    .B1(_01696_),
    .B2(_01700_),
    .A2(_01647_),
    .A1(\core.lsu.dreg[3] ));
 sg13g2_nand2_1 _07238_ (.Y(_01702_),
    .A(\core.e2m_addr[7] ),
    .B(_01693_));
 sg13g2_xor2_1 _07239_ (.B(_01702_),
    .A(_01650_),
    .X(_01703_));
 sg13g2_nor4_1 _07240_ (.A(_01697_),
    .B(_01699_),
    .C(_01701_),
    .D(_01703_),
    .Y(_01704_));
 sg13g2_a21oi_1 _07241_ (.A1(_01695_),
    .A2(_01704_),
    .Y(_01705_),
    .B1(_01690_));
 sg13g2_nand2b_1 _07242_ (.Y(_01706_),
    .B(net3332),
    .A_N(_01705_));
 sg13g2_and2_2 _07243_ (.A(_01644_),
    .B(_01706_),
    .X(_01707_));
 sg13g2_nand2_1 _07244_ (.Y(_01708_),
    .A(_01644_),
    .B(_01706_));
 sg13g2_nor2b_2 _07245_ (.A(net3502),
    .B_N(net3501),
    .Y(_01709_));
 sg13g2_nand2b_1 _07246_ (.Y(_01710_),
    .B(\core.work.state[1] ),
    .A_N(net3502));
 sg13g2_nor2_2 _07247_ (.A(\core.work.op[4] ),
    .B(\core.work.alu.is_mem ),
    .Y(_01711_));
 sg13g2_and3_2 _07248_ (.X(_01712_),
    .A(net3441),
    .B(\core.work.alu.ls_size_b ),
    .C(_01711_));
 sg13g2_nand3_1 _07249_ (.B(\core.work.alu.ls_size_b ),
    .C(_01711_),
    .A(net3441),
    .Y(_01713_));
 sg13g2_nor2_2 _07250_ (.A(_00629_),
    .B(net3440),
    .Y(_01714_));
 sg13g2_nand2b_1 _07251_ (.Y(_01715_),
    .B(\core.work.alu.is_sign ),
    .A_N(net3440));
 sg13g2_nor2_2 _07252_ (.A(_01713_),
    .B(_01715_),
    .Y(_01716_));
 sg13g2_nand2_2 _07253_ (.Y(_01717_),
    .A(_01712_),
    .B(_01714_));
 sg13g2_and2_2 _07254_ (.A(_01312_),
    .B(_01711_),
    .X(_01718_));
 sg13g2_nand2_1 _07255_ (.Y(_01719_),
    .A(_01312_),
    .B(_01711_));
 sg13g2_and2_2 _07256_ (.A(_01298_),
    .B(_01711_),
    .X(_01720_));
 sg13g2_nand2_1 _07257_ (.Y(_01721_),
    .A(_01308_),
    .B(_01720_));
 sg13g2_o21ai_1 _07258_ (.B1(_01721_),
    .Y(_01722_),
    .A1(_01309_),
    .A2(_01719_));
 sg13g2_nand2b_1 _07259_ (.Y(_01723_),
    .B(_01717_),
    .A_N(_01722_));
 sg13g2_o21ai_1 _07260_ (.B1(_01707_),
    .Y(_01724_),
    .A1(net3298),
    .A2(_01723_));
 sg13g2_and2_2 _07261_ (.A(net3497),
    .B(_01691_),
    .X(_01725_));
 sg13g2_nand2b_1 _07262_ (.Y(_01726_),
    .B(net3331),
    .A_N(net3028));
 sg13g2_nor2_1 _07263_ (.A(net3037),
    .B(_01685_),
    .Y(_01727_));
 sg13g2_nand2_1 _07264_ (.Y(_01728_),
    .A(net3034),
    .B(_01686_));
 sg13g2_mux2_1 _07265_ (.A0(_00033_),
    .A1(_00106_),
    .S(_01665_),
    .X(_01729_));
 sg13g2_a221oi_1 _07266_ (.B2(_01729_),
    .C1(_01669_),
    .B1(_01727_),
    .A1(_00107_),
    .Y(_01730_),
    .A2(_01685_));
 sg13g2_nand2_1 _07267_ (.Y(_01731_),
    .A(net3465),
    .B(\core.work.registers.genblk1[1].latch[1] ));
 sg13g2_nand2_1 _07268_ (.Y(_01732_),
    .A(net3457),
    .B(net3465));
 sg13g2_nand2_2 _07269_ (.Y(_01733_),
    .A(_00617_),
    .B(net3455));
 sg13g2_nor2_1 _07270_ (.A(_01732_),
    .B(_01733_),
    .Y(_01734_));
 sg13g2_nand2_2 _07271_ (.Y(_01735_),
    .A(net3453),
    .B(net3455));
 sg13g2_nand2_2 _07272_ (.Y(_01736_),
    .A(net3457),
    .B(_00622_));
 sg13g2_nor2_1 _07273_ (.A(_01735_),
    .B(_01736_),
    .Y(_01737_));
 sg13g2_nor3_1 _07274_ (.A(net3453),
    .B(net3455),
    .C(_01736_),
    .Y(_01738_));
 sg13g2_nor3_1 _07275_ (.A(net3453),
    .B(net3455),
    .C(_01732_),
    .Y(_01739_));
 sg13g2_nand2_1 _07276_ (.Y(_01740_),
    .A(_00620_),
    .B(net3465));
 sg13g2_nor2_1 _07277_ (.A(_01735_),
    .B(_01740_),
    .Y(_01741_));
 sg13g2_nand2b_1 _07278_ (.Y(_01742_),
    .B(net3453),
    .A_N(net3455));
 sg13g2_nor2_1 _07279_ (.A(_01732_),
    .B(_01742_),
    .Y(_01743_));
 sg13g2_nor2_1 _07280_ (.A(_01733_),
    .B(_01740_),
    .Y(_01744_));
 sg13g2_nor2_1 _07281_ (.A(_01740_),
    .B(_01742_),
    .Y(_01745_));
 sg13g2_nor2_1 _07282_ (.A(_01732_),
    .B(_01735_),
    .Y(_01746_));
 sg13g2_nor3_1 _07283_ (.A(net3457),
    .B(net3465),
    .C(_01742_),
    .Y(_01747_));
 sg13g2_nor2_1 _07284_ (.A(_01733_),
    .B(_01736_),
    .Y(_01748_));
 sg13g2_nor2_1 _07285_ (.A(_01736_),
    .B(_01742_),
    .Y(_01749_));
 sg13g2_nand2_1 _07286_ (.Y(_01750_),
    .A(\core.work.registers.genblk1[10].latch[1] ),
    .B(net2991));
 sg13g2_nor3_1 _07287_ (.A(net3457),
    .B(net3465),
    .C(_01733_),
    .Y(_01751_));
 sg13g2_nor3_1 _07288_ (.A(net3457),
    .B(net3464),
    .C(_01735_),
    .Y(_01752_));
 sg13g2_a22oi_1 _07289_ (.Y(_01753_),
    .B1(net2996),
    .B2(\core.work.registers.genblk1[6].latch[1] ),
    .A2(net3026),
    .A1(\core.work.registers.genblk1[7].latch[1] ));
 sg13g2_a22oi_1 _07290_ (.Y(_01754_),
    .B1(net3001),
    .B2(\core.work.registers.genblk1[9].latch[1] ),
    .A2(net3011),
    .A1(\core.work.registers.genblk1[13].latch[1] ));
 sg13g2_a21oi_1 _07291_ (.A1(\core.work.registers.genblk1[15].latch[1] ),
    .A2(net3182),
    .Y(_01755_),
    .B1(net3319));
 sg13g2_a22oi_1 _07292_ (.Y(_01756_),
    .B1(net2986),
    .B2(\core.work.registers.genblk1[4].latch[1] ),
    .A2(net3187),
    .A1(\core.work.registers.genblk1[11].latch[1] ));
 sg13g2_a22oi_1 _07293_ (.Y(_01757_),
    .B1(net3176),
    .B2(\core.work.registers.genblk1[8].latch[1] ),
    .A2(net3016),
    .A1(\core.work.registers.genblk1[2].latch[1] ));
 sg13g2_nand4_1 _07294_ (.B(_01755_),
    .C(_01756_),
    .A(_01753_),
    .Y(_01758_),
    .D(_01757_));
 sg13g2_a22oi_1 _07295_ (.Y(_01759_),
    .B1(net3006),
    .B2(\core.work.registers.genblk1[5].latch[1] ),
    .A2(net3192),
    .A1(\core.work.registers.genblk1[3].latch[1] ));
 sg13g2_a22oi_1 _07296_ (.Y(_01760_),
    .B1(net3172),
    .B2(\core.work.registers.genblk1[12].latch[1] ),
    .A2(net3021),
    .A1(\core.work.registers.genblk1[14].latch[1] ));
 sg13g2_nand4_1 _07297_ (.B(_01754_),
    .C(_01759_),
    .A(_01750_),
    .Y(_01761_),
    .D(_01760_));
 sg13g2_nor2_1 _07298_ (.A(_01758_),
    .B(_01761_),
    .Y(_01762_));
 sg13g2_a21oi_2 _07299_ (.B1(_01762_),
    .Y(_01763_),
    .A2(_01731_),
    .A1(net3319));
 sg13g2_o21ai_1 _07300_ (.B1(_01763_),
    .Y(_01764_),
    .A1(_01671_),
    .A2(_01730_));
 sg13g2_a22oi_1 _07301_ (.Y(_01765_),
    .B1(_01730_),
    .B2(net3035),
    .A2(net2923),
    .A1(_00640_));
 sg13g2_a21oi_1 _07302_ (.A1(_01764_),
    .A2(_01765_),
    .Y(_01766_),
    .B1(net2910));
 sg13g2_nor2_1 _07303_ (.A(net3331),
    .B(net3303),
    .Y(_01767_));
 sg13g2_nand2_1 _07304_ (.Y(_01768_),
    .A(net3329),
    .B(net3298));
 sg13g2_a221oi_1 _07305_ (.B2(\core.f2e_addr[1] ),
    .C1(_01766_),
    .B1(net3167),
    .A1(_00590_),
    .Y(_01769_),
    .A2(net3308));
 sg13g2_nand2_1 _07306_ (.Y(_01770_),
    .A(net3561),
    .B(net2778));
 sg13g2_o21ai_1 _07307_ (.B1(_01770_),
    .Y(_00265_),
    .A1(net2778),
    .A2(_01769_));
 sg13g2_nand2_1 _07308_ (.Y(_01771_),
    .A(net3464),
    .B(\core.work.registers.genblk1[1].latch[2] ));
 sg13g2_nand2_1 _07309_ (.Y(_01772_),
    .A(\core.work.registers.genblk1[8].latch[2] ),
    .B(net3176));
 sg13g2_a22oi_1 _07310_ (.Y(_01773_),
    .B1(net2996),
    .B2(\core.work.registers.genblk1[6].latch[2] ),
    .A2(net3182),
    .A1(\core.work.registers.genblk1[15].latch[2] ));
 sg13g2_a21oi_1 _07311_ (.A1(\core.work.registers.genblk1[4].latch[2] ),
    .A2(net2986),
    .Y(_01774_),
    .B1(net3318));
 sg13g2_a22oi_1 _07312_ (.Y(_01775_),
    .B1(net3171),
    .B2(\core.work.registers.genblk1[12].latch[2] ),
    .A2(net3021),
    .A1(\core.work.registers.genblk1[14].latch[2] ));
 sg13g2_a22oi_1 _07313_ (.Y(_01776_),
    .B1(net3186),
    .B2(\core.work.registers.genblk1[11].latch[2] ),
    .A2(net3191),
    .A1(\core.work.registers.genblk1[3].latch[2] ));
 sg13g2_nand4_1 _07314_ (.B(_01774_),
    .C(_01775_),
    .A(_01773_),
    .Y(_01777_),
    .D(_01776_));
 sg13g2_a22oi_1 _07315_ (.Y(_01778_),
    .B1(net2991),
    .B2(\core.work.registers.genblk1[10].latch[2] ),
    .A2(net3005),
    .A1(\core.work.registers.genblk1[5].latch[2] ));
 sg13g2_a22oi_1 _07316_ (.Y(_01779_),
    .B1(net3000),
    .B2(\core.work.registers.genblk1[9].latch[2] ),
    .A2(net3025),
    .A1(\core.work.registers.genblk1[7].latch[2] ));
 sg13g2_a22oi_1 _07317_ (.Y(_01780_),
    .B1(net3011),
    .B2(\core.work.registers.genblk1[13].latch[2] ),
    .A2(net3015),
    .A1(\core.work.registers.genblk1[2].latch[2] ));
 sg13g2_nand4_1 _07318_ (.B(_01778_),
    .C(_01779_),
    .A(_01772_),
    .Y(_01781_),
    .D(_01780_));
 sg13g2_nor2_1 _07319_ (.A(_01777_),
    .B(_01781_),
    .Y(_01782_));
 sg13g2_a21oi_2 _07320_ (.B1(_01782_),
    .Y(_01783_),
    .A2(_01771_),
    .A1(net3317));
 sg13g2_mux2_1 _07321_ (.A0(_00036_),
    .A1(_00108_),
    .S(_01665_),
    .X(_01784_));
 sg13g2_a221oi_1 _07322_ (.B2(_01784_),
    .C1(_01669_),
    .B1(_01727_),
    .A1(\core.work.inst_was_short ),
    .Y(_01785_),
    .A2(_01685_));
 sg13g2_o21ai_1 _07323_ (.B1(_01783_),
    .Y(_01786_),
    .A1(_01671_),
    .A2(_01785_));
 sg13g2_a22oi_1 _07324_ (.Y(_01787_),
    .B1(_01785_),
    .B2(net3035),
    .A2(net2923),
    .A1(_00642_));
 sg13g2_a21oi_1 _07325_ (.A1(_01786_),
    .A2(_01787_),
    .Y(_01788_),
    .B1(net2910));
 sg13g2_xor2_1 _07326_ (.B(net3557),
    .A(net3561),
    .X(_01789_));
 sg13g2_a21oi_2 _07327_ (.B1(_01788_),
    .Y(_01790_),
    .A2(net3168),
    .A1(\core.f2e_addr[2] ));
 sg13g2_o21ai_1 _07328_ (.B1(_01790_),
    .Y(_01791_),
    .A1(net3302),
    .A2(_01789_));
 sg13g2_mux2_1 _07329_ (.A0(_01791_),
    .A1(net3557),
    .S(net2777),
    .X(_00266_));
 sg13g2_nand2_1 _07330_ (.Y(_01792_),
    .A(net3554),
    .B(net2777));
 sg13g2_nand2_1 _07331_ (.Y(_01793_),
    .A(net3464),
    .B(\core.work.registers.genblk1[1].latch[3] ));
 sg13g2_a22oi_1 _07332_ (.Y(_01794_),
    .B1(net3182),
    .B2(\core.work.registers.genblk1[15].latch[3] ),
    .A2(net3187),
    .A1(\core.work.registers.genblk1[11].latch[3] ));
 sg13g2_nand2_1 _07333_ (.Y(_01795_),
    .A(\core.work.registers.genblk1[6].latch[3] ),
    .B(net2995));
 sg13g2_a22oi_1 _07334_ (.Y(_01796_),
    .B1(net3001),
    .B2(\core.work.registers.genblk1[9].latch[3] ),
    .A2(net3191),
    .A1(\core.work.registers.genblk1[3].latch[3] ));
 sg13g2_a21oi_1 _07335_ (.A1(\core.work.registers.genblk1[4].latch[3] ),
    .A2(net2986),
    .Y(_01797_),
    .B1(net3317));
 sg13g2_a22oi_1 _07336_ (.Y(_01798_),
    .B1(net2990),
    .B2(\core.work.registers.genblk1[10].latch[3] ),
    .A2(net3021),
    .A1(\core.work.registers.genblk1[14].latch[3] ));
 sg13g2_nand4_1 _07337_ (.B(_01796_),
    .C(_01797_),
    .A(_01794_),
    .Y(_01799_),
    .D(_01798_));
 sg13g2_a22oi_1 _07338_ (.Y(_01800_),
    .B1(net3006),
    .B2(\core.work.registers.genblk1[5].latch[3] ),
    .A2(net3015),
    .A1(\core.work.registers.genblk1[2].latch[3] ));
 sg13g2_a22oi_1 _07339_ (.Y(_01801_),
    .B1(net3176),
    .B2(\core.work.registers.genblk1[8].latch[3] ),
    .A2(net3026),
    .A1(\core.work.registers.genblk1[7].latch[3] ));
 sg13g2_a22oi_1 _07340_ (.Y(_01802_),
    .B1(net3172),
    .B2(\core.work.registers.genblk1[12].latch[3] ),
    .A2(net3011),
    .A1(\core.work.registers.genblk1[13].latch[3] ));
 sg13g2_nand4_1 _07341_ (.B(_01800_),
    .C(_01801_),
    .A(_01795_),
    .Y(_01803_),
    .D(_01802_));
 sg13g2_nor2_1 _07342_ (.A(_01799_),
    .B(_01803_),
    .Y(_01804_));
 sg13g2_a21oi_2 _07343_ (.B1(_01804_),
    .Y(_01805_),
    .A2(_01793_),
    .A1(net3317));
 sg13g2_nor2b_1 _07344_ (.A(_01665_),
    .B_N(_00038_),
    .Y(_01806_));
 sg13g2_a21oi_1 _07345_ (.A1(_00110_),
    .A2(_01665_),
    .Y(_01807_),
    .B1(_01806_));
 sg13g2_nand2_1 _07346_ (.Y(_01808_),
    .A(net3452),
    .B(net2923));
 sg13g2_a221oi_1 _07347_ (.B2(net2908),
    .C1(net3031),
    .B1(_01807_),
    .A1(net3037),
    .Y(_01809_),
    .A2(_01805_));
 sg13g2_o21ai_1 _07348_ (.B1(_01808_),
    .Y(_01810_),
    .A1(_01672_),
    .A2(_01805_));
 sg13g2_nor3_1 _07349_ (.A(net2910),
    .B(_01809_),
    .C(_01810_),
    .Y(_01811_));
 sg13g2_nor2_1 _07350_ (.A(net3559),
    .B(net3551),
    .Y(_01812_));
 sg13g2_o21ai_1 _07351_ (.B1(_00109_),
    .Y(_01813_),
    .A1(net3562),
    .A2(net3559));
 sg13g2_a21oi_1 _07352_ (.A1(_00590_),
    .A2(net3296),
    .Y(_01814_),
    .B1(net3301));
 sg13g2_a221oi_1 _07353_ (.B2(_01814_),
    .C1(_01811_),
    .B1(_01813_),
    .A1(net622),
    .Y(_01815_),
    .A2(net3167));
 sg13g2_o21ai_1 _07354_ (.B1(_01792_),
    .Y(_00267_),
    .A1(net2777),
    .A2(_01815_));
 sg13g2_a21oi_1 _07355_ (.A1(_00040_),
    .A2(net2923),
    .Y(_01816_),
    .B1(net2910));
 sg13g2_nand2_1 _07356_ (.Y(_01817_),
    .A(net3464),
    .B(\core.work.registers.genblk1[1].latch[4] ));
 sg13g2_nand2_1 _07357_ (.Y(_01818_),
    .A(\core.work.registers.genblk1[11].latch[4] ),
    .B(net3187));
 sg13g2_a22oi_1 _07358_ (.Y(_01819_),
    .B1(net2991),
    .B2(\core.work.registers.genblk1[10].latch[4] ),
    .A2(net3016),
    .A1(\core.work.registers.genblk1[2].latch[4] ));
 sg13g2_a22oi_1 _07359_ (.Y(_01820_),
    .B1(net2985),
    .B2(\core.work.registers.genblk1[4].latch[4] ),
    .A2(net3181),
    .A1(\core.work.registers.genblk1[15].latch[4] ));
 sg13g2_a21oi_1 _07360_ (.A1(\core.work.registers.genblk1[14].latch[4] ),
    .A2(net3021),
    .Y(_01821_),
    .B1(net3317));
 sg13g2_a22oi_1 _07361_ (.Y(_01822_),
    .B1(net2996),
    .B2(\core.work.registers.genblk1[6].latch[4] ),
    .A2(net3010),
    .A1(\core.work.registers.genblk1[13].latch[4] ));
 sg13g2_nand3_1 _07362_ (.B(_01821_),
    .C(_01822_),
    .A(_01819_),
    .Y(_01823_));
 sg13g2_a221oi_1 _07363_ (.B2(\core.work.registers.genblk1[9].latch[4] ),
    .C1(_01823_),
    .B1(net3001),
    .A1(\core.work.registers.genblk1[5].latch[4] ),
    .Y(_01824_),
    .A2(net3006));
 sg13g2_a22oi_1 _07364_ (.Y(_01825_),
    .B1(net3172),
    .B2(\core.work.registers.genblk1[12].latch[4] ),
    .A2(net3176),
    .A1(\core.work.registers.genblk1[8].latch[4] ));
 sg13g2_nand3_1 _07365_ (.B(_01820_),
    .C(_01825_),
    .A(_01818_),
    .Y(_01826_));
 sg13g2_a221oi_1 _07366_ (.B2(\core.work.registers.genblk1[3].latch[4] ),
    .C1(_01826_),
    .B1(net3192),
    .A1(\core.work.registers.genblk1[7].latch[4] ),
    .Y(_01827_),
    .A2(net3026));
 sg13g2_a22oi_1 _07367_ (.Y(_01828_),
    .B1(_01824_),
    .B2(_01827_),
    .A2(_01817_),
    .A1(net3319));
 sg13g2_mux2_1 _07368_ (.A0(_00040_),
    .A1(_00111_),
    .S(_01665_),
    .X(_01829_));
 sg13g2_o21ai_1 _07369_ (.B1(_01670_),
    .Y(_01830_),
    .A1(net2906),
    .A2(_01829_));
 sg13g2_a21oi_1 _07370_ (.A1(_01672_),
    .A2(_01830_),
    .Y(_01831_),
    .B1(_01828_));
 sg13g2_o21ai_1 _07371_ (.B1(_01816_),
    .Y(_01832_),
    .A1(net3037),
    .A2(_01830_));
 sg13g2_nor2_1 _07372_ (.A(net3553),
    .B(net3557),
    .Y(_01833_));
 sg13g2_or2_2 _07373_ (.X(_01834_),
    .B(net3558),
    .A(net3552));
 sg13g2_nor2_1 _07374_ (.A(net3562),
    .B(_01834_),
    .Y(_01835_));
 sg13g2_xnor2_1 _07375_ (.Y(_01836_),
    .A(net3544),
    .B(_01835_));
 sg13g2_a22oi_1 _07376_ (.Y(_01837_),
    .B1(_01836_),
    .B2(net3308),
    .A2(net3167),
    .A1(net3564));
 sg13g2_o21ai_1 _07377_ (.B1(_01837_),
    .Y(_01838_),
    .A1(_01831_),
    .A2(_01832_));
 sg13g2_nor2_1 _07378_ (.A(net2778),
    .B(_01838_),
    .Y(_01839_));
 sg13g2_a21oi_1 _07379_ (.A1(_00596_),
    .A2(net2778),
    .Y(_00268_),
    .B1(_01839_));
 sg13g2_nand2_1 _07380_ (.Y(_01840_),
    .A(net3462),
    .B(\core.work.registers.genblk1[1].latch[5] ));
 sg13g2_nand2_1 _07381_ (.Y(_01841_),
    .A(\core.work.registers.genblk1[14].latch[5] ),
    .B(net3019));
 sg13g2_a21oi_1 _07382_ (.A1(\core.work.registers.genblk1[6].latch[5] ),
    .A2(net2994),
    .Y(_01842_),
    .B1(net3313));
 sg13g2_a22oi_1 _07383_ (.Y(_01843_),
    .B1(net3009),
    .B2(\core.work.registers.genblk1[13].latch[5] ),
    .A2(net3017),
    .A1(\core.work.registers.genblk1[2].latch[5] ));
 sg13g2_a22oi_1 _07384_ (.Y(_01844_),
    .B1(net2984),
    .B2(\core.work.registers.genblk1[4].latch[5] ),
    .A2(net2999),
    .A1(\core.work.registers.genblk1[9].latch[5] ));
 sg13g2_a22oi_1 _07385_ (.Y(_01845_),
    .B1(net3175),
    .B2(\core.work.registers.genblk1[8].latch[5] ),
    .A2(net3004),
    .A1(\core.work.registers.genblk1[5].latch[5] ));
 sg13g2_nand4_1 _07386_ (.B(_01843_),
    .C(_01844_),
    .A(_01842_),
    .Y(_01846_),
    .D(_01845_));
 sg13g2_a22oi_1 _07387_ (.Y(_01847_),
    .B1(net3185),
    .B2(\core.work.registers.genblk1[11].latch[5] ),
    .A2(net3190),
    .A1(\core.work.registers.genblk1[3].latch[5] ));
 sg13g2_a22oi_1 _07388_ (.Y(_01848_),
    .B1(net2989),
    .B2(\core.work.registers.genblk1[10].latch[5] ),
    .A2(net3027),
    .A1(\core.work.registers.genblk1[7].latch[5] ));
 sg13g2_a22oi_1 _07389_ (.Y(_01849_),
    .B1(net3170),
    .B2(\core.work.registers.genblk1[12].latch[5] ),
    .A2(net3180),
    .A1(\core.work.registers.genblk1[15].latch[5] ));
 sg13g2_nand4_1 _07390_ (.B(_01847_),
    .C(_01848_),
    .A(_01841_),
    .Y(_01850_),
    .D(_01849_));
 sg13g2_nor2_2 _07391_ (.A(_01846_),
    .B(_01850_),
    .Y(_01851_));
 sg13g2_a21oi_2 _07392_ (.B1(_01851_),
    .Y(_01852_),
    .A2(_01840_),
    .A1(net3315));
 sg13g2_nand2_1 _07393_ (.Y(_01853_),
    .A(net3037),
    .B(_01852_));
 sg13g2_o21ai_1 _07394_ (.B1(_01670_),
    .Y(_01854_),
    .A1(_00041_),
    .A2(net2905));
 sg13g2_o21ai_1 _07395_ (.B1(_01854_),
    .Y(_01855_),
    .A1(_01672_),
    .A2(_01852_));
 sg13g2_a221oi_1 _07396_ (.B2(_01855_),
    .C1(net2911),
    .B1(_01853_),
    .A1(_00041_),
    .Y(_01856_),
    .A2(net2922));
 sg13g2_nor3_1 _07397_ (.A(net3562),
    .B(net3548),
    .C(_01834_),
    .Y(_01857_));
 sg13g2_xnor2_1 _07398_ (.Y(_01858_),
    .A(_00112_),
    .B(_01857_));
 sg13g2_a221oi_1 _07399_ (.B2(net3308),
    .C1(_01856_),
    .B1(_01858_),
    .A1(\core.f2e_addr[5] ),
    .Y(_01859_),
    .A2(net3167));
 sg13g2_nand2_1 _07400_ (.Y(_01860_),
    .A(net3543),
    .B(net2777));
 sg13g2_o21ai_1 _07401_ (.B1(_01860_),
    .Y(_00269_),
    .A1(net2777),
    .A2(_01859_));
 sg13g2_nand2_1 _07402_ (.Y(_01861_),
    .A(net3464),
    .B(\core.work.registers.genblk1[1].latch[6] ));
 sg13g2_nand2_1 _07403_ (.Y(_01862_),
    .A(\core.work.registers.genblk1[14].latch[6] ),
    .B(net3021));
 sg13g2_a22oi_1 _07404_ (.Y(_01863_),
    .B1(net2991),
    .B2(\core.work.registers.genblk1[10].latch[6] ),
    .A2(net3006),
    .A1(\core.work.registers.genblk1[5].latch[6] ));
 sg13g2_a21oi_1 _07405_ (.A1(\core.work.registers.genblk1[7].latch[6] ),
    .A2(net3026),
    .Y(_01864_),
    .B1(net3318));
 sg13g2_a22oi_1 _07406_ (.Y(_01865_),
    .B1(net3182),
    .B2(\core.work.registers.genblk1[15].latch[6] ),
    .A2(net3192),
    .A1(\core.work.registers.genblk1[3].latch[6] ));
 sg13g2_a22oi_1 _07407_ (.Y(_01866_),
    .B1(net2986),
    .B2(\core.work.registers.genblk1[4].latch[6] ),
    .A2(net3177),
    .A1(\core.work.registers.genblk1[8].latch[6] ));
 sg13g2_nand4_1 _07408_ (.B(_01864_),
    .C(_01865_),
    .A(_01863_),
    .Y(_01867_),
    .D(_01866_));
 sg13g2_a22oi_1 _07409_ (.Y(_01868_),
    .B1(net2996),
    .B2(\core.work.registers.genblk1[6].latch[6] ),
    .A2(net3187),
    .A1(\core.work.registers.genblk1[11].latch[6] ));
 sg13g2_a22oi_1 _07410_ (.Y(_01869_),
    .B1(net3172),
    .B2(\core.work.registers.genblk1[12].latch[6] ),
    .A2(net3001),
    .A1(\core.work.registers.genblk1[9].latch[6] ));
 sg13g2_a22oi_1 _07411_ (.Y(_01870_),
    .B1(net3011),
    .B2(\core.work.registers.genblk1[13].latch[6] ),
    .A2(net3016),
    .A1(\core.work.registers.genblk1[2].latch[6] ));
 sg13g2_nand4_1 _07412_ (.B(_01868_),
    .C(_01869_),
    .A(_01862_),
    .Y(_01871_),
    .D(_01870_));
 sg13g2_nor2_1 _07413_ (.A(_01867_),
    .B(_01871_),
    .Y(_01872_));
 sg13g2_a21oi_2 _07414_ (.B1(_01872_),
    .Y(_01873_),
    .A2(_01861_),
    .A1(net3317));
 sg13g2_a21oi_1 _07415_ (.A1(_00044_),
    .A2(_01670_),
    .Y(_01874_),
    .B1(net2906));
 sg13g2_a21oi_1 _07416_ (.A1(_01672_),
    .A2(_01874_),
    .Y(_01875_),
    .B1(_01873_));
 sg13g2_a21oi_1 _07417_ (.A1(_00044_),
    .A2(net2922),
    .Y(_01876_),
    .B1(net2910));
 sg13g2_o21ai_1 _07418_ (.B1(_01876_),
    .Y(_01877_),
    .A1(net3037),
    .A2(_01874_));
 sg13g2_nor4_2 _07419_ (.A(net3562),
    .B(net3543),
    .C(net3549),
    .Y(_01878_),
    .D(_01834_));
 sg13g2_xnor2_1 _07420_ (.Y(_01879_),
    .A(_00113_),
    .B(_01878_));
 sg13g2_a22oi_1 _07421_ (.Y(_01880_),
    .B1(_01879_),
    .B2(net3308),
    .A2(net3167),
    .A1(\core.f2e_addr[6] ));
 sg13g2_o21ai_1 _07422_ (.B1(_01880_),
    .Y(_01881_),
    .A1(_01875_),
    .A2(_01877_));
 sg13g2_mux2_1 _07423_ (.A0(_01881_),
    .A1(net842),
    .S(net2777),
    .X(_00270_));
 sg13g2_nor2_2 _07424_ (.A(_01671_),
    .B(net2907),
    .Y(_01882_));
 sg13g2_nand2_1 _07425_ (.Y(_01883_),
    .A(net3464),
    .B(\core.work.registers.genblk1[1].latch[7] ));
 sg13g2_nand2_1 _07426_ (.Y(_01884_),
    .A(\core.work.registers.genblk1[13].latch[7] ),
    .B(net3010));
 sg13g2_a21oi_1 _07427_ (.A1(\core.work.registers.genblk1[9].latch[7] ),
    .A2(net3000),
    .Y(_01885_),
    .B1(net3315));
 sg13g2_a22oi_1 _07428_ (.Y(_01886_),
    .B1(net2995),
    .B2(\core.work.registers.genblk1[6].latch[7] ),
    .A2(net3025),
    .A1(\core.work.registers.genblk1[7].latch[7] ));
 sg13g2_a22oi_1 _07429_ (.Y(_01887_),
    .B1(net2985),
    .B2(\core.work.registers.genblk1[4].latch[7] ),
    .A2(net3020),
    .A1(\core.work.registers.genblk1[14].latch[7] ));
 sg13g2_nand3_1 _07430_ (.B(_01886_),
    .C(_01887_),
    .A(_01885_),
    .Y(_01888_));
 sg13g2_a221oi_1 _07431_ (.B2(\core.work.registers.genblk1[12].latch[7] ),
    .C1(_01888_),
    .B1(net3171),
    .A1(\core.work.registers.genblk1[3].latch[7] ),
    .Y(_01889_),
    .A2(net3191));
 sg13g2_a22oi_1 _07432_ (.Y(_01890_),
    .B1(net3182),
    .B2(\core.work.registers.genblk1[15].latch[7] ),
    .A2(net3187),
    .A1(\core.work.registers.genblk1[11].latch[7] ));
 sg13g2_a22oi_1 _07433_ (.Y(_01891_),
    .B1(net2990),
    .B2(\core.work.registers.genblk1[10].latch[7] ),
    .A2(net3005),
    .A1(\core.work.registers.genblk1[5].latch[7] ));
 sg13g2_nand3_1 _07434_ (.B(_01890_),
    .C(_01891_),
    .A(_01884_),
    .Y(_01892_));
 sg13g2_a221oi_1 _07435_ (.B2(\core.work.registers.genblk1[8].latch[7] ),
    .C1(_01892_),
    .B1(net3176),
    .A1(\core.work.registers.genblk1[2].latch[7] ),
    .Y(_01893_),
    .A2(net3016));
 sg13g2_a22oi_1 _07436_ (.Y(_01894_),
    .B1(_01889_),
    .B2(_01893_),
    .A2(_01883_),
    .A1(net3317));
 sg13g2_a22oi_1 _07437_ (.Y(_01895_),
    .B1(_01894_),
    .B2(_01673_),
    .A2(_01882_),
    .A1(_00645_));
 sg13g2_nor2b_1 _07438_ (.A(\core.work.alu.sval2[6] ),
    .B_N(_01878_),
    .Y(_01896_));
 sg13g2_xnor2_1 _07439_ (.Y(_01897_),
    .A(_00114_),
    .B(_01896_));
 sg13g2_a21oi_1 _07440_ (.A1(net3308),
    .A2(_01897_),
    .Y(_01898_),
    .B1(net3167));
 sg13g2_o21ai_1 _07441_ (.B1(_01898_),
    .Y(_01899_),
    .A1(net2910),
    .A2(_01895_));
 sg13g2_o21ai_1 _07442_ (.B1(_01899_),
    .Y(_01900_),
    .A1(net3563),
    .A2(net3161));
 sg13g2_nand2_1 _07443_ (.Y(_01901_),
    .A(net699),
    .B(net2777));
 sg13g2_o21ai_1 _07444_ (.B1(_01901_),
    .Y(_00271_),
    .A1(net2777),
    .A2(_01900_));
 sg13g2_nand2_1 _07445_ (.Y(_01902_),
    .A(net3462),
    .B(\core.work.registers.genblk1[1].latch[8] ));
 sg13g2_nand2_1 _07446_ (.Y(_01903_),
    .A(\core.work.registers.genblk1[8].latch[8] ),
    .B(net3175));
 sg13g2_a21oi_1 _07447_ (.A1(\core.work.registers.genblk1[6].latch[8] ),
    .A2(net2994),
    .Y(_01904_),
    .B1(net3314));
 sg13g2_a22oi_1 _07448_ (.Y(_01905_),
    .B1(net2984),
    .B2(\core.work.registers.genblk1[4].latch[8] ),
    .A2(net3024),
    .A1(\core.work.registers.genblk1[7].latch[8] ));
 sg13g2_a22oi_1 _07449_ (.Y(_01906_),
    .B1(net2999),
    .B2(\core.work.registers.genblk1[9].latch[8] ),
    .A2(net3188),
    .A1(\core.work.registers.genblk1[11].latch[8] ));
 sg13g2_nand3_1 _07450_ (.B(_01905_),
    .C(_01906_),
    .A(_01904_),
    .Y(_01907_));
 sg13g2_a221oi_1 _07451_ (.B2(\core.work.registers.genblk1[3].latch[8] ),
    .C1(_01907_),
    .B1(net3190),
    .A1(\core.work.registers.genblk1[2].latch[8] ),
    .Y(_01908_),
    .A2(net3014));
 sg13g2_a22oi_1 _07452_ (.Y(_01909_),
    .B1(net3170),
    .B2(\core.work.registers.genblk1[12].latch[8] ),
    .A2(net3009),
    .A1(\core.work.registers.genblk1[13].latch[8] ));
 sg13g2_a22oi_1 _07453_ (.Y(_01910_),
    .B1(net3183),
    .B2(\core.work.registers.genblk1[15].latch[8] ),
    .A2(net3004),
    .A1(\core.work.registers.genblk1[5].latch[8] ));
 sg13g2_nand3_1 _07454_ (.B(_01909_),
    .C(_01910_),
    .A(_01903_),
    .Y(_01911_));
 sg13g2_a221oi_1 _07455_ (.B2(\core.work.registers.genblk1[10].latch[8] ),
    .C1(_01911_),
    .B1(net2989),
    .A1(\core.work.registers.genblk1[14].latch[8] ),
    .Y(_01912_),
    .A2(net3020));
 sg13g2_a22oi_1 _07456_ (.Y(_01913_),
    .B1(_01908_),
    .B2(_01912_),
    .A2(_01902_),
    .A1(net3314));
 sg13g2_a22oi_1 _07457_ (.Y(_01914_),
    .B1(_01913_),
    .B2(_01673_),
    .A2(_01882_),
    .A1(_00646_));
 sg13g2_nor2b_2 _07458_ (.A(\core.work.alu.sval2[7] ),
    .B_N(_01896_),
    .Y(_01915_));
 sg13g2_xnor2_1 _07459_ (.Y(_01916_),
    .A(_00115_),
    .B(_01915_));
 sg13g2_a21oi_1 _07460_ (.A1(net3306),
    .A2(_01916_),
    .Y(_01917_),
    .B1(net3166));
 sg13g2_o21ai_1 _07461_ (.B1(_01917_),
    .Y(_01918_),
    .A1(net2910),
    .A2(_01914_));
 sg13g2_o21ai_1 _07462_ (.B1(_01918_),
    .Y(_01919_),
    .A1(\core.f2e_addr[8] ),
    .A2(net3161));
 sg13g2_nand2_1 _07463_ (.Y(_01920_),
    .A(net702),
    .B(net2774));
 sg13g2_o21ai_1 _07464_ (.B1(_01920_),
    .Y(_00272_),
    .A1(net2780),
    .A2(_01919_));
 sg13g2_nand2_1 _07465_ (.Y(_01921_),
    .A(net3467),
    .B(\core.work.registers.genblk1[1].latch[9] ));
 sg13g2_a22oi_1 _07466_ (.Y(_01922_),
    .B1(net2990),
    .B2(\core.work.registers.genblk1[10].latch[9] ),
    .A2(net2995),
    .A1(\core.work.registers.genblk1[6].latch[9] ));
 sg13g2_nand2_1 _07467_ (.Y(_01923_),
    .A(\core.work.registers.genblk1[8].latch[9] ),
    .B(net3177));
 sg13g2_a21oi_1 _07468_ (.A1(\core.work.registers.genblk1[9].latch[9] ),
    .A2(net3000),
    .Y(_01924_),
    .B1(net3316));
 sg13g2_a22oi_1 _07469_ (.Y(_01925_),
    .B1(net3010),
    .B2(\core.work.registers.genblk1[13].latch[9] ),
    .A2(net3020),
    .A1(\core.work.registers.genblk1[14].latch[9] ));
 sg13g2_nand3_1 _07470_ (.B(_01924_),
    .C(_01925_),
    .A(_01922_),
    .Y(_01926_));
 sg13g2_a221oi_1 _07471_ (.B2(\core.work.registers.genblk1[4].latch[9] ),
    .C1(_01926_),
    .B1(net2985),
    .A1(\core.work.registers.genblk1[2].latch[9] ),
    .Y(_01927_),
    .A2(net3015));
 sg13g2_a22oi_1 _07472_ (.Y(_01928_),
    .B1(net3171),
    .B2(\core.work.registers.genblk1[12].latch[9] ),
    .A2(net3005),
    .A1(\core.work.registers.genblk1[5].latch[9] ));
 sg13g2_a22oi_1 _07473_ (.Y(_01929_),
    .B1(net3181),
    .B2(\core.work.registers.genblk1[15].latch[9] ),
    .A2(net3025),
    .A1(\core.work.registers.genblk1[7].latch[9] ));
 sg13g2_nand3_1 _07474_ (.B(_01928_),
    .C(_01929_),
    .A(_01923_),
    .Y(_01930_));
 sg13g2_a221oi_1 _07475_ (.B2(\core.work.registers.genblk1[11].latch[9] ),
    .C1(_01930_),
    .B1(net3186),
    .A1(\core.work.registers.genblk1[3].latch[9] ),
    .Y(_01931_),
    .A2(net3191));
 sg13g2_a22oi_1 _07476_ (.Y(_01932_),
    .B1(_01927_),
    .B2(_01931_),
    .A2(_01921_),
    .A1(net3316));
 sg13g2_a22oi_1 _07477_ (.Y(_01933_),
    .B1(_01932_),
    .B2(_01673_),
    .A2(_01882_),
    .A1(_00647_));
 sg13g2_nand2b_2 _07478_ (.Y(_01934_),
    .B(_01915_),
    .A_N(\core.work.alu.sval2[8] ));
 sg13g2_xnor2_1 _07479_ (.Y(_01935_),
    .A(_00720_),
    .B(_01934_));
 sg13g2_a22oi_1 _07480_ (.Y(_01936_),
    .B1(_01935_),
    .B2(net3306),
    .A2(net3166),
    .A1(\core.f2e_addr[9] ));
 sg13g2_o21ai_1 _07481_ (.B1(_01936_),
    .Y(_01937_),
    .A1(net2911),
    .A2(_01933_));
 sg13g2_mux2_1 _07482_ (.A0(_01937_),
    .A1(net3542),
    .S(net2774),
    .X(_00273_));
 sg13g2_nor2_1 _07483_ (.A(net3542),
    .B(_01934_),
    .Y(_01938_));
 sg13g2_xnor2_1 _07484_ (.Y(_01939_),
    .A(_00117_),
    .B(_01938_));
 sg13g2_nand2_1 _07485_ (.Y(_01940_),
    .A(net3463),
    .B(\core.work.registers.genblk1[1].latch[10] ));
 sg13g2_a22oi_1 _07486_ (.Y(_01941_),
    .B1(net2997),
    .B2(\core.work.registers.genblk1[6].latch[10] ),
    .A2(net3017),
    .A1(\core.work.registers.genblk1[2].latch[10] ));
 sg13g2_nand2_1 _07487_ (.Y(_01942_),
    .A(\core.work.registers.genblk1[4].latch[10] ),
    .B(net2987));
 sg13g2_a22oi_1 _07488_ (.Y(_01943_),
    .B1(net3178),
    .B2(\core.work.registers.genblk1[8].latch[10] ),
    .A2(net3193),
    .A1(\core.work.registers.genblk1[3].latch[10] ));
 sg13g2_a22oi_1 _07489_ (.Y(_01944_),
    .B1(net3173),
    .B2(\core.work.registers.genblk1[12].latch[10] ),
    .A2(net3183),
    .A1(\core.work.registers.genblk1[15].latch[10] ));
 sg13g2_a21oi_1 _07490_ (.A1(\core.work.registers.genblk1[11].latch[10] ),
    .A2(net3188),
    .Y(_01945_),
    .B1(net3320));
 sg13g2_a22oi_1 _07491_ (.Y(_01946_),
    .B1(net3022),
    .B2(\core.work.registers.genblk1[14].latch[10] ),
    .A2(net3027),
    .A1(\core.work.registers.genblk1[7].latch[10] ));
 sg13g2_nand4_1 _07492_ (.B(_01944_),
    .C(_01945_),
    .A(_01941_),
    .Y(_01947_),
    .D(_01946_));
 sg13g2_a22oi_1 _07493_ (.Y(_01948_),
    .B1(net2992),
    .B2(\core.work.registers.genblk1[10].latch[10] ),
    .A2(net3002),
    .A1(\core.work.registers.genblk1[9].latch[10] ));
 sg13g2_a22oi_1 _07494_ (.Y(_01949_),
    .B1(net3007),
    .B2(\core.work.registers.genblk1[5].latch[10] ),
    .A2(net3012),
    .A1(\core.work.registers.genblk1[13].latch[10] ));
 sg13g2_nand4_1 _07495_ (.B(_01943_),
    .C(_01948_),
    .A(_01942_),
    .Y(_01950_),
    .D(_01949_));
 sg13g2_nor2_1 _07496_ (.A(_01947_),
    .B(_01950_),
    .Y(_01951_));
 sg13g2_a21oi_2 _07497_ (.B1(_01951_),
    .Y(_01952_),
    .A2(_01940_),
    .A1(net3314));
 sg13g2_a22oi_1 _07498_ (.Y(_01953_),
    .B1(_01952_),
    .B2(_01673_),
    .A2(_01882_),
    .A1(_00648_));
 sg13g2_a22oi_1 _07499_ (.Y(_01954_),
    .B1(_01939_),
    .B2(net3306),
    .A2(net3166),
    .A1(net759));
 sg13g2_o21ai_1 _07500_ (.B1(_01954_),
    .Y(_01955_),
    .A1(net2909),
    .A2(_01953_));
 sg13g2_nor2_1 _07501_ (.A(net2774),
    .B(_01955_),
    .Y(_01956_));
 sg13g2_a21oi_1 _07502_ (.A1(_00602_),
    .A2(net2774),
    .Y(_00274_),
    .B1(_01956_));
 sg13g2_nand2_1 _07503_ (.Y(_01957_),
    .A(net749),
    .B(net2774));
 sg13g2_nor3_2 _07504_ (.A(\core.work.alu.sval2[10] ),
    .B(net3542),
    .C(_01934_),
    .Y(_01958_));
 sg13g2_xnor2_1 _07505_ (.Y(_01959_),
    .A(_00118_),
    .B(_01958_));
 sg13g2_nand2_1 _07506_ (.Y(_01960_),
    .A(net3461),
    .B(\core.work.registers.genblk1[1].latch[11] ));
 sg13g2_nand2_1 _07507_ (.Y(_01961_),
    .A(\core.work.registers.genblk1[13].latch[11] ),
    .B(net3009));
 sg13g2_a22oi_1 _07508_ (.Y(_01962_),
    .B1(net2994),
    .B2(\core.work.registers.genblk1[6].latch[11] ),
    .A2(net3014),
    .A1(\core.work.registers.genblk1[2].latch[11] ));
 sg13g2_a21oi_1 _07509_ (.A1(\core.work.registers.genblk1[11].latch[11] ),
    .A2(net3185),
    .Y(_01963_),
    .B1(net3311));
 sg13g2_a22oi_1 _07510_ (.Y(_01964_),
    .B1(net3170),
    .B2(\core.work.registers.genblk1[12].latch[11] ),
    .A2(net3019),
    .A1(\core.work.registers.genblk1[14].latch[11] ));
 sg13g2_a22oi_1 _07511_ (.Y(_01965_),
    .B1(net3004),
    .B2(\core.work.registers.genblk1[5].latch[11] ),
    .A2(net3190),
    .A1(\core.work.registers.genblk1[3].latch[11] ));
 sg13g2_nand4_1 _07512_ (.B(_01963_),
    .C(_01964_),
    .A(_01962_),
    .Y(_01966_),
    .D(_01965_));
 sg13g2_a22oi_1 _07513_ (.Y(_01967_),
    .B1(net3180),
    .B2(\core.work.registers.genblk1[15].latch[11] ),
    .A2(net2999),
    .A1(\core.work.registers.genblk1[9].latch[11] ));
 sg13g2_a22oi_1 _07514_ (.Y(_01968_),
    .B1(net2983),
    .B2(\core.work.registers.genblk1[4].latch[11] ),
    .A2(net2989),
    .A1(\core.work.registers.genblk1[10].latch[11] ));
 sg13g2_a22oi_1 _07515_ (.Y(_01969_),
    .B1(net3174),
    .B2(\core.work.registers.genblk1[8].latch[11] ),
    .A2(net3023),
    .A1(\core.work.registers.genblk1[7].latch[11] ));
 sg13g2_nand4_1 _07516_ (.B(_01967_),
    .C(_01968_),
    .A(_01961_),
    .Y(_01970_),
    .D(_01969_));
 sg13g2_nor2_1 _07517_ (.A(_01966_),
    .B(_01970_),
    .Y(_01971_));
 sg13g2_a21oi_2 _07518_ (.B1(_01971_),
    .Y(_01972_),
    .A2(_01960_),
    .A1(net3312));
 sg13g2_a22oi_1 _07519_ (.Y(_01973_),
    .B1(_01972_),
    .B2(_01673_),
    .A2(_01882_),
    .A1(net3361));
 sg13g2_nor2_1 _07520_ (.A(net2909),
    .B(_01973_),
    .Y(_01974_));
 sg13g2_a221oi_1 _07521_ (.B2(net3305),
    .C1(_01974_),
    .B1(_01959_),
    .A1(net685),
    .Y(_01975_),
    .A2(net3166));
 sg13g2_o21ai_1 _07522_ (.B1(_01957_),
    .Y(_00275_),
    .A1(net2774),
    .A2(_01975_));
 sg13g2_nand2b_2 _07523_ (.Y(_01976_),
    .B(_01958_),
    .A_N(\core.work.alu.sval2[11] ));
 sg13g2_xnor2_1 _07524_ (.Y(_01977_),
    .A(_00722_),
    .B(_01976_));
 sg13g2_a21oi_2 _07525_ (.B1(_01685_),
    .Y(_01978_),
    .A2(net3035),
    .A1(net3442));
 sg13g2_nand2_1 _07526_ (.Y(_01979_),
    .A(net3462),
    .B(\core.work.registers.genblk1[1].latch[12] ));
 sg13g2_a21oi_1 _07527_ (.A1(\core.work.registers.genblk1[10].latch[12] ),
    .A2(net2992),
    .Y(_01980_),
    .B1(net3314));
 sg13g2_nand2_1 _07528_ (.Y(_01981_),
    .A(\core.work.registers.genblk1[5].latch[12] ),
    .B(net3007));
 sg13g2_a22oi_1 _07529_ (.Y(_01982_),
    .B1(net2987),
    .B2(\core.work.registers.genblk1[4].latch[12] ),
    .A2(net3012),
    .A1(\core.work.registers.genblk1[13].latch[12] ));
 sg13g2_a22oi_1 _07530_ (.Y(_01983_),
    .B1(net2999),
    .B2(\core.work.registers.genblk1[9].latch[12] ),
    .A2(net3019),
    .A1(\core.work.registers.genblk1[14].latch[12] ));
 sg13g2_a22oi_1 _07531_ (.Y(_01984_),
    .B1(net3193),
    .B2(\core.work.registers.genblk1[3].latch[12] ),
    .A2(net3014),
    .A1(\core.work.registers.genblk1[2].latch[12] ));
 sg13g2_a22oi_1 _07532_ (.Y(_01985_),
    .B1(net3175),
    .B2(\core.work.registers.genblk1[8].latch[12] ),
    .A2(net3024),
    .A1(\core.work.registers.genblk1[7].latch[12] ));
 sg13g2_a22oi_1 _07533_ (.Y(_01986_),
    .B1(net2994),
    .B2(\core.work.registers.genblk1[6].latch[12] ),
    .A2(net3185),
    .A1(\core.work.registers.genblk1[11].latch[12] ));
 sg13g2_nand4_1 _07534_ (.B(_01984_),
    .C(_01985_),
    .A(_01980_),
    .Y(_01987_),
    .D(_01986_));
 sg13g2_a22oi_1 _07535_ (.Y(_01988_),
    .B1(net3170),
    .B2(\core.work.registers.genblk1[12].latch[12] ),
    .A2(net3180),
    .A1(\core.work.registers.genblk1[15].latch[12] ));
 sg13g2_nand4_1 _07536_ (.B(_01982_),
    .C(_01983_),
    .A(_01981_),
    .Y(_01989_),
    .D(_01988_));
 sg13g2_nor2_1 _07537_ (.A(_01987_),
    .B(_01989_),
    .Y(_01990_));
 sg13g2_a21oi_2 _07538_ (.B1(_01990_),
    .Y(_01991_),
    .A2(_01979_),
    .A1(net3313));
 sg13g2_o21ai_1 _07539_ (.B1(net2895),
    .Y(_01992_),
    .A1(net3034),
    .A2(_01991_));
 sg13g2_nand2_1 _07540_ (.Y(_01993_),
    .A(net3480),
    .B(net3482));
 sg13g2_a21o_1 _07541_ (.A2(_01993_),
    .A1(net3484),
    .B1(net3442),
    .X(_01994_));
 sg13g2_o21ai_1 _07542_ (.B1(net3031),
    .Y(_01995_),
    .A1(net3492),
    .A2(_01994_));
 sg13g2_a21oi_1 _07543_ (.A1(net3490),
    .A2(_01991_),
    .Y(_01996_),
    .B1(net2892));
 sg13g2_nand2b_1 _07544_ (.Y(_01997_),
    .B(net3332),
    .A_N(_00120_));
 sg13g2_a221oi_1 _07545_ (.B2(net2909),
    .C1(_01996_),
    .B1(_01997_),
    .A1(net3196),
    .Y(_01998_),
    .A2(_01992_));
 sg13g2_a221oi_1 _07546_ (.B2(net3304),
    .C1(_01998_),
    .B1(_01977_),
    .A1(\core.f2e_addr[12] ),
    .Y(_01999_),
    .A2(net3165));
 sg13g2_nand2_1 _07547_ (.Y(_02000_),
    .A(net3541),
    .B(net2770));
 sg13g2_o21ai_1 _07548_ (.B1(_02000_),
    .Y(_00276_),
    .A1(net2771),
    .A2(_01999_));
 sg13g2_nor2_1 _07549_ (.A(net3541),
    .B(_01976_),
    .Y(_02001_));
 sg13g2_xnor2_1 _07550_ (.Y(_02002_),
    .A(_00121_),
    .B(_02001_));
 sg13g2_nand2_1 _07551_ (.Y(_02003_),
    .A(net3462),
    .B(\core.work.registers.genblk1[1].latch[13] ));
 sg13g2_nand2_1 _07552_ (.Y(_02004_),
    .A(\core.work.registers.genblk1[9].latch[13] ),
    .B(net2999));
 sg13g2_a22oi_1 _07553_ (.Y(_02005_),
    .B1(net2997),
    .B2(\core.work.registers.genblk1[6].latch[13] ),
    .A2(net3024),
    .A1(\core.work.registers.genblk1[7].latch[13] ));
 sg13g2_a21oi_1 _07554_ (.A1(\core.work.registers.genblk1[12].latch[13] ),
    .A2(net3170),
    .Y(_02006_),
    .B1(net3313));
 sg13g2_a22oi_1 _07555_ (.Y(_02007_),
    .B1(net3014),
    .B2(\core.work.registers.genblk1[2].latch[13] ),
    .A2(net3019),
    .A1(\core.work.registers.genblk1[14].latch[13] ));
 sg13g2_a22oi_1 _07556_ (.Y(_02008_),
    .B1(net2989),
    .B2(\core.work.registers.genblk1[10].latch[13] ),
    .A2(net3004),
    .A1(\core.work.registers.genblk1[5].latch[13] ));
 sg13g2_a22oi_1 _07557_ (.Y(_02009_),
    .B1(net3175),
    .B2(\core.work.registers.genblk1[8].latch[13] ),
    .A2(net3180),
    .A1(\core.work.registers.genblk1[15].latch[13] ));
 sg13g2_nand4_1 _07558_ (.B(_02007_),
    .C(_02008_),
    .A(_02006_),
    .Y(_02010_),
    .D(_02009_));
 sg13g2_a22oi_1 _07559_ (.Y(_02011_),
    .B1(net2984),
    .B2(\core.work.registers.genblk1[4].latch[13] ),
    .A2(net3009),
    .A1(\core.work.registers.genblk1[13].latch[13] ));
 sg13g2_a22oi_1 _07560_ (.Y(_02012_),
    .B1(net3185),
    .B2(\core.work.registers.genblk1[11].latch[13] ),
    .A2(net3190),
    .A1(\core.work.registers.genblk1[3].latch[13] ));
 sg13g2_nand4_1 _07561_ (.B(_02005_),
    .C(_02011_),
    .A(_02004_),
    .Y(_02013_),
    .D(_02012_));
 sg13g2_nor2_2 _07562_ (.A(_02010_),
    .B(_02013_),
    .Y(_02014_));
 sg13g2_a21oi_2 _07563_ (.B1(_02014_),
    .Y(_02015_),
    .A2(_02003_),
    .A1(net3313));
 sg13g2_o21ai_1 _07564_ (.B1(net2895),
    .Y(_02016_),
    .A1(net3034),
    .A2(_02015_));
 sg13g2_a21oi_1 _07565_ (.A1(net3490),
    .A2(_02015_),
    .Y(_02017_),
    .B1(net2892));
 sg13g2_nand2b_1 _07566_ (.Y(_02018_),
    .B(net3332),
    .A_N(_00122_));
 sg13g2_a221oi_1 _07567_ (.B2(net2909),
    .C1(_02017_),
    .B1(_02018_),
    .A1(net3196),
    .Y(_02019_),
    .A2(_02016_));
 sg13g2_a221oi_1 _07568_ (.B2(net3306),
    .C1(_02019_),
    .B1(_02002_),
    .A1(\core.f2e_addr[13] ),
    .Y(_02020_),
    .A2(net3165));
 sg13g2_nand2_1 _07569_ (.Y(_02021_),
    .A(net740),
    .B(net2774));
 sg13g2_o21ai_1 _07570_ (.B1(_02021_),
    .Y(_00277_),
    .A1(net2774),
    .A2(_02020_));
 sg13g2_nor3_2 _07571_ (.A(\core.work.alu.sval2[13] ),
    .B(net3541),
    .C(_01976_),
    .Y(_02022_));
 sg13g2_xnor2_1 _07572_ (.Y(_02023_),
    .A(net896),
    .B(_02022_));
 sg13g2_nand2_1 _07573_ (.Y(_02024_),
    .A(net3463),
    .B(\core.work.registers.genblk1[1].latch[14] ));
 sg13g2_nand2_1 _07574_ (.Y(_02025_),
    .A(\core.work.registers.genblk1[5].latch[14] ),
    .B(net3007));
 sg13g2_a22oi_1 _07575_ (.Y(_02026_),
    .B1(net3002),
    .B2(\core.work.registers.genblk1[9].latch[14] ),
    .A2(net3027),
    .A1(\core.work.registers.genblk1[7].latch[14] ));
 sg13g2_a22oi_1 _07576_ (.Y(_02027_),
    .B1(net3178),
    .B2(\core.work.registers.genblk1[8].latch[14] ),
    .A2(net3188),
    .A1(\core.work.registers.genblk1[11].latch[14] ));
 sg13g2_a22oi_1 _07577_ (.Y(_02028_),
    .B1(net2992),
    .B2(\core.work.registers.genblk1[10].latch[14] ),
    .A2(net3183),
    .A1(\core.work.registers.genblk1[15].latch[14] ));
 sg13g2_a21oi_1 _07578_ (.A1(\core.work.registers.genblk1[4].latch[14] ),
    .A2(net2987),
    .Y(_02029_),
    .B1(net3313));
 sg13g2_a22oi_1 _07579_ (.Y(_02030_),
    .B1(net2997),
    .B2(\core.work.registers.genblk1[6].latch[14] ),
    .A2(net3022),
    .A1(\core.work.registers.genblk1[14].latch[14] ));
 sg13g2_a22oi_1 _07580_ (.Y(_02031_),
    .B1(net3173),
    .B2(\core.work.registers.genblk1[12].latch[14] ),
    .A2(net3193),
    .A1(\core.work.registers.genblk1[3].latch[14] ));
 sg13g2_nand4_1 _07581_ (.B(_02029_),
    .C(_02030_),
    .A(_02028_),
    .Y(_02032_),
    .D(_02031_));
 sg13g2_a22oi_1 _07582_ (.Y(_02033_),
    .B1(net3012),
    .B2(\core.work.registers.genblk1[13].latch[14] ),
    .A2(net3017),
    .A1(\core.work.registers.genblk1[2].latch[14] ));
 sg13g2_nand4_1 _07583_ (.B(_02026_),
    .C(_02027_),
    .A(_02025_),
    .Y(_02034_),
    .D(_02033_));
 sg13g2_nor2_1 _07584_ (.A(_02032_),
    .B(_02034_),
    .Y(_02035_));
 sg13g2_a21oi_2 _07585_ (.B1(_02035_),
    .Y(_02036_),
    .A2(_02024_),
    .A1(net3314));
 sg13g2_o21ai_1 _07586_ (.B1(net2895),
    .Y(_02037_),
    .A1(net3032),
    .A2(_02036_));
 sg13g2_a21oi_1 _07587_ (.A1(net3490),
    .A2(_02036_),
    .Y(_02038_),
    .B1(net2892));
 sg13g2_nand2b_1 _07588_ (.Y(_02039_),
    .B(net3331),
    .A_N(_00124_));
 sg13g2_a221oi_1 _07589_ (.B2(net2909),
    .C1(_02038_),
    .B1(_02039_),
    .A1(net3194),
    .Y(_02040_),
    .A2(_02037_));
 sg13g2_a221oi_1 _07590_ (.B2(net3303),
    .C1(_02040_),
    .B1(_02023_),
    .A1(\core.f2e_addr[14] ),
    .Y(_02041_),
    .A2(net3165));
 sg13g2_nand2_1 _07591_ (.Y(_02042_),
    .A(net776),
    .B(net2770));
 sg13g2_o21ai_1 _07592_ (.B1(_02042_),
    .Y(_00278_),
    .A1(net2771),
    .A2(_02041_));
 sg13g2_nand2b_2 _07593_ (.Y(_02043_),
    .B(_02022_),
    .A_N(\core.work.alu.sval2[14] ));
 sg13g2_xor2_1 _07594_ (.B(_02043_),
    .A(_00125_),
    .X(_02044_));
 sg13g2_nand2_1 _07595_ (.Y(_02045_),
    .A(net3461),
    .B(\core.work.registers.genblk1[1].latch[15] ));
 sg13g2_nand2_1 _07596_ (.Y(_02046_),
    .A(\core.work.registers.genblk1[14].latch[15] ),
    .B(net3018));
 sg13g2_a22oi_1 _07597_ (.Y(_02047_),
    .B1(net2984),
    .B2(\core.work.registers.genblk1[4].latch[15] ),
    .A2(net3189),
    .A1(\core.work.registers.genblk1[3].latch[15] ));
 sg13g2_a21oi_1 _07598_ (.A1(\core.work.registers.genblk1[10].latch[15] ),
    .A2(net2988),
    .Y(_02048_),
    .B1(net3312));
 sg13g2_a22oi_1 _07599_ (.Y(_02049_),
    .B1(net2993),
    .B2(\core.work.registers.genblk1[6].latch[15] ),
    .A2(net3174),
    .A1(\core.work.registers.genblk1[8].latch[15] ));
 sg13g2_a22oi_1 _07600_ (.Y(_02050_),
    .B1(net3179),
    .B2(\core.work.registers.genblk1[15].latch[15] ),
    .A2(net3184),
    .A1(\core.work.registers.genblk1[11].latch[15] ));
 sg13g2_nand4_1 _07601_ (.B(_02048_),
    .C(_02049_),
    .A(_02047_),
    .Y(_02051_),
    .D(_02050_));
 sg13g2_a22oi_1 _07602_ (.Y(_02052_),
    .B1(net3169),
    .B2(\core.work.registers.genblk1[12].latch[15] ),
    .A2(net2998),
    .A1(\core.work.registers.genblk1[9].latch[15] ));
 sg13g2_a22oi_1 _07603_ (.Y(_02053_),
    .B1(net3008),
    .B2(\core.work.registers.genblk1[13].latch[15] ),
    .A2(net3013),
    .A1(\core.work.registers.genblk1[2].latch[15] ));
 sg13g2_a22oi_1 _07604_ (.Y(_02054_),
    .B1(net3003),
    .B2(\core.work.registers.genblk1[5].latch[15] ),
    .A2(net3023),
    .A1(\core.work.registers.genblk1[7].latch[15] ));
 sg13g2_nand4_1 _07605_ (.B(_02052_),
    .C(_02053_),
    .A(_02046_),
    .Y(_02055_),
    .D(_02054_));
 sg13g2_nor2_2 _07606_ (.A(_02051_),
    .B(_02055_),
    .Y(_02056_));
 sg13g2_a21oi_2 _07607_ (.B1(_02056_),
    .Y(_02057_),
    .A2(_02045_),
    .A1(net3311));
 sg13g2_o21ai_1 _07608_ (.B1(net2895),
    .Y(_02058_),
    .A1(net3032),
    .A2(_02057_));
 sg13g2_a21oi_1 _07609_ (.A1(net3490),
    .A2(_02057_),
    .Y(_02059_),
    .B1(net2892));
 sg13g2_nand2b_1 _07610_ (.Y(_02060_),
    .B(net3331),
    .A_N(_00126_));
 sg13g2_a221oi_1 _07611_ (.B2(net2909),
    .C1(_02059_),
    .B1(_02060_),
    .A1(net3194),
    .Y(_02061_),
    .A2(_02058_));
 sg13g2_a221oi_1 _07612_ (.B2(net3303),
    .C1(_02061_),
    .B1(_02044_),
    .A1(\core.f2e_addr[15] ),
    .Y(_02062_),
    .A2(net3165));
 sg13g2_nand2_1 _07613_ (.Y(_02063_),
    .A(net772),
    .B(net2770));
 sg13g2_o21ai_1 _07614_ (.B1(_02063_),
    .Y(_00279_),
    .A1(net2770),
    .A2(_02062_));
 sg13g2_and2_1 _07615_ (.A(net3331),
    .B(_01705_),
    .X(_02064_));
 sg13g2_nand3_1 _07616_ (.B(net2908),
    .C(_02064_),
    .A(net3195),
    .Y(_02065_));
 sg13g2_o21ai_1 _07617_ (.B1(_02065_),
    .Y(_00280_),
    .A1(_00630_),
    .A2(net2787));
 sg13g2_nand2b_2 _07618_ (.Y(_02066_),
    .B(_00598_),
    .A_N(_02043_));
 sg13g2_nor2_2 _07619_ (.A(net784),
    .B(_02066_),
    .Y(_02067_));
 sg13g2_nand3_1 _07620_ (.B(_00627_),
    .C(_02067_),
    .A(_00625_),
    .Y(_02068_));
 sg13g2_inv_1 _07621_ (.Y(_02069_),
    .A(_02068_));
 sg13g2_nor4_2 _07622_ (.A(\core.work.alu.sval2[22] ),
    .B(\core.work.alu.sval2[21] ),
    .C(net3530),
    .Y(_02070_),
    .D(net3531));
 sg13g2_nand2_2 _07623_ (.Y(_02071_),
    .A(_02069_),
    .B(_02070_));
 sg13g2_nor4_2 _07624_ (.A(\core.work.alu.sval2[26] ),
    .B(net3536),
    .C(net3533),
    .Y(_02072_),
    .D(net3534));
 sg13g2_nand3_1 _07625_ (.B(_02070_),
    .C(_02072_),
    .A(_02069_),
    .Y(_02073_));
 sg13g2_nor2_1 _07626_ (.A(net3537),
    .B(_02073_),
    .Y(_02074_));
 sg13g2_nor3_2 _07627_ (.A(\core.work.alu.sval2[28] ),
    .B(net3537),
    .C(_02073_),
    .Y(_02075_));
 sg13g2_nor2_1 _07628_ (.A(net3297),
    .B(_02075_),
    .Y(_02076_));
 sg13g2_o21ai_1 _07629_ (.B1(net3540),
    .Y(_02077_),
    .A1(net2770),
    .A2(_02076_));
 sg13g2_nand2_1 _07630_ (.Y(_02078_),
    .A(net3463),
    .B(\core.work.registers.genblk1[1].latch[29] ));
 sg13g2_nand2_1 _07631_ (.Y(_02079_),
    .A(\core.work.registers.genblk1[4].latch[29] ),
    .B(net2983));
 sg13g2_a21oi_1 _07632_ (.A1(\core.work.registers.genblk1[6].latch[29] ),
    .A2(net2993),
    .Y(_02080_),
    .B1(net3310));
 sg13g2_a22oi_1 _07633_ (.Y(_02081_),
    .B1(net3003),
    .B2(\core.work.registers.genblk1[5].latch[29] ),
    .A2(net3013),
    .A1(\core.work.registers.genblk1[2].latch[29] ));
 sg13g2_a22oi_1 _07634_ (.Y(_02082_),
    .B1(net3184),
    .B2(\core.work.registers.genblk1[11].latch[29] ),
    .A2(net3023),
    .A1(\core.work.registers.genblk1[7].latch[29] ));
 sg13g2_a22oi_1 _07635_ (.Y(_02083_),
    .B1(net3179),
    .B2(\core.work.registers.genblk1[15].latch[29] ),
    .A2(net3018),
    .A1(\core.work.registers.genblk1[14].latch[29] ));
 sg13g2_nand4_1 _07636_ (.B(_02081_),
    .C(_02082_),
    .A(_02080_),
    .Y(_02084_),
    .D(_02083_));
 sg13g2_a22oi_1 _07637_ (.Y(_02085_),
    .B1(net3174),
    .B2(\core.work.registers.genblk1[8].latch[29] ),
    .A2(net2998),
    .A1(\core.work.registers.genblk1[9].latch[29] ));
 sg13g2_a22oi_1 _07638_ (.Y(_02086_),
    .B1(net3169),
    .B2(\core.work.registers.genblk1[12].latch[29] ),
    .A2(net2988),
    .A1(\core.work.registers.genblk1[10].latch[29] ));
 sg13g2_a22oi_1 _07639_ (.Y(_02087_),
    .B1(net3008),
    .B2(\core.work.registers.genblk1[13].latch[29] ),
    .A2(net3189),
    .A1(\core.work.registers.genblk1[3].latch[29] ));
 sg13g2_nand4_1 _07640_ (.B(_02085_),
    .C(_02086_),
    .A(_02079_),
    .Y(_02088_),
    .D(_02087_));
 sg13g2_nor2_2 _07641_ (.A(_02084_),
    .B(_02088_),
    .Y(_02089_));
 sg13g2_a21oi_2 _07642_ (.B1(_02089_),
    .Y(_02090_),
    .A2(_02078_),
    .A1(net3311));
 sg13g2_o21ai_1 _07643_ (.B1(net2894),
    .Y(_02091_),
    .A1(net3033),
    .A2(_02090_));
 sg13g2_a21oi_1 _07644_ (.A1(net3489),
    .A2(_02090_),
    .Y(_02092_),
    .B1(net2891));
 sg13g2_a221oi_1 _07645_ (.B2(net3195),
    .C1(_02092_),
    .B1(_02091_),
    .A1(_00049_),
    .Y(_02093_),
    .A2(net3028));
 sg13g2_nor2_1 _07646_ (.A(net3540),
    .B(net3297),
    .Y(_02094_));
 sg13g2_a22oi_1 _07647_ (.Y(_02095_),
    .B1(_02094_),
    .B2(_02075_),
    .A2(_02093_),
    .A1(net3332));
 sg13g2_o21ai_1 _07648_ (.B1(_02077_),
    .Y(_00281_),
    .A1(net2770),
    .A2(_02095_));
 sg13g2_nand3_1 _07649_ (.B(_00608_),
    .C(_02075_),
    .A(_00606_),
    .Y(_02096_));
 sg13g2_a21oi_1 _07650_ (.A1(net663),
    .A2(_02096_),
    .Y(_02097_),
    .B1(_01710_));
 sg13g2_o21ai_1 _07651_ (.B1(_02097_),
    .Y(_02098_),
    .A1(net663),
    .A2(_02096_));
 sg13g2_nand2_1 _07652_ (.Y(_02099_),
    .A(net3463),
    .B(\core.work.registers.genblk1[1].latch[31] ));
 sg13g2_nand2_1 _07653_ (.Y(_02100_),
    .A(\core.work.registers.genblk1[8].latch[31] ),
    .B(net3174));
 sg13g2_a21oi_1 _07654_ (.A1(\core.work.registers.genblk1[13].latch[31] ),
    .A2(net3008),
    .Y(_02101_),
    .B1(net3311));
 sg13g2_a22oi_1 _07655_ (.Y(_02102_),
    .B1(net2993),
    .B2(\core.work.registers.genblk1[6].latch[31] ),
    .A2(net3189),
    .A1(\core.work.registers.genblk1[3].latch[31] ));
 sg13g2_a22oi_1 _07656_ (.Y(_02103_),
    .B1(net2988),
    .B2(\core.work.registers.genblk1[10].latch[31] ),
    .A2(net2998),
    .A1(\core.work.registers.genblk1[9].latch[31] ));
 sg13g2_nand3_1 _07657_ (.B(_02102_),
    .C(_02103_),
    .A(_02101_),
    .Y(_02104_));
 sg13g2_a221oi_1 _07658_ (.B2(\core.work.registers.genblk1[12].latch[31] ),
    .C1(_02104_),
    .B1(net3169),
    .A1(\core.work.registers.genblk1[4].latch[31] ),
    .Y(_02105_),
    .A2(net2983));
 sg13g2_a22oi_1 _07659_ (.Y(_02106_),
    .B1(net3179),
    .B2(\core.work.registers.genblk1[15].latch[31] ),
    .A2(net3023),
    .A1(\core.work.registers.genblk1[7].latch[31] ));
 sg13g2_a22oi_1 _07660_ (.Y(_02107_),
    .B1(net3013),
    .B2(\core.work.registers.genblk1[2].latch[31] ),
    .A2(net3018),
    .A1(\core.work.registers.genblk1[14].latch[31] ));
 sg13g2_nand3_1 _07661_ (.B(_02106_),
    .C(_02107_),
    .A(_02100_),
    .Y(_02108_));
 sg13g2_a221oi_1 _07662_ (.B2(\core.work.registers.genblk1[5].latch[31] ),
    .C1(_02108_),
    .B1(net3003),
    .A1(\core.work.registers.genblk1[11].latch[31] ),
    .Y(_02109_),
    .A2(net3184));
 sg13g2_a22oi_1 _07663_ (.Y(_02110_),
    .B1(_02105_),
    .B2(_02109_),
    .A2(_02099_),
    .A1(net3311));
 sg13g2_o21ai_1 _07664_ (.B1(net2895),
    .Y(_02111_),
    .A1(net3034),
    .A2(_02110_));
 sg13g2_a21oi_1 _07665_ (.A1(net3490),
    .A2(_02110_),
    .Y(_02112_),
    .B1(net2892));
 sg13g2_a21oi_1 _07666_ (.A1(_01670_),
    .A2(_02111_),
    .Y(_02113_),
    .B1(_02112_));
 sg13g2_a21oi_1 _07667_ (.A1(net3331),
    .A2(_02113_),
    .Y(_02114_),
    .B1(net2771));
 sg13g2_a22oi_1 _07668_ (.Y(_00282_),
    .B1(net664),
    .B2(_02114_),
    .A2(net2771),
    .A1(_00604_));
 sg13g2_o21ai_1 _07669_ (.B1(net816),
    .Y(_02115_),
    .A1(\core.work.state[1] ),
    .A2(_01708_));
 sg13g2_nand2_1 _07670_ (.Y(_02116_),
    .A(net3464),
    .B(\core.work.registers.genblk1[1].latch[0] ));
 sg13g2_nand2_1 _07671_ (.Y(_02117_),
    .A(\core.work.registers.genblk1[13].latch[0] ),
    .B(net3010));
 sg13g2_a22oi_1 _07672_ (.Y(_02118_),
    .B1(net3186),
    .B2(\core.work.registers.genblk1[11].latch[0] ),
    .A2(net3192),
    .A1(\core.work.registers.genblk1[3].latch[0] ));
 sg13g2_a21oi_1 _07673_ (.A1(\core.work.registers.genblk1[12].latch[0] ),
    .A2(net3171),
    .Y(_02119_),
    .B1(net3318));
 sg13g2_a22oi_1 _07674_ (.Y(_02120_),
    .B1(net3176),
    .B2(\core.work.registers.genblk1[8].latch[0] ),
    .A2(net3006),
    .A1(\core.work.registers.genblk1[5].latch[0] ));
 sg13g2_a22oi_1 _07675_ (.Y(_02121_),
    .B1(net3016),
    .B2(\core.work.registers.genblk1[2].latch[0] ),
    .A2(net3021),
    .A1(\core.work.registers.genblk1[14].latch[0] ));
 sg13g2_nand4_1 _07676_ (.B(_02119_),
    .C(_02120_),
    .A(_02118_),
    .Y(_02122_),
    .D(_02121_));
 sg13g2_a22oi_1 _07677_ (.Y(_02123_),
    .B1(net3001),
    .B2(\core.work.registers.genblk1[9].latch[0] ),
    .A2(net3026),
    .A1(\core.work.registers.genblk1[7].latch[0] ));
 sg13g2_a22oi_1 _07678_ (.Y(_02124_),
    .B1(net2985),
    .B2(\core.work.registers.genblk1[4].latch[0] ),
    .A2(net2991),
    .A1(\core.work.registers.genblk1[10].latch[0] ));
 sg13g2_a22oi_1 _07679_ (.Y(_02125_),
    .B1(net2996),
    .B2(\core.work.registers.genblk1[6].latch[0] ),
    .A2(net3181),
    .A1(\core.work.registers.genblk1[15].latch[0] ));
 sg13g2_nand4_1 _07680_ (.B(_02123_),
    .C(_02124_),
    .A(_02117_),
    .Y(_02126_),
    .D(_02125_));
 sg13g2_nor2_1 _07681_ (.A(_02122_),
    .B(_02126_),
    .Y(_02127_));
 sg13g2_a21oi_2 _07682_ (.B1(_02127_),
    .Y(_02128_),
    .A2(_02116_),
    .A1(net3317));
 sg13g2_inv_1 _07683_ (.Y(_02129_),
    .A(_02128_));
 sg13g2_a21oi_1 _07684_ (.A1(net3493),
    .A2(_02129_),
    .Y(_02130_),
    .B1(net3330));
 sg13g2_mux2_1 _07685_ (.A0(net3460),
    .A1(_00154_),
    .S(_01665_),
    .X(_02131_));
 sg13g2_or2_1 _07686_ (.X(_02132_),
    .B(net3030),
    .A(_01685_));
 sg13g2_nor2_1 _07687_ (.A(_01685_),
    .B(net2910),
    .Y(_02133_));
 sg13g2_nand2b_2 _07688_ (.Y(_02134_),
    .B(_01686_),
    .A_N(net2909));
 sg13g2_a221oi_1 _07689_ (.B2(net2908),
    .C1(_02134_),
    .B1(_02131_),
    .A1(_01673_),
    .Y(_02135_),
    .A2(_02129_));
 sg13g2_a21oi_1 _07690_ (.A1(net3031),
    .A2(_02130_),
    .Y(_02136_),
    .B1(_02135_));
 sg13g2_a21oi_1 _07691_ (.A1(net3460),
    .A2(net2922),
    .Y(_02137_),
    .B1(_02136_));
 sg13g2_nand2_1 _07692_ (.Y(_02138_),
    .A(_01707_),
    .B(_02137_));
 sg13g2_nand2_2 _07693_ (.Y(_00283_),
    .A(net817),
    .B(_02138_));
 sg13g2_nand2_1 _07694_ (.Y(_02139_),
    .A(_00051_),
    .B(_02075_));
 sg13g2_a21oi_1 _07695_ (.A1(net679),
    .A2(_02139_),
    .Y(_02140_),
    .B1(net3297));
 sg13g2_o21ai_1 _07696_ (.B1(_02140_),
    .Y(_02141_),
    .A1(net679),
    .A2(_02139_));
 sg13g2_nand2_1 _07697_ (.Y(_02142_),
    .A(net3461),
    .B(\core.work.registers.genblk1[1].latch[30] ));
 sg13g2_nand2_1 _07698_ (.Y(_02143_),
    .A(\core.work.registers.genblk1[8].latch[30] ),
    .B(net3174));
 sg13g2_a21oi_1 _07699_ (.A1(\core.work.registers.genblk1[4].latch[30] ),
    .A2(net2983),
    .Y(_02144_),
    .B1(net3310));
 sg13g2_a22oi_1 _07700_ (.Y(_02145_),
    .B1(net3169),
    .B2(\core.work.registers.genblk1[12].latch[30] ),
    .A2(net3018),
    .A1(\core.work.registers.genblk1[14].latch[30] ));
 sg13g2_a22oi_1 _07701_ (.Y(_02146_),
    .B1(net2993),
    .B2(\core.work.registers.genblk1[6].latch[30] ),
    .A2(net3189),
    .A1(\core.work.registers.genblk1[3].latch[30] ));
 sg13g2_nand3_1 _07702_ (.B(_02145_),
    .C(_02146_),
    .A(_02144_),
    .Y(_02147_));
 sg13g2_a221oi_1 _07703_ (.B2(\core.work.registers.genblk1[10].latch[30] ),
    .C1(_02147_),
    .B1(net2988),
    .A1(\core.work.registers.genblk1[15].latch[30] ),
    .Y(_02148_),
    .A2(net3179));
 sg13g2_a22oi_1 _07704_ (.Y(_02149_),
    .B1(net2998),
    .B2(\core.work.registers.genblk1[9].latch[30] ),
    .A2(net3023),
    .A1(\core.work.registers.genblk1[7].latch[30] ));
 sg13g2_a22oi_1 _07705_ (.Y(_02150_),
    .B1(net3003),
    .B2(\core.work.registers.genblk1[5].latch[30] ),
    .A2(net3184),
    .A1(\core.work.registers.genblk1[11].latch[30] ));
 sg13g2_nand3_1 _07706_ (.B(_02149_),
    .C(_02150_),
    .A(_02143_),
    .Y(_02151_));
 sg13g2_a221oi_1 _07707_ (.B2(\core.work.registers.genblk1[13].latch[30] ),
    .C1(_02151_),
    .B1(net3008),
    .A1(\core.work.registers.genblk1[2].latch[30] ),
    .Y(_02152_),
    .A2(net3013));
 sg13g2_a22oi_1 _07708_ (.Y(_02153_),
    .B1(_02148_),
    .B2(_02152_),
    .A2(_02142_),
    .A1(net3310));
 sg13g2_o21ai_1 _07709_ (.B1(net2895),
    .Y(_02154_),
    .A1(net3033),
    .A2(_02153_));
 sg13g2_a21oi_1 _07710_ (.A1(_00052_),
    .A2(net3029),
    .Y(_02155_),
    .B1(net3329));
 sg13g2_a21oi_1 _07711_ (.A1(net3490),
    .A2(_02153_),
    .Y(_02156_),
    .B1(net2892));
 sg13g2_a21oi_1 _07712_ (.A1(net3194),
    .A2(_02154_),
    .Y(_02157_),
    .B1(_02156_));
 sg13g2_a21oi_1 _07713_ (.A1(_02155_),
    .A2(_02157_),
    .Y(_02158_),
    .B1(net2770));
 sg13g2_a22oi_1 _07714_ (.Y(_00284_),
    .B1(net680),
    .B2(_02158_),
    .A2(net2770),
    .A1(_00606_));
 sg13g2_xnor2_1 _07715_ (.Y(_02159_),
    .A(_00047_),
    .B(_02074_));
 sg13g2_nand2_1 _07716_ (.Y(_02160_),
    .A(net3461),
    .B(\core.work.registers.genblk1[1].latch[28] ));
 sg13g2_nand2_1 _07717_ (.Y(_02161_),
    .A(\core.work.registers.genblk1[6].latch[28] ),
    .B(net2993));
 sg13g2_a22oi_1 _07718_ (.Y(_02162_),
    .B1(net3179),
    .B2(\core.work.registers.genblk1[15].latch[28] ),
    .A2(net3023),
    .A1(\core.work.registers.genblk1[7].latch[28] ));
 sg13g2_a21oi_1 _07719_ (.A1(\core.work.registers.genblk1[12].latch[28] ),
    .A2(net3169),
    .Y(_02163_),
    .B1(net3310));
 sg13g2_a22oi_1 _07720_ (.Y(_02164_),
    .B1(net3013),
    .B2(\core.work.registers.genblk1[2].latch[28] ),
    .A2(net3018),
    .A1(\core.work.registers.genblk1[14].latch[28] ));
 sg13g2_a22oi_1 _07721_ (.Y(_02165_),
    .B1(net3184),
    .B2(\core.work.registers.genblk1[11].latch[28] ),
    .A2(net3189),
    .A1(\core.work.registers.genblk1[3].latch[28] ));
 sg13g2_nand4_1 _07722_ (.B(_02163_),
    .C(_02164_),
    .A(_02162_),
    .Y(_02166_),
    .D(_02165_));
 sg13g2_a22oi_1 _07723_ (.Y(_02167_),
    .B1(net2983),
    .B2(\core.work.registers.genblk1[4].latch[28] ),
    .A2(net2998),
    .A1(\core.work.registers.genblk1[9].latch[28] ));
 sg13g2_a22oi_1 _07724_ (.Y(_02168_),
    .B1(net3174),
    .B2(\core.work.registers.genblk1[8].latch[28] ),
    .A2(net3003),
    .A1(\core.work.registers.genblk1[5].latch[28] ));
 sg13g2_a22oi_1 _07725_ (.Y(_02169_),
    .B1(net2988),
    .B2(\core.work.registers.genblk1[10].latch[28] ),
    .A2(net3008),
    .A1(\core.work.registers.genblk1[13].latch[28] ));
 sg13g2_nand4_1 _07726_ (.B(_02167_),
    .C(_02168_),
    .A(_02161_),
    .Y(_02170_),
    .D(_02169_));
 sg13g2_nor2_2 _07727_ (.A(_02166_),
    .B(_02170_),
    .Y(_02171_));
 sg13g2_a21oi_2 _07728_ (.B1(_02171_),
    .Y(_02172_),
    .A2(_02160_),
    .A1(net3311));
 sg13g2_o21ai_1 _07729_ (.B1(net2894),
    .Y(_02173_),
    .A1(net3032),
    .A2(_02172_));
 sg13g2_a21oi_1 _07730_ (.A1(_00048_),
    .A2(net3028),
    .Y(_02174_),
    .B1(net3329));
 sg13g2_a21oi_1 _07731_ (.A1(net3489),
    .A2(_02172_),
    .Y(_02175_),
    .B1(net2891));
 sg13g2_a21oi_1 _07732_ (.A1(net3194),
    .A2(_02173_),
    .Y(_02176_),
    .B1(_02175_));
 sg13g2_a221oi_1 _07733_ (.B2(_02176_),
    .C1(net2769),
    .B1(_02174_),
    .A1(net3304),
    .Y(_02177_),
    .A2(_02159_));
 sg13g2_a21oi_1 _07734_ (.A1(_00610_),
    .A2(net2769),
    .Y(_00285_),
    .B1(_02177_));
 sg13g2_xor2_1 _07735_ (.B(_02073_),
    .A(net810),
    .X(_02178_));
 sg13g2_nand2_1 _07736_ (.Y(_02179_),
    .A(net3461),
    .B(\core.work.registers.genblk1[1].latch[27] ));
 sg13g2_a21oi_1 _07737_ (.A1(\core.work.registers.genblk1[12].latch[27] ),
    .A2(net3169),
    .Y(_02180_),
    .B1(net3310));
 sg13g2_nand2_1 _07738_ (.Y(_02181_),
    .A(\core.work.registers.genblk1[13].latch[27] ),
    .B(net3008));
 sg13g2_a22oi_1 _07739_ (.Y(_02182_),
    .B1(net3189),
    .B2(\core.work.registers.genblk1[3].latch[27] ),
    .A2(net3013),
    .A1(\core.work.registers.genblk1[2].latch[27] ));
 sg13g2_a22oi_1 _07740_ (.Y(_02183_),
    .B1(net2988),
    .B2(\core.work.registers.genblk1[10].latch[27] ),
    .A2(net3179),
    .A1(\core.work.registers.genblk1[15].latch[27] ));
 sg13g2_a22oi_1 _07741_ (.Y(_02184_),
    .B1(net2983),
    .B2(\core.work.registers.genblk1[4].latch[27] ),
    .A2(net3175),
    .A1(\core.work.registers.genblk1[8].latch[27] ));
 sg13g2_nand4_1 _07742_ (.B(_02182_),
    .C(_02183_),
    .A(_02180_),
    .Y(_02185_),
    .D(_02184_));
 sg13g2_a22oi_1 _07743_ (.Y(_02186_),
    .B1(net2998),
    .B2(\core.work.registers.genblk1[9].latch[27] ),
    .A2(net3024),
    .A1(\core.work.registers.genblk1[7].latch[27] ));
 sg13g2_a22oi_1 _07744_ (.Y(_02187_),
    .B1(net2993),
    .B2(\core.work.registers.genblk1[6].latch[27] ),
    .A2(net3018),
    .A1(\core.work.registers.genblk1[14].latch[27] ));
 sg13g2_a22oi_1 _07745_ (.Y(_02188_),
    .B1(net3003),
    .B2(\core.work.registers.genblk1[5].latch[27] ),
    .A2(net3184),
    .A1(\core.work.registers.genblk1[11].latch[27] ));
 sg13g2_nand4_1 _07746_ (.B(_02186_),
    .C(_02187_),
    .A(_02181_),
    .Y(_02189_),
    .D(_02188_));
 sg13g2_nor2_2 _07747_ (.A(_02185_),
    .B(_02189_),
    .Y(_02190_));
 sg13g2_a21oi_2 _07748_ (.B1(_02190_),
    .Y(_02191_),
    .A2(_02179_),
    .A1(net3311));
 sg13g2_o21ai_1 _07749_ (.B1(net2894),
    .Y(_02192_),
    .A1(net3032),
    .A2(_02191_));
 sg13g2_a21oi_1 _07750_ (.A1(_00046_),
    .A2(net3028),
    .Y(_02193_),
    .B1(net3330));
 sg13g2_a21oi_1 _07751_ (.A1(net3489),
    .A2(_02191_),
    .Y(_02194_),
    .B1(net2891));
 sg13g2_a21oi_1 _07752_ (.A1(net3194),
    .A2(_02192_),
    .Y(_02195_),
    .B1(_02194_));
 sg13g2_a22oi_1 _07753_ (.Y(_02196_),
    .B1(_02193_),
    .B2(_02195_),
    .A2(_02178_),
    .A1(net3304));
 sg13g2_nand2_1 _07754_ (.Y(_02197_),
    .A(net3537),
    .B(net2772));
 sg13g2_o21ai_1 _07755_ (.B1(_02197_),
    .Y(_00286_),
    .A1(net2769),
    .A2(net811));
 sg13g2_nor2_1 _07756_ (.A(net3534),
    .B(_02071_),
    .Y(_02198_));
 sg13g2_nor3_1 _07757_ (.A(\core.work.alu.sval2[24] ),
    .B(net3534),
    .C(_02071_),
    .Y(_02199_));
 sg13g2_nand2_1 _07758_ (.Y(_02200_),
    .A(_00043_),
    .B(_02199_));
 sg13g2_xor2_1 _07759_ (.B(_02200_),
    .A(_00042_),
    .X(_02201_));
 sg13g2_nand2_1 _07760_ (.Y(_02202_),
    .A(net3461),
    .B(\core.work.registers.genblk1[1].latch[26] ));
 sg13g2_nand2_1 _07761_ (.Y(_02203_),
    .A(\core.work.registers.genblk1[6].latch[26] ),
    .B(net2993));
 sg13g2_a22oi_1 _07762_ (.Y(_02204_),
    .B1(net3189),
    .B2(\core.work.registers.genblk1[3].latch[26] ),
    .A2(net3013),
    .A1(\core.work.registers.genblk1[2].latch[26] ));
 sg13g2_a21oi_1 _07763_ (.A1(\core.work.registers.genblk1[7].latch[26] ),
    .A2(net3023),
    .Y(_02205_),
    .B1(net3310));
 sg13g2_a22oi_1 _07764_ (.Y(_02206_),
    .B1(net3179),
    .B2(\core.work.registers.genblk1[15].latch[26] ),
    .A2(net3184),
    .A1(\core.work.registers.genblk1[11].latch[26] ));
 sg13g2_a22oi_1 _07765_ (.Y(_02207_),
    .B1(net2983),
    .B2(\core.work.registers.genblk1[4].latch[26] ),
    .A2(net3018),
    .A1(\core.work.registers.genblk1[14].latch[26] ));
 sg13g2_nand4_1 _07766_ (.B(_02205_),
    .C(_02206_),
    .A(_02204_),
    .Y(_02208_),
    .D(_02207_));
 sg13g2_a22oi_1 _07767_ (.Y(_02209_),
    .B1(net2988),
    .B2(\core.work.registers.genblk1[10].latch[26] ),
    .A2(net3008),
    .A1(\core.work.registers.genblk1[13].latch[26] ));
 sg13g2_a22oi_1 _07768_ (.Y(_02210_),
    .B1(net3169),
    .B2(\core.work.registers.genblk1[12].latch[26] ),
    .A2(net3003),
    .A1(\core.work.registers.genblk1[5].latch[26] ));
 sg13g2_a22oi_1 _07769_ (.Y(_02211_),
    .B1(net3174),
    .B2(\core.work.registers.genblk1[8].latch[26] ),
    .A2(net2998),
    .A1(\core.work.registers.genblk1[9].latch[26] ));
 sg13g2_nand4_1 _07770_ (.B(_02209_),
    .C(_02210_),
    .A(_02203_),
    .Y(_02212_),
    .D(_02211_));
 sg13g2_nor2_2 _07771_ (.A(_02208_),
    .B(_02212_),
    .Y(_02213_));
 sg13g2_a21oi_2 _07772_ (.B1(_02213_),
    .Y(_02214_),
    .A2(_02202_),
    .A1(net3311));
 sg13g2_o21ai_1 _07773_ (.B1(net2895),
    .Y(_02215_),
    .A1(net3033),
    .A2(_02214_));
 sg13g2_nand2_1 _07774_ (.Y(_02216_),
    .A(net3195),
    .B(_02215_));
 sg13g2_a21oi_1 _07775_ (.A1(net3491),
    .A2(_02214_),
    .Y(_02217_),
    .B1(net2892));
 sg13g2_a21oi_1 _07776_ (.A1(_00044_),
    .A2(net3028),
    .Y(_02218_),
    .B1(net3330));
 sg13g2_nor2b_1 _07777_ (.A(_02217_),
    .B_N(_02218_),
    .Y(_02219_));
 sg13g2_a221oi_1 _07778_ (.B2(_02219_),
    .C1(net2769),
    .B1(_02216_),
    .A1(net3304),
    .Y(_02220_),
    .A2(_02201_));
 sg13g2_a21oi_1 _07779_ (.A1(_00612_),
    .A2(net2769),
    .Y(_00287_),
    .B1(_02220_));
 sg13g2_nor2_1 _07780_ (.A(net3298),
    .B(_02199_),
    .Y(_02221_));
 sg13g2_o21ai_1 _07781_ (.B1(net3536),
    .Y(_02222_),
    .A1(net2773),
    .A2(_02221_));
 sg13g2_nand2_1 _07782_ (.Y(_02223_),
    .A(net3462),
    .B(\core.work.registers.genblk1[1].latch[25] ));
 sg13g2_nand2_1 _07783_ (.Y(_02224_),
    .A(\core.work.registers.genblk1[5].latch[25] ),
    .B(net3004));
 sg13g2_a22oi_1 _07784_ (.Y(_02225_),
    .B1(net2989),
    .B2(\core.work.registers.genblk1[10].latch[25] ),
    .A2(net3014),
    .A1(\core.work.registers.genblk1[2].latch[25] ));
 sg13g2_a22oi_1 _07785_ (.Y(_02226_),
    .B1(net2984),
    .B2(\core.work.registers.genblk1[4].latch[25] ),
    .A2(net3190),
    .A1(\core.work.registers.genblk1[3].latch[25] ));
 sg13g2_a21oi_1 _07786_ (.A1(\core.work.registers.genblk1[7].latch[25] ),
    .A2(net3024),
    .Y(_02227_),
    .B1(net3313));
 sg13g2_a22oi_1 _07787_ (.Y(_02228_),
    .B1(net3185),
    .B2(\core.work.registers.genblk1[11].latch[25] ),
    .A2(net3019),
    .A1(\core.work.registers.genblk1[14].latch[25] ));
 sg13g2_nand4_1 _07788_ (.B(_02226_),
    .C(_02227_),
    .A(_02225_),
    .Y(_02229_),
    .D(_02228_));
 sg13g2_a22oi_1 _07789_ (.Y(_02230_),
    .B1(net2994),
    .B2(\core.work.registers.genblk1[6].latch[25] ),
    .A2(net3009),
    .A1(\core.work.registers.genblk1[13].latch[25] ));
 sg13g2_a22oi_1 _07790_ (.Y(_02231_),
    .B1(net3173),
    .B2(\core.work.registers.genblk1[12].latch[25] ),
    .A2(net3180),
    .A1(\core.work.registers.genblk1[15].latch[25] ));
 sg13g2_a22oi_1 _07791_ (.Y(_02232_),
    .B1(net3178),
    .B2(\core.work.registers.genblk1[8].latch[25] ),
    .A2(net3002),
    .A1(\core.work.registers.genblk1[9].latch[25] ));
 sg13g2_nand4_1 _07792_ (.B(_02230_),
    .C(_02231_),
    .A(_02224_),
    .Y(_02233_),
    .D(_02232_));
 sg13g2_nor2_1 _07793_ (.A(_02229_),
    .B(_02233_),
    .Y(_02234_));
 sg13g2_a21oi_2 _07794_ (.B1(_02234_),
    .Y(_02235_),
    .A2(_02223_),
    .A1(net3313));
 sg13g2_o21ai_1 _07795_ (.B1(net2894),
    .Y(_02236_),
    .A1(net3032),
    .A2(_02235_));
 sg13g2_a21oi_1 _07796_ (.A1(net3489),
    .A2(_02235_),
    .Y(_02237_),
    .B1(net2891));
 sg13g2_nand2b_1 _07797_ (.Y(_02238_),
    .B(net3331),
    .A_N(_00041_));
 sg13g2_a221oi_1 _07798_ (.B2(net2909),
    .C1(_02237_),
    .B1(_02238_),
    .A1(net3194),
    .Y(_02239_),
    .A2(_02236_));
 sg13g2_nor3_1 _07799_ (.A(net3536),
    .B(net3533),
    .C(net3297),
    .Y(_02240_));
 sg13g2_a21oi_1 _07800_ (.A1(_02198_),
    .A2(_02240_),
    .Y(_02241_),
    .B1(_02239_));
 sg13g2_o21ai_1 _07801_ (.B1(net839),
    .Y(_00288_),
    .A1(net2773),
    .A2(_02241_));
 sg13g2_xnor2_1 _07802_ (.Y(_02242_),
    .A(_00635_),
    .B(_02066_));
 sg13g2_nand2_1 _07803_ (.Y(_02243_),
    .A(net3467),
    .B(\core.work.registers.genblk1[1].latch[16] ));
 sg13g2_nand2_1 _07804_ (.Y(_02244_),
    .A(\core.work.registers.genblk1[7].latch[16] ),
    .B(net3025));
 sg13g2_a22oi_1 _07805_ (.Y(_02245_),
    .B1(net2990),
    .B2(\core.work.registers.genblk1[10].latch[16] ),
    .A2(net3181),
    .A1(\core.work.registers.genblk1[15].latch[16] ));
 sg13g2_a21oi_1 _07806_ (.A1(\core.work.registers.genblk1[14].latch[16] ),
    .A2(net3020),
    .Y(_02246_),
    .B1(net3315));
 sg13g2_a22oi_1 _07807_ (.Y(_02247_),
    .B1(net3186),
    .B2(\core.work.registers.genblk1[11].latch[16] ),
    .A2(net3191),
    .A1(\core.work.registers.genblk1[3].latch[16] ));
 sg13g2_a22oi_1 _07808_ (.Y(_02248_),
    .B1(net2985),
    .B2(\core.work.registers.genblk1[4].latch[16] ),
    .A2(net3177),
    .A1(\core.work.registers.genblk1[8].latch[16] ));
 sg13g2_nand4_1 _07809_ (.B(_02246_),
    .C(_02247_),
    .A(_02245_),
    .Y(_02249_),
    .D(_02248_));
 sg13g2_a22oi_1 _07810_ (.Y(_02250_),
    .B1(net2995),
    .B2(\core.work.registers.genblk1[6].latch[16] ),
    .A2(net3000),
    .A1(\core.work.registers.genblk1[9].latch[16] ));
 sg13g2_a22oi_1 _07811_ (.Y(_02251_),
    .B1(net3171),
    .B2(\core.work.registers.genblk1[12].latch[16] ),
    .A2(net3005),
    .A1(\core.work.registers.genblk1[5].latch[16] ));
 sg13g2_a22oi_1 _07812_ (.Y(_02252_),
    .B1(net3010),
    .B2(\core.work.registers.genblk1[13].latch[16] ),
    .A2(net3015),
    .A1(\core.work.registers.genblk1[2].latch[16] ));
 sg13g2_nand4_1 _07813_ (.B(_02250_),
    .C(_02251_),
    .A(_02244_),
    .Y(_02253_),
    .D(_02252_));
 sg13g2_nor2_2 _07814_ (.A(_02249_),
    .B(_02253_),
    .Y(_02254_));
 sg13g2_a21oi_2 _07815_ (.B1(_02254_),
    .Y(_02255_),
    .A2(_02243_),
    .A1(net3315));
 sg13g2_o21ai_1 _07816_ (.B1(net2896),
    .Y(_02256_),
    .A1(net3036),
    .A2(_02255_));
 sg13g2_a21oi_1 _07817_ (.A1(_00023_),
    .A2(net3030),
    .Y(_02257_),
    .B1(net3330));
 sg13g2_a21oi_1 _07818_ (.A1(net3494),
    .A2(_02255_),
    .Y(_02258_),
    .B1(net2893));
 sg13g2_a21oi_1 _07819_ (.A1(net3196),
    .A2(_02256_),
    .Y(_02259_),
    .B1(_02258_));
 sg13g2_a22oi_1 _07820_ (.Y(_02260_),
    .B1(_02257_),
    .B2(_02259_),
    .A2(_02242_),
    .A1(net3309));
 sg13g2_nand2_1 _07821_ (.Y(_02261_),
    .A(net3535),
    .B(net2776));
 sg13g2_o21ai_1 _07822_ (.B1(_02261_),
    .Y(_00289_),
    .A1(net2776),
    .A2(_02260_));
 sg13g2_nor2_1 _07823_ (.A(net3531),
    .B(_02068_),
    .Y(_02262_));
 sg13g2_nor3_1 _07824_ (.A(net3530),
    .B(net3531),
    .C(_02068_),
    .Y(_02263_));
 sg13g2_nor2_1 _07825_ (.A(net3299),
    .B(_02263_),
    .Y(_02264_));
 sg13g2_o21ai_1 _07826_ (.B1(net778),
    .Y(_02265_),
    .A1(net2775),
    .A2(_02264_));
 sg13g2_nand2_1 _07827_ (.Y(_02266_),
    .A(net3462),
    .B(\core.work.registers.genblk1[1].latch[21] ));
 sg13g2_a21oi_1 _07828_ (.A1(\core.work.registers.genblk1[9].latch[21] ),
    .A2(net2999),
    .Y(_02267_),
    .B1(net3313));
 sg13g2_nand2_1 _07829_ (.Y(_02268_),
    .A(\core.work.registers.genblk1[15].latch[21] ),
    .B(net3180));
 sg13g2_a22oi_1 _07830_ (.Y(_02269_),
    .B1(net3004),
    .B2(\core.work.registers.genblk1[5].latch[21] ),
    .A2(net3014),
    .A1(\core.work.registers.genblk1[2].latch[21] ));
 sg13g2_a22oi_1 _07831_ (.Y(_02270_),
    .B1(net2989),
    .B2(\core.work.registers.genblk1[10].latch[21] ),
    .A2(net3019),
    .A1(\core.work.registers.genblk1[14].latch[21] ));
 sg13g2_a22oi_1 _07832_ (.Y(_02271_),
    .B1(net3170),
    .B2(\core.work.registers.genblk1[12].latch[21] ),
    .A2(net3185),
    .A1(\core.work.registers.genblk1[11].latch[21] ));
 sg13g2_a22oi_1 _07833_ (.Y(_02272_),
    .B1(net3190),
    .B2(\core.work.registers.genblk1[3].latch[21] ),
    .A2(net3024),
    .A1(\core.work.registers.genblk1[7].latch[21] ));
 sg13g2_nand4_1 _07834_ (.B(_02270_),
    .C(_02271_),
    .A(_02267_),
    .Y(_02273_),
    .D(_02272_));
 sg13g2_a22oi_1 _07835_ (.Y(_02274_),
    .B1(net2984),
    .B2(\core.work.registers.genblk1[4].latch[21] ),
    .A2(net3175),
    .A1(\core.work.registers.genblk1[8].latch[21] ));
 sg13g2_a22oi_1 _07836_ (.Y(_02275_),
    .B1(net2994),
    .B2(\core.work.registers.genblk1[6].latch[21] ),
    .A2(net3009),
    .A1(\core.work.registers.genblk1[13].latch[21] ));
 sg13g2_nand4_1 _07837_ (.B(_02269_),
    .C(_02274_),
    .A(_02268_),
    .Y(_02276_),
    .D(_02275_));
 sg13g2_nor2_2 _07838_ (.A(_02273_),
    .B(_02276_),
    .Y(_02277_));
 sg13g2_a21oi_2 _07839_ (.B1(_02277_),
    .Y(_02278_),
    .A2(_02266_),
    .A1(net3314));
 sg13g2_o21ai_1 _07840_ (.B1(net2896),
    .Y(_02279_),
    .A1(net3036),
    .A2(_02278_));
 sg13g2_a21oi_1 _07841_ (.A1(net3494),
    .A2(_02278_),
    .Y(_02280_),
    .B1(net2893));
 sg13g2_a221oi_1 _07842_ (.B2(net3196),
    .C1(_02280_),
    .B1(_02279_),
    .A1(_00033_),
    .Y(_02281_),
    .A2(net3030));
 sg13g2_nor4_1 _07843_ (.A(\core.work.alu.sval2[21] ),
    .B(net3530),
    .C(net3531),
    .D(net3299),
    .Y(_02282_));
 sg13g2_a22oi_1 _07844_ (.Y(_02283_),
    .B1(_02282_),
    .B2(_02069_),
    .A2(_02281_),
    .A1(_01645_));
 sg13g2_o21ai_1 _07845_ (.B1(_02265_),
    .Y(_00290_),
    .A1(net2775),
    .A2(_02283_));
 sg13g2_nand2_1 _07846_ (.Y(_02284_),
    .A(_00035_),
    .B(_02263_));
 sg13g2_a21oi_1 _07847_ (.A1(net682),
    .A2(_02284_),
    .Y(_02285_),
    .B1(net3299));
 sg13g2_o21ai_1 _07848_ (.B1(_02285_),
    .Y(_02286_),
    .A1(net682),
    .A2(_02284_));
 sg13g2_nand2_1 _07849_ (.Y(_02287_),
    .A(net3461),
    .B(\core.work.registers.genblk1[1].latch[22] ));
 sg13g2_nand2_1 _07850_ (.Y(_02288_),
    .A(\core.work.registers.genblk1[14].latch[22] ),
    .B(net3019));
 sg13g2_a22oi_1 _07851_ (.Y(_02289_),
    .B1(net2989),
    .B2(\core.work.registers.genblk1[10].latch[22] ),
    .A2(net3014),
    .A1(\core.work.registers.genblk1[2].latch[22] ));
 sg13g2_a22oi_1 _07852_ (.Y(_02290_),
    .B1(net3175),
    .B2(\core.work.registers.genblk1[8].latch[22] ),
    .A2(net3190),
    .A1(\core.work.registers.genblk1[3].latch[22] ));
 sg13g2_a21oi_1 _07853_ (.A1(\core.work.registers.genblk1[7].latch[22] ),
    .A2(net3024),
    .Y(_02291_),
    .B1(net3312));
 sg13g2_nand3_1 _07854_ (.B(_02290_),
    .C(_02291_),
    .A(_02289_),
    .Y(_02292_));
 sg13g2_a221oi_1 _07855_ (.B2(\core.work.registers.genblk1[5].latch[22] ),
    .C1(_02292_),
    .B1(net3004),
    .A1(\core.work.registers.genblk1[11].latch[22] ),
    .Y(_02293_),
    .A2(net3185));
 sg13g2_a22oi_1 _07856_ (.Y(_02294_),
    .B1(net3170),
    .B2(\core.work.registers.genblk1[12].latch[22] ),
    .A2(net3180),
    .A1(\core.work.registers.genblk1[15].latch[22] ));
 sg13g2_a22oi_1 _07857_ (.Y(_02295_),
    .B1(net2994),
    .B2(\core.work.registers.genblk1[6].latch[22] ),
    .A2(net2999),
    .A1(\core.work.registers.genblk1[9].latch[22] ));
 sg13g2_nand3_1 _07858_ (.B(_02294_),
    .C(_02295_),
    .A(_02288_),
    .Y(_02296_));
 sg13g2_a221oi_1 _07859_ (.B2(\core.work.registers.genblk1[4].latch[22] ),
    .C1(_02296_),
    .B1(net2984),
    .A1(\core.work.registers.genblk1[13].latch[22] ),
    .Y(_02297_),
    .A2(net3009));
 sg13g2_a22oi_1 _07860_ (.Y(_02298_),
    .B1(_02293_),
    .B2(_02297_),
    .A2(_02287_),
    .A1(net3312));
 sg13g2_o21ai_1 _07861_ (.B1(net2894),
    .Y(_02299_),
    .A1(net3032),
    .A2(_02298_));
 sg13g2_a21oi_1 _07862_ (.A1(net3489),
    .A2(_02298_),
    .Y(_02300_),
    .B1(net2891));
 sg13g2_a21oi_1 _07863_ (.A1(_00036_),
    .A2(net3028),
    .Y(_02301_),
    .B1(_02300_));
 sg13g2_nand2_1 _07864_ (.Y(_02302_),
    .A(net3331),
    .B(_02301_));
 sg13g2_a21oi_1 _07865_ (.A1(net3194),
    .A2(_02299_),
    .Y(_02303_),
    .B1(_02302_));
 sg13g2_nor2_1 _07866_ (.A(net2769),
    .B(_02303_),
    .Y(_02304_));
 sg13g2_a22oi_1 _07867_ (.Y(_00291_),
    .B1(net683),
    .B2(_02304_),
    .A2(net2775),
    .A1(_00618_));
 sg13g2_xnor2_1 _07868_ (.Y(_02305_),
    .A(_00643_),
    .B(_02071_));
 sg13g2_nand2_1 _07869_ (.Y(_02306_),
    .A(net3461),
    .B(\core.work.registers.genblk1[1].latch[23] ));
 sg13g2_nand2_1 _07870_ (.Y(_02307_),
    .A(\core.work.registers.genblk1[2].latch[23] ),
    .B(net3013));
 sg13g2_a21oi_1 _07871_ (.A1(\core.work.registers.genblk1[4].latch[23] ),
    .A2(net2983),
    .Y(_02308_),
    .B1(net3310));
 sg13g2_a22oi_1 _07872_ (.Y(_02309_),
    .B1(net3174),
    .B2(\core.work.registers.genblk1[8].latch[23] ),
    .A2(net3008),
    .A1(\core.work.registers.genblk1[13].latch[23] ));
 sg13g2_a22oi_1 _07873_ (.Y(_02310_),
    .B1(net2988),
    .B2(\core.work.registers.genblk1[10].latch[23] ),
    .A2(net2993),
    .A1(\core.work.registers.genblk1[6].latch[23] ));
 sg13g2_nand3_1 _07874_ (.B(_02309_),
    .C(_02310_),
    .A(_02308_),
    .Y(_02311_));
 sg13g2_a221oi_1 _07875_ (.B2(\core.work.registers.genblk1[12].latch[23] ),
    .C1(_02311_),
    .B1(net3169),
    .A1(\core.work.registers.genblk1[11].latch[23] ),
    .Y(_02312_),
    .A2(net3184));
 sg13g2_a22oi_1 _07876_ (.Y(_02313_),
    .B1(net2998),
    .B2(\core.work.registers.genblk1[9].latch[23] ),
    .A2(net3023),
    .A1(\core.work.registers.genblk1[7].latch[23] ));
 sg13g2_a22oi_1 _07877_ (.Y(_02314_),
    .B1(net3179),
    .B2(\core.work.registers.genblk1[15].latch[23] ),
    .A2(net3003),
    .A1(\core.work.registers.genblk1[5].latch[23] ));
 sg13g2_nand3_1 _07878_ (.B(_02313_),
    .C(_02314_),
    .A(_02307_),
    .Y(_02315_));
 sg13g2_a221oi_1 _07879_ (.B2(\core.work.registers.genblk1[3].latch[23] ),
    .C1(_02315_),
    .B1(net3189),
    .A1(\core.work.registers.genblk1[14].latch[23] ),
    .Y(_02316_),
    .A2(net3018));
 sg13g2_a22oi_1 _07880_ (.Y(_02317_),
    .B1(_02312_),
    .B2(_02316_),
    .A2(_02306_),
    .A1(net3310));
 sg13g2_o21ai_1 _07881_ (.B1(net2894),
    .Y(_02318_),
    .A1(net3032),
    .A2(_02317_));
 sg13g2_a21oi_2 _07882_ (.B1(_01646_),
    .Y(_02319_),
    .A2(_01725_),
    .A1(net3452));
 sg13g2_a21oi_1 _07883_ (.A1(net3489),
    .A2(_02317_),
    .Y(_02320_),
    .B1(net2891));
 sg13g2_a21oi_2 _07884_ (.B1(_02320_),
    .Y(_02321_),
    .A2(_02318_),
    .A1(net3194));
 sg13g2_a221oi_1 _07885_ (.B2(_02321_),
    .C1(net2773),
    .B1(_02319_),
    .A1(net3309),
    .Y(_02322_),
    .A2(_02305_));
 sg13g2_a21oi_1 _07886_ (.A1(_00616_),
    .A2(net2773),
    .Y(_00292_),
    .B1(net860));
 sg13g2_xnor2_1 _07887_ (.Y(_02323_),
    .A(_00039_),
    .B(_02198_));
 sg13g2_nand2_1 _07888_ (.Y(_02324_),
    .A(net3467),
    .B(\core.work.registers.genblk1[1].latch[24] ));
 sg13g2_nand2_1 _07889_ (.Y(_02325_),
    .A(\core.work.registers.genblk1[10].latch[24] ),
    .B(net2990));
 sg13g2_a22oi_1 _07890_ (.Y(_02326_),
    .B1(net3015),
    .B2(\core.work.registers.genblk1[2].latch[24] ),
    .A2(net3025),
    .A1(\core.work.registers.genblk1[7].latch[24] ));
 sg13g2_a22oi_1 _07891_ (.Y(_02327_),
    .B1(net3171),
    .B2(\core.work.registers.genblk1[12].latch[24] ),
    .A2(net2985),
    .A1(\core.work.registers.genblk1[4].latch[24] ));
 sg13g2_a21oi_1 _07892_ (.A1(\core.work.registers.genblk1[13].latch[24] ),
    .A2(net3010),
    .Y(_02328_),
    .B1(net3315));
 sg13g2_a22oi_1 _07893_ (.Y(_02329_),
    .B1(net2995),
    .B2(\core.work.registers.genblk1[6].latch[24] ),
    .A2(net3020),
    .A1(\core.work.registers.genblk1[14].latch[24] ));
 sg13g2_a22oi_1 _07894_ (.Y(_02330_),
    .B1(net3177),
    .B2(\core.work.registers.genblk1[8].latch[24] ),
    .A2(net3000),
    .A1(\core.work.registers.genblk1[9].latch[24] ));
 sg13g2_nand4_1 _07895_ (.B(_02328_),
    .C(_02329_),
    .A(_02327_),
    .Y(_02331_),
    .D(_02330_));
 sg13g2_a22oi_1 _07896_ (.Y(_02332_),
    .B1(net3181),
    .B2(\core.work.registers.genblk1[15].latch[24] ),
    .A2(net3191),
    .A1(\core.work.registers.genblk1[3].latch[24] ));
 sg13g2_a22oi_1 _07897_ (.Y(_02333_),
    .B1(net3005),
    .B2(\core.work.registers.genblk1[5].latch[24] ),
    .A2(net3186),
    .A1(\core.work.registers.genblk1[11].latch[24] ));
 sg13g2_nand4_1 _07898_ (.B(_02326_),
    .C(_02332_),
    .A(_02325_),
    .Y(_02334_),
    .D(_02333_));
 sg13g2_nor2_1 _07899_ (.A(_02331_),
    .B(_02334_),
    .Y(_02335_));
 sg13g2_a21oi_2 _07900_ (.B1(_02335_),
    .Y(_02336_),
    .A2(_02324_),
    .A1(net3316));
 sg13g2_o21ai_1 _07901_ (.B1(net2894),
    .Y(_02337_),
    .A1(net3033),
    .A2(_02336_));
 sg13g2_a21oi_1 _07902_ (.A1(_00040_),
    .A2(net3028),
    .Y(_02338_),
    .B1(net3329));
 sg13g2_a21oi_1 _07903_ (.A1(net3491),
    .A2(_02336_),
    .Y(_02339_),
    .B1(net2891));
 sg13g2_a21oi_1 _07904_ (.A1(_01692_),
    .A2(_02337_),
    .Y(_02340_),
    .B1(_02339_));
 sg13g2_a221oi_1 _07905_ (.B2(_02340_),
    .C1(net2769),
    .B1(_02338_),
    .A1(net3304),
    .Y(_02341_),
    .A2(_02323_));
 sg13g2_a21oi_1 _07906_ (.A1(_00614_),
    .A2(net2773),
    .Y(_00293_),
    .B1(_02341_));
 sg13g2_nor2_1 _07907_ (.A(net3300),
    .B(_02067_),
    .Y(_02342_));
 sg13g2_o21ai_1 _07908_ (.B1(net3532),
    .Y(_02343_),
    .A1(net2776),
    .A2(_02342_));
 sg13g2_nand2_1 _07909_ (.Y(_02344_),
    .A(net3464),
    .B(\core.work.registers.genblk1[1].latch[17] ));
 sg13g2_nand2_1 _07910_ (.Y(_02345_),
    .A(\core.work.registers.genblk1[8].latch[17] ),
    .B(net3176));
 sg13g2_a22oi_1 _07911_ (.Y(_02346_),
    .B1(net2995),
    .B2(\core.work.registers.genblk1[6].latch[17] ),
    .A2(net3025),
    .A1(\core.work.registers.genblk1[7].latch[17] ));
 sg13g2_a21oi_1 _07912_ (.A1(\core.work.registers.genblk1[2].latch[17] ),
    .A2(net3015),
    .Y(_02347_),
    .B1(net3315));
 sg13g2_a22oi_1 _07913_ (.Y(_02348_),
    .B1(net3000),
    .B2(\core.work.registers.genblk1[9].latch[17] ),
    .A2(net3020),
    .A1(\core.work.registers.genblk1[14].latch[17] ));
 sg13g2_a22oi_1 _07914_ (.Y(_02349_),
    .B1(net3172),
    .B2(\core.work.registers.genblk1[12].latch[17] ),
    .A2(net3192),
    .A1(\core.work.registers.genblk1[3].latch[17] ));
 sg13g2_nand3_1 _07915_ (.B(_02348_),
    .C(_02349_),
    .A(_02347_),
    .Y(_02350_));
 sg13g2_a221oi_1 _07916_ (.B2(\core.work.registers.genblk1[10].latch[17] ),
    .C1(_02350_),
    .B1(net2990),
    .A1(\core.work.registers.genblk1[15].latch[17] ),
    .Y(_02351_),
    .A2(net3181));
 sg13g2_a22oi_1 _07917_ (.Y(_02352_),
    .B1(net3005),
    .B2(\core.work.registers.genblk1[5].latch[17] ),
    .A2(net3186),
    .A1(\core.work.registers.genblk1[11].latch[17] ));
 sg13g2_nand3_1 _07918_ (.B(_02346_),
    .C(_02352_),
    .A(_02345_),
    .Y(_02353_));
 sg13g2_a221oi_1 _07919_ (.B2(\core.work.registers.genblk1[4].latch[17] ),
    .C1(_02353_),
    .B1(net2986),
    .A1(\core.work.registers.genblk1[13].latch[17] ),
    .Y(_02354_),
    .A2(net3011));
 sg13g2_a22oi_1 _07920_ (.Y(_02355_),
    .B1(_02351_),
    .B2(_02354_),
    .A2(_02344_),
    .A1(net3317));
 sg13g2_o21ai_1 _07921_ (.B1(net2896),
    .Y(_02356_),
    .A1(net3036),
    .A2(_02355_));
 sg13g2_a21oi_1 _07922_ (.A1(net3494),
    .A2(_02355_),
    .Y(_02357_),
    .B1(net2893));
 sg13g2_a221oi_1 _07923_ (.B2(net3196),
    .C1(_02357_),
    .B1(_02356_),
    .A1(_00025_),
    .Y(_02358_),
    .A2(net3030));
 sg13g2_nor2_1 _07924_ (.A(net3532),
    .B(net3300),
    .Y(_02359_));
 sg13g2_a22oi_1 _07925_ (.Y(_02360_),
    .B1(_02359_),
    .B2(_02067_),
    .A2(_02358_),
    .A1(_01645_));
 sg13g2_o21ai_1 _07926_ (.B1(_02343_),
    .Y(_00294_),
    .A1(net2775),
    .A2(_02360_));
 sg13g2_nand2_1 _07927_ (.Y(_02361_),
    .A(_00027_),
    .B(_02067_));
 sg13g2_o21ai_1 _07928_ (.B1(net3309),
    .Y(_02362_),
    .A1(net709),
    .A2(_02361_));
 sg13g2_a21o_1 _07929_ (.A2(_02361_),
    .A1(net709),
    .B1(_02362_),
    .X(_02363_));
 sg13g2_nand2_1 _07930_ (.Y(_02364_),
    .A(net3467),
    .B(\core.work.registers.genblk1[1].latch[18] ));
 sg13g2_nand2_1 _07931_ (.Y(_02365_),
    .A(\core.work.registers.genblk1[7].latch[18] ),
    .B(net3025));
 sg13g2_a22oi_1 _07932_ (.Y(_02366_),
    .B1(net2990),
    .B2(\core.work.registers.genblk1[10].latch[18] ),
    .A2(net3000),
    .A1(\core.work.registers.genblk1[9].latch[18] ));
 sg13g2_a22oi_1 _07933_ (.Y(_02367_),
    .B1(net3171),
    .B2(\core.work.registers.genblk1[12].latch[18] ),
    .A2(net3177),
    .A1(\core.work.registers.genblk1[8].latch[18] ));
 sg13g2_a22oi_1 _07934_ (.Y(_02368_),
    .B1(net2995),
    .B2(\core.work.registers.genblk1[6].latch[18] ),
    .A2(net3191),
    .A1(\core.work.registers.genblk1[3].latch[18] ));
 sg13g2_a21oi_1 _07935_ (.A1(\core.work.registers.genblk1[14].latch[18] ),
    .A2(net3020),
    .Y(_02369_),
    .B1(net3315));
 sg13g2_a22oi_1 _07936_ (.Y(_02370_),
    .B1(net3005),
    .B2(\core.work.registers.genblk1[5].latch[18] ),
    .A2(net3010),
    .A1(\core.work.registers.genblk1[13].latch[18] ));
 sg13g2_nand4_1 _07937_ (.B(_02367_),
    .C(_02369_),
    .A(_02366_),
    .Y(_02371_),
    .D(_02370_));
 sg13g2_a22oi_1 _07938_ (.Y(_02372_),
    .B1(net2985),
    .B2(\core.work.registers.genblk1[4].latch[18] ),
    .A2(net3181),
    .A1(\core.work.registers.genblk1[15].latch[18] ));
 sg13g2_a22oi_1 _07939_ (.Y(_02373_),
    .B1(net3186),
    .B2(\core.work.registers.genblk1[11].latch[18] ),
    .A2(net3015),
    .A1(\core.work.registers.genblk1[2].latch[18] ));
 sg13g2_nand4_1 _07940_ (.B(_02368_),
    .C(_02372_),
    .A(_02365_),
    .Y(_02374_),
    .D(_02373_));
 sg13g2_nor2_2 _07941_ (.A(_02371_),
    .B(_02374_),
    .Y(_02375_));
 sg13g2_a21oi_2 _07942_ (.B1(_02375_),
    .Y(_02376_),
    .A2(_02364_),
    .A1(net3316));
 sg13g2_o21ai_1 _07943_ (.B1(net2894),
    .Y(_02377_),
    .A1(net3032),
    .A2(_02376_));
 sg13g2_a21oi_1 _07944_ (.A1(_00028_),
    .A2(net3028),
    .Y(_02378_),
    .B1(net3329));
 sg13g2_a21oi_1 _07945_ (.A1(net3489),
    .A2(_02376_),
    .Y(_02379_),
    .B1(net2891));
 sg13g2_a21oi_1 _07946_ (.A1(net3195),
    .A2(_02377_),
    .Y(_02380_),
    .B1(_02379_));
 sg13g2_a21oi_2 _07947_ (.B1(net2769),
    .Y(_02381_),
    .A2(_02380_),
    .A1(_02378_));
 sg13g2_a22oi_1 _07948_ (.Y(_00295_),
    .B1(net710),
    .B2(_02381_),
    .A2(net2775),
    .A1(_00625_));
 sg13g2_a21oi_1 _07949_ (.A1(net721),
    .A2(_02068_),
    .Y(_02382_),
    .B1(net3300));
 sg13g2_o21ai_1 _07950_ (.B1(_02382_),
    .Y(_02383_),
    .A1(net721),
    .A2(_02068_));
 sg13g2_nand2_1 _07951_ (.Y(_02384_),
    .A(net3466),
    .B(\core.work.registers.genblk1[1].latch[19] ));
 sg13g2_nand2_1 _07952_ (.Y(_02385_),
    .A(\core.work.registers.genblk1[13].latch[19] ),
    .B(net3011));
 sg13g2_a22oi_1 _07953_ (.Y(_02386_),
    .B1(net3172),
    .B2(\core.work.registers.genblk1[12].latch[19] ),
    .A2(net2996),
    .A1(\core.work.registers.genblk1[6].latch[19] ));
 sg13g2_a22oi_1 _07954_ (.Y(_02387_),
    .B1(net2986),
    .B2(\core.work.registers.genblk1[4].latch[19] ),
    .A2(net3006),
    .A1(\core.work.registers.genblk1[5].latch[19] ));
 sg13g2_a21oi_1 _07955_ (.A1(\core.work.registers.genblk1[10].latch[19] ),
    .A2(net2991),
    .Y(_02388_),
    .B1(net3318));
 sg13g2_a22oi_1 _07956_ (.Y(_02389_),
    .B1(net3016),
    .B2(\core.work.registers.genblk1[2].latch[19] ),
    .A2(net3026),
    .A1(\core.work.registers.genblk1[7].latch[19] ));
 sg13g2_a22oi_1 _07957_ (.Y(_02390_),
    .B1(net3176),
    .B2(\core.work.registers.genblk1[8].latch[19] ),
    .A2(net3021),
    .A1(\core.work.registers.genblk1[14].latch[19] ));
 sg13g2_nand4_1 _07958_ (.B(_02388_),
    .C(_02389_),
    .A(_02387_),
    .Y(_02391_),
    .D(_02390_));
 sg13g2_a22oi_1 _07959_ (.Y(_02392_),
    .B1(net3182),
    .B2(\core.work.registers.genblk1[15].latch[19] ),
    .A2(net3187),
    .A1(\core.work.registers.genblk1[11].latch[19] ));
 sg13g2_a22oi_1 _07960_ (.Y(_02393_),
    .B1(net3001),
    .B2(\core.work.registers.genblk1[9].latch[19] ),
    .A2(net3192),
    .A1(\core.work.registers.genblk1[3].latch[19] ));
 sg13g2_nand4_1 _07961_ (.B(_02386_),
    .C(_02392_),
    .A(_02385_),
    .Y(_02394_),
    .D(_02393_));
 sg13g2_nor2_1 _07962_ (.A(_02391_),
    .B(_02394_),
    .Y(_02395_));
 sg13g2_a21oi_2 _07963_ (.B1(_02395_),
    .Y(_02396_),
    .A2(_02384_),
    .A1(net3318));
 sg13g2_o21ai_1 _07964_ (.B1(net2896),
    .Y(_02397_),
    .A1(net3036),
    .A2(_02396_));
 sg13g2_a21oi_1 _07965_ (.A1(_00030_),
    .A2(net3030),
    .Y(_02398_),
    .B1(net3330));
 sg13g2_a21oi_1 _07966_ (.A1(net3494),
    .A2(_02396_),
    .Y(_02399_),
    .B1(net2893));
 sg13g2_a21oi_1 _07967_ (.A1(net3196),
    .A2(_02397_),
    .Y(_02400_),
    .B1(_02399_));
 sg13g2_a21oi_1 _07968_ (.A1(_02398_),
    .A2(_02400_),
    .Y(_02401_),
    .B1(net2775));
 sg13g2_a22oi_1 _07969_ (.Y(_00296_),
    .B1(_02383_),
    .B2(_02401_),
    .A2(net2775),
    .A1(_00624_));
 sg13g2_xnor2_1 _07970_ (.Y(_02402_),
    .A(_00031_),
    .B(_02262_));
 sg13g2_nand2_1 _07971_ (.Y(_02403_),
    .A(net3467),
    .B(\core.work.registers.genblk1[1].latch[20] ));
 sg13g2_nand2_1 _07972_ (.Y(_02404_),
    .A(\core.work.registers.genblk1[9].latch[20] ),
    .B(net3000));
 sg13g2_a22oi_1 _07973_ (.Y(_02405_),
    .B1(net3171),
    .B2(\core.work.registers.genblk1[12].latch[20] ),
    .A2(net2995),
    .A1(\core.work.registers.genblk1[6].latch[20] ));
 sg13g2_a21oi_1 _07974_ (.A1(\core.work.registers.genblk1[2].latch[20] ),
    .A2(net3015),
    .Y(_02406_),
    .B1(net3315));
 sg13g2_a22oi_1 _07975_ (.Y(_02407_),
    .B1(net2985),
    .B2(\core.work.registers.genblk1[4].latch[20] ),
    .A2(net3010),
    .A1(\core.work.registers.genblk1[13].latch[20] ));
 sg13g2_a22oi_1 _07976_ (.Y(_02408_),
    .B1(net3181),
    .B2(\core.work.registers.genblk1[15].latch[20] ),
    .A2(net3020),
    .A1(\core.work.registers.genblk1[14].latch[20] ));
 sg13g2_nand3_1 _07977_ (.B(_02407_),
    .C(_02408_),
    .A(_02406_),
    .Y(_02409_));
 sg13g2_a221oi_1 _07978_ (.B2(\core.work.registers.genblk1[11].latch[20] ),
    .C1(_02409_),
    .B1(net3186),
    .A1(\core.work.registers.genblk1[7].latch[20] ),
    .Y(_02410_),
    .A2(net3025));
 sg13g2_a22oi_1 _07979_ (.Y(_02411_),
    .B1(net2990),
    .B2(\core.work.registers.genblk1[10].latch[20] ),
    .A2(net3191),
    .A1(\core.work.registers.genblk1[3].latch[20] ));
 sg13g2_nand3_1 _07980_ (.B(_02405_),
    .C(_02411_),
    .A(_02404_),
    .Y(_02412_));
 sg13g2_a221oi_1 _07981_ (.B2(\core.work.registers.genblk1[8].latch[20] ),
    .C1(_02412_),
    .B1(net3177),
    .A1(\core.work.registers.genblk1[5].latch[20] ),
    .Y(_02413_),
    .A2(net3005));
 sg13g2_a22oi_1 _07982_ (.Y(_02414_),
    .B1(_02410_),
    .B2(_02413_),
    .A2(_02403_),
    .A1(net3316));
 sg13g2_o21ai_1 _07983_ (.B1(net2896),
    .Y(_02415_),
    .A1(net3036),
    .A2(_02414_));
 sg13g2_a21oi_1 _07984_ (.A1(_00032_),
    .A2(net3030),
    .Y(_02416_),
    .B1(net3330));
 sg13g2_a21oi_1 _07985_ (.A1(net3494),
    .A2(_02414_),
    .Y(_02417_),
    .B1(net2893));
 sg13g2_a21oi_1 _07986_ (.A1(net3196),
    .A2(_02415_),
    .Y(_02418_),
    .B1(_02417_));
 sg13g2_a221oi_1 _07987_ (.B2(_02418_),
    .C1(net2776),
    .B1(_02416_),
    .A1(net3309),
    .Y(_02419_),
    .A2(_02402_));
 sg13g2_a21oi_1 _07988_ (.A1(_00621_),
    .A2(net2775),
    .Y(_00297_),
    .B1(_02419_));
 sg13g2_nor2_1 _07989_ (.A(_01327_),
    .B(_01371_),
    .Y(_02420_));
 sg13g2_nand2b_1 _07990_ (.Y(_02421_),
    .B(net2737),
    .A_N(_01138_));
 sg13g2_nand3_1 _07991_ (.B(_00986_),
    .C(_01330_),
    .A(net3565),
    .Y(_02422_));
 sg13g2_a21oi_1 _07992_ (.A1(_01331_),
    .A2(_02422_),
    .Y(_02423_),
    .B1(net2737));
 sg13g2_nor3_1 _07993_ (.A(net2737),
    .B(_01327_),
    .C(net3042),
    .Y(_02424_));
 sg13g2_nor3_2 _07994_ (.A(_01138_),
    .B(_02423_),
    .C(_02424_),
    .Y(_02425_));
 sg13g2_a21oi_1 _07995_ (.A1(net2886),
    .A2(_02425_),
    .Y(_02426_),
    .B1(net364));
 sg13g2_a21o_1 _07996_ (.A2(net2886),
    .A1(net3529),
    .B1(net2737),
    .X(_02427_));
 sg13g2_a21oi_1 _07997_ (.A1(_02425_),
    .A2(_02427_),
    .Y(_00298_),
    .B1(_02426_));
 sg13g2_nand2_2 _07998_ (.Y(_02428_),
    .A(\core.lsu.state[0] ),
    .B(\core.lsu.state[1] ));
 sg13g2_nor2_2 _07999_ (.A(_00021_),
    .B(_02428_),
    .Y(_02429_));
 sg13g2_o21ai_1 _08000_ (.B1(_02429_),
    .Y(_02430_),
    .A1(\core.lsu.dreg[0] ),
    .A2(\core.lsu.dreg[3] ));
 sg13g2_o21ai_1 _08001_ (.B1(_02429_),
    .Y(_02431_),
    .A1(\core.lsu.dreg[1] ),
    .A2(\core.lsu.dreg[2] ));
 sg13g2_and2_2 _08002_ (.A(_02430_),
    .B(_02431_),
    .X(_02432_));
 sg13g2_inv_1 _08003_ (.Y(_02433_),
    .A(net2871));
 sg13g2_nand4_1 _08004_ (.B(\core.work.state[0] ),
    .C(_01314_),
    .A(net3501),
    .Y(_02434_),
    .D(_01718_));
 sg13g2_nor2_2 _08005_ (.A(_02433_),
    .B(_02434_),
    .Y(_02435_));
 sg13g2_nor4_2 _08006_ (.A(\core.work.dreg[1] ),
    .B(\core.work.dreg[0] ),
    .C(\core.work.dreg[3] ),
    .Y(_02436_),
    .D(\core.work.dreg[2] ));
 sg13g2_inv_1 _08007_ (.Y(_02437_),
    .A(_02436_));
 sg13g2_o21ai_1 _08008_ (.B1(net2871),
    .Y(_02438_),
    .A1(_02434_),
    .A2(_02436_));
 sg13g2_nor2_1 _08009_ (.A(\core.work.registers.state[2] ),
    .B(_00735_),
    .Y(_02439_));
 sg13g2_and3_2 _08010_ (.X(_02440_),
    .A(net3581),
    .B(_02438_),
    .C(_02439_));
 sg13g2_a22oi_1 _08011_ (.Y(_02441_),
    .B1(_02435_),
    .B2(\core.work.dreg[0] ),
    .A2(_02429_),
    .A1(\core.lsu.dreg[0] ));
 sg13g2_nor2_1 _08012_ (.A(net526),
    .B(net2808),
    .Y(_02442_));
 sg13g2_a21oi_1 _08013_ (.A1(net2808),
    .A2(_02441_),
    .Y(_00299_),
    .B1(_02442_));
 sg13g2_nor2_1 _08014_ (.A(net568),
    .B(net2808),
    .Y(_02443_));
 sg13g2_a22oi_1 _08015_ (.Y(_02444_),
    .B1(_02435_),
    .B2(net562),
    .A2(_02429_),
    .A1(\core.lsu.dreg[1] ));
 sg13g2_a21oi_1 _08016_ (.A1(net2808),
    .A2(_02444_),
    .Y(_00300_),
    .B1(_02443_));
 sg13g2_nor2_1 _08017_ (.A(net671),
    .B(net2808),
    .Y(_02445_));
 sg13g2_a22oi_1 _08018_ (.Y(_02446_),
    .B1(_02435_),
    .B2(net392),
    .A2(_02429_),
    .A1(\core.lsu.dreg[2] ));
 sg13g2_a21oi_1 _08019_ (.A1(net2808),
    .A2(_02446_),
    .Y(_00301_),
    .B1(_02445_));
 sg13g2_a22oi_1 _08020_ (.Y(_02447_),
    .B1(_02435_),
    .B2(net414),
    .A2(_02429_),
    .A1(\core.lsu.dreg[3] ));
 sg13g2_nor2_1 _08021_ (.A(net690),
    .B(net2808),
    .Y(_02448_));
 sg13g2_a21oi_1 _08022_ (.A1(net2808),
    .A2(_02447_),
    .Y(_00302_),
    .B1(_02448_));
 sg13g2_a21oi_1 _08023_ (.A1(net513),
    .A2(net3298),
    .Y(_02449_),
    .B1(net2787));
 sg13g2_a21oi_1 _08024_ (.A1(net2908),
    .A2(net2787),
    .Y(_00303_),
    .B1(_02449_));
 sg13g2_nor2_1 _08025_ (.A(net3344),
    .B(net2884),
    .Y(_02450_));
 sg13g2_a21o_1 _08026_ (.A2(net2886),
    .A1(net3529),
    .B1(net2839),
    .X(_02451_));
 sg13g2_nand3_1 _08027_ (.B(_02425_),
    .C(_02451_),
    .A(net3528),
    .Y(_02452_));
 sg13g2_a21o_1 _08028_ (.A2(_02451_),
    .A1(_02425_),
    .B1(net3528),
    .X(_02453_));
 sg13g2_and3_1 _08029_ (.X(_00304_),
    .A(_02421_),
    .B(_02452_),
    .C(_02453_));
 sg13g2_nand2_1 _08030_ (.Y(_02454_),
    .A(net3528),
    .B(net3529));
 sg13g2_nor2_1 _08031_ (.A(net3527),
    .B(_02454_),
    .Y(_02455_));
 sg13g2_and2_1 _08032_ (.A(net3527),
    .B(_02454_),
    .X(_02456_));
 sg13g2_o21ai_1 _08033_ (.B1(net2886),
    .Y(_02457_),
    .A1(net3159),
    .A2(_02456_));
 sg13g2_nand2_1 _08034_ (.Y(_02458_),
    .A(_01326_),
    .B(_01371_));
 sg13g2_o21ai_1 _08035_ (.B1(_02458_),
    .Y(_02459_),
    .A1(_01146_),
    .A2(net3348));
 sg13g2_o21ai_1 _08036_ (.B1(_02459_),
    .Y(_02460_),
    .A1(_01323_),
    .A2(_01371_));
 sg13g2_a21oi_1 _08037_ (.A1(_02457_),
    .A2(_02460_),
    .Y(_02461_),
    .B1(net2737));
 sg13g2_nand2_1 _08038_ (.Y(_02462_),
    .A(_02425_),
    .B(_02461_));
 sg13g2_o21ai_1 _08039_ (.B1(_02462_),
    .Y(_00305_),
    .A1(_00580_),
    .A2(_02425_));
 sg13g2_nand2b_1 _08040_ (.Y(_02463_),
    .B(net678),
    .A_N(net3574));
 sg13g2_nor2b_1 _08041_ (.A(_00991_),
    .B_N(_01544_),
    .Y(_02464_));
 sg13g2_nand2b_2 _08042_ (.Y(_02465_),
    .B(net3574),
    .A_N(_02464_));
 sg13g2_xnor2_1 _08043_ (.Y(_02466_),
    .A(net678),
    .B(net3572));
 sg13g2_o21ai_1 _08044_ (.B1(_02463_),
    .Y(_00306_),
    .A1(_02465_),
    .A2(_02466_));
 sg13g2_nand2b_1 _08045_ (.Y(_02467_),
    .B(\core.fetch.spi_reader.counter[1] ),
    .A_N(net3574));
 sg13g2_nor2_1 _08046_ (.A(net3572),
    .B(net365),
    .Y(_02468_));
 sg13g2_xnor2_1 _08047_ (.Y(_02469_),
    .A(\core.fetch.spi_reader.counter[1] ),
    .B(\core.fetch.spi_reader.counter[0] ));
 sg13g2_a21oi_1 _08048_ (.A1(net3572),
    .A2(_02469_),
    .Y(_02470_),
    .B1(_02468_));
 sg13g2_o21ai_1 _08049_ (.B1(_02467_),
    .Y(_00307_),
    .A1(_02465_),
    .A2(_02470_));
 sg13g2_nand2b_1 _08050_ (.Y(_02471_),
    .B(\core.fetch.spi_reader.counter[2] ),
    .A_N(net3574));
 sg13g2_nand2_2 _08051_ (.Y(_02472_),
    .A(net3572),
    .B(_00983_));
 sg13g2_xnor2_1 _08052_ (.Y(_02473_),
    .A(net431),
    .B(_02472_));
 sg13g2_o21ai_1 _08053_ (.B1(_02471_),
    .Y(_00308_),
    .A1(_02465_),
    .A2(_02473_));
 sg13g2_nand2b_1 _08054_ (.Y(_02474_),
    .B(net433),
    .A_N(net3574));
 sg13g2_nor2_1 _08055_ (.A(\core.fetch.spi_reader.counter[2] ),
    .B(_02472_),
    .Y(_02475_));
 sg13g2_xnor2_1 _08056_ (.Y(_02476_),
    .A(_00165_),
    .B(_02475_));
 sg13g2_nor2_1 _08057_ (.A(net3565),
    .B(_02476_),
    .Y(_02477_));
 sg13g2_nor2_1 _08058_ (.A(_00833_),
    .B(_00942_),
    .Y(_02478_));
 sg13g2_nand4_1 _08059_ (.B(_00978_),
    .C(_01462_),
    .A(net3565),
    .Y(_02479_),
    .D(_02478_));
 sg13g2_nor2b_1 _08060_ (.A(_02477_),
    .B_N(_02479_),
    .Y(_02480_));
 sg13g2_o21ai_1 _08061_ (.B1(_02476_),
    .Y(_02481_),
    .A1(_00990_),
    .A2(_01543_));
 sg13g2_nand2_1 _08062_ (.Y(_02482_),
    .A(_00988_),
    .B(_02481_));
 sg13g2_a221oi_1 _08063_ (.B2(_00748_),
    .C1(_02482_),
    .B1(_02480_),
    .A1(net3200),
    .Y(_02483_),
    .A2(_01543_));
 sg13g2_o21ai_1 _08064_ (.B1(net3575),
    .Y(_02484_),
    .A1(_00988_),
    .A2(_02476_));
 sg13g2_o21ai_1 _08065_ (.B1(_02474_),
    .Y(_00309_),
    .A1(_02483_),
    .A2(_02484_));
 sg13g2_nor3_1 _08066_ (.A(\core.fetch.spi_reader.counter[3] ),
    .B(\core.fetch.spi_reader.counter[2] ),
    .C(_02472_),
    .Y(_02485_));
 sg13g2_xor2_1 _08067_ (.B(_02485_),
    .A(_00166_),
    .X(_02486_));
 sg13g2_nand2_1 _08068_ (.Y(_02487_),
    .A(_00833_),
    .B(_00834_));
 sg13g2_nor3_1 _08069_ (.A(net3362),
    .B(_00749_),
    .C(_00835_),
    .Y(_02488_));
 sg13g2_nand4_1 _08070_ (.B(_01462_),
    .C(_02487_),
    .A(_00978_),
    .Y(_02489_),
    .D(_02488_));
 sg13g2_o21ai_1 _08071_ (.B1(_02489_),
    .Y(_02490_),
    .A1(_02464_),
    .A2(_02486_));
 sg13g2_mux2_1 _08072_ (.A0(net376),
    .A1(_02490_),
    .S(net3574),
    .X(_00310_));
 sg13g2_nand2b_1 _08073_ (.Y(_02491_),
    .B(net425),
    .A_N(net3574));
 sg13g2_nor2_1 _08074_ (.A(_00982_),
    .B(_02472_),
    .Y(_02492_));
 sg13g2_xor2_1 _08075_ (.B(_02492_),
    .A(_00167_),
    .X(_02493_));
 sg13g2_o21ai_1 _08076_ (.B1(_02491_),
    .Y(_00311_),
    .A1(_02465_),
    .A2(_02493_));
 sg13g2_nand2_2 _08077_ (.Y(_02494_),
    .A(net3588),
    .B(_00001_));
 sg13g2_nor2_1 _08078_ (.A(net823),
    .B(net2864),
    .Y(_02495_));
 sg13g2_a21oi_1 _08079_ (.A1(_00652_),
    .A2(net2868),
    .Y(_00312_),
    .B1(_02495_));
 sg13g2_nand2_1 _08080_ (.Y(_02496_),
    .A(net395),
    .B(net2865));
 sg13g2_o21ai_1 _08081_ (.B1(_02496_),
    .Y(_00313_),
    .A1(_00591_),
    .A2(net2866));
 sg13g2_mux2_1 _08082_ (.A0(net3498),
    .A1(net814),
    .S(net2866),
    .X(_00314_));
 sg13g2_nor2_1 _08083_ (.A(net3496),
    .B(net2868),
    .Y(_02497_));
 sg13g2_a21oi_1 _08084_ (.A1(_00653_),
    .A2(net2868),
    .Y(_00315_),
    .B1(_02497_));
 sg13g2_nor2_1 _08085_ (.A(net3495),
    .B(net2866),
    .Y(_02498_));
 sg13g2_a21oi_1 _08086_ (.A1(_00654_),
    .A2(net2866),
    .Y(_00316_),
    .B1(_02498_));
 sg13g2_nand2_1 _08087_ (.Y(_02499_),
    .A(net447),
    .B(net2865));
 sg13g2_o21ai_1 _08088_ (.B1(_02499_),
    .Y(_00317_),
    .A1(_00595_),
    .A2(net2865));
 sg13g2_nand2_1 _08089_ (.Y(_02500_),
    .A(net381),
    .B(net2865));
 sg13g2_o21ai_1 _08090_ (.B1(_02500_),
    .Y(_00318_),
    .A1(_00594_),
    .A2(net2866));
 sg13g2_nand2_1 _08091_ (.Y(_02501_),
    .A(net369),
    .B(net2865));
 sg13g2_o21ai_1 _08092_ (.B1(_02501_),
    .Y(_00319_),
    .A1(_00593_),
    .A2(net2865));
 sg13g2_nor2_1 _08093_ (.A(\core.e2m_addr[8] ),
    .B(net2866),
    .Y(_02502_));
 sg13g2_a21oi_1 _08094_ (.A1(_00655_),
    .A2(net2865),
    .Y(_00320_),
    .B1(_02502_));
 sg13g2_mux2_1 _08095_ (.A0(net3488),
    .A1(net734),
    .S(net2865),
    .X(_00321_));
 sg13g2_mux2_1 _08096_ (.A0(net3487),
    .A1(\core.fetch.rd_addr_i[10] ),
    .S(net2867),
    .X(_00322_));
 sg13g2_mux2_1 _08097_ (.A0(\core.e2m_addr[11] ),
    .A1(net632),
    .S(net2867),
    .X(_00323_));
 sg13g2_nand2_1 _08098_ (.Y(_02503_),
    .A(net3525),
    .B(net2864));
 sg13g2_o21ai_1 _08099_ (.B1(_02503_),
    .Y(_00324_),
    .A1(_00601_),
    .A2(net2864));
 sg13g2_mux2_1 _08100_ (.A0(net3483),
    .A1(net630),
    .S(net2864),
    .X(_00325_));
 sg13g2_nand2_1 _08101_ (.Y(_02504_),
    .A(net378),
    .B(net2864));
 sg13g2_o21ai_1 _08102_ (.B1(_02504_),
    .Y(_00326_),
    .A1(_00600_),
    .A2(net2864));
 sg13g2_nand2_1 _08103_ (.Y(_02505_),
    .A(net375),
    .B(net2864));
 sg13g2_o21ai_1 _08104_ (.B1(_02505_),
    .Y(_00327_),
    .A1(_00599_),
    .A2(net2864));
 sg13g2_nor4_1 _08105_ (.A(\core.fetch.rd_addr_i[5] ),
    .B(\core.fetch.rd_addr_i[4] ),
    .C(\core.fetch.rd_addr_i[7] ),
    .D(\core.fetch.rd_addr_i[6] ),
    .Y(_02506_));
 sg13g2_nor4_1 _08106_ (.A(net3526),
    .B(\core.fetch.rd_addr_i[0] ),
    .C(\core.fetch.rd_addr_i[3] ),
    .D(\core.fetch.rd_addr_i[2] ),
    .Y(_02507_));
 sg13g2_or2_1 _08107_ (.X(_02508_),
    .B(\core.fetch.rd_addr_i[8] ),
    .A(\core.fetch.rd_addr_i[9] ));
 sg13g2_nor4_1 _08108_ (.A(\core.fetch.rd_addr_i[13] ),
    .B(net3525),
    .C(\core.fetch.rd_addr_i[15] ),
    .D(\core.fetch.rd_addr_i[14] ),
    .Y(_02509_));
 sg13g2_nand3_1 _08109_ (.B(_02507_),
    .C(_02509_),
    .A(_02506_),
    .Y(_02510_));
 sg13g2_nor4_2 _08110_ (.A(net632),
    .B(\core.fetch.rd_addr_i[10] ),
    .C(_02508_),
    .Y(_02511_),
    .D(_02510_));
 sg13g2_nand3_1 _08111_ (.B(\core.fetch.rd_addr_i[3] ),
    .C(\core.fetch.rd_addr_i[2] ),
    .A(net3526),
    .Y(_02512_));
 sg13g2_nor3_1 _08112_ (.A(net3523),
    .B(_00652_),
    .C(_02512_),
    .Y(_02513_));
 sg13g2_nand4_1 _08113_ (.B(net3525),
    .C(\core.fetch.rd_addr_i[15] ),
    .A(\core.fetch.rd_addr_i[13] ),
    .Y(_02514_),
    .D(\core.fetch.rd_addr_i[14] ));
 sg13g2_nor3_2 _08114_ (.A(_00751_),
    .B(_00753_),
    .C(_02514_),
    .Y(_02515_));
 sg13g2_nor3_2 _08115_ (.A(_00751_),
    .B(_00753_),
    .C(_02514_),
    .Y(_02516_));
 sg13g2_and2_1 _08116_ (.A(_02513_),
    .B(_02516_),
    .X(_02517_));
 sg13g2_or2_1 _08117_ (.X(_02518_),
    .B(net2979),
    .A(net2982));
 sg13g2_nor4_1 _08118_ (.A(net3523),
    .B(\core.lsu.is_half ),
    .C(net3526),
    .D(_00652_),
    .Y(_02519_));
 sg13g2_nor4_2 _08119_ (.A(net3523),
    .B(\core.lsu.is_half ),
    .C(\core.fetch.rd_addr_i[0] ),
    .Y(_02520_),
    .D(_02512_));
 sg13g2_nand2_1 _08120_ (.Y(_02521_),
    .A(_02516_),
    .B(_02520_));
 sg13g2_inv_1 _08121_ (.Y(_02522_),
    .A(net2978));
 sg13g2_and4_1 _08122_ (.A(\core.fetch.rd_addr_i[3] ),
    .B(\core.fetch.rd_addr_i[2] ),
    .C(_02516_),
    .D(_02519_),
    .X(_02523_));
 sg13g2_nor3_2 _08123_ (.A(net2862),
    .B(_02522_),
    .C(net2976),
    .Y(_02524_));
 sg13g2_nor2_1 _08124_ (.A(_00634_),
    .B(_02428_),
    .Y(_02525_));
 sg13g2_nor4_2 _08125_ (.A(_00634_),
    .B(_00059_),
    .C(_02428_),
    .Y(_02526_),
    .D(_02524_));
 sg13g2_nand2b_1 _08126_ (.Y(_02527_),
    .B(_02521_),
    .A_N(\core.gpio.stray_data_i[24] ));
 sg13g2_o21ai_1 _08127_ (.B1(_02527_),
    .Y(_02528_),
    .A1(\core.gpio.stray_data_i[16] ),
    .A2(net2977));
 sg13g2_a22oi_1 _08128_ (.Y(_02529_),
    .B1(net2979),
    .B2(\core.gpio.stray_data_i[8] ),
    .A2(net2981),
    .A1(\core.gpio.stray_data_i[0] ));
 sg13g2_o21ai_1 _08129_ (.B1(_02529_),
    .Y(_02530_),
    .A1(_02518_),
    .A2(_02528_));
 sg13g2_mux2_1 _08130_ (.A0(net661),
    .A1(_02530_),
    .S(_02526_),
    .X(_00328_));
 sg13g2_nand2b_1 _08131_ (.Y(_02531_),
    .B(net2977),
    .A_N(\core.gpio.stray_data_i[25] ));
 sg13g2_o21ai_1 _08132_ (.B1(_02531_),
    .Y(_02532_),
    .A1(\core.gpio.stray_data_i[17] ),
    .A2(net2977));
 sg13g2_a22oi_1 _08133_ (.Y(_02533_),
    .B1(net2979),
    .B2(\core.gpio.stray_data_i[9] ),
    .A2(net2981),
    .A1(\core.gpio.stray_data_i[1] ));
 sg13g2_o21ai_1 _08134_ (.B1(_02533_),
    .Y(_02534_),
    .A1(net2862),
    .A2(_02532_));
 sg13g2_mux2_1 _08135_ (.A0(net567),
    .A1(_02534_),
    .S(_02526_),
    .X(_00329_));
 sg13g2_nand2b_1 _08136_ (.Y(_02535_),
    .B(net2977),
    .A_N(\core.gpio.stray_data_i[26] ));
 sg13g2_o21ai_1 _08137_ (.B1(_02535_),
    .Y(_02536_),
    .A1(\core.gpio.stray_data_i[18] ),
    .A2(net2977));
 sg13g2_a22oi_1 _08138_ (.Y(_02537_),
    .B1(net2979),
    .B2(\core.gpio.stray_data_i[10] ),
    .A2(net2982),
    .A1(\core.gpio.stray_data_i[2] ));
 sg13g2_o21ai_1 _08139_ (.B1(_02537_),
    .Y(_02538_),
    .A1(net2862),
    .A2(_02536_));
 sg13g2_mux2_1 _08140_ (.A0(net611),
    .A1(_02538_),
    .S(_02526_),
    .X(_00330_));
 sg13g2_nand2b_1 _08141_ (.Y(_02539_),
    .B(net2977),
    .A_N(\core.gpio.stray_data_i[27] ));
 sg13g2_o21ai_1 _08142_ (.B1(_02539_),
    .Y(_02540_),
    .A1(\core.gpio.stray_data_i[19] ),
    .A2(_02521_));
 sg13g2_a22oi_1 _08143_ (.Y(_02541_),
    .B1(net2979),
    .B2(\core.gpio.stray_data_i[11] ),
    .A2(net2981),
    .A1(net899));
 sg13g2_o21ai_1 _08144_ (.B1(_02541_),
    .Y(_02542_),
    .A1(net2862),
    .A2(_02540_));
 sg13g2_mux2_1 _08145_ (.A0(net660),
    .A1(_02542_),
    .S(_02526_),
    .X(_00331_));
 sg13g2_nand2b_1 _08146_ (.Y(_02543_),
    .B(net2977),
    .A_N(\core.gpio.stray_data_i[28] ));
 sg13g2_o21ai_1 _08147_ (.B1(_02543_),
    .Y(_02544_),
    .A1(\core.gpio.stray_data_i[20] ),
    .A2(net2977));
 sg13g2_a22oi_1 _08148_ (.Y(_02545_),
    .B1(net2979),
    .B2(\core.gpio.stray_data_i[12] ),
    .A2(net2981),
    .A1(\core.gpio.stray_data_i[4] ));
 sg13g2_o21ai_1 _08149_ (.B1(_02545_),
    .Y(_02546_),
    .A1(net2862),
    .A2(_02544_));
 sg13g2_mux2_1 _08150_ (.A0(net639),
    .A1(_02546_),
    .S(_02526_),
    .X(_00332_));
 sg13g2_nand2b_1 _08151_ (.Y(_02547_),
    .B(net2978),
    .A_N(\core.gpio.stray_data_i[29] ));
 sg13g2_o21ai_1 _08152_ (.B1(_02547_),
    .Y(_02548_),
    .A1(\core.gpio.stray_data_i[21] ),
    .A2(net2978));
 sg13g2_a22oi_1 _08153_ (.Y(_02549_),
    .B1(net2980),
    .B2(\core.gpio.stray_data_i[13] ),
    .A2(net2982),
    .A1(\core.gpio.stray_data_i[5] ));
 sg13g2_o21ai_1 _08154_ (.B1(_02549_),
    .Y(_02550_),
    .A1(net2862),
    .A2(_02548_));
 sg13g2_mux2_1 _08155_ (.A0(net608),
    .A1(_02550_),
    .S(_02526_),
    .X(_00333_));
 sg13g2_nand2b_1 _08156_ (.Y(_02551_),
    .B(net2978),
    .A_N(\core.gpio.stray_data_i[30] ));
 sg13g2_o21ai_1 _08157_ (.B1(_02551_),
    .Y(_02552_),
    .A1(\core.gpio.stray_data_i[22] ),
    .A2(net2978));
 sg13g2_a22oi_1 _08158_ (.Y(_02553_),
    .B1(net2980),
    .B2(\core.gpio.stray_data_i[14] ),
    .A2(net2982),
    .A1(\core.gpio.stray_data_i[6] ));
 sg13g2_o21ai_1 _08159_ (.B1(_02553_),
    .Y(_02554_),
    .A1(net2862),
    .A2(_02552_));
 sg13g2_mux2_1 _08160_ (.A0(net638),
    .A1(_02554_),
    .S(_02526_),
    .X(_00334_));
 sg13g2_nand2b_1 _08161_ (.Y(_02555_),
    .B(net2978),
    .A_N(\core.gpio.stray_data_i[31] ));
 sg13g2_o21ai_1 _08162_ (.B1(_02555_),
    .Y(_02556_),
    .A1(\core.gpio.stray_data_i[23] ),
    .A2(net2978));
 sg13g2_a22oi_1 _08163_ (.Y(_02557_),
    .B1(net2980),
    .B2(\core.gpio.stray_data_i[15] ),
    .A2(net2982),
    .A1(\core.gpio.stray_data_i[7] ));
 sg13g2_o21ai_1 _08164_ (.B1(_02557_),
    .Y(_02558_),
    .A1(net2862),
    .A2(_02556_));
 sg13g2_mux2_1 _08165_ (.A0(net589),
    .A1(_02558_),
    .S(_02526_),
    .X(_00335_));
 sg13g2_nor2_1 _08166_ (.A(net3446),
    .B(net3447),
    .Y(_02559_));
 sg13g2_nor3_2 _08167_ (.A(net3443),
    .B(net3446),
    .C(net3447),
    .Y(_02560_));
 sg13g2_nand2_1 _08168_ (.Y(_02561_),
    .A(_00607_),
    .B(_02560_));
 sg13g2_or4_2 _08169_ (.A(net3448),
    .B(\core.e2m_addr[26] ),
    .C(net3451),
    .D(_02561_),
    .X(_02562_));
 sg13g2_nor3_1 _08170_ (.A(net3448),
    .B(\core.e2m_addr[26] ),
    .C(net3449),
    .Y(_02563_));
 sg13g2_nand2_2 _08171_ (.Y(_02564_),
    .A(_02560_),
    .B(_02563_));
 sg13g2_nor2_2 _08172_ (.A(net3444),
    .B(_02564_),
    .Y(_02565_));
 sg13g2_nand2_1 _08173_ (.Y(_02566_),
    .A(net3451),
    .B(_02565_));
 sg13g2_inv_1 _08174_ (.Y(_02567_),
    .A(_02566_));
 sg13g2_o21ai_1 _08175_ (.B1(_01128_),
    .Y(_02568_),
    .A1(net3440),
    .A2(_02437_));
 sg13g2_nor2b_1 _08176_ (.A(net3451),
    .B_N(net3440),
    .Y(_02569_));
 sg13g2_a221oi_1 _08177_ (.B2(_02565_),
    .C1(_02568_),
    .B1(_02569_),
    .A1(_02562_),
    .Y(_02570_),
    .A2(_02566_));
 sg13g2_a21oi_2 _08178_ (.B1(_01143_),
    .Y(_02571_),
    .A2(_01136_),
    .A1(net3358));
 sg13g2_and2_1 _08179_ (.A(\core.lsu.state[2] ),
    .B(_01125_),
    .X(_02572_));
 sg13g2_nand2_1 _08180_ (.Y(_02573_),
    .A(\core.lsu.state[2] ),
    .B(_01125_));
 sg13g2_nor3_1 _08181_ (.A(\core.lsu.spi.counter[3] ),
    .B(\core.lsu.spi.counter[2] ),
    .C(\core.lsu.spi.counter[4] ),
    .Y(_02574_));
 sg13g2_nor2_1 _08182_ (.A(\core.lsu.spi.counter[1] ),
    .B(\core.lsu.spi.counter[5] ),
    .Y(_02575_));
 sg13g2_nand2_1 _08183_ (.Y(_02576_),
    .A(_02574_),
    .B(_02575_));
 sg13g2_nor2_2 _08184_ (.A(\core.lsu.spi.counter[0] ),
    .B(_02576_),
    .Y(_02577_));
 sg13g2_nor2_1 _08185_ (.A(_00585_),
    .B(_00999_),
    .Y(_02578_));
 sg13g2_nand2_1 _08186_ (.Y(_02579_),
    .A(\core.lsu.spi.state[2] ),
    .B(_00998_));
 sg13g2_nand3_1 _08187_ (.B(_02577_),
    .C(net2975),
    .A(\core.lsu.spi_valid ),
    .Y(_02580_));
 sg13g2_nand2_1 _08188_ (.Y(_02581_),
    .A(net3155),
    .B(_02580_));
 sg13g2_nand2_1 _08189_ (.Y(_02582_),
    .A(\core.work.registers.state[1] ),
    .B(\core.work.registers.state[0] ));
 sg13g2_nand3_1 _08190_ (.B(\core.work.registers.state[0] ),
    .C(_00058_),
    .A(\core.work.registers.state[1] ),
    .Y(_02583_));
 sg13g2_nand2_1 _08191_ (.Y(_02584_),
    .A(_01140_),
    .B(net3151));
 sg13g2_and4_1 _08192_ (.A(_01126_),
    .B(_01140_),
    .C(_02428_),
    .D(net3151),
    .X(_02585_));
 sg13g2_a21oi_1 _08193_ (.A1(_02429_),
    .A2(_02583_),
    .Y(_02586_),
    .B1(_02585_));
 sg13g2_xnor2_1 _08194_ (.Y(_02587_),
    .A(_00056_),
    .B(net3351));
 sg13g2_nor2_1 _08195_ (.A(net3518),
    .B(\core.lsu.write_index[2] ),
    .Y(_02588_));
 sg13g2_nor2b_1 _08196_ (.A(\core.lsu.write_index[2] ),
    .B_N(net3518),
    .Y(_02589_));
 sg13g2_xnor2_1 _08197_ (.Y(_02590_),
    .A(net3523),
    .B(net3517));
 sg13g2_nor4_2 _08198_ (.A(\core.lsu.write_index[2] ),
    .B(_02580_),
    .C(_02587_),
    .Y(_02591_),
    .D(_02590_));
 sg13g2_o21ai_1 _08199_ (.B1(_02586_),
    .Y(_02592_),
    .A1(net3151),
    .A2(_02591_));
 sg13g2_nor2_1 _08200_ (.A(_02571_),
    .B(_02592_),
    .Y(_02593_));
 sg13g2_o21ai_1 _08201_ (.B1(_02593_),
    .Y(_02594_),
    .A1(_01126_),
    .A2(_02570_));
 sg13g2_a21oi_1 _08202_ (.A1(_00059_),
    .A2(_02584_),
    .Y(_02595_),
    .B1(net3201));
 sg13g2_or2_1 _08203_ (.X(_02596_),
    .B(_02584_),
    .A(_02429_));
 sg13g2_nor2_1 _08204_ (.A(_02562_),
    .B(_02596_),
    .Y(_02597_));
 sg13g2_nand2_1 _08205_ (.Y(_02598_),
    .A(net3449),
    .B(_02597_));
 sg13g2_nand2_1 _08206_ (.Y(_02599_),
    .A(_02595_),
    .B(_02598_));
 sg13g2_mux2_1 _08207_ (.A0(_02599_),
    .A1(net736),
    .S(_02594_),
    .X(_00336_));
 sg13g2_o21ai_1 _08208_ (.B1(_02595_),
    .Y(_02600_),
    .A1(_02567_),
    .A2(_02596_));
 sg13g2_mux2_1 _08209_ (.A0(_02600_),
    .A1(net691),
    .S(_02594_),
    .X(_00337_));
 sg13g2_o21ai_1 _08210_ (.B1(_02595_),
    .Y(_02601_),
    .A1(_02566_),
    .A2(_02596_));
 sg13g2_mux2_1 _08211_ (.A0(_02601_),
    .A1(net590),
    .S(_02594_),
    .X(_00338_));
 sg13g2_mux2_1 _08212_ (.A0(net3440),
    .A1(net849),
    .S(net2863),
    .X(_00339_));
 sg13g2_nand2_1 _08213_ (.Y(_02602_),
    .A(net399),
    .B(net2863));
 sg13g2_o21ai_1 _08214_ (.B1(_02602_),
    .Y(_00340_),
    .A1(_00629_),
    .A2(net2863));
 sg13g2_mux2_1 _08215_ (.A0(net438),
    .A1(\core.lsu.is_half ),
    .S(_02494_),
    .X(_00341_));
 sg13g2_nand2_1 _08216_ (.Y(_02603_),
    .A(net3590),
    .B(net3156));
 sg13g2_nor3_1 _08217_ (.A(_00018_),
    .B(_02580_),
    .C(_02603_),
    .Y(_02604_));
 sg13g2_a21oi_1 _08218_ (.A1(_00579_),
    .A2(_02603_),
    .Y(_00342_),
    .B1(_02604_));
 sg13g2_mux2_1 _08219_ (.A0(net840),
    .A1(net3523),
    .S(net2863),
    .X(_00343_));
 sg13g2_o21ai_1 _08220_ (.B1(_02581_),
    .Y(_02605_),
    .A1(_01126_),
    .A2(_01128_));
 sg13g2_inv_1 _08221_ (.Y(_02606_),
    .A(_02605_));
 sg13g2_o21ai_1 _08222_ (.B1(net3589),
    .Y(_02607_),
    .A1(_01125_),
    .A2(_01141_));
 sg13g2_nor3_2 _08223_ (.A(_02571_),
    .B(_02605_),
    .C(_02607_),
    .Y(_02608_));
 sg13g2_or3_1 _08224_ (.A(_02571_),
    .B(_02605_),
    .C(_02607_),
    .X(_02609_));
 sg13g2_nor3_2 _08225_ (.A(net3517),
    .B(net3515),
    .C(\core.lsu.write_index[2] ),
    .Y(_02610_));
 sg13g2_o21ai_1 _08226_ (.B1(_02608_),
    .Y(_02611_),
    .A1(net3152),
    .A2(_02610_));
 sg13g2_nand2_1 _08227_ (.Y(_02612_),
    .A(net725),
    .B(_02611_));
 sg13g2_nor3_1 _08228_ (.A(net3203),
    .B(net3157),
    .C(net3155),
    .Y(_02613_));
 sg13g2_and2_2 _08229_ (.A(net1),
    .B(_02525_),
    .X(_02614_));
 sg13g2_and2_2 _08230_ (.A(net3155),
    .B(_02610_),
    .X(_02615_));
 sg13g2_a22oi_1 _08231_ (.Y(_02616_),
    .B1(_02615_),
    .B2(\core.lsu.spi.buffer[0] ),
    .A2(net3205),
    .A1(\core.fetch.data[0] ));
 sg13g2_inv_1 _08232_ (.Y(_02617_),
    .A(_02616_));
 sg13g2_a221oi_1 _08233_ (.B2(net2981),
    .C1(_02617_),
    .B1(_02614_),
    .A1(net468),
    .Y(_02618_),
    .A2(net2970));
 sg13g2_o21ai_1 _08234_ (.B1(_02612_),
    .Y(_00344_),
    .A1(net2804),
    .A2(_02618_));
 sg13g2_and2_1 _08235_ (.A(net2),
    .B(net3157),
    .X(_02619_));
 sg13g2_nand2_1 _08236_ (.Y(_02620_),
    .A(net2981),
    .B(_02619_));
 sg13g2_a221oi_1 _08237_ (.B2(\core.lsu.spi.buffer[1] ),
    .C1(net2970),
    .B1(_02615_),
    .A1(\core.fetch.data[1] ),
    .Y(_02621_),
    .A2(net3205));
 sg13g2_a221oi_1 _08238_ (.B2(_02621_),
    .C1(net2804),
    .B1(_02620_),
    .A1(_00709_),
    .Y(_02622_),
    .A2(net2970));
 sg13g2_a21o_1 _08239_ (.A2(_02611_),
    .A1(net787),
    .B1(_02622_),
    .X(_00345_));
 sg13g2_nand2_1 _08240_ (.Y(_02623_),
    .A(net696),
    .B(_02611_));
 sg13g2_and2_2 _08241_ (.A(net3),
    .B(net3157),
    .X(_02624_));
 sg13g2_a22oi_1 _08242_ (.Y(_02625_),
    .B1(_02615_),
    .B2(\core.lsu.spi.buffer[2] ),
    .A2(net3205),
    .A1(\core.fetch.data[2] ));
 sg13g2_inv_1 _08243_ (.Y(_02626_),
    .A(_02625_));
 sg13g2_a221oi_1 _08244_ (.B2(_02511_),
    .C1(_02626_),
    .B1(_02624_),
    .A1(net629),
    .Y(_02627_),
    .A2(net2971));
 sg13g2_o21ai_1 _08245_ (.B1(_02623_),
    .Y(_00346_),
    .A1(net2804),
    .A2(_02627_));
 sg13g2_and2_2 _08246_ (.A(net4),
    .B(net3157),
    .X(_02628_));
 sg13g2_nand2_1 _08247_ (.Y(_02629_),
    .A(net2981),
    .B(_02628_));
 sg13g2_a221oi_1 _08248_ (.B2(\core.lsu.spi.buffer[3] ),
    .C1(net2970),
    .B1(_02615_),
    .A1(\core.fetch.data[3] ),
    .Y(_02630_),
    .A2(net3205));
 sg13g2_a221oi_1 _08249_ (.B2(_02630_),
    .C1(net2804),
    .B1(_02629_),
    .A1(_00710_),
    .Y(_02631_),
    .A2(net2970));
 sg13g2_a21o_1 _08250_ (.A2(_02611_),
    .A1(net668),
    .B1(_02631_),
    .X(_00347_));
 sg13g2_and2_2 _08251_ (.A(net5),
    .B(net3157),
    .X(_02632_));
 sg13g2_nand2_1 _08252_ (.Y(_02633_),
    .A(net2981),
    .B(_02632_));
 sg13g2_a221oi_1 _08253_ (.B2(\core.lsu.spi.buffer[4] ),
    .C1(net2970),
    .B1(_02615_),
    .A1(\core.fetch.data[4] ),
    .Y(_02634_),
    .A2(net3205));
 sg13g2_a221oi_1 _08254_ (.B2(_02634_),
    .C1(net2804),
    .B1(_02633_),
    .A1(_00711_),
    .Y(_02635_),
    .A2(net2970));
 sg13g2_a21o_1 _08255_ (.A2(_02611_),
    .A1(net735),
    .B1(_02635_),
    .X(_00348_));
 sg13g2_and2_1 _08256_ (.A(net6),
    .B(net3157),
    .X(_02636_));
 sg13g2_nand2_1 _08257_ (.Y(_02637_),
    .A(net2982),
    .B(_02636_));
 sg13g2_a221oi_1 _08258_ (.B2(\core.lsu.spi.buffer[5] ),
    .C1(net2972),
    .B1(_02615_),
    .A1(\core.fetch.data[5] ),
    .Y(_02638_),
    .A2(net3202));
 sg13g2_a221oi_1 _08259_ (.B2(_02638_),
    .C1(net2802),
    .B1(_02637_),
    .A1(_00712_),
    .Y(_02639_),
    .A2(net2972));
 sg13g2_a21o_1 _08260_ (.A2(_02611_),
    .A1(net687),
    .B1(_02639_),
    .X(_00349_));
 sg13g2_and2_1 _08261_ (.A(net7),
    .B(net3157),
    .X(_02640_));
 sg13g2_o21ai_1 _08262_ (.B1(net3153),
    .Y(_02641_),
    .A1(\core.gpio.stray_data_i[6] ),
    .A2(_02610_));
 sg13g2_a21oi_1 _08263_ (.A1(_00728_),
    .A2(_02610_),
    .Y(_02642_),
    .B1(_02641_));
 sg13g2_a221oi_1 _08264_ (.B2(_02640_),
    .C1(_02642_),
    .B1(net2982),
    .A1(net442),
    .Y(_02643_),
    .A2(net3203));
 sg13g2_a21oi_1 _08265_ (.A1(net517),
    .A2(net2971),
    .Y(_02644_),
    .B1(net2804));
 sg13g2_a22oi_1 _08266_ (.Y(_00350_),
    .B1(_02643_),
    .B2(_02644_),
    .A2(net2804),
    .A1(_00729_));
 sg13g2_and2_1 _08267_ (.A(net8),
    .B(net3157),
    .X(_02645_));
 sg13g2_nand2_1 _08268_ (.Y(_02646_),
    .A(net2982),
    .B(_02645_));
 sg13g2_and2_1 _08269_ (.A(\core.lsu.spi.buffer[7] ),
    .B(net3153),
    .X(_02647_));
 sg13g2_a221oi_1 _08270_ (.B2(_02647_),
    .C1(net2967),
    .B1(_02610_),
    .A1(net455),
    .Y(_02648_),
    .A2(net3202));
 sg13g2_a221oi_1 _08271_ (.B2(_02648_),
    .C1(net2802),
    .B1(_02646_),
    .A1(_00713_),
    .Y(_02649_),
    .A2(net2967));
 sg13g2_a21o_1 _08272_ (.A2(_02611_),
    .A1(net693),
    .B1(_02649_),
    .X(_00351_));
 sg13g2_nand2b_2 _08273_ (.Y(_02650_),
    .B(_02589_),
    .A_N(net3516));
 sg13g2_a22oi_1 _08274_ (.Y(_02651_),
    .B1(net2969),
    .B2(net560),
    .A2(net3204),
    .A1(\core.fetch.data[8] ));
 sg13g2_mux2_1 _08275_ (.A0(\core.lsu.spi.buffer[0] ),
    .A1(\core.gpio.stray_data_i[8] ),
    .S(_02650_),
    .X(_02652_));
 sg13g2_a22oi_1 _08276_ (.Y(_02653_),
    .B1(_02652_),
    .B2(net3156),
    .A2(_02614_),
    .A1(net2979));
 sg13g2_a21oi_1 _08277_ (.A1(_02651_),
    .A2(_02653_),
    .Y(_02654_),
    .B1(net2806));
 sg13g2_a21o_1 _08278_ (.A2(net2803),
    .A1(net733),
    .B1(_02654_),
    .X(_00352_));
 sg13g2_a22oi_1 _08279_ (.Y(_02655_),
    .B1(net2969),
    .B2(\core.e2m_data[9] ),
    .A2(net3204),
    .A1(\core.fetch.data[9] ));
 sg13g2_mux2_1 _08280_ (.A0(\core.lsu.spi.buffer[1] ),
    .A1(\core.gpio.stray_data_i[9] ),
    .S(_02650_),
    .X(_02656_));
 sg13g2_a22oi_1 _08281_ (.Y(_02657_),
    .B1(_02656_),
    .B2(net3156),
    .A2(_02619_),
    .A1(net2979));
 sg13g2_a21oi_1 _08282_ (.A1(_02655_),
    .A2(_02657_),
    .Y(_02658_),
    .B1(net2805));
 sg13g2_a21o_1 _08283_ (.A2(net2804),
    .A1(net726),
    .B1(_02658_),
    .X(_00353_));
 sg13g2_a22oi_1 _08284_ (.Y(_02659_),
    .B1(net2968),
    .B2(net542),
    .A2(net3201),
    .A1(net504));
 sg13g2_mux2_1 _08285_ (.A0(\core.lsu.spi.buffer[2] ),
    .A1(\core.gpio.stray_data_i[10] ),
    .S(_02650_),
    .X(_02660_));
 sg13g2_a22oi_1 _08286_ (.Y(_02661_),
    .B1(_02660_),
    .B2(net3155),
    .A2(_02624_),
    .A1(net2980));
 sg13g2_a21oi_1 _08287_ (.A1(_02659_),
    .A2(_02661_),
    .Y(_02662_),
    .B1(net2802));
 sg13g2_a21o_1 _08288_ (.A2(net2802),
    .A1(net728),
    .B1(_02662_),
    .X(_00354_));
 sg13g2_a22oi_1 _08289_ (.Y(_02663_),
    .B1(net2971),
    .B2(\core.e2m_data[11] ),
    .A2(net3205),
    .A1(\core.fetch.data[11] ));
 sg13g2_mux2_1 _08290_ (.A0(\core.lsu.spi.buffer[3] ),
    .A1(\core.gpio.stray_data_i[11] ),
    .S(_02650_),
    .X(_02664_));
 sg13g2_a22oi_1 _08291_ (.Y(_02665_),
    .B1(_02664_),
    .B2(net3156),
    .A2(_02628_),
    .A1(_02517_));
 sg13g2_a21oi_1 _08292_ (.A1(_02663_),
    .A2(_02665_),
    .Y(_02666_),
    .B1(net2805));
 sg13g2_a21o_1 _08293_ (.A2(net2805),
    .A1(net719),
    .B1(_02666_),
    .X(_00355_));
 sg13g2_a22oi_1 _08294_ (.Y(_02667_),
    .B1(net2969),
    .B2(\core.e2m_data[12] ),
    .A2(net3205),
    .A1(\core.fetch.data[12] ));
 sg13g2_mux2_1 _08295_ (.A0(\core.lsu.spi.buffer[4] ),
    .A1(\core.gpio.stray_data_i[12] ),
    .S(_02650_),
    .X(_02668_));
 sg13g2_a22oi_1 _08296_ (.Y(_02669_),
    .B1(_02668_),
    .B2(net3156),
    .A2(_02632_),
    .A1(_02517_));
 sg13g2_a21oi_1 _08297_ (.A1(_02667_),
    .A2(_02669_),
    .Y(_02670_),
    .B1(net2803));
 sg13g2_a21o_1 _08298_ (.A2(net2805),
    .A1(net713),
    .B1(_02670_),
    .X(_00356_));
 sg13g2_a22oi_1 _08299_ (.Y(_02671_),
    .B1(net2968),
    .B2(net604),
    .A2(net3201),
    .A1(net397));
 sg13g2_mux2_1 _08300_ (.A0(\core.lsu.spi.buffer[5] ),
    .A1(\core.gpio.stray_data_i[13] ),
    .S(_02650_),
    .X(_02672_));
 sg13g2_a22oi_1 _08301_ (.Y(_02673_),
    .B1(_02672_),
    .B2(net3154),
    .A2(_02636_),
    .A1(net2980));
 sg13g2_a21oi_1 _08302_ (.A1(_02671_),
    .A2(_02673_),
    .Y(_02674_),
    .B1(net2800));
 sg13g2_a21o_1 _08303_ (.A2(net2799),
    .A1(net753),
    .B1(_02674_),
    .X(_00357_));
 sg13g2_a22oi_1 _08304_ (.Y(_02675_),
    .B1(net2968),
    .B2(\core.e2m_data[14] ),
    .A2(net3201),
    .A1(\core.fetch.data[14] ));
 sg13g2_mux2_1 _08305_ (.A0(\core.lsu.spi.buffer[6] ),
    .A1(\core.gpio.stray_data_i[14] ),
    .S(_02650_),
    .X(_02676_));
 sg13g2_a22oi_1 _08306_ (.Y(_02677_),
    .B1(_02676_),
    .B2(net3153),
    .A2(_02640_),
    .A1(net2980));
 sg13g2_a21oi_1 _08307_ (.A1(_02675_),
    .A2(_02677_),
    .Y(_02678_),
    .B1(net2802));
 sg13g2_a21o_1 _08308_ (.A2(net2802),
    .A1(net723),
    .B1(_02678_),
    .X(_00358_));
 sg13g2_a22oi_1 _08309_ (.Y(_02679_),
    .B1(net2968),
    .B2(net617),
    .A2(net3201),
    .A1(net522));
 sg13g2_mux2_1 _08310_ (.A0(\core.lsu.spi.buffer[7] ),
    .A1(\core.gpio.stray_data_i[15] ),
    .S(_02650_),
    .X(_02680_));
 sg13g2_a22oi_1 _08311_ (.Y(_02681_),
    .B1(_02680_),
    .B2(net3153),
    .A2(_02645_),
    .A1(net2980));
 sg13g2_a21oi_1 _08312_ (.A1(_02679_),
    .A2(_02681_),
    .Y(_02682_),
    .B1(net2801));
 sg13g2_a21o_1 _08313_ (.A2(net2798),
    .A1(net700),
    .B1(_02682_),
    .X(_00359_));
 sg13g2_and2_2 _08314_ (.A(net3515),
    .B(_02588_),
    .X(_02683_));
 sg13g2_nand2_2 _08315_ (.Y(_02684_),
    .A(net3515),
    .B(_02588_));
 sg13g2_o21ai_1 _08316_ (.B1(_02608_),
    .Y(_02685_),
    .A1(net3152),
    .A2(_02683_));
 sg13g2_nand3_1 _08317_ (.B(_02520_),
    .C(_02614_),
    .A(_02515_),
    .Y(_02686_));
 sg13g2_nor3_1 _08318_ (.A(_00133_),
    .B(net3152),
    .C(_02684_),
    .Y(_02687_));
 sg13g2_a221oi_1 _08319_ (.B2(\core.e2m_data[16] ),
    .C1(_02687_),
    .B1(net2969),
    .A1(\core.fetch.data[16] ),
    .Y(_02688_),
    .A2(net3204));
 sg13g2_a21oi_1 _08320_ (.A1(_02686_),
    .A2(_02688_),
    .Y(_02689_),
    .B1(net2803));
 sg13g2_a21o_1 _08321_ (.A2(_02685_),
    .A1(net651),
    .B1(_02689_),
    .X(_00360_));
 sg13g2_nor2_1 _08322_ (.A(\core.gpio.stray_data_i[17] ),
    .B(_02683_),
    .Y(_02690_));
 sg13g2_a22oi_1 _08323_ (.Y(_02691_),
    .B1(net2969),
    .B2(net489),
    .A2(net3204),
    .A1(\core.fetch.data[17] ));
 sg13g2_a21oi_1 _08324_ (.A1(_00134_),
    .A2(_02683_),
    .Y(_02692_),
    .B1(_02690_));
 sg13g2_a22oi_1 _08325_ (.Y(_02693_),
    .B1(_02692_),
    .B2(net3154),
    .A2(_02619_),
    .A1(_02522_));
 sg13g2_a21oi_1 _08326_ (.A1(_02691_),
    .A2(_02693_),
    .Y(_02694_),
    .B1(net2806));
 sg13g2_a21o_1 _08327_ (.A2(net2803),
    .A1(net760),
    .B1(_02694_),
    .X(_00361_));
 sg13g2_nand3_1 _08328_ (.B(_02520_),
    .C(_02624_),
    .A(_02515_),
    .Y(_02695_));
 sg13g2_nor3_1 _08329_ (.A(_00135_),
    .B(net3151),
    .C(_02684_),
    .Y(_02696_));
 sg13g2_a221oi_1 _08330_ (.B2(net475),
    .C1(_02696_),
    .B1(net2969),
    .A1(\core.fetch.data[18] ),
    .Y(_02697_),
    .A2(net3204));
 sg13g2_a21oi_1 _08331_ (.A1(_02695_),
    .A2(_02697_),
    .Y(_02698_),
    .B1(net2803));
 sg13g2_a21o_1 _08332_ (.A2(_02685_),
    .A1(net649),
    .B1(_02698_),
    .X(_00362_));
 sg13g2_nand3_1 _08333_ (.B(_02520_),
    .C(_02628_),
    .A(_02515_),
    .Y(_02699_));
 sg13g2_nor3_1 _08334_ (.A(_00136_),
    .B(net3151),
    .C(_02684_),
    .Y(_02700_));
 sg13g2_a221oi_1 _08335_ (.B2(net467),
    .C1(_02700_),
    .B1(net2969),
    .A1(\core.fetch.data[19] ),
    .Y(_02701_),
    .A2(net3204));
 sg13g2_a21oi_1 _08336_ (.A1(_02699_),
    .A2(_02701_),
    .Y(_02702_),
    .B1(net2803));
 sg13g2_a21o_1 _08337_ (.A2(_02685_),
    .A1(net673),
    .B1(_02702_),
    .X(_00363_));
 sg13g2_nand3_1 _08338_ (.B(_02520_),
    .C(_02632_),
    .A(_02515_),
    .Y(_02703_));
 sg13g2_nor3_1 _08339_ (.A(_00137_),
    .B(net3151),
    .C(_02684_),
    .Y(_02704_));
 sg13g2_a221oi_1 _08340_ (.B2(net488),
    .C1(_02704_),
    .B1(net2969),
    .A1(\core.fetch.data[20] ),
    .Y(_02705_),
    .A2(net3204));
 sg13g2_nand2_1 _08341_ (.Y(_02706_),
    .A(_02703_),
    .B(_02705_));
 sg13g2_a22oi_1 _08342_ (.Y(_02707_),
    .B1(_02706_),
    .B2(_02608_),
    .A2(_02685_),
    .A1(net625));
 sg13g2_inv_1 _08343_ (.Y(_00364_),
    .A(_02707_));
 sg13g2_nor2_1 _08344_ (.A(\core.gpio.stray_data_i[21] ),
    .B(_02683_),
    .Y(_02708_));
 sg13g2_a22oi_1 _08345_ (.Y(_02709_),
    .B1(net2968),
    .B2(net491),
    .A2(net3203),
    .A1(\core.fetch.data[21] ));
 sg13g2_a21oi_1 _08346_ (.A1(_00138_),
    .A2(_02683_),
    .Y(_02710_),
    .B1(_02708_));
 sg13g2_a22oi_1 _08347_ (.Y(_02711_),
    .B1(_02710_),
    .B2(net3154),
    .A2(_02636_),
    .A1(_02522_));
 sg13g2_a21oi_1 _08348_ (.A1(_02709_),
    .A2(_02711_),
    .Y(_02712_),
    .B1(net2807));
 sg13g2_a21o_1 _08349_ (.A2(net2800),
    .A1(net747),
    .B1(_02712_),
    .X(_00365_));
 sg13g2_nor2_1 _08350_ (.A(\core.gpio.stray_data_i[22] ),
    .B(_02683_),
    .Y(_02713_));
 sg13g2_a22oi_1 _08351_ (.Y(_02714_),
    .B1(net2968),
    .B2(net483),
    .A2(net3201),
    .A1(\core.fetch.data[22] ));
 sg13g2_a21oi_1 _08352_ (.A1(_00139_),
    .A2(_02683_),
    .Y(_02715_),
    .B1(_02713_));
 sg13g2_a22oi_1 _08353_ (.Y(_02716_),
    .B1(_02715_),
    .B2(net3153),
    .A2(_02640_),
    .A1(_02522_));
 sg13g2_a21oi_1 _08354_ (.A1(_02714_),
    .A2(_02716_),
    .Y(_02717_),
    .B1(net2799));
 sg13g2_a21o_1 _08355_ (.A2(net2798),
    .A1(net754),
    .B1(_02717_),
    .X(_00366_));
 sg13g2_nand3_1 _08356_ (.B(_02520_),
    .C(_02645_),
    .A(_02515_),
    .Y(_02718_));
 sg13g2_nor3_2 _08357_ (.A(_00140_),
    .B(net3151),
    .C(_02684_),
    .Y(_02719_));
 sg13g2_a221oi_1 _08358_ (.B2(\core.e2m_data[23] ),
    .C1(_02719_),
    .B1(net2968),
    .A1(\core.fetch.data[23] ),
    .Y(_02720_),
    .A2(net3201));
 sg13g2_a21oi_1 _08359_ (.A1(_02718_),
    .A2(_02720_),
    .Y(_02721_),
    .B1(net2802));
 sg13g2_a21o_1 _08360_ (.A2(_02685_),
    .A1(net675),
    .B1(_02721_),
    .X(_00367_));
 sg13g2_nand2_1 _08361_ (.Y(_02722_),
    .A(net3518),
    .B(net3515));
 sg13g2_nor2_1 _08362_ (.A(\core.lsu.write_index[2] ),
    .B(_02722_),
    .Y(_02723_));
 sg13g2_a22oi_1 _08363_ (.Y(_02724_),
    .B1(net2970),
    .B2(net413),
    .A2(net3204),
    .A1(net464));
 sg13g2_mux2_1 _08364_ (.A0(\core.gpio.stray_data_i[24] ),
    .A1(\core.lsu.spi.buffer[0] ),
    .S(net3146),
    .X(_02725_));
 sg13g2_a22oi_1 _08365_ (.Y(_02726_),
    .B1(_02725_),
    .B2(net3156),
    .A2(_02614_),
    .A1(_02523_));
 sg13g2_a21oi_1 _08366_ (.A1(_02724_),
    .A2(_02726_),
    .Y(_02727_),
    .B1(net2803));
 sg13g2_a21o_1 _08367_ (.A2(net2803),
    .A1(net614),
    .B1(_02727_),
    .X(_00368_));
 sg13g2_a22oi_1 _08368_ (.Y(_02728_),
    .B1(net2968),
    .B2(\core.e2m_data[25] ),
    .A2(net3201),
    .A1(\core.fetch.data[25] ));
 sg13g2_o21ai_1 _08369_ (.B1(net3156),
    .Y(_02729_),
    .A1(\core.gpio.stray_data_i[25] ),
    .A2(net3145));
 sg13g2_a21oi_1 _08370_ (.A1(_00724_),
    .A2(net3146),
    .Y(_02730_),
    .B1(_02729_));
 sg13g2_a21oi_1 _08371_ (.A1(net2976),
    .A2(_02619_),
    .Y(_02731_),
    .B1(_02730_));
 sg13g2_a21oi_1 _08372_ (.A1(_02728_),
    .A2(_02731_),
    .Y(_02732_),
    .B1(net2802));
 sg13g2_a21o_1 _08373_ (.A2(net2806),
    .A1(net786),
    .B1(_02732_),
    .X(_00369_));
 sg13g2_a22oi_1 _08374_ (.Y(_02733_),
    .B1(net2967),
    .B2(net493),
    .A2(net3202),
    .A1(net404));
 sg13g2_mux2_1 _08375_ (.A0(\core.gpio.stray_data_i[26] ),
    .A1(\core.lsu.spi.buffer[2] ),
    .S(net3145),
    .X(_02734_));
 sg13g2_a22oi_1 _08376_ (.Y(_02735_),
    .B1(_02734_),
    .B2(net3155),
    .A2(_02624_),
    .A1(net2976));
 sg13g2_a21oi_1 _08377_ (.A1(_02733_),
    .A2(_02735_),
    .Y(_02736_),
    .B1(net2801));
 sg13g2_a21o_1 _08378_ (.A2(net2801),
    .A1(net701),
    .B1(_02736_),
    .X(_00370_));
 sg13g2_a22oi_1 _08379_ (.Y(_02737_),
    .B1(net2967),
    .B2(net529),
    .A2(net3202),
    .A1(\core.fetch.data[27] ));
 sg13g2_o21ai_1 _08380_ (.B1(net3154),
    .Y(_02738_),
    .A1(\core.gpio.stray_data_i[27] ),
    .A2(net3146));
 sg13g2_a21oi_1 _08381_ (.A1(_00725_),
    .A2(net3146),
    .Y(_02739_),
    .B1(_02738_));
 sg13g2_a21oi_1 _08382_ (.A1(net2976),
    .A2(_02628_),
    .Y(_02740_),
    .B1(_02739_));
 sg13g2_a21oi_1 _08383_ (.A1(_02737_),
    .A2(_02740_),
    .Y(_02741_),
    .B1(net2798));
 sg13g2_a21o_1 _08384_ (.A2(net2798),
    .A1(net767),
    .B1(_02741_),
    .X(_00371_));
 sg13g2_a22oi_1 _08385_ (.Y(_02742_),
    .B1(net2967),
    .B2(net662),
    .A2(net3202),
    .A1(net367));
 sg13g2_o21ai_1 _08386_ (.B1(net3154),
    .Y(_02743_),
    .A1(\core.gpio.stray_data_i[28] ),
    .A2(net3145));
 sg13g2_a21oi_1 _08387_ (.A1(_00726_),
    .A2(net3146),
    .Y(_02744_),
    .B1(_02743_));
 sg13g2_a21oi_1 _08388_ (.A1(net2976),
    .A2(_02632_),
    .Y(_02745_),
    .B1(_02744_));
 sg13g2_a21oi_1 _08389_ (.A1(_02742_),
    .A2(_02745_),
    .Y(_02746_),
    .B1(net2798));
 sg13g2_a21o_1 _08390_ (.A2(net2799),
    .A1(net802),
    .B1(_02746_),
    .X(_00372_));
 sg13g2_a22oi_1 _08391_ (.Y(_02747_),
    .B1(net2967),
    .B2(net512),
    .A2(net3202),
    .A1(net388));
 sg13g2_o21ai_1 _08392_ (.B1(net3153),
    .Y(_02748_),
    .A1(\core.gpio.stray_data_i[29] ),
    .A2(net3145));
 sg13g2_a21oi_1 _08393_ (.A1(_00727_),
    .A2(net3145),
    .Y(_02749_),
    .B1(_02748_));
 sg13g2_a21oi_1 _08394_ (.A1(net2976),
    .A2(_02636_),
    .Y(_02750_),
    .B1(_02749_));
 sg13g2_a21oi_1 _08395_ (.A1(_02747_),
    .A2(_02750_),
    .Y(_02751_),
    .B1(net2799));
 sg13g2_a21o_1 _08396_ (.A2(net2799),
    .A1(net766),
    .B1(_02751_),
    .X(_00373_));
 sg13g2_a22oi_1 _08397_ (.Y(_02752_),
    .B1(net2967),
    .B2(net592),
    .A2(net3202),
    .A1(net423));
 sg13g2_o21ai_1 _08398_ (.B1(net3153),
    .Y(_02753_),
    .A1(\core.gpio.stray_data_i[30] ),
    .A2(net3145));
 sg13g2_a21oi_1 _08399_ (.A1(_00728_),
    .A2(net3145),
    .Y(_02754_),
    .B1(_02753_));
 sg13g2_a21oi_1 _08400_ (.A1(net2976),
    .A2(_02640_),
    .Y(_02755_),
    .B1(_02754_));
 sg13g2_a21oi_1 _08401_ (.A1(_02752_),
    .A2(_02755_),
    .Y(_02756_),
    .B1(net2798));
 sg13g2_a21o_1 _08402_ (.A2(net2799),
    .A1(net768),
    .B1(_02756_),
    .X(_00374_));
 sg13g2_a22oi_1 _08403_ (.Y(_02757_),
    .B1(net2967),
    .B2(\core.e2m_data[31] ),
    .A2(net3202),
    .A1(net416));
 sg13g2_mux2_1 _08404_ (.A0(\core.gpio.stray_data_i[31] ),
    .A1(\core.lsu.spi.buffer[7] ),
    .S(net3145),
    .X(_02758_));
 sg13g2_a22oi_1 _08405_ (.Y(_02759_),
    .B1(_02758_),
    .B2(net3153),
    .A2(_02645_),
    .A1(net2976));
 sg13g2_a21oi_1 _08406_ (.A1(_02757_),
    .A2(_02759_),
    .Y(_02760_),
    .B1(net2798));
 sg13g2_a21o_1 _08407_ (.A2(net2798),
    .A1(net667),
    .B1(_02760_),
    .X(_00375_));
 sg13g2_mux2_1 _08408_ (.A0(net541),
    .A1(net559),
    .S(net2863),
    .X(_00376_));
 sg13g2_mux2_1 _08409_ (.A0(net562),
    .A1(net572),
    .S(net2863),
    .X(_00377_));
 sg13g2_mux2_1 _08410_ (.A0(net392),
    .A1(\core.lsu.dreg[2] ),
    .S(net2863),
    .X(_00378_));
 sg13g2_mux2_1 _08411_ (.A0(net414),
    .A1(\core.lsu.dreg[3] ),
    .S(net2863),
    .X(_00379_));
 sg13g2_nand2_1 _08412_ (.Y(_02761_),
    .A(\core.lsu.spi.cs ),
    .B(net359));
 sg13g2_nand2_1 _08413_ (.Y(_02762_),
    .A(net3522),
    .B(_00666_));
 sg13g2_o21ai_1 _08414_ (.B1(_02762_),
    .Y(_00380_),
    .A1(_02577_),
    .A2(net360));
 sg13g2_and2_2 _08415_ (.A(net3592),
    .B(\core.lsu.spi.cs ),
    .X(_02763_));
 sg13g2_nand2_1 _08416_ (.Y(_02764_),
    .A(net3593),
    .B(\core.lsu.spi.cs ));
 sg13g2_nor3_1 _08417_ (.A(net3521),
    .B(_02577_),
    .C(net3293),
    .Y(_02765_));
 sg13g2_mux2_1 _08418_ (.A0(net435),
    .A1(net10),
    .S(_02765_),
    .X(_00381_));
 sg13g2_or2_1 _08419_ (.X(_00382_),
    .B(_01002_),
    .A(net461));
 sg13g2_nor2b_1 _08420_ (.A(net3522),
    .B_N(\core.lsu.spi.buffer[0] ),
    .Y(_02766_));
 sg13g2_a21oi_2 _08421_ (.B1(_02766_),
    .Y(_02767_),
    .A2(\core.lsu.spi.cache_bit ),
    .A1(net3522));
 sg13g2_nand2_1 _08422_ (.Y(_02768_),
    .A(_01017_),
    .B(_01022_));
 sg13g2_xor2_1 _08423_ (.B(_01055_),
    .A(_00085_),
    .X(_02769_));
 sg13g2_nand4_1 _08424_ (.B(_01108_),
    .C(_01110_),
    .A(_01057_),
    .Y(_02770_),
    .D(_02769_));
 sg13g2_nor4_1 _08425_ (.A(_01048_),
    .B(_01060_),
    .C(_01106_),
    .D(_02770_),
    .Y(_02771_));
 sg13g2_nand3_1 _08426_ (.B(_00084_),
    .C(_00998_),
    .A(\core.lsu.spi_valid ),
    .Y(_02772_));
 sg13g2_mux4_1 _08427_ (.S0(net3519),
    .A0(\core.gpio.stray_data_i[0] ),
    .A1(\core.gpio.stray_data_i[8] ),
    .A2(\core.gpio.stray_data_i[16] ),
    .A3(\core.gpio.stray_data_i[24] ),
    .S1(net3516),
    .X(_02773_));
 sg13g2_nand2_2 _08428_ (.Y(_02774_),
    .A(net3514),
    .B(_02773_));
 sg13g2_or2_1 _08429_ (.X(_02775_),
    .B(_02768_),
    .A(_01101_));
 sg13g2_nand3_1 _08430_ (.B(_01103_),
    .C(_02771_),
    .A(_01072_),
    .Y(_02776_));
 sg13g2_nor4_1 _08431_ (.A(_01032_),
    .B(_01038_),
    .C(_02775_),
    .D(_02776_),
    .Y(_02777_));
 sg13g2_a21oi_1 _08432_ (.A1(_02774_),
    .A2(net2768),
    .Y(_02778_),
    .B1(_02772_));
 sg13g2_nor2_2 _08433_ (.A(_01124_),
    .B(net2768),
    .Y(_02779_));
 sg13g2_a22oi_1 _08434_ (.Y(_02780_),
    .B1(_02767_),
    .B2(_02779_),
    .A2(_01124_),
    .A1(\core.gpio.stray_wr_i ));
 sg13g2_nand2_1 _08435_ (.Y(_02781_),
    .A(_02778_),
    .B(_02780_));
 sg13g2_nand3_1 _08436_ (.B(\core.lsu.spi.state[0] ),
    .C(_00585_),
    .A(\core.lsu.spi.state[1] ),
    .Y(_02782_));
 sg13g2_inv_1 _08437_ (.Y(_02783_),
    .A(net3144));
 sg13g2_nor2_1 _08438_ (.A(\core.lsu.spi.state[1] ),
    .B(_00584_),
    .Y(_02784_));
 sg13g2_nand2_1 _08439_ (.Y(_02785_),
    .A(_00583_),
    .B(\core.lsu.spi.state[0] ));
 sg13g2_nor2_2 _08440_ (.A(\core.lsu.spi.state[2] ),
    .B(_02785_),
    .Y(_02786_));
 sg13g2_nand2_2 _08441_ (.Y(_02787_),
    .A(_00585_),
    .B(_02784_));
 sg13g2_and3_2 _08442_ (.X(_02788_),
    .A(\core.lsu.spi.state[1] ),
    .B(_00584_),
    .C(_00084_));
 sg13g2_nand3_1 _08443_ (.B(_00584_),
    .C(_00084_),
    .A(\core.lsu.spi.state[1] ),
    .Y(_02789_));
 sg13g2_o21ai_1 _08444_ (.B1(_02789_),
    .Y(_02790_),
    .A1(_00584_),
    .A2(\core.lsu.spi.state[2] ));
 sg13g2_nor2b_2 _08445_ (.A(_02790_),
    .B_N(_01000_),
    .Y(_02791_));
 sg13g2_nand2b_1 _08446_ (.Y(_02792_),
    .B(\core.lsu.spi.counter[0] ),
    .A_N(net3522));
 sg13g2_nand3_1 _08447_ (.B(_02575_),
    .C(_02792_),
    .A(_02574_),
    .Y(_02793_));
 sg13g2_nor2_1 _08448_ (.A(_02774_),
    .B(_02782_),
    .Y(_02794_));
 sg13g2_nand2_2 _08449_ (.Y(_02795_),
    .A(_02790_),
    .B(net3143));
 sg13g2_nor2_1 _08450_ (.A(_00095_),
    .B(_02787_),
    .Y(_02796_));
 sg13g2_nor2_1 _08451_ (.A(_00085_),
    .B(_02789_),
    .Y(_02797_));
 sg13g2_nor2_1 _08452_ (.A(\core.lsu.spi_valid ),
    .B(_01000_),
    .Y(_02798_));
 sg13g2_nand3_1 _08453_ (.B(_00084_),
    .C(_00998_),
    .A(_00579_),
    .Y(_02799_));
 sg13g2_nor2_1 _08454_ (.A(_02767_),
    .B(_02799_),
    .Y(_02800_));
 sg13g2_nor3_1 _08455_ (.A(_02794_),
    .B(_02796_),
    .C(_02797_),
    .Y(_02801_));
 sg13g2_a22oi_1 _08456_ (.Y(_02802_),
    .B1(_02795_),
    .B2(_02801_),
    .A2(net3143),
    .A1(_02767_));
 sg13g2_nor2_2 _08457_ (.A(_02791_),
    .B(_02798_),
    .Y(_02803_));
 sg13g2_nor3_1 _08458_ (.A(_02791_),
    .B(_02800_),
    .C(_02802_),
    .Y(_02804_));
 sg13g2_a221oi_1 _08459_ (.B2(_02781_),
    .C1(net3293),
    .B1(_02804_),
    .A1(_02767_),
    .Y(_02805_),
    .A2(_02791_));
 sg13g2_a21o_1 _08460_ (.A2(net3294),
    .A1(net729),
    .B1(_02805_),
    .X(_00383_));
 sg13g2_mux2_1 _08461_ (.A0(_00134_),
    .A1(_00133_),
    .S(\core.lsu.spi.sck ),
    .X(_02806_));
 sg13g2_mux4_1 _08462_ (.S0(net3519),
    .A0(\core.gpio.stray_data_i[1] ),
    .A1(\core.gpio.stray_data_i[9] ),
    .A2(\core.gpio.stray_data_i[17] ),
    .A3(\core.gpio.stray_data_i[25] ),
    .S1(net3516),
    .X(_02807_));
 sg13g2_nand2_1 _08463_ (.Y(_02808_),
    .A(net3514),
    .B(_02807_));
 sg13g2_a221oi_1 _08464_ (.B2(net2768),
    .C1(_02772_),
    .B1(_02808_),
    .A1(_02779_),
    .Y(_02809_),
    .A2(_02806_));
 sg13g2_o21ai_1 _08465_ (.B1(_02763_),
    .Y(_02810_),
    .A1(_02803_),
    .A2(_02806_));
 sg13g2_or2_1 _08466_ (.X(_02811_),
    .B(_02808_),
    .A(net3144));
 sg13g2_o21ai_1 _08467_ (.B1(_02795_),
    .Y(_02812_),
    .A1(_00094_),
    .A2(_02787_));
 sg13g2_a21oi_1 _08468_ (.A1(\core.lsu.spi.addr[1] ),
    .A2(_02788_),
    .Y(_02813_),
    .B1(_02812_));
 sg13g2_a22oi_1 _08469_ (.Y(_02814_),
    .B1(_02811_),
    .B2(_02813_),
    .A2(_02806_),
    .A1(net3142));
 sg13g2_nor3_1 _08470_ (.A(_02809_),
    .B(_02810_),
    .C(_02814_),
    .Y(_02815_));
 sg13g2_a21oi_1 _08471_ (.A1(_00724_),
    .A2(net3293),
    .Y(_00384_),
    .B1(_02815_));
 sg13g2_mux4_1 _08472_ (.S0(net3518),
    .A0(\core.gpio.stray_data_i[2] ),
    .A1(\core.gpio.stray_data_i[10] ),
    .A2(\core.gpio.stray_data_i[18] ),
    .A3(\core.gpio.stray_data_i[26] ),
    .S1(net3516),
    .X(_02816_));
 sg13g2_and2_1 _08473_ (.A(net3514),
    .B(_02816_),
    .X(_02817_));
 sg13g2_mux2_1 _08474_ (.A0(_00135_),
    .A1(_00134_),
    .S(\core.lsu.spi.sck ),
    .X(_02818_));
 sg13g2_inv_1 _08475_ (.Y(_02819_),
    .A(_02818_));
 sg13g2_a22oi_1 _08476_ (.Y(_02820_),
    .B1(_02819_),
    .B2(_02779_),
    .A2(_02817_),
    .A1(net2768));
 sg13g2_o21ai_1 _08477_ (.B1(_02795_),
    .Y(_02821_),
    .A1(_00086_),
    .A2(_02789_));
 sg13g2_a221oi_1 _08478_ (.B2(_02783_),
    .C1(_02821_),
    .B1(_02817_),
    .A1(_00674_),
    .Y(_02822_),
    .A2(_02786_));
 sg13g2_a21oi_1 _08479_ (.A1(net3143),
    .A2(_02818_),
    .Y(_02823_),
    .B1(_02822_));
 sg13g2_nor2_1 _08480_ (.A(_02799_),
    .B(_02818_),
    .Y(_02824_));
 sg13g2_nor3_1 _08481_ (.A(_02791_),
    .B(_02823_),
    .C(_02824_),
    .Y(_02825_));
 sg13g2_o21ai_1 _08482_ (.B1(_02825_),
    .Y(_02826_),
    .A1(_02772_),
    .A2(_02820_));
 sg13g2_a21oi_1 _08483_ (.A1(_02791_),
    .A2(_02818_),
    .Y(_02827_),
    .B1(net3294));
 sg13g2_a22oi_1 _08484_ (.Y(_02828_),
    .B1(_02826_),
    .B2(_02827_),
    .A2(net3294),
    .A1(net641));
 sg13g2_inv_1 _08485_ (.Y(_00385_),
    .A(_02828_));
 sg13g2_nor2_2 _08486_ (.A(_01124_),
    .B(_02772_),
    .Y(_02829_));
 sg13g2_inv_1 _08487_ (.Y(_02830_),
    .A(_02829_));
 sg13g2_mux4_1 _08488_ (.S0(net3519),
    .A0(\core.gpio.stray_data_i[3] ),
    .A1(\core.gpio.stray_data_i[11] ),
    .A2(\core.gpio.stray_data_i[19] ),
    .A3(\core.gpio.stray_data_i[27] ),
    .S1(net3516),
    .X(_02831_));
 sg13g2_nand2_1 _08489_ (.Y(_02832_),
    .A(net3514),
    .B(_02831_));
 sg13g2_mux2_1 _08490_ (.A0(_00136_),
    .A1(_00135_),
    .S(net3522),
    .X(_02833_));
 sg13g2_nand2b_1 _08491_ (.Y(_02834_),
    .B(_02833_),
    .A_N(net2768));
 sg13g2_nand2_1 _08492_ (.Y(_02835_),
    .A(net2767),
    .B(_02832_));
 sg13g2_nand3_1 _08493_ (.B(_02834_),
    .C(_02835_),
    .A(_02829_),
    .Y(_02836_));
 sg13g2_or2_1 _08494_ (.X(_02837_),
    .B(_02832_),
    .A(net3144));
 sg13g2_a22oi_1 _08495_ (.Y(_02838_),
    .B1(_02788_),
    .B2(\core.lsu.spi.addr[3] ),
    .A2(_02786_),
    .A1(\core.lsu.spi.addr[11] ));
 sg13g2_a21oi_1 _08496_ (.A1(_02837_),
    .A2(_02838_),
    .Y(_02839_),
    .B1(net3142));
 sg13g2_a21oi_1 _08497_ (.A1(_02795_),
    .A2(_02803_),
    .Y(_02840_),
    .B1(_02833_));
 sg13g2_nor3_1 _08498_ (.A(net3294),
    .B(_02839_),
    .C(_02840_),
    .Y(_02841_));
 sg13g2_a22oi_1 _08499_ (.Y(_00386_),
    .B1(_02836_),
    .B2(_02841_),
    .A2(net3293),
    .A1(_00725_));
 sg13g2_mux4_1 _08500_ (.S0(net3519),
    .A0(\core.gpio.stray_data_i[4] ),
    .A1(\core.gpio.stray_data_i[12] ),
    .A2(\core.gpio.stray_data_i[20] ),
    .A3(\core.gpio.stray_data_i[28] ),
    .S1(net3516),
    .X(_02842_));
 sg13g2_nand2_2 _08501_ (.Y(_02843_),
    .A(net3514),
    .B(_02842_));
 sg13g2_mux2_1 _08502_ (.A0(_00137_),
    .A1(_00136_),
    .S(net3521),
    .X(_02844_));
 sg13g2_nand2b_1 _08503_ (.Y(_02845_),
    .B(_02844_),
    .A_N(net2767));
 sg13g2_nand2_1 _08504_ (.Y(_02846_),
    .A(net2767),
    .B(_02843_));
 sg13g2_nand3_1 _08505_ (.B(_02845_),
    .C(_02846_),
    .A(_02829_),
    .Y(_02847_));
 sg13g2_o21ai_1 _08506_ (.B1(_02763_),
    .Y(_02848_),
    .A1(_02803_),
    .A2(_02844_));
 sg13g2_nor2_1 _08507_ (.A(_02782_),
    .B(_02843_),
    .Y(_02849_));
 sg13g2_nor2_1 _08508_ (.A(_00092_),
    .B(_02787_),
    .Y(_02850_));
 sg13g2_nor2_1 _08509_ (.A(_00089_),
    .B(_02789_),
    .Y(_02851_));
 sg13g2_nor3_1 _08510_ (.A(_02849_),
    .B(_02850_),
    .C(_02851_),
    .Y(_02852_));
 sg13g2_a22oi_1 _08511_ (.Y(_02853_),
    .B1(_02852_),
    .B2(_02795_),
    .A2(_02844_),
    .A1(net3142));
 sg13g2_nor2_1 _08512_ (.A(_02848_),
    .B(_02853_),
    .Y(_02854_));
 sg13g2_a22oi_1 _08513_ (.Y(_00387_),
    .B1(_02847_),
    .B2(_02854_),
    .A2(net3293),
    .A1(_00726_));
 sg13g2_mux4_1 _08514_ (.S0(net3517),
    .A0(\core.gpio.stray_data_i[5] ),
    .A1(\core.gpio.stray_data_i[13] ),
    .A2(\core.gpio.stray_data_i[21] ),
    .A3(\core.gpio.stray_data_i[29] ),
    .S1(net3515),
    .X(_02855_));
 sg13g2_nand2_1 _08515_ (.Y(_02856_),
    .A(_00057_),
    .B(_02855_));
 sg13g2_mux2_1 _08516_ (.A0(_00138_),
    .A1(_00137_),
    .S(net3521),
    .X(_02857_));
 sg13g2_nand2b_1 _08517_ (.Y(_02858_),
    .B(_02857_),
    .A_N(net2767));
 sg13g2_nand2_1 _08518_ (.Y(_02859_),
    .A(net2767),
    .B(_02856_));
 sg13g2_nand3_1 _08519_ (.B(_02858_),
    .C(_02859_),
    .A(_02829_),
    .Y(_02860_));
 sg13g2_o21ai_1 _08520_ (.B1(_02763_),
    .Y(_02861_),
    .A1(_02803_),
    .A2(_02857_));
 sg13g2_nor2_1 _08521_ (.A(net3144),
    .B(_02856_),
    .Y(_02862_));
 sg13g2_a221oi_1 _08522_ (.B2(_00668_),
    .C1(_02862_),
    .B1(_02788_),
    .A1(\core.lsu.spi.addr[13] ),
    .Y(_02863_),
    .A2(_02786_));
 sg13g2_a22oi_1 _08523_ (.Y(_02864_),
    .B1(_02863_),
    .B2(_02795_),
    .A2(_02857_),
    .A1(net3142));
 sg13g2_nor2_1 _08524_ (.A(_02861_),
    .B(_02864_),
    .Y(_02865_));
 sg13g2_a22oi_1 _08525_ (.Y(_00388_),
    .B1(_02860_),
    .B2(_02865_),
    .A2(net3293),
    .A1(_00727_));
 sg13g2_mux4_1 _08526_ (.S0(net3517),
    .A0(\core.gpio.stray_data_i[6] ),
    .A1(\core.gpio.stray_data_i[14] ),
    .A2(\core.gpio.stray_data_i[22] ),
    .A3(\core.gpio.stray_data_i[30] ),
    .S1(net3515),
    .X(_02866_));
 sg13g2_nand2_2 _08527_ (.Y(_02867_),
    .A(net3514),
    .B(_02866_));
 sg13g2_mux2_1 _08528_ (.A0(_00139_),
    .A1(_00138_),
    .S(net3521),
    .X(_02868_));
 sg13g2_nand2b_1 _08529_ (.Y(_02869_),
    .B(_02868_),
    .A_N(net2767));
 sg13g2_nand2_1 _08530_ (.Y(_02870_),
    .A(net2767),
    .B(_02867_));
 sg13g2_nand3_1 _08531_ (.B(_02869_),
    .C(_02870_),
    .A(_02829_),
    .Y(_02871_));
 sg13g2_o21ai_1 _08532_ (.B1(_02763_),
    .Y(_02872_),
    .A1(_02803_),
    .A2(_02868_));
 sg13g2_nor2_1 _08533_ (.A(net3144),
    .B(_02867_),
    .Y(_02873_));
 sg13g2_nor2_1 _08534_ (.A(_00087_),
    .B(_02789_),
    .Y(_02874_));
 sg13g2_nor2_1 _08535_ (.A(_00091_),
    .B(_02787_),
    .Y(_02875_));
 sg13g2_nor3_2 _08536_ (.A(_02873_),
    .B(_02874_),
    .C(_02875_),
    .Y(_02876_));
 sg13g2_a22oi_1 _08537_ (.Y(_02877_),
    .B1(_02876_),
    .B2(_02795_),
    .A2(_02868_),
    .A1(net3142));
 sg13g2_nor2_1 _08538_ (.A(_02872_),
    .B(_02877_),
    .Y(_02878_));
 sg13g2_a22oi_1 _08539_ (.Y(_00389_),
    .B1(_02871_),
    .B2(_02878_),
    .A2(net3293),
    .A1(_00728_));
 sg13g2_mux4_1 _08540_ (.S0(net3517),
    .A0(\core.gpio.stray_data_i[7] ),
    .A1(\core.gpio.stray_data_i[15] ),
    .A2(\core.gpio.stray_data_i[23] ),
    .A3(\core.gpio.stray_data_i[31] ),
    .S1(net3515),
    .X(_02879_));
 sg13g2_nand2_1 _08541_ (.Y(_02880_),
    .A(_00057_),
    .B(_02879_));
 sg13g2_mux2_1 _08542_ (.A0(_00140_),
    .A1(_00139_),
    .S(net3521),
    .X(_02881_));
 sg13g2_mux2_1 _08543_ (.A0(_02881_),
    .A1(_02880_),
    .S(net2767),
    .X(_02882_));
 sg13g2_nor2_1 _08544_ (.A(net3144),
    .B(_02880_),
    .Y(_02883_));
 sg13g2_nor2_1 _08545_ (.A(_02799_),
    .B(_02881_),
    .Y(_02884_));
 sg13g2_a221oi_1 _08546_ (.B2(net3520),
    .C1(_02883_),
    .B1(_02788_),
    .A1(_00670_),
    .Y(_02885_),
    .A2(_02786_));
 sg13g2_a22oi_1 _08547_ (.Y(_02886_),
    .B1(_02885_),
    .B2(_02795_),
    .A2(_02881_),
    .A1(net3142));
 sg13g2_nor3_1 _08548_ (.A(_02791_),
    .B(_02884_),
    .C(_02886_),
    .Y(_02887_));
 sg13g2_o21ai_1 _08549_ (.B1(_02887_),
    .Y(_02888_),
    .A1(_02830_),
    .A2(_02882_));
 sg13g2_a21oi_1 _08550_ (.A1(_02791_),
    .A2(_02881_),
    .Y(_02889_),
    .B1(net3293));
 sg13g2_a22oi_1 _08551_ (.Y(_02890_),
    .B1(_02888_),
    .B2(_02889_),
    .A2(net3294),
    .A1(net677));
 sg13g2_inv_1 _08552_ (.Y(_00390_),
    .A(_02890_));
 sg13g2_o21ai_1 _08553_ (.B1(_02772_),
    .Y(_02891_),
    .A1(_00084_),
    .A2(net3150));
 sg13g2_o21ai_1 _08554_ (.B1(net2975),
    .Y(_02892_),
    .A1(_00587_),
    .A2(net3143));
 sg13g2_nand3_1 _08555_ (.B(_02891_),
    .C(_02892_),
    .A(_02763_),
    .Y(_02893_));
 sg13g2_a21oi_1 _08556_ (.A1(_01001_),
    .A2(net2768),
    .Y(_02894_),
    .B1(_02893_));
 sg13g2_nand2b_1 _08557_ (.Y(_02895_),
    .B(net3150),
    .A_N(_01055_));
 sg13g2_o21ai_1 _08558_ (.B1(_02895_),
    .Y(_02896_),
    .A1(_00085_),
    .A2(net3150));
 sg13g2_nor2_1 _08559_ (.A(net481),
    .B(net2757),
    .Y(_02897_));
 sg13g2_a21oi_1 _08560_ (.A1(net2757),
    .A2(_02896_),
    .Y(_00391_),
    .B1(_02897_));
 sg13g2_nor2_1 _08561_ (.A(net672),
    .B(net2757),
    .Y(_02898_));
 sg13g2_nand2_1 _08562_ (.Y(_02899_),
    .A(\core.lsu.spi.addr[0] ),
    .B(\core.lsu.spi.addr[1] ));
 sg13g2_or2_1 _08563_ (.X(_02900_),
    .B(\core.lsu.spi.addr[1] ),
    .A(\core.lsu.spi.addr[0] ));
 sg13g2_and3_1 _08564_ (.X(_02901_),
    .A(net2973),
    .B(_02899_),
    .C(_02900_));
 sg13g2_a21oi_1 _08565_ (.A1(_01053_),
    .A2(net3150),
    .Y(_02902_),
    .B1(_02901_));
 sg13g2_a21oi_1 _08566_ (.A1(net2757),
    .A2(_02902_),
    .Y(_00392_),
    .B1(_02898_));
 sg13g2_xnor2_1 _08567_ (.Y(_02903_),
    .A(\core.lsu.spi.addr[2] ),
    .B(_02899_));
 sg13g2_nand2_1 _08568_ (.Y(_02904_),
    .A(_01059_),
    .B(net3150));
 sg13g2_o21ai_1 _08569_ (.B1(_02904_),
    .Y(_02905_),
    .A1(net3150),
    .A2(_02903_));
 sg13g2_nor2_1 _08570_ (.A(net551),
    .B(net2757),
    .Y(_02906_));
 sg13g2_a21oi_1 _08571_ (.A1(net2757),
    .A2(_02905_),
    .Y(_00393_),
    .B1(_02906_));
 sg13g2_nor2_1 _08572_ (.A(_01050_),
    .B(net2973),
    .Y(_02907_));
 sg13g2_nor2_1 _08573_ (.A(_00086_),
    .B(_02899_),
    .Y(_02908_));
 sg13g2_xnor2_1 _08574_ (.Y(_02909_),
    .A(\core.lsu.spi.addr[3] ),
    .B(_02908_));
 sg13g2_a21oi_1 _08575_ (.A1(net2973),
    .A2(_02909_),
    .Y(_02910_),
    .B1(_02907_));
 sg13g2_mux2_1 _08576_ (.A0(net716),
    .A1(_02910_),
    .S(net2757),
    .X(_00394_));
 sg13g2_nand4_1 _08577_ (.B(\core.lsu.spi.addr[1] ),
    .C(\core.lsu.spi.addr[3] ),
    .A(\core.lsu.spi.addr[0] ),
    .Y(_02911_),
    .D(\core.lsu.spi.addr[2] ));
 sg13g2_inv_1 _08578_ (.Y(_02912_),
    .A(_02911_));
 sg13g2_xor2_1 _08579_ (.B(_02911_),
    .A(\core.lsu.spi.addr[4] ),
    .X(_02913_));
 sg13g2_nand2_1 _08580_ (.Y(_02914_),
    .A(net2974),
    .B(_02913_));
 sg13g2_o21ai_1 _08581_ (.B1(_02914_),
    .Y(_02915_),
    .A1(_01046_),
    .A2(net2973));
 sg13g2_nor2_1 _08582_ (.A(net509),
    .B(net2760),
    .Y(_02916_));
 sg13g2_a21oi_1 _08583_ (.A1(net2760),
    .A2(_02915_),
    .Y(_00395_),
    .B1(_02916_));
 sg13g2_nor2_1 _08584_ (.A(_00089_),
    .B(_02911_),
    .Y(_02917_));
 sg13g2_xnor2_1 _08585_ (.Y(_02918_),
    .A(net556),
    .B(_02917_));
 sg13g2_nor2_1 _08586_ (.A(net3149),
    .B(_02918_),
    .Y(_02919_));
 sg13g2_a21oi_1 _08587_ (.A1(_01044_),
    .A2(net3149),
    .Y(_02920_),
    .B1(_02919_));
 sg13g2_nor2_1 _08588_ (.A(net556),
    .B(net2757),
    .Y(_02921_));
 sg13g2_a21oi_1 _08589_ (.A1(net2758),
    .A2(_02920_),
    .Y(_00396_),
    .B1(_02921_));
 sg13g2_nand3_1 _08590_ (.B(\core.lsu.spi.addr[4] ),
    .C(_02912_),
    .A(\core.lsu.spi.addr[5] ),
    .Y(_02922_));
 sg13g2_and2_1 _08591_ (.A(_00667_),
    .B(_02922_),
    .X(_02923_));
 sg13g2_nor2_1 _08592_ (.A(_00667_),
    .B(_02922_),
    .Y(_02924_));
 sg13g2_nor3_1 _08593_ (.A(net3148),
    .B(_02923_),
    .C(_02924_),
    .Y(_02925_));
 sg13g2_and2_1 _08594_ (.A(_01071_),
    .B(net3147),
    .X(_02926_));
 sg13g2_o21ai_1 _08595_ (.B1(net2760),
    .Y(_02927_),
    .A1(_02925_),
    .A2(_02926_));
 sg13g2_o21ai_1 _08596_ (.B1(_02927_),
    .Y(_00397_),
    .A1(_00667_),
    .A2(net2760));
 sg13g2_nor2_1 _08597_ (.A(_00087_),
    .B(_02922_),
    .Y(_02928_));
 sg13g2_xor2_1 _08598_ (.B(_02928_),
    .A(net3520),
    .X(_02929_));
 sg13g2_nand2_1 _08599_ (.Y(_02930_),
    .A(_01041_),
    .B(net3148));
 sg13g2_o21ai_1 _08600_ (.B1(_02930_),
    .Y(_02931_),
    .A1(net3147),
    .A2(_02929_));
 sg13g2_nor2_1 _08601_ (.A(net3520),
    .B(net2760),
    .Y(_02932_));
 sg13g2_a21oi_1 _08602_ (.A1(net2760),
    .A2(_02931_),
    .Y(_00398_),
    .B1(_02932_));
 sg13g2_nand2_1 _08603_ (.Y(_02933_),
    .A(_01036_),
    .B(net3148));
 sg13g2_nand2_1 _08604_ (.Y(_02934_),
    .A(net3520),
    .B(_02924_));
 sg13g2_xnor2_1 _08605_ (.Y(_02935_),
    .A(net558),
    .B(_02934_));
 sg13g2_o21ai_1 _08606_ (.B1(_02933_),
    .Y(_02936_),
    .A1(net3148),
    .A2(_02935_));
 sg13g2_nor2_1 _08607_ (.A(net558),
    .B(net2760),
    .Y(_02937_));
 sg13g2_a21oi_1 _08608_ (.A1(net2760),
    .A2(_02936_),
    .Y(_00399_),
    .B1(_02937_));
 sg13g2_nor2_1 _08609_ (.A(_00095_),
    .B(_02934_),
    .Y(_02938_));
 sg13g2_xnor2_1 _08610_ (.Y(_02939_),
    .A(net578),
    .B(_02938_));
 sg13g2_nor2_1 _08611_ (.A(_01033_),
    .B(net2974),
    .Y(_02940_));
 sg13g2_a21oi_1 _08612_ (.A1(net2974),
    .A2(_02939_),
    .Y(_02941_),
    .B1(_02940_));
 sg13g2_nand2_1 _08613_ (.Y(_02942_),
    .A(net2761),
    .B(_02941_));
 sg13g2_o21ai_1 _08614_ (.B1(_02942_),
    .Y(_00400_),
    .A1(_00675_),
    .A2(net2761));
 sg13g2_nand4_1 _08615_ (.B(\core.lsu.spi.addr[9] ),
    .C(\core.lsu.spi.addr[8] ),
    .A(net3520),
    .Y(_02943_),
    .D(_02924_));
 sg13g2_nor2_1 _08616_ (.A(_00673_),
    .B(_02943_),
    .Y(_02944_));
 sg13g2_xnor2_1 _08617_ (.Y(_02945_),
    .A(_00673_),
    .B(_02943_));
 sg13g2_nand2_1 _08618_ (.Y(_02946_),
    .A(_01030_),
    .B(net3147));
 sg13g2_o21ai_1 _08619_ (.B1(_02946_),
    .Y(_02947_),
    .A1(net3147),
    .A2(_02945_));
 sg13g2_nand2_1 _08620_ (.Y(_02948_),
    .A(net2759),
    .B(_02947_));
 sg13g2_o21ai_1 _08621_ (.B1(_02948_),
    .Y(_00401_),
    .A1(_00673_),
    .A2(net2759));
 sg13g2_nor2_1 _08622_ (.A(_00093_),
    .B(_02943_),
    .Y(_02949_));
 sg13g2_xnor2_1 _08623_ (.Y(_02950_),
    .A(\core.lsu.spi.addr[11] ),
    .B(_02949_));
 sg13g2_nor2_1 _08624_ (.A(net3147),
    .B(_02950_),
    .Y(_02951_));
 sg13g2_a21oi_1 _08625_ (.A1(_01025_),
    .A2(net3147),
    .Y(_02952_),
    .B1(_02951_));
 sg13g2_nor2_1 _08626_ (.A(net779),
    .B(net2759),
    .Y(_02953_));
 sg13g2_a21oi_1 _08627_ (.A1(net2759),
    .A2(_02952_),
    .Y(_00402_),
    .B1(_02953_));
 sg13g2_nand2_1 _08628_ (.Y(_02954_),
    .A(\core.lsu.spi.addr[11] ),
    .B(_02944_));
 sg13g2_nand2_1 _08629_ (.Y(_02955_),
    .A(_01020_),
    .B(net3147));
 sg13g2_xnor2_1 _08630_ (.Y(_02956_),
    .A(net561),
    .B(_02954_));
 sg13g2_o21ai_1 _08631_ (.B1(_02955_),
    .Y(_02957_),
    .A1(net3147),
    .A2(_02956_));
 sg13g2_nor2_1 _08632_ (.A(net561),
    .B(net2759),
    .Y(_02958_));
 sg13g2_a21oi_1 _08633_ (.A1(net2759),
    .A2(_02957_),
    .Y(_00403_),
    .B1(_02958_));
 sg13g2_nor2_1 _08634_ (.A(_00092_),
    .B(_02954_),
    .Y(_02959_));
 sg13g2_xnor2_1 _08635_ (.Y(_02960_),
    .A(\core.lsu.spi.addr[13] ),
    .B(_02959_));
 sg13g2_nor2_1 _08636_ (.A(_01018_),
    .B(net2974),
    .Y(_02961_));
 sg13g2_a21oi_1 _08637_ (.A1(net2974),
    .A2(_02960_),
    .Y(_02962_),
    .B1(_02961_));
 sg13g2_nand2_1 _08638_ (.Y(_02963_),
    .A(net2761),
    .B(_02962_));
 sg13g2_o21ai_1 _08639_ (.B1(_02963_),
    .Y(_00404_),
    .A1(_00672_),
    .A2(net2759));
 sg13g2_nor2_1 _08640_ (.A(_01016_),
    .B(net2973),
    .Y(_02964_));
 sg13g2_nand4_1 _08641_ (.B(\core.lsu.spi.addr[12] ),
    .C(\core.lsu.spi.addr[11] ),
    .A(\core.lsu.spi.addr[13] ),
    .Y(_02965_),
    .D(_02944_));
 sg13g2_xnor2_1 _08642_ (.Y(_02966_),
    .A(_00671_),
    .B(_02965_));
 sg13g2_a21oi_1 _08643_ (.A1(net2973),
    .A2(_02966_),
    .Y(_02967_),
    .B1(_02964_));
 sg13g2_nand2_1 _08644_ (.Y(_02968_),
    .A(net2759),
    .B(_02967_));
 sg13g2_o21ai_1 _08645_ (.B1(_02968_),
    .Y(_00405_),
    .A1(_00671_),
    .A2(net2758));
 sg13g2_nor2_1 _08646_ (.A(_00091_),
    .B(_02965_),
    .Y(_02969_));
 sg13g2_nand3_1 _08647_ (.B(net2973),
    .C(_02969_),
    .A(net372),
    .Y(_02970_));
 sg13g2_o21ai_1 _08648_ (.B1(_02970_),
    .Y(_02971_),
    .A1(_01100_),
    .A2(net2973));
 sg13g2_o21ai_1 _08649_ (.B1(net2758),
    .Y(_02972_),
    .A1(net3149),
    .A2(_02969_));
 sg13g2_a22oi_1 _08650_ (.Y(_00406_),
    .B1(_02972_),
    .B2(_00669_),
    .A2(_02971_),
    .A1(net2758));
 sg13g2_o21ai_1 _08651_ (.B1(net3144),
    .Y(_02973_),
    .A1(_00585_),
    .A2(_02785_));
 sg13g2_nand3_1 _08652_ (.B(_02785_),
    .C(_02789_),
    .A(net3144),
    .Y(_02974_));
 sg13g2_nor2_1 _08653_ (.A(net2975),
    .B(_02974_),
    .Y(_02975_));
 sg13g2_a221oi_1 _08654_ (.B2(_01000_),
    .C1(_02798_),
    .B1(_02975_),
    .A1(net3143),
    .Y(_02976_),
    .A2(_02974_));
 sg13g2_nand3_1 _08655_ (.B(_02892_),
    .C(_02976_),
    .A(\core.lsu.spi.cs ),
    .Y(_02977_));
 sg13g2_nand2b_1 _08656_ (.Y(_02978_),
    .B(_02975_),
    .A_N(net2768));
 sg13g2_nor2_1 _08657_ (.A(_02788_),
    .B(_02977_),
    .Y(_02979_));
 sg13g2_a22oi_1 _08658_ (.Y(_00407_),
    .B1(_02978_),
    .B2(_02979_),
    .A2(_02977_),
    .A1(_00584_));
 sg13g2_nor3_1 _08659_ (.A(_02786_),
    .B(_02788_),
    .C(_02977_),
    .Y(_02980_));
 sg13g2_a21oi_1 _08660_ (.A1(_00583_),
    .A2(_02977_),
    .Y(_00408_),
    .B1(_02980_));
 sg13g2_nor2_1 _08661_ (.A(_02973_),
    .B(_02977_),
    .Y(_02981_));
 sg13g2_nand2b_1 _08662_ (.Y(_02982_),
    .B(_02975_),
    .A_N(_01124_));
 sg13g2_a22oi_1 _08663_ (.Y(_00409_),
    .B1(_02981_),
    .B2(_02982_),
    .A2(_02977_),
    .A1(_00585_));
 sg13g2_a21oi_2 _08664_ (.B1(_02605_),
    .Y(_02983_),
    .A2(net3151),
    .A1(_01126_));
 sg13g2_a21oi_1 _08665_ (.A1(net3155),
    .A2(_02606_),
    .Y(_02984_),
    .B1(net3517));
 sg13g2_a21oi_1 _08666_ (.A1(net3517),
    .A2(_02983_),
    .Y(_00410_),
    .B1(_02984_));
 sg13g2_a21oi_1 _08667_ (.A1(net3517),
    .A2(_02983_),
    .Y(_02985_),
    .B1(net3515));
 sg13g2_nand2_1 _08668_ (.Y(_02986_),
    .A(net3155),
    .B(_02722_));
 sg13g2_a21oi_1 _08669_ (.A1(_02983_),
    .A2(_02986_),
    .Y(_00411_),
    .B1(_02985_));
 sg13g2_a21oi_1 _08670_ (.A1(net3514),
    .A2(_02722_),
    .Y(_02987_),
    .B1(net3152));
 sg13g2_o21ai_1 _08671_ (.B1(_02987_),
    .Y(_02988_),
    .A1(net3514),
    .A2(_02722_));
 sg13g2_nor2_1 _08672_ (.A(net880),
    .B(_02983_),
    .Y(_02989_));
 sg13g2_a21oi_1 _08673_ (.A1(_02983_),
    .A2(_02988_),
    .Y(_00412_),
    .B1(_02989_));
 sg13g2_nor2_1 _08674_ (.A(_00084_),
    .B(_02784_),
    .Y(_02990_));
 sg13g2_a21oi_1 _08675_ (.A1(_00999_),
    .A2(net3142),
    .Y(_02991_),
    .B1(_02990_));
 sg13g2_nand2_1 _08676_ (.Y(_02992_),
    .A(_02799_),
    .B(_02991_));
 sg13g2_nand2_2 _08677_ (.Y(_02993_),
    .A(\core.lsu.spi.cs ),
    .B(_02992_));
 sg13g2_xnor2_1 _08678_ (.Y(_02994_),
    .A(net653),
    .B(net3521));
 sg13g2_nand2_1 _08679_ (.Y(_02995_),
    .A(net653),
    .B(_00666_));
 sg13g2_o21ai_1 _08680_ (.B1(_02995_),
    .Y(_00413_),
    .A1(_02993_),
    .A2(_02994_));
 sg13g2_nand2_1 _08681_ (.Y(_02996_),
    .A(\core.lsu.spi.counter[1] ),
    .B(_00666_));
 sg13g2_nor2_1 _08682_ (.A(net3521),
    .B(net406),
    .Y(_02997_));
 sg13g2_nor2_1 _08683_ (.A(\core.lsu.spi.counter[1] ),
    .B(\core.lsu.spi.counter[0] ),
    .Y(_02998_));
 sg13g2_xnor2_1 _08684_ (.Y(_02999_),
    .A(\core.lsu.spi.counter[1] ),
    .B(\core.lsu.spi.counter[0] ));
 sg13g2_a21oi_1 _08685_ (.A1(net3521),
    .A2(_02999_),
    .Y(_03000_),
    .B1(_02997_));
 sg13g2_o21ai_1 _08686_ (.B1(_02996_),
    .Y(_00414_),
    .A1(_02993_),
    .A2(net407));
 sg13g2_nand2_1 _08687_ (.Y(_03001_),
    .A(net379),
    .B(_00666_));
 sg13g2_nand2_1 _08688_ (.Y(_03002_),
    .A(net3522),
    .B(_02998_));
 sg13g2_xnor2_1 _08689_ (.Y(_03003_),
    .A(_00129_),
    .B(_03002_));
 sg13g2_o21ai_1 _08690_ (.B1(_03001_),
    .Y(_00415_),
    .A1(_02993_),
    .A2(_03003_));
 sg13g2_a21oi_1 _08691_ (.A1(_02769_),
    .A2(_02779_),
    .Y(_03004_),
    .B1(_02772_));
 sg13g2_or2_1 _08692_ (.X(_03005_),
    .B(_03002_),
    .A(\core.lsu.spi.counter[2] ));
 sg13g2_xnor2_1 _08693_ (.Y(_03006_),
    .A(_00130_),
    .B(_03005_));
 sg13g2_nor2_1 _08694_ (.A(_00998_),
    .B(net3142),
    .Y(_03007_));
 sg13g2_a21oi_1 _08695_ (.A1(_00998_),
    .A2(_02799_),
    .Y(_03008_),
    .B1(_03006_));
 sg13g2_nor4_1 _08696_ (.A(_02990_),
    .B(_03004_),
    .C(_03007_),
    .D(_03008_),
    .Y(_03009_));
 sg13g2_a21oi_1 _08697_ (.A1(_02990_),
    .A2(_03006_),
    .Y(_03010_),
    .B1(_03009_));
 sg13g2_mux2_1 _08698_ (.A0(net484),
    .A1(_03010_),
    .S(\core.lsu.spi.cs ),
    .X(_00416_));
 sg13g2_xor2_1 _08699_ (.B(_01057_),
    .A(_01056_),
    .X(_03011_));
 sg13g2_nor2_1 _08700_ (.A(\core.lsu.spi.counter[3] ),
    .B(_03005_),
    .Y(_03012_));
 sg13g2_xnor2_1 _08701_ (.Y(_03013_),
    .A(_00131_),
    .B(_03012_));
 sg13g2_a221oi_1 _08702_ (.B2(_02992_),
    .C1(_00666_),
    .B1(_03013_),
    .A1(_02829_),
    .Y(_03014_),
    .A2(_03011_));
 sg13g2_a21oi_1 _08703_ (.A1(_00586_),
    .A2(_00666_),
    .Y(_00417_),
    .B1(_03014_));
 sg13g2_nand2_1 _08704_ (.Y(_03015_),
    .A(_00586_),
    .B(_03012_));
 sg13g2_xnor2_1 _08705_ (.Y(_03016_),
    .A(_00132_),
    .B(_03015_));
 sg13g2_nand2_1 _08706_ (.Y(_03017_),
    .A(net362),
    .B(_00666_));
 sg13g2_o21ai_1 _08707_ (.B1(_03017_),
    .Y(_00418_),
    .A1(_02993_),
    .A2(_03016_));
 sg13g2_nand2_1 _08708_ (.Y(_03018_),
    .A(net3585),
    .B(net2736));
 sg13g2_nor4_1 _08709_ (.A(_01138_),
    .B(_02423_),
    .C(_02424_),
    .D(_03018_),
    .Y(_03019_));
 sg13g2_nor2_1 _08710_ (.A(net3513),
    .B(net2717),
    .Y(_03020_));
 sg13g2_nor4_2 _08711_ (.A(net3527),
    .B(net3528),
    .C(net3529),
    .Y(_03021_),
    .D(_00656_));
 sg13g2_nor2_1 _08712_ (.A(net3513),
    .B(net3140),
    .Y(_03022_));
 sg13g2_a21oi_2 _08713_ (.B1(_03022_),
    .Y(_03023_),
    .A2(net3140),
    .A1(net477));
 sg13g2_nor2_1 _08714_ (.A(\core.f2e_inst[16] ),
    .B(net3340),
    .Y(_03024_));
 sg13g2_a221oi_1 _08715_ (.B2(net3040),
    .C1(_03024_),
    .B1(net3043),
    .A1(_00676_),
    .Y(_03025_),
    .A2(net3340));
 sg13g2_a21oi_1 _08716_ (.A1(net2880),
    .A2(_03023_),
    .Y(_03026_),
    .B1(_03025_));
 sg13g2_a21oi_1 _08717_ (.A1(net2715),
    .A2(_03026_),
    .Y(_00419_),
    .B1(_03020_));
 sg13g2_nor2_1 _08718_ (.A(net3512),
    .B(net2717),
    .Y(_03027_));
 sg13g2_nor2_1 _08719_ (.A(net3512),
    .B(net3140),
    .Y(_03028_));
 sg13g2_a21oi_2 _08720_ (.B1(_03028_),
    .Y(_03029_),
    .A2(net3140),
    .A1(_00097_));
 sg13g2_nor2_1 _08721_ (.A(\core.f2e_inst[17] ),
    .B(net3340),
    .Y(_03030_));
 sg13g2_a221oi_1 _08722_ (.B2(net3040),
    .C1(_03030_),
    .B1(net3043),
    .A1(_00677_),
    .Y(_03031_),
    .A2(net3340));
 sg13g2_a21oi_1 _08723_ (.A1(net2880),
    .A2(_03029_),
    .Y(_03032_),
    .B1(_03031_));
 sg13g2_a21oi_1 _08724_ (.A1(net2717),
    .A2(_03032_),
    .Y(_00420_),
    .B1(_03027_));
 sg13g2_nor2_1 _08725_ (.A(net656),
    .B(net2727),
    .Y(_03033_));
 sg13g2_nor2_1 _08726_ (.A(\core.f2e_inst[2] ),
    .B(_03021_),
    .Y(_03034_));
 sg13g2_a21oi_1 _08727_ (.A1(net601),
    .A2(net3140),
    .Y(_03035_),
    .B1(_03034_));
 sg13g2_nor2_1 _08728_ (.A(net585),
    .B(net3339),
    .Y(_03036_));
 sg13g2_a221oi_1 _08729_ (.B2(net3041),
    .C1(_03036_),
    .B1(net3044),
    .A1(_00678_),
    .Y(_03037_),
    .A2(net3339));
 sg13g2_a21oi_1 _08730_ (.A1(net2884),
    .A2(_03035_),
    .Y(_03038_),
    .B1(_03037_));
 sg13g2_a21oi_1 _08731_ (.A1(net2727),
    .A2(_03038_),
    .Y(_00421_),
    .B1(_03033_));
 sg13g2_nor2_1 _08732_ (.A(net658),
    .B(net2717),
    .Y(_03039_));
 sg13g2_nor2_1 _08733_ (.A(\core.f2e_inst[3] ),
    .B(net3141),
    .Y(_03040_));
 sg13g2_a21oi_1 _08734_ (.A1(net452),
    .A2(net3140),
    .Y(_03041_),
    .B1(_03040_));
 sg13g2_nor2_1 _08735_ (.A(\core.f2e_inst[19] ),
    .B(net3342),
    .Y(_03042_));
 sg13g2_a221oi_1 _08736_ (.B2(net3040),
    .C1(_03042_),
    .B1(net3043),
    .A1(_00682_),
    .Y(_03043_),
    .A2(net3342));
 sg13g2_a21oi_1 _08737_ (.A1(net2882),
    .A2(_03041_),
    .Y(_03044_),
    .B1(_03043_));
 sg13g2_a21oi_1 _08738_ (.A1(net2717),
    .A2(_03044_),
    .Y(_00422_),
    .B1(_03039_));
 sg13g2_nor2_1 _08739_ (.A(net712),
    .B(net2728),
    .Y(_03045_));
 sg13g2_nor2_1 _08740_ (.A(\core.f2e_inst[4] ),
    .B(net3141),
    .Y(_03046_));
 sg13g2_a21oi_1 _08741_ (.A1(net500),
    .A2(net3141),
    .Y(_03047_),
    .B1(_03046_));
 sg13g2_nor2_1 _08742_ (.A(net543),
    .B(net3344),
    .Y(_03048_));
 sg13g2_a221oi_1 _08743_ (.B2(net3042),
    .C1(_03048_),
    .B1(net3044),
    .A1(_00685_),
    .Y(_03049_),
    .A2(net3344));
 sg13g2_a21oi_1 _08744_ (.A1(net2886),
    .A2(_03047_),
    .Y(_03050_),
    .B1(_03049_));
 sg13g2_a21oi_1 _08745_ (.A1(net2728),
    .A2(_03050_),
    .Y(_00423_),
    .B1(_03045_));
 sg13g2_nor2_1 _08746_ (.A(net3511),
    .B(net2727),
    .Y(_03051_));
 sg13g2_nor2_1 _08747_ (.A(net3511),
    .B(net3141),
    .Y(_03052_));
 sg13g2_a21oi_1 _08748_ (.A1(net421),
    .A2(net3141),
    .Y(_03053_),
    .B1(_03052_));
 sg13g2_nor2_1 _08749_ (.A(net581),
    .B(net3339),
    .Y(_03054_));
 sg13g2_a221oi_1 _08750_ (.B2(net3041),
    .C1(_03054_),
    .B1(net3044),
    .A1(_00687_),
    .Y(_03055_),
    .A2(net3335));
 sg13g2_a21oi_1 _08751_ (.A1(net2887),
    .A2(_03053_),
    .Y(_03056_),
    .B1(_03055_));
 sg13g2_a21oi_1 _08752_ (.A1(net2727),
    .A2(_03056_),
    .Y(_00424_),
    .B1(_03051_));
 sg13g2_nor2_1 _08753_ (.A(net3510),
    .B(net2727),
    .Y(_03057_));
 sg13g2_nor2_1 _08754_ (.A(net3510),
    .B(net3141),
    .Y(_03058_));
 sg13g2_a21oi_1 _08755_ (.A1(net429),
    .A2(net3141),
    .Y(_03059_),
    .B1(_03058_));
 sg13g2_nor2_1 _08756_ (.A(\core.f2e_inst[22] ),
    .B(net3344),
    .Y(_03060_));
 sg13g2_a221oi_1 _08757_ (.B2(net3041),
    .C1(_03060_),
    .B1(net3044),
    .A1(_00690_),
    .Y(_03061_),
    .A2(net3344));
 sg13g2_a21oi_1 _08758_ (.A1(net2887),
    .A2(_03059_),
    .Y(_03062_),
    .B1(_03061_));
 sg13g2_a21oi_1 _08759_ (.A1(net2727),
    .A2(_03062_),
    .Y(_00425_),
    .B1(_03057_));
 sg13g2_nor2_1 _08760_ (.A(net706),
    .B(net2721),
    .Y(_03063_));
 sg13g2_nor2_1 _08761_ (.A(\core.f2e_inst[7] ),
    .B(net3140),
    .Y(_03064_));
 sg13g2_a21oi_1 _08762_ (.A1(net411),
    .A2(net3140),
    .Y(_03065_),
    .B1(_03064_));
 sg13g2_nor2_1 _08763_ (.A(\core.f2e_inst[23] ),
    .B(net3344),
    .Y(_03066_));
 sg13g2_a221oi_1 _08764_ (.B2(net3041),
    .C1(_03066_),
    .B1(net3044),
    .A1(_00692_),
    .Y(_03067_),
    .A2(net3344));
 sg13g2_a21oi_1 _08765_ (.A1(net2884),
    .A2(_03065_),
    .Y(_03068_),
    .B1(_03067_));
 sg13g2_a21oi_1 _08766_ (.A1(net2721),
    .A2(_03068_),
    .Y(_00426_),
    .B1(_03063_));
 sg13g2_nor2_1 _08767_ (.A(net582),
    .B(net2725),
    .Y(_03069_));
 sg13g2_nand4_1 _08768_ (.B(_00581_),
    .C(net3529),
    .A(_00580_),
    .Y(_03070_),
    .D(_00656_));
 sg13g2_nor2_1 _08769_ (.A(net3570),
    .B(net3138),
    .Y(_03071_));
 sg13g2_a21oi_1 _08770_ (.A1(_00695_),
    .A2(net3138),
    .Y(_03072_),
    .B1(_03071_));
 sg13g2_nor2_1 _08771_ (.A(net555),
    .B(net3341),
    .Y(_03073_));
 sg13g2_a221oi_1 _08772_ (.B2(net3040),
    .C1(_03073_),
    .B1(net3043),
    .A1(_00694_),
    .Y(_03074_),
    .A2(net3341));
 sg13g2_a21oi_1 _08773_ (.A1(net2888),
    .A2(_03072_),
    .Y(_03075_),
    .B1(_03074_));
 sg13g2_a21oi_1 _08774_ (.A1(net2724),
    .A2(_03075_),
    .Y(_00427_),
    .B1(_03069_));
 sg13g2_nor2_1 _08775_ (.A(net722),
    .B(net2724),
    .Y(_03076_));
 sg13g2_mux2_1 _08776_ (.A0(net3569),
    .A1(\core.f2e_inst[9] ),
    .S(net3138),
    .X(_03077_));
 sg13g2_nor2_1 _08777_ (.A(net605),
    .B(net3340),
    .Y(_03078_));
 sg13g2_a221oi_1 _08778_ (.B2(net3040),
    .C1(_03078_),
    .B1(net3043),
    .A1(_00696_),
    .Y(_03079_),
    .A2(net3340));
 sg13g2_a21oi_1 _08779_ (.A1(net2882),
    .A2(_03077_),
    .Y(_03080_),
    .B1(_03079_));
 sg13g2_a21oi_1 _08780_ (.A1(net2724),
    .A2(_03080_),
    .Y(_00428_),
    .B1(_03076_));
 sg13g2_nor2_1 _08781_ (.A(net3509),
    .B(net2728),
    .Y(_03081_));
 sg13g2_mux2_1 _08782_ (.A0(\core.fetch.cmd_data[2] ),
    .A1(net3509),
    .S(net3139),
    .X(_03082_));
 sg13g2_nor2_1 _08783_ (.A(net518),
    .B(net3347),
    .Y(_03083_));
 sg13g2_a221oi_1 _08784_ (.B2(net3042),
    .C1(_03083_),
    .B1(net3045),
    .A1(_00697_),
    .Y(_03084_),
    .A2(net3347));
 sg13g2_a21oi_1 _08785_ (.A1(net2886),
    .A2(_03082_),
    .Y(_03085_),
    .B1(_03084_));
 sg13g2_a21oi_1 _08786_ (.A1(net2728),
    .A2(_03085_),
    .Y(_00429_),
    .B1(_03081_));
 sg13g2_nor2_1 _08787_ (.A(net689),
    .B(net2725),
    .Y(_03086_));
 sg13g2_nor2_1 _08788_ (.A(\core.fetch.cmd_data[3] ),
    .B(net3138),
    .Y(_03087_));
 sg13g2_a21oi_1 _08789_ (.A1(_00699_),
    .A2(net3138),
    .Y(_03088_),
    .B1(_03087_));
 sg13g2_nor2_1 _08790_ (.A(net603),
    .B(net3341),
    .Y(_03089_));
 sg13g2_a221oi_1 _08791_ (.B2(net3040),
    .C1(_03089_),
    .B1(net3043),
    .A1(_00698_),
    .Y(_03090_),
    .A2(net3341));
 sg13g2_a21oi_1 _08792_ (.A1(net2888),
    .A2(_03088_),
    .Y(_03091_),
    .B1(_03090_));
 sg13g2_a21oi_1 _08793_ (.A1(net2725),
    .A2(_03091_),
    .Y(_00430_),
    .B1(_03086_));
 sg13g2_nor2_1 _08794_ (.A(net3507),
    .B(net2724),
    .Y(_03092_));
 sg13g2_nor2_1 _08795_ (.A(\core.fetch.cmd_data[4] ),
    .B(net3139),
    .Y(_03093_));
 sg13g2_a21oi_1 _08796_ (.A1(_00701_),
    .A2(net3139),
    .Y(_03094_),
    .B1(_03093_));
 sg13g2_nor2_1 _08797_ (.A(net498),
    .B(net3342),
    .Y(_03095_));
 sg13g2_a221oi_1 _08798_ (.B2(net3041),
    .C1(_03095_),
    .B1(net3043),
    .A1(_00700_),
    .Y(_03096_),
    .A2(net3342));
 sg13g2_a21oi_1 _08799_ (.A1(net2888),
    .A2(_03094_),
    .Y(_03097_),
    .B1(_03096_));
 sg13g2_a21oi_1 _08800_ (.A1(net2725),
    .A2(_03097_),
    .Y(_00431_),
    .B1(_03092_));
 sg13g2_nor2_1 _08801_ (.A(net3505),
    .B(net2724),
    .Y(_03098_));
 sg13g2_mux2_1 _08802_ (.A0(\core.fetch.cmd_data[5] ),
    .A1(net3505),
    .S(net3138),
    .X(_03099_));
 sg13g2_nor2_1 _08803_ (.A(net545),
    .B(net3340),
    .Y(_03100_));
 sg13g2_a221oi_1 _08804_ (.B2(net3040),
    .C1(_03100_),
    .B1(net3043),
    .A1(_00702_),
    .Y(_03101_),
    .A2(net3340));
 sg13g2_a21oi_1 _08805_ (.A1(net2882),
    .A2(_03099_),
    .Y(_03102_),
    .B1(_03101_));
 sg13g2_a21oi_1 _08806_ (.A1(net2724),
    .A2(_03102_),
    .Y(_00432_),
    .B1(_03098_));
 sg13g2_nor2_1 _08807_ (.A(net715),
    .B(net2726),
    .Y(_03103_));
 sg13g2_nor2_1 _08808_ (.A(\core.fetch.cmd_data[6] ),
    .B(net3139),
    .Y(_03104_));
 sg13g2_a21oi_1 _08809_ (.A1(_00705_),
    .A2(net3138),
    .Y(_03105_),
    .B1(_03104_));
 sg13g2_nor2_1 _08810_ (.A(net574),
    .B(net3335),
    .Y(_03106_));
 sg13g2_a221oi_1 _08811_ (.B2(net3041),
    .C1(_03106_),
    .B1(net3045),
    .A1(_00703_),
    .Y(_03107_),
    .A2(net3335));
 sg13g2_a21oi_1 _08812_ (.A1(net2888),
    .A2(_03105_),
    .Y(_03108_),
    .B1(_03107_));
 sg13g2_a21oi_1 _08813_ (.A1(net2725),
    .A2(_03108_),
    .Y(_00433_),
    .B1(_03103_));
 sg13g2_nor2_1 _08814_ (.A(net794),
    .B(net2726),
    .Y(_03109_));
 sg13g2_nor2_1 _08815_ (.A(\core.fetch.cmd_data[7] ),
    .B(net3139),
    .Y(_03110_));
 sg13g2_a21oi_1 _08816_ (.A1(_00708_),
    .A2(net3138),
    .Y(_03111_),
    .B1(_03110_));
 sg13g2_nor2_1 _08817_ (.A(net534),
    .B(net3335),
    .Y(_03112_));
 sg13g2_a221oi_1 _08818_ (.B2(net3040),
    .C1(_03112_),
    .B1(net3045),
    .A1(_00706_),
    .Y(_03113_),
    .A2(net3335));
 sg13g2_a21oi_1 _08819_ (.A1(net2888),
    .A2(_03111_),
    .Y(_03114_),
    .B1(_03113_));
 sg13g2_a21oi_1 _08820_ (.A1(net2726),
    .A2(_03114_),
    .Y(_00434_),
    .B1(_03109_));
 sg13g2_nor3_1 _08821_ (.A(net3527),
    .B(_00581_),
    .C(net3529),
    .Y(_03115_));
 sg13g2_mux2_1 _08822_ (.A0(\core.f2e_inst[16] ),
    .A1(net3570),
    .S(net3136),
    .X(_03116_));
 sg13g2_a22oi_1 _08823_ (.Y(_03117_),
    .B1(_03116_),
    .B2(net2880),
    .A2(net2837),
    .A1(net472));
 sg13g2_nor2_1 _08824_ (.A(\core.f2e_inst[16] ),
    .B(net2715),
    .Y(_03118_));
 sg13g2_a21oi_1 _08825_ (.A1(net2715),
    .A2(net473),
    .Y(_00435_),
    .B1(_03118_));
 sg13g2_nor2_1 _08826_ (.A(\core.f2e_inst[17] ),
    .B(net2714),
    .Y(_03119_));
 sg13g2_mux2_1 _08827_ (.A0(\core.f2e_inst[17] ),
    .A1(net3569),
    .S(net3136),
    .X(_03120_));
 sg13g2_a22oi_1 _08828_ (.Y(_03121_),
    .B1(_03120_),
    .B2(net2880),
    .A2(net2837),
    .A1(net506));
 sg13g2_a21oi_1 _08829_ (.A1(net2714),
    .A2(net507),
    .Y(_00436_),
    .B1(_03119_));
 sg13g2_o21ai_1 _08830_ (.B1(net2883),
    .Y(_03122_),
    .A1(net450),
    .A2(net3137));
 sg13g2_a21oi_1 _08831_ (.A1(_00681_),
    .A2(net3136),
    .Y(_03123_),
    .B1(_03122_));
 sg13g2_a21oi_1 _08832_ (.A1(\core.fetch.inst[34] ),
    .A2(net2837),
    .Y(_03124_),
    .B1(_03123_));
 sg13g2_nor2_1 _08833_ (.A(net450),
    .B(net2723),
    .Y(_03125_));
 sg13g2_a21oi_1 _08834_ (.A1(net2720),
    .A2(_03124_),
    .Y(_00437_),
    .B1(_03125_));
 sg13g2_mux2_1 _08835_ (.A0(\core.f2e_inst[19] ),
    .A1(\core.fetch.cmd_data[3] ),
    .S(net3136),
    .X(_03126_));
 sg13g2_a22oi_1 _08836_ (.Y(_03127_),
    .B1(_03126_),
    .B2(net2881),
    .A2(net2837),
    .A1(net531));
 sg13g2_nor2_1 _08837_ (.A(\core.f2e_inst[19] ),
    .B(net2716),
    .Y(_03128_));
 sg13g2_a21oi_1 _08838_ (.A1(net2716),
    .A2(net532),
    .Y(_00438_),
    .B1(_03128_));
 sg13g2_nor2_1 _08839_ (.A(net543),
    .B(net2728),
    .Y(_03129_));
 sg13g2_nor2_1 _08840_ (.A(net543),
    .B(net3137),
    .Y(_03130_));
 sg13g2_a21oi_1 _08841_ (.A1(_00686_),
    .A2(net3137),
    .Y(_03131_),
    .B1(_03130_));
 sg13g2_a22oi_1 _08842_ (.Y(_03132_),
    .B1(_03131_),
    .B2(net2886),
    .A2(net2839),
    .A1(net520));
 sg13g2_a21oi_1 _08843_ (.A1(net2728),
    .A2(_03132_),
    .Y(_00439_),
    .B1(_03129_));
 sg13g2_nor2_1 _08844_ (.A(net419),
    .B(net2721),
    .Y(_03133_));
 sg13g2_nor2_1 _08845_ (.A(net419),
    .B(net3136),
    .Y(_03134_));
 sg13g2_a21oi_1 _08846_ (.A1(_00689_),
    .A2(net3136),
    .Y(_03135_),
    .B1(_03134_));
 sg13g2_a22oi_1 _08847_ (.Y(_03136_),
    .B1(_03135_),
    .B2(net2884),
    .A2(net2838),
    .A1(\core.fetch.inst[37] ));
 sg13g2_a21oi_1 _08848_ (.A1(net2722),
    .A2(_03136_),
    .Y(_00440_),
    .B1(_03133_));
 sg13g2_nor2_1 _08849_ (.A(\core.f2e_inst[22] ),
    .B(net2729),
    .Y(_03137_));
 sg13g2_nor2_1 _08850_ (.A(\core.f2e_inst[22] ),
    .B(net3137),
    .Y(_03138_));
 sg13g2_a21oi_1 _08851_ (.A1(_00691_),
    .A2(net3137),
    .Y(_03139_),
    .B1(_03138_));
 sg13g2_a22oi_1 _08852_ (.Y(_03140_),
    .B1(_03139_),
    .B2(net2887),
    .A2(net2839),
    .A1(net536));
 sg13g2_a21oi_1 _08853_ (.A1(net2729),
    .A2(net537),
    .Y(_00441_),
    .B1(_03137_));
 sg13g2_o21ai_1 _08854_ (.B1(net2884),
    .Y(_03141_),
    .A1(\core.f2e_inst[23] ),
    .A2(net3136));
 sg13g2_a21oi_1 _08855_ (.A1(_00693_),
    .A2(net3136),
    .Y(_03142_),
    .B1(_03141_));
 sg13g2_a21oi_1 _08856_ (.A1(net539),
    .A2(net2838),
    .Y(_03143_),
    .B1(_03142_));
 sg13g2_nor2_1 _08857_ (.A(\core.f2e_inst[23] ),
    .B(net2723),
    .Y(_03144_));
 sg13g2_a21oi_1 _08858_ (.A1(net2723),
    .A2(_03143_),
    .Y(_00442_),
    .B1(_03144_));
 sg13g2_mux2_1 _08859_ (.A0(net555),
    .A1(net3570),
    .S(net3158),
    .X(_03145_));
 sg13g2_a22oi_1 _08860_ (.Y(_03146_),
    .B1(_03145_),
    .B2(net2888),
    .A2(net2839),
    .A1(net528));
 sg13g2_nor2_1 _08861_ (.A(net555),
    .B(net2724),
    .Y(_03147_));
 sg13g2_a21oi_1 _08862_ (.A1(net2724),
    .A2(_03146_),
    .Y(_00443_),
    .B1(_03147_));
 sg13g2_mux2_1 _08863_ (.A0(\core.f2e_inst[25] ),
    .A1(net3569),
    .S(net3158),
    .X(_03148_));
 sg13g2_a22oi_1 _08864_ (.Y(_03149_),
    .B1(_03148_),
    .B2(net2880),
    .A2(net2837),
    .A1(net524));
 sg13g2_nor2_1 _08865_ (.A(net605),
    .B(net2714),
    .Y(_03150_));
 sg13g2_a21oi_1 _08866_ (.A1(net2714),
    .A2(_03149_),
    .Y(_00444_),
    .B1(_03150_));
 sg13g2_o21ai_1 _08867_ (.B1(net2887),
    .Y(_03151_),
    .A1(net518),
    .A2(net3159));
 sg13g2_a21oi_1 _08868_ (.A1(_00681_),
    .A2(net3159),
    .Y(_03152_),
    .B1(_03151_));
 sg13g2_a21oi_1 _08869_ (.A1(\core.fetch.inst[42] ),
    .A2(net2839),
    .Y(_03153_),
    .B1(_03152_));
 sg13g2_nor2_1 _08870_ (.A(net518),
    .B(net2728),
    .Y(_03154_));
 sg13g2_a21oi_1 _08871_ (.A1(net2728),
    .A2(_03153_),
    .Y(_00445_),
    .B1(_03154_));
 sg13g2_mux2_1 _08872_ (.A0(net603),
    .A1(\core.fetch.cmd_data[3] ),
    .S(net3158),
    .X(_03155_));
 sg13g2_a22oi_1 _08873_ (.Y(_03156_),
    .B1(_03155_),
    .B2(net2882),
    .A2(net2837),
    .A1(net564));
 sg13g2_nor2_1 _08874_ (.A(net603),
    .B(net2717),
    .Y(_03157_));
 sg13g2_a21oi_1 _08875_ (.A1(net2718),
    .A2(_03156_),
    .Y(_00446_),
    .B1(_03157_));
 sg13g2_o21ai_1 _08876_ (.B1(net2885),
    .Y(_03158_),
    .A1(net498),
    .A2(net3159));
 sg13g2_a21oi_1 _08877_ (.A1(_00686_),
    .A2(net3158),
    .Y(_03159_),
    .B1(_03158_));
 sg13g2_a21oi_1 _08878_ (.A1(\core.fetch.inst[44] ),
    .A2(net2838),
    .Y(_03160_),
    .B1(_03159_));
 sg13g2_nor2_1 _08879_ (.A(net498),
    .B(net2721),
    .Y(_03161_));
 sg13g2_a21oi_1 _08880_ (.A1(net2721),
    .A2(_03160_),
    .Y(_00447_),
    .B1(_03161_));
 sg13g2_o21ai_1 _08881_ (.B1(net2881),
    .Y(_03162_),
    .A1(net545),
    .A2(net3158));
 sg13g2_a21oi_1 _08882_ (.A1(_00689_),
    .A2(net3158),
    .Y(_03163_),
    .B1(_03162_));
 sg13g2_a21oi_1 _08883_ (.A1(net530),
    .A2(net2837),
    .Y(_03164_),
    .B1(_03163_));
 sg13g2_nor2_1 _08884_ (.A(net545),
    .B(net2716),
    .Y(_03165_));
 sg13g2_a21oi_1 _08885_ (.A1(net2716),
    .A2(_03164_),
    .Y(_00448_),
    .B1(_03165_));
 sg13g2_o21ai_1 _08886_ (.B1(net2883),
    .Y(_03166_),
    .A1(net486),
    .A2(net3159));
 sg13g2_a21oi_1 _08887_ (.A1(_00691_),
    .A2(net3158),
    .Y(_03167_),
    .B1(_03166_));
 sg13g2_a21oi_1 _08888_ (.A1(\core.fetch.inst[46] ),
    .A2(net2838),
    .Y(_03168_),
    .B1(_03167_));
 sg13g2_nor2_1 _08889_ (.A(net486),
    .B(net2720),
    .Y(_03169_));
 sg13g2_a21oi_1 _08890_ (.A1(net2720),
    .A2(_03168_),
    .Y(_00449_),
    .B1(_03169_));
 sg13g2_o21ai_1 _08891_ (.B1(net2883),
    .Y(_03170_),
    .A1(net448),
    .A2(net3158));
 sg13g2_a21oi_1 _08892_ (.A1(_00693_),
    .A2(net3159),
    .Y(_03171_),
    .B1(_03170_));
 sg13g2_a21oi_1 _08893_ (.A1(\core.fetch.inst[47] ),
    .A2(net2837),
    .Y(_03172_),
    .B1(_03171_));
 sg13g2_nor2_1 _08894_ (.A(net448),
    .B(net2719),
    .Y(_03173_));
 sg13g2_a21oi_1 _08895_ (.A1(net2719),
    .A2(_03172_),
    .Y(_00450_),
    .B1(_03173_));
 sg13g2_nand2_1 _08896_ (.Y(_03174_),
    .A(net3338),
    .B(_01327_));
 sg13g2_a21oi_1 _08897_ (.A1(net2736),
    .A2(_03174_),
    .Y(_03175_),
    .B1(_01138_));
 sg13g2_nand2_1 _08898_ (.Y(_03176_),
    .A(net2736),
    .B(_01571_));
 sg13g2_o21ai_1 _08899_ (.B1(_03176_),
    .Y(_03177_),
    .A1(_00709_),
    .A2(net2736));
 sg13g2_mux2_1 _08900_ (.A0(net3503),
    .A1(_03177_),
    .S(_03175_),
    .X(_00451_));
 sg13g2_nand3b_1 _08901_ (.B(_01124_),
    .C(_02763_),
    .Y(_03178_),
    .A_N(_02772_));
 sg13g2_mux2_1 _08902_ (.A0(\core.gpio.stray_wr_i ),
    .A1(net502),
    .S(_03178_),
    .X(_00452_));
 sg13g2_a21oi_1 _08903_ (.A1(net3562),
    .A2(_00596_),
    .Y(_03179_),
    .B1(net3545));
 sg13g2_and2_1 _08904_ (.A(net3538),
    .B(net3560),
    .X(_03180_));
 sg13g2_nand2_1 _08905_ (.Y(_03181_),
    .A(net3539),
    .B(net3562));
 sg13g2_nor3_2 _08906_ (.A(_01834_),
    .B(_03179_),
    .C(net3291),
    .Y(_03182_));
 sg13g2_nand3b_1 _08907_ (.B(net3308),
    .C(_01723_),
    .Y(_03183_),
    .A_N(_03182_));
 sg13g2_nor3_2 _08908_ (.A(\core.work.registers.state[1] ),
    .B(_00651_),
    .C(_00058_),
    .Y(_03184_));
 sg13g2_o21ai_1 _08909_ (.B1(_00055_),
    .Y(_03185_),
    .A1(_02436_),
    .A2(_03184_));
 sg13g2_a21oi_1 _08910_ (.A1(\core.work.alu.is_mem ),
    .A2(\core.lsu.accept ),
    .Y(_03186_),
    .B1(_01127_));
 sg13g2_a22oi_1 _08911_ (.Y(_03187_),
    .B1(_03185_),
    .B2(_03186_),
    .A2(_01326_),
    .A1(_01323_));
 sg13g2_nand3_1 _08912_ (.B(_03183_),
    .C(_03187_),
    .A(net3502),
    .Y(_03188_));
 sg13g2_nand3_1 _08913_ (.B(_03183_),
    .C(_03188_),
    .A(_01643_),
    .Y(_03189_));
 sg13g2_nand2_1 _08914_ (.Y(_00453_),
    .A(_01706_),
    .B(_03189_));
 sg13g2_a21o_1 _08915_ (.A2(_03188_),
    .A1(net3501),
    .B1(net2787),
    .X(_00454_));
 sg13g2_nor2_1 _08916_ (.A(net541),
    .B(net2786),
    .Y(_03190_));
 sg13g2_a21oi_1 _08917_ (.A1(_01702_),
    .A2(net2786),
    .Y(_00455_),
    .B1(_03190_));
 sg13g2_nor2_1 _08918_ (.A(net562),
    .B(net2786),
    .Y(_03191_));
 sg13g2_a21oi_1 _08919_ (.A1(_01698_),
    .A2(net2786),
    .Y(_00456_),
    .B1(_03191_));
 sg13g2_nor2_1 _08920_ (.A(net392),
    .B(net2786),
    .Y(_03192_));
 sg13g2_a21oi_1 _08921_ (.A1(_01694_),
    .A2(net2786),
    .Y(_00457_),
    .B1(_03192_));
 sg13g2_nor2_1 _08922_ (.A(net414),
    .B(net2786),
    .Y(_03193_));
 sg13g2_a21oi_1 _08923_ (.A1(_01696_),
    .A2(net2786),
    .Y(_00458_),
    .B1(_03193_));
 sg13g2_nand2_2 _08924_ (.Y(_03194_),
    .A(net3586),
    .B(net2787));
 sg13g2_nand2_1 _08925_ (.Y(_03195_),
    .A(net468),
    .B(net2781));
 sg13g2_nor2_1 _08926_ (.A(_01691_),
    .B(_03194_),
    .Y(_03196_));
 sg13g2_nand3_1 _08927_ (.B(net3195),
    .C(net2787),
    .A(net3588),
    .Y(_03197_));
 sg13g2_nand2_1 _08928_ (.Y(_03198_),
    .A(net3476),
    .B(\core.work.registers.genblk1[1].latch[0] ));
 sg13g2_nor2b_1 _08929_ (.A(net3469),
    .B_N(net3468),
    .Y(_03199_));
 sg13g2_nor2b_1 _08930_ (.A(net3476),
    .B_N(net3471),
    .Y(_03200_));
 sg13g2_and2_1 _08931_ (.A(_03199_),
    .B(_03200_),
    .X(_03201_));
 sg13g2_nor2_1 _08932_ (.A(net3476),
    .B(net3471),
    .Y(_03202_));
 sg13g2_and2_1 _08933_ (.A(_03199_),
    .B(_03202_),
    .X(_03203_));
 sg13g2_and2_1 _08934_ (.A(net3477),
    .B(net3471),
    .X(_03204_));
 sg13g2_nor2b_2 _08935_ (.A(net3468),
    .B_N(net3469),
    .Y(_03205_));
 sg13g2_and2_1 _08936_ (.A(_03204_),
    .B(_03205_),
    .X(_03206_));
 sg13g2_and2_1 _08937_ (.A(_03202_),
    .B(_03205_),
    .X(_03207_));
 sg13g2_and2_1 _08938_ (.A(_01655_),
    .B(_03200_),
    .X(_03208_));
 sg13g2_nand2_1 _08939_ (.Y(_03209_),
    .A(\core.work.registers.genblk1[2].latch[0] ),
    .B(net3114));
 sg13g2_and2_1 _08940_ (.A(_03200_),
    .B(_03205_),
    .X(_03210_));
 sg13g2_and2_1 _08941_ (.A(net3468),
    .B(net3469),
    .X(_03211_));
 sg13g2_and2_1 _08942_ (.A(_03200_),
    .B(_03211_),
    .X(_03212_));
 sg13g2_and2_1 _08943_ (.A(_03199_),
    .B(_03204_),
    .X(_03213_));
 sg13g2_and2_1 _08944_ (.A(_03202_),
    .B(_03211_),
    .X(_03214_));
 sg13g2_a22oi_1 _08945_ (.Y(_03215_),
    .B1(net3094),
    .B2(\core.work.registers.genblk1[12].latch[0] ),
    .A2(net3098),
    .A1(\core.work.registers.genblk1[11].latch[0] ));
 sg13g2_and2_1 _08946_ (.A(_01655_),
    .B(_03204_),
    .X(_03216_));
 sg13g2_nor2b_1 _08947_ (.A(net3471),
    .B_N(net3476),
    .Y(_03217_));
 sg13g2_and2_1 _08948_ (.A(_03205_),
    .B(_03217_),
    .X(_03218_));
 sg13g2_and2_1 _08949_ (.A(_03199_),
    .B(_03217_),
    .X(_03219_));
 sg13g2_and2_1 _08950_ (.A(_03204_),
    .B(_03211_),
    .X(_03220_));
 sg13g2_and2_1 _08951_ (.A(_03211_),
    .B(_03217_),
    .X(_03221_));
 sg13g2_a22oi_1 _08952_ (.Y(_03222_),
    .B1(net3123),
    .B2(\core.work.registers.genblk1[7].latch[0] ),
    .A2(net3134),
    .A1(\core.work.registers.genblk1[10].latch[0] ));
 sg13g2_a21oi_1 _08953_ (.A1(\core.work.registers.genblk1[8].latch[0] ),
    .A2(net3128),
    .Y(_03223_),
    .B1(net3326));
 sg13g2_a22oi_1 _08954_ (.Y(_03224_),
    .B1(net3073),
    .B2(\core.work.registers.genblk1[15].latch[0] ),
    .A2(net3089),
    .A1(\core.work.registers.genblk1[3].latch[0] ));
 sg13g2_and4_1 _08955_ (.A(_03215_),
    .B(_03222_),
    .C(_03223_),
    .D(_03224_),
    .X(_03225_));
 sg13g2_a22oi_1 _08956_ (.Y(_03226_),
    .B1(net3109),
    .B2(\core.work.registers.genblk1[6].latch[0] ),
    .A2(net3118),
    .A1(\core.work.registers.genblk1[4].latch[0] ));
 sg13g2_a22oi_1 _08957_ (.Y(_03227_),
    .B1(net3084),
    .B2(\core.work.registers.genblk1[5].latch[0] ),
    .A2(net3104),
    .A1(\core.work.registers.genblk1[14].latch[0] ));
 sg13g2_a22oi_1 _08958_ (.Y(_03228_),
    .B1(net3068),
    .B2(\core.work.registers.genblk1[13].latch[0] ),
    .A2(net3079),
    .A1(\core.work.registers.genblk1[9].latch[0] ));
 sg13g2_and4_1 _08959_ (.A(_03209_),
    .B(_03226_),
    .C(_03227_),
    .D(_03228_),
    .X(_03229_));
 sg13g2_a22oi_1 _08960_ (.Y(_03230_),
    .B1(_03225_),
    .B2(_03229_),
    .A2(_03198_),
    .A1(net3326));
 sg13g2_nand2b_1 _08961_ (.Y(_03231_),
    .B(net3460),
    .A_N(_03230_));
 sg13g2_nand2_1 _08962_ (.Y(_03232_),
    .A(net2919),
    .B(_03230_));
 sg13g2_nor2_1 _08963_ (.A(net3460),
    .B(_03232_),
    .Y(_03233_));
 sg13g2_nand3b_1 _08964_ (.B(net2919),
    .C(_03230_),
    .Y(_03234_),
    .A_N(net3460));
 sg13g2_nor2_1 _08965_ (.A(net2912),
    .B(_03233_),
    .Y(_03235_));
 sg13g2_a22oi_1 _08966_ (.Y(_03236_),
    .B1(_03231_),
    .B2(_03235_),
    .A2(_02128_),
    .A1(net2908));
 sg13g2_o21ai_1 _08967_ (.B1(_03195_),
    .Y(_00459_),
    .A1(_03197_),
    .A2(_03236_));
 sg13g2_nor2_1 _08968_ (.A(net2907),
    .B(_01763_),
    .Y(_03237_));
 sg13g2_nand2_1 _08969_ (.Y(_03238_),
    .A(_00640_),
    .B(net3035));
 sg13g2_o21ai_1 _08970_ (.B1(_03238_),
    .Y(_03239_),
    .A1(_00106_),
    .A2(net3036));
 sg13g2_nand2_1 _08971_ (.Y(_03240_),
    .A(\core.work.registers.genblk1[8].latch[1] ),
    .B(net3128));
 sg13g2_a22oi_1 _08972_ (.Y(_03241_),
    .B1(net3114),
    .B2(\core.work.registers.genblk1[2].latch[1] ),
    .A2(net3119),
    .A1(\core.work.registers.genblk1[4].latch[1] ));
 sg13g2_a22oi_1 _08973_ (.Y(_03242_),
    .B1(net3068),
    .B2(\core.work.registers.genblk1[13].latch[1] ),
    .A2(net3104),
    .A1(\core.work.registers.genblk1[14].latch[1] ));
 sg13g2_a21oi_1 _08974_ (.A1(\core.work.registers.genblk1[12].latch[1] ),
    .A2(net3094),
    .Y(_03243_),
    .B1(net3327));
 sg13g2_a22oi_1 _08975_ (.Y(_03244_),
    .B1(net3079),
    .B2(\core.work.registers.genblk1[9].latch[1] ),
    .A2(net3109),
    .A1(\core.work.registers.genblk1[6].latch[1] ));
 sg13g2_a22oi_1 _08976_ (.Y(_03245_),
    .B1(net3089),
    .B2(\core.work.registers.genblk1[3].latch[1] ),
    .A2(net3099),
    .A1(\core.work.registers.genblk1[11].latch[1] ));
 sg13g2_and4_1 _08977_ (.A(_03241_),
    .B(_03243_),
    .C(_03244_),
    .D(_03245_),
    .X(_03246_));
 sg13g2_a22oi_1 _08978_ (.Y(_03247_),
    .B1(net3084),
    .B2(\core.work.registers.genblk1[5].latch[1] ),
    .A2(net3123),
    .A1(\core.work.registers.genblk1[7].latch[1] ));
 sg13g2_a22oi_1 _08979_ (.Y(_03248_),
    .B1(net3074),
    .B2(\core.work.registers.genblk1[15].latch[1] ),
    .A2(net3134),
    .A1(\core.work.registers.genblk1[10].latch[1] ));
 sg13g2_and4_1 _08980_ (.A(_03240_),
    .B(_03242_),
    .C(_03247_),
    .D(_03248_),
    .X(_03249_));
 sg13g2_nand2_1 _08981_ (.Y(_03250_),
    .A(net3476),
    .B(\core.work.registers.genblk1[1].latch[1] ));
 sg13g2_a22oi_1 _08982_ (.Y(_03251_),
    .B1(_03250_),
    .B2(net3327),
    .A2(_03249_),
    .A1(_03246_));
 sg13g2_a221oi_1 _08983_ (.B2(net3327),
    .C1(net2912),
    .B1(_03250_),
    .A1(_03246_),
    .Y(_03252_),
    .A2(_03249_));
 sg13g2_nor2_1 _08984_ (.A(_00143_),
    .B(net2919),
    .Y(_03253_));
 sg13g2_o21ai_1 _08985_ (.B1(_03239_),
    .Y(_03254_),
    .A1(_03252_),
    .A2(_03253_));
 sg13g2_nor3_1 _08986_ (.A(_03239_),
    .B(_03252_),
    .C(_03253_),
    .Y(_03255_));
 sg13g2_or3_1 _08987_ (.A(_03239_),
    .B(_03252_),
    .C(_03253_),
    .X(_03256_));
 sg13g2_and2_1 _08988_ (.A(_03254_),
    .B(_03256_),
    .X(_03257_));
 sg13g2_xnor2_1 _08989_ (.Y(_03258_),
    .A(_03233_),
    .B(_03257_));
 sg13g2_a21oi_1 _08990_ (.A1(net2907),
    .A2(_03258_),
    .Y(_03259_),
    .B1(_03237_));
 sg13g2_a22oi_1 _08991_ (.Y(_03260_),
    .B1(net2766),
    .B2(_03259_),
    .A2(net2785),
    .A1(net374));
 sg13g2_inv_1 _08992_ (.Y(_00460_),
    .A(_03260_));
 sg13g2_o21ai_1 _08993_ (.B1(_03254_),
    .Y(_03261_),
    .A1(_03234_),
    .A2(_03255_));
 sg13g2_nand2_1 _08994_ (.Y(_03262_),
    .A(_00108_),
    .B(net3038));
 sg13g2_o21ai_1 _08995_ (.B1(_03262_),
    .Y(_03263_),
    .A1(_00642_),
    .A2(net3037));
 sg13g2_nand2_1 _08996_ (.Y(_03264_),
    .A(net3476),
    .B(\core.work.registers.genblk1[1].latch[2] ));
 sg13g2_nand2_1 _08997_ (.Y(_03265_),
    .A(\core.work.registers.genblk1[8].latch[2] ),
    .B(net3128));
 sg13g2_a21oi_1 _08998_ (.A1(\core.work.registers.genblk1[14].latch[2] ),
    .A2(net3103),
    .Y(_03266_),
    .B1(net3326));
 sg13g2_a22oi_1 _08999_ (.Y(_03267_),
    .B1(net3083),
    .B2(\core.work.registers.genblk1[5].latch[2] ),
    .A2(net3118),
    .A1(\core.work.registers.genblk1[4].latch[2] ));
 sg13g2_a22oi_1 _09000_ (.Y(_03268_),
    .B1(net3108),
    .B2(\core.work.registers.genblk1[6].latch[2] ),
    .A2(net3133),
    .A1(\core.work.registers.genblk1[10].latch[2] ));
 sg13g2_a22oi_1 _09001_ (.Y(_03269_),
    .B1(net3073),
    .B2(\core.work.registers.genblk1[15].latch[2] ),
    .A2(net3088),
    .A1(\core.work.registers.genblk1[3].latch[2] ));
 sg13g2_and4_1 _09002_ (.A(_03266_),
    .B(_03267_),
    .C(_03268_),
    .D(_03269_),
    .X(_03270_));
 sg13g2_a22oi_1 _09003_ (.Y(_03271_),
    .B1(net3094),
    .B2(\core.work.registers.genblk1[12].latch[2] ),
    .A2(net3123),
    .A1(\core.work.registers.genblk1[7].latch[2] ));
 sg13g2_a22oi_1 _09004_ (.Y(_03272_),
    .B1(net3068),
    .B2(\core.work.registers.genblk1[13].latch[2] ),
    .A2(net3098),
    .A1(\core.work.registers.genblk1[11].latch[2] ));
 sg13g2_a22oi_1 _09005_ (.Y(_03273_),
    .B1(net3078),
    .B2(\core.work.registers.genblk1[9].latch[2] ),
    .A2(net3114),
    .A1(\core.work.registers.genblk1[2].latch[2] ));
 sg13g2_and4_1 _09006_ (.A(_03265_),
    .B(_03271_),
    .C(_03272_),
    .D(_03273_),
    .X(_03274_));
 sg13g2_a22oi_1 _09007_ (.Y(_03275_),
    .B1(_03270_),
    .B2(_03274_),
    .A2(_03264_),
    .A1(net3325));
 sg13g2_nand2_1 _09008_ (.Y(_03276_),
    .A(net3556),
    .B(net2912));
 sg13g2_o21ai_1 _09009_ (.B1(_03276_),
    .Y(_03277_),
    .A1(_01688_),
    .A2(_03275_));
 sg13g2_nor2_1 _09010_ (.A(_03263_),
    .B(_03277_),
    .Y(_03278_));
 sg13g2_xor2_1 _09011_ (.B(_03277_),
    .A(_03263_),
    .X(_03279_));
 sg13g2_xnor2_1 _09012_ (.Y(_03280_),
    .A(_03261_),
    .B(_03279_));
 sg13g2_o21ai_1 _09013_ (.B1(net2766),
    .Y(_03281_),
    .A1(net2907),
    .A2(_01783_));
 sg13g2_a21oi_1 _09014_ (.A1(net2907),
    .A2(_03280_),
    .Y(_03282_),
    .B1(_03281_));
 sg13g2_a21o_1 _09015_ (.A2(net2785),
    .A1(net629),
    .B1(_03282_),
    .X(_00461_));
 sg13g2_nand2_1 _09016_ (.Y(_03283_),
    .A(net457),
    .B(net2785));
 sg13g2_a21oi_1 _09017_ (.A1(_03261_),
    .A2(_03279_),
    .Y(_03284_),
    .B1(_03278_));
 sg13g2_nand2_1 _09018_ (.Y(_03285_),
    .A(net3452),
    .B(net3035));
 sg13g2_o21ai_1 _09019_ (.B1(_03285_),
    .Y(_03286_),
    .A1(_00714_),
    .A2(net3035));
 sg13g2_nand2_1 _09020_ (.Y(_03287_),
    .A(net3477),
    .B(\core.work.registers.genblk1[1].latch[3] ));
 sg13g2_a22oi_1 _09021_ (.Y(_03288_),
    .B1(net3108),
    .B2(\core.work.registers.genblk1[6].latch[3] ),
    .A2(net3123),
    .A1(\core.work.registers.genblk1[7].latch[3] ));
 sg13g2_nand2_1 _09022_ (.Y(_03289_),
    .A(\core.work.registers.genblk1[8].latch[3] ),
    .B(net3128));
 sg13g2_a22oi_1 _09023_ (.Y(_03290_),
    .B1(net3093),
    .B2(\core.work.registers.genblk1[12].latch[3] ),
    .A2(net3113),
    .A1(\core.work.registers.genblk1[2].latch[3] ));
 sg13g2_a21oi_1 _09024_ (.A1(\core.work.registers.genblk1[3].latch[3] ),
    .A2(net3088),
    .Y(_03291_),
    .B1(net3325));
 sg13g2_a22oi_1 _09025_ (.Y(_03292_),
    .B1(net3079),
    .B2(\core.work.registers.genblk1[9].latch[3] ),
    .A2(net3103),
    .A1(\core.work.registers.genblk1[14].latch[3] ));
 sg13g2_nand3_1 _09026_ (.B(_03291_),
    .C(_03292_),
    .A(_03290_),
    .Y(_03293_));
 sg13g2_a221oi_1 _09027_ (.B2(\core.work.registers.genblk1[15].latch[3] ),
    .C1(_03293_),
    .B1(net3074),
    .A1(\core.work.registers.genblk1[11].latch[3] ),
    .Y(_03294_),
    .A2(net3099));
 sg13g2_a22oi_1 _09028_ (.Y(_03295_),
    .B1(net3084),
    .B2(\core.work.registers.genblk1[5].latch[3] ),
    .A2(net3134),
    .A1(\core.work.registers.genblk1[10].latch[3] ));
 sg13g2_nand3_1 _09029_ (.B(_03289_),
    .C(_03295_),
    .A(_03288_),
    .Y(_03296_));
 sg13g2_a221oi_1 _09030_ (.B2(\core.work.registers.genblk1[13].latch[3] ),
    .C1(_03296_),
    .B1(net3068),
    .A1(\core.work.registers.genblk1[4].latch[3] ),
    .Y(_03297_),
    .A2(net3119));
 sg13g2_a22oi_1 _09031_ (.Y(_03298_),
    .B1(_03294_),
    .B2(_03297_),
    .A2(_03287_),
    .A1(net3325));
 sg13g2_nor2_1 _09032_ (.A(net3551),
    .B(net2919),
    .Y(_03299_));
 sg13g2_a21oi_1 _09033_ (.A1(net2919),
    .A2(_03298_),
    .Y(_03300_),
    .B1(_03299_));
 sg13g2_or2_1 _09034_ (.X(_03301_),
    .B(_03300_),
    .A(_03286_));
 sg13g2_xnor2_1 _09035_ (.Y(_03302_),
    .A(_03286_),
    .B(_03300_));
 sg13g2_xor2_1 _09036_ (.B(_03302_),
    .A(_03284_),
    .X(_03303_));
 sg13g2_nor2_1 _09037_ (.A(net2906),
    .B(_01805_),
    .Y(_03304_));
 sg13g2_o21ai_1 _09038_ (.B1(net2766),
    .Y(_03305_),
    .A1(net2908),
    .A2(_03303_));
 sg13g2_o21ai_1 _09039_ (.B1(_03283_),
    .Y(_00462_),
    .A1(_03304_),
    .A2(_03305_));
 sg13g2_nand2_1 _09040_ (.Y(_03306_),
    .A(net463),
    .B(net2785));
 sg13g2_o21ai_1 _09041_ (.B1(_03301_),
    .Y(_03307_),
    .A1(_03284_),
    .A2(_03302_));
 sg13g2_nor2_1 _09042_ (.A(_00040_),
    .B(net3037),
    .Y(_03308_));
 sg13g2_a21oi_1 _09043_ (.A1(_00715_),
    .A2(net3037),
    .Y(_03309_),
    .B1(_03308_));
 sg13g2_nand2_1 _09044_ (.Y(_03310_),
    .A(net3477),
    .B(\core.work.registers.genblk1[1].latch[4] ));
 sg13g2_nand2_1 _09045_ (.Y(_03311_),
    .A(\core.work.registers.genblk1[8].latch[4] ),
    .B(net3128));
 sg13g2_a22oi_1 _09046_ (.Y(_03312_),
    .B1(net3074),
    .B2(\core.work.registers.genblk1[15].latch[4] ),
    .A2(net3094),
    .A1(\core.work.registers.genblk1[12].latch[4] ));
 sg13g2_a22oi_1 _09047_ (.Y(_03313_),
    .B1(net3089),
    .B2(\core.work.registers.genblk1[3].latch[4] ),
    .A2(net3114),
    .A1(\core.work.registers.genblk1[2].latch[4] ));
 sg13g2_a21oi_1 _09048_ (.A1(\core.work.registers.genblk1[7].latch[4] ),
    .A2(net3123),
    .Y(_03314_),
    .B1(net3325));
 sg13g2_a22oi_1 _09049_ (.Y(_03315_),
    .B1(net3079),
    .B2(\core.work.registers.genblk1[9].latch[4] ),
    .A2(net3134),
    .A1(\core.work.registers.genblk1[10].latch[4] ));
 sg13g2_and4_1 _09050_ (.A(_03312_),
    .B(_03313_),
    .C(_03314_),
    .D(_03315_),
    .X(_03316_));
 sg13g2_a22oi_1 _09051_ (.Y(_03317_),
    .B1(net3084),
    .B2(\core.work.registers.genblk1[5].latch[4] ),
    .A2(net3099),
    .A1(\core.work.registers.genblk1[11].latch[4] ));
 sg13g2_a22oi_1 _09052_ (.Y(_03318_),
    .B1(net3068),
    .B2(\core.work.registers.genblk1[13].latch[4] ),
    .A2(net3109),
    .A1(\core.work.registers.genblk1[6].latch[4] ));
 sg13g2_a22oi_1 _09053_ (.Y(_03319_),
    .B1(net3104),
    .B2(\core.work.registers.genblk1[14].latch[4] ),
    .A2(net3119),
    .A1(\core.work.registers.genblk1[4].latch[4] ));
 sg13g2_and4_1 _09054_ (.A(_03311_),
    .B(_03317_),
    .C(_03318_),
    .D(_03319_),
    .X(_03320_));
 sg13g2_a22oi_1 _09055_ (.Y(_03321_),
    .B1(_03316_),
    .B2(_03320_),
    .A2(_03310_),
    .A1(net3325));
 sg13g2_nor2_1 _09056_ (.A(_00054_),
    .B(net2920),
    .Y(_03322_));
 sg13g2_a21oi_2 _09057_ (.B1(_03322_),
    .Y(_03323_),
    .A2(_03321_),
    .A1(net2920));
 sg13g2_nor2_1 _09058_ (.A(_03309_),
    .B(_03323_),
    .Y(_03324_));
 sg13g2_xor2_1 _09059_ (.B(_03323_),
    .A(_03309_),
    .X(_03325_));
 sg13g2_xnor2_1 _09060_ (.Y(_03326_),
    .A(_03307_),
    .B(_03325_));
 sg13g2_and2_1 _09061_ (.A(net2905),
    .B(_03326_),
    .X(_03327_));
 sg13g2_o21ai_1 _09062_ (.B1(net2766),
    .Y(_03328_),
    .A1(net2905),
    .A2(_01828_));
 sg13g2_o21ai_1 _09063_ (.B1(_03306_),
    .Y(_00463_),
    .A1(_03327_),
    .A2(_03328_));
 sg13g2_nand2_1 _09064_ (.Y(_03329_),
    .A(net3474),
    .B(\core.work.registers.genblk1[1].latch[5] ));
 sg13g2_nand2_1 _09065_ (.Y(_03330_),
    .A(\core.work.registers.genblk1[4].latch[5] ),
    .B(net3117));
 sg13g2_a22oi_1 _09066_ (.Y(_03331_),
    .B1(net3067),
    .B2(\core.work.registers.genblk1[13].latch[5] ),
    .A2(net3082),
    .A1(\core.work.registers.genblk1[5].latch[5] ));
 sg13g2_a22oi_1 _09067_ (.Y(_03332_),
    .B1(net3092),
    .B2(\core.work.registers.genblk1[12].latch[5] ),
    .A2(net3097),
    .A1(\core.work.registers.genblk1[11].latch[5] ));
 sg13g2_a21oi_1 _09068_ (.A1(\core.work.registers.genblk1[6].latch[5] ),
    .A2(net3107),
    .Y(_03333_),
    .B1(net3322));
 sg13g2_a22oi_1 _09069_ (.Y(_03334_),
    .B1(net3087),
    .B2(\core.work.registers.genblk1[3].latch[5] ),
    .A2(net3127),
    .A1(\core.work.registers.genblk1[8].latch[5] ));
 sg13g2_and4_1 _09070_ (.A(_03331_),
    .B(_03332_),
    .C(_03333_),
    .D(_03334_),
    .X(_03335_));
 sg13g2_a22oi_1 _09071_ (.Y(_03336_),
    .B1(net3102),
    .B2(\core.work.registers.genblk1[14].latch[5] ),
    .A2(net3132),
    .A1(\core.work.registers.genblk1[10].latch[5] ));
 sg13g2_a22oi_1 _09072_ (.Y(_03337_),
    .B1(net3072),
    .B2(\core.work.registers.genblk1[15].latch[5] ),
    .A2(net3112),
    .A1(\core.work.registers.genblk1[2].latch[5] ));
 sg13g2_a22oi_1 _09073_ (.Y(_03338_),
    .B1(net3077),
    .B2(\core.work.registers.genblk1[9].latch[5] ),
    .A2(net3122),
    .A1(\core.work.registers.genblk1[7].latch[5] ));
 sg13g2_and4_1 _09074_ (.A(_03330_),
    .B(_03336_),
    .C(_03337_),
    .D(_03338_),
    .X(_03339_));
 sg13g2_a22oi_1 _09075_ (.Y(_03340_),
    .B1(_03335_),
    .B2(_03339_),
    .A2(_03329_),
    .A1(net3322));
 sg13g2_mux2_2 _09076_ (.A0(_00716_),
    .A1(_03340_),
    .S(net2919),
    .X(_03341_));
 sg13g2_or2_1 _09077_ (.X(_03342_),
    .B(_03341_),
    .A(net3449));
 sg13g2_and2_1 _09078_ (.A(net3450),
    .B(_03341_),
    .X(_03343_));
 sg13g2_xor2_1 _09079_ (.B(_03341_),
    .A(net3449),
    .X(_03344_));
 sg13g2_a21oi_1 _09080_ (.A1(_03307_),
    .A2(_03325_),
    .Y(_03345_),
    .B1(_03324_));
 sg13g2_xor2_1 _09081_ (.B(_03345_),
    .A(_03344_),
    .X(_03346_));
 sg13g2_o21ai_1 _09082_ (.B1(net2766),
    .Y(_03347_),
    .A1(net2905),
    .A2(_01852_));
 sg13g2_a21oi_1 _09083_ (.A1(net2905),
    .A2(_03346_),
    .Y(_03348_),
    .B1(_03347_));
 sg13g2_a21o_1 _09084_ (.A2(net2785),
    .A1(net546),
    .B1(_03348_),
    .X(_00464_));
 sg13g2_and2_1 _09085_ (.A(_03325_),
    .B(_03344_),
    .X(_03349_));
 sg13g2_nand2_1 _09086_ (.Y(_03350_),
    .A(_03307_),
    .B(_03349_));
 sg13g2_a21oi_1 _09087_ (.A1(_03324_),
    .A2(_03342_),
    .Y(_03351_),
    .B1(_03343_));
 sg13g2_nand2_1 _09088_ (.Y(_03352_),
    .A(_03350_),
    .B(_03351_));
 sg13g2_a21o_1 _09089_ (.A2(\core.work.registers.genblk1[1].latch[6] ),
    .A1(net3476),
    .B1(net3199),
    .X(_03353_));
 sg13g2_nand2_1 _09090_ (.Y(_03354_),
    .A(\core.work.registers.genblk1[6].latch[6] ),
    .B(net3109));
 sg13g2_a22oi_1 _09091_ (.Y(_03355_),
    .B1(net3089),
    .B2(\core.work.registers.genblk1[3].latch[6] ),
    .A2(net3124),
    .A1(\core.work.registers.genblk1[7].latch[6] ));
 sg13g2_a22oi_1 _09092_ (.Y(_03356_),
    .B1(net3084),
    .B2(\core.work.registers.genblk1[5].latch[6] ),
    .A2(net3119),
    .A1(\core.work.registers.genblk1[4].latch[6] ));
 sg13g2_a21oi_1 _09093_ (.A1(\core.work.registers.genblk1[14].latch[6] ),
    .A2(net3104),
    .Y(_03357_),
    .B1(net3326));
 sg13g2_a22oi_1 _09094_ (.Y(_03358_),
    .B1(net3074),
    .B2(\core.work.registers.genblk1[15].latch[6] ),
    .A2(net3079),
    .A1(\core.work.registers.genblk1[9].latch[6] ));
 sg13g2_a22oi_1 _09095_ (.Y(_03359_),
    .B1(net3128),
    .B2(\core.work.registers.genblk1[8].latch[6] ),
    .A2(net3134),
    .A1(\core.work.registers.genblk1[10].latch[6] ));
 sg13g2_a22oi_1 _09096_ (.Y(_03360_),
    .B1(net3094),
    .B2(\core.work.registers.genblk1[12].latch[6] ),
    .A2(net3114),
    .A1(\core.work.registers.genblk1[2].latch[6] ));
 sg13g2_nand4_1 _09097_ (.B(_03358_),
    .C(_03359_),
    .A(_03357_),
    .Y(_03361_),
    .D(_03360_));
 sg13g2_a22oi_1 _09098_ (.Y(_03362_),
    .B1(net3069),
    .B2(\core.work.registers.genblk1[13].latch[6] ),
    .A2(net3099),
    .A1(\core.work.registers.genblk1[11].latch[6] ));
 sg13g2_nand4_1 _09099_ (.B(_03355_),
    .C(_03356_),
    .A(_03354_),
    .Y(_03363_),
    .D(_03362_));
 sg13g2_o21ai_1 _09100_ (.B1(_03353_),
    .Y(_03364_),
    .A1(_03361_),
    .A2(_03363_));
 sg13g2_nor2_1 _09101_ (.A(_00717_),
    .B(net2919),
    .Y(_03365_));
 sg13g2_a21oi_2 _09102_ (.B1(_03365_),
    .Y(_03366_),
    .A2(_03364_),
    .A1(net2919));
 sg13g2_xnor2_1 _09103_ (.Y(_03367_),
    .A(_00613_),
    .B(_03366_));
 sg13g2_xnor2_1 _09104_ (.Y(_03368_),
    .A(_03352_),
    .B(_03367_));
 sg13g2_o21ai_1 _09105_ (.B1(net2766),
    .Y(_03369_),
    .A1(net2906),
    .A2(_01873_));
 sg13g2_a21oi_1 _09106_ (.A1(net2905),
    .A2(_03368_),
    .Y(_03370_),
    .B1(_03369_));
 sg13g2_a21o_1 _09107_ (.A2(net2785),
    .A1(net517),
    .B1(_03370_),
    .X(_00465_));
 sg13g2_nor2b_1 _09108_ (.A(_00044_),
    .B_N(_03366_),
    .Y(_03371_));
 sg13g2_a21oi_1 _09109_ (.A1(_03352_),
    .A2(_03367_),
    .Y(_03372_),
    .B1(_03371_));
 sg13g2_nand2_1 _09110_ (.Y(_03373_),
    .A(net3477),
    .B(\core.work.registers.genblk1[1].latch[7] ));
 sg13g2_a22oi_1 _09111_ (.Y(_03374_),
    .B1(net3074),
    .B2(\core.work.registers.genblk1[15].latch[7] ),
    .A2(net3078),
    .A1(\core.work.registers.genblk1[9].latch[7] ));
 sg13g2_a22oi_1 _09112_ (.Y(_03375_),
    .B1(net3083),
    .B2(\core.work.registers.genblk1[5].latch[7] ),
    .A2(net3088),
    .A1(\core.work.registers.genblk1[3].latch[7] ));
 sg13g2_a22oi_1 _09113_ (.Y(_03376_),
    .B1(net3118),
    .B2(\core.work.registers.genblk1[4].latch[7] ),
    .A2(net3133),
    .A1(\core.work.registers.genblk1[10].latch[7] ));
 sg13g2_nand2_1 _09114_ (.Y(_03377_),
    .A(\core.work.registers.genblk1[8].latch[7] ),
    .B(net3128));
 sg13g2_a22oi_1 _09115_ (.Y(_03378_),
    .B1(net3093),
    .B2(\core.work.registers.genblk1[12].latch[7] ),
    .A2(net3103),
    .A1(\core.work.registers.genblk1[14].latch[7] ));
 sg13g2_a21oi_1 _09116_ (.A1(\core.work.registers.genblk1[11].latch[7] ),
    .A2(net3099),
    .Y(_03379_),
    .B1(net3325));
 sg13g2_a22oi_1 _09117_ (.Y(_03380_),
    .B1(net3108),
    .B2(\core.work.registers.genblk1[6].latch[7] ),
    .A2(net3113),
    .A1(\core.work.registers.genblk1[2].latch[7] ));
 sg13g2_and4_1 _09118_ (.A(_03375_),
    .B(_03378_),
    .C(_03379_),
    .D(_03380_),
    .X(_03381_));
 sg13g2_a22oi_1 _09119_ (.Y(_03382_),
    .B1(net3068),
    .B2(\core.work.registers.genblk1[13].latch[7] ),
    .A2(net3123),
    .A1(\core.work.registers.genblk1[7].latch[7] ));
 sg13g2_and4_1 _09120_ (.A(_03374_),
    .B(_03376_),
    .C(_03377_),
    .D(_03382_),
    .X(_03383_));
 sg13g2_a22oi_1 _09121_ (.Y(_03384_),
    .B1(_03381_),
    .B2(_03383_),
    .A2(_03373_),
    .A1(net3325));
 sg13g2_mux2_1 _09122_ (.A0(_00718_),
    .A1(_03384_),
    .S(net2920),
    .X(_03385_));
 sg13g2_nand2b_1 _09123_ (.Y(_03386_),
    .B(_00611_),
    .A_N(_03385_));
 sg13g2_inv_1 _09124_ (.Y(_03387_),
    .A(_03386_));
 sg13g2_and2_1 _09125_ (.A(\core.e2m_addr[27] ),
    .B(_03385_),
    .X(_03388_));
 sg13g2_nor2_1 _09126_ (.A(_03387_),
    .B(_03388_),
    .Y(_03389_));
 sg13g2_xor2_1 _09127_ (.B(_03389_),
    .A(_03372_),
    .X(_03390_));
 sg13g2_o21ai_1 _09128_ (.B1(net2766),
    .Y(_03391_),
    .A1(net2905),
    .A2(_01894_));
 sg13g2_a21oi_1 _09129_ (.A1(net2905),
    .A2(_03390_),
    .Y(_03392_),
    .B1(_03391_));
 sg13g2_a21o_1 _09130_ (.A2(net2785),
    .A1(net454),
    .B1(_03392_),
    .X(_00466_));
 sg13g2_a21oi_1 _09131_ (.A1(_03371_),
    .A2(_03386_),
    .Y(_03393_),
    .B1(_03388_));
 sg13g2_nand2_1 _09132_ (.Y(_03394_),
    .A(_03367_),
    .B(_03386_));
 sg13g2_and2_1 _09133_ (.A(_03393_),
    .B(_03394_),
    .X(_03395_));
 sg13g2_nand2_1 _09134_ (.Y(_03396_),
    .A(_03351_),
    .B(_03393_));
 sg13g2_a21oi_2 _09135_ (.B1(_03396_),
    .Y(_03397_),
    .A2(_03349_),
    .A1(_03307_));
 sg13g2_or2_1 _09136_ (.X(_03398_),
    .B(_03397_),
    .A(_03395_));
 sg13g2_a21oi_1 _09137_ (.A1(net3474),
    .A2(\core.work.registers.genblk1[1].latch[8] ),
    .Y(_03399_),
    .B1(net3199));
 sg13g2_nand2_1 _09138_ (.Y(_03400_),
    .A(\core.work.registers.genblk1[10].latch[8] ),
    .B(net3132));
 sg13g2_a22oi_1 _09139_ (.Y(_03401_),
    .B1(net3072),
    .B2(\core.work.registers.genblk1[15].latch[8] ),
    .A2(net3120),
    .A1(\core.work.registers.genblk1[4].latch[8] ));
 sg13g2_a22oi_1 _09140_ (.Y(_03402_),
    .B1(net3080),
    .B2(\core.work.registers.genblk1[9].latch[8] ),
    .A2(net3087),
    .A1(\core.work.registers.genblk1[3].latch[8] ));
 sg13g2_a21oi_1 _09141_ (.A1(\core.work.registers.genblk1[8].latch[8] ),
    .A2(net3127),
    .Y(_03403_),
    .B1(net3322));
 sg13g2_a22oi_1 _09142_ (.Y(_03404_),
    .B1(net3100),
    .B2(\core.work.registers.genblk1[11].latch[8] ),
    .A2(net3115),
    .A1(\core.work.registers.genblk1[2].latch[8] ));
 sg13g2_a22oi_1 _09143_ (.Y(_03405_),
    .B1(net3067),
    .B2(\core.work.registers.genblk1[13].latch[8] ),
    .A2(net3082),
    .A1(\core.work.registers.genblk1[5].latch[8] ));
 sg13g2_nand4_1 _09144_ (.B(_03403_),
    .C(_03404_),
    .A(_03402_),
    .Y(_03406_),
    .D(_03405_));
 sg13g2_a22oi_1 _09145_ (.Y(_03407_),
    .B1(net3093),
    .B2(\core.work.registers.genblk1[12].latch[8] ),
    .A2(net3102),
    .A1(\core.work.registers.genblk1[14].latch[8] ));
 sg13g2_a22oi_1 _09146_ (.Y(_03408_),
    .B1(net3107),
    .B2(\core.work.registers.genblk1[6].latch[8] ),
    .A2(net3122),
    .A1(\core.work.registers.genblk1[7].latch[8] ));
 sg13g2_nand4_1 _09147_ (.B(_03401_),
    .C(_03407_),
    .A(_03400_),
    .Y(_03409_),
    .D(_03408_));
 sg13g2_nor2_1 _09148_ (.A(_03406_),
    .B(_03409_),
    .Y(_03410_));
 sg13g2_nor2_2 _09149_ (.A(_03399_),
    .B(_03410_),
    .Y(_03411_));
 sg13g2_nor2_1 _09150_ (.A(_00115_),
    .B(net2918),
    .Y(_03412_));
 sg13g2_a21oi_1 _09151_ (.A1(net2921),
    .A2(_03411_),
    .Y(_03413_),
    .B1(_03412_));
 sg13g2_xnor2_1 _09152_ (.Y(_03414_),
    .A(\core.e2m_addr[28] ),
    .B(_03413_));
 sg13g2_nor2b_1 _09153_ (.A(_03398_),
    .B_N(_03414_),
    .Y(_03415_));
 sg13g2_xor2_1 _09154_ (.B(_03414_),
    .A(_03398_),
    .X(_03416_));
 sg13g2_o21ai_1 _09155_ (.B1(net2765),
    .Y(_03417_),
    .A1(net2903),
    .A2(_01913_));
 sg13g2_a21oi_1 _09156_ (.A1(net2903),
    .A2(_03416_),
    .Y(_03418_),
    .B1(_03417_));
 sg13g2_a21o_1 _09157_ (.A2(net2782),
    .A1(net560),
    .B1(_03418_),
    .X(_00467_));
 sg13g2_nand2_1 _09158_ (.Y(_03419_),
    .A(_00116_),
    .B(net2912));
 sg13g2_a21oi_1 _09159_ (.A1(net3479),
    .A2(\core.work.registers.genblk1[1].latch[9] ),
    .Y(_03420_),
    .B1(net3199));
 sg13g2_nand2_1 _09160_ (.Y(_03421_),
    .A(\core.work.registers.genblk1[10].latch[9] ),
    .B(net3133));
 sg13g2_a22oi_1 _09161_ (.Y(_03422_),
    .B1(net3093),
    .B2(\core.work.registers.genblk1[12].latch[9] ),
    .A2(net3108),
    .A1(\core.work.registers.genblk1[6].latch[9] ));
 sg13g2_a21oi_1 _09162_ (.A1(\core.work.registers.genblk1[14].latch[9] ),
    .A2(net3103),
    .Y(_03423_),
    .B1(net3328));
 sg13g2_a22oi_1 _09163_ (.Y(_03424_),
    .B1(net3073),
    .B2(\core.work.registers.genblk1[15].latch[9] ),
    .A2(net3129),
    .A1(\core.work.registers.genblk1[8].latch[9] ));
 sg13g2_a22oi_1 _09164_ (.Y(_03425_),
    .B1(net3078),
    .B2(\core.work.registers.genblk1[9].latch[9] ),
    .A2(net3113),
    .A1(\core.work.registers.genblk1[2].latch[9] ));
 sg13g2_nand4_1 _09165_ (.B(_03423_),
    .C(_03424_),
    .A(_03422_),
    .Y(_03426_),
    .D(_03425_));
 sg13g2_a22oi_1 _09166_ (.Y(_03427_),
    .B1(net3088),
    .B2(\core.work.registers.genblk1[3].latch[9] ),
    .A2(net3098),
    .A1(\core.work.registers.genblk1[11].latch[9] ));
 sg13g2_a22oi_1 _09167_ (.Y(_03428_),
    .B1(net3069),
    .B2(\core.work.registers.genblk1[13].latch[9] ),
    .A2(net3118),
    .A1(\core.work.registers.genblk1[4].latch[9] ));
 sg13g2_a22oi_1 _09168_ (.Y(_03429_),
    .B1(net3083),
    .B2(\core.work.registers.genblk1[5].latch[9] ),
    .A2(net3124),
    .A1(\core.work.registers.genblk1[7].latch[9] ));
 sg13g2_nand4_1 _09169_ (.B(_03427_),
    .C(_03428_),
    .A(_03421_),
    .Y(_03430_),
    .D(_03429_));
 sg13g2_nor2_1 _09170_ (.A(_03426_),
    .B(_03430_),
    .Y(_03431_));
 sg13g2_nor2_2 _09171_ (.A(_03420_),
    .B(_03431_),
    .Y(_03432_));
 sg13g2_nand2b_1 _09172_ (.Y(_03433_),
    .B(net2918),
    .A_N(_03432_));
 sg13g2_a21oi_1 _09173_ (.A1(_03419_),
    .A2(_03433_),
    .Y(_03434_),
    .B1(net3445));
 sg13g2_a21o_1 _09174_ (.A2(_03433_),
    .A1(_03419_),
    .B1(net3445),
    .X(_03435_));
 sg13g2_and3_1 _09175_ (.X(_03436_),
    .A(net3445),
    .B(_03419_),
    .C(_03433_));
 sg13g2_inv_1 _09176_ (.Y(_03437_),
    .A(_03436_));
 sg13g2_nor2_1 _09177_ (.A(_03434_),
    .B(_03436_),
    .Y(_03438_));
 sg13g2_nor2_1 _09178_ (.A(_00048_),
    .B(_03413_),
    .Y(_03439_));
 sg13g2_nor2_1 _09179_ (.A(_03415_),
    .B(_03439_),
    .Y(_03440_));
 sg13g2_xor2_1 _09180_ (.B(_03440_),
    .A(_03438_),
    .X(_03441_));
 sg13g2_o21ai_1 _09181_ (.B1(net2765),
    .Y(_03442_),
    .A1(net2903),
    .A2(_01932_));
 sg13g2_a21oi_1 _09182_ (.A1(net2903),
    .A2(_03441_),
    .Y(_03443_),
    .B1(_03442_));
 sg13g2_a21o_1 _09183_ (.A2(net2781),
    .A1(net635),
    .B1(_03443_),
    .X(_00468_));
 sg13g2_a21oi_1 _09184_ (.A1(_03437_),
    .A2(_03440_),
    .Y(_03444_),
    .B1(_03434_));
 sg13g2_nand2_1 _09185_ (.Y(_03445_),
    .A(net3474),
    .B(\core.work.registers.genblk1[1].latch[10] ));
 sg13g2_nand2_1 _09186_ (.Y(_03446_),
    .A(\core.work.registers.genblk1[12].latch[10] ),
    .B(net3095));
 sg13g2_a21oi_1 _09187_ (.A1(\core.work.registers.genblk1[13].latch[10] ),
    .A2(net3070),
    .Y(_03447_),
    .B1(net3323));
 sg13g2_a22oi_1 _09188_ (.Y(_03448_),
    .B1(net3115),
    .B2(\core.work.registers.genblk1[2].latch[10] ),
    .A2(net3130),
    .A1(\core.work.registers.genblk1[8].latch[10] ));
 sg13g2_a22oi_1 _09189_ (.Y(_03449_),
    .B1(net3075),
    .B2(\core.work.registers.genblk1[15].latch[10] ),
    .A2(net3100),
    .A1(\core.work.registers.genblk1[11].latch[10] ));
 sg13g2_nand3_1 _09190_ (.B(_03448_),
    .C(_03449_),
    .A(_03447_),
    .Y(_03450_));
 sg13g2_a221oi_1 _09191_ (.B2(\core.work.registers.genblk1[3].latch[10] ),
    .C1(_03450_),
    .B1(net3090),
    .A1(\core.work.registers.genblk1[4].latch[10] ),
    .Y(_03451_),
    .A2(net3120));
 sg13g2_a22oi_1 _09192_ (.Y(_03452_),
    .B1(net3110),
    .B2(\core.work.registers.genblk1[6].latch[10] ),
    .A2(net3125),
    .A1(\core.work.registers.genblk1[7].latch[10] ));
 sg13g2_a22oi_1 _09193_ (.Y(_03453_),
    .B1(net3080),
    .B2(\core.work.registers.genblk1[9].latch[10] ),
    .A2(net3085),
    .A1(\core.work.registers.genblk1[5].latch[10] ));
 sg13g2_nand3_1 _09194_ (.B(_03452_),
    .C(_03453_),
    .A(_03446_),
    .Y(_03454_));
 sg13g2_a221oi_1 _09195_ (.B2(\core.work.registers.genblk1[14].latch[10] ),
    .C1(_03454_),
    .B1(net3105),
    .A1(\core.work.registers.genblk1[10].latch[10] ),
    .Y(_03455_),
    .A2(net3135));
 sg13g2_a22oi_1 _09196_ (.Y(_03456_),
    .B1(_03451_),
    .B2(_03455_),
    .A2(_03445_),
    .A1(net3323));
 sg13g2_nor2_1 _09197_ (.A(_00117_),
    .B(net2918),
    .Y(_03457_));
 sg13g2_a21oi_1 _09198_ (.A1(net2918),
    .A2(_03456_),
    .Y(_03458_),
    .B1(_03457_));
 sg13g2_xnor2_1 _09199_ (.Y(_03459_),
    .A(\core.e2m_addr[30] ),
    .B(_03458_));
 sg13g2_xnor2_1 _09200_ (.Y(_03460_),
    .A(_03444_),
    .B(_03459_));
 sg13g2_o21ai_1 _09201_ (.B1(net2765),
    .Y(_03461_),
    .A1(net2903),
    .A2(_01952_));
 sg13g2_a21oi_1 _09202_ (.A1(net2904),
    .A2(_03460_),
    .Y(_03462_),
    .B1(_03461_));
 sg13g2_a21o_1 _09203_ (.A2(net2781),
    .A1(net542),
    .B1(_03462_),
    .X(_00469_));
 sg13g2_and2_2 _09204_ (.A(net3496),
    .B(_01685_),
    .X(_03463_));
 sg13g2_nor2_1 _09205_ (.A(net3361),
    .B(net2861),
    .Y(_03464_));
 sg13g2_a21oi_1 _09206_ (.A1(net3460),
    .A2(_03463_),
    .Y(_03465_),
    .B1(_03464_));
 sg13g2_nor2_1 _09207_ (.A(_00154_),
    .B(net3035),
    .Y(_03466_));
 sg13g2_a21oi_1 _09208_ (.A1(net3034),
    .A2(_03465_),
    .Y(_03467_),
    .B1(_03466_));
 sg13g2_nand2_1 _09209_ (.Y(_03468_),
    .A(net3473),
    .B(\core.work.registers.genblk1[1].latch[11] ));
 sg13g2_nand2_1 _09210_ (.Y(_03469_),
    .A(\core.work.registers.genblk1[14].latch[11] ),
    .B(net3102));
 sg13g2_a22oi_1 _09211_ (.Y(_03470_),
    .B1(net3082),
    .B2(\core.work.registers.genblk1[5].latch[11] ),
    .A2(net3107),
    .A1(\core.work.registers.genblk1[6].latch[11] ));
 sg13g2_a21oi_1 _09212_ (.A1(\core.work.registers.genblk1[10].latch[11] ),
    .A2(net3131),
    .Y(_03471_),
    .B1(net3324));
 sg13g2_a22oi_1 _09213_ (.Y(_03472_),
    .B1(net3076),
    .B2(\core.work.registers.genblk1[9].latch[11] ),
    .A2(net3121),
    .A1(\core.work.registers.genblk1[7].latch[11] ));
 sg13g2_a22oi_1 _09214_ (.Y(_03473_),
    .B1(net3116),
    .B2(\core.work.registers.genblk1[4].latch[11] ),
    .A2(net3126),
    .A1(\core.work.registers.genblk1[8].latch[11] ));
 sg13g2_nand3_1 _09215_ (.B(_03472_),
    .C(_03473_),
    .A(_03471_),
    .Y(_03474_));
 sg13g2_a221oi_1 _09216_ (.B2(\core.work.registers.genblk1[3].latch[11] ),
    .C1(_03474_),
    .B1(net3087),
    .A1(\core.work.registers.genblk1[2].latch[11] ),
    .Y(_03475_),
    .A2(net3112));
 sg13g2_a22oi_1 _09217_ (.Y(_03476_),
    .B1(net3067),
    .B2(\core.work.registers.genblk1[13].latch[11] ),
    .A2(net3097),
    .A1(\core.work.registers.genblk1[11].latch[11] ));
 sg13g2_nand3_1 _09218_ (.B(_03470_),
    .C(_03476_),
    .A(_03469_),
    .Y(_03477_));
 sg13g2_a221oi_1 _09219_ (.B2(\core.work.registers.genblk1[15].latch[11] ),
    .C1(_03477_),
    .B1(net3072),
    .A1(\core.work.registers.genblk1[12].latch[11] ),
    .Y(_03478_),
    .A2(net3092));
 sg13g2_a22oi_1 _09220_ (.Y(_03479_),
    .B1(_03475_),
    .B2(_03478_),
    .A2(_03468_),
    .A1(net3324));
 sg13g2_nand2_1 _09221_ (.Y(_03480_),
    .A(net2918),
    .B(_03479_));
 sg13g2_o21ai_1 _09222_ (.B1(_03480_),
    .Y(_03481_),
    .A1(_00118_),
    .A2(net2918));
 sg13g2_nand2b_1 _09223_ (.Y(_03482_),
    .B(_03467_),
    .A_N(_03481_));
 sg13g2_nand2b_1 _09224_ (.Y(_03483_),
    .B(_03481_),
    .A_N(_03467_));
 sg13g2_xnor2_1 _09225_ (.Y(_03484_),
    .A(_03467_),
    .B(_03481_));
 sg13g2_nor2_1 _09226_ (.A(_00052_),
    .B(_03458_),
    .Y(_03485_));
 sg13g2_a21oi_1 _09227_ (.A1(_03444_),
    .A2(_03459_),
    .Y(_03486_),
    .B1(_03485_));
 sg13g2_xor2_1 _09228_ (.B(_03486_),
    .A(_03484_),
    .X(_03487_));
 sg13g2_o21ai_1 _09229_ (.B1(net2765),
    .Y(_03488_),
    .A1(net2903),
    .A2(_01972_));
 sg13g2_a21oi_1 _09230_ (.A1(net2904),
    .A2(_03487_),
    .Y(_03489_),
    .B1(_03488_));
 sg13g2_a21o_1 _09231_ (.A2(net2781),
    .A1(net619),
    .B1(_03489_),
    .X(_00470_));
 sg13g2_nand4_1 _09232_ (.B(_03438_),
    .C(_03459_),
    .A(_03414_),
    .Y(_03490_),
    .D(_03484_));
 sg13g2_nor3_2 _09233_ (.A(_03395_),
    .B(_03397_),
    .C(_03490_),
    .Y(_03491_));
 sg13g2_a21o_1 _09234_ (.A2(_03439_),
    .A1(_03435_),
    .B1(_03436_),
    .X(_03492_));
 sg13g2_nand3_1 _09235_ (.B(_03484_),
    .C(_03492_),
    .A(_03459_),
    .Y(_03493_));
 sg13g2_nand2_1 _09236_ (.Y(_03494_),
    .A(_03482_),
    .B(_03485_));
 sg13g2_nand3_1 _09237_ (.B(_03493_),
    .C(_03494_),
    .A(_03483_),
    .Y(_03495_));
 sg13g2_or2_1 _09238_ (.X(_03496_),
    .B(_03495_),
    .A(_03491_));
 sg13g2_a21o_1 _09239_ (.A2(net2861),
    .A1(_00120_),
    .B1(net2836),
    .X(_03497_));
 sg13g2_a21oi_1 _09240_ (.A1(net3474),
    .A2(\core.work.registers.genblk1[1].latch[12] ),
    .Y(_03498_),
    .B1(net3199));
 sg13g2_a22oi_1 _09241_ (.Y(_03499_),
    .B1(net3070),
    .B2(\core.work.registers.genblk1[13].latch[12] ),
    .A2(net3075),
    .A1(\core.work.registers.genblk1[15].latch[12] ));
 sg13g2_nand2_1 _09242_ (.Y(_03500_),
    .A(\core.work.registers.genblk1[12].latch[12] ),
    .B(net3092));
 sg13g2_a22oi_1 _09243_ (.Y(_03501_),
    .B1(net3085),
    .B2(\core.work.registers.genblk1[5].latch[12] ),
    .A2(net3112),
    .A1(\core.work.registers.genblk1[2].latch[12] ));
 sg13g2_a22oi_1 _09244_ (.Y(_03502_),
    .B1(net3090),
    .B2(\core.work.registers.genblk1[3].latch[12] ),
    .A2(net3117),
    .A1(\core.work.registers.genblk1[4].latch[12] ));
 sg13g2_a21oi_1 _09245_ (.A1(\core.work.registers.genblk1[11].latch[12] ),
    .A2(net3097),
    .Y(_03503_),
    .B1(net3322));
 sg13g2_a22oi_1 _09246_ (.Y(_03504_),
    .B1(net3077),
    .B2(\core.work.registers.genblk1[9].latch[12] ),
    .A2(net3135),
    .A1(\core.work.registers.genblk1[10].latch[12] ));
 sg13g2_nand4_1 _09247_ (.B(_03502_),
    .C(_03503_),
    .A(_03499_),
    .Y(_03505_),
    .D(_03504_));
 sg13g2_a22oi_1 _09248_ (.Y(_03506_),
    .B1(net3125),
    .B2(\core.work.registers.genblk1[7].latch[12] ),
    .A2(net3130),
    .A1(\core.work.registers.genblk1[8].latch[12] ));
 sg13g2_a22oi_1 _09249_ (.Y(_03507_),
    .B1(net3105),
    .B2(\core.work.registers.genblk1[14].latch[12] ),
    .A2(net3107),
    .A1(\core.work.registers.genblk1[6].latch[12] ));
 sg13g2_nand4_1 _09250_ (.B(_03501_),
    .C(_03506_),
    .A(_03500_),
    .Y(_03508_),
    .D(_03507_));
 sg13g2_nor2_1 _09251_ (.A(_03505_),
    .B(_03508_),
    .Y(_03509_));
 sg13g2_nor2_2 _09252_ (.A(_03498_),
    .B(_03509_),
    .Y(_03510_));
 sg13g2_nand2_1 _09253_ (.Y(_03511_),
    .A(net2916),
    .B(_03510_));
 sg13g2_o21ai_1 _09254_ (.B1(_03511_),
    .Y(_03512_),
    .A1(_00119_),
    .A2(net2916));
 sg13g2_nor2b_1 _09255_ (.A(_03497_),
    .B_N(_03512_),
    .Y(_03513_));
 sg13g2_xor2_1 _09256_ (.B(_03512_),
    .A(_03497_),
    .X(_03514_));
 sg13g2_nor2b_1 _09257_ (.A(_03514_),
    .B_N(_03496_),
    .Y(_03515_));
 sg13g2_xor2_1 _09258_ (.B(_03514_),
    .A(_03496_),
    .X(_03516_));
 sg13g2_o21ai_1 _09259_ (.B1(net2764),
    .Y(_03517_),
    .A1(net2901),
    .A2(_01991_));
 sg13g2_a21oi_2 _09260_ (.B1(_03517_),
    .Y(_03518_),
    .A2(_03516_),
    .A1(net2901));
 sg13g2_a21o_1 _09261_ (.A2(net2781),
    .A1(net521),
    .B1(_03518_),
    .X(_00471_));
 sg13g2_a21o_1 _09262_ (.A2(net2861),
    .A1(_00122_),
    .B1(net2836),
    .X(_03519_));
 sg13g2_a21oi_1 _09263_ (.A1(net3474),
    .A2(\core.work.registers.genblk1[1].latch[13] ),
    .Y(_03520_),
    .B1(net3198));
 sg13g2_nand2_1 _09264_ (.Y(_03521_),
    .A(\core.work.registers.genblk1[6].latch[13] ),
    .B(net3110));
 sg13g2_a22oi_1 _09265_ (.Y(_03522_),
    .B1(net3067),
    .B2(\core.work.registers.genblk1[13].latch[13] ),
    .A2(net3122),
    .A1(\core.work.registers.genblk1[7].latch[13] ));
 sg13g2_a22oi_1 _09266_ (.Y(_03523_),
    .B1(net3087),
    .B2(\core.work.registers.genblk1[3].latch[13] ),
    .A2(net3112),
    .A1(\core.work.registers.genblk1[2].latch[13] ));
 sg13g2_a21oi_1 _09267_ (.A1(\core.work.registers.genblk1[12].latch[13] ),
    .A2(net3092),
    .Y(_03524_),
    .B1(net3322));
 sg13g2_a22oi_1 _09268_ (.Y(_03525_),
    .B1(net3072),
    .B2(\core.work.registers.genblk1[15].latch[13] ),
    .A2(net3097),
    .A1(\core.work.registers.genblk1[11].latch[13] ));
 sg13g2_a22oi_1 _09269_ (.Y(_03526_),
    .B1(net3117),
    .B2(\core.work.registers.genblk1[4].latch[13] ),
    .A2(net3127),
    .A1(\core.work.registers.genblk1[8].latch[13] ));
 sg13g2_nand4_1 _09270_ (.B(_03524_),
    .C(_03525_),
    .A(_03523_),
    .Y(_03527_),
    .D(_03526_));
 sg13g2_a22oi_1 _09271_ (.Y(_03528_),
    .B1(net3077),
    .B2(\core.work.registers.genblk1[9].latch[13] ),
    .A2(net3082),
    .A1(\core.work.registers.genblk1[5].latch[13] ));
 sg13g2_a22oi_1 _09272_ (.Y(_03529_),
    .B1(net3102),
    .B2(\core.work.registers.genblk1[14].latch[13] ),
    .A2(net3132),
    .A1(\core.work.registers.genblk1[10].latch[13] ));
 sg13g2_nand4_1 _09273_ (.B(_03522_),
    .C(_03528_),
    .A(_03521_),
    .Y(_03530_),
    .D(_03529_));
 sg13g2_nor2_2 _09274_ (.A(_03527_),
    .B(_03530_),
    .Y(_03531_));
 sg13g2_nor2_2 _09275_ (.A(_03520_),
    .B(_03531_),
    .Y(_03532_));
 sg13g2_nand2_1 _09276_ (.Y(_03533_),
    .A(net2915),
    .B(_03532_));
 sg13g2_nand2b_1 _09277_ (.Y(_03534_),
    .B(net2912),
    .A_N(_00121_));
 sg13g2_and3_1 _09278_ (.X(_03535_),
    .A(_03519_),
    .B(_03533_),
    .C(_03534_));
 sg13g2_nand3_1 _09279_ (.B(_03533_),
    .C(_03534_),
    .A(_03519_),
    .Y(_03536_));
 sg13g2_a21oi_1 _09280_ (.A1(_03533_),
    .A2(_03534_),
    .Y(_03537_),
    .B1(_03519_));
 sg13g2_or2_1 _09281_ (.X(_03538_),
    .B(_03537_),
    .A(_03535_));
 sg13g2_nor2_1 _09282_ (.A(_03513_),
    .B(_03515_),
    .Y(_03539_));
 sg13g2_xnor2_1 _09283_ (.Y(_03540_),
    .A(_03538_),
    .B(_03539_));
 sg13g2_o21ai_1 _09284_ (.B1(net2763),
    .Y(_03541_),
    .A1(net2899),
    .A2(_02015_));
 sg13g2_a21oi_2 _09285_ (.B1(_03541_),
    .Y(_03542_),
    .A2(_03540_),
    .A1(net2899));
 sg13g2_a21o_1 _09286_ (.A2(net2783),
    .A1(net597),
    .B1(_03542_),
    .X(_00472_));
 sg13g2_a21oi_1 _09287_ (.A1(_00124_),
    .A2(net2861),
    .Y(_03543_),
    .B1(net2836));
 sg13g2_a21oi_1 _09288_ (.A1(net3474),
    .A2(\core.work.registers.genblk1[1].latch[14] ),
    .Y(_03544_),
    .B1(net3198));
 sg13g2_a21oi_1 _09289_ (.A1(\core.work.registers.genblk1[14].latch[14] ),
    .A2(net3105),
    .Y(_03545_),
    .B1(net3323));
 sg13g2_nand2_1 _09290_ (.Y(_03546_),
    .A(\core.work.registers.genblk1[7].latch[14] ),
    .B(net3125));
 sg13g2_a22oi_1 _09291_ (.Y(_03547_),
    .B1(net3090),
    .B2(\core.work.registers.genblk1[3].latch[14] ),
    .A2(net3095),
    .A1(\core.work.registers.genblk1[12].latch[14] ));
 sg13g2_a22oi_1 _09292_ (.Y(_03548_),
    .B1(net3075),
    .B2(\core.work.registers.genblk1[15].latch[14] ),
    .A2(net3110),
    .A1(\core.work.registers.genblk1[6].latch[14] ));
 sg13g2_a22oi_1 _09293_ (.Y(_03549_),
    .B1(net3070),
    .B2(\core.work.registers.genblk1[13].latch[14] ),
    .A2(net3120),
    .A1(\core.work.registers.genblk1[4].latch[14] ));
 sg13g2_a22oi_1 _09294_ (.Y(_03550_),
    .B1(net3080),
    .B2(\core.work.registers.genblk1[9].latch[14] ),
    .A2(net3085),
    .A1(\core.work.registers.genblk1[5].latch[14] ));
 sg13g2_a22oi_1 _09295_ (.Y(_03551_),
    .B1(net3130),
    .B2(\core.work.registers.genblk1[8].latch[14] ),
    .A2(net3135),
    .A1(\core.work.registers.genblk1[10].latch[14] ));
 sg13g2_nand4_1 _09296_ (.B(_03549_),
    .C(_03550_),
    .A(_03545_),
    .Y(_03552_),
    .D(_03551_));
 sg13g2_a22oi_1 _09297_ (.Y(_03553_),
    .B1(net3100),
    .B2(\core.work.registers.genblk1[11].latch[14] ),
    .A2(net3115),
    .A1(\core.work.registers.genblk1[2].latch[14] ));
 sg13g2_nand4_1 _09298_ (.B(_03547_),
    .C(_03548_),
    .A(_03546_),
    .Y(_03554_),
    .D(_03553_));
 sg13g2_nor2_1 _09299_ (.A(_03552_),
    .B(_03554_),
    .Y(_03555_));
 sg13g2_nor2_2 _09300_ (.A(_03544_),
    .B(_03555_),
    .Y(_03556_));
 sg13g2_nand2_1 _09301_ (.Y(_03557_),
    .A(net2916),
    .B(_03556_));
 sg13g2_o21ai_1 _09302_ (.B1(_03557_),
    .Y(_03558_),
    .A1(_00123_),
    .A2(net2916));
 sg13g2_and2_1 _09303_ (.A(_03543_),
    .B(_03558_),
    .X(_03559_));
 sg13g2_inv_1 _09304_ (.Y(_03560_),
    .A(_03559_));
 sg13g2_xnor2_1 _09305_ (.Y(_03561_),
    .A(_03543_),
    .B(_03558_));
 sg13g2_a21o_1 _09306_ (.A2(_03536_),
    .A1(_03513_),
    .B1(_03537_),
    .X(_03562_));
 sg13g2_nor2_1 _09307_ (.A(_03514_),
    .B(_03538_),
    .Y(_03563_));
 sg13g2_a21oi_1 _09308_ (.A1(_03496_),
    .A2(_03563_),
    .Y(_03564_),
    .B1(_03562_));
 sg13g2_xnor2_1 _09309_ (.Y(_03565_),
    .A(_03561_),
    .B(_03564_));
 sg13g2_o21ai_1 _09310_ (.B1(net2763),
    .Y(_03566_),
    .A1(net2902),
    .A2(_02036_));
 sg13g2_a21oi_2 _09311_ (.B1(_03566_),
    .Y(_03567_),
    .A2(_03565_),
    .A1(net2899));
 sg13g2_a21o_1 _09312_ (.A2(net2783),
    .A1(net644),
    .B1(_03567_),
    .X(_00473_));
 sg13g2_a21o_1 _09313_ (.A2(net2861),
    .A1(_00126_),
    .B1(net2836),
    .X(_03568_));
 sg13g2_nand2_1 _09314_ (.Y(_03569_),
    .A(_00125_),
    .B(net2912));
 sg13g2_a21oi_1 _09315_ (.A1(net3473),
    .A2(\core.work.registers.genblk1[1].latch[15] ),
    .Y(_03570_),
    .B1(net3197));
 sg13g2_nand2_1 _09316_ (.Y(_03571_),
    .A(\core.work.registers.genblk1[10].latch[15] ),
    .B(net3132));
 sg13g2_a22oi_1 _09317_ (.Y(_03572_),
    .B1(net3081),
    .B2(\core.work.registers.genblk1[5].latch[15] ),
    .A2(net3127),
    .A1(\core.work.registers.genblk1[8].latch[15] ));
 sg13g2_a21oi_1 _09318_ (.A1(\core.work.registers.genblk1[9].latch[15] ),
    .A2(net3076),
    .Y(_03573_),
    .B1(net3321));
 sg13g2_a22oi_1 _09319_ (.Y(_03574_),
    .B1(net3091),
    .B2(\core.work.registers.genblk1[12].latch[15] ),
    .A2(net3096),
    .A1(\core.work.registers.genblk1[11].latch[15] ));
 sg13g2_a22oi_1 _09320_ (.Y(_03575_),
    .B1(net3071),
    .B2(\core.work.registers.genblk1[15].latch[15] ),
    .A2(net3122),
    .A1(\core.work.registers.genblk1[7].latch[15] ));
 sg13g2_nand4_1 _09321_ (.B(_03573_),
    .C(_03574_),
    .A(_03572_),
    .Y(_03576_),
    .D(_03575_));
 sg13g2_a22oi_1 _09322_ (.Y(_03577_),
    .B1(net3101),
    .B2(\core.work.registers.genblk1[14].latch[15] ),
    .A2(net3111),
    .A1(\core.work.registers.genblk1[2].latch[15] ));
 sg13g2_a22oi_1 _09323_ (.Y(_03578_),
    .B1(net3086),
    .B2(\core.work.registers.genblk1[3].latch[15] ),
    .A2(net3106),
    .A1(\core.work.registers.genblk1[6].latch[15] ));
 sg13g2_a22oi_1 _09324_ (.Y(_03579_),
    .B1(net3066),
    .B2(\core.work.registers.genblk1[13].latch[15] ),
    .A2(net3116),
    .A1(\core.work.registers.genblk1[4].latch[15] ));
 sg13g2_nand4_1 _09325_ (.B(_03577_),
    .C(_03578_),
    .A(_03571_),
    .Y(_03580_),
    .D(_03579_));
 sg13g2_nor2_2 _09326_ (.A(_03576_),
    .B(_03580_),
    .Y(_03581_));
 sg13g2_nor2_2 _09327_ (.A(_03570_),
    .B(_03581_),
    .Y(_03582_));
 sg13g2_o21ai_1 _09328_ (.B1(_03569_),
    .Y(_03583_),
    .A1(net2912),
    .A2(_03582_));
 sg13g2_nand2_1 _09329_ (.Y(_03584_),
    .A(_03568_),
    .B(_03583_));
 sg13g2_nor2_1 _09330_ (.A(_03568_),
    .B(_03583_),
    .Y(_03585_));
 sg13g2_xnor2_1 _09331_ (.Y(_03586_),
    .A(_03568_),
    .B(_03583_));
 sg13g2_o21ai_1 _09332_ (.B1(_03560_),
    .Y(_03587_),
    .A1(_03561_),
    .A2(_03564_));
 sg13g2_xor2_1 _09333_ (.B(_03587_),
    .A(_03586_),
    .X(_03588_));
 sg13g2_o21ai_1 _09334_ (.B1(net2763),
    .Y(_03589_),
    .A1(net2899),
    .A2(_02057_));
 sg13g2_a21oi_2 _09335_ (.B1(_03589_),
    .Y(_03590_),
    .A2(_03588_),
    .A1(net2899));
 sg13g2_a21o_1 _09336_ (.A2(net2783),
    .A1(net617),
    .B1(_03590_),
    .X(_00474_));
 sg13g2_nor2_1 _09337_ (.A(_03561_),
    .B(_03586_),
    .Y(_03591_));
 sg13g2_and2_1 _09338_ (.A(_03563_),
    .B(_03591_),
    .X(_03592_));
 sg13g2_o21ai_1 _09339_ (.B1(_03592_),
    .Y(_03593_),
    .A1(_03491_),
    .A2(_03495_));
 sg13g2_a221oi_1 _09340_ (.B2(_03562_),
    .C1(_03585_),
    .B1(_03591_),
    .A1(_03559_),
    .Y(_03594_),
    .A2(_03584_));
 sg13g2_and2_1 _09341_ (.A(_03593_),
    .B(_03594_),
    .X(_03595_));
 sg13g2_a21oi_1 _09342_ (.A1(_00023_),
    .A2(net2861),
    .Y(_03596_),
    .B1(net2836));
 sg13g2_a21oi_1 _09343_ (.A1(net3479),
    .A2(\core.work.registers.genblk1[1].latch[16] ),
    .Y(_03597_),
    .B1(net3199));
 sg13g2_nand2_1 _09344_ (.Y(_03598_),
    .A(\core.work.registers.genblk1[7].latch[16] ),
    .B(net3124));
 sg13g2_a22oi_1 _09345_ (.Y(_03599_),
    .B1(net3073),
    .B2(\core.work.registers.genblk1[15].latch[16] ),
    .A2(net3093),
    .A1(\core.work.registers.genblk1[12].latch[16] ));
 sg13g2_a22oi_1 _09346_ (.Y(_03600_),
    .B1(net3088),
    .B2(\core.work.registers.genblk1[3].latch[16] ),
    .A2(net3113),
    .A1(\core.work.registers.genblk1[2].latch[16] ));
 sg13g2_a21oi_1 _09347_ (.A1(\core.work.registers.genblk1[5].latch[16] ),
    .A2(net3083),
    .Y(_03601_),
    .B1(net3328));
 sg13g2_a22oi_1 _09348_ (.Y(_03602_),
    .B1(net3103),
    .B2(\core.work.registers.genblk1[14].latch[16] ),
    .A2(net3129),
    .A1(\core.work.registers.genblk1[8].latch[16] ));
 sg13g2_a22oi_1 _09349_ (.Y(_03603_),
    .B1(net3108),
    .B2(\core.work.registers.genblk1[6].latch[16] ),
    .A2(net3133),
    .A1(\core.work.registers.genblk1[10].latch[16] ));
 sg13g2_nand4_1 _09350_ (.B(_03601_),
    .C(_03602_),
    .A(_03600_),
    .Y(_03604_),
    .D(_03603_));
 sg13g2_a22oi_1 _09351_ (.Y(_03605_),
    .B1(net3069),
    .B2(\core.work.registers.genblk1[13].latch[16] ),
    .A2(net3098),
    .A1(\core.work.registers.genblk1[11].latch[16] ));
 sg13g2_a22oi_1 _09352_ (.Y(_03606_),
    .B1(net3078),
    .B2(\core.work.registers.genblk1[9].latch[16] ),
    .A2(net3118),
    .A1(\core.work.registers.genblk1[4].latch[16] ));
 sg13g2_nand4_1 _09353_ (.B(_03599_),
    .C(_03605_),
    .A(_03598_),
    .Y(_03607_),
    .D(_03606_));
 sg13g2_nor2_2 _09354_ (.A(_03604_),
    .B(_03607_),
    .Y(_03608_));
 sg13g2_nor2_2 _09355_ (.A(_03597_),
    .B(_03608_),
    .Y(_03609_));
 sg13g2_nand3_1 _09356_ (.B(_03596_),
    .C(_03609_),
    .A(net2917),
    .Y(_03610_));
 sg13g2_a21o_1 _09357_ (.A2(_03609_),
    .A1(net2917),
    .B1(_03596_),
    .X(_03611_));
 sg13g2_and2_1 _09358_ (.A(_03610_),
    .B(_03611_),
    .X(_03612_));
 sg13g2_nand2b_1 _09359_ (.Y(_03613_),
    .B(_03612_),
    .A_N(_03595_));
 sg13g2_xor2_1 _09360_ (.B(_03612_),
    .A(_03595_),
    .X(_03614_));
 sg13g2_o21ai_1 _09361_ (.B1(net2764),
    .Y(_03615_),
    .A1(net2900),
    .A2(_02255_));
 sg13g2_a21oi_2 _09362_ (.B1(_03615_),
    .Y(_03616_),
    .A2(_03614_),
    .A1(net2900));
 sg13g2_a21o_1 _09363_ (.A2(net2782),
    .A1(net444),
    .B1(_03616_),
    .X(_00475_));
 sg13g2_a21oi_1 _09364_ (.A1(_00025_),
    .A2(_03463_),
    .Y(_03617_),
    .B1(net2836));
 sg13g2_a21oi_1 _09365_ (.A1(net3477),
    .A2(\core.work.registers.genblk1[1].latch[17] ),
    .Y(_03618_),
    .B1(_01657_));
 sg13g2_nand2_1 _09366_ (.Y(_03619_),
    .A(\core.work.registers.genblk1[9].latch[17] ),
    .B(net3078));
 sg13g2_a22oi_1 _09367_ (.Y(_03620_),
    .B1(net3123),
    .B2(\core.work.registers.genblk1[7].latch[17] ),
    .A2(net3128),
    .A1(\core.work.registers.genblk1[8].latch[17] ));
 sg13g2_a22oi_1 _09368_ (.Y(_03621_),
    .B1(net3089),
    .B2(\core.work.registers.genblk1[3].latch[17] ),
    .A2(net3119),
    .A1(\core.work.registers.genblk1[4].latch[17] ));
 sg13g2_a22oi_1 _09369_ (.Y(_03622_),
    .B1(net3068),
    .B2(\core.work.registers.genblk1[13].latch[17] ),
    .A2(net3109),
    .A1(\core.work.registers.genblk1[6].latch[17] ));
 sg13g2_a21oi_1 _09370_ (.A1(\core.work.registers.genblk1[14].latch[17] ),
    .A2(net3104),
    .Y(_03623_),
    .B1(net3325));
 sg13g2_a22oi_1 _09371_ (.Y(_03624_),
    .B1(net3094),
    .B2(\core.work.registers.genblk1[12].latch[17] ),
    .A2(net3133),
    .A1(\core.work.registers.genblk1[10].latch[17] ));
 sg13g2_nand4_1 _09372_ (.B(_03622_),
    .C(_03623_),
    .A(_03621_),
    .Y(_03625_),
    .D(_03624_));
 sg13g2_a22oi_1 _09373_ (.Y(_03626_),
    .B1(net3083),
    .B2(\core.work.registers.genblk1[5].latch[17] ),
    .A2(net3098),
    .A1(\core.work.registers.genblk1[11].latch[17] ));
 sg13g2_a22oi_1 _09374_ (.Y(_03627_),
    .B1(net3073),
    .B2(\core.work.registers.genblk1[15].latch[17] ),
    .A2(net3113),
    .A1(\core.work.registers.genblk1[2].latch[17] ));
 sg13g2_nand4_1 _09375_ (.B(_03620_),
    .C(_03626_),
    .A(_03619_),
    .Y(_03628_),
    .D(_03627_));
 sg13g2_nor2_2 _09376_ (.A(_03625_),
    .B(_03628_),
    .Y(_03629_));
 sg13g2_nor2_2 _09377_ (.A(_03618_),
    .B(_03629_),
    .Y(_03630_));
 sg13g2_nand3_1 _09378_ (.B(_03617_),
    .C(_03630_),
    .A(net2916),
    .Y(_03631_));
 sg13g2_a21o_1 _09379_ (.A2(_03630_),
    .A1(net2916),
    .B1(_03617_),
    .X(_03632_));
 sg13g2_and2_1 _09380_ (.A(_03631_),
    .B(_03632_),
    .X(_03633_));
 sg13g2_nand2_1 _09381_ (.Y(_03634_),
    .A(_03610_),
    .B(_03613_));
 sg13g2_xnor2_1 _09382_ (.Y(_03635_),
    .A(_03633_),
    .B(_03634_));
 sg13g2_o21ai_1 _09383_ (.B1(net2764),
    .Y(_03636_),
    .A1(net2900),
    .A2(_02355_));
 sg13g2_a21oi_2 _09384_ (.B1(_03636_),
    .Y(_03637_),
    .A2(_03635_),
    .A1(net2900));
 sg13g2_a21o_1 _09385_ (.A2(net2781),
    .A1(net489),
    .B1(_03637_),
    .X(_00476_));
 sg13g2_a21oi_1 _09386_ (.A1(_00028_),
    .A2(net2861),
    .Y(_03638_),
    .B1(net2836));
 sg13g2_a21oi_1 _09387_ (.A1(net3479),
    .A2(\core.work.registers.genblk1[1].latch[18] ),
    .Y(_03639_),
    .B1(net3199));
 sg13g2_nand2_1 _09388_ (.Y(_03640_),
    .A(\core.work.registers.genblk1[6].latch[18] ),
    .B(net3108));
 sg13g2_a22oi_1 _09389_ (.Y(_03641_),
    .B1(net3113),
    .B2(\core.work.registers.genblk1[2].latch[18] ),
    .A2(net3118),
    .A1(\core.work.registers.genblk1[4].latch[18] ));
 sg13g2_a21oi_1 _09390_ (.A1(\core.work.registers.genblk1[13].latch[18] ),
    .A2(net3069),
    .Y(_03642_),
    .B1(net3328));
 sg13g2_a22oi_1 _09391_ (.Y(_03643_),
    .B1(net3124),
    .B2(\core.work.registers.genblk1[7].latch[18] ),
    .A2(net3133),
    .A1(\core.work.registers.genblk1[10].latch[18] ));
 sg13g2_a22oi_1 _09392_ (.Y(_03644_),
    .B1(net3078),
    .B2(\core.work.registers.genblk1[9].latch[18] ),
    .A2(net3093),
    .A1(\core.work.registers.genblk1[12].latch[18] ));
 sg13g2_nand4_1 _09393_ (.B(_03642_),
    .C(_03643_),
    .A(_03641_),
    .Y(_03645_),
    .D(_03644_));
 sg13g2_a22oi_1 _09394_ (.Y(_03646_),
    .B1(net3098),
    .B2(\core.work.registers.genblk1[11].latch[18] ),
    .A2(net3103),
    .A1(\core.work.registers.genblk1[14].latch[18] ));
 sg13g2_a22oi_1 _09395_ (.Y(_03647_),
    .B1(net3083),
    .B2(\core.work.registers.genblk1[5].latch[18] ),
    .A2(net3129),
    .A1(\core.work.registers.genblk1[8].latch[18] ));
 sg13g2_a22oi_1 _09396_ (.Y(_03648_),
    .B1(net3073),
    .B2(\core.work.registers.genblk1[15].latch[18] ),
    .A2(net3088),
    .A1(\core.work.registers.genblk1[3].latch[18] ));
 sg13g2_nand4_1 _09397_ (.B(_03646_),
    .C(_03647_),
    .A(_03640_),
    .Y(_03649_),
    .D(_03648_));
 sg13g2_nor2_2 _09398_ (.A(_03645_),
    .B(_03649_),
    .Y(_03650_));
 sg13g2_nor2_2 _09399_ (.A(_03639_),
    .B(_03650_),
    .Y(_03651_));
 sg13g2_and3_1 _09400_ (.X(_03652_),
    .A(net2917),
    .B(_03638_),
    .C(_03651_));
 sg13g2_a21oi_1 _09401_ (.A1(net2916),
    .A2(_03651_),
    .Y(_03653_),
    .B1(_03638_));
 sg13g2_nor2_1 _09402_ (.A(_03652_),
    .B(_03653_),
    .Y(_03654_));
 sg13g2_nand2_1 _09403_ (.Y(_03655_),
    .A(_03610_),
    .B(_03631_));
 sg13g2_inv_1 _09404_ (.Y(_03656_),
    .A(_03655_));
 sg13g2_nand2_1 _09405_ (.Y(_03657_),
    .A(_03612_),
    .B(_03633_));
 sg13g2_o21ai_1 _09406_ (.B1(_03656_),
    .Y(_03658_),
    .A1(_03595_),
    .A2(_03657_));
 sg13g2_xnor2_1 _09407_ (.Y(_03659_),
    .A(_03654_),
    .B(_03658_));
 sg13g2_o21ai_1 _09408_ (.B1(net2764),
    .Y(_03660_),
    .A1(net2901),
    .A2(_02376_));
 sg13g2_a21oi_2 _09409_ (.B1(_03660_),
    .Y(_03661_),
    .A2(_03659_),
    .A1(net2900));
 sg13g2_a21o_1 _09410_ (.A2(net2781),
    .A1(net475),
    .B1(_03661_),
    .X(_00477_));
 sg13g2_a21oi_1 _09411_ (.A1(_00030_),
    .A2(net2861),
    .Y(_03662_),
    .B1(net2836));
 sg13g2_nand2_1 _09412_ (.Y(_03663_),
    .A(net3476),
    .B(\core.work.registers.genblk1[1].latch[19] ));
 sg13g2_nand2_1 _09413_ (.Y(_03664_),
    .A(\core.work.registers.genblk1[13].latch[19] ),
    .B(net3068));
 sg13g2_a22oi_1 _09414_ (.Y(_03665_),
    .B1(net3084),
    .B2(\core.work.registers.genblk1[5].latch[19] ),
    .A2(net3089),
    .A1(\core.work.registers.genblk1[3].latch[19] ));
 sg13g2_a21oi_1 _09415_ (.A1(\core.work.registers.genblk1[11].latch[19] ),
    .A2(net3099),
    .Y(_03666_),
    .B1(net3326));
 sg13g2_a22oi_1 _09416_ (.Y(_03667_),
    .B1(net3094),
    .B2(\core.work.registers.genblk1[12].latch[19] ),
    .A2(net3104),
    .A1(\core.work.registers.genblk1[14].latch[19] ));
 sg13g2_nand3_1 _09417_ (.B(_03666_),
    .C(_03667_),
    .A(_03665_),
    .Y(_03668_));
 sg13g2_a221oi_1 _09418_ (.B2(\core.work.registers.genblk1[6].latch[19] ),
    .C1(_03668_),
    .B1(net3109),
    .A1(\core.work.registers.genblk1[2].latch[19] ),
    .Y(_03669_),
    .A2(net3114));
 sg13g2_a22oi_1 _09419_ (.Y(_03670_),
    .B1(net3119),
    .B2(\core.work.registers.genblk1[4].latch[19] ),
    .A2(net3134),
    .A1(\core.work.registers.genblk1[10].latch[19] ));
 sg13g2_a22oi_1 _09420_ (.Y(_03671_),
    .B1(net3123),
    .B2(\core.work.registers.genblk1[7].latch[19] ),
    .A2(net3129),
    .A1(\core.work.registers.genblk1[8].latch[19] ));
 sg13g2_nand3_1 _09421_ (.B(_03670_),
    .C(_03671_),
    .A(_03664_),
    .Y(_03672_));
 sg13g2_a221oi_1 _09422_ (.B2(\core.work.registers.genblk1[15].latch[19] ),
    .C1(_03672_),
    .B1(net3074),
    .A1(\core.work.registers.genblk1[9].latch[19] ),
    .Y(_03673_),
    .A2(net3079));
 sg13g2_a22oi_1 _09423_ (.Y(_03674_),
    .B1(_03669_),
    .B2(_03673_),
    .A2(_03663_),
    .A1(net3326));
 sg13g2_and3_1 _09424_ (.X(_03675_),
    .A(net2917),
    .B(_03662_),
    .C(_03674_));
 sg13g2_a21oi_1 _09425_ (.A1(net2917),
    .A2(_03674_),
    .Y(_03676_),
    .B1(_03662_));
 sg13g2_nor2_1 _09426_ (.A(_03675_),
    .B(_03676_),
    .Y(_03677_));
 sg13g2_a21oi_1 _09427_ (.A1(_03654_),
    .A2(_03658_),
    .Y(_03678_),
    .B1(_03652_));
 sg13g2_xor2_1 _09428_ (.B(_03678_),
    .A(_03677_),
    .X(_03679_));
 sg13g2_o21ai_1 _09429_ (.B1(net2764),
    .Y(_03680_),
    .A1(net2901),
    .A2(_02396_));
 sg13g2_a21oi_2 _09430_ (.B1(_03680_),
    .Y(_03681_),
    .A2(_03679_),
    .A1(net2901));
 sg13g2_a21o_1 _09431_ (.A2(net2782),
    .A1(net467),
    .B1(_03681_),
    .X(_00478_));
 sg13g2_nor3_1 _09432_ (.A(_03652_),
    .B(_03655_),
    .C(_03675_),
    .Y(_03682_));
 sg13g2_inv_1 _09433_ (.Y(_03683_),
    .A(_03682_));
 sg13g2_nand4_1 _09434_ (.B(_03633_),
    .C(_03654_),
    .A(_03612_),
    .Y(_03684_),
    .D(_03677_));
 sg13g2_a21oi_1 _09435_ (.A1(_03593_),
    .A2(_03594_),
    .Y(_03685_),
    .B1(_03684_));
 sg13g2_nor2_1 _09436_ (.A(_03683_),
    .B(_03685_),
    .Y(_03686_));
 sg13g2_a21oi_1 _09437_ (.A1(net3479),
    .A2(\core.work.registers.genblk1[1].latch[20] ),
    .Y(_03687_),
    .B1(net3199));
 sg13g2_nand2_1 _09438_ (.Y(_03688_),
    .A(\core.work.registers.genblk1[10].latch[20] ),
    .B(net3133));
 sg13g2_a22oi_1 _09439_ (.Y(_03689_),
    .B1(net3083),
    .B2(\core.work.registers.genblk1[5].latch[20] ),
    .A2(net3113),
    .A1(\core.work.registers.genblk1[2].latch[20] ));
 sg13g2_a22oi_1 _09440_ (.Y(_03690_),
    .B1(net3093),
    .B2(\core.work.registers.genblk1[12].latch[20] ),
    .A2(net3118),
    .A1(\core.work.registers.genblk1[4].latch[20] ));
 sg13g2_a21oi_1 _09441_ (.A1(\core.work.registers.genblk1[15].latch[20] ),
    .A2(net3073),
    .Y(_03691_),
    .B1(net3328));
 sg13g2_a22oi_1 _09442_ (.Y(_03692_),
    .B1(net3098),
    .B2(\core.work.registers.genblk1[11].latch[20] ),
    .A2(net3103),
    .A1(\core.work.registers.genblk1[14].latch[20] ));
 sg13g2_a22oi_1 _09443_ (.Y(_03693_),
    .B1(net3069),
    .B2(\core.work.registers.genblk1[13].latch[20] ),
    .A2(net3078),
    .A1(\core.work.registers.genblk1[9].latch[20] ));
 sg13g2_nand4_1 _09444_ (.B(_03691_),
    .C(_03692_),
    .A(_03690_),
    .Y(_03694_),
    .D(_03693_));
 sg13g2_a22oi_1 _09445_ (.Y(_03695_),
    .B1(net3108),
    .B2(\core.work.registers.genblk1[6].latch[20] ),
    .A2(net3124),
    .A1(\core.work.registers.genblk1[7].latch[20] ));
 sg13g2_a22oi_1 _09446_ (.Y(_03696_),
    .B1(net3088),
    .B2(\core.work.registers.genblk1[3].latch[20] ),
    .A2(net3129),
    .A1(\core.work.registers.genblk1[8].latch[20] ));
 sg13g2_nand4_1 _09447_ (.B(_03689_),
    .C(_03695_),
    .A(_03688_),
    .Y(_03697_),
    .D(_03696_));
 sg13g2_nor2_1 _09448_ (.A(_03694_),
    .B(_03697_),
    .Y(_03698_));
 sg13g2_nor2_2 _09449_ (.A(_03687_),
    .B(_03698_),
    .Y(_03699_));
 sg13g2_nand2_1 _09450_ (.Y(_03700_),
    .A(net2916),
    .B(_03699_));
 sg13g2_xnor2_1 _09451_ (.Y(_03701_),
    .A(net3442),
    .B(_03700_));
 sg13g2_inv_1 _09452_ (.Y(_03702_),
    .A(_03701_));
 sg13g2_o21ai_1 _09453_ (.B1(_03702_),
    .Y(_03703_),
    .A1(_03683_),
    .A2(_03685_));
 sg13g2_xnor2_1 _09454_ (.Y(_03704_),
    .A(_03686_),
    .B(_03701_));
 sg13g2_o21ai_1 _09455_ (.B1(net2764),
    .Y(_03705_),
    .A1(net2900),
    .A2(_02414_));
 sg13g2_a21oi_2 _09456_ (.B1(_03705_),
    .Y(_03706_),
    .A2(_03704_),
    .A1(net2900));
 sg13g2_a21o_1 _09457_ (.A2(net2782),
    .A1(net488),
    .B1(_03706_),
    .X(_00479_));
 sg13g2_a21oi_1 _09458_ (.A1(net3474),
    .A2(\core.work.registers.genblk1[1].latch[21] ),
    .Y(_03707_),
    .B1(net3198));
 sg13g2_nand2_1 _09459_ (.Y(_03708_),
    .A(\core.work.registers.genblk1[8].latch[21] ),
    .B(net3127));
 sg13g2_a21oi_1 _09460_ (.A1(\core.work.registers.genblk1[13].latch[21] ),
    .A2(net3067),
    .Y(_03709_),
    .B1(net3322));
 sg13g2_a22oi_1 _09461_ (.Y(_03710_),
    .B1(net3077),
    .B2(\core.work.registers.genblk1[9].latch[21] ),
    .A2(net3122),
    .A1(\core.work.registers.genblk1[7].latch[21] ));
 sg13g2_a22oi_1 _09462_ (.Y(_03711_),
    .B1(net3097),
    .B2(\core.work.registers.genblk1[11].latch[21] ),
    .A2(net3117),
    .A1(\core.work.registers.genblk1[4].latch[21] ));
 sg13g2_a22oi_1 _09463_ (.Y(_03712_),
    .B1(net3112),
    .B2(\core.work.registers.genblk1[2].latch[21] ),
    .A2(net3132),
    .A1(\core.work.registers.genblk1[10].latch[21] ));
 sg13g2_nand4_1 _09464_ (.B(_03710_),
    .C(_03711_),
    .A(_03709_),
    .Y(_03713_),
    .D(_03712_));
 sg13g2_a22oi_1 _09465_ (.Y(_03714_),
    .B1(net3087),
    .B2(\core.work.registers.genblk1[3].latch[21] ),
    .A2(net3107),
    .A1(\core.work.registers.genblk1[6].latch[21] ));
 sg13g2_a22oi_1 _09466_ (.Y(_03715_),
    .B1(net3072),
    .B2(\core.work.registers.genblk1[15].latch[21] ),
    .A2(net3092),
    .A1(\core.work.registers.genblk1[12].latch[21] ));
 sg13g2_a22oi_1 _09467_ (.Y(_03716_),
    .B1(net3082),
    .B2(\core.work.registers.genblk1[5].latch[21] ),
    .A2(net3102),
    .A1(\core.work.registers.genblk1[14].latch[21] ));
 sg13g2_nand4_1 _09468_ (.B(_03714_),
    .C(_03715_),
    .A(_03708_),
    .Y(_03717_),
    .D(_03716_));
 sg13g2_nor2_2 _09469_ (.A(_03713_),
    .B(_03717_),
    .Y(_03718_));
 sg13g2_nor2_2 _09470_ (.A(_03707_),
    .B(_03718_),
    .Y(_03719_));
 sg13g2_nand2_1 _09471_ (.Y(_03720_),
    .A(net2915),
    .B(_03719_));
 sg13g2_nand2_1 _09472_ (.Y(_03721_),
    .A(net3442),
    .B(_03720_));
 sg13g2_nor2_1 _09473_ (.A(_00605_),
    .B(_03700_),
    .Y(_03722_));
 sg13g2_inv_1 _09474_ (.Y(_03723_),
    .A(_03722_));
 sg13g2_nand2_1 _09475_ (.Y(_03724_),
    .A(_03703_),
    .B(_03723_));
 sg13g2_nor2_1 _09476_ (.A(net3442),
    .B(_03720_),
    .Y(_03725_));
 sg13g2_inv_1 _09477_ (.Y(_03726_),
    .A(_03725_));
 sg13g2_nand3_1 _09478_ (.B(_03723_),
    .C(_03726_),
    .A(_03703_),
    .Y(_03727_));
 sg13g2_and2_1 _09479_ (.A(_03721_),
    .B(_03726_),
    .X(_03728_));
 sg13g2_xnor2_1 _09480_ (.Y(_03729_),
    .A(_03724_),
    .B(_03728_));
 sg13g2_o21ai_1 _09481_ (.B1(net2762),
    .Y(_03730_),
    .A1(net2899),
    .A2(_02278_));
 sg13g2_a21oi_2 _09482_ (.B1(_03730_),
    .Y(_03731_),
    .A2(_03729_),
    .A1(net2899));
 sg13g2_a21o_1 _09483_ (.A2(net2783),
    .A1(net491),
    .B1(_03731_),
    .X(_00480_));
 sg13g2_nand2_1 _09484_ (.Y(_03732_),
    .A(_03721_),
    .B(_03727_));
 sg13g2_a21oi_1 _09485_ (.A1(net3473),
    .A2(\core.work.registers.genblk1[1].latch[22] ),
    .Y(_03733_),
    .B1(net3198));
 sg13g2_nand2_1 _09486_ (.Y(_03734_),
    .A(\core.work.registers.genblk1[10].latch[22] ),
    .B(net3132));
 sg13g2_a22oi_1 _09487_ (.Y(_03735_),
    .B1(net3072),
    .B2(\core.work.registers.genblk1[15].latch[22] ),
    .A2(net3112),
    .A1(\core.work.registers.genblk1[2].latch[22] ));
 sg13g2_a22oi_1 _09488_ (.Y(_03736_),
    .B1(net3087),
    .B2(\core.work.registers.genblk1[3].latch[22] ),
    .A2(net3102),
    .A1(\core.work.registers.genblk1[14].latch[22] ));
 sg13g2_a22oi_1 _09489_ (.Y(_03737_),
    .B1(net3092),
    .B2(\core.work.registers.genblk1[12].latch[22] ),
    .A2(net3107),
    .A1(\core.work.registers.genblk1[6].latch[22] ));
 sg13g2_a21oi_1 _09490_ (.A1(\core.work.registers.genblk1[8].latch[22] ),
    .A2(net3127),
    .Y(_03738_),
    .B1(net3321));
 sg13g2_a22oi_1 _09491_ (.Y(_03739_),
    .B1(net3077),
    .B2(\core.work.registers.genblk1[9].latch[22] ),
    .A2(net3082),
    .A1(\core.work.registers.genblk1[5].latch[22] ));
 sg13g2_a22oi_1 _09492_ (.Y(_03740_),
    .B1(net3097),
    .B2(\core.work.registers.genblk1[11].latch[22] ),
    .A2(net3122),
    .A1(\core.work.registers.genblk1[7].latch[22] ));
 sg13g2_nand4_1 _09493_ (.B(_03738_),
    .C(_03739_),
    .A(_03737_),
    .Y(_03741_),
    .D(_03740_));
 sg13g2_a22oi_1 _09494_ (.Y(_03742_),
    .B1(net3067),
    .B2(\core.work.registers.genblk1[13].latch[22] ),
    .A2(net3117),
    .A1(\core.work.registers.genblk1[4].latch[22] ));
 sg13g2_nand4_1 _09495_ (.B(_03735_),
    .C(_03736_),
    .A(_03734_),
    .Y(_03743_),
    .D(_03742_));
 sg13g2_nor2_1 _09496_ (.A(_03741_),
    .B(_03743_),
    .Y(_03744_));
 sg13g2_nor2_2 _09497_ (.A(_03733_),
    .B(_03744_),
    .Y(_03745_));
 sg13g2_nand2_1 _09498_ (.Y(_03746_),
    .A(net2913),
    .B(_03745_));
 sg13g2_xnor2_1 _09499_ (.Y(_03747_),
    .A(net3359),
    .B(_03746_));
 sg13g2_nand3_1 _09500_ (.B(_03727_),
    .C(_03747_),
    .A(_03721_),
    .Y(_03748_));
 sg13g2_xor2_1 _09501_ (.B(_03747_),
    .A(_03732_),
    .X(_03749_));
 sg13g2_o21ai_1 _09502_ (.B1(net2762),
    .Y(_03750_),
    .A1(net2897),
    .A2(_02298_));
 sg13g2_a21oi_2 _09503_ (.B1(_03750_),
    .Y(_03751_),
    .A2(_03749_),
    .A1(net2898));
 sg13g2_a21o_1 _09504_ (.A2(net2784),
    .A1(net483),
    .B1(_03751_),
    .X(_00481_));
 sg13g2_nand2_1 _09505_ (.Y(_03752_),
    .A(net584),
    .B(net2784));
 sg13g2_a21oi_1 _09506_ (.A1(net3473),
    .A2(\core.work.registers.genblk1[1].latch[23] ),
    .Y(_03753_),
    .B1(net3197));
 sg13g2_a22oi_1 _09507_ (.Y(_03754_),
    .B1(net3106),
    .B2(\core.work.registers.genblk1[6].latch[23] ),
    .A2(net3126),
    .A1(\core.work.registers.genblk1[8].latch[23] ));
 sg13g2_nand2_1 _09508_ (.Y(_03755_),
    .A(\core.work.registers.genblk1[10].latch[23] ),
    .B(net3131));
 sg13g2_a22oi_1 _09509_ (.Y(_03756_),
    .B1(net3101),
    .B2(\core.work.registers.genblk1[14].latch[23] ),
    .A2(net3121),
    .A1(\core.work.registers.genblk1[7].latch[23] ));
 sg13g2_a22oi_1 _09510_ (.Y(_03757_),
    .B1(net3111),
    .B2(\core.work.registers.genblk1[2].latch[23] ),
    .A2(net3116),
    .A1(\core.work.registers.genblk1[4].latch[23] ));
 sg13g2_a21oi_1 _09511_ (.A1(\core.work.registers.genblk1[3].latch[23] ),
    .A2(net3086),
    .Y(_03758_),
    .B1(net3321));
 sg13g2_a22oi_1 _09512_ (.Y(_03759_),
    .B1(net3066),
    .B2(\core.work.registers.genblk1[13].latch[23] ),
    .A2(net3076),
    .A1(\core.work.registers.genblk1[9].latch[23] ));
 sg13g2_a22oi_1 _09513_ (.Y(_03760_),
    .B1(net3071),
    .B2(\core.work.registers.genblk1[15].latch[23] ),
    .A2(net3096),
    .A1(\core.work.registers.genblk1[11].latch[23] ));
 sg13g2_nand4_1 _09514_ (.B(_03758_),
    .C(_03759_),
    .A(_03757_),
    .Y(_03761_),
    .D(_03760_));
 sg13g2_a22oi_1 _09515_ (.Y(_03762_),
    .B1(net3081),
    .B2(\core.work.registers.genblk1[5].latch[23] ),
    .A2(net3091),
    .A1(\core.work.registers.genblk1[12].latch[23] ));
 sg13g2_nand4_1 _09516_ (.B(_03755_),
    .C(_03756_),
    .A(_03754_),
    .Y(_03763_),
    .D(_03762_));
 sg13g2_nor2_2 _09517_ (.A(_03761_),
    .B(_03763_),
    .Y(_03764_));
 sg13g2_nor2_2 _09518_ (.A(_03753_),
    .B(_03764_),
    .Y(_03765_));
 sg13g2_nand2_1 _09519_ (.Y(_03766_),
    .A(net2914),
    .B(_03765_));
 sg13g2_nand3_1 _09520_ (.B(net2913),
    .C(_03765_),
    .A(net3359),
    .Y(_03767_));
 sg13g2_xnor2_1 _09521_ (.Y(_03768_),
    .A(net3360),
    .B(_03766_));
 sg13g2_nor2_1 _09522_ (.A(_00605_),
    .B(_03746_),
    .Y(_03769_));
 sg13g2_inv_1 _09523_ (.Y(_03770_),
    .A(_03769_));
 sg13g2_and3_1 _09524_ (.X(_03771_),
    .A(_03748_),
    .B(_03768_),
    .C(_03770_));
 sg13g2_a21oi_1 _09525_ (.A1(_03748_),
    .A2(_03770_),
    .Y(_03772_),
    .B1(_03768_));
 sg13g2_nor3_1 _09526_ (.A(net2908),
    .B(_03771_),
    .C(_03772_),
    .Y(_03773_));
 sg13g2_o21ai_1 _09527_ (.B1(net2762),
    .Y(_03774_),
    .A1(net2898),
    .A2(_02317_));
 sg13g2_o21ai_1 _09528_ (.B1(_03752_),
    .Y(_00482_),
    .A1(_03773_),
    .A2(_03774_));
 sg13g2_nand3_1 _09529_ (.B(_03747_),
    .C(_03768_),
    .A(_03721_),
    .Y(_03775_));
 sg13g2_nor4_1 _09530_ (.A(_03684_),
    .B(_03701_),
    .C(_03725_),
    .D(_03775_),
    .Y(_03776_));
 sg13g2_inv_1 _09531_ (.Y(_03777_),
    .A(_03776_));
 sg13g2_a21oi_2 _09532_ (.B1(_03777_),
    .Y(_03778_),
    .A2(_03594_),
    .A1(_03593_));
 sg13g2_nor2_1 _09533_ (.A(_03722_),
    .B(_03725_),
    .Y(_03779_));
 sg13g2_o21ai_1 _09534_ (.B1(_03779_),
    .Y(_03780_),
    .A1(_03682_),
    .A2(_03701_));
 sg13g2_nand2b_1 _09535_ (.Y(_03781_),
    .B(_03780_),
    .A_N(_03775_));
 sg13g2_a21o_1 _09536_ (.A2(_03766_),
    .A1(net3442),
    .B1(_03770_),
    .X(_03782_));
 sg13g2_nand3_1 _09537_ (.B(_03781_),
    .C(_03782_),
    .A(_03767_),
    .Y(_03783_));
 sg13g2_a21oi_1 _09538_ (.A1(net3479),
    .A2(\core.work.registers.genblk1[1].latch[24] ),
    .Y(_03784_),
    .B1(net3199));
 sg13g2_nand2_1 _09539_ (.Y(_03785_),
    .A(\core.work.registers.genblk1[5].latch[24] ),
    .B(net3083));
 sg13g2_a22oi_1 _09540_ (.Y(_03786_),
    .B1(net3073),
    .B2(\core.work.registers.genblk1[15].latch[24] ),
    .A2(net3093),
    .A1(\core.work.registers.genblk1[12].latch[24] ));
 sg13g2_a22oi_1 _09541_ (.Y(_03787_),
    .B1(net3108),
    .B2(\core.work.registers.genblk1[6].latch[24] ),
    .A2(net3113),
    .A1(\core.work.registers.genblk1[2].latch[24] ));
 sg13g2_a22oi_1 _09542_ (.Y(_03788_),
    .B1(net3078),
    .B2(\core.work.registers.genblk1[9].latch[24] ),
    .A2(net3129),
    .A1(\core.work.registers.genblk1[8].latch[24] ));
 sg13g2_a21oi_1 _09543_ (.A1(\core.work.registers.genblk1[7].latch[24] ),
    .A2(net3124),
    .Y(_03789_),
    .B1(net3328));
 sg13g2_a22oi_1 _09544_ (.Y(_03790_),
    .B1(net3103),
    .B2(\core.work.registers.genblk1[14].latch[24] ),
    .A2(net3118),
    .A1(\core.work.registers.genblk1[4].latch[24] ));
 sg13g2_nand4_1 _09545_ (.B(_03788_),
    .C(_03789_),
    .A(_03787_),
    .Y(_03791_),
    .D(_03790_));
 sg13g2_a22oi_1 _09546_ (.Y(_03792_),
    .B1(net3069),
    .B2(\core.work.registers.genblk1[13].latch[24] ),
    .A2(net3098),
    .A1(\core.work.registers.genblk1[11].latch[24] ));
 sg13g2_a22oi_1 _09547_ (.Y(_03793_),
    .B1(net3088),
    .B2(\core.work.registers.genblk1[3].latch[24] ),
    .A2(net3133),
    .A1(\core.work.registers.genblk1[10].latch[24] ));
 sg13g2_nand4_1 _09548_ (.B(_03786_),
    .C(_03792_),
    .A(_03785_),
    .Y(_03794_),
    .D(_03793_));
 sg13g2_nor2_1 _09549_ (.A(_03791_),
    .B(_03794_),
    .Y(_03795_));
 sg13g2_nor2_2 _09550_ (.A(_03784_),
    .B(_03795_),
    .Y(_03796_));
 sg13g2_nand2_2 _09551_ (.Y(_03797_),
    .A(net2915),
    .B(_03796_));
 sg13g2_inv_1 _09552_ (.Y(_03798_),
    .A(_03797_));
 sg13g2_xnor2_1 _09553_ (.Y(_03799_),
    .A(net3360),
    .B(_03797_));
 sg13g2_o21ai_1 _09554_ (.B1(_03799_),
    .Y(_03800_),
    .A1(_03778_),
    .A2(_03783_));
 sg13g2_inv_1 _09555_ (.Y(_03801_),
    .A(_03800_));
 sg13g2_nor3_1 _09556_ (.A(_03778_),
    .B(_03783_),
    .C(_03799_),
    .Y(_03802_));
 sg13g2_o21ai_1 _09557_ (.B1(net2897),
    .Y(_03803_),
    .A1(_03801_),
    .A2(_03802_));
 sg13g2_o21ai_1 _09558_ (.B1(_03803_),
    .Y(_03804_),
    .A1(net2900),
    .A2(_02336_));
 sg13g2_nand2_1 _09559_ (.Y(_03805_),
    .A(net413),
    .B(net2781));
 sg13g2_o21ai_1 _09560_ (.B1(_03805_),
    .Y(_00483_),
    .A1(_03197_),
    .A2(_03804_));
 sg13g2_o21ai_1 _09561_ (.B1(_03800_),
    .Y(_03806_),
    .A1(_00605_),
    .A2(_03797_));
 sg13g2_nand2_1 _09562_ (.Y(_03807_),
    .A(net3474),
    .B(\core.work.registers.genblk1[1].latch[25] ));
 sg13g2_nand2_1 _09563_ (.Y(_03808_),
    .A(\core.work.registers.genblk1[2].latch[25] ),
    .B(net3112));
 sg13g2_a22oi_1 _09564_ (.Y(_03809_),
    .B1(net3082),
    .B2(\core.work.registers.genblk1[5].latch[25] ),
    .A2(net3092),
    .A1(\core.work.registers.genblk1[12].latch[25] ));
 sg13g2_a22oi_1 _09565_ (.Y(_03810_),
    .B1(net3067),
    .B2(\core.work.registers.genblk1[13].latch[25] ),
    .A2(net3087),
    .A1(\core.work.registers.genblk1[3].latch[25] ));
 sg13g2_a21oi_1 _09566_ (.A1(\core.work.registers.genblk1[14].latch[25] ),
    .A2(net3102),
    .Y(_03811_),
    .B1(net3322));
 sg13g2_a22oi_1 _09567_ (.Y(_03812_),
    .B1(net3122),
    .B2(\core.work.registers.genblk1[7].latch[25] ),
    .A2(net3127),
    .A1(\core.work.registers.genblk1[8].latch[25] ));
 sg13g2_a22oi_1 _09568_ (.Y(_03813_),
    .B1(net3077),
    .B2(\core.work.registers.genblk1[9].latch[25] ),
    .A2(net3107),
    .A1(\core.work.registers.genblk1[6].latch[25] ));
 sg13g2_nand3_1 _09569_ (.B(_03812_),
    .C(_03813_),
    .A(_03811_),
    .Y(_03814_));
 sg13g2_a221oi_1 _09570_ (.B2(\core.work.registers.genblk1[15].latch[25] ),
    .C1(_03814_),
    .B1(net3072),
    .A1(\core.work.registers.genblk1[11].latch[25] ),
    .Y(_03815_),
    .A2(net3097));
 sg13g2_nand3_1 _09571_ (.B(_03809_),
    .C(_03810_),
    .A(_03808_),
    .Y(_03816_));
 sg13g2_a221oi_1 _09572_ (.B2(\core.work.registers.genblk1[4].latch[25] ),
    .C1(_03816_),
    .B1(net3117),
    .A1(\core.work.registers.genblk1[10].latch[25] ),
    .Y(_03817_),
    .A2(net3132));
 sg13g2_a22oi_1 _09573_ (.Y(_03818_),
    .B1(_03815_),
    .B2(_03817_),
    .A2(_03807_),
    .A1(net3322));
 sg13g2_a21oi_1 _09574_ (.A1(net2914),
    .A2(_03818_),
    .Y(_03819_),
    .B1(net3359));
 sg13g2_and3_1 _09575_ (.X(_03820_),
    .A(net3360),
    .B(net2913),
    .C(_03818_));
 sg13g2_nor2_1 _09576_ (.A(_03819_),
    .B(_03820_),
    .Y(_03821_));
 sg13g2_xnor2_1 _09577_ (.Y(_03822_),
    .A(_03806_),
    .B(_03821_));
 sg13g2_o21ai_1 _09578_ (.B1(net2762),
    .Y(_03823_),
    .A1(net2898),
    .A2(_02235_));
 sg13g2_a21oi_2 _09579_ (.B1(_03823_),
    .Y(_03824_),
    .A2(_03822_),
    .A1(net2898));
 sg13g2_a21o_1 _09580_ (.A2(net2783),
    .A1(net476),
    .B1(_03824_),
    .X(_00484_));
 sg13g2_a21oi_1 _09581_ (.A1(net3473),
    .A2(\core.work.registers.genblk1[1].latch[26] ),
    .Y(_03825_),
    .B1(net3197));
 sg13g2_a22oi_1 _09582_ (.Y(_03826_),
    .B1(net3096),
    .B2(\core.work.registers.genblk1[11].latch[26] ),
    .A2(net3126),
    .A1(\core.work.registers.genblk1[8].latch[26] ));
 sg13g2_a22oi_1 _09583_ (.Y(_03827_),
    .B1(net3091),
    .B2(\core.work.registers.genblk1[12].latch[26] ),
    .A2(net3131),
    .A1(\core.work.registers.genblk1[10].latch[26] ));
 sg13g2_a21oi_1 _09584_ (.A1(\core.work.registers.genblk1[14].latch[26] ),
    .A2(net3101),
    .Y(_03828_),
    .B1(net3321));
 sg13g2_a22oi_1 _09585_ (.Y(_03829_),
    .B1(net3081),
    .B2(\core.work.registers.genblk1[5].latch[26] ),
    .A2(net3116),
    .A1(\core.work.registers.genblk1[4].latch[26] ));
 sg13g2_nand4_1 _09586_ (.B(_03827_),
    .C(_03828_),
    .A(_03826_),
    .Y(_03830_),
    .D(_03829_));
 sg13g2_nand2_1 _09587_ (.Y(_03831_),
    .A(\core.work.registers.genblk1[7].latch[26] ),
    .B(net3121));
 sg13g2_a22oi_1 _09588_ (.Y(_03832_),
    .B1(net3076),
    .B2(\core.work.registers.genblk1[9].latch[26] ),
    .A2(net3086),
    .A1(\core.work.registers.genblk1[3].latch[26] ));
 sg13g2_a22oi_1 _09589_ (.Y(_03833_),
    .B1(net3066),
    .B2(\core.work.registers.genblk1[13].latch[26] ),
    .A2(net3111),
    .A1(\core.work.registers.genblk1[2].latch[26] ));
 sg13g2_a22oi_1 _09590_ (.Y(_03834_),
    .B1(net3071),
    .B2(\core.work.registers.genblk1[15].latch[26] ),
    .A2(net3106),
    .A1(\core.work.registers.genblk1[6].latch[26] ));
 sg13g2_nand4_1 _09591_ (.B(_03832_),
    .C(_03833_),
    .A(_03831_),
    .Y(_03835_),
    .D(_03834_));
 sg13g2_nor2_2 _09592_ (.A(_03830_),
    .B(_03835_),
    .Y(_03836_));
 sg13g2_nor2_1 _09593_ (.A(_03825_),
    .B(_03836_),
    .Y(_03837_));
 sg13g2_nand2_1 _09594_ (.Y(_03838_),
    .A(net2913),
    .B(_03837_));
 sg13g2_inv_1 _09595_ (.Y(_03839_),
    .A(_03838_));
 sg13g2_xnor2_1 _09596_ (.Y(_03840_),
    .A(net3359),
    .B(_03838_));
 sg13g2_a21oi_1 _09597_ (.A1(net3443),
    .A2(_03798_),
    .Y(_03841_),
    .B1(_03820_));
 sg13g2_a21oi_1 _09598_ (.A1(_03800_),
    .A2(_03841_),
    .Y(_03842_),
    .B1(_03819_));
 sg13g2_xnor2_1 _09599_ (.Y(_03843_),
    .A(_03840_),
    .B(_03842_));
 sg13g2_o21ai_1 _09600_ (.B1(net2762),
    .Y(_03844_),
    .A1(net2897),
    .A2(_02214_));
 sg13g2_a21oi_2 _09601_ (.B1(_03844_),
    .Y(_03845_),
    .A2(_03843_),
    .A1(net2897));
 sg13g2_a21o_1 _09602_ (.A2(net2783),
    .A1(net493),
    .B1(_03845_),
    .X(_00485_));
 sg13g2_a22oi_1 _09603_ (.Y(_03846_),
    .B1(_03840_),
    .B2(_03842_),
    .A2(_03839_),
    .A1(net3443));
 sg13g2_a21oi_1 _09604_ (.A1(net3473),
    .A2(\core.work.registers.genblk1[1].latch[27] ),
    .Y(_03847_),
    .B1(net3197));
 sg13g2_nand2_1 _09605_ (.Y(_03848_),
    .A(\core.work.registers.genblk1[12].latch[27] ),
    .B(net3091));
 sg13g2_a22oi_1 _09606_ (.Y(_03849_),
    .B1(net3081),
    .B2(\core.work.registers.genblk1[5].latch[27] ),
    .A2(net3106),
    .A1(\core.work.registers.genblk1[6].latch[27] ));
 sg13g2_a21oi_1 _09607_ (.A1(\core.work.registers.genblk1[4].latch[27] ),
    .A2(net3117),
    .Y(_03850_),
    .B1(net3321));
 sg13g2_a22oi_1 _09608_ (.Y(_03851_),
    .B1(net3066),
    .B2(\core.work.registers.genblk1[13].latch[27] ),
    .A2(net3111),
    .A1(\core.work.registers.genblk1[2].latch[27] ));
 sg13g2_a22oi_1 _09609_ (.Y(_03852_),
    .B1(net3101),
    .B2(\core.work.registers.genblk1[14].latch[27] ),
    .A2(net3131),
    .A1(\core.work.registers.genblk1[10].latch[27] ));
 sg13g2_a22oi_1 _09610_ (.Y(_03853_),
    .B1(net3071),
    .B2(\core.work.registers.genblk1[15].latch[27] ),
    .A2(net3077),
    .A1(\core.work.registers.genblk1[9].latch[27] ));
 sg13g2_nand4_1 _09611_ (.B(_03851_),
    .C(_03852_),
    .A(_03850_),
    .Y(_03854_),
    .D(_03853_));
 sg13g2_a22oi_1 _09612_ (.Y(_03855_),
    .B1(net3086),
    .B2(\core.work.registers.genblk1[3].latch[27] ),
    .A2(net3096),
    .A1(\core.work.registers.genblk1[11].latch[27] ));
 sg13g2_a22oi_1 _09613_ (.Y(_03856_),
    .B1(net3121),
    .B2(\core.work.registers.genblk1[7].latch[27] ),
    .A2(net3126),
    .A1(\core.work.registers.genblk1[8].latch[27] ));
 sg13g2_nand4_1 _09614_ (.B(_03849_),
    .C(_03855_),
    .A(_03848_),
    .Y(_03857_),
    .D(_03856_));
 sg13g2_nor2_2 _09615_ (.A(_03854_),
    .B(_03857_),
    .Y(_03858_));
 sg13g2_nor2_2 _09616_ (.A(_03847_),
    .B(_03858_),
    .Y(_03859_));
 sg13g2_nand2_1 _09617_ (.Y(_03860_),
    .A(net2913),
    .B(_03859_));
 sg13g2_xnor2_1 _09618_ (.Y(_03861_),
    .A(net3359),
    .B(_03860_));
 sg13g2_xor2_1 _09619_ (.B(_03861_),
    .A(_03846_),
    .X(_03862_));
 sg13g2_o21ai_1 _09620_ (.B1(net2762),
    .Y(_03863_),
    .A1(net2897),
    .A2(_02191_));
 sg13g2_a21oi_2 _09621_ (.B1(_03863_),
    .Y(_03864_),
    .A2(_03862_),
    .A1(net2897));
 sg13g2_a21o_1 _09622_ (.A2(net2783),
    .A1(net529),
    .B1(_03864_),
    .X(_00486_));
 sg13g2_nand2_1 _09623_ (.Y(_03865_),
    .A(_03840_),
    .B(_03861_));
 sg13g2_and4_1 _09624_ (.A(_03799_),
    .B(_03821_),
    .C(_03840_),
    .D(_03861_),
    .X(_03866_));
 sg13g2_o21ai_1 _09625_ (.B1(_03866_),
    .Y(_03867_),
    .A1(_03778_),
    .A2(_03783_));
 sg13g2_nor3_1 _09626_ (.A(_03819_),
    .B(_03841_),
    .C(_03865_),
    .Y(_03868_));
 sg13g2_o21ai_1 _09627_ (.B1(_03860_),
    .Y(_03869_),
    .A1(net3442),
    .A2(_03838_));
 sg13g2_a21oi_1 _09628_ (.A1(net3443),
    .A2(_03869_),
    .Y(_03870_),
    .B1(_03868_));
 sg13g2_nand2_1 _09629_ (.Y(_03871_),
    .A(_03867_),
    .B(_03870_));
 sg13g2_a21oi_1 _09630_ (.A1(net3475),
    .A2(\core.work.registers.genblk1[1].latch[28] ),
    .Y(_03872_),
    .B1(net3197));
 sg13g2_nand2_1 _09631_ (.Y(_03873_),
    .A(\core.work.registers.genblk1[4].latch[28] ),
    .B(net3116));
 sg13g2_a22oi_1 _09632_ (.Y(_03874_),
    .B1(net3086),
    .B2(\core.work.registers.genblk1[3].latch[28] ),
    .A2(net3111),
    .A1(\core.work.registers.genblk1[2].latch[28] ));
 sg13g2_a21oi_1 _09633_ (.A1(\core.work.registers.genblk1[6].latch[28] ),
    .A2(net3106),
    .Y(_03875_),
    .B1(net3321));
 sg13g2_a22oi_1 _09634_ (.Y(_03876_),
    .B1(net3071),
    .B2(\core.work.registers.genblk1[15].latch[28] ),
    .A2(net3091),
    .A1(\core.work.registers.genblk1[12].latch[28] ));
 sg13g2_a22oi_1 _09635_ (.Y(_03877_),
    .B1(net3076),
    .B2(\core.work.registers.genblk1[9].latch[28] ),
    .A2(net3081),
    .A1(\core.work.registers.genblk1[5].latch[28] ));
 sg13g2_a22oi_1 _09636_ (.Y(_03878_),
    .B1(net3121),
    .B2(\core.work.registers.genblk1[7].latch[28] ),
    .A2(net3126),
    .A1(\core.work.registers.genblk1[8].latch[28] ));
 sg13g2_nand4_1 _09637_ (.B(_03876_),
    .C(_03877_),
    .A(_03875_),
    .Y(_03879_),
    .D(_03878_));
 sg13g2_a22oi_1 _09638_ (.Y(_03880_),
    .B1(net3066),
    .B2(\core.work.registers.genblk1[13].latch[28] ),
    .A2(net3131),
    .A1(\core.work.registers.genblk1[10].latch[28] ));
 sg13g2_a22oi_1 _09639_ (.Y(_03881_),
    .B1(net3096),
    .B2(\core.work.registers.genblk1[11].latch[28] ),
    .A2(net3101),
    .A1(\core.work.registers.genblk1[14].latch[28] ));
 sg13g2_nand4_1 _09640_ (.B(_03874_),
    .C(_03880_),
    .A(_03873_),
    .Y(_03882_),
    .D(_03881_));
 sg13g2_nor2_2 _09641_ (.A(_03879_),
    .B(_03882_),
    .Y(_03883_));
 sg13g2_nor2_2 _09642_ (.A(_03872_),
    .B(_03883_),
    .Y(_03884_));
 sg13g2_nand2_1 _09643_ (.Y(_03885_),
    .A(net2913),
    .B(_03884_));
 sg13g2_inv_1 _09644_ (.Y(_03886_),
    .A(_03885_));
 sg13g2_nand2_1 _09645_ (.Y(_03887_),
    .A(net3359),
    .B(_03886_));
 sg13g2_xnor2_1 _09646_ (.Y(_03888_),
    .A(net3359),
    .B(_03885_));
 sg13g2_xnor2_1 _09647_ (.Y(_03889_),
    .A(_03871_),
    .B(_03888_));
 sg13g2_o21ai_1 _09648_ (.B1(net2762),
    .Y(_03890_),
    .A1(net2897),
    .A2(_02172_));
 sg13g2_a21oi_1 _09649_ (.A1(net2897),
    .A2(_03889_),
    .Y(_03891_),
    .B1(_03890_));
 sg13g2_a21o_1 _09650_ (.A2(net2784),
    .A1(net662),
    .B1(_03891_),
    .X(_00487_));
 sg13g2_a22oi_1 _09651_ (.Y(_03892_),
    .B1(_03888_),
    .B2(_03871_),
    .A2(_03886_),
    .A1(net3443));
 sg13g2_a21oi_1 _09652_ (.A1(net3475),
    .A2(\core.work.registers.genblk1[1].latch[29] ),
    .Y(_03893_),
    .B1(net3197));
 sg13g2_nand2_1 _09653_ (.Y(_03894_),
    .A(\core.work.registers.genblk1[13].latch[29] ),
    .B(net3066));
 sg13g2_a21oi_1 _09654_ (.A1(\core.work.registers.genblk1[6].latch[29] ),
    .A2(net3106),
    .Y(_03895_),
    .B1(net3321));
 sg13g2_a22oi_1 _09655_ (.Y(_03896_),
    .B1(net3081),
    .B2(\core.work.registers.genblk1[5].latch[29] ),
    .A2(net3086),
    .A1(\core.work.registers.genblk1[3].latch[29] ));
 sg13g2_a22oi_1 _09656_ (.Y(_03897_),
    .B1(net3076),
    .B2(\core.work.registers.genblk1[9].latch[29] ),
    .A2(net3121),
    .A1(\core.work.registers.genblk1[7].latch[29] ));
 sg13g2_a22oi_1 _09657_ (.Y(_03898_),
    .B1(net3096),
    .B2(\core.work.registers.genblk1[11].latch[29] ),
    .A2(net3116),
    .A1(\core.work.registers.genblk1[4].latch[29] ));
 sg13g2_nand4_1 _09658_ (.B(_03896_),
    .C(_03897_),
    .A(_03895_),
    .Y(_03899_),
    .D(_03898_));
 sg13g2_a22oi_1 _09659_ (.Y(_03900_),
    .B1(net3091),
    .B2(\core.work.registers.genblk1[12].latch[29] ),
    .A2(net3101),
    .A1(\core.work.registers.genblk1[14].latch[29] ));
 sg13g2_a22oi_1 _09660_ (.Y(_03901_),
    .B1(net3111),
    .B2(\core.work.registers.genblk1[2].latch[29] ),
    .A2(net3126),
    .A1(\core.work.registers.genblk1[8].latch[29] ));
 sg13g2_a22oi_1 _09661_ (.Y(_03902_),
    .B1(net3071),
    .B2(\core.work.registers.genblk1[15].latch[29] ),
    .A2(net3131),
    .A1(\core.work.registers.genblk1[10].latch[29] ));
 sg13g2_nand4_1 _09662_ (.B(_03900_),
    .C(_03901_),
    .A(_03894_),
    .Y(_03903_),
    .D(_03902_));
 sg13g2_nor2_2 _09663_ (.A(_03899_),
    .B(_03903_),
    .Y(_03904_));
 sg13g2_nor2_1 _09664_ (.A(_03893_),
    .B(_03904_),
    .Y(_03905_));
 sg13g2_nand2_1 _09665_ (.Y(_03906_),
    .A(net2913),
    .B(_03905_));
 sg13g2_xnor2_1 _09666_ (.Y(_03907_),
    .A(net3359),
    .B(_03906_));
 sg13g2_xor2_1 _09667_ (.B(_03907_),
    .A(_03892_),
    .X(_03908_));
 sg13g2_o21ai_1 _09668_ (.B1(net2762),
    .Y(_03909_),
    .A1(net2898),
    .A2(_02090_));
 sg13g2_a21oi_2 _09669_ (.B1(_03909_),
    .Y(_03910_),
    .A2(_03908_),
    .A1(net2898));
 sg13g2_a21o_1 _09670_ (.A2(net2783),
    .A1(net512),
    .B1(_03910_),
    .X(_00488_));
 sg13g2_and2_1 _09671_ (.A(_03888_),
    .B(_03907_),
    .X(_03911_));
 sg13g2_inv_1 _09672_ (.Y(_03912_),
    .A(_03911_));
 sg13g2_a21oi_1 _09673_ (.A1(_03867_),
    .A2(_03870_),
    .Y(_03913_),
    .B1(_03912_));
 sg13g2_a21oi_1 _09674_ (.A1(_03887_),
    .A2(_03906_),
    .Y(_03914_),
    .B1(_00605_));
 sg13g2_nor2_1 _09675_ (.A(_03913_),
    .B(_03914_),
    .Y(_03915_));
 sg13g2_a21oi_1 _09676_ (.A1(net3473),
    .A2(\core.work.registers.genblk1[1].latch[30] ),
    .Y(_03916_),
    .B1(net3197));
 sg13g2_a22oi_1 _09677_ (.Y(_03917_),
    .B1(net3096),
    .B2(\core.work.registers.genblk1[11].latch[30] ),
    .A2(net3121),
    .A1(\core.work.registers.genblk1[7].latch[30] ));
 sg13g2_nand2_1 _09678_ (.Y(_03918_),
    .A(\core.work.registers.genblk1[6].latch[30] ),
    .B(net3106));
 sg13g2_a22oi_1 _09679_ (.Y(_03919_),
    .B1(net3081),
    .B2(\core.work.registers.genblk1[5].latch[30] ),
    .A2(net3131),
    .A1(\core.work.registers.genblk1[10].latch[30] ));
 sg13g2_a22oi_1 _09680_ (.Y(_03920_),
    .B1(net3086),
    .B2(\core.work.registers.genblk1[3].latch[30] ),
    .A2(net3116),
    .A1(\core.work.registers.genblk1[4].latch[30] ));
 sg13g2_a22oi_1 _09681_ (.Y(_03921_),
    .B1(net3076),
    .B2(\core.work.registers.genblk1[9].latch[30] ),
    .A2(net3091),
    .A1(\core.work.registers.genblk1[12].latch[30] ));
 sg13g2_a21oi_1 _09682_ (.A1(\core.work.registers.genblk1[8].latch[30] ),
    .A2(net3126),
    .Y(_03922_),
    .B1(net3321));
 sg13g2_a22oi_1 _09683_ (.Y(_03923_),
    .B1(net3101),
    .B2(\core.work.registers.genblk1[14].latch[30] ),
    .A2(net3111),
    .A1(\core.work.registers.genblk1[2].latch[30] ));
 sg13g2_nand4_1 _09684_ (.B(_03921_),
    .C(_03922_),
    .A(_03920_),
    .Y(_03924_),
    .D(_03923_));
 sg13g2_a22oi_1 _09685_ (.Y(_03925_),
    .B1(net3066),
    .B2(\core.work.registers.genblk1[13].latch[30] ),
    .A2(net3071),
    .A1(\core.work.registers.genblk1[15].latch[30] ));
 sg13g2_nand4_1 _09686_ (.B(_03918_),
    .C(_03919_),
    .A(_03917_),
    .Y(_03926_),
    .D(_03925_));
 sg13g2_nor2_1 _09687_ (.A(_03924_),
    .B(_03926_),
    .Y(_03927_));
 sg13g2_nor2_2 _09688_ (.A(_03916_),
    .B(_03927_),
    .Y(_03928_));
 sg13g2_nand2_1 _09689_ (.Y(_03929_),
    .A(net2913),
    .B(_03928_));
 sg13g2_xnor2_1 _09690_ (.Y(_03930_),
    .A(net3360),
    .B(_03929_));
 sg13g2_o21ai_1 _09691_ (.B1(_03930_),
    .Y(_03931_),
    .A1(_03913_),
    .A2(_03914_));
 sg13g2_xor2_1 _09692_ (.B(_03930_),
    .A(_03915_),
    .X(_03932_));
 sg13g2_o21ai_1 _09693_ (.B1(net2763),
    .Y(_03933_),
    .A1(net2898),
    .A2(_02153_));
 sg13g2_a21oi_2 _09694_ (.B1(_03933_),
    .Y(_03934_),
    .A2(_03932_),
    .A1(net2902));
 sg13g2_a21o_1 _09695_ (.A2(net2784),
    .A1(net592),
    .B1(_03934_),
    .X(_00489_));
 sg13g2_nand2_1 _09696_ (.Y(_03935_),
    .A(net621),
    .B(net2784));
 sg13g2_nand3_1 _09697_ (.B(net2914),
    .C(_03928_),
    .A(net3443),
    .Y(_03936_));
 sg13g2_a21oi_1 _09698_ (.A1(net3475),
    .A2(\core.work.registers.genblk1[1].latch[31] ),
    .Y(_03937_),
    .B1(net3197));
 sg13g2_a22oi_1 _09699_ (.Y(_03938_),
    .B1(net3091),
    .B2(\core.work.registers.genblk1[12].latch[31] ),
    .A2(net3116),
    .A1(\core.work.registers.genblk1[4].latch[31] ));
 sg13g2_nand2_1 _09700_ (.Y(_03939_),
    .A(\core.work.registers.genblk1[3].latch[31] ),
    .B(net3086));
 sg13g2_a22oi_1 _09701_ (.Y(_03940_),
    .B1(net3081),
    .B2(\core.work.registers.genblk1[5].latch[31] ),
    .A2(net3106),
    .A1(\core.work.registers.genblk1[6].latch[31] ));
 sg13g2_a22oi_1 _09702_ (.Y(_03941_),
    .B1(net3111),
    .B2(\core.work.registers.genblk1[2].latch[31] ),
    .A2(net3121),
    .A1(\core.work.registers.genblk1[7].latch[31] ));
 sg13g2_a21oi_1 _09703_ (.A1(\core.work.registers.genblk1[14].latch[31] ),
    .A2(net3101),
    .Y(_03942_),
    .B1(net3324));
 sg13g2_a22oi_1 _09704_ (.Y(_03943_),
    .B1(net3066),
    .B2(\core.work.registers.genblk1[13].latch[31] ),
    .A2(net3126),
    .A1(\core.work.registers.genblk1[8].latch[31] ));
 sg13g2_nand4_1 _09705_ (.B(_03941_),
    .C(_03942_),
    .A(_03940_),
    .Y(_03944_),
    .D(_03943_));
 sg13g2_a22oi_1 _09706_ (.Y(_03945_),
    .B1(net3076),
    .B2(\core.work.registers.genblk1[9].latch[31] ),
    .A2(net3096),
    .A1(\core.work.registers.genblk1[11].latch[31] ));
 sg13g2_a22oi_1 _09707_ (.Y(_03946_),
    .B1(net3071),
    .B2(\core.work.registers.genblk1[15].latch[31] ),
    .A2(net3131),
    .A1(\core.work.registers.genblk1[10].latch[31] ));
 sg13g2_nand4_1 _09708_ (.B(_03939_),
    .C(_03945_),
    .A(_03938_),
    .Y(_03947_),
    .D(_03946_));
 sg13g2_nor2_1 _09709_ (.A(_03944_),
    .B(_03947_),
    .Y(_03948_));
 sg13g2_nor2_2 _09710_ (.A(_03937_),
    .B(_03948_),
    .Y(_03949_));
 sg13g2_nand2_1 _09711_ (.Y(_03950_),
    .A(net2914),
    .B(_03949_));
 sg13g2_xnor2_1 _09712_ (.Y(_03951_),
    .A(net3360),
    .B(_03950_));
 sg13g2_and3_1 _09713_ (.X(_03952_),
    .A(_03931_),
    .B(_03936_),
    .C(_03951_));
 sg13g2_a21oi_1 _09714_ (.A1(_03931_),
    .A2(_03936_),
    .Y(_03953_),
    .B1(_03951_));
 sg13g2_nor3_1 _09715_ (.A(net2908),
    .B(_03952_),
    .C(_03953_),
    .Y(_03954_));
 sg13g2_o21ai_1 _09716_ (.B1(net2763),
    .Y(_03955_),
    .A1(net2902),
    .A2(_02110_));
 sg13g2_o21ai_1 _09717_ (.B1(_03935_),
    .Y(_00490_),
    .A1(_03954_),
    .A2(_03955_));
 sg13g2_mux2_1 _09718_ (.A0(net458),
    .A1(_01325_),
    .S(_01327_),
    .X(_00491_));
 sg13g2_nor4_2 _09719_ (.A(net3538),
    .B(\core.work.alu.sval2[31] ),
    .C(\core.work.alu.sval2[18] ),
    .Y(_03956_),
    .D(\core.work.alu.sval2[17] ));
 sg13g2_nor4_2 _09720_ (.A(\core.work.alu.sval2[30] ),
    .B(net3540),
    .C(\core.work.alu.sval2[28] ),
    .Y(_03957_),
    .D(\core.work.alu.sval2[27] ));
 sg13g2_nand4_1 _09721_ (.B(_02072_),
    .C(_03956_),
    .A(_02070_),
    .Y(_03958_),
    .D(_03957_));
 sg13g2_nor3_2 _09722_ (.A(net3535),
    .B(_02066_),
    .C(_03958_),
    .Y(_03959_));
 sg13g2_o21ai_1 _09723_ (.B1(_03959_),
    .Y(_03960_),
    .A1(_01309_),
    .A2(_01713_));
 sg13g2_nor2b_2 _09724_ (.A(_01301_),
    .B_N(_01711_),
    .Y(_03961_));
 sg13g2_nand2b_1 _09725_ (.Y(_03962_),
    .B(_01711_),
    .A_N(_01301_));
 sg13g2_a21o_1 _09726_ (.A2(_03961_),
    .A1(_01308_),
    .B1(_03959_),
    .X(_03963_));
 sg13g2_nand3_1 _09727_ (.B(_03960_),
    .C(_03963_),
    .A(net3305),
    .Y(_03964_));
 sg13g2_nand2_1 _09728_ (.Y(_03965_),
    .A(_01707_),
    .B(_03964_));
 sg13g2_nor2_1 _09729_ (.A(_01715_),
    .B(_03962_),
    .Y(_03966_));
 sg13g2_nand2b_1 _09730_ (.Y(_03967_),
    .B(_03966_),
    .A_N(_01295_));
 sg13g2_nand3_1 _09731_ (.B(_01714_),
    .C(_01720_),
    .A(_01290_),
    .Y(_03968_));
 sg13g2_nor2_1 _09732_ (.A(_01297_),
    .B(_03962_),
    .Y(_03969_));
 sg13g2_a21oi_2 _09733_ (.B1(net2959),
    .Y(_03970_),
    .A2(_01718_),
    .A1(_01714_));
 sg13g2_a21o_1 _09734_ (.A2(_01718_),
    .A1(_01714_),
    .B1(net2959),
    .X(_03971_));
 sg13g2_nor2_1 _09735_ (.A(net3538),
    .B(net3560),
    .Y(_03972_));
 sg13g2_nand3_1 _09736_ (.B(_01833_),
    .C(net3290),
    .A(net3545),
    .Y(_03973_));
 sg13g2_nand2_1 _09737_ (.Y(_03974_),
    .A(net2963),
    .B(_03973_));
 sg13g2_o21ai_1 _09738_ (.B1(_03974_),
    .Y(_03975_),
    .A1(net3538),
    .A2(net2966));
 sg13g2_o21ai_1 _09739_ (.B1(net2858),
    .Y(_03976_),
    .A1(_00141_),
    .A2(_03975_));
 sg13g2_and2_1 _09740_ (.A(_01314_),
    .B(_03961_),
    .X(_03977_));
 sg13g2_nand2_2 _09741_ (.Y(_03978_),
    .A(_01314_),
    .B(_03961_));
 sg13g2_nor3_1 _09742_ (.A(_01308_),
    .B(_01713_),
    .C(_01714_),
    .Y(_03979_));
 sg13g2_o21ai_1 _09743_ (.B1(_01712_),
    .Y(_03980_),
    .A1(_01296_),
    .A2(_01314_));
 sg13g2_nor2_1 _09744_ (.A(_01297_),
    .B(_01719_),
    .Y(_03981_));
 sg13g2_a21oi_1 _09745_ (.A1(_03973_),
    .A2(net2939),
    .Y(_03982_),
    .B1(net2951));
 sg13g2_o21ai_1 _09746_ (.B1(_03982_),
    .Y(_03983_),
    .A1(_00144_),
    .A2(_03978_));
 sg13g2_nor2b_1 _09747_ (.A(net3560),
    .B_N(net3538),
    .Y(_03984_));
 sg13g2_nand2_1 _09748_ (.Y(_03985_),
    .A(net3539),
    .B(_00590_));
 sg13g2_and3_1 _09749_ (.X(_03986_),
    .A(net3546),
    .B(net3295),
    .C(net3288));
 sg13g2_nand3_1 _09750_ (.B(net3295),
    .C(net3287),
    .A(net3546),
    .Y(_03987_));
 sg13g2_and2_2 _09751_ (.A(_00143_),
    .B(_03182_),
    .X(_03988_));
 sg13g2_nand2_1 _09752_ (.Y(_03989_),
    .A(_00143_),
    .B(_03182_));
 sg13g2_nor2_2 _09753_ (.A(_01717_),
    .B(_03989_),
    .Y(_03990_));
 sg13g2_nand2_1 _09754_ (.Y(_03991_),
    .A(_01716_),
    .B(_03988_));
 sg13g2_a21oi_1 _09755_ (.A1(net3059),
    .A2(_03990_),
    .Y(_03992_),
    .B1(_03983_));
 sg13g2_nor2_2 _09756_ (.A(_01297_),
    .B(_01713_),
    .Y(_03993_));
 sg13g2_nand2_2 _09757_ (.Y(_03994_),
    .A(_01296_),
    .B(_01712_));
 sg13g2_a21oi_1 _09758_ (.A1(_03973_),
    .A2(net2935),
    .Y(_03995_),
    .B1(net2947));
 sg13g2_o21ai_1 _09759_ (.B1(_03995_),
    .Y(_03996_),
    .A1(net3538),
    .A2(net2935));
 sg13g2_o21ai_1 _09760_ (.B1(_03996_),
    .Y(_03997_),
    .A1(_03970_),
    .A2(_03975_));
 sg13g2_inv_1 _09761_ (.Y(_03998_),
    .A(_03997_));
 sg13g2_a22oi_1 _09762_ (.Y(_03999_),
    .B1(_03998_),
    .B2(_00141_),
    .A2(_03992_),
    .A1(_03976_));
 sg13g2_nor2_2 _09763_ (.A(net2955),
    .B(net2940),
    .Y(_04000_));
 sg13g2_nand3_1 _09764_ (.B(_01308_),
    .C(_01711_),
    .A(net3441),
    .Y(_04001_));
 sg13g2_nand3_1 _09765_ (.B(_04000_),
    .C(_04001_),
    .A(net2860),
    .Y(_04002_));
 sg13g2_a21oi_1 _09766_ (.A1(_01309_),
    .A2(_01720_),
    .Y(_04003_),
    .B1(_03966_));
 sg13g2_nor2_1 _09767_ (.A(_01723_),
    .B(_04002_),
    .Y(_04004_));
 sg13g2_and3_2 _09768_ (.X(_04005_),
    .A(net2943),
    .B(_04003_),
    .C(_04004_));
 sg13g2_nand3_1 _09769_ (.B(_04003_),
    .C(_04004_),
    .A(net2943),
    .Y(_04006_));
 sg13g2_nor2_1 _09770_ (.A(_00145_),
    .B(net3059),
    .Y(_04007_));
 sg13g2_a21oi_1 _09771_ (.A1(_00730_),
    .A2(net3059),
    .Y(_04008_),
    .B1(_04007_));
 sg13g2_nand2_1 _09772_ (.Y(_04009_),
    .A(_01722_),
    .B(_03988_));
 sg13g2_inv_2 _09773_ (.Y(_04010_),
    .A(net2831));
 sg13g2_and2_2 _09774_ (.A(_01314_),
    .B(_01720_),
    .X(_04011_));
 sg13g2_nand2_2 _09775_ (.Y(_04012_),
    .A(_01314_),
    .B(_01720_));
 sg13g2_nand2b_1 _09776_ (.Y(_04013_),
    .B(net3058),
    .A_N(_00147_));
 sg13g2_o21ai_1 _09777_ (.B1(_04013_),
    .Y(_04014_),
    .A1(_00146_),
    .A2(net3058));
 sg13g2_and2_2 _09778_ (.A(_01722_),
    .B(_03989_),
    .X(_04015_));
 sg13g2_nand2_1 _09779_ (.Y(_04016_),
    .A(_01722_),
    .B(net2853));
 sg13g2_a22oi_1 _09780_ (.Y(_04017_),
    .B1(_04014_),
    .B2(_04015_),
    .A2(net2927),
    .A1(_01303_));
 sg13g2_o21ai_1 _09781_ (.B1(_04017_),
    .Y(_04018_),
    .A1(_04008_),
    .A2(net2832));
 sg13g2_nand2_1 _09782_ (.Y(_04019_),
    .A(_01296_),
    .B(_01720_));
 sg13g2_nand2_1 _09783_ (.Y(_04020_),
    .A(net3483),
    .B(net3287));
 sg13g2_nand2_1 _09784_ (.Y(_04021_),
    .A(net3478),
    .B(net3291));
 sg13g2_nor2_1 _09785_ (.A(net3539),
    .B(_00590_),
    .Y(_04022_));
 sg13g2_nand2b_1 _09786_ (.Y(_04023_),
    .B(net3562),
    .A_N(net3539));
 sg13g2_a22oi_1 _09787_ (.Y(_04024_),
    .B1(net3053),
    .B2(net3481),
    .A2(net3289),
    .A1(net3485));
 sg13g2_nand4_1 _09788_ (.B(_04020_),
    .C(_04021_),
    .A(net3558),
    .Y(_04025_),
    .D(_04024_));
 sg13g2_nand2_1 _09789_ (.Y(_04026_),
    .A(net3488),
    .B(net3287));
 sg13g2_a21oi_1 _09790_ (.A1(\core.e2m_addr[8] ),
    .A2(net3290),
    .Y(_04027_),
    .B1(net3558));
 sg13g2_a22oi_1 _09791_ (.Y(_04028_),
    .B1(net3054),
    .B2(net3487),
    .A2(net3291),
    .A1(\core.e2m_addr[11] ));
 sg13g2_nand3_1 _09792_ (.B(_04027_),
    .C(_04028_),
    .A(_04026_),
    .Y(_04029_));
 sg13g2_nand3_1 _09793_ (.B(_04025_),
    .C(_04029_),
    .A(net3552),
    .Y(_04030_));
 sg13g2_nand2_2 _09794_ (.Y(_04031_),
    .A(_00592_),
    .B(net3558));
 sg13g2_a22oi_1 _09795_ (.Y(_04032_),
    .B1(net3290),
    .B2(net3495),
    .A2(net3291),
    .A1(\core.e2m_addr[7] ));
 sg13g2_a22oi_1 _09796_ (.Y(_04033_),
    .B1(net3053),
    .B2(\core.e2m_addr[6] ),
    .A2(net3287),
    .A1(net3493));
 sg13g2_a21oi_1 _09797_ (.A1(_04032_),
    .A2(_04033_),
    .Y(_04034_),
    .B1(_04031_));
 sg13g2_a22oi_1 _09798_ (.Y(_04035_),
    .B1(net3289),
    .B2(net3500),
    .A2(net3292),
    .A1(net3496));
 sg13g2_a22oi_1 _09799_ (.Y(_04036_),
    .B1(net3054),
    .B2(net3497),
    .A2(net3287),
    .A1(net3499));
 sg13g2_a21oi_1 _09800_ (.A1(_04035_),
    .A2(_04036_),
    .Y(_04037_),
    .B1(_01834_));
 sg13g2_nand2_1 _09801_ (.Y(_04038_),
    .A(net3451),
    .B(net3289));
 sg13g2_a21oi_1 _09802_ (.A1(\core.e2m_addr[27] ),
    .A2(net3292),
    .Y(_04039_),
    .B1(net3559));
 sg13g2_a22oi_1 _09803_ (.Y(_04040_),
    .B1(net3053),
    .B2(\core.e2m_addr[26] ),
    .A2(net3288),
    .A1(net3450));
 sg13g2_nand3_1 _09804_ (.B(_04039_),
    .C(_04040_),
    .A(_04038_),
    .Y(_04041_));
 sg13g2_nand2_1 _09805_ (.Y(_04042_),
    .A(net3445),
    .B(net3288));
 sg13g2_nand2_1 _09806_ (.Y(_04043_),
    .A(net3447),
    .B(net3289));
 sg13g2_a22oi_1 _09807_ (.Y(_04044_),
    .B1(net3053),
    .B2(net3444),
    .A2(net3292),
    .A1(\core.e2m_addr[31] ));
 sg13g2_nand4_1 _09808_ (.B(_04042_),
    .C(_04043_),
    .A(net3559),
    .Y(_04045_),
    .D(_04044_));
 sg13g2_nand3_1 _09809_ (.B(_04041_),
    .C(_04045_),
    .A(net3554),
    .Y(_04046_));
 sg13g2_a22oi_1 _09810_ (.Y(_04047_),
    .B1(net3053),
    .B2(net3456),
    .A2(net3291),
    .A1(net3454));
 sg13g2_a22oi_1 _09811_ (.Y(_04048_),
    .B1(net3287),
    .B2(net3458),
    .A2(net3289),
    .A1(net3466));
 sg13g2_a21oi_1 _09812_ (.A1(_04047_),
    .A2(_04048_),
    .Y(_04049_),
    .B1(_04031_));
 sg13g2_a22oi_1 _09813_ (.Y(_04050_),
    .B1(net3287),
    .B2(net3469),
    .A2(net3289),
    .A1(net3471));
 sg13g2_a22oi_1 _09814_ (.Y(_04051_),
    .B1(net3053),
    .B2(net3468),
    .A2(net3291),
    .A1(\core.e2m_addr[19] ));
 sg13g2_a21oi_1 _09815_ (.A1(_04050_),
    .A2(_04051_),
    .Y(_04052_),
    .B1(_01834_));
 sg13g2_nor3_1 _09816_ (.A(_00596_),
    .B(_04049_),
    .C(_04052_),
    .Y(_04053_));
 sg13g2_nor3_1 _09817_ (.A(net3549),
    .B(_04034_),
    .C(_04037_),
    .Y(_04054_));
 sg13g2_a221oi_1 _09818_ (.B2(_04030_),
    .C1(_04019_),
    .B1(_04054_),
    .A1(_04046_),
    .Y(_04055_),
    .A2(_04053_));
 sg13g2_nor4_1 _09819_ (.A(_03999_),
    .B(net2795),
    .C(_04018_),
    .D(_04055_),
    .Y(_04056_));
 sg13g2_nand3_1 _09820_ (.B(_03968_),
    .C(_04056_),
    .A(_03967_),
    .Y(_04057_));
 sg13g2_o21ai_1 _09821_ (.B1(net3309),
    .Y(_04058_),
    .A1(_01303_),
    .A2(net2791));
 sg13g2_nand2b_1 _09822_ (.Y(_04059_),
    .B(_04057_),
    .A_N(_04058_));
 sg13g2_nand3_1 _09823_ (.B(net3161),
    .C(_03964_),
    .A(_01707_),
    .Y(_04060_));
 sg13g2_a21oi_1 _09824_ (.A1(net2843),
    .A2(_03230_),
    .Y(_04061_),
    .B1(_04060_));
 sg13g2_a22oi_1 _09825_ (.Y(_00492_),
    .B1(_04059_),
    .B2(_04061_),
    .A2(net2750),
    .A1(_00589_));
 sg13g2_nand2b_1 _09826_ (.Y(_04062_),
    .B(_03251_),
    .A_N(net2890));
 sg13g2_a21oi_1 _09827_ (.A1(net3493),
    .A2(_01686_),
    .Y(_04063_),
    .B1(_00143_));
 sg13g2_a21oi_1 _09828_ (.A1(net2890),
    .A2(_04063_),
    .Y(_04064_),
    .B1(net3330));
 sg13g2_a21oi_2 _09829_ (.B1(_01709_),
    .Y(_04065_),
    .A2(_04064_),
    .A1(_04062_));
 sg13g2_a21oi_1 _09830_ (.A1(_00141_),
    .A2(net3065),
    .Y(_04066_),
    .B1(_01717_));
 sg13g2_nand2_1 _09831_ (.Y(_04067_),
    .A(_00147_),
    .B(net3065));
 sg13g2_a21oi_1 _09832_ (.A1(_01722_),
    .A2(_04067_),
    .Y(_04068_),
    .B1(_04066_));
 sg13g2_nand2_1 _09833_ (.Y(_04069_),
    .A(_00145_),
    .B(net3058));
 sg13g2_nand2_1 _09834_ (.Y(_04070_),
    .A(_00148_),
    .B(net3065));
 sg13g2_nand2_1 _09835_ (.Y(_04071_),
    .A(_00146_),
    .B(net3058));
 sg13g2_nand2_1 _09836_ (.Y(_04072_),
    .A(_04070_),
    .B(_04071_));
 sg13g2_nor2_1 _09837_ (.A(net2827),
    .B(_04072_),
    .Y(_04073_));
 sg13g2_nand2_1 _09838_ (.Y(_04074_),
    .A(net2964),
    .B(net3065));
 sg13g2_o21ai_1 _09839_ (.B1(_04074_),
    .Y(_04075_),
    .A1(_00590_),
    .A2(net2964));
 sg13g2_nand2b_1 _09840_ (.Y(_04076_),
    .B(_00145_),
    .A_N(_04075_));
 sg13g2_a21oi_1 _09841_ (.A1(_00731_),
    .A2(_04075_),
    .Y(_04077_),
    .B1(net2859));
 sg13g2_o21ai_1 _09842_ (.B1(net2947),
    .Y(_04078_),
    .A1(_00143_),
    .A2(_03978_));
 sg13g2_a21oi_1 _09843_ (.A1(net2940),
    .A2(net3059),
    .Y(_04079_),
    .B1(_04078_));
 sg13g2_nor2_1 _09844_ (.A(_00145_),
    .B(_04079_),
    .Y(_04080_));
 sg13g2_a21oi_1 _09845_ (.A1(net3058),
    .A2(net2935),
    .Y(_04081_),
    .B1(net2947));
 sg13g2_o21ai_1 _09846_ (.B1(_04081_),
    .Y(_04082_),
    .A1(net3561),
    .A2(net2935));
 sg13g2_xnor2_1 _09847_ (.Y(_04083_),
    .A(_01204_),
    .B(_01205_));
 sg13g2_o21ai_1 _09848_ (.B1(_04082_),
    .Y(_04084_),
    .A1(net2924),
    .A2(_04083_));
 sg13g2_nor4_1 _09849_ (.A(net2796),
    .B(_04073_),
    .C(_04080_),
    .D(_04084_),
    .Y(_04085_));
 sg13g2_nor2b_1 _09850_ (.A(_04068_),
    .B_N(_04069_),
    .Y(_04086_));
 sg13g2_a22oi_1 _09851_ (.Y(_04087_),
    .B1(_04086_),
    .B2(_03988_),
    .A2(_04077_),
    .A1(_04076_));
 sg13g2_nand2_1 _09852_ (.Y(_04088_),
    .A(net3539),
    .B(net3500));
 sg13g2_xor2_1 _09853_ (.B(_04088_),
    .A(_01204_),
    .X(_04089_));
 sg13g2_a221oi_1 _09854_ (.B2(net2796),
    .C1(net3301),
    .B1(_04089_),
    .A1(_04085_),
    .Y(_04090_),
    .A2(_04087_));
 sg13g2_nor3_1 _09855_ (.A(net2749),
    .B(_04065_),
    .C(_04090_),
    .Y(_04091_));
 sg13g2_a21oi_1 _09856_ (.A1(_00591_),
    .A2(net2749),
    .Y(_00493_),
    .B1(_04091_));
 sg13g2_nand2_1 _09857_ (.Y(_04092_),
    .A(_01716_),
    .B(net2853));
 sg13g2_nor3_1 _09858_ (.A(_00141_),
    .B(net3065),
    .C(net2824),
    .Y(_04093_));
 sg13g2_a21o_1 _09859_ (.A2(_04014_),
    .A1(_04010_),
    .B1(_04093_),
    .X(_04094_));
 sg13g2_xor2_1 _09860_ (.B(_01209_),
    .A(_01206_),
    .X(_04095_));
 sg13g2_nand2_1 _09861_ (.Y(_04096_),
    .A(_04011_),
    .B(_04095_));
 sg13g2_nand3_1 _09862_ (.B(net3295),
    .C(net3054),
    .A(net3545),
    .Y(_04097_));
 sg13g2_o21ai_1 _09863_ (.B1(net2948),
    .Y(_04098_),
    .A1(net3556),
    .A2(net2953));
 sg13g2_a21oi_1 _09864_ (.A1(net2940),
    .A2(_04097_),
    .Y(_04099_),
    .B1(_04098_));
 sg13g2_o21ai_1 _09865_ (.B1(_04096_),
    .Y(_04100_),
    .A1(_00147_),
    .A2(_04099_));
 sg13g2_nor3_1 _09866_ (.A(net2795),
    .B(_04094_),
    .C(_04100_),
    .Y(_04101_));
 sg13g2_nor2_1 _09867_ (.A(net3557),
    .B(net2964),
    .Y(_04102_));
 sg13g2_a21oi_1 _09868_ (.A1(net2964),
    .A2(_04097_),
    .Y(_04103_),
    .B1(_04102_));
 sg13g2_xnor2_1 _09869_ (.Y(_04104_),
    .A(_00147_),
    .B(_04103_));
 sg13g2_nor2_1 _09870_ (.A(net3557),
    .B(net2935),
    .Y(_04105_));
 sg13g2_a21oi_1 _09871_ (.A1(net2935),
    .A2(_04097_),
    .Y(_04106_),
    .B1(_04105_));
 sg13g2_nand2_1 _09872_ (.Y(_04107_),
    .A(_00153_),
    .B(net3065));
 sg13g2_nand2_1 _09873_ (.Y(_04108_),
    .A(_00148_),
    .B(net3058));
 sg13g2_nand2_1 _09874_ (.Y(_04109_),
    .A(_04107_),
    .B(_04108_));
 sg13g2_nor2b_1 _09875_ (.A(_04007_),
    .B_N(_04013_),
    .Y(_04110_));
 sg13g2_nand2b_1 _09876_ (.Y(_04111_),
    .B(_03990_),
    .A_N(_04110_));
 sg13g2_o21ai_1 _09877_ (.B1(_04111_),
    .Y(_04112_),
    .A1(net2827),
    .A2(_04109_));
 sg13g2_a221oi_1 _09878_ (.B2(net2951),
    .C1(_04112_),
    .B1(_04106_),
    .A1(net2857),
    .Y(_04113_),
    .A2(_04104_));
 sg13g2_o21ai_1 _09879_ (.B1(_01202_),
    .Y(_04114_),
    .A1(_01203_),
    .A2(_04088_));
 sg13g2_xor2_1 _09880_ (.B(_04114_),
    .A(_01209_),
    .X(_04115_));
 sg13g2_a221oi_1 _09881_ (.B2(net2795),
    .C1(net3302),
    .B1(_04115_),
    .A1(_04101_),
    .Y(_04116_),
    .A2(_04113_));
 sg13g2_nor2_1 _09882_ (.A(net2890),
    .B(_03275_),
    .Y(_04117_));
 sg13g2_a21o_1 _09883_ (.A2(net3029),
    .A1(net3490),
    .B1(net3329),
    .X(_04118_));
 sg13g2_a21oi_2 _09884_ (.B1(net3329),
    .Y(_04119_),
    .A2(net3029),
    .A1(net3492));
 sg13g2_a21oi_1 _09885_ (.A1(net3555),
    .A2(_02134_),
    .Y(_04120_),
    .B1(_04117_));
 sg13g2_nand2_2 _09886_ (.Y(_04121_),
    .A(\core.f2e_inst[0] ),
    .B(_00582_));
 sg13g2_and2_1 _09887_ (.A(net3504),
    .B(\core.f2e_inst[14] ),
    .X(_04122_));
 sg13g2_nand4_1 _09888_ (.B(_00582_),
    .C(_00151_),
    .A(\core.f2e_inst[0] ),
    .Y(_04123_),
    .D(_04122_));
 sg13g2_inv_1 _09889_ (.Y(_04124_),
    .A(_04123_));
 sg13g2_nor3_1 _09890_ (.A(\core.f2e_inst[7] ),
    .B(_00695_),
    .C(\core.f2e_inst[9] ),
    .Y(_04125_));
 sg13g2_nand3b_1 _09891_ (.B(_00152_),
    .C(_04125_),
    .Y(_04126_),
    .A_N(net3508));
 sg13g2_nand2_1 _09892_ (.Y(_04127_),
    .A(_04124_),
    .B(_04126_));
 sg13g2_nand2_1 _09893_ (.Y(_04128_),
    .A(net3504),
    .B(_00705_));
 sg13g2_nor3_2 _09894_ (.A(\core.f2e_inst[15] ),
    .B(_04121_),
    .C(_04128_),
    .Y(_04129_));
 sg13g2_nor3_2 _09895_ (.A(_00151_),
    .B(_04121_),
    .C(_04128_),
    .Y(_04130_));
 sg13g2_nor2_2 _09896_ (.A(_04129_),
    .B(_04130_),
    .Y(_04131_));
 sg13g2_nand3_1 _09897_ (.B(net2852),
    .C(_04131_),
    .A(net3337),
    .Y(_04132_));
 sg13g2_nor2_1 _09898_ (.A(\core.f2e_inst[4] ),
    .B(net3511),
    .Y(_04133_));
 sg13g2_nand4_1 _09899_ (.B(_00683_),
    .C(_00150_),
    .A(_00680_),
    .Y(_04134_),
    .D(_04133_));
 sg13g2_nor3_2 _09900_ (.A(net3513),
    .B(_00582_),
    .C(net3504),
    .Y(_04135_));
 sg13g2_nor2_1 _09901_ (.A(\core.f2e_inst[14] ),
    .B(_00708_),
    .Y(_04136_));
 sg13g2_and2_2 _09902_ (.A(_04135_),
    .B(_04136_),
    .X(_04137_));
 sg13g2_nand2b_1 _09903_ (.Y(_04138_),
    .B(_04137_),
    .A_N(_04134_));
 sg13g2_nand2b_2 _09904_ (.Y(_04139_),
    .B(_00701_),
    .A_N(_04138_));
 sg13g2_a21oi_1 _09905_ (.A1(net3507),
    .A2(net3506),
    .Y(_04140_),
    .B1(_04138_));
 sg13g2_nor2_1 _09906_ (.A(_04132_),
    .B(_04140_),
    .Y(_04141_));
 sg13g2_a21oi_2 _09907_ (.B1(_04141_),
    .Y(_04142_),
    .A2(net3347),
    .A1(_00680_));
 sg13g2_a221oi_1 _09908_ (.B2(net3167),
    .C1(_04116_),
    .B1(_04142_),
    .A1(_04119_),
    .Y(_04143_),
    .A2(_04120_));
 sg13g2_nand2_1 _09909_ (.Y(_04144_),
    .A(net3497),
    .B(net2749));
 sg13g2_o21ai_1 _09910_ (.B1(_04144_),
    .Y(_00494_),
    .A1(net2749),
    .A2(_04143_));
 sg13g2_nand2_1 _09911_ (.Y(_04145_),
    .A(net3496),
    .B(net2749));
 sg13g2_xor2_1 _09912_ (.B(_01210_),
    .A(_01199_),
    .X(_04146_));
 sg13g2_nand2_1 _09913_ (.Y(_04147_),
    .A(_00020_),
    .B(net3064));
 sg13g2_nand2_1 _09914_ (.Y(_04148_),
    .A(_00153_),
    .B(net3058));
 sg13g2_nand2_1 _09915_ (.Y(_04149_),
    .A(_04147_),
    .B(_04148_));
 sg13g2_nor2_1 _09916_ (.A(net2827),
    .B(_04149_),
    .Y(_04150_));
 sg13g2_nand3_1 _09917_ (.B(net3295),
    .C(net3291),
    .A(net3545),
    .Y(_04151_));
 sg13g2_a21oi_1 _09918_ (.A1(net2936),
    .A2(_04151_),
    .Y(_04152_),
    .B1(net2947));
 sg13g2_o21ai_1 _09919_ (.B1(_04152_),
    .Y(_04153_),
    .A1(net3552),
    .A2(net2935));
 sg13g2_o21ai_1 _09920_ (.B1(_04153_),
    .Y(_04154_),
    .A1(net2832),
    .A2(_04072_));
 sg13g2_o21ai_1 _09921_ (.B1(net2947),
    .Y(_04155_),
    .A1(net3551),
    .A2(net2953));
 sg13g2_a21oi_1 _09922_ (.A1(net2940),
    .A2(_04151_),
    .Y(_04156_),
    .B1(_04155_));
 sg13g2_o21ai_1 _09923_ (.B1(net2791),
    .Y(_04157_),
    .A1(_00146_),
    .A2(_04156_));
 sg13g2_nor2_1 _09924_ (.A(net3552),
    .B(net2964),
    .Y(_04158_));
 sg13g2_a21oi_1 _09925_ (.A1(net2964),
    .A2(_04151_),
    .Y(_04159_),
    .B1(_04158_));
 sg13g2_a21oi_1 _09926_ (.A1(_00732_),
    .A2(_04159_),
    .Y(_04160_),
    .B1(net2859));
 sg13g2_o21ai_1 _09927_ (.B1(_04160_),
    .Y(_04161_),
    .A1(_00732_),
    .A2(_04159_));
 sg13g2_a21oi_1 _09928_ (.A1(_04067_),
    .A2(_04071_),
    .Y(_04162_),
    .B1(net2853));
 sg13g2_a21oi_1 _09929_ (.A1(_04066_),
    .A2(_04069_),
    .Y(_04163_),
    .B1(_03990_));
 sg13g2_o21ai_1 _09930_ (.B1(_04161_),
    .Y(_04164_),
    .A1(_04162_),
    .A2(_04163_));
 sg13g2_nor4_1 _09931_ (.A(_04150_),
    .B(_04154_),
    .C(_04157_),
    .D(_04164_),
    .Y(_04165_));
 sg13g2_o21ai_1 _09932_ (.B1(_04165_),
    .Y(_04166_),
    .A1(net2924),
    .A2(_04146_));
 sg13g2_a21oi_1 _09933_ (.A1(_01208_),
    .A2(_04114_),
    .Y(_04167_),
    .B1(_01207_));
 sg13g2_xnor2_1 _09934_ (.Y(_04168_),
    .A(_01199_),
    .B(_04167_));
 sg13g2_a21oi_1 _09935_ (.A1(net2795),
    .A2(_04168_),
    .Y(_04169_),
    .B1(net3302));
 sg13g2_nand2_2 _09936_ (.Y(_04170_),
    .A(net2890),
    .B(_04119_));
 sg13g2_o21ai_1 _09937_ (.B1(_04131_),
    .Y(_04171_),
    .A1(_00683_),
    .A2(net3338));
 sg13g2_a22oi_1 _09938_ (.Y(_04172_),
    .B1(_04171_),
    .B2(net3167),
    .A2(_03298_),
    .A1(net2843));
 sg13g2_o21ai_1 _09939_ (.B1(_04172_),
    .Y(_04173_),
    .A1(net3551),
    .A2(_04170_));
 sg13g2_a21oi_1 _09940_ (.A1(_04166_),
    .A2(_04169_),
    .Y(_04174_),
    .B1(_04173_));
 sg13g2_o21ai_1 _09941_ (.B1(_04145_),
    .Y(_00495_),
    .A1(net2749),
    .A2(_04174_));
 sg13g2_xor2_1 _09942_ (.B(_01213_),
    .A(_01197_),
    .X(_04175_));
 sg13g2_nor4_2 _09943_ (.A(net3538),
    .B(net3560),
    .C(net3552),
    .Y(_04176_),
    .D(net3556));
 sg13g2_inv_1 _09944_ (.Y(_04177_),
    .A(_04176_));
 sg13g2_nand2_1 _09945_ (.Y(_04178_),
    .A(net3545),
    .B(_04176_));
 sg13g2_nand2_1 _09946_ (.Y(_04179_),
    .A(net2964),
    .B(_04178_));
 sg13g2_o21ai_1 _09947_ (.B1(_04179_),
    .Y(_04180_),
    .A1(net3549),
    .A2(net2965));
 sg13g2_a21oi_1 _09948_ (.A1(_00148_),
    .A2(_04180_),
    .Y(_04181_),
    .B1(net2859));
 sg13g2_o21ai_1 _09949_ (.B1(_04181_),
    .Y(_04182_),
    .A1(_00148_),
    .A2(_04180_));
 sg13g2_o21ai_1 _09950_ (.B1(net2951),
    .Y(_04183_),
    .A1(net3549),
    .A2(net2936));
 sg13g2_a21o_1 _09951_ (.A2(_04178_),
    .A1(net2935),
    .B1(_04183_),
    .X(_04184_));
 sg13g2_nor2_1 _09952_ (.A(net3545),
    .B(_04000_),
    .Y(_04185_));
 sg13g2_a21oi_1 _09953_ (.A1(net2940),
    .A2(_04177_),
    .Y(_04186_),
    .B1(_04185_));
 sg13g2_a22oi_1 _09954_ (.Y(_04187_),
    .B1(_04186_),
    .B2(net2947),
    .A2(_04184_),
    .A1(_00148_));
 sg13g2_nor2_1 _09955_ (.A(net2832),
    .B(_04109_),
    .Y(_04188_));
 sg13g2_nand2_1 _09956_ (.Y(_04189_),
    .A(_00020_),
    .B(net3060));
 sg13g2_nand2_1 _09957_ (.Y(_04190_),
    .A(_00154_),
    .B(net3065));
 sg13g2_nand2_1 _09958_ (.Y(_04191_),
    .A(_04189_),
    .B(_04190_));
 sg13g2_nor2_1 _09959_ (.A(net2826),
    .B(_04191_),
    .Y(_04192_));
 sg13g2_o21ai_1 _09960_ (.B1(_04108_),
    .Y(_04193_),
    .A1(_00732_),
    .A2(net3058));
 sg13g2_inv_1 _09961_ (.Y(_04194_),
    .A(_04193_));
 sg13g2_nor4_1 _09962_ (.A(net2796),
    .B(_04187_),
    .C(_04188_),
    .D(_04192_),
    .Y(_04195_));
 sg13g2_o21ai_1 _09963_ (.B1(_04182_),
    .Y(_04196_),
    .A1(net2824),
    .A2(_04110_));
 sg13g2_a221oi_1 _09964_ (.B2(_03990_),
    .C1(_04196_),
    .B1(_04194_),
    .A1(net2927),
    .Y(_04197_),
    .A2(_04175_));
 sg13g2_o21ai_1 _09965_ (.B1(_01198_),
    .Y(_04198_),
    .A1(_01199_),
    .A2(_04167_));
 sg13g2_xnor2_1 _09966_ (.Y(_04199_),
    .A(_01197_),
    .B(_04198_));
 sg13g2_a221oi_1 _09967_ (.B2(net2795),
    .C1(net3301),
    .B1(_04199_),
    .A1(_04195_),
    .Y(_04200_),
    .A2(_04197_));
 sg13g2_nand2_1 _09968_ (.Y(_04201_),
    .A(net2844),
    .B(_03321_));
 sg13g2_o21ai_1 _09969_ (.B1(_04201_),
    .Y(_04202_),
    .A1(net3546),
    .A2(_04170_));
 sg13g2_nor2_1 _09970_ (.A(net3504),
    .B(_04121_),
    .Y(_04203_));
 sg13g2_and2_1 _09971_ (.A(_04136_),
    .B(_04203_),
    .X(_04204_));
 sg13g2_nand2_2 _09972_ (.Y(_04205_),
    .A(_04136_),
    .B(_04203_));
 sg13g2_nor3_2 _09973_ (.A(_00705_),
    .B(_00151_),
    .C(_04121_),
    .Y(_04206_));
 sg13g2_or3_2 _09974_ (.A(_00705_),
    .B(_00151_),
    .C(_04121_),
    .X(_04207_));
 sg13g2_nand2b_1 _09975_ (.Y(_04208_),
    .B(\core.f2e_inst[14] ),
    .A_N(net3513));
 sg13g2_nor4_2 _09976_ (.A(net3512),
    .B(net3505),
    .C(\core.f2e_inst[15] ),
    .Y(_04209_),
    .D(_04208_));
 sg13g2_nor4_2 _09977_ (.A(net3512),
    .B(net3504),
    .C(_00151_),
    .Y(_04210_),
    .D(_04208_));
 sg13g2_nor2_1 _09978_ (.A(_04209_),
    .B(_04210_),
    .Y(_04211_));
 sg13g2_and2_1 _09979_ (.A(_04207_),
    .B(_04211_),
    .X(_04212_));
 sg13g2_nand2_1 _09980_ (.Y(_04213_),
    .A(net2851),
    .B(_04212_));
 sg13g2_nand2_2 _09981_ (.Y(_04214_),
    .A(\core.f2e_inst[14] ),
    .B(_04135_));
 sg13g2_nor2_2 _09982_ (.A(_00151_),
    .B(_04214_),
    .Y(_04215_));
 sg13g2_nor3_2 _09983_ (.A(net3504),
    .B(\core.f2e_inst[15] ),
    .C(_04121_),
    .Y(_04216_));
 sg13g2_and2_1 _09984_ (.A(_00708_),
    .B(_04135_),
    .X(_04217_));
 sg13g2_nor2_1 _09985_ (.A(_04216_),
    .B(_04217_),
    .Y(_04218_));
 sg13g2_nand2b_1 _09986_ (.Y(_04219_),
    .B(_04218_),
    .A_N(_04215_));
 sg13g2_nor4_2 _09987_ (.A(_04124_),
    .B(_04137_),
    .C(_04213_),
    .Y(_04220_),
    .D(_04219_));
 sg13g2_nand2_2 _09988_ (.Y(_04221_),
    .A(_04131_),
    .B(_04220_));
 sg13g2_nand2_2 _09989_ (.Y(_04222_),
    .A(_04134_),
    .B(_04137_));
 sg13g2_or2_1 _09990_ (.X(_04223_),
    .B(_04222_),
    .A(net3506));
 sg13g2_and2_2 _09991_ (.A(net2851),
    .B(_04223_),
    .X(_04224_));
 sg13g2_nand2_1 _09992_ (.Y(_04225_),
    .A(_04123_),
    .B(_04224_));
 sg13g2_nor2_2 _09993_ (.A(net3507),
    .B(_04222_),
    .Y(_04226_));
 sg13g2_and2_1 _09994_ (.A(_00705_),
    .B(_04217_),
    .X(_04227_));
 sg13g2_nor4_2 _09995_ (.A(_04216_),
    .B(_04225_),
    .C(_04226_),
    .Y(_04228_),
    .D(_04227_));
 sg13g2_o21ai_1 _09996_ (.B1(net3162),
    .Y(_04229_),
    .A1(\core.f2e_inst[4] ),
    .A2(net3337));
 sg13g2_a21oi_2 _09997_ (.B1(_04229_),
    .Y(_04230_),
    .A2(_04228_),
    .A1(_04221_));
 sg13g2_nor4_1 _09998_ (.A(net2748),
    .B(_04200_),
    .C(_04202_),
    .D(_04230_),
    .Y(_04231_));
 sg13g2_a21oi_1 _09999_ (.A1(_00597_),
    .A2(net2748),
    .Y(_00496_),
    .B1(_04231_));
 sg13g2_a21oi_1 _10000_ (.A1(_01197_),
    .A2(_04198_),
    .Y(_04232_),
    .B1(_01196_));
 sg13g2_xnor2_1 _10001_ (.Y(_04233_),
    .A(_01194_),
    .B(_04232_));
 sg13g2_nor3_2 _10002_ (.A(net3552),
    .B(net3555),
    .C(_03985_),
    .Y(_04234_));
 sg13g2_nand2_2 _10003_ (.Y(_04235_),
    .A(net3545),
    .B(_04234_));
 sg13g2_nand2_1 _10004_ (.Y(_04236_),
    .A(net2965),
    .B(_04235_));
 sg13g2_o21ai_1 _10005_ (.B1(_04236_),
    .Y(_04237_),
    .A1(net3543),
    .A2(net2964));
 sg13g2_o21ai_1 _10006_ (.B1(net2858),
    .Y(_04238_),
    .A1(_00153_),
    .A2(_04237_));
 sg13g2_a21oi_1 _10007_ (.A1(_00153_),
    .A2(_04237_),
    .Y(_04239_),
    .B1(_04238_));
 sg13g2_a22oi_1 _10008_ (.Y(_04240_),
    .B1(net2940),
    .B2(_04235_),
    .A2(net2955),
    .A1(_00716_));
 sg13g2_a21oi_1 _10009_ (.A1(net3543),
    .A2(net2929),
    .Y(_04241_),
    .B1(_00733_));
 sg13g2_o21ai_1 _10010_ (.B1(_04241_),
    .Y(_04242_),
    .A1(_03994_),
    .A2(_04235_));
 sg13g2_o21ai_1 _10011_ (.B1(net2947),
    .Y(_04243_),
    .A1(_00153_),
    .A2(_04240_));
 sg13g2_nand2_1 _10012_ (.Y(_04244_),
    .A(_04242_),
    .B(_04243_));
 sg13g2_nand4_1 _10013_ (.B(net2853),
    .C(_04067_),
    .A(_01716_),
    .Y(_04245_),
    .D(_04071_));
 sg13g2_nand2_1 _10014_ (.Y(_04246_),
    .A(_00154_),
    .B(net3060));
 sg13g2_nand2_1 _10015_ (.Y(_04247_),
    .A(_00106_),
    .B(net3063));
 sg13g2_nand2_1 _10016_ (.Y(_04248_),
    .A(_04246_),
    .B(_04247_));
 sg13g2_nor2_1 _10017_ (.A(net2827),
    .B(_04248_),
    .Y(_04249_));
 sg13g2_nand2_1 _10018_ (.Y(_04250_),
    .A(_04070_),
    .B(_04148_));
 sg13g2_o21ai_1 _10019_ (.B1(_04245_),
    .Y(_04251_),
    .A1(_03991_),
    .A2(_04250_));
 sg13g2_o21ai_1 _10020_ (.B1(_04244_),
    .Y(_04252_),
    .A1(net2832),
    .A2(_04149_));
 sg13g2_nor4_1 _10021_ (.A(_04239_),
    .B(_04249_),
    .C(_04251_),
    .D(_04252_),
    .Y(_04253_));
 sg13g2_xnor2_1 _10022_ (.Y(_04254_),
    .A(_01194_),
    .B(_01215_));
 sg13g2_a22oi_1 _10023_ (.Y(_04255_),
    .B1(_04254_),
    .B2(net2927),
    .A2(_04233_),
    .A1(net2795));
 sg13g2_a21oi_1 _10024_ (.A1(_04253_),
    .A2(_04255_),
    .Y(_04256_),
    .B1(net3301));
 sg13g2_nand2_1 _10025_ (.Y(_04257_),
    .A(net2843),
    .B(_03340_));
 sg13g2_nor2_1 _10026_ (.A(_00699_),
    .B(_04205_),
    .Y(_04258_));
 sg13g2_a21oi_1 _10027_ (.A1(net3509),
    .A2(_04258_),
    .Y(_04259_),
    .B1(_04210_));
 sg13g2_nor4_1 _10028_ (.A(_04132_),
    .B(_04137_),
    .C(_04206_),
    .D(_04215_),
    .Y(_04260_));
 sg13g2_o21ai_1 _10029_ (.B1(net3163),
    .Y(_04261_),
    .A1(\core.f2e_inst[5] ),
    .A2(net3336));
 sg13g2_a21oi_2 _10030_ (.B1(_04261_),
    .Y(_04262_),
    .A2(_04260_),
    .A1(_04259_));
 sg13g2_o21ai_1 _10031_ (.B1(_04257_),
    .Y(_04263_),
    .A1(net882),
    .A2(_04170_));
 sg13g2_nor4_1 _10032_ (.A(net2748),
    .B(_04256_),
    .C(_04262_),
    .D(_04263_),
    .Y(_04264_));
 sg13g2_a21oi_1 _10033_ (.A1(_00595_),
    .A2(net2748),
    .Y(_00497_),
    .B1(_04264_));
 sg13g2_xnor2_1 _10034_ (.Y(_04265_),
    .A(_01216_),
    .B(_01217_));
 sg13g2_nor3_2 _10035_ (.A(net3552),
    .B(net3555),
    .C(_04023_),
    .Y(_04266_));
 sg13g2_nand2_1 _10036_ (.Y(_04267_),
    .A(net3546),
    .B(_04266_));
 sg13g2_nor2_1 _10037_ (.A(\core.work.alu.sval2[6] ),
    .B(net2965),
    .Y(_04268_));
 sg13g2_a21oi_1 _10038_ (.A1(net2965),
    .A2(_04267_),
    .Y(_04269_),
    .B1(_04268_));
 sg13g2_xnor2_1 _10039_ (.Y(_04270_),
    .A(_00020_),
    .B(_04269_));
 sg13g2_nand2_1 _10040_ (.Y(_04271_),
    .A(_04107_),
    .B(_04189_));
 sg13g2_nor2_1 _10041_ (.A(net2835),
    .B(_04271_),
    .Y(_04272_));
 sg13g2_nor2_1 _10042_ (.A(net2832),
    .B(_04191_),
    .Y(_04273_));
 sg13g2_nand2_1 _10043_ (.Y(_04274_),
    .A(_00108_),
    .B(net3063));
 sg13g2_nand2_1 _10044_ (.Y(_04275_),
    .A(_00106_),
    .B(net3057));
 sg13g2_nand2_1 _10045_ (.Y(_04276_),
    .A(_04274_),
    .B(_04275_));
 sg13g2_nor2_1 _10046_ (.A(net2824),
    .B(_04193_),
    .Y(_04277_));
 sg13g2_a22oi_1 _10047_ (.Y(_04278_),
    .B1(net2940),
    .B2(_04267_),
    .A2(net2955),
    .A1(_00717_));
 sg13g2_or2_1 _10048_ (.X(_04279_),
    .B(_04278_),
    .A(_00020_));
 sg13g2_nor2_1 _10049_ (.A(net2929),
    .B(_04267_),
    .Y(_04280_));
 sg13g2_a21oi_1 _10050_ (.A1(\core.work.alu.sval2[6] ),
    .A2(net2929),
    .Y(_04281_),
    .B1(_04280_));
 sg13g2_a22oi_1 _10051_ (.Y(_04282_),
    .B1(_04281_),
    .B2(_00020_),
    .A2(_04279_),
    .A1(net2947));
 sg13g2_nor2_1 _10052_ (.A(net2795),
    .B(_04277_),
    .Y(_04283_));
 sg13g2_nor3_1 _10053_ (.A(_04272_),
    .B(_04273_),
    .C(_04282_),
    .Y(_04284_));
 sg13g2_o21ai_1 _10054_ (.B1(_04283_),
    .Y(_04285_),
    .A1(net2827),
    .A2(_04276_));
 sg13g2_a221oi_1 _10055_ (.B2(net2858),
    .C1(_04285_),
    .B1(_04270_),
    .A1(net2927),
    .Y(_04286_),
    .A2(_04265_));
 sg13g2_a221oi_1 _10056_ (.B2(_04198_),
    .C1(_01196_),
    .B1(_01197_),
    .A1(net3543),
    .Y(_04287_),
    .A2(net3493));
 sg13g2_nor3_1 _10057_ (.A(_01193_),
    .B(_01218_),
    .C(_04287_),
    .Y(_04288_));
 sg13g2_o21ai_1 _10058_ (.B1(_01218_),
    .Y(_04289_),
    .A1(_01193_),
    .A2(_04287_));
 sg13g2_nand2b_1 _10059_ (.Y(_04290_),
    .B(_04289_),
    .A_N(_04288_));
 sg13g2_a221oi_1 _10060_ (.B2(net2795),
    .C1(net3301),
    .B1(_04290_),
    .A1(_04284_),
    .Y(_04291_),
    .A2(_04286_));
 sg13g2_or2_1 _10061_ (.X(_04292_),
    .B(_03364_),
    .A(_02134_));
 sg13g2_nand2_1 _10062_ (.Y(_04293_),
    .A(_04131_),
    .B(_04207_));
 sg13g2_nor3_1 _10063_ (.A(net3347),
    .B(_04140_),
    .C(_04293_),
    .Y(_04294_));
 sg13g2_o21ai_1 _10064_ (.B1(net3163),
    .Y(_04295_),
    .A1(net3510),
    .A2(net3338));
 sg13g2_nor2_2 _10065_ (.A(_04294_),
    .B(_04295_),
    .Y(_04296_));
 sg13g2_o21ai_1 _10066_ (.B1(_04292_),
    .Y(_04297_),
    .A1(net855),
    .A2(_04170_));
 sg13g2_nor4_1 _10067_ (.A(net2748),
    .B(_04291_),
    .C(_04296_),
    .D(_04297_),
    .Y(_04298_));
 sg13g2_a21oi_1 _10068_ (.A1(_00594_),
    .A2(net2748),
    .Y(_00498_),
    .B1(_04298_));
 sg13g2_nor3_1 _10069_ (.A(_01190_),
    .B(_01191_),
    .C(_01219_),
    .Y(_04299_));
 sg13g2_nand2_1 _10070_ (.Y(_04300_),
    .A(_01221_),
    .B(net2927));
 sg13g2_nor2_1 _10071_ (.A(_04299_),
    .B(_04300_),
    .Y(_04301_));
 sg13g2_nor3_2 _10072_ (.A(net3552),
    .B(net3555),
    .C(_03181_),
    .Y(_04302_));
 sg13g2_nand2_1 _10073_ (.Y(_04303_),
    .A(net3546),
    .B(_04302_));
 sg13g2_nand2_1 _10074_ (.Y(_04304_),
    .A(net2965),
    .B(_04303_));
 sg13g2_o21ai_1 _10075_ (.B1(_04304_),
    .Y(_04305_),
    .A1(\core.work.alu.sval2[7] ),
    .A2(net2965));
 sg13g2_o21ai_1 _10076_ (.B1(net2857),
    .Y(_04306_),
    .A1(_00154_),
    .A2(_04305_));
 sg13g2_a21oi_1 _10077_ (.A1(_00154_),
    .A2(_04305_),
    .Y(_04307_),
    .B1(_04306_));
 sg13g2_nand2_1 _10078_ (.Y(_04308_),
    .A(_00110_),
    .B(net3063));
 sg13g2_nand2_1 _10079_ (.Y(_04309_),
    .A(_00108_),
    .B(net3057));
 sg13g2_nand3_1 _10080_ (.B(_04308_),
    .C(_04309_),
    .A(_04015_),
    .Y(_04310_));
 sg13g2_o21ai_1 _10081_ (.B1(_04310_),
    .Y(_04311_),
    .A1(net2832),
    .A2(_04248_));
 sg13g2_nand3_1 _10082_ (.B(_04147_),
    .C(_04246_),
    .A(_03990_),
    .Y(_04312_));
 sg13g2_o21ai_1 _10083_ (.B1(_04312_),
    .Y(_04313_),
    .A1(net2824),
    .A2(_04250_));
 sg13g2_a22oi_1 _10084_ (.Y(_04314_),
    .B1(net2940),
    .B2(_04303_),
    .A2(net2954),
    .A1(_00718_));
 sg13g2_o21ai_1 _10085_ (.B1(_00154_),
    .Y(_04315_),
    .A1(net2929),
    .A2(_04303_));
 sg13g2_a21o_1 _10086_ (.A2(net2929),
    .A1(\core.work.alu.sval2[7] ),
    .B1(_04315_),
    .X(_04316_));
 sg13g2_a21oi_1 _10087_ (.A1(net2951),
    .A2(_04316_),
    .Y(_04317_),
    .B1(_04311_));
 sg13g2_o21ai_1 _10088_ (.B1(net2790),
    .Y(_04318_),
    .A1(_00154_),
    .A2(_04314_));
 sg13g2_nor4_1 _10089_ (.A(_04301_),
    .B(_04307_),
    .C(_04313_),
    .D(_04318_),
    .Y(_04319_));
 sg13g2_a21oi_1 _10090_ (.A1(\core.work.alu.sval2[6] ),
    .A2(\core.e2m_addr[6] ),
    .Y(_04320_),
    .B1(_04288_));
 sg13g2_xnor2_1 _10091_ (.Y(_04321_),
    .A(_01190_),
    .B(_04320_));
 sg13g2_a221oi_1 _10092_ (.B2(net2796),
    .C1(net3301),
    .B1(_04321_),
    .A1(_04317_),
    .Y(_04322_),
    .A2(_04319_));
 sg13g2_nand2_1 _10093_ (.Y(_04323_),
    .A(net3336),
    .B(_04218_));
 sg13g2_a21oi_2 _10094_ (.B1(_04209_),
    .Y(_04324_),
    .A2(_04220_),
    .A1(_04131_));
 sg13g2_a21oi_1 _10095_ (.A1(\core.f2e_inst[12] ),
    .A2(_04206_),
    .Y(_04325_),
    .B1(_04129_));
 sg13g2_o21ai_1 _10096_ (.B1(_04325_),
    .Y(_04326_),
    .A1(net3506),
    .A2(_04138_));
 sg13g2_and2_1 _10097_ (.A(net2852),
    .B(_04205_),
    .X(_04327_));
 sg13g2_a21oi_1 _10098_ (.A1(_04222_),
    .A2(_04327_),
    .Y(_04328_),
    .B1(_00155_));
 sg13g2_nor2_1 _10099_ (.A(_04326_),
    .B(_04328_),
    .Y(_04329_));
 sg13g2_o21ai_1 _10100_ (.B1(_04329_),
    .Y(_04330_),
    .A1(_00680_),
    .A2(_04324_));
 sg13g2_a22oi_1 _10101_ (.Y(_04331_),
    .B1(_04330_),
    .B2(net3337),
    .A2(_04323_),
    .A1(\core.f2e_inst[7] ));
 sg13g2_nor2_2 _10102_ (.A(net3160),
    .B(_04331_),
    .Y(_04332_));
 sg13g2_nand2_1 _10103_ (.Y(_04333_),
    .A(net2843),
    .B(_03384_));
 sg13g2_nor2_1 _10104_ (.A(net803),
    .B(_04170_),
    .Y(_04334_));
 sg13g2_nor4_1 _10105_ (.A(net2748),
    .B(_04322_),
    .C(_04332_),
    .D(_04334_),
    .Y(_04335_));
 sg13g2_a22oi_1 _10106_ (.Y(_00499_),
    .B1(_04333_),
    .B2(_04335_),
    .A2(net2748),
    .A1(_00593_));
 sg13g2_nand3_1 _10107_ (.B(net3296),
    .C(net3289),
    .A(net3544),
    .Y(_04336_));
 sg13g2_nand2_1 _10108_ (.Y(_04337_),
    .A(net2960),
    .B(_04336_));
 sg13g2_o21ai_1 _10109_ (.B1(_04337_),
    .Y(_04338_),
    .A1(\core.work.alu.sval2[8] ),
    .A2(net2960));
 sg13g2_xnor2_1 _10110_ (.Y(_04339_),
    .A(_00106_),
    .B(_04338_));
 sg13g2_nand2_1 _10111_ (.Y(_04340_),
    .A(_00111_),
    .B(net3063));
 sg13g2_nand2_1 _10112_ (.Y(_04341_),
    .A(_00110_),
    .B(net3057));
 sg13g2_nand2_1 _10113_ (.Y(_04342_),
    .A(_04340_),
    .B(_04341_));
 sg13g2_nor2_1 _10114_ (.A(net2828),
    .B(_04342_),
    .Y(_04343_));
 sg13g2_nor2_1 _10115_ (.A(net2829),
    .B(_04276_),
    .Y(_04344_));
 sg13g2_nor2_1 _10116_ (.A(net2824),
    .B(_04271_),
    .Y(_04345_));
 sg13g2_nand2_1 _10117_ (.Y(_04346_),
    .A(_04190_),
    .B(_04275_));
 sg13g2_nor2_1 _10118_ (.A(net2834),
    .B(_04346_),
    .Y(_04347_));
 sg13g2_a22oi_1 _10119_ (.Y(_04348_),
    .B1(net2938),
    .B2(_04336_),
    .A2(net2954),
    .A1(_00719_));
 sg13g2_nor2_1 _10120_ (.A(net2928),
    .B(_04336_),
    .Y(_04349_));
 sg13g2_a21oi_1 _10121_ (.A1(\core.work.alu.sval2[8] ),
    .A2(net2928),
    .Y(_04350_),
    .B1(_04349_));
 sg13g2_a21oi_1 _10122_ (.A1(_00106_),
    .A2(_04350_),
    .Y(_04351_),
    .B1(net2944));
 sg13g2_o21ai_1 _10123_ (.B1(net2789),
    .Y(_04352_),
    .A1(_00106_),
    .A2(_04348_));
 sg13g2_nor3_1 _10124_ (.A(_04345_),
    .B(_04347_),
    .C(_04352_),
    .Y(_04353_));
 sg13g2_o21ai_1 _10125_ (.B1(_04353_),
    .Y(_04354_),
    .A1(net2860),
    .A2(_04339_));
 sg13g2_nor4_1 _10126_ (.A(_04343_),
    .B(_04344_),
    .C(_04351_),
    .D(_04354_),
    .Y(_04355_));
 sg13g2_nand2b_1 _10127_ (.Y(_04356_),
    .B(_01222_),
    .A_N(_01176_));
 sg13g2_nand2_1 _10128_ (.Y(_04357_),
    .A(_01176_),
    .B(_01223_));
 sg13g2_nand3_1 _10129_ (.B(_04356_),
    .C(_04357_),
    .A(net2926),
    .Y(_04358_));
 sg13g2_nand2_1 _10130_ (.Y(_04359_),
    .A(\core.e2m_addr[7] ),
    .B(\core.work.alu.sval2[7] ));
 sg13g2_o21ai_1 _10131_ (.B1(_04359_),
    .Y(_04360_),
    .A1(_01190_),
    .A2(_04320_));
 sg13g2_nand2b_1 _10132_ (.Y(_04361_),
    .B(_04360_),
    .A_N(_01176_));
 sg13g2_xor2_1 _10133_ (.B(_04360_),
    .A(_01176_),
    .X(_04362_));
 sg13g2_a22oi_1 _10134_ (.Y(_04363_),
    .B1(_04362_),
    .B2(net2793),
    .A2(_04358_),
    .A1(_04355_));
 sg13g2_nand2_1 _10135_ (.Y(_04364_),
    .A(net3308),
    .B(_04363_));
 sg13g2_nor2_1 _10136_ (.A(net2889),
    .B(_03411_),
    .Y(_04365_));
 sg13g2_a21oi_1 _10137_ (.A1(_00115_),
    .A2(net2840),
    .Y(_04366_),
    .B1(_04365_));
 sg13g2_nand2_1 _10138_ (.Y(_04367_),
    .A(_04207_),
    .B(_04324_));
 sg13g2_nand3_1 _10139_ (.B(net3337),
    .C(_04367_),
    .A(\core.f2e_inst[3] ),
    .Y(_04368_));
 sg13g2_nand2b_1 _10140_ (.Y(_04369_),
    .B(_04225_),
    .A_N(_00156_));
 sg13g2_or2_2 _10141_ (.X(_04370_),
    .B(_04126_),
    .A(_04123_));
 sg13g2_o21ai_1 _10142_ (.B1(\core.f2e_inst[8] ),
    .Y(_04371_),
    .A1(_04226_),
    .A2(_04323_));
 sg13g2_nand4_1 _10143_ (.B(_04369_),
    .C(_04370_),
    .A(_04368_),
    .Y(_04372_),
    .D(_04371_));
 sg13g2_a221oi_1 _10144_ (.B2(net3164),
    .C1(net2747),
    .B1(_04372_),
    .A1(_04119_),
    .Y(_04373_),
    .A2(_04366_));
 sg13g2_a22oi_1 _10145_ (.Y(_00500_),
    .B1(_04364_),
    .B2(_04373_),
    .A2(net2751),
    .A1(_00603_));
 sg13g2_nand2b_1 _10146_ (.Y(_04374_),
    .B(_04357_),
    .A_N(_01229_));
 sg13g2_xnor2_1 _10147_ (.Y(_04375_),
    .A(_01174_),
    .B(_04374_));
 sg13g2_nand3_1 _10148_ (.B(net3296),
    .C(net3288),
    .A(net3544),
    .Y(_04376_));
 sg13g2_nand2_1 _10149_ (.Y(_04377_),
    .A(net2959),
    .B(_04376_));
 sg13g2_o21ai_1 _10150_ (.B1(_04377_),
    .Y(_04378_),
    .A1(\core.work.alu.sval2[9] ),
    .A2(net2959));
 sg13g2_o21ai_1 _10151_ (.B1(net2856),
    .Y(_04379_),
    .A1(_00108_),
    .A2(_04378_));
 sg13g2_a21oi_1 _10152_ (.A1(_00108_),
    .A2(_04378_),
    .Y(_04380_),
    .B1(_04379_));
 sg13g2_nand3_1 _10153_ (.B(_04308_),
    .C(_04309_),
    .A(_04010_),
    .Y(_04381_));
 sg13g2_nand2_1 _10154_ (.Y(_04382_),
    .A(_04247_),
    .B(_04309_));
 sg13g2_o21ai_1 _10155_ (.B1(_04381_),
    .Y(_04383_),
    .A1(net2834),
    .A2(_04382_));
 sg13g2_nand4_1 _10156_ (.B(net2853),
    .C(_04147_),
    .A(_01716_),
    .Y(_04384_),
    .D(_04246_));
 sg13g2_nand2_1 _10157_ (.Y(_04385_),
    .A(_00120_),
    .B(net3063));
 sg13g2_nand2_1 _10158_ (.Y(_04386_),
    .A(_00111_),
    .B(net3057));
 sg13g2_nand2_1 _10159_ (.Y(_04387_),
    .A(_04385_),
    .B(_04386_));
 sg13g2_o21ai_1 _10160_ (.B1(_04384_),
    .Y(_04388_),
    .A1(net2828),
    .A2(_04387_));
 sg13g2_a22oi_1 _10161_ (.Y(_04389_),
    .B1(net2938),
    .B2(_04376_),
    .A2(net2954),
    .A1(_00720_));
 sg13g2_nor2_1 _10162_ (.A(net2929),
    .B(_04376_),
    .Y(_04390_));
 sg13g2_a21oi_1 _10163_ (.A1(net3542),
    .A2(net2929),
    .Y(_04391_),
    .B1(_04390_));
 sg13g2_a21oi_1 _10164_ (.A1(_00108_),
    .A2(_04391_),
    .Y(_04392_),
    .B1(net2943));
 sg13g2_nor2_1 _10165_ (.A(net2793),
    .B(_04392_),
    .Y(_04393_));
 sg13g2_o21ai_1 _10166_ (.B1(_04393_),
    .Y(_04394_),
    .A1(_00108_),
    .A2(_04389_));
 sg13g2_nor4_1 _10167_ (.A(_04380_),
    .B(_04383_),
    .C(_04388_),
    .D(_04394_),
    .Y(_04395_));
 sg13g2_o21ai_1 _10168_ (.B1(_04395_),
    .Y(_04396_),
    .A1(net2924),
    .A2(_04375_));
 sg13g2_nand2_1 _10169_ (.Y(_04397_),
    .A(_01175_),
    .B(_04361_));
 sg13g2_a21oi_1 _10170_ (.A1(_01174_),
    .A2(_04397_),
    .Y(_04398_),
    .B1(net2789));
 sg13g2_o21ai_1 _10171_ (.B1(_04398_),
    .Y(_04399_),
    .A1(_01174_),
    .A2(_04397_));
 sg13g2_nand3_1 _10172_ (.B(_04396_),
    .C(_04399_),
    .A(net3308),
    .Y(_04400_));
 sg13g2_nor2_1 _10173_ (.A(net2889),
    .B(_03432_),
    .Y(_04401_));
 sg13g2_a21oi_1 _10174_ (.A1(_00116_),
    .A2(net2840),
    .Y(_04402_),
    .B1(_04401_));
 sg13g2_a21oi_1 _10175_ (.A1(_04119_),
    .A2(_04402_),
    .Y(_04403_),
    .B1(net3165));
 sg13g2_nand3_1 _10176_ (.B(net3336),
    .C(_04367_),
    .A(\core.f2e_inst[4] ),
    .Y(_04404_));
 sg13g2_nor3_1 _10177_ (.A(net3345),
    .B(_04219_),
    .C(_04226_),
    .Y(_04405_));
 sg13g2_nand2b_1 _10178_ (.Y(_04406_),
    .B(\core.f2e_inst[9] ),
    .A_N(_04405_));
 sg13g2_a21o_1 _10179_ (.A2(_04327_),
    .A1(_04223_),
    .B1(_00157_),
    .X(_04407_));
 sg13g2_a21oi_1 _10180_ (.A1(\core.f2e_inst[6] ),
    .A2(_04210_),
    .Y(_04408_),
    .B1(net3160));
 sg13g2_nand4_1 _10181_ (.B(_04406_),
    .C(_04407_),
    .A(_04404_),
    .Y(_04409_),
    .D(_04408_));
 sg13g2_a21oi_1 _10182_ (.A1(_04400_),
    .A2(_04403_),
    .Y(_04410_),
    .B1(net2747));
 sg13g2_a22oi_1 _10183_ (.Y(_04411_),
    .B1(_04409_),
    .B2(_04410_),
    .A2(net2747),
    .A1(net3488));
 sg13g2_inv_1 _10184_ (.Y(_00501_),
    .A(_04411_));
 sg13g2_a21oi_1 _10185_ (.A1(_01174_),
    .A2(_04374_),
    .Y(_04412_),
    .B1(_01231_));
 sg13g2_xnor2_1 _10186_ (.Y(_04413_),
    .A(_01167_),
    .B(_04412_));
 sg13g2_nor2_1 _10187_ (.A(\core.work.alu.sval2[10] ),
    .B(net2960),
    .Y(_04414_));
 sg13g2_nand3_1 _10188_ (.B(_01812_),
    .C(net3053),
    .A(net3544),
    .Y(_04415_));
 sg13g2_a21oi_1 _10189_ (.A1(net2960),
    .A2(_04415_),
    .Y(_04416_),
    .B1(_04414_));
 sg13g2_a21o_1 _10190_ (.A2(_04416_),
    .A1(_00714_),
    .B1(net2860),
    .X(_04417_));
 sg13g2_o21ai_1 _10191_ (.B1(net2944),
    .Y(_04418_),
    .A1(_00117_),
    .A2(net2953));
 sg13g2_a21oi_1 _10192_ (.A1(net2938),
    .A2(_04415_),
    .Y(_04419_),
    .B1(_04418_));
 sg13g2_a21oi_1 _10193_ (.A1(net2932),
    .A2(_04415_),
    .Y(_04420_),
    .B1(net2943));
 sg13g2_o21ai_1 _10194_ (.B1(_04420_),
    .Y(_04421_),
    .A1(\core.work.alu.sval2[10] ),
    .A2(net2932));
 sg13g2_a21oi_1 _10195_ (.A1(net2856),
    .A2(_04416_),
    .Y(_04422_),
    .B1(_00714_));
 sg13g2_a22oi_1 _10196_ (.Y(_04423_),
    .B1(_04421_),
    .B2(_04422_),
    .A2(_04419_),
    .A1(_04417_));
 sg13g2_or2_1 _10197_ (.X(_04424_),
    .B(_04346_),
    .A(net2822));
 sg13g2_nand2_1 _10198_ (.Y(_04425_),
    .A(_00120_),
    .B(net3057));
 sg13g2_nand2_1 _10199_ (.Y(_04426_),
    .A(_00122_),
    .B(net3061));
 sg13g2_nand2_1 _10200_ (.Y(_04427_),
    .A(_04425_),
    .B(_04426_));
 sg13g2_o21ai_1 _10201_ (.B1(_04424_),
    .Y(_04428_),
    .A1(net2828),
    .A2(_04427_));
 sg13g2_nand2_1 _10202_ (.Y(_04429_),
    .A(_04274_),
    .B(_04341_));
 sg13g2_nor2_1 _10203_ (.A(net2830),
    .B(_04342_),
    .Y(_04430_));
 sg13g2_o21ai_1 _10204_ (.B1(net2789),
    .Y(_04431_),
    .A1(net2834),
    .A2(_04429_));
 sg13g2_nor4_2 _10205_ (.A(_04423_),
    .B(_04428_),
    .C(_04430_),
    .Y(_04432_),
    .D(_04431_));
 sg13g2_o21ai_1 _10206_ (.B1(_04432_),
    .Y(_04433_),
    .A1(net2924),
    .A2(_04413_));
 sg13g2_o21ai_1 _10207_ (.B1(_01173_),
    .Y(_04434_),
    .A1(_01172_),
    .A2(_01175_));
 sg13g2_nor2_1 _10208_ (.A(_01174_),
    .B(_01176_),
    .Y(_04435_));
 sg13g2_a21oi_1 _10209_ (.A1(_04360_),
    .A2(_04435_),
    .Y(_04436_),
    .B1(_04434_));
 sg13g2_xnor2_1 _10210_ (.Y(_04437_),
    .A(_01168_),
    .B(_04436_));
 sg13g2_a21oi_1 _10211_ (.A1(net2793),
    .A2(_04437_),
    .Y(_04438_),
    .B1(net3298));
 sg13g2_nor2_1 _10212_ (.A(net2889),
    .B(_03456_),
    .Y(_04439_));
 sg13g2_a21oi_1 _10213_ (.A1(_00117_),
    .A2(net2840),
    .Y(_04440_),
    .B1(_04439_));
 sg13g2_a221oi_1 _10214_ (.B2(_04119_),
    .C1(net3165),
    .B1(_04440_),
    .A1(_04433_),
    .Y(_04441_),
    .A2(_04438_));
 sg13g2_a21oi_1 _10215_ (.A1(net2852),
    .A2(_04223_),
    .Y(_04442_),
    .B1(_00158_));
 sg13g2_a21oi_1 _10216_ (.A1(net3509),
    .A2(_04226_),
    .Y(_04443_),
    .B1(_04442_));
 sg13g2_nand3_1 _10217_ (.B(_04324_),
    .C(_04443_),
    .A(net2851),
    .Y(_04444_));
 sg13g2_or2_1 _10218_ (.X(_04445_),
    .B(_04216_),
    .A(_04210_));
 sg13g2_nor2_1 _10219_ (.A(\core.f2e_inst[15] ),
    .B(_04214_),
    .Y(_04446_));
 sg13g2_a21oi_1 _10220_ (.A1(\core.f2e_inst[15] ),
    .A2(_00151_),
    .Y(_04447_),
    .B1(_04214_));
 sg13g2_nor2_1 _10221_ (.A(_04445_),
    .B(_04447_),
    .Y(_04448_));
 sg13g2_nor2_1 _10222_ (.A(\core.f2e_inst[14] ),
    .B(_04218_),
    .Y(_04449_));
 sg13g2_nor3_1 _10223_ (.A(net3345),
    .B(_04206_),
    .C(_04449_),
    .Y(_04450_));
 sg13g2_o21ai_1 _10224_ (.B1(_04450_),
    .Y(_04451_),
    .A1(_00705_),
    .A2(_04448_));
 sg13g2_a221oi_1 _10225_ (.B2(net3509),
    .C1(net3160),
    .B1(_04451_),
    .A1(net3337),
    .Y(_04452_),
    .A2(_04444_));
 sg13g2_nor3_1 _10226_ (.A(net2747),
    .B(_04441_),
    .C(_04452_),
    .Y(_04453_));
 sg13g2_a21o_1 _10227_ (.A2(net2747),
    .A1(net3486),
    .B1(_04453_),
    .X(_00502_));
 sg13g2_o21ai_1 _10228_ (.B1(_01230_),
    .Y(_04454_),
    .A1(_01167_),
    .A2(_04412_));
 sg13g2_xnor2_1 _10229_ (.Y(_04455_),
    .A(_01171_),
    .B(_04454_));
 sg13g2_nand2_1 _10230_ (.Y(_04456_),
    .A(_00122_),
    .B(net3055));
 sg13g2_nand2_1 _10231_ (.Y(_04457_),
    .A(_00124_),
    .B(net3062));
 sg13g2_nand2_1 _10232_ (.Y(_04458_),
    .A(_04456_),
    .B(_04457_));
 sg13g2_nand2_1 _10233_ (.Y(_04459_),
    .A(_04308_),
    .B(_04386_));
 sg13g2_nor2_1 _10234_ (.A(net2834),
    .B(_04459_),
    .Y(_04460_));
 sg13g2_nor2_1 _10235_ (.A(net2830),
    .B(_04387_),
    .Y(_04461_));
 sg13g2_nand3_1 _10236_ (.B(net3296),
    .C(net3292),
    .A(net3544),
    .Y(_04462_));
 sg13g2_a22oi_1 _10237_ (.Y(_04463_),
    .B1(net2938),
    .B2(_04462_),
    .A2(net2954),
    .A1(_00721_));
 sg13g2_a21oi_1 _10238_ (.A1(net2932),
    .A2(_04462_),
    .Y(_04464_),
    .B1(net2943));
 sg13g2_o21ai_1 _10239_ (.B1(_04464_),
    .Y(_04465_),
    .A1(\core.work.alu.sval2[11] ),
    .A2(net2932));
 sg13g2_a22oi_1 _10240_ (.Y(_04466_),
    .B1(_04465_),
    .B2(_00111_),
    .A2(_04463_),
    .A1(net2943));
 sg13g2_nor2_1 _10241_ (.A(\core.work.alu.sval2[11] ),
    .B(net2959),
    .Y(_04467_));
 sg13g2_a21oi_1 _10242_ (.A1(net2959),
    .A2(_04462_),
    .Y(_04468_),
    .B1(_04467_));
 sg13g2_a21oi_1 _10243_ (.A1(_00715_),
    .A2(_04468_),
    .Y(_04469_),
    .B1(net2860));
 sg13g2_o21ai_1 _10244_ (.B1(_04469_),
    .Y(_04470_),
    .A1(_00715_),
    .A2(_04468_));
 sg13g2_nor2_1 _10245_ (.A(_04460_),
    .B(_04461_),
    .Y(_04471_));
 sg13g2_o21ai_1 _10246_ (.B1(_04471_),
    .Y(_04472_),
    .A1(net2822),
    .A2(_04382_));
 sg13g2_o21ai_1 _10247_ (.B1(_04470_),
    .Y(_04473_),
    .A1(net2825),
    .A2(_04458_));
 sg13g2_nor4_1 _10248_ (.A(net2793),
    .B(_04466_),
    .C(_04472_),
    .D(_04473_),
    .Y(_04474_));
 sg13g2_o21ai_1 _10249_ (.B1(_04474_),
    .Y(_04475_),
    .A1(net2924),
    .A2(_04455_));
 sg13g2_o21ai_1 _10250_ (.B1(_01166_),
    .Y(_04476_),
    .A1(_01168_),
    .A2(_04436_));
 sg13g2_a21oi_1 _10251_ (.A1(_01171_),
    .A2(_04476_),
    .Y(_04477_),
    .B1(net2789));
 sg13g2_o21ai_1 _10252_ (.B1(_04477_),
    .Y(_04478_),
    .A1(_01171_),
    .A2(_04476_));
 sg13g2_nand3_1 _10253_ (.B(_04475_),
    .C(_04478_),
    .A(net3305),
    .Y(_04479_));
 sg13g2_nor2_1 _10254_ (.A(net2889),
    .B(_03479_),
    .Y(_04480_));
 sg13g2_a21oi_1 _10255_ (.A1(_00118_),
    .A2(net2840),
    .Y(_04481_),
    .B1(_04480_));
 sg13g2_a21oi_1 _10256_ (.A1(_04119_),
    .A2(_04481_),
    .Y(_04482_),
    .B1(_01767_));
 sg13g2_o21ai_1 _10257_ (.B1(\core.f2e_inst[11] ),
    .Y(_04483_),
    .A1(_04226_),
    .A2(_04451_));
 sg13g2_a21oi_1 _10258_ (.A1(_04123_),
    .A2(_04223_),
    .Y(_04484_),
    .B1(_00152_));
 sg13g2_nor2_1 _10259_ (.A(net3160),
    .B(_04484_),
    .Y(_04485_));
 sg13g2_a221oi_1 _10260_ (.B2(_04485_),
    .C1(net2744),
    .B1(_04483_),
    .A1(_04479_),
    .Y(_04486_),
    .A2(_04482_));
 sg13g2_a21o_1 _10261_ (.A2(net2747),
    .A1(net876),
    .B1(_04486_),
    .X(_00503_));
 sg13g2_o21ai_1 _10262_ (.B1(_01170_),
    .Y(_04487_),
    .A1(_01166_),
    .A2(_01169_));
 sg13g2_nor2_1 _10263_ (.A(_01168_),
    .B(_01171_),
    .Y(_04488_));
 sg13g2_and2_1 _10264_ (.A(_04435_),
    .B(_04488_),
    .X(_04489_));
 sg13g2_a221oi_1 _10265_ (.B2(_04360_),
    .C1(_04487_),
    .B1(_04489_),
    .A1(_04434_),
    .Y(_04490_),
    .A2(_04488_));
 sg13g2_xor2_1 _10266_ (.B(_04490_),
    .A(_01187_),
    .X(_04491_));
 sg13g2_nor2_1 _10267_ (.A(net2789),
    .B(_04491_),
    .Y(_04492_));
 sg13g2_a21o_1 _10268_ (.A2(_01223_),
    .A1(_01177_),
    .B1(_01234_),
    .X(_04493_));
 sg13g2_nand2_1 _10269_ (.Y(_04494_),
    .A(_01187_),
    .B(_04493_));
 sg13g2_xnor2_1 _10270_ (.Y(_04495_),
    .A(_01187_),
    .B(_04493_));
 sg13g2_nor2_1 _10271_ (.A(\core.work.alu.sval2[12] ),
    .B(net2957),
    .Y(_04496_));
 sg13g2_nor4_2 _10272_ (.A(net3539),
    .B(net3562),
    .C(net3551),
    .Y(_04497_),
    .D(net3555));
 sg13g2_nand2_1 _10273_ (.Y(_04498_),
    .A(net3544),
    .B(_04497_));
 sg13g2_a21oi_1 _10274_ (.A1(net2957),
    .A2(_04498_),
    .Y(_04499_),
    .B1(_04496_));
 sg13g2_xnor2_1 _10275_ (.Y(_04500_),
    .A(_00120_),
    .B(_04499_));
 sg13g2_nor2_1 _10276_ (.A(net2830),
    .B(_04427_),
    .Y(_04501_));
 sg13g2_nand2_1 _10277_ (.Y(_04502_),
    .A(_00126_),
    .B(net3064));
 sg13g2_nand2_1 _10278_ (.Y(_04503_),
    .A(_00124_),
    .B(net3056));
 sg13g2_nand2_1 _10279_ (.Y(_04504_),
    .A(_04502_),
    .B(_04503_));
 sg13g2_nor2_1 _10280_ (.A(net2825),
    .B(_04504_),
    .Y(_04505_));
 sg13g2_a22oi_1 _10281_ (.Y(_04506_),
    .B1(net2938),
    .B2(_04498_),
    .A2(net2954),
    .A1(_00722_));
 sg13g2_a21oi_1 _10282_ (.A1(net2943),
    .A2(_04506_),
    .Y(_04507_),
    .B1(_00120_));
 sg13g2_nand2_1 _10283_ (.Y(_04508_),
    .A(_04340_),
    .B(_04425_));
 sg13g2_o21ai_1 _10284_ (.B1(net2950),
    .Y(_04509_),
    .A1(net3541),
    .A2(net2932));
 sg13g2_a21oi_1 _10285_ (.A1(net2931),
    .A2(_04498_),
    .Y(_04510_),
    .B1(_04509_));
 sg13g2_o21ai_1 _10286_ (.B1(net2789),
    .Y(_04511_),
    .A1(net2822),
    .A2(_04429_));
 sg13g2_nor2_1 _10287_ (.A(_04505_),
    .B(_04510_),
    .Y(_04512_));
 sg13g2_o21ai_1 _10288_ (.B1(_04512_),
    .Y(_04513_),
    .A1(net2833),
    .A2(_04508_));
 sg13g2_a21oi_1 _10289_ (.A1(net2855),
    .A2(_04500_),
    .Y(_04514_),
    .B1(_04513_));
 sg13g2_o21ai_1 _10290_ (.B1(_04514_),
    .Y(_04515_),
    .A1(net2924),
    .A2(_04495_));
 sg13g2_nor4_1 _10291_ (.A(_04501_),
    .B(_04507_),
    .C(_04511_),
    .D(_04515_),
    .Y(_04516_));
 sg13g2_nor3_2 _10292_ (.A(net3301),
    .B(_04492_),
    .C(_04516_),
    .Y(_04517_));
 sg13g2_o21ai_1 _10293_ (.B1(\core.f2e_inst[12] ),
    .Y(_04518_),
    .A1(_04129_),
    .A2(_04130_));
 sg13g2_nand2_2 _10294_ (.Y(_04519_),
    .A(net3336),
    .B(_04518_));
 sg13g2_nand2_1 _10295_ (.Y(_04520_),
    .A(net3511),
    .B(net3506));
 sg13g2_nand3_1 _10296_ (.B(net3510),
    .C(net3506),
    .A(net3511),
    .Y(_04521_));
 sg13g2_nand3_1 _10297_ (.B(\core.f2e_inst[11] ),
    .C(_04521_),
    .A(net3508),
    .Y(_04522_));
 sg13g2_nand2_1 _10298_ (.Y(_04523_),
    .A(net3504),
    .B(_04206_));
 sg13g2_a21oi_1 _10299_ (.A1(_04204_),
    .A2(_04522_),
    .Y(_04524_),
    .B1(_04227_));
 sg13g2_o21ai_1 _10300_ (.B1(_04523_),
    .Y(_04525_),
    .A1(_00159_),
    .A2(_04127_));
 sg13g2_nor2_1 _10301_ (.A(_04519_),
    .B(_04525_),
    .Y(_04526_));
 sg13g2_a221oi_1 _10302_ (.B2(_04526_),
    .C1(net3160),
    .B1(_04524_),
    .A1(_00701_),
    .Y(_04527_),
    .A2(net3346));
 sg13g2_o21ai_1 _10303_ (.B1(net2840),
    .Y(_04528_),
    .A1(net765),
    .A2(_04118_));
 sg13g2_o21ai_1 _10304_ (.B1(_04528_),
    .Y(_04529_),
    .A1(net2889),
    .A2(_03510_));
 sg13g2_nor3_1 _10305_ (.A(net2746),
    .B(_04517_),
    .C(_04527_),
    .Y(_04530_));
 sg13g2_a22oi_1 _10306_ (.Y(_00504_),
    .B1(_04529_),
    .B2(_04530_),
    .A2(net2746),
    .A1(_00601_));
 sg13g2_o21ai_1 _10307_ (.B1(_01186_),
    .Y(_04531_),
    .A1(_01187_),
    .A2(_04490_));
 sg13g2_xnor2_1 _10308_ (.Y(_04532_),
    .A(_01185_),
    .B(_04531_));
 sg13g2_nand3_1 _10309_ (.B(_01227_),
    .C(_04494_),
    .A(_01184_),
    .Y(_04533_));
 sg13g2_a21o_1 _10310_ (.A2(_04494_),
    .A1(_01227_),
    .B1(_01184_),
    .X(_04534_));
 sg13g2_and2_1 _10311_ (.A(_04533_),
    .B(_04534_),
    .X(_04535_));
 sg13g2_nand2_1 _10312_ (.Y(_04536_),
    .A(_00126_),
    .B(net3056));
 sg13g2_nand2_1 _10313_ (.Y(_04537_),
    .A(_00023_),
    .B(net3064));
 sg13g2_nand2_1 _10314_ (.Y(_04538_),
    .A(_04536_),
    .B(_04537_));
 sg13g2_nor2_1 _10315_ (.A(net2825),
    .B(_04538_),
    .Y(_04539_));
 sg13g2_nand2_1 _10316_ (.Y(_04540_),
    .A(_04385_),
    .B(_04456_));
 sg13g2_nor2_1 _10317_ (.A(net2833),
    .B(_04540_),
    .Y(_04541_));
 sg13g2_nor2_1 _10318_ (.A(net2829),
    .B(_04458_),
    .Y(_04542_));
 sg13g2_nor3_2 _10319_ (.A(net3551),
    .B(net3555),
    .C(_03985_),
    .Y(_04543_));
 sg13g2_nand2_1 _10320_ (.Y(_04544_),
    .A(net3544),
    .B(_04543_));
 sg13g2_o21ai_1 _10321_ (.B1(net2943),
    .Y(_04545_),
    .A1(_00121_),
    .A2(net2952));
 sg13g2_a21oi_1 _10322_ (.A1(net2941),
    .A2(_04544_),
    .Y(_04546_),
    .B1(_04545_));
 sg13g2_nor2_1 _10323_ (.A(net2822),
    .B(_04459_),
    .Y(_04547_));
 sg13g2_o21ai_1 _10324_ (.B1(net2950),
    .Y(_04548_),
    .A1(\core.work.alu.sval2[13] ),
    .A2(net2932));
 sg13g2_a21oi_1 _10325_ (.A1(net2932),
    .A2(_04544_),
    .Y(_04549_),
    .B1(_04548_));
 sg13g2_nor3_1 _10326_ (.A(net2793),
    .B(_04547_),
    .C(_04549_),
    .Y(_04550_));
 sg13g2_o21ai_1 _10327_ (.B1(_04550_),
    .Y(_04551_),
    .A1(_00122_),
    .A2(_04546_));
 sg13g2_nor4_1 _10328_ (.A(_04539_),
    .B(_04541_),
    .C(_04542_),
    .D(_04551_),
    .Y(_04552_));
 sg13g2_nor2_1 _10329_ (.A(\core.work.alu.sval2[13] ),
    .B(net2959),
    .Y(_04553_));
 sg13g2_a21oi_1 _10330_ (.A1(net2959),
    .A2(_04544_),
    .Y(_04554_),
    .B1(_04553_));
 sg13g2_xnor2_1 _10331_ (.Y(_04555_),
    .A(_00122_),
    .B(_04554_));
 sg13g2_a22oi_1 _10332_ (.Y(_04556_),
    .B1(_04555_),
    .B2(net2854),
    .A2(_04535_),
    .A1(net2926));
 sg13g2_a21oi_1 _10333_ (.A1(_04552_),
    .A2(_04556_),
    .Y(_04557_),
    .B1(net3301));
 sg13g2_o21ai_1 _10334_ (.B1(_04557_),
    .Y(_04558_),
    .A1(net2788),
    .A2(_04532_));
 sg13g2_nor2_1 _10335_ (.A(net2889),
    .B(_03532_),
    .Y(_04559_));
 sg13g2_a21oi_1 _10336_ (.A1(_00121_),
    .A2(net2840),
    .Y(_04560_),
    .B1(_04559_));
 sg13g2_a21oi_1 _10337_ (.A1(_04119_),
    .A2(_04560_),
    .Y(_04561_),
    .B1(net3164));
 sg13g2_nand3b_1 _10338_ (.B(net3510),
    .C(_00701_),
    .Y(_04562_),
    .A_N(net3511));
 sg13g2_nand3_1 _10339_ (.B(_04521_),
    .C(_04562_),
    .A(net3508),
    .Y(_04563_));
 sg13g2_nand2_1 _10340_ (.Y(_04564_),
    .A(_04258_),
    .B(_04563_));
 sg13g2_o21ai_1 _10341_ (.B1(_04564_),
    .Y(_04565_),
    .A1(_00160_),
    .A2(net2852));
 sg13g2_inv_1 _10342_ (.Y(_04566_),
    .A(_04565_));
 sg13g2_nand4_1 _10343_ (.B(_04214_),
    .C(_04518_),
    .A(_04211_),
    .Y(_04567_),
    .D(_04566_));
 sg13g2_a22oi_1 _10344_ (.Y(_04568_),
    .B1(_04221_),
    .B2(_04567_),
    .A2(net3346),
    .A1(net3504));
 sg13g2_a221oi_1 _10345_ (.B2(net3164),
    .C1(net2743),
    .B1(_04568_),
    .A1(_04558_),
    .Y(_04569_),
    .A2(_04561_));
 sg13g2_a21o_1 _10346_ (.A2(net2743),
    .A1(net3482),
    .B1(_04569_),
    .X(_00505_));
 sg13g2_o21ai_1 _10347_ (.B1(_01183_),
    .Y(_04570_),
    .A1(_01182_),
    .A2(_01186_));
 sg13g2_nor2_1 _10348_ (.A(_01185_),
    .B(_01187_),
    .Y(_04571_));
 sg13g2_nand2b_1 _10349_ (.Y(_04572_),
    .B(_04571_),
    .A_N(_04490_));
 sg13g2_nand2b_1 _10350_ (.Y(_04573_),
    .B(_04572_),
    .A_N(_04570_));
 sg13g2_nand2_1 _10351_ (.Y(_04574_),
    .A(_01180_),
    .B(_04573_));
 sg13g2_xnor2_1 _10352_ (.Y(_04575_),
    .A(_01180_),
    .B(_04573_));
 sg13g2_nor2_1 _10353_ (.A(\core.work.alu.sval2[14] ),
    .B(net2958),
    .Y(_04576_));
 sg13g2_nor3_2 _10354_ (.A(net3551),
    .B(net3555),
    .C(_04023_),
    .Y(_04577_));
 sg13g2_nand2_1 _10355_ (.Y(_04578_),
    .A(net3544),
    .B(_04577_));
 sg13g2_a21oi_1 _10356_ (.A1(net2958),
    .A2(_04578_),
    .Y(_04579_),
    .B1(_04576_));
 sg13g2_xnor2_1 _10357_ (.Y(_04580_),
    .A(_00124_),
    .B(_04579_));
 sg13g2_a22oi_1 _10358_ (.Y(_04581_),
    .B1(net2938),
    .B2(_04578_),
    .A2(net2954),
    .A1(_00723_));
 sg13g2_nand2_1 _10359_ (.Y(_04582_),
    .A(_00025_),
    .B(net3064));
 sg13g2_nand2_1 _10360_ (.Y(_04583_),
    .A(_00023_),
    .B(net3060));
 sg13g2_nand2_1 _10361_ (.Y(_04584_),
    .A(_04582_),
    .B(_04583_));
 sg13g2_nor2_1 _10362_ (.A(net2826),
    .B(_04584_),
    .Y(_04585_));
 sg13g2_nand2_1 _10363_ (.Y(_04586_),
    .A(_04426_),
    .B(_04503_));
 sg13g2_nor2_1 _10364_ (.A(net2834),
    .B(_04586_),
    .Y(_04587_));
 sg13g2_a21oi_1 _10365_ (.A1(net2942),
    .A2(_04581_),
    .Y(_04588_),
    .B1(_00124_));
 sg13g2_o21ai_1 _10366_ (.B1(net2949),
    .Y(_04589_),
    .A1(\core.work.alu.sval2[14] ),
    .A2(net2931));
 sg13g2_a21oi_1 _10367_ (.A1(net2931),
    .A2(_04578_),
    .Y(_04590_),
    .B1(_04589_));
 sg13g2_nand2_1 _10368_ (.Y(_04591_),
    .A(_01226_),
    .B(_04534_));
 sg13g2_nand2b_1 _10369_ (.Y(_04592_),
    .B(_04591_),
    .A_N(_01180_));
 sg13g2_o21ai_1 _10370_ (.B1(net2788),
    .Y(_04593_),
    .A1(net2829),
    .A2(_04504_));
 sg13g2_nor3_1 _10371_ (.A(_04587_),
    .B(_04588_),
    .C(_04593_),
    .Y(_04594_));
 sg13g2_nor2_1 _10372_ (.A(_04585_),
    .B(_04590_),
    .Y(_04595_));
 sg13g2_o21ai_1 _10373_ (.B1(_04595_),
    .Y(_04596_),
    .A1(net2821),
    .A2(_04508_));
 sg13g2_xnor2_1 _10374_ (.Y(_04597_),
    .A(_01180_),
    .B(_04591_));
 sg13g2_a221oi_1 _10375_ (.B2(net2925),
    .C1(_04596_),
    .B1(_04597_),
    .A1(net2854),
    .Y(_04598_),
    .A2(_04580_));
 sg13g2_a22oi_1 _10376_ (.Y(_04599_),
    .B1(_04594_),
    .B2(_04598_),
    .A2(_04575_),
    .A1(net2793));
 sg13g2_o21ai_1 _10377_ (.B1(net2840),
    .Y(_04600_),
    .A1(net850),
    .A2(_04118_));
 sg13g2_o21ai_1 _10378_ (.B1(_04600_),
    .Y(_04601_),
    .A1(net2889),
    .A2(_03556_));
 sg13g2_and4_1 _10379_ (.A(net3508),
    .B(\core.f2e_inst[11] ),
    .C(_04520_),
    .D(_04562_),
    .X(_04602_));
 sg13g2_nor2_1 _10380_ (.A(net2851),
    .B(_04602_),
    .Y(_04603_));
 sg13g2_nor2_1 _10381_ (.A(_00161_),
    .B(net2852),
    .Y(_04604_));
 sg13g2_nor3_1 _10382_ (.A(_04519_),
    .B(_04603_),
    .C(_04604_),
    .Y(_04605_));
 sg13g2_a21oi_1 _10383_ (.A1(_00705_),
    .A2(net3345),
    .Y(_04606_),
    .B1(_04605_));
 sg13g2_a221oi_1 _10384_ (.B2(net3164),
    .C1(net2743),
    .B1(_04606_),
    .A1(net3303),
    .Y(_04607_),
    .A2(_04599_));
 sg13g2_a22oi_1 _10385_ (.Y(_00506_),
    .B1(_04601_),
    .B2(_04607_),
    .A2(net2743),
    .A1(_00600_));
 sg13g2_nand2_1 _10386_ (.Y(_04608_),
    .A(\core.work.alu.sval2[14] ),
    .B(net3481));
 sg13g2_nand2_1 _10387_ (.Y(_04609_),
    .A(_04574_),
    .B(_04608_));
 sg13g2_xnor2_1 _10388_ (.Y(_04610_),
    .A(_01178_),
    .B(_04609_));
 sg13g2_nand2_1 _10389_ (.Y(_04611_),
    .A(_01179_),
    .B(_04592_));
 sg13g2_xor2_1 _10390_ (.B(_04611_),
    .A(_01178_),
    .X(_04612_));
 sg13g2_nand2_1 _10391_ (.Y(_04613_),
    .A(_04457_),
    .B(_04536_));
 sg13g2_nor2_1 _10392_ (.A(net2835),
    .B(_04613_),
    .Y(_04614_));
 sg13g2_or2_1 _10393_ (.X(_04615_),
    .B(_04538_),
    .A(net2831));
 sg13g2_o21ai_1 _10394_ (.B1(_04615_),
    .Y(_04616_),
    .A1(net2823),
    .A2(_04540_));
 sg13g2_nor3_2 _10395_ (.A(net3551),
    .B(net3555),
    .C(_03181_),
    .Y(_04617_));
 sg13g2_nand2_1 _10396_ (.Y(_04618_),
    .A(net3545),
    .B(_04617_));
 sg13g2_o21ai_1 _10397_ (.B1(net2946),
    .Y(_04619_),
    .A1(_00125_),
    .A2(_03978_));
 sg13g2_a21oi_1 _10398_ (.A1(net2939),
    .A2(_04618_),
    .Y(_04620_),
    .B1(_04619_));
 sg13g2_nor2_1 _10399_ (.A(_00126_),
    .B(_04620_),
    .Y(_04621_));
 sg13g2_nand2_1 _10400_ (.Y(_04622_),
    .A(_00028_),
    .B(net3064));
 sg13g2_nand2_1 _10401_ (.Y(_04623_),
    .A(_00025_),
    .B(net3060));
 sg13g2_nand2_1 _10402_ (.Y(_04624_),
    .A(_04622_),
    .B(_04623_));
 sg13g2_o21ai_1 _10403_ (.B1(net2951),
    .Y(_04625_),
    .A1(\core.work.alu.sval2[15] ),
    .A2(net2934));
 sg13g2_a21o_1 _10404_ (.A2(_04618_),
    .A1(net2934),
    .B1(_04625_),
    .X(_04626_));
 sg13g2_o21ai_1 _10405_ (.B1(_04626_),
    .Y(_04627_),
    .A1(net2826),
    .A2(_04624_));
 sg13g2_nor4_1 _10406_ (.A(_04614_),
    .B(_04616_),
    .C(_04621_),
    .D(_04627_),
    .Y(_04628_));
 sg13g2_nand2_1 _10407_ (.Y(_04629_),
    .A(net2963),
    .B(_04618_));
 sg13g2_o21ai_1 _10408_ (.B1(_04629_),
    .Y(_04630_),
    .A1(\core.work.alu.sval2[15] ),
    .A2(net2963));
 sg13g2_xnor2_1 _10409_ (.Y(_04631_),
    .A(_00126_),
    .B(_04630_));
 sg13g2_o21ai_1 _10410_ (.B1(_04628_),
    .Y(_04632_),
    .A1(net2859),
    .A2(_04631_));
 sg13g2_a221oi_1 _10411_ (.B2(net2927),
    .C1(_04632_),
    .B1(_04612_),
    .A1(net2794),
    .Y(_04633_),
    .A2(_04610_));
 sg13g2_nand2b_1 _10412_ (.Y(_04634_),
    .B(net3309),
    .A_N(_04633_));
 sg13g2_a21oi_1 _10413_ (.A1(net3507),
    .A2(_04137_),
    .Y(_04635_),
    .B1(_04449_));
 sg13g2_inv_1 _10414_ (.Y(_04636_),
    .A(_04635_));
 sg13g2_nand2_1 _10415_ (.Y(_04637_),
    .A(_04212_),
    .B(_04635_));
 sg13g2_nand2_1 _10416_ (.Y(_04638_),
    .A(\core.f2e_inst[7] ),
    .B(_04637_));
 sg13g2_a21oi_1 _10417_ (.A1(_04139_),
    .A2(_04205_),
    .Y(_04639_),
    .B1(_00155_));
 sg13g2_nor2_1 _10418_ (.A(_00162_),
    .B(net2852),
    .Y(_04640_));
 sg13g2_nor3_1 _10419_ (.A(_04519_),
    .B(_04639_),
    .C(_04640_),
    .Y(_04641_));
 sg13g2_a22oi_1 _10420_ (.Y(_04642_),
    .B1(_04638_),
    .B2(_04641_),
    .A2(net3345),
    .A1(_00708_));
 sg13g2_nor2_1 _10421_ (.A(net2889),
    .B(_03582_),
    .Y(_04643_));
 sg13g2_a21oi_1 _10422_ (.A1(_00125_),
    .A2(net2840),
    .Y(_04644_),
    .B1(_04643_));
 sg13g2_a221oi_1 _10423_ (.B2(_04119_),
    .C1(net2745),
    .B1(_04644_),
    .A1(net3164),
    .Y(_04645_),
    .A2(_04642_));
 sg13g2_a22oi_1 _10424_ (.Y(_00507_),
    .B1(_04634_),
    .B2(_04645_),
    .A2(net2750),
    .A1(_00599_));
 sg13g2_nand2_1 _10425_ (.Y(_04646_),
    .A(net3472),
    .B(net2745));
 sg13g2_nor2b_1 _10426_ (.A(_01178_),
    .B_N(_01180_),
    .Y(_04647_));
 sg13g2_nand2_1 _10427_ (.Y(_04648_),
    .A(_04571_),
    .B(_04647_));
 sg13g2_a21oi_1 _10428_ (.A1(_00598_),
    .A2(_00599_),
    .Y(_04649_),
    .B1(_04608_));
 sg13g2_a221oi_1 _10429_ (.B2(_04647_),
    .C1(_04649_),
    .B1(_04570_),
    .A1(\core.work.alu.sval2[15] ),
    .Y(_04650_),
    .A2(net3478));
 sg13g2_o21ai_1 _10430_ (.B1(_04650_),
    .Y(_04651_),
    .A1(_04490_),
    .A2(_04648_));
 sg13g2_nand2_1 _10431_ (.Y(_04652_),
    .A(_01163_),
    .B(_04651_));
 sg13g2_xnor2_1 _10432_ (.Y(_04653_),
    .A(_01163_),
    .B(_04651_));
 sg13g2_xor2_1 _10433_ (.B(_01240_),
    .A(_01163_),
    .X(_04654_));
 sg13g2_nand3_1 _10434_ (.B(net3295),
    .C(net3290),
    .A(net3548),
    .Y(_04655_));
 sg13g2_nand2_1 _10435_ (.Y(_04656_),
    .A(net2962),
    .B(_04655_));
 sg13g2_o21ai_1 _10436_ (.B1(_04656_),
    .Y(_04657_),
    .A1(net3535),
    .A2(net2962));
 sg13g2_o21ai_1 _10437_ (.B1(net2857),
    .Y(_04658_),
    .A1(_00023_),
    .A2(_04657_));
 sg13g2_a22oi_1 _10438_ (.Y(_04659_),
    .B1(net2939),
    .B2(_04655_),
    .A2(net2955),
    .A1(_00635_));
 sg13g2_nand3_1 _10439_ (.B(_04658_),
    .C(_04659_),
    .A(net2946),
    .Y(_04660_));
 sg13g2_a21oi_1 _10440_ (.A1(net2933),
    .A2(_04655_),
    .Y(_04661_),
    .B1(net2945));
 sg13g2_o21ai_1 _10441_ (.B1(_04661_),
    .Y(_04662_),
    .A1(net3535),
    .A2(net2933));
 sg13g2_and2_1 _10442_ (.A(_00023_),
    .B(_04662_),
    .X(_04663_));
 sg13g2_o21ai_1 _10443_ (.B1(_04663_),
    .Y(_04664_),
    .A1(net2859),
    .A2(_04657_));
 sg13g2_nand2_1 _10444_ (.Y(_04665_),
    .A(_04502_),
    .B(_04583_));
 sg13g2_nor2_1 _10445_ (.A(net2835),
    .B(_04665_),
    .Y(_04666_));
 sg13g2_or2_1 _10446_ (.X(_04667_),
    .B(_04584_),
    .A(net2831));
 sg13g2_nand2_1 _10447_ (.Y(_04668_),
    .A(_00030_),
    .B(net3064));
 sg13g2_nand2_1 _10448_ (.Y(_04669_),
    .A(_00028_),
    .B(net3060));
 sg13g2_nand2_1 _10449_ (.Y(_04670_),
    .A(_04668_),
    .B(_04669_));
 sg13g2_o21ai_1 _10450_ (.B1(net2790),
    .Y(_04671_),
    .A1(net2826),
    .A2(_04670_));
 sg13g2_o21ai_1 _10451_ (.B1(_04667_),
    .Y(_04672_),
    .A1(net2823),
    .A2(_04586_));
 sg13g2_a21oi_1 _10452_ (.A1(_04660_),
    .A2(_04664_),
    .Y(_04673_),
    .B1(_04672_));
 sg13g2_o21ai_1 _10453_ (.B1(_04673_),
    .Y(_04674_),
    .A1(_04012_),
    .A2(_04654_));
 sg13g2_nor3_1 _10454_ (.A(_04666_),
    .B(_04671_),
    .C(_04674_),
    .Y(_04675_));
 sg13g2_a21oi_2 _10455_ (.B1(_04675_),
    .Y(_04676_),
    .A2(_04653_),
    .A1(net2797));
 sg13g2_a221oi_1 _10456_ (.B2(net3303),
    .C1(net3165),
    .B1(_04676_),
    .A1(net2842),
    .Y(_04677_),
    .A2(_03609_));
 sg13g2_a21oi_1 _10457_ (.A1(_00150_),
    .A2(_04126_),
    .Y(_04678_),
    .B1(_04123_));
 sg13g2_nor3_1 _10458_ (.A(_04447_),
    .B(_04519_),
    .C(_04678_),
    .Y(_04679_));
 sg13g2_a21oi_1 _10459_ (.A1(_04139_),
    .A2(net2851),
    .Y(_04680_),
    .B1(_00156_));
 sg13g2_a21oi_1 _10460_ (.A1(\core.f2e_inst[8] ),
    .A2(_04637_),
    .Y(_04681_),
    .B1(_04680_));
 sg13g2_nand3_1 _10461_ (.B(_04679_),
    .C(_04681_),
    .A(_04221_),
    .Y(_04682_));
 sg13g2_o21ai_1 _10462_ (.B1(_04682_),
    .Y(_04683_),
    .A1(\core.f2e_inst[16] ),
    .A2(net3336));
 sg13g2_a21o_1 _10463_ (.A2(_04683_),
    .A1(net3162),
    .B1(net2742),
    .X(_04684_));
 sg13g2_o21ai_1 _10464_ (.B1(_04646_),
    .Y(_00508_),
    .A1(_04677_),
    .A2(_04684_));
 sg13g2_nand2_1 _10465_ (.Y(_04685_),
    .A(_01162_),
    .B(_04652_));
 sg13g2_xnor2_1 _10466_ (.Y(_04686_),
    .A(_01164_),
    .B(_04685_));
 sg13g2_o21ai_1 _10467_ (.B1(_01241_),
    .Y(_04687_),
    .A1(_01163_),
    .A2(_01239_));
 sg13g2_xnor2_1 _10468_ (.Y(_04688_),
    .A(_01164_),
    .B(_04687_));
 sg13g2_nand3_1 _10469_ (.B(net3295),
    .C(net3287),
    .A(net3548),
    .Y(_04689_));
 sg13g2_nand2_1 _10470_ (.Y(_04690_),
    .A(net2962),
    .B(_04689_));
 sg13g2_o21ai_1 _10471_ (.B1(_04690_),
    .Y(_04691_),
    .A1(net3532),
    .A2(net2962));
 sg13g2_o21ai_1 _10472_ (.B1(net2857),
    .Y(_04692_),
    .A1(_00025_),
    .A2(_04691_));
 sg13g2_a22oi_1 _10473_ (.Y(_04693_),
    .B1(net2939),
    .B2(_04689_),
    .A2(net2955),
    .A1(_00637_));
 sg13g2_nand3_1 _10474_ (.B(_04692_),
    .C(_04693_),
    .A(net2945),
    .Y(_04694_));
 sg13g2_a21oi_1 _10475_ (.A1(net2933),
    .A2(_04689_),
    .Y(_04695_),
    .B1(net2945));
 sg13g2_o21ai_1 _10476_ (.B1(_04695_),
    .Y(_04696_),
    .A1(\core.work.alu.sval2[17] ),
    .A2(net2933));
 sg13g2_and2_1 _10477_ (.A(_00025_),
    .B(_04696_),
    .X(_04697_));
 sg13g2_o21ai_1 _10478_ (.B1(_04697_),
    .Y(_04698_),
    .A1(net2859),
    .A2(_04691_));
 sg13g2_nand2_1 _10479_ (.Y(_04699_),
    .A(net3460),
    .B(net3064));
 sg13g2_nand2_1 _10480_ (.Y(_04700_),
    .A(_00030_),
    .B(net3060));
 sg13g2_nand2_1 _10481_ (.Y(_04701_),
    .A(_04699_),
    .B(_04700_));
 sg13g2_nor2_1 _10482_ (.A(net2826),
    .B(_04701_),
    .Y(_04702_));
 sg13g2_nand2_1 _10483_ (.Y(_04703_),
    .A(_04537_),
    .B(_04623_));
 sg13g2_nor2_1 _10484_ (.A(net2823),
    .B(_04613_),
    .Y(_04704_));
 sg13g2_or2_1 _10485_ (.X(_04705_),
    .B(_04624_),
    .A(net2831));
 sg13g2_nor3_1 _10486_ (.A(net2794),
    .B(_04702_),
    .C(_04704_),
    .Y(_04706_));
 sg13g2_o21ai_1 _10487_ (.B1(_04705_),
    .Y(_04707_),
    .A1(net2835),
    .A2(_04703_));
 sg13g2_a221oi_1 _10488_ (.B2(_04698_),
    .C1(_04707_),
    .B1(_04694_),
    .A1(net2927),
    .Y(_04708_),
    .A2(_04688_));
 sg13g2_a221oi_1 _10489_ (.B2(_04708_),
    .C1(net3299),
    .B1(_04706_),
    .A1(net2797),
    .Y(_04709_),
    .A2(_04686_));
 sg13g2_nor2_1 _10490_ (.A(net3506),
    .B(_04123_),
    .Y(_04710_));
 sg13g2_nor2_1 _10491_ (.A(_00149_),
    .B(net2852),
    .Y(_04711_));
 sg13g2_or2_1 _10492_ (.X(_04712_),
    .B(_04711_),
    .A(_04519_));
 sg13g2_a21o_1 _10493_ (.A2(net2851),
    .A1(_04139_),
    .B1(_00157_),
    .X(_04713_));
 sg13g2_a21oi_1 _10494_ (.A1(\core.f2e_inst[9] ),
    .A2(_04637_),
    .Y(_04714_),
    .B1(_04712_));
 sg13g2_o21ai_1 _10495_ (.B1(net3162),
    .Y(_04715_),
    .A1(\core.f2e_inst[17] ),
    .A2(net3335));
 sg13g2_a21oi_2 _10496_ (.B1(_04715_),
    .Y(_04716_),
    .A2(_04714_),
    .A1(_04713_));
 sg13g2_a21oi_1 _10497_ (.A1(net2843),
    .A2(_03630_),
    .Y(_04717_),
    .B1(_04709_));
 sg13g2_nor2_2 _10498_ (.A(net2744),
    .B(_04716_),
    .Y(_04718_));
 sg13g2_a22oi_1 _10499_ (.Y(_00509_),
    .B1(_04717_),
    .B2(_04718_),
    .A2(net2750),
    .A1(_00628_));
 sg13g2_nor2_1 _10500_ (.A(net3532),
    .B(net3469),
    .Y(_04719_));
 sg13g2_a22oi_1 _10501_ (.Y(_04720_),
    .B1(net3535),
    .B2(net3471),
    .A2(net3469),
    .A1(net3532));
 sg13g2_nor2_1 _10502_ (.A(_04719_),
    .B(_04720_),
    .Y(_04721_));
 sg13g2_a21oi_1 _10503_ (.A1(_04652_),
    .A2(_04720_),
    .Y(_04722_),
    .B1(_04719_));
 sg13g2_xnor2_1 _10504_ (.Y(_04723_),
    .A(_01159_),
    .B(_04722_));
 sg13g2_a21oi_1 _10505_ (.A1(_01159_),
    .A2(_01243_),
    .Y(_04724_),
    .B1(_04012_));
 sg13g2_o21ai_1 _10506_ (.B1(_04724_),
    .Y(_04725_),
    .A1(_01159_),
    .A2(_01243_));
 sg13g2_nor2_1 _10507_ (.A(\core.work.alu.sval2[18] ),
    .B(net2962),
    .Y(_04726_));
 sg13g2_nand3_1 _10508_ (.B(net3295),
    .C(net3054),
    .A(net3548),
    .Y(_04727_));
 sg13g2_a21oi_1 _10509_ (.A1(net2962),
    .A2(_04727_),
    .Y(_04728_),
    .B1(_04726_));
 sg13g2_a21o_1 _10510_ (.A2(_04728_),
    .A1(_00638_),
    .B1(net2859),
    .X(_04729_));
 sg13g2_o21ai_1 _10511_ (.B1(net2945),
    .Y(_04730_),
    .A1(_00026_),
    .A2(net2953));
 sg13g2_a21oi_1 _10512_ (.A1(net2939),
    .A2(_04727_),
    .Y(_04731_),
    .B1(_04730_));
 sg13g2_a21oi_1 _10513_ (.A1(net2933),
    .A2(_04727_),
    .Y(_04732_),
    .B1(net2945));
 sg13g2_o21ai_1 _10514_ (.B1(_04732_),
    .Y(_04733_),
    .A1(\core.work.alu.sval2[18] ),
    .A2(net2934));
 sg13g2_a21oi_1 _10515_ (.A1(net2857),
    .A2(_04728_),
    .Y(_04734_),
    .B1(_00638_));
 sg13g2_a22oi_1 _10516_ (.Y(_04735_),
    .B1(_04733_),
    .B2(_04734_),
    .A2(_04731_),
    .A1(_04729_));
 sg13g2_nor2_1 _10517_ (.A(net2823),
    .B(_04665_),
    .Y(_04736_));
 sg13g2_nand2_1 _10518_ (.Y(_04737_),
    .A(_00033_),
    .B(net3064));
 sg13g2_nand2_1 _10519_ (.Y(_04738_),
    .A(net3460),
    .B(net3060));
 sg13g2_nand2_1 _10520_ (.Y(_04739_),
    .A(_04737_),
    .B(_04738_));
 sg13g2_nand2_1 _10521_ (.Y(_04740_),
    .A(_04582_),
    .B(_04669_));
 sg13g2_or2_1 _10522_ (.X(_04741_),
    .B(_04740_),
    .A(net2835));
 sg13g2_o21ai_1 _10523_ (.B1(net2790),
    .Y(_04742_),
    .A1(net2831),
    .A2(_04670_));
 sg13g2_o21ai_1 _10524_ (.B1(_04741_),
    .Y(_04743_),
    .A1(net2826),
    .A2(_04739_));
 sg13g2_nor4_1 _10525_ (.A(_04735_),
    .B(_04736_),
    .C(_04742_),
    .D(_04743_),
    .Y(_04744_));
 sg13g2_a22oi_1 _10526_ (.Y(_04745_),
    .B1(_04725_),
    .B2(_04744_),
    .A2(_04723_),
    .A1(net2794));
 sg13g2_nand2_1 _10527_ (.Y(_04746_),
    .A(net3309),
    .B(_04745_));
 sg13g2_nor2_1 _10528_ (.A(_00158_),
    .B(_04139_),
    .Y(_04747_));
 sg13g2_a21oi_1 _10529_ (.A1(net3508),
    .A2(_04636_),
    .Y(_04748_),
    .B1(_04747_));
 sg13g2_nor2_1 _10530_ (.A(_04213_),
    .B(_04712_),
    .Y(_04749_));
 sg13g2_a22oi_1 _10531_ (.Y(_04750_),
    .B1(_04748_),
    .B2(_04749_),
    .A2(net3343),
    .A1(_00678_));
 sg13g2_a221oi_1 _10532_ (.B2(net3165),
    .C1(net2745),
    .B1(_04750_),
    .A1(net2842),
    .Y(_04751_),
    .A2(_03651_));
 sg13g2_a22oi_1 _10533_ (.Y(_00510_),
    .B1(_04746_),
    .B2(_04751_),
    .A2(net2750),
    .A1(_00626_));
 sg13g2_a21oi_1 _10534_ (.A1(_01159_),
    .A2(_04722_),
    .Y(_04752_),
    .B1(_01158_));
 sg13g2_xor2_1 _10535_ (.B(_04752_),
    .A(_01157_),
    .X(_04753_));
 sg13g2_o21ai_1 _10536_ (.B1(_01244_),
    .Y(_04754_),
    .A1(_01159_),
    .A2(_01243_));
 sg13g2_xor2_1 _10537_ (.B(_04754_),
    .A(_01157_),
    .X(_04755_));
 sg13g2_nand3_1 _10538_ (.B(net3295),
    .C(net3291),
    .A(net3548),
    .Y(_04756_));
 sg13g2_nor2_1 _10539_ (.A(\core.work.alu.sval2[19] ),
    .B(net2962),
    .Y(_04757_));
 sg13g2_a21oi_1 _10540_ (.A1(net2962),
    .A2(_04756_),
    .Y(_04758_),
    .B1(_04757_));
 sg13g2_a21o_1 _10541_ (.A2(_04758_),
    .A1(_00639_),
    .B1(net2859),
    .X(_04759_));
 sg13g2_o21ai_1 _10542_ (.B1(net2945),
    .Y(_04760_),
    .A1(_00029_),
    .A2(net2953));
 sg13g2_a21oi_1 _10543_ (.A1(net2939),
    .A2(_04756_),
    .Y(_04761_),
    .B1(_04760_));
 sg13g2_a21oi_1 _10544_ (.A1(net2933),
    .A2(_04756_),
    .Y(_04762_),
    .B1(net2945));
 sg13g2_o21ai_1 _10545_ (.B1(_04762_),
    .Y(_04763_),
    .A1(\core.work.alu.sval2[19] ),
    .A2(net2933));
 sg13g2_a21oi_1 _10546_ (.A1(net2857),
    .A2(_04758_),
    .Y(_04764_),
    .B1(_00639_));
 sg13g2_a22oi_1 _10547_ (.Y(_04765_),
    .B1(_04763_),
    .B2(_04764_),
    .A2(_04761_),
    .A1(_04759_));
 sg13g2_or2_1 _10548_ (.X(_04766_),
    .B(_04703_),
    .A(net2823));
 sg13g2_o21ai_1 _10549_ (.B1(_04766_),
    .Y(_04767_),
    .A1(net2831),
    .A2(_04701_));
 sg13g2_nand2_1 _10550_ (.Y(_04768_),
    .A(_04622_),
    .B(_04700_));
 sg13g2_nand2_1 _10551_ (.Y(_04769_),
    .A(_00036_),
    .B(net3062));
 sg13g2_nand2_1 _10552_ (.Y(_04770_),
    .A(_00033_),
    .B(net3056));
 sg13g2_nand2_1 _10553_ (.Y(_04771_),
    .A(_04769_),
    .B(_04770_));
 sg13g2_or2_1 _10554_ (.X(_04772_),
    .B(_04771_),
    .A(net2826));
 sg13g2_o21ai_1 _10555_ (.B1(_04772_),
    .Y(_04773_),
    .A1(net2835),
    .A2(_04768_));
 sg13g2_nor4_1 _10556_ (.A(net2794),
    .B(_04765_),
    .C(_04767_),
    .D(_04773_),
    .Y(_04774_));
 sg13g2_o21ai_1 _10557_ (.B1(_04774_),
    .Y(_04775_),
    .A1(_04012_),
    .A2(_04755_));
 sg13g2_a21oi_1 _10558_ (.A1(net2794),
    .A2(_04753_),
    .Y(_04776_),
    .B1(net3299));
 sg13g2_a22oi_1 _10559_ (.Y(_04777_),
    .B1(_04775_),
    .B2(_04776_),
    .A2(_03674_),
    .A1(net2843));
 sg13g2_a21oi_1 _10560_ (.A1(\core.f2e_inst[11] ),
    .A2(_04636_),
    .Y(_04778_),
    .B1(_04712_));
 sg13g2_o21ai_1 _10561_ (.B1(_04778_),
    .Y(_04779_),
    .A1(_00152_),
    .A2(_04139_));
 sg13g2_o21ai_1 _10562_ (.B1(_04779_),
    .Y(_04780_),
    .A1(\core.f2e_inst[19] ),
    .A2(net3335));
 sg13g2_nor3_2 _10563_ (.A(net3161),
    .B(net2744),
    .C(_04780_),
    .Y(_04781_));
 sg13g2_a21oi_1 _10564_ (.A1(net824),
    .A2(net2750),
    .Y(_04782_),
    .B1(_04781_));
 sg13g2_o21ai_1 _10565_ (.B1(_04782_),
    .Y(_00511_),
    .A1(_04060_),
    .A2(_04777_));
 sg13g2_and2_1 _10566_ (.A(_01157_),
    .B(_01159_),
    .X(_04783_));
 sg13g2_and3_1 _10567_ (.X(_04784_),
    .A(_01163_),
    .B(_01164_),
    .C(_04783_));
 sg13g2_a21oi_1 _10568_ (.A1(\core.e2m_addr[19] ),
    .A2(net3531),
    .Y(_04785_),
    .B1(_01158_));
 sg13g2_a21oi_1 _10569_ (.A1(_00623_),
    .A2(_00624_),
    .Y(_04786_),
    .B1(_04785_));
 sg13g2_a221oi_1 _10570_ (.B2(_04651_),
    .C1(_04786_),
    .B1(_04784_),
    .A1(_04721_),
    .Y(_04787_),
    .A2(_04783_));
 sg13g2_or2_1 _10571_ (.X(_04788_),
    .B(_04787_),
    .A(_01153_));
 sg13g2_xnor2_1 _10572_ (.Y(_04789_),
    .A(_01153_),
    .B(_04787_));
 sg13g2_nor2_1 _10573_ (.A(_01153_),
    .B(_01247_),
    .Y(_04790_));
 sg13g2_nand2_1 _10574_ (.Y(_04791_),
    .A(_01153_),
    .B(_01247_));
 sg13g2_nand2_1 _10575_ (.Y(_04792_),
    .A(net3452),
    .B(net3062));
 sg13g2_nand2_1 _10576_ (.Y(_04793_),
    .A(_00036_),
    .B(net3056));
 sg13g2_nand2_1 _10577_ (.Y(_04794_),
    .A(_04792_),
    .B(_04793_));
 sg13g2_nor2_1 _10578_ (.A(net2826),
    .B(_04794_),
    .Y(_04795_));
 sg13g2_nand2_1 _10579_ (.Y(_04796_),
    .A(_04668_),
    .B(_04738_));
 sg13g2_nor2_1 _10580_ (.A(net2835),
    .B(_04796_),
    .Y(_04797_));
 sg13g2_nor2_1 _10581_ (.A(net2832),
    .B(_04739_),
    .Y(_04798_));
 sg13g2_nand2_2 _10582_ (.Y(_04799_),
    .A(net3548),
    .B(_04176_));
 sg13g2_o21ai_1 _10583_ (.B1(net2945),
    .Y(_04800_),
    .A1(_00031_),
    .A2(net2953));
 sg13g2_a21oi_1 _10584_ (.A1(net2939),
    .A2(_04799_),
    .Y(_04801_),
    .B1(_04800_));
 sg13g2_nor2_1 _10585_ (.A(net2823),
    .B(_04740_),
    .Y(_04802_));
 sg13g2_o21ai_1 _10586_ (.B1(net2951),
    .Y(_04803_),
    .A1(net3530),
    .A2(net2934));
 sg13g2_a21oi_1 _10587_ (.A1(net2933),
    .A2(_04799_),
    .Y(_04804_),
    .B1(_04803_));
 sg13g2_nor3_1 _10588_ (.A(net2794),
    .B(_04802_),
    .C(_04804_),
    .Y(_04805_));
 sg13g2_o21ai_1 _10589_ (.B1(_04805_),
    .Y(_04806_),
    .A1(_00032_),
    .A2(_04801_));
 sg13g2_nor4_1 _10590_ (.A(_04795_),
    .B(_04797_),
    .C(_04798_),
    .D(_04806_),
    .Y(_04807_));
 sg13g2_nor2_1 _10591_ (.A(net3530),
    .B(net2963),
    .Y(_04808_));
 sg13g2_a21oi_1 _10592_ (.A1(net2963),
    .A2(_04799_),
    .Y(_04809_),
    .B1(_04808_));
 sg13g2_xnor2_1 _10593_ (.Y(_04810_),
    .A(_00032_),
    .B(_04809_));
 sg13g2_nor2_1 _10594_ (.A(net2924),
    .B(_04790_),
    .Y(_04811_));
 sg13g2_a22oi_1 _10595_ (.Y(_04812_),
    .B1(_04811_),
    .B2(_04791_),
    .A2(_04810_),
    .A1(net2857));
 sg13g2_a221oi_1 _10596_ (.B2(_04812_),
    .C1(net3300),
    .B1(_04807_),
    .A1(net2794),
    .Y(_04813_),
    .A2(_04789_));
 sg13g2_or4_1 _10597_ (.A(_04215_),
    .B(_04226_),
    .C(_04227_),
    .D(_04445_),
    .X(_04814_));
 sg13g2_a21oi_1 _10598_ (.A1(\core.f2e_inst[2] ),
    .A2(_04814_),
    .Y(_04815_),
    .B1(_04712_));
 sg13g2_o21ai_1 _10599_ (.B1(_04815_),
    .Y(_04816_),
    .A1(_00159_),
    .A2(_04224_));
 sg13g2_o21ai_1 _10600_ (.B1(net3163),
    .Y(_04817_),
    .A1(\core.f2e_inst[20] ),
    .A2(net3338));
 sg13g2_inv_1 _10601_ (.Y(_04818_),
    .A(_04817_));
 sg13g2_a21oi_2 _10602_ (.B1(net2744),
    .Y(_04819_),
    .A2(_04818_),
    .A1(_04816_));
 sg13g2_a21oi_1 _10603_ (.A1(net2843),
    .A2(_03699_),
    .Y(_04820_),
    .B1(_04813_));
 sg13g2_a22oi_1 _10604_ (.Y(_00512_),
    .B1(_04819_),
    .B2(_04820_),
    .A2(net2750),
    .A1(_00622_));
 sg13g2_o21ai_1 _10605_ (.B1(_04788_),
    .Y(_04821_),
    .A1(_00621_),
    .A2(_00622_));
 sg13g2_xor2_1 _10606_ (.B(_04821_),
    .A(_01154_),
    .X(_04822_));
 sg13g2_nand2b_1 _10607_ (.Y(_04823_),
    .B(_04791_),
    .A_N(_01248_));
 sg13g2_xnor2_1 _10608_ (.Y(_04824_),
    .A(_01154_),
    .B(_04823_));
 sg13g2_nor2_1 _10609_ (.A(net2924),
    .B(_04824_),
    .Y(_04825_));
 sg13g2_nor2_1 _10610_ (.A(\core.work.alu.sval2[21] ),
    .B(net2963),
    .Y(_04826_));
 sg13g2_nand2_2 _10611_ (.Y(_04827_),
    .A(net3548),
    .B(_04234_));
 sg13g2_a21oi_1 _10612_ (.A1(net2963),
    .A2(_04827_),
    .Y(_04828_),
    .B1(_04826_));
 sg13g2_o21ai_1 _10613_ (.B1(net2857),
    .Y(_04829_),
    .A1(_00640_),
    .A2(_04828_));
 sg13g2_a21oi_1 _10614_ (.A1(_00640_),
    .A2(_04828_),
    .Y(_04830_),
    .B1(_04829_));
 sg13g2_a22oi_1 _10615_ (.Y(_04831_),
    .B1(net2939),
    .B2(_04827_),
    .A2(net2955),
    .A1(_00641_));
 sg13g2_a21oi_1 _10616_ (.A1(net2946),
    .A2(_04831_),
    .Y(_04832_),
    .B1(_00033_));
 sg13g2_nor2_1 _10617_ (.A(net2831),
    .B(_04771_),
    .Y(_04833_));
 sg13g2_o21ai_1 _10618_ (.B1(net2790),
    .Y(_04834_),
    .A1(net2823),
    .A2(_04768_));
 sg13g2_nor3_1 _10619_ (.A(_04832_),
    .B(_04833_),
    .C(_04834_),
    .Y(_04835_));
 sg13g2_o21ai_1 _10620_ (.B1(net2951),
    .Y(_04836_),
    .A1(\core.work.alu.sval2[21] ),
    .A2(net2934));
 sg13g2_a21oi_1 _10621_ (.A1(net2934),
    .A2(_04827_),
    .Y(_04837_),
    .B1(_04836_));
 sg13g2_nand2_1 _10622_ (.Y(_04838_),
    .A(_00040_),
    .B(net3062));
 sg13g2_nand2_1 _10623_ (.Y(_04839_),
    .A(net3452),
    .B(net3056));
 sg13g2_nand2_1 _10624_ (.Y(_04840_),
    .A(_04838_),
    .B(_04839_));
 sg13g2_nand3_1 _10625_ (.B(_04699_),
    .C(_04770_),
    .A(_03990_),
    .Y(_04841_));
 sg13g2_o21ai_1 _10626_ (.B1(_04841_),
    .Y(_04842_),
    .A1(net2825),
    .A2(_04840_));
 sg13g2_nor4_1 _10627_ (.A(_04825_),
    .B(_04830_),
    .C(_04837_),
    .D(_04842_),
    .Y(_04843_));
 sg13g2_a221oi_1 _10628_ (.B2(_04843_),
    .C1(net3299),
    .B1(_04835_),
    .A1(net2794),
    .Y(_04844_),
    .A2(_04822_));
 sg13g2_nor2_1 _10629_ (.A(_04130_),
    .B(_04226_),
    .Y(_04845_));
 sg13g2_nor3_1 _10630_ (.A(\core.f2e_inst[15] ),
    .B(_04121_),
    .C(_04122_),
    .Y(_04846_));
 sg13g2_nor4_1 _10631_ (.A(_04210_),
    .B(_04215_),
    .C(_04227_),
    .D(_04846_),
    .Y(_04847_));
 sg13g2_a21oi_1 _10632_ (.A1(_04845_),
    .A2(_04847_),
    .Y(_04848_),
    .B1(_00683_));
 sg13g2_nor2_1 _10633_ (.A(_00160_),
    .B(_04224_),
    .Y(_04849_));
 sg13g2_or4_1 _10634_ (.A(net3346),
    .B(_04711_),
    .C(_04848_),
    .D(_04849_),
    .X(_04850_));
 sg13g2_a21oi_2 _10635_ (.B1(net3160),
    .Y(_04851_),
    .A2(net3347),
    .A1(_00687_));
 sg13g2_a21oi_1 _10636_ (.A1(net2843),
    .A2(_03719_),
    .Y(_04852_),
    .B1(_04844_));
 sg13g2_a21oi_2 _10637_ (.B1(net2744),
    .Y(_04853_),
    .A2(_04851_),
    .A1(_04850_));
 sg13g2_a22oi_1 _10638_ (.Y(_00513_),
    .B1(_04852_),
    .B2(_04853_),
    .A2(net2751),
    .A1(_00620_));
 sg13g2_a22oi_1 _10639_ (.Y(_04854_),
    .B1(net3530),
    .B2(net3465),
    .A2(net3457),
    .A1(\core.work.alu.sval2[21] ));
 sg13g2_a21oi_1 _10640_ (.A1(_00619_),
    .A2(_00620_),
    .Y(_04855_),
    .B1(_04854_));
 sg13g2_inv_1 _10641_ (.Y(_04856_),
    .A(_04855_));
 sg13g2_o21ai_1 _10642_ (.B1(_04856_),
    .Y(_04857_),
    .A1(_01154_),
    .A2(_04788_));
 sg13g2_xor2_1 _10643_ (.B(_04857_),
    .A(_01151_),
    .X(_04858_));
 sg13g2_a21oi_1 _10644_ (.A1(_01249_),
    .A2(_04791_),
    .Y(_04859_),
    .B1(_01250_));
 sg13g2_nand2b_1 _10645_ (.Y(_04860_),
    .B(_04859_),
    .A_N(_01151_));
 sg13g2_xnor2_1 _10646_ (.Y(_04861_),
    .A(_01151_),
    .B(_04859_));
 sg13g2_nor2_1 _10647_ (.A(\core.work.alu.sval2[22] ),
    .B(net2958),
    .Y(_04862_));
 sg13g2_nand2_2 _10648_ (.Y(_04863_),
    .A(net3548),
    .B(_04266_));
 sg13g2_a21oi_1 _10649_ (.A1(net2958),
    .A2(_04863_),
    .Y(_04864_),
    .B1(_04862_));
 sg13g2_xnor2_1 _10650_ (.Y(_04865_),
    .A(_00036_),
    .B(_04864_));
 sg13g2_nor2_1 _10651_ (.A(net2823),
    .B(_04796_),
    .Y(_04866_));
 sg13g2_nor2_1 _10652_ (.A(\core.work.alu.sval2[22] ),
    .B(net2931),
    .Y(_04867_));
 sg13g2_a21oi_1 _10653_ (.A1(net2931),
    .A2(_04863_),
    .Y(_04868_),
    .B1(_04867_));
 sg13g2_a21oi_1 _10654_ (.A1(net2937),
    .A2(_04863_),
    .Y(_04869_),
    .B1(net2949));
 sg13g2_o21ai_1 _10655_ (.B1(_04869_),
    .Y(_04870_),
    .A1(_00034_),
    .A2(net2952));
 sg13g2_nand2_1 _10656_ (.Y(_04871_),
    .A(_04737_),
    .B(_04793_));
 sg13g2_nor2_1 _10657_ (.A(net2835),
    .B(_04871_),
    .Y(_04872_));
 sg13g2_nand2_1 _10658_ (.Y(_04873_),
    .A(_00040_),
    .B(net3055));
 sg13g2_nand2_1 _10659_ (.Y(_04874_),
    .A(_00041_),
    .B(net3061));
 sg13g2_nand2_1 _10660_ (.Y(_04875_),
    .A(_04873_),
    .B(_04874_));
 sg13g2_o21ai_1 _10661_ (.B1(net2790),
    .Y(_04876_),
    .A1(net2831),
    .A2(_04794_));
 sg13g2_nor3_1 _10662_ (.A(_04866_),
    .B(_04872_),
    .C(_04876_),
    .Y(_04877_));
 sg13g2_a22oi_1 _10663_ (.Y(_04878_),
    .B1(_04870_),
    .B2(_00642_),
    .A2(_04868_),
    .A1(net2950));
 sg13g2_o21ai_1 _10664_ (.B1(_04878_),
    .Y(_04879_),
    .A1(net2825),
    .A2(_04875_));
 sg13g2_a221oi_1 _10665_ (.B2(net2855),
    .C1(_04879_),
    .B1(_04865_),
    .A1(net2927),
    .Y(_04880_),
    .A2(_04861_));
 sg13g2_a21oi_1 _10666_ (.A1(_04877_),
    .A2(_04880_),
    .Y(_04881_),
    .B1(net3299));
 sg13g2_o21ai_1 _10667_ (.B1(_04881_),
    .Y(_04882_),
    .A1(net2790),
    .A2(_04858_));
 sg13g2_a21oi_1 _10668_ (.A1(net2841),
    .A2(_03745_),
    .Y(_04883_),
    .B1(net3163));
 sg13g2_nand3b_1 _10669_ (.B(net3510),
    .C(net3336),
    .Y(_04884_),
    .A_N(_04324_));
 sg13g2_nor3_1 _10670_ (.A(_04215_),
    .B(_04217_),
    .C(_04846_),
    .Y(_04885_));
 sg13g2_nand3b_1 _10671_ (.B(_04845_),
    .C(_04885_),
    .Y(_04886_),
    .A_N(_04210_));
 sg13g2_o21ai_1 _10672_ (.B1(net3162),
    .Y(_04887_),
    .A1(net3506),
    .A2(net2852));
 sg13g2_a21oi_1 _10673_ (.A1(\core.f2e_inst[22] ),
    .A2(net3343),
    .Y(_04888_),
    .B1(_04887_));
 sg13g2_o21ai_1 _10674_ (.B1(_04888_),
    .Y(_04889_),
    .A1(_00161_),
    .A2(_04224_));
 sg13g2_a21oi_1 _10675_ (.A1(\core.f2e_inst[4] ),
    .A2(_04886_),
    .Y(_04890_),
    .B1(_04889_));
 sg13g2_a221oi_1 _10676_ (.B2(_04890_),
    .C1(net2742),
    .B1(_04884_),
    .A1(_04882_),
    .Y(_04891_),
    .A2(_04883_));
 sg13g2_a21o_1 _10677_ (.A2(net2742),
    .A1(net3456),
    .B1(_04891_),
    .X(_00514_));
 sg13g2_a21oi_1 _10678_ (.A1(_01151_),
    .A2(_04857_),
    .Y(_04892_),
    .B1(_01150_));
 sg13g2_xnor2_1 _10679_ (.Y(_04893_),
    .A(_01149_),
    .B(_04892_));
 sg13g2_nand2_1 _10680_ (.Y(_04894_),
    .A(_01252_),
    .B(_04860_));
 sg13g2_xnor2_1 _10681_ (.Y(_04895_),
    .A(_01149_),
    .B(_04894_));
 sg13g2_nand2_2 _10682_ (.Y(_04896_),
    .A(net3550),
    .B(_04302_));
 sg13g2_o21ai_1 _10683_ (.B1(net3452),
    .Y(_04897_),
    .A1(_03994_),
    .A2(_04896_));
 sg13g2_a21oi_1 _10684_ (.A1(\core.work.alu.sval2[23] ),
    .A2(_03994_),
    .Y(_04898_),
    .B1(_04897_));
 sg13g2_a22oi_1 _10685_ (.Y(_04899_),
    .B1(net2938),
    .B2(_04896_),
    .A2(net2954),
    .A1(_00643_));
 sg13g2_or2_1 _10686_ (.X(_04900_),
    .B(_04840_),
    .A(net2829));
 sg13g2_nand2_1 _10687_ (.Y(_04901_),
    .A(_00044_),
    .B(net3061));
 sg13g2_nand2_1 _10688_ (.Y(_04902_),
    .A(_00041_),
    .B(net3055));
 sg13g2_nand2_1 _10689_ (.Y(_04903_),
    .A(_04901_),
    .B(_04902_));
 sg13g2_o21ai_1 _10690_ (.B1(_04900_),
    .Y(_04904_),
    .A1(net2825),
    .A2(_04903_));
 sg13g2_nand4_1 _10691_ (.B(net2853),
    .C(_04699_),
    .A(_01716_),
    .Y(_04905_),
    .D(_04770_));
 sg13g2_nand2_1 _10692_ (.Y(_04906_),
    .A(_04769_),
    .B(_04839_));
 sg13g2_o21ai_1 _10693_ (.B1(_04905_),
    .Y(_04907_),
    .A1(net2834),
    .A2(_04906_));
 sg13g2_o21ai_1 _10694_ (.B1(net2788),
    .Y(_04908_),
    .A1(net3452),
    .A2(_04899_));
 sg13g2_nor2_1 _10695_ (.A(net2944),
    .B(_04898_),
    .Y(_04909_));
 sg13g2_nor4_1 _10696_ (.A(_04904_),
    .B(_04907_),
    .C(_04908_),
    .D(_04909_),
    .Y(_04910_));
 sg13g2_nor2_1 _10697_ (.A(\core.work.alu.sval2[23] ),
    .B(net2961),
    .Y(_04911_));
 sg13g2_a21oi_1 _10698_ (.A1(net2958),
    .A2(_04896_),
    .Y(_04912_),
    .B1(_04911_));
 sg13g2_xnor2_1 _10699_ (.Y(_04913_),
    .A(net3452),
    .B(_04912_));
 sg13g2_a22oi_1 _10700_ (.Y(_04914_),
    .B1(_04913_),
    .B2(net2855),
    .A2(_04895_),
    .A1(net2926));
 sg13g2_a21oi_1 _10701_ (.A1(_04910_),
    .A2(_04914_),
    .Y(_04915_),
    .B1(net3299));
 sg13g2_o21ai_1 _10702_ (.B1(_04915_),
    .Y(_04916_),
    .A1(net2790),
    .A2(_04893_));
 sg13g2_a21oi_1 _10703_ (.A1(net2841),
    .A2(_03765_),
    .Y(_04917_),
    .B1(net3162));
 sg13g2_nand3_1 _10704_ (.B(_04845_),
    .C(_04885_),
    .A(_04221_),
    .Y(_04918_));
 sg13g2_nand3_1 _10705_ (.B(net3336),
    .C(_04918_),
    .A(net3511),
    .Y(_04919_));
 sg13g2_nor2_1 _10706_ (.A(_00162_),
    .B(_04224_),
    .Y(_04920_));
 sg13g2_a22oi_1 _10707_ (.Y(_04921_),
    .B1(_04209_),
    .B2(net3509),
    .A2(net3347),
    .A1(\core.f2e_inst[23] ));
 sg13g2_nand2_1 _10708_ (.Y(_04922_),
    .A(_04259_),
    .B(_04921_));
 sg13g2_nor3_2 _10709_ (.A(_04887_),
    .B(_04920_),
    .C(_04922_),
    .Y(_04923_));
 sg13g2_a22oi_1 _10710_ (.Y(_04924_),
    .B1(_04919_),
    .B2(_04923_),
    .A2(_04917_),
    .A1(_04916_));
 sg13g2_mux2_1 _10711_ (.A0(_04924_),
    .A1(net3454),
    .S(net2742),
    .X(_00515_));
 sg13g2_and2_1 _10712_ (.A(_01149_),
    .B(_01151_),
    .X(_04925_));
 sg13g2_nor2_1 _10713_ (.A(_01153_),
    .B(_01154_),
    .Y(_04926_));
 sg13g2_nand2_1 _10714_ (.Y(_04927_),
    .A(_04925_),
    .B(_04926_));
 sg13g2_o21ai_1 _10715_ (.B1(_01150_),
    .Y(_04928_),
    .A1(net3534),
    .A2(net3453));
 sg13g2_inv_1 _10716_ (.Y(_04929_),
    .A(_04928_));
 sg13g2_a221oi_1 _10717_ (.B2(_04925_),
    .C1(_04929_),
    .B1(_04855_),
    .A1(net3534),
    .Y(_04930_),
    .A2(net3453));
 sg13g2_o21ai_1 _10718_ (.B1(_04930_),
    .Y(_04931_),
    .A1(_04787_),
    .A2(_04927_));
 sg13g2_nand2_1 _10719_ (.Y(_04932_),
    .A(_01263_),
    .B(_04931_));
 sg13g2_xnor2_1 _10720_ (.Y(_04933_),
    .A(_01263_),
    .B(_04931_));
 sg13g2_nor2_1 _10721_ (.A(_01255_),
    .B(_01263_),
    .Y(_04934_));
 sg13g2_nand3_1 _10722_ (.B(net3296),
    .C(net3289),
    .A(net3547),
    .Y(_04935_));
 sg13g2_nor2_1 _10723_ (.A(net3533),
    .B(net2956),
    .Y(_04936_));
 sg13g2_a21oi_1 _10724_ (.A1(net2961),
    .A2(_04935_),
    .Y(_04937_),
    .B1(_04936_));
 sg13g2_xnor2_1 _10725_ (.Y(_04938_),
    .A(_00040_),
    .B(_04937_));
 sg13g2_nand2_1 _10726_ (.Y(_04939_),
    .A(_00044_),
    .B(net3055));
 sg13g2_nand2_1 _10727_ (.Y(_04940_),
    .A(_00046_),
    .B(net3061));
 sg13g2_nand2_1 _10728_ (.Y(_04941_),
    .A(_04939_),
    .B(_04940_));
 sg13g2_nor2_1 _10729_ (.A(net2825),
    .B(_04941_),
    .Y(_04942_));
 sg13g2_o21ai_1 _10730_ (.B1(net2949),
    .Y(_04943_),
    .A1(net3533),
    .A2(net2930));
 sg13g2_a21oi_1 _10731_ (.A1(net2930),
    .A2(_04935_),
    .Y(_04944_),
    .B1(_04943_));
 sg13g2_nor2_1 _10732_ (.A(net2829),
    .B(_04875_),
    .Y(_04945_));
 sg13g2_o21ai_1 _10733_ (.B1(net2942),
    .Y(_04946_),
    .A1(_00039_),
    .A2(net2952));
 sg13g2_a21oi_1 _10734_ (.A1(net2937),
    .A2(_04935_),
    .Y(_04947_),
    .B1(_04946_));
 sg13g2_nand2_1 _10735_ (.Y(_04948_),
    .A(_04792_),
    .B(_04873_));
 sg13g2_nor2_1 _10736_ (.A(net2833),
    .B(_04948_),
    .Y(_04949_));
 sg13g2_nor2_1 _10737_ (.A(_04942_),
    .B(_04945_),
    .Y(_04950_));
 sg13g2_o21ai_1 _10738_ (.B1(net2790),
    .Y(_04951_),
    .A1(net2821),
    .A2(_04871_));
 sg13g2_nor3_1 _10739_ (.A(_04944_),
    .B(_04949_),
    .C(_04951_),
    .Y(_04952_));
 sg13g2_o21ai_1 _10740_ (.B1(_04950_),
    .Y(_04953_),
    .A1(_00040_),
    .A2(_04947_));
 sg13g2_xor2_1 _10741_ (.B(_01263_),
    .A(_01255_),
    .X(_04954_));
 sg13g2_a221oi_1 _10742_ (.B2(net2926),
    .C1(_04953_),
    .B1(_04954_),
    .A1(net2855),
    .Y(_04955_),
    .A2(_04938_));
 sg13g2_a22oi_1 _10743_ (.Y(_04956_),
    .B1(_04952_),
    .B2(_04955_),
    .A2(_04933_),
    .A1(net2793));
 sg13g2_a221oi_1 _10744_ (.B2(net3303),
    .C1(net3164),
    .B1(_04956_),
    .A1(net2842),
    .Y(_04957_),
    .A2(_03796_));
 sg13g2_nor2_1 _10745_ (.A(_00699_),
    .B(net3345),
    .Y(_04958_));
 sg13g2_o21ai_1 _10746_ (.B1(_04958_),
    .Y(_04959_),
    .A1(_04209_),
    .A2(_04220_));
 sg13g2_nand3_1 _10747_ (.B(_00699_),
    .C(_04204_),
    .A(net3508),
    .Y(_04960_));
 sg13g2_a21oi_1 _10748_ (.A1(net3507),
    .A2(_04137_),
    .Y(_04961_),
    .B1(_04219_));
 sg13g2_nand3_1 _10749_ (.B(_04960_),
    .C(_04961_),
    .A(_04222_),
    .Y(_04962_));
 sg13g2_o21ai_1 _10750_ (.B1(_04370_),
    .Y(_04963_),
    .A1(net3508),
    .A2(net2851));
 sg13g2_nand2b_1 _10751_ (.Y(_04964_),
    .B(_04963_),
    .A_N(_00150_));
 sg13g2_a21oi_1 _10752_ (.A1(\core.f2e_inst[24] ),
    .A2(net3343),
    .Y(_04965_),
    .B1(_04887_));
 sg13g2_nand3_1 _10753_ (.B(_04964_),
    .C(_04965_),
    .A(_04959_),
    .Y(_04966_));
 sg13g2_a21oi_2 _10754_ (.B1(_04966_),
    .Y(_04967_),
    .A2(_04962_),
    .A1(net3510));
 sg13g2_nor3_1 _10755_ (.A(net2745),
    .B(_04957_),
    .C(_04967_),
    .Y(_04968_));
 sg13g2_a21o_1 _10756_ (.A2(net2745),
    .A1(net3451),
    .B1(_04968_),
    .X(_00516_));
 sg13g2_o21ai_1 _10757_ (.B1(_04932_),
    .Y(_04969_),
    .A1(_00614_),
    .A2(_00615_));
 sg13g2_xnor2_1 _10758_ (.Y(_04970_),
    .A(_01266_),
    .B(_04969_));
 sg13g2_nor2_1 _10759_ (.A(_01262_),
    .B(_04934_),
    .Y(_04971_));
 sg13g2_xor2_1 _10760_ (.B(_04971_),
    .A(_01266_),
    .X(_04972_));
 sg13g2_nand3_1 _10761_ (.B(net3296),
    .C(net3288),
    .A(net3547),
    .Y(_04973_));
 sg13g2_nor2_1 _10762_ (.A(\core.work.alu.sval2[25] ),
    .B(net2956),
    .Y(_04974_));
 sg13g2_a21oi_1 _10763_ (.A1(net2957),
    .A2(_04973_),
    .Y(_04975_),
    .B1(_04974_));
 sg13g2_xnor2_1 _10764_ (.Y(_04976_),
    .A(_00041_),
    .B(_04975_));
 sg13g2_nor2_1 _10765_ (.A(net2829),
    .B(_04903_),
    .Y(_04977_));
 sg13g2_nor2_1 _10766_ (.A(_00048_),
    .B(net3055),
    .Y(_04978_));
 sg13g2_nor2_1 _10767_ (.A(_00046_),
    .B(net3061),
    .Y(_04979_));
 sg13g2_o21ai_1 _10768_ (.B1(_04015_),
    .Y(_04980_),
    .A1(_04978_),
    .A2(_04979_));
 sg13g2_nand2_1 _10769_ (.Y(_04981_),
    .A(_04838_),
    .B(_04902_));
 sg13g2_nor2_1 _10770_ (.A(net2928),
    .B(_04973_),
    .Y(_04982_));
 sg13g2_a21oi_1 _10771_ (.A1(net3536),
    .A2(net2928),
    .Y(_04983_),
    .B1(_04982_));
 sg13g2_a21oi_1 _10772_ (.A1(_00041_),
    .A2(_04983_),
    .Y(_04984_),
    .B1(net2942));
 sg13g2_a22oi_1 _10773_ (.Y(_04985_),
    .B1(net2937),
    .B2(_04973_),
    .A2(net2954),
    .A1(_00644_));
 sg13g2_nor2_1 _10774_ (.A(_00041_),
    .B(_04985_),
    .Y(_04986_));
 sg13g2_nor4_1 _10775_ (.A(net2792),
    .B(_04977_),
    .C(_04984_),
    .D(_04986_),
    .Y(_04987_));
 sg13g2_o21ai_1 _10776_ (.B1(_04980_),
    .Y(_04988_),
    .A1(net2822),
    .A2(_04906_));
 sg13g2_inv_1 _10777_ (.Y(_04989_),
    .A(_04988_));
 sg13g2_o21ai_1 _10778_ (.B1(_04989_),
    .Y(_04990_),
    .A1(net2833),
    .A2(_04981_));
 sg13g2_a221oi_1 _10779_ (.B2(net2854),
    .C1(_04990_),
    .B1(_04976_),
    .A1(net2925),
    .Y(_04991_),
    .A2(_04972_));
 sg13g2_a221oi_1 _10780_ (.B2(_04991_),
    .C1(net3297),
    .B1(_04987_),
    .A1(net2792),
    .Y(_04992_),
    .A2(_04970_));
 sg13g2_a221oi_1 _10781_ (.B2(_03818_),
    .C1(_04992_),
    .B1(net2842),
    .A1(net3329),
    .Y(_04993_),
    .A2(net3297));
 sg13g2_a221oi_1 _10782_ (.B2(_04448_),
    .C1(_00701_),
    .B1(_04324_),
    .A1(net3513),
    .Y(_04994_),
    .A2(net3512));
 sg13g2_or4_1 _10783_ (.A(net3508),
    .B(_00699_),
    .C(net3506),
    .D(net2851),
    .X(_04995_));
 sg13g2_a21oi_1 _10784_ (.A1(_04131_),
    .A2(_04207_),
    .Y(_04996_),
    .B1(_00680_));
 sg13g2_a21oi_1 _10785_ (.A1(\core.f2e_inst[25] ),
    .A2(net3345),
    .Y(_04997_),
    .B1(net3160));
 sg13g2_nand2b_1 _10786_ (.Y(_04998_),
    .B(_04995_),
    .A_N(_04711_));
 sg13g2_o21ai_1 _10787_ (.B1(_04997_),
    .Y(_04999_),
    .A1(_00159_),
    .A2(_04370_));
 sg13g2_nor4_2 _10788_ (.A(_04994_),
    .B(_04996_),
    .C(_04998_),
    .Y(_05000_),
    .D(_04999_));
 sg13g2_nor3_1 _10789_ (.A(net2745),
    .B(_04993_),
    .C(_05000_),
    .Y(_05001_));
 sg13g2_a21o_1 _10790_ (.A2(net2745),
    .A1(net3449),
    .B1(_05001_),
    .X(_00517_));
 sg13g2_nor2_1 _10791_ (.A(net3536),
    .B(net3450),
    .Y(_05002_));
 sg13g2_a22oi_1 _10792_ (.Y(_05003_),
    .B1(net3533),
    .B2(net3451),
    .A2(net3450),
    .A1(net3536));
 sg13g2_nor2_1 _10793_ (.A(_05002_),
    .B(_05003_),
    .Y(_05004_));
 sg13g2_a21oi_2 _10794_ (.B1(_05002_),
    .Y(_05005_),
    .A2(_05003_),
    .A1(_04932_));
 sg13g2_xnor2_1 _10795_ (.Y(_05006_),
    .A(_01260_),
    .B(_05005_));
 sg13g2_o21ai_1 _10796_ (.B1(_01264_),
    .Y(_05007_),
    .A1(_01262_),
    .A2(_04934_));
 sg13g2_nand3_1 _10797_ (.B(_01265_),
    .C(_05007_),
    .A(_01260_),
    .Y(_05008_));
 sg13g2_a21o_1 _10798_ (.A2(_05007_),
    .A1(_01265_),
    .B1(_01260_),
    .X(_05009_));
 sg13g2_nand3_1 _10799_ (.B(_05008_),
    .C(_05009_),
    .A(net2925),
    .Y(_05010_));
 sg13g2_nand3_1 _10800_ (.B(net3296),
    .C(net3053),
    .A(net3547),
    .Y(_05011_));
 sg13g2_nand2_1 _10801_ (.Y(_05012_),
    .A(net2956),
    .B(_05011_));
 sg13g2_o21ai_1 _10802_ (.B1(_05012_),
    .Y(_05013_),
    .A1(\core.work.alu.sval2[26] ),
    .A2(net2956));
 sg13g2_o21ai_1 _10803_ (.B1(net2854),
    .Y(_05014_),
    .A1(_00044_),
    .A2(_05013_));
 sg13g2_o21ai_1 _10804_ (.B1(net2942),
    .Y(_05015_),
    .A1(_00042_),
    .A2(net2952));
 sg13g2_a21oi_1 _10805_ (.A1(net2937),
    .A2(_05011_),
    .Y(_05016_),
    .B1(_05015_));
 sg13g2_a21oi_1 _10806_ (.A1(net2930),
    .A2(_05011_),
    .Y(_05017_),
    .B1(net2942));
 sg13g2_o21ai_1 _10807_ (.B1(_05017_),
    .Y(_05018_),
    .A1(\core.work.alu.sval2[26] ),
    .A2(net2930));
 sg13g2_o21ai_1 _10808_ (.B1(_00044_),
    .Y(_05019_),
    .A1(net2860),
    .A2(_05013_));
 sg13g2_inv_1 _10809_ (.Y(_05020_),
    .A(_05019_));
 sg13g2_a22oi_1 _10810_ (.Y(_05021_),
    .B1(_05018_),
    .B2(_05020_),
    .A2(_05016_),
    .A1(_05014_));
 sg13g2_nor2_1 _10811_ (.A(net2829),
    .B(_04941_),
    .Y(_05022_));
 sg13g2_nand2_1 _10812_ (.Y(_05023_),
    .A(_00048_),
    .B(net3055));
 sg13g2_nand2_1 _10813_ (.Y(_05024_),
    .A(_00049_),
    .B(net3061));
 sg13g2_nand2_1 _10814_ (.Y(_05025_),
    .A(_05023_),
    .B(_05024_));
 sg13g2_or2_1 _10815_ (.X(_05026_),
    .B(_04948_),
    .A(net2821));
 sg13g2_nand2_1 _10816_ (.Y(_05027_),
    .A(_04874_),
    .B(_04939_));
 sg13g2_o21ai_1 _10817_ (.B1(net2788),
    .Y(_05028_),
    .A1(net2833),
    .A2(_05027_));
 sg13g2_o21ai_1 _10818_ (.B1(_05026_),
    .Y(_05029_),
    .A1(net2825),
    .A2(_05025_));
 sg13g2_nor4_1 _10819_ (.A(_05021_),
    .B(_05022_),
    .C(_05028_),
    .D(_05029_),
    .Y(_05030_));
 sg13g2_a221oi_1 _10820_ (.B2(_05030_),
    .C1(net3298),
    .B1(_05010_),
    .A1(net2792),
    .Y(_05031_),
    .A2(_05006_));
 sg13g2_a21oi_1 _10821_ (.A1(_04131_),
    .A2(_04220_),
    .Y(_05032_),
    .B1(_04215_));
 sg13g2_o21ai_1 _10822_ (.B1(\core.f2e_inst[7] ),
    .Y(_05033_),
    .A1(_04215_),
    .A2(_04220_));
 sg13g2_a21o_1 _10823_ (.A2(_04216_),
    .A1(net3507),
    .B1(_04998_),
    .X(_05034_));
 sg13g2_nor2b_1 _10824_ (.A(_04212_),
    .B_N(net3511),
    .Y(_05035_));
 sg13g2_a21oi_1 _10825_ (.A1(\core.f2e_inst[2] ),
    .A2(_04446_),
    .Y(_05036_),
    .B1(net3348));
 sg13g2_o21ai_1 _10826_ (.B1(_05036_),
    .Y(_05037_),
    .A1(_00162_),
    .A2(_04370_));
 sg13g2_nor3_1 _10827_ (.A(_05034_),
    .B(_05035_),
    .C(_05037_),
    .Y(_05038_));
 sg13g2_o21ai_1 _10828_ (.B1(net3163),
    .Y(_05039_),
    .A1(\core.f2e_inst[26] ),
    .A2(net3337));
 sg13g2_a21oi_2 _10829_ (.B1(_05039_),
    .Y(_05040_),
    .A2(_05038_),
    .A1(_05033_));
 sg13g2_nand2_1 _10830_ (.Y(_05041_),
    .A(net2841),
    .B(_03837_));
 sg13g2_nor3_1 _10831_ (.A(net2746),
    .B(_05031_),
    .C(_05040_),
    .Y(_05042_));
 sg13g2_a22oi_1 _10832_ (.Y(_00518_),
    .B1(_05041_),
    .B2(_05042_),
    .A2(net2746),
    .A1(_00613_));
 sg13g2_nor2_1 _10833_ (.A(_00612_),
    .B(_00613_),
    .Y(_05043_));
 sg13g2_a21oi_1 _10834_ (.A1(_01260_),
    .A2(_05005_),
    .Y(_05044_),
    .B1(_05043_));
 sg13g2_xor2_1 _10835_ (.B(_05044_),
    .A(_01258_),
    .X(_05045_));
 sg13g2_nand2b_1 _10836_ (.Y(_05046_),
    .B(_05009_),
    .A_N(_01259_));
 sg13g2_xnor2_1 _10837_ (.Y(_05047_),
    .A(_01258_),
    .B(_05046_));
 sg13g2_nand3_1 _10838_ (.B(net3296),
    .C(net3292),
    .A(net3547),
    .Y(_05048_));
 sg13g2_nor2_1 _10839_ (.A(net3537),
    .B(net2956),
    .Y(_05049_));
 sg13g2_a21oi_1 _10840_ (.A1(net2956),
    .A2(_05048_),
    .Y(_05050_),
    .B1(_05049_));
 sg13g2_a21o_1 _10841_ (.A2(_05050_),
    .A1(_00645_),
    .B1(net2860),
    .X(_05051_));
 sg13g2_o21ai_1 _10842_ (.B1(net2942),
    .Y(_05052_),
    .A1(_00045_),
    .A2(net2952));
 sg13g2_a21oi_1 _10843_ (.A1(net2937),
    .A2(_05048_),
    .Y(_05053_),
    .B1(_05052_));
 sg13g2_o21ai_1 _10844_ (.B1(net2949),
    .Y(_05054_),
    .A1(net3537),
    .A2(net2930));
 sg13g2_a21oi_1 _10845_ (.A1(net2930),
    .A2(_05048_),
    .Y(_05055_),
    .B1(_05054_));
 sg13g2_a21oi_1 _10846_ (.A1(net2854),
    .A2(_05050_),
    .Y(_05056_),
    .B1(_05055_));
 sg13g2_a22oi_1 _10847_ (.Y(_05057_),
    .B1(_05056_),
    .B2(_00046_),
    .A2(_05053_),
    .A1(_05051_));
 sg13g2_o21ai_1 _10848_ (.B1(_04901_),
    .Y(_05058_),
    .A1(_00645_),
    .A2(net3061));
 sg13g2_nor2_1 _10849_ (.A(_00052_),
    .B(net3055),
    .Y(_05059_));
 sg13g2_nor2_1 _10850_ (.A(_00049_),
    .B(net3061),
    .Y(_05060_));
 sg13g2_o21ai_1 _10851_ (.B1(_04015_),
    .Y(_05061_),
    .A1(_05059_),
    .A2(_05060_));
 sg13g2_o21ai_1 _10852_ (.B1(_05061_),
    .Y(_05062_),
    .A1(net2833),
    .A2(_05058_));
 sg13g2_o21ai_1 _10853_ (.B1(_04010_),
    .Y(_05063_),
    .A1(_04978_),
    .A2(_04979_));
 sg13g2_o21ai_1 _10854_ (.B1(_05063_),
    .Y(_05064_),
    .A1(net2821),
    .A2(_04981_));
 sg13g2_or4_1 _10855_ (.A(net2792),
    .B(_05057_),
    .C(_05062_),
    .D(_05064_),
    .X(_05065_));
 sg13g2_a21oi_1 _10856_ (.A1(net2925),
    .A2(_05047_),
    .Y(_05066_),
    .B1(_05065_));
 sg13g2_a21oi_2 _10857_ (.B1(_05066_),
    .Y(_05067_),
    .A2(_05045_),
    .A1(net2792));
 sg13g2_a221oi_1 _10858_ (.B2(net3303),
    .C1(net3164),
    .B1(_05067_),
    .A1(net2841),
    .Y(_05068_),
    .A2(_03859_));
 sg13g2_nor3_1 _10859_ (.A(_00695_),
    .B(net3345),
    .C(_05032_),
    .Y(_05069_));
 sg13g2_and2_1 _10860_ (.A(net3510),
    .B(_04293_),
    .X(_05070_));
 sg13g2_a221oi_1 _10861_ (.B2(\core.f2e_inst[3] ),
    .C1(net3160),
    .B1(_04446_),
    .A1(\core.f2e_inst[27] ),
    .Y(_05071_),
    .A2(net3345));
 sg13g2_o21ai_1 _10862_ (.B1(_05071_),
    .Y(_05072_),
    .A1(_00160_),
    .A2(_04370_));
 sg13g2_nor4_1 _10863_ (.A(_05034_),
    .B(_05069_),
    .C(_05070_),
    .D(_05072_),
    .Y(_05073_));
 sg13g2_or2_1 _10864_ (.X(_05074_),
    .B(_05073_),
    .A(net2742));
 sg13g2_nand2_1 _10865_ (.Y(_05075_),
    .A(net3448),
    .B(net2744));
 sg13g2_o21ai_1 _10866_ (.B1(_05075_),
    .Y(_00519_),
    .A1(_05068_),
    .A2(_05074_));
 sg13g2_and2_1 _10867_ (.A(_01258_),
    .B(_01260_),
    .X(_05076_));
 sg13g2_nand4_1 _10868_ (.B(_01266_),
    .C(_04931_),
    .A(_01263_),
    .Y(_05077_),
    .D(_05076_));
 sg13g2_nand2_1 _10869_ (.Y(_05078_),
    .A(net3537),
    .B(net3448));
 sg13g2_o21ai_1 _10870_ (.B1(_05043_),
    .Y(_05079_),
    .A1(\core.work.alu.sval2[27] ),
    .A2(net3448));
 sg13g2_nand3_1 _10871_ (.B(_01260_),
    .C(_05004_),
    .A(_01258_),
    .Y(_05080_));
 sg13g2_nand4_1 _10872_ (.B(_05078_),
    .C(_05079_),
    .A(_05077_),
    .Y(_05081_),
    .D(_05080_));
 sg13g2_nand2_1 _10873_ (.Y(_05082_),
    .A(_01283_),
    .B(_05081_));
 sg13g2_xnor2_1 _10874_ (.Y(_05083_),
    .A(_01284_),
    .B(_05081_));
 sg13g2_xnor2_1 _10875_ (.Y(_05084_),
    .A(_01272_),
    .B(_01283_));
 sg13g2_nor2_1 _10876_ (.A(net2829),
    .B(_05025_),
    .Y(_05085_));
 sg13g2_nor2_1 _10877_ (.A(net2821),
    .B(_05027_),
    .Y(_05086_));
 sg13g2_nor2_1 _10878_ (.A(_05085_),
    .B(_05086_),
    .Y(_05087_));
 sg13g2_nand2_1 _10879_ (.Y(_05088_),
    .A(_04940_),
    .B(_05023_));
 sg13g2_nand2_1 _10880_ (.Y(_05089_),
    .A(net3547),
    .B(_04497_));
 sg13g2_o21ai_1 _10881_ (.B1(net2942),
    .Y(_05090_),
    .A1(_00047_),
    .A2(net2952));
 sg13g2_a21oi_1 _10882_ (.A1(net2937),
    .A2(_05089_),
    .Y(_05091_),
    .B1(_05090_));
 sg13g2_nand2_1 _10883_ (.Y(_05092_),
    .A(_00052_),
    .B(net3055));
 sg13g2_nand2_1 _10884_ (.Y(_05093_),
    .A(_00024_),
    .B(net3062));
 sg13g2_nand3_1 _10885_ (.B(_05092_),
    .C(_05093_),
    .A(_04015_),
    .Y(_05094_));
 sg13g2_o21ai_1 _10886_ (.B1(net2949),
    .Y(_05095_),
    .A1(\core.work.alu.sval2[28] ),
    .A2(net2930));
 sg13g2_a21oi_1 _10887_ (.A1(net2930),
    .A2(_05089_),
    .Y(_05096_),
    .B1(_05095_));
 sg13g2_o21ai_1 _10888_ (.B1(_05087_),
    .Y(_05097_),
    .A1(_00048_),
    .A2(_05091_));
 sg13g2_o21ai_1 _10889_ (.B1(_05094_),
    .Y(_05098_),
    .A1(net2833),
    .A2(_05088_));
 sg13g2_nor4_1 _10890_ (.A(net2792),
    .B(_05096_),
    .C(_05097_),
    .D(_05098_),
    .Y(_05099_));
 sg13g2_nor2_1 _10891_ (.A(\core.work.alu.sval2[28] ),
    .B(net2956),
    .Y(_05100_));
 sg13g2_a21oi_1 _10892_ (.A1(net2956),
    .A2(_05089_),
    .Y(_05101_),
    .B1(_05100_));
 sg13g2_xnor2_1 _10893_ (.Y(_05102_),
    .A(_00048_),
    .B(_05101_));
 sg13g2_a22oi_1 _10894_ (.Y(_05103_),
    .B1(_05102_),
    .B2(net2854),
    .A2(_05084_),
    .A1(net2925));
 sg13g2_a21oi_1 _10895_ (.A1(_05099_),
    .A2(_05103_),
    .Y(_05104_),
    .B1(net3297));
 sg13g2_o21ai_1 _10896_ (.B1(_05104_),
    .Y(_05105_),
    .A1(net2788),
    .A2(_05083_));
 sg13g2_a21oi_1 _10897_ (.A1(net2841),
    .A2(_03884_),
    .Y(_05106_),
    .B1(net3163));
 sg13g2_nand3_1 _10898_ (.B(net3336),
    .C(_04220_),
    .A(net897),
    .Y(_05107_));
 sg13g2_o21ai_1 _10899_ (.B1(net3507),
    .Y(_05108_),
    .A1(_04206_),
    .A2(_04216_));
 sg13g2_nand2_1 _10900_ (.Y(_05109_),
    .A(_04995_),
    .B(_05108_));
 sg13g2_nand2_1 _10901_ (.Y(_05110_),
    .A(\core.f2e_inst[28] ),
    .B(net3342));
 sg13g2_o21ai_1 _10902_ (.B1(_05110_),
    .Y(_05111_),
    .A1(_00161_),
    .A2(_04370_));
 sg13g2_nor3_1 _10903_ (.A(_04887_),
    .B(_05109_),
    .C(_05111_),
    .Y(_05112_));
 sg13g2_a221oi_1 _10904_ (.B2(_05112_),
    .C1(net2742),
    .B1(_05107_),
    .A1(_05105_),
    .Y(_05113_),
    .A2(_05106_));
 sg13g2_a21o_1 _10905_ (.A2(net2742),
    .A1(net3447),
    .B1(_05113_),
    .X(_00520_));
 sg13g2_nand2_1 _10906_ (.Y(_05114_),
    .A(_01282_),
    .B(_05082_));
 sg13g2_xnor2_1 _10907_ (.Y(_05115_),
    .A(_01280_),
    .B(_05114_));
 sg13g2_nand2_1 _10908_ (.Y(_05116_),
    .A(_01286_),
    .B(_01291_));
 sg13g2_xnor2_1 _10909_ (.Y(_05117_),
    .A(_01281_),
    .B(_05116_));
 sg13g2_nand2_1 _10910_ (.Y(_05118_),
    .A(net2925),
    .B(_05117_));
 sg13g2_nor2_1 _10911_ (.A(net3540),
    .B(net2958),
    .Y(_05119_));
 sg13g2_nand2_1 _10912_ (.Y(_05120_),
    .A(net3547),
    .B(_04543_));
 sg13g2_a21oi_1 _10913_ (.A1(net2958),
    .A2(_05120_),
    .Y(_05121_),
    .B1(_05119_));
 sg13g2_xnor2_1 _10914_ (.Y(_05122_),
    .A(_00049_),
    .B(_05121_));
 sg13g2_nor3_1 _10915_ (.A(net2853),
    .B(_05059_),
    .C(_05060_),
    .Y(_05123_));
 sg13g2_nor4_1 _10916_ (.A(_00024_),
    .B(_01309_),
    .C(_01719_),
    .D(net3063),
    .Y(_05124_));
 sg13g2_o21ai_1 _10917_ (.B1(net2830),
    .Y(_05125_),
    .A1(_00024_),
    .A2(_01721_));
 sg13g2_nor2_1 _10918_ (.A(_05124_),
    .B(_05125_),
    .Y(_05126_));
 sg13g2_o21ai_1 _10919_ (.B1(net2949),
    .Y(_05127_),
    .A1(net3540),
    .A2(net2931));
 sg13g2_a21oi_1 _10920_ (.A1(net2931),
    .A2(_05120_),
    .Y(_05128_),
    .B1(_05127_));
 sg13g2_nor2_1 _10921_ (.A(_04978_),
    .B(_05060_),
    .Y(_05129_));
 sg13g2_nor2_1 _10922_ (.A(net2833),
    .B(_05129_),
    .Y(_05130_));
 sg13g2_nor2_1 _10923_ (.A(net2821),
    .B(_05058_),
    .Y(_05131_));
 sg13g2_o21ai_1 _10924_ (.B1(net2942),
    .Y(_05132_),
    .A1(_00051_),
    .A2(net2952));
 sg13g2_a21oi_1 _10925_ (.A1(net2937),
    .A2(_05120_),
    .Y(_05133_),
    .B1(_05132_));
 sg13g2_o21ai_1 _10926_ (.B1(net2788),
    .Y(_05134_),
    .A1(_00049_),
    .A2(_05133_));
 sg13g2_nor4_1 _10927_ (.A(_05128_),
    .B(_05130_),
    .C(_05131_),
    .D(_05134_),
    .Y(_05135_));
 sg13g2_o21ai_1 _10928_ (.B1(_05135_),
    .Y(_05136_),
    .A1(_05123_),
    .A2(_05126_));
 sg13g2_a21oi_1 _10929_ (.A1(net2854),
    .A2(_05122_),
    .Y(_05137_),
    .B1(_05136_));
 sg13g2_a21oi_1 _10930_ (.A1(_05118_),
    .A2(_05137_),
    .Y(_05138_),
    .B1(net3297));
 sg13g2_o21ai_1 _10931_ (.B1(_05138_),
    .Y(_05139_),
    .A1(net2788),
    .A2(_05115_));
 sg13g2_nand2_1 _10932_ (.Y(_05140_),
    .A(net2841),
    .B(_03905_));
 sg13g2_or2_1 _10933_ (.X(_05141_),
    .B(_05109_),
    .A(_04710_));
 sg13g2_nor2_1 _10934_ (.A(net3346),
    .B(_05141_),
    .Y(_05142_));
 sg13g2_a221oi_1 _10935_ (.B2(_04220_),
    .C1(_05141_),
    .B1(net3509),
    .A1(net3513),
    .Y(_05143_),
    .A2(net3512));
 sg13g2_o21ai_1 _10936_ (.B1(net3162),
    .Y(_05144_),
    .A1(\core.f2e_inst[29] ),
    .A2(net3335));
 sg13g2_o21ai_1 _10937_ (.B1(_05140_),
    .Y(_05145_),
    .A1(_05143_),
    .A2(_05144_));
 sg13g2_nor2_1 _10938_ (.A(net2743),
    .B(_05145_),
    .Y(_05146_));
 sg13g2_a22oi_1 _10939_ (.Y(_00521_),
    .B1(_05139_),
    .B2(_05146_),
    .A2(net2745),
    .A1(_00609_));
 sg13g2_nor2_1 _10940_ (.A(_01280_),
    .B(_01284_),
    .Y(_05147_));
 sg13g2_a21oi_1 _10941_ (.A1(_00608_),
    .A2(_00609_),
    .Y(_05148_),
    .B1(_01282_));
 sg13g2_a221oi_1 _10942_ (.B2(_05147_),
    .C1(_05148_),
    .B1(_05081_),
    .A1(\core.work.alu.sval2[29] ),
    .Y(_05149_),
    .A2(net3445));
 sg13g2_xnor2_1 _10943_ (.Y(_05150_),
    .A(_01275_),
    .B(_05149_));
 sg13g2_xnor2_1 _10944_ (.Y(_05151_),
    .A(_01275_),
    .B(_01293_));
 sg13g2_nor2_1 _10945_ (.A(\core.work.alu.sval2[30] ),
    .B(net2957),
    .Y(_05152_));
 sg13g2_nand2_1 _10946_ (.Y(_05153_),
    .A(net3547),
    .B(_04577_));
 sg13g2_a21oi_1 _10947_ (.A1(net2957),
    .A2(_05153_),
    .Y(_05154_),
    .B1(_05152_));
 sg13g2_nand2b_1 _10948_ (.Y(_05155_),
    .B(_00052_),
    .A_N(_05154_));
 sg13g2_a21oi_1 _10949_ (.A1(_00648_),
    .A2(_05154_),
    .Y(_05156_),
    .B1(net2860));
 sg13g2_a21oi_1 _10950_ (.A1(\core.work.alu.sval2[30] ),
    .A2(net2928),
    .Y(_05157_),
    .B1(_00648_));
 sg13g2_o21ai_1 _10951_ (.B1(_05157_),
    .Y(_05158_),
    .A1(net2928),
    .A2(_05153_));
 sg13g2_nand2_1 _10952_ (.Y(_05159_),
    .A(net2937),
    .B(_05153_));
 sg13g2_o21ai_1 _10953_ (.B1(_05159_),
    .Y(_05160_),
    .A1(_00050_),
    .A2(net2953));
 sg13g2_a22oi_1 _10954_ (.Y(_05161_),
    .B1(_05160_),
    .B2(_00648_),
    .A2(_05158_),
    .A1(net2949));
 sg13g2_a21o_1 _10955_ (.A2(_05093_),
    .A1(_05092_),
    .B1(net2853),
    .X(_05162_));
 sg13g2_and2_1 _10956_ (.A(_03990_),
    .B(_05024_),
    .X(_05163_));
 sg13g2_a221oi_1 _10957_ (.B2(_05092_),
    .C1(net2792),
    .B1(_05163_),
    .A1(_05125_),
    .Y(_05164_),
    .A2(_05162_));
 sg13g2_o21ai_1 _10958_ (.B1(_05161_),
    .Y(_05165_),
    .A1(net2821),
    .A2(_05088_));
 sg13g2_a221oi_1 _10959_ (.B2(_05156_),
    .C1(_05165_),
    .B1(_05155_),
    .A1(net2925),
    .Y(_05166_),
    .A2(_05151_));
 sg13g2_a22oi_1 _10960_ (.Y(_05167_),
    .B1(_05164_),
    .B2(_05166_),
    .A2(_05150_),
    .A1(net2792));
 sg13g2_nand2_1 _10961_ (.Y(_05168_),
    .A(net3303),
    .B(_05167_));
 sg13g2_o21ai_1 _10962_ (.B1(_04960_),
    .Y(_05169_),
    .A1(_00695_),
    .A2(_04131_));
 sg13g2_a21oi_1 _10963_ (.A1(_04204_),
    .A2(_04602_),
    .Y(_05170_),
    .B1(_05169_));
 sg13g2_a22oi_1 _10964_ (.Y(_05171_),
    .B1(_05142_),
    .B2(_05170_),
    .A2(net3346),
    .A1(_00703_));
 sg13g2_a221oi_1 _10965_ (.B2(net3162),
    .C1(net2743),
    .B1(_05171_),
    .A1(net2841),
    .Y(_05172_),
    .A2(_03928_));
 sg13g2_a22oi_1 _10966_ (.Y(_00522_),
    .B1(_05168_),
    .B2(_05172_),
    .A2(net2746),
    .A1(_00607_));
 sg13g2_nand2_1 _10967_ (.Y(_05173_),
    .A(\core.work.alu.sval2[30] ),
    .B(net3444));
 sg13g2_o21ai_1 _10968_ (.B1(_05173_),
    .Y(_05174_),
    .A1(_01275_),
    .A2(_05149_));
 sg13g2_xor2_1 _10969_ (.B(_05174_),
    .A(_01273_),
    .X(_05175_));
 sg13g2_nand2_1 _10970_ (.Y(_05176_),
    .A(net3547),
    .B(_04617_));
 sg13g2_nand2_1 _10971_ (.Y(_05177_),
    .A(net2957),
    .B(_05176_));
 sg13g2_o21ai_1 _10972_ (.B1(_05177_),
    .Y(_05178_),
    .A1(\core.work.alu.sval2[31] ),
    .A2(net2957));
 sg13g2_xnor2_1 _10973_ (.Y(_05179_),
    .A(net3361),
    .B(_05178_));
 sg13g2_a21o_1 _10974_ (.A2(net3056),
    .A1(net3361),
    .B1(_05059_),
    .X(_05180_));
 sg13g2_a22oi_1 _10975_ (.Y(_05181_),
    .B1(net2941),
    .B2(_05176_),
    .A2(_01720_),
    .A1(_01308_));
 sg13g2_o21ai_1 _10976_ (.B1(_05181_),
    .Y(_05182_),
    .A1(_00053_),
    .A2(net2952));
 sg13g2_a21oi_1 _10977_ (.A1(\core.work.alu.sval2[31] ),
    .A2(net2928),
    .Y(_05183_),
    .B1(net3361));
 sg13g2_o21ai_1 _10978_ (.B1(_05183_),
    .Y(_05184_),
    .A1(net2928),
    .A2(_05176_));
 sg13g2_a22oi_1 _10979_ (.Y(_05185_),
    .B1(_05184_),
    .B2(net2949),
    .A2(_05180_),
    .A1(_03990_));
 sg13g2_a221oi_1 _10980_ (.B2(net3361),
    .C1(_04005_),
    .B1(_05182_),
    .A1(_03988_),
    .Y(_05186_),
    .A2(_05124_));
 sg13g2_o21ai_1 _10981_ (.B1(_05185_),
    .Y(_05187_),
    .A1(net2821),
    .A2(_05129_));
 sg13g2_xnor2_1 _10982_ (.Y(_05188_),
    .A(_01273_),
    .B(_01294_));
 sg13g2_a221oi_1 _10983_ (.B2(net2925),
    .C1(_05187_),
    .B1(_05188_),
    .A1(net2854),
    .Y(_05189_),
    .A2(_05179_));
 sg13g2_a21oi_1 _10984_ (.A1(_05186_),
    .A2(_05189_),
    .Y(_05190_),
    .B1(net3298));
 sg13g2_o21ai_1 _10985_ (.B1(_05190_),
    .Y(_05191_),
    .A1(net2788),
    .A2(_05175_));
 sg13g2_nor2_1 _10986_ (.A(_04519_),
    .B(_05141_),
    .Y(_05192_));
 sg13g2_a21oi_1 _10987_ (.A1(_00706_),
    .A2(net3348),
    .Y(_05193_),
    .B1(_05192_));
 sg13g2_a221oi_1 _10988_ (.B2(net3162),
    .C1(net2743),
    .B1(_05193_),
    .A1(net2841),
    .Y(_05194_),
    .A2(_03949_));
 sg13g2_a22oi_1 _10989_ (.Y(_00523_),
    .B1(_05191_),
    .B2(_05194_),
    .A2(net2742),
    .A1(_00605_));
 sg13g2_and2_1 _10990_ (.A(_00055_),
    .B(net3305),
    .X(_05195_));
 sg13g2_o21ai_1 _10991_ (.B1(_03183_),
    .Y(_05196_),
    .A1(net2787),
    .A2(_05195_));
 sg13g2_nor2_1 _10992_ (.A(net3480),
    .B(net2922),
    .Y(_05197_));
 sg13g2_a22oi_1 _10993_ (.Y(_05198_),
    .B1(_02565_),
    .B2(_05197_),
    .A2(net2922),
    .A1(_00124_));
 sg13g2_nor2_1 _10994_ (.A(net2922),
    .B(_02565_),
    .Y(_05199_));
 sg13g2_nand2b_1 _10995_ (.Y(_05200_),
    .B(net3482),
    .A_N(_05198_));
 sg13g2_nor2_2 _10996_ (.A(net3483),
    .B(net3484),
    .Y(_05201_));
 sg13g2_nand2_1 _10997_ (.Y(_05202_),
    .A(net3480),
    .B(_05201_));
 sg13g2_o21ai_1 _10998_ (.B1(_05200_),
    .Y(_05203_),
    .A1(_05199_),
    .A2(_05202_));
 sg13g2_nor2_1 _10999_ (.A(net3482),
    .B(_00601_),
    .Y(_05204_));
 sg13g2_nand2b_1 _11000_ (.Y(_05205_),
    .B(net3484),
    .A_N(net3482));
 sg13g2_a22oi_1 _11001_ (.Y(_05206_),
    .B1(_05204_),
    .B2(net3480),
    .A2(_05201_),
    .A1(_05197_));
 sg13g2_nor3_1 _11002_ (.A(_00600_),
    .B(_02564_),
    .C(_05205_),
    .Y(_05207_));
 sg13g2_nor2_1 _11003_ (.A(_02564_),
    .B(_05206_),
    .Y(_05208_));
 sg13g2_nand4_1 _11004_ (.B(net3448),
    .C(\core.e2m_addr[26] ),
    .A(net3480),
    .Y(_05209_),
    .D(net3449));
 sg13g2_nor3_1 _11005_ (.A(net2922),
    .B(_02561_),
    .C(_05209_),
    .Y(_05210_));
 sg13g2_nand2_1 _11006_ (.Y(_05211_),
    .A(net3484),
    .B(_05210_));
 sg13g2_o21ai_1 _11007_ (.B1(_05211_),
    .Y(_05212_),
    .A1(_01993_),
    .A2(_05199_));
 sg13g2_nand3_1 _11008_ (.B(net2922),
    .C(_05201_),
    .A(_00124_),
    .Y(_05213_));
 sg13g2_nor3_1 _11009_ (.A(net3480),
    .B(_00609_),
    .C(net3447),
    .Y(_05214_));
 sg13g2_nand2_1 _11010_ (.Y(_05215_),
    .A(_00605_),
    .B(_05204_));
 sg13g2_nor4_1 _11011_ (.A(_00611_),
    .B(\core.e2m_addr[26] ),
    .C(net3449),
    .D(_05215_),
    .Y(_05216_));
 sg13g2_nand3_1 _11012_ (.B(_02559_),
    .C(_05216_),
    .A(net3444),
    .Y(_05217_));
 sg13g2_nand2_1 _11013_ (.Y(_05218_),
    .A(_05214_),
    .B(_05216_));
 sg13g2_inv_1 _11014_ (.Y(_05219_),
    .A(_05218_));
 sg13g2_nand2_1 _11015_ (.Y(_05220_),
    .A(_05217_),
    .B(_05218_));
 sg13g2_nand3_1 _11016_ (.B(_05217_),
    .C(_05218_),
    .A(_05213_),
    .Y(_05221_));
 sg13g2_nor4_2 _11017_ (.A(_05203_),
    .B(_05208_),
    .C(_05212_),
    .Y(_05222_),
    .D(_05221_));
 sg13g2_or2_1 _11018_ (.X(_05223_),
    .B(_05217_),
    .A(_00600_));
 sg13g2_nand2_1 _11019_ (.Y(_05224_),
    .A(_00607_),
    .B(_05219_));
 sg13g2_o21ai_1 _11020_ (.B1(_00601_),
    .Y(_05225_),
    .A1(_01993_),
    .A2(_05199_));
 sg13g2_a21oi_1 _11021_ (.A1(net3482),
    .A2(_05210_),
    .Y(_05226_),
    .B1(_00601_));
 sg13g2_nand2_1 _11022_ (.Y(_05227_),
    .A(_05200_),
    .B(_05226_));
 sg13g2_nand2_1 _11023_ (.Y(_05228_),
    .A(_05225_),
    .B(_05227_));
 sg13g2_nand4_1 _11024_ (.B(_05223_),
    .C(_05224_),
    .A(net3031),
    .Y(_05229_),
    .D(_05228_));
 sg13g2_a21o_1 _11025_ (.A2(_05208_),
    .A1(net3444),
    .B1(_05229_),
    .X(_05230_));
 sg13g2_nor2_1 _11026_ (.A(net3484),
    .B(net3034),
    .Y(_05231_));
 sg13g2_o21ai_1 _11027_ (.B1(_01686_),
    .Y(_05232_),
    .A1(net3038),
    .A2(_05201_));
 sg13g2_o21ai_1 _11028_ (.B1(net3195),
    .Y(_05233_),
    .A1(_05231_),
    .A2(_05232_));
 sg13g2_o21ai_1 _11029_ (.B1(_05233_),
    .Y(_05234_),
    .A1(_05222_),
    .A2(_05230_));
 sg13g2_nor4_1 _11030_ (.A(net3305),
    .B(net3029),
    .C(_05196_),
    .D(_05234_),
    .Y(_05235_));
 sg13g2_a21o_1 _11031_ (.A2(_05196_),
    .A1(net840),
    .B1(_05235_),
    .X(_00524_));
 sg13g2_o21ai_1 _11032_ (.B1(net3031),
    .Y(_05236_),
    .A1(net3484),
    .A2(_05200_));
 sg13g2_nor4_1 _11033_ (.A(_05212_),
    .B(_05219_),
    .C(_05222_),
    .D(_05236_),
    .Y(_05237_));
 sg13g2_nand2_1 _11034_ (.Y(_05238_),
    .A(net3482),
    .B(_01686_));
 sg13g2_a22oi_1 _11035_ (.Y(_05239_),
    .B1(_05238_),
    .B2(net2903),
    .A2(_05205_),
    .A1(net3034));
 sg13g2_nor3_1 _11036_ (.A(net3305),
    .B(net3029),
    .C(_05237_),
    .Y(_05240_));
 sg13g2_o21ai_1 _11037_ (.B1(_05240_),
    .Y(_05241_),
    .A1(net3031),
    .A2(_05239_));
 sg13g2_nand2_1 _11038_ (.Y(_05242_),
    .A(net3441),
    .B(_05196_));
 sg13g2_o21ai_1 _11039_ (.B1(_05242_),
    .Y(_00525_),
    .A1(_05196_),
    .A2(_05241_));
 sg13g2_nor4_1 _11040_ (.A(_01670_),
    .B(_05203_),
    .C(_05220_),
    .D(_05222_),
    .Y(_05243_));
 sg13g2_a21oi_1 _11041_ (.A1(net3481),
    .A2(net3038),
    .Y(_05244_),
    .B1(net3031));
 sg13g2_o21ai_1 _11042_ (.B1(_05244_),
    .Y(_05245_),
    .A1(net3481),
    .A2(net2903));
 sg13g2_nor3_1 _11043_ (.A(net3305),
    .B(net3029),
    .C(_05243_),
    .Y(_05246_));
 sg13g2_a21oi_1 _11044_ (.A1(_05245_),
    .A2(_05246_),
    .Y(_05247_),
    .B1(_05196_));
 sg13g2_a21oi_1 _11045_ (.A1(_00629_),
    .A2(_05196_),
    .Y(_00526_),
    .B1(_05247_));
 sg13g2_nor3_1 _11046_ (.A(_01670_),
    .B(_05207_),
    .C(_05220_),
    .Y(_05248_));
 sg13g2_and2_1 _11047_ (.A(_05211_),
    .B(_05248_),
    .X(_05249_));
 sg13g2_nor4_1 _11048_ (.A(_01684_),
    .B(net3305),
    .C(_05196_),
    .D(_05249_),
    .Y(_05250_));
 sg13g2_a21o_1 _11049_ (.A2(_05196_),
    .A1(net3440),
    .B1(_05250_),
    .X(_00527_));
 sg13g2_nor3_1 _11050_ (.A(_00580_),
    .B(net3528),
    .C(net3529),
    .Y(_05251_));
 sg13g2_nand2_1 _11051_ (.Y(_05252_),
    .A(net3570),
    .B(net3052));
 sg13g2_o21ai_1 _11052_ (.B1(_05252_),
    .Y(_05253_),
    .A1(_00676_),
    .A2(net3052));
 sg13g2_nand3_1 _11053_ (.B(net2715),
    .C(_05253_),
    .A(net2880),
    .Y(_05254_));
 sg13g2_o21ai_1 _11054_ (.B1(_05254_),
    .Y(_00528_),
    .A1(_00676_),
    .A2(net2714));
 sg13g2_nand2_1 _11055_ (.Y(_05255_),
    .A(net3569),
    .B(net3052));
 sg13g2_o21ai_1 _11056_ (.B1(_05255_),
    .Y(_05256_),
    .A1(_00677_),
    .A2(net3052));
 sg13g2_nand3_1 _11057_ (.B(net2715),
    .C(_05256_),
    .A(net2880),
    .Y(_05257_));
 sg13g2_o21ai_1 _11058_ (.B1(_05257_),
    .Y(_00529_),
    .A1(_00677_),
    .A2(net2714));
 sg13g2_nand2_1 _11059_ (.Y(_05258_),
    .A(\core.fetch.cmd_data[2] ),
    .B(net3051));
 sg13g2_o21ai_1 _11060_ (.B1(_05258_),
    .Y(_05259_),
    .A1(_00679_),
    .A2(net3051));
 sg13g2_nand3_1 _11061_ (.B(net2720),
    .C(_05259_),
    .A(net2883),
    .Y(_05260_));
 sg13g2_o21ai_1 _11062_ (.B1(_05260_),
    .Y(_00530_),
    .A1(_00679_),
    .A2(net2720));
 sg13g2_nand2_1 _11063_ (.Y(_05261_),
    .A(\core.fetch.cmd_data[3] ),
    .B(net3052));
 sg13g2_o21ai_1 _11064_ (.B1(_05261_),
    .Y(_05262_),
    .A1(_00682_),
    .A2(net3052));
 sg13g2_nand3_1 _11065_ (.B(net2719),
    .C(_05262_),
    .A(net2883),
    .Y(_05263_));
 sg13g2_o21ai_1 _11066_ (.B1(_05263_),
    .Y(_00531_),
    .A1(_00682_),
    .A2(net2719));
 sg13g2_nand2_1 _11067_ (.Y(_05264_),
    .A(\core.fetch.cmd_data[4] ),
    .B(net3052));
 sg13g2_o21ai_1 _11068_ (.B1(_05264_),
    .Y(_05265_),
    .A1(_00685_),
    .A2(_05251_));
 sg13g2_nand3_1 _11069_ (.B(net2727),
    .C(_05265_),
    .A(net2887),
    .Y(_05266_));
 sg13g2_o21ai_1 _11070_ (.B1(_05266_),
    .Y(_00532_),
    .A1(_00685_),
    .A2(net2727));
 sg13g2_nand2_1 _11071_ (.Y(_05267_),
    .A(\core.fetch.cmd_data[5] ),
    .B(net3051));
 sg13g2_o21ai_1 _11072_ (.B1(_05267_),
    .Y(_05268_),
    .A1(_00688_),
    .A2(net3051));
 sg13g2_nand3_1 _11073_ (.B(net2721),
    .C(_05268_),
    .A(net2883),
    .Y(_05269_));
 sg13g2_o21ai_1 _11074_ (.B1(_05269_),
    .Y(_00533_),
    .A1(_00688_),
    .A2(net2722));
 sg13g2_nand2_1 _11075_ (.Y(_05270_),
    .A(\core.fetch.cmd_data[6] ),
    .B(net3051));
 sg13g2_o21ai_1 _11076_ (.B1(net566),
    .Y(_05271_),
    .A1(_00690_),
    .A2(net3051));
 sg13g2_nand3_1 _11077_ (.B(net2722),
    .C(_05271_),
    .A(net2885),
    .Y(_05272_));
 sg13g2_o21ai_1 _11078_ (.B1(_05272_),
    .Y(_00534_),
    .A1(_00690_),
    .A2(net2722));
 sg13g2_nand2_1 _11079_ (.Y(_05273_),
    .A(net607),
    .B(net3051));
 sg13g2_o21ai_1 _11080_ (.B1(_05273_),
    .Y(_05274_),
    .A1(_00692_),
    .A2(net3051));
 sg13g2_nand3_1 _11081_ (.B(net2720),
    .C(_05274_),
    .A(net2884),
    .Y(_05275_));
 sg13g2_o21ai_1 _11082_ (.B1(_05275_),
    .Y(_00535_),
    .A1(_00692_),
    .A2(net2720));
 sg13g2_nand3_1 _11083_ (.B(_00581_),
    .C(net3529),
    .A(net3527),
    .Y(_05276_));
 sg13g2_nor2_1 _11084_ (.A(net3570),
    .B(net3048),
    .Y(_05277_));
 sg13g2_a21oi_1 _11085_ (.A1(_00694_),
    .A2(net3048),
    .Y(_05278_),
    .B1(_05277_));
 sg13g2_nand3_1 _11086_ (.B(net2717),
    .C(_05278_),
    .A(net2882),
    .Y(_05279_));
 sg13g2_o21ai_1 _11087_ (.B1(_05279_),
    .Y(_00536_),
    .A1(_00694_),
    .A2(net2717));
 sg13g2_nor2_1 _11088_ (.A(net3569),
    .B(net3048),
    .Y(_05280_));
 sg13g2_a21oi_1 _11089_ (.A1(_00696_),
    .A2(net3048),
    .Y(_05281_),
    .B1(_05280_));
 sg13g2_nand3_1 _11090_ (.B(net2714),
    .C(_05281_),
    .A(net2880),
    .Y(_05282_));
 sg13g2_o21ai_1 _11091_ (.B1(_05282_),
    .Y(_00537_),
    .A1(_00696_),
    .A2(net2714));
 sg13g2_nor2_1 _11092_ (.A(\core.fetch.cmd_data[2] ),
    .B(net3050),
    .Y(_05283_));
 sg13g2_a21oi_1 _11093_ (.A1(_00697_),
    .A2(net3050),
    .Y(_05284_),
    .B1(_05283_));
 sg13g2_nand3_1 _11094_ (.B(net2729),
    .C(_05284_),
    .A(net2886),
    .Y(_05285_));
 sg13g2_o21ai_1 _11095_ (.B1(_05285_),
    .Y(_00538_),
    .A1(_00697_),
    .A2(net2729));
 sg13g2_nor2_1 _11096_ (.A(\core.fetch.cmd_data[3] ),
    .B(net3048),
    .Y(_05286_));
 sg13g2_a21oi_1 _11097_ (.A1(_00698_),
    .A2(net3048),
    .Y(_05287_),
    .B1(_05286_));
 sg13g2_nand3_1 _11098_ (.B(net2718),
    .C(_05287_),
    .A(net2881),
    .Y(_05288_));
 sg13g2_o21ai_1 _11099_ (.B1(_05288_),
    .Y(_00539_),
    .A1(_00698_),
    .A2(net2716));
 sg13g2_nor2_1 _11100_ (.A(\core.fetch.cmd_data[4] ),
    .B(net3049),
    .Y(_05289_));
 sg13g2_a21oi_1 _11101_ (.A1(_00700_),
    .A2(net3049),
    .Y(_05290_),
    .B1(_05289_));
 sg13g2_nand3_1 _11102_ (.B(net2721),
    .C(_05290_),
    .A(net2884),
    .Y(_05291_));
 sg13g2_o21ai_1 _11103_ (.B1(_05291_),
    .Y(_00540_),
    .A1(_00700_),
    .A2(net2721));
 sg13g2_nor2_1 _11104_ (.A(\core.fetch.cmd_data[5] ),
    .B(net3048),
    .Y(_05292_));
 sg13g2_a21oi_1 _11105_ (.A1(_00702_),
    .A2(net3048),
    .Y(_05293_),
    .B1(_05292_));
 sg13g2_nand3_1 _11106_ (.B(net2716),
    .C(_05293_),
    .A(net2881),
    .Y(_05294_));
 sg13g2_o21ai_1 _11107_ (.B1(_05294_),
    .Y(_00541_),
    .A1(_00702_),
    .A2(net2716));
 sg13g2_nor2_1 _11108_ (.A(\core.fetch.cmd_data[6] ),
    .B(net3049),
    .Y(_05295_));
 sg13g2_a21oi_1 _11109_ (.A1(_00704_),
    .A2(net3049),
    .Y(_05296_),
    .B1(_05295_));
 sg13g2_nand3_1 _11110_ (.B(net2719),
    .C(_05296_),
    .A(net2883),
    .Y(_05297_));
 sg13g2_o21ai_1 _11111_ (.B1(_05297_),
    .Y(_00542_),
    .A1(_00704_),
    .A2(net2719));
 sg13g2_nor2_1 _11112_ (.A(\core.fetch.cmd_data[7] ),
    .B(net3049),
    .Y(_05298_));
 sg13g2_a21oi_1 _11113_ (.A1(_00707_),
    .A2(net3049),
    .Y(_05299_),
    .B1(_05298_));
 sg13g2_nand3_1 _11114_ (.B(net2719),
    .C(_05299_),
    .A(net2883),
    .Y(_05300_));
 sg13g2_o21ai_1 _11115_ (.B1(_05300_),
    .Y(_00543_),
    .A1(_00707_),
    .A2(net2719));
 sg13g2_mux2_1 _11116_ (.A0(_02582_),
    .A1(\core.work.registers.state[1] ),
    .S(\core.work.registers.state[2] ),
    .X(_05301_));
 sg13g2_inv_1 _11117_ (.Y(_05302_),
    .A(_05301_));
 sg13g2_and2_1 _11118_ (.A(_00734_),
    .B(_05301_),
    .X(_05303_));
 sg13g2_nor2b_1 _11119_ (.A(_02438_),
    .B_N(_02439_),
    .Y(_05304_));
 sg13g2_a21oi_2 _11120_ (.B1(_05304_),
    .Y(_05305_),
    .A2(_05303_),
    .A1(_00735_));
 sg13g2_o21ai_1 _11121_ (.B1(_00737_),
    .Y(_00544_),
    .A1(_00651_),
    .A2(_05305_));
 sg13g2_o21ai_1 _11122_ (.B1(_00734_),
    .Y(_05306_),
    .A1(net2875),
    .A2(_05302_));
 sg13g2_mux2_1 _11123_ (.A0(net742),
    .A1(_05306_),
    .S(_05305_),
    .X(_00545_));
 sg13g2_nand2_1 _11124_ (.Y(_05307_),
    .A(net2875),
    .B(_05303_));
 sg13g2_nand2_1 _11125_ (.Y(_05308_),
    .A(_00736_),
    .B(_05307_));
 sg13g2_mux2_1 _11126_ (.A0(net544),
    .A1(_05308_),
    .S(_05305_),
    .X(_00546_));
 sg13g2_nor2b_1 _11127_ (.A(net2879),
    .B_N(\core.gpio.stray_data_i[0] ),
    .Y(_05309_));
 sg13g2_a21oi_2 _11128_ (.B1(_05309_),
    .Y(_05310_),
    .A2(net2878),
    .A1(net895));
 sg13g2_nor2_1 _11129_ (.A(net514),
    .B(net2819),
    .Y(_05311_));
 sg13g2_a21oi_1 _11130_ (.A1(net2818),
    .A2(_05310_),
    .Y(_00547_),
    .B1(_05311_));
 sg13g2_nor2b_1 _11131_ (.A(net2879),
    .B_N(\core.gpio.stray_data_i[1] ),
    .Y(_05312_));
 sg13g2_a21oi_2 _11132_ (.B1(_05312_),
    .Y(_05313_),
    .A2(net2878),
    .A1(net744));
 sg13g2_nor2_1 _11133_ (.A(net3437),
    .B(net2818),
    .Y(_05314_));
 sg13g2_a21oi_1 _11134_ (.A1(net2818),
    .A2(_05313_),
    .Y(_00548_),
    .B1(_05314_));
 sg13g2_nor2b_1 _11135_ (.A(net2879),
    .B_N(\core.gpio.stray_data_i[2] ),
    .Y(_05315_));
 sg13g2_a21oi_2 _11136_ (.B1(_05315_),
    .Y(_05316_),
    .A2(net2878),
    .A1(net3498));
 sg13g2_nor2_1 _11137_ (.A(net3435),
    .B(net2819),
    .Y(_05317_));
 sg13g2_a21oi_1 _11138_ (.A1(net2819),
    .A2(_05316_),
    .Y(_00549_),
    .B1(_05317_));
 sg13g2_nor2b_1 _11139_ (.A(net2877),
    .B_N(net668),
    .Y(_05318_));
 sg13g2_a21oi_2 _11140_ (.B1(_05318_),
    .Y(_05319_),
    .A2(net2877),
    .A1(net3496));
 sg13g2_nor2_1 _11141_ (.A(net694),
    .B(net2818),
    .Y(_05320_));
 sg13g2_a21oi_1 _11142_ (.A1(net2816),
    .A2(_05319_),
    .Y(_00550_),
    .B1(_05320_));
 sg13g2_nor2b_1 _11143_ (.A(net2878),
    .B_N(\core.gpio.stray_data_i[4] ),
    .Y(_05321_));
 sg13g2_a21oi_2 _11144_ (.B1(_05321_),
    .Y(_05322_),
    .A2(net2878),
    .A1(net3495));
 sg13g2_nor2_1 _11145_ (.A(net3431),
    .B(net2818),
    .Y(_05323_));
 sg13g2_a21oi_1 _11146_ (.A1(net2818),
    .A2(_05322_),
    .Y(_00551_),
    .B1(_05323_));
 sg13g2_nor2b_2 _11147_ (.A(net2873),
    .B_N(\core.gpio.stray_data_i[5] ),
    .Y(_05324_));
 sg13g2_a21oi_1 _11148_ (.A1(net3489),
    .A2(net2872),
    .Y(_05325_),
    .B1(_05324_));
 sg13g2_nor2_1 _11149_ (.A(net576),
    .B(net2813),
    .Y(_05326_));
 sg13g2_a21oi_1 _11150_ (.A1(net2815),
    .A2(_05325_),
    .Y(_00552_),
    .B1(_05326_));
 sg13g2_nor2b_1 _11151_ (.A(net2878),
    .B_N(\core.gpio.stray_data_i[6] ),
    .Y(_05327_));
 sg13g2_a21oi_2 _11152_ (.B1(_05327_),
    .Y(_05328_),
    .A2(net2878),
    .A1(\core.e2m_addr[6] ));
 sg13g2_nor2_1 _11153_ (.A(net525),
    .B(net2818),
    .Y(_05329_));
 sg13g2_a21oi_1 _11154_ (.A1(net2818),
    .A2(_05328_),
    .Y(_00553_),
    .B1(_05329_));
 sg13g2_nor2b_1 _11155_ (.A(net2873),
    .B_N(\core.gpio.stray_data_i[7] ),
    .Y(_05330_));
 sg13g2_a21oi_2 _11156_ (.B1(_05330_),
    .Y(_05331_),
    .A2(net2873),
    .A1(\core.e2m_addr[7] ));
 sg13g2_nor2_1 _11157_ (.A(net394),
    .B(net2817),
    .Y(_05332_));
 sg13g2_a21oi_1 _11158_ (.A1(net2817),
    .A2(_05331_),
    .Y(_00554_),
    .B1(_05332_));
 sg13g2_nand3_1 _11159_ (.B(\core.gpio.stray_data_i[7] ),
    .C(\core.lsu.is_signed ),
    .A(net3524),
    .Y(_05333_));
 sg13g2_nand2b_1 _11160_ (.Y(_05334_),
    .B(\core.gpio.stray_data_i[8] ),
    .A_N(net3523));
 sg13g2_a21oi_1 _11161_ (.A1(_05333_),
    .A2(_05334_),
    .Y(_05335_),
    .B1(net2874));
 sg13g2_a21oi_2 _11162_ (.B1(_05335_),
    .Y(_05336_),
    .A2(net2874),
    .A1(\core.e2m_addr[8] ));
 sg13g2_nor2_1 _11163_ (.A(net3422),
    .B(net2815),
    .Y(_05337_));
 sg13g2_a21oi_1 _11164_ (.A1(net2813),
    .A2(_05336_),
    .Y(_00555_),
    .B1(_05337_));
 sg13g2_nand2b_1 _11165_ (.Y(_05338_),
    .B(\core.gpio.stray_data_i[9] ),
    .A_N(\core.lsu.is_byte ));
 sg13g2_a21oi_1 _11166_ (.A1(net3286),
    .A2(_05338_),
    .Y(_05339_),
    .B1(net2876));
 sg13g2_a21oi_2 _11167_ (.B1(_05339_),
    .Y(_05340_),
    .A2(net2876),
    .A1(net3488));
 sg13g2_nor2_1 _11168_ (.A(net3419),
    .B(net2816),
    .Y(_05341_));
 sg13g2_a21oi_1 _11169_ (.A1(net2816),
    .A2(_05340_),
    .Y(_00556_),
    .B1(_05341_));
 sg13g2_nand2b_1 _11170_ (.Y(_05342_),
    .B(\core.gpio.stray_data_i[10] ),
    .A_N(net3524));
 sg13g2_a21oi_1 _11171_ (.A1(net3286),
    .A2(_05342_),
    .Y(_05343_),
    .B1(net2873));
 sg13g2_a21oi_2 _11172_ (.B1(_05343_),
    .Y(_05344_),
    .A2(net2874),
    .A1(net3486));
 sg13g2_nor2_1 _11173_ (.A(net3418),
    .B(net2814),
    .Y(_05345_));
 sg13g2_a21oi_1 _11174_ (.A1(net2814),
    .A2(_05344_),
    .Y(_00557_),
    .B1(_05345_));
 sg13g2_nand2b_1 _11175_ (.Y(_05346_),
    .B(\core.gpio.stray_data_i[11] ),
    .A_N(net3523));
 sg13g2_a21oi_1 _11176_ (.A1(net3286),
    .A2(_05346_),
    .Y(_05347_),
    .B1(net2873));
 sg13g2_a21oi_2 _11177_ (.B1(_05347_),
    .Y(_05348_),
    .A2(net2873),
    .A1(\core.e2m_addr[11] ));
 sg13g2_nor2_1 _11178_ (.A(net3416),
    .B(net2811),
    .Y(_05349_));
 sg13g2_a21oi_1 _11179_ (.A1(net2811),
    .A2(_05348_),
    .Y(_00558_),
    .B1(_05349_));
 sg13g2_nand2b_1 _11180_ (.Y(_05350_),
    .B(\core.gpio.stray_data_i[12] ),
    .A_N(net3523));
 sg13g2_a21oi_2 _11181_ (.B1(net2876),
    .Y(_05351_),
    .A2(_05350_),
    .A1(net3286));
 sg13g2_a21oi_2 _11182_ (.B1(_05351_),
    .Y(_05352_),
    .A2(net2872),
    .A1(net3484));
 sg13g2_nor2_1 _11183_ (.A(net583),
    .B(net2813),
    .Y(_05353_));
 sg13g2_a21oi_1 _11184_ (.A1(net2813),
    .A2(_05352_),
    .Y(_00559_),
    .B1(_05353_));
 sg13g2_nand2b_1 _11185_ (.Y(_05354_),
    .B(\core.gpio.stray_data_i[13] ),
    .A_N(net3524));
 sg13g2_a21oi_2 _11186_ (.B1(net2874),
    .Y(_05355_),
    .A2(_05354_),
    .A1(net3286));
 sg13g2_a21oi_2 _11187_ (.B1(_05355_),
    .Y(_05356_),
    .A2(net2874),
    .A1(net3482));
 sg13g2_nor2_1 _11188_ (.A(net511),
    .B(net2814),
    .Y(_05357_));
 sg13g2_a21oi_1 _11189_ (.A1(net2814),
    .A2(_05356_),
    .Y(_00560_),
    .B1(_05357_));
 sg13g2_nand2b_1 _11190_ (.Y(_05358_),
    .B(\core.gpio.stray_data_i[14] ),
    .A_N(net3524));
 sg13g2_a21oi_2 _11191_ (.B1(net2873),
    .Y(_05359_),
    .A2(_05358_),
    .A1(net3286));
 sg13g2_a21oi_2 _11192_ (.B1(_05359_),
    .Y(_05360_),
    .A2(net2872),
    .A1(net3480));
 sg13g2_nor2_1 _11193_ (.A(net3409),
    .B(net2814),
    .Y(_05361_));
 sg13g2_a21oi_1 _11194_ (.A1(net2814),
    .A2(_05360_),
    .Y(_00561_),
    .B1(_05361_));
 sg13g2_nand2b_1 _11195_ (.Y(_05362_),
    .B(\core.gpio.stray_data_i[15] ),
    .A_N(net3524));
 sg13g2_a21oi_2 _11196_ (.B1(net2874),
    .Y(_05363_),
    .A2(_05362_),
    .A1(net3286));
 sg13g2_a21oi_1 _11197_ (.A1(net3473),
    .A2(net2875),
    .Y(_05364_),
    .B1(_05363_));
 sg13g2_nor2_1 _11198_ (.A(net3407),
    .B(net2810),
    .Y(_05365_));
 sg13g2_a21oi_1 _11199_ (.A1(net2810),
    .A2(_05364_),
    .Y(_00562_),
    .B1(_05365_));
 sg13g2_nand2_1 _11200_ (.Y(_05366_),
    .A(\core.lsu.is_half ),
    .B(\core.lsu.is_signed ));
 sg13g2_o21ai_1 _11201_ (.B1(net3286),
    .Y(_05367_),
    .A1(_05362_),
    .A2(_05366_));
 sg13g2_a21oi_2 _11202_ (.B1(_05367_),
    .Y(_05368_),
    .A2(_01132_),
    .A1(\core.gpio.stray_data_i[16] ));
 sg13g2_nor2_2 _11203_ (.A(net2876),
    .B(_05368_),
    .Y(_05369_));
 sg13g2_a21oi_1 _11204_ (.A1(net3472),
    .A2(net2877),
    .Y(_05370_),
    .B1(_05369_));
 sg13g2_nor2_1 _11205_ (.A(net3404),
    .B(net2816),
    .Y(_05371_));
 sg13g2_a21oi_1 _11206_ (.A1(net2816),
    .A2(_05370_),
    .Y(_00563_),
    .B1(_05371_));
 sg13g2_a21oi_2 _11207_ (.B1(net3047),
    .Y(_05372_),
    .A2(net3351),
    .A1(\core.gpio.stray_data_i[17] ));
 sg13g2_nor2_2 _11208_ (.A(net2876),
    .B(_05372_),
    .Y(_05373_));
 sg13g2_a21oi_1 _11209_ (.A1(net3470),
    .A2(net2877),
    .Y(_05374_),
    .B1(_05373_));
 sg13g2_nor2_1 _11210_ (.A(net599),
    .B(net2816),
    .Y(_05375_));
 sg13g2_a21oi_1 _11211_ (.A1(net2817),
    .A2(_05374_),
    .Y(_00564_),
    .B1(_05375_));
 sg13g2_a21oi_2 _11212_ (.B1(net3047),
    .Y(_05376_),
    .A2(net3351),
    .A1(\core.gpio.stray_data_i[18] ));
 sg13g2_nor2_2 _11213_ (.A(net2873),
    .B(_05376_),
    .Y(_05377_));
 sg13g2_a21oi_1 _11214_ (.A1(net3468),
    .A2(net2872),
    .Y(_05378_),
    .B1(_05377_));
 sg13g2_nor2_1 _11215_ (.A(net648),
    .B(net2813),
    .Y(_05379_));
 sg13g2_a21oi_1 _11216_ (.A1(net2813),
    .A2(_05378_),
    .Y(_00565_),
    .B1(_05379_));
 sg13g2_a21oi_2 _11217_ (.B1(net3047),
    .Y(_05380_),
    .A2(net3351),
    .A1(\core.gpio.stray_data_i[19] ));
 sg13g2_nor2_2 _11218_ (.A(net2878),
    .B(_05380_),
    .Y(_05381_));
 sg13g2_a21oi_2 _11219_ (.B1(_05381_),
    .Y(_05382_),
    .A2(net2879),
    .A1(\core.e2m_addr[19] ));
 sg13g2_nor2_1 _11220_ (.A(net409),
    .B(net2819),
    .Y(_05383_));
 sg13g2_a21oi_1 _11221_ (.A1(net2819),
    .A2(_05382_),
    .Y(_00566_),
    .B1(_05383_));
 sg13g2_a21oi_2 _11222_ (.B1(net3047),
    .Y(_05384_),
    .A2(net3351),
    .A1(\core.gpio.stray_data_i[20] ));
 sg13g2_nor2_2 _11223_ (.A(net2876),
    .B(_05384_),
    .Y(_05385_));
 sg13g2_a21oi_1 _11224_ (.A1(net3467),
    .A2(net2877),
    .Y(_05386_),
    .B1(_05385_));
 sg13g2_nor2_1 _11225_ (.A(net3394),
    .B(net2817),
    .Y(_05387_));
 sg13g2_a21oi_1 _11226_ (.A1(net2817),
    .A2(_05386_),
    .Y(_00567_),
    .B1(_05387_));
 sg13g2_a21oi_2 _11227_ (.B1(net3047),
    .Y(_05388_),
    .A2(net3351),
    .A1(\core.gpio.stray_data_i[21] ));
 sg13g2_nor2_1 _11228_ (.A(net2870),
    .B(_05388_),
    .Y(_05389_));
 sg13g2_a21oi_1 _11229_ (.A1(net3459),
    .A2(net2872),
    .Y(_05390_),
    .B1(_05389_));
 sg13g2_nor2_1 _11230_ (.A(net3392),
    .B(net2813),
    .Y(_05391_));
 sg13g2_a21oi_1 _11231_ (.A1(net2813),
    .A2(_05390_),
    .Y(_00568_),
    .B1(_05391_));
 sg13g2_a21oi_2 _11232_ (.B1(net3046),
    .Y(_05392_),
    .A2(net3350),
    .A1(\core.gpio.stray_data_i[22] ));
 sg13g2_nor2_1 _11233_ (.A(net2869),
    .B(_05392_),
    .Y(_05393_));
 sg13g2_a21oi_2 _11234_ (.B1(_05393_),
    .Y(_05394_),
    .A2(net2869),
    .A1(net3456));
 sg13g2_nor2_1 _11235_ (.A(net440),
    .B(net2811),
    .Y(_05395_));
 sg13g2_a21oi_1 _11236_ (.A1(net2811),
    .A2(_05394_),
    .Y(_00569_),
    .B1(_05395_));
 sg13g2_a21oi_2 _11237_ (.B1(net3046),
    .Y(_05396_),
    .A2(net3350),
    .A1(\core.gpio.stray_data_i[23] ));
 sg13g2_nor2_1 _11238_ (.A(net2869),
    .B(_05396_),
    .Y(_05397_));
 sg13g2_a21oi_1 _11239_ (.A1(net3454),
    .A2(net2875),
    .Y(_05398_),
    .B1(_05397_));
 sg13g2_nor2_1 _11240_ (.A(net403),
    .B(net2810),
    .Y(_05399_));
 sg13g2_a21oi_1 _11241_ (.A1(net2810),
    .A2(_05398_),
    .Y(_00570_),
    .B1(_05399_));
 sg13g2_a21oi_1 _11242_ (.A1(\core.gpio.stray_data_i[24] ),
    .A2(_01132_),
    .Y(_05400_),
    .B1(net3047));
 sg13g2_nor2_1 _11243_ (.A(net2876),
    .B(_05400_),
    .Y(_05401_));
 sg13g2_a21oi_2 _11244_ (.B1(_05401_),
    .Y(_05402_),
    .A2(net2876),
    .A1(net3451));
 sg13g2_nor2_1 _11245_ (.A(net3384),
    .B(net2816),
    .Y(_05403_));
 sg13g2_a21oi_1 _11246_ (.A1(net2816),
    .A2(_05402_),
    .Y(_00571_),
    .B1(_05403_));
 sg13g2_a21oi_2 _11247_ (.B1(net3047),
    .Y(_05404_),
    .A2(net3351),
    .A1(\core.gpio.stray_data_i[25] ));
 sg13g2_nor2_1 _11248_ (.A(net2872),
    .B(_05404_),
    .Y(_05405_));
 sg13g2_a21oi_1 _11249_ (.A1(net3449),
    .A2(net2872),
    .Y(_05406_),
    .B1(_05405_));
 sg13g2_nor2_1 _11250_ (.A(net3381),
    .B(net2814),
    .Y(_05407_));
 sg13g2_a21oi_1 _11251_ (.A1(net2814),
    .A2(_05406_),
    .Y(_00572_),
    .B1(_05407_));
 sg13g2_a21oi_2 _11252_ (.B1(net3046),
    .Y(_05408_),
    .A2(net3350),
    .A1(\core.gpio.stray_data_i[26] ));
 sg13g2_nor2_1 _11253_ (.A(net2869),
    .B(_05408_),
    .Y(_05409_));
 sg13g2_a21oi_2 _11254_ (.B1(_05409_),
    .Y(_05410_),
    .A2(net2870),
    .A1(\core.e2m_addr[26] ));
 sg13g2_nor2_1 _11255_ (.A(net647),
    .B(net2810),
    .Y(_05411_));
 sg13g2_a21oi_1 _11256_ (.A1(net2810),
    .A2(_05410_),
    .Y(_00573_),
    .B1(_05411_));
 sg13g2_a21oi_2 _11257_ (.B1(net3046),
    .Y(_05412_),
    .A2(net3350),
    .A1(\core.gpio.stray_data_i[27] ));
 sg13g2_nor2_1 _11258_ (.A(net2870),
    .B(_05412_),
    .Y(_05413_));
 sg13g2_a21oi_2 _11259_ (.B1(_05413_),
    .Y(_05414_),
    .A2(net2870),
    .A1(net3448));
 sg13g2_nor2_1 _11260_ (.A(net595),
    .B(net2811),
    .Y(_05415_));
 sg13g2_a21oi_1 _11261_ (.A1(net2811),
    .A2(_05414_),
    .Y(_00574_),
    .B1(_05415_));
 sg13g2_a21oi_2 _11262_ (.B1(net3046),
    .Y(_05416_),
    .A2(net3350),
    .A1(\core.gpio.stray_data_i[28] ));
 sg13g2_nor2_1 _11263_ (.A(net2869),
    .B(_05416_),
    .Y(_05417_));
 sg13g2_a21oi_2 _11264_ (.B1(_05417_),
    .Y(_05418_),
    .A2(net2869),
    .A1(net3447));
 sg13g2_nor2_1 _11265_ (.A(net620),
    .B(net2809),
    .Y(_05419_));
 sg13g2_a21oi_1 _11266_ (.A1(net2809),
    .A2(_05418_),
    .Y(_00575_),
    .B1(_05419_));
 sg13g2_a21oi_2 _11267_ (.B1(net3046),
    .Y(_05420_),
    .A2(net3350),
    .A1(\core.gpio.stray_data_i[29] ));
 sg13g2_nor2_1 _11268_ (.A(net2871),
    .B(_05420_),
    .Y(_05421_));
 sg13g2_a21oi_2 _11269_ (.B1(_05421_),
    .Y(_05422_),
    .A2(net2871),
    .A1(net3446));
 sg13g2_nor2_1 _11270_ (.A(net626),
    .B(net2809),
    .Y(_05423_));
 sg13g2_a21oi_1 _11271_ (.A1(net2809),
    .A2(_05422_),
    .Y(_00576_),
    .B1(_05423_));
 sg13g2_a21oi_2 _11272_ (.B1(net3046),
    .Y(_05424_),
    .A2(net3350),
    .A1(\core.gpio.stray_data_i[30] ));
 sg13g2_nor2_1 _11273_ (.A(net2874),
    .B(_05424_),
    .Y(_05425_));
 sg13g2_a21oi_2 _11274_ (.B1(_05425_),
    .Y(_05426_),
    .A2(net2871),
    .A1(net3444));
 sg13g2_nor2_1 _11275_ (.A(net3368),
    .B(net2810),
    .Y(_05427_));
 sg13g2_a21oi_1 _11276_ (.A1(net2810),
    .A2(_05426_),
    .Y(_00577_),
    .B1(_05427_));
 sg13g2_a21oi_2 _11277_ (.B1(net3046),
    .Y(_05428_),
    .A2(net3350),
    .A1(\core.gpio.stray_data_i[31] ));
 sg13g2_nor2_1 _11278_ (.A(net2869),
    .B(_05428_),
    .Y(_05429_));
 sg13g2_a21oi_2 _11279_ (.B1(_05429_),
    .Y(_05430_),
    .A2(net2869),
    .A1(net3443));
 sg13g2_nor2_1 _11280_ (.A(net3365),
    .B(net2809),
    .Y(_05431_));
 sg13g2_a21oi_1 _11281_ (.A1(net2809),
    .A2(_05430_),
    .Y(_00578_),
    .B1(_05431_));
 sg13g2_inv_1 _11283__3 (.Y(net343),
    .A(clknet_2_0__leaf_clk));
 sg13g2_inv_1 _11284__4 (.Y(net344),
    .A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 _11285__5 (.Y(net345),
    .A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 _11286__6 (.Y(net346),
    .A(clknet_2_3__leaf_clk));
 sg13g2_inv_1 _11287__7 (.Y(net347),
    .A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 _11288__8 (.Y(net348),
    .A(clknet_2_3__leaf_clk));
 sg13g2_inv_1 _11289__9 (.Y(net349),
    .A(clknet_2_0__leaf_clk));
 sg13g2_inv_1 _11290__10 (.Y(net350),
    .A(clknet_2_3__leaf_clk));
 sg13g2_inv_1 _11291__11 (.Y(net351),
    .A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 _11292__12 (.Y(net352),
    .A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 _11293__13 (.Y(net353),
    .A(clknet_2_0__leaf_clk));
 sg13g2_inv_1 _11294__14 (.Y(net354),
    .A(clknet_2_0__leaf_clk));
 sg13g2_inv_1 _11295__15 (.Y(net355),
    .A(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbp_1 _11296_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3585),
    .D(_00183_),
    .Q_N(_05691_),
    .Q(\core.fetch.state[0] ));
 sg13g2_dfrbp_1 _11297_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3586),
    .D(_00184_),
    .Q_N(_05690_),
    .Q(\core.fetch.state[1] ));
 sg13g2_dfrbp_1 _11298_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net332),
    .D(_00185_),
    .Q_N(_05689_),
    .Q(\core.fetch.data[0] ));
 sg13g2_dfrbp_1 _11299_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net331),
    .D(_00186_),
    .Q_N(_05688_),
    .Q(\core.fetch.data[1] ));
 sg13g2_dfrbp_1 _11300_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net330),
    .D(net570),
    .Q_N(_05687_),
    .Q(\core.fetch.data[2] ));
 sg13g2_dfrbp_1 _11301_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net329),
    .D(net466),
    .Q_N(_05686_),
    .Q(\core.fetch.data[3] ));
 sg13g2_dfrbp_1 _11302_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net328),
    .D(net594),
    .Q_N(_05685_),
    .Q(\core.fetch.data[4] ));
 sg13g2_dfrbp_1 _11303_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net327),
    .D(net402),
    .Q_N(_05684_),
    .Q(\core.fetch.data[5] ));
 sg13g2_dfrbp_1 _11304_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net326),
    .D(net443),
    .Q_N(_05683_),
    .Q(\core.fetch.data[6] ));
 sg13g2_dfrbp_1 _11305_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net325),
    .D(net456),
    .Q_N(_05682_),
    .Q(\core.fetch.data[7] ));
 sg13g2_dfrbp_1 _11306_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net324),
    .D(_00193_),
    .Q_N(_05681_),
    .Q(\core.fetch.data[8] ));
 sg13g2_dfrbp_1 _11307_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net323),
    .D(net480),
    .Q_N(_05680_),
    .Q(\core.fetch.data[9] ));
 sg13g2_dfrbp_1 _11308_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net322),
    .D(net505),
    .Q_N(_05679_),
    .Q(\core.fetch.data[10] ));
 sg13g2_dfrbp_1 _11309_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net321),
    .D(_00196_),
    .Q_N(_05678_),
    .Q(\core.fetch.data[11] ));
 sg13g2_dfrbp_1 _11310_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net320),
    .D(net643),
    .Q_N(_05677_),
    .Q(\core.fetch.data[12] ));
 sg13g2_dfrbp_1 _11311_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net319),
    .D(net398),
    .Q_N(_05676_),
    .Q(\core.fetch.data[13] ));
 sg13g2_dfrbp_1 _11312_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net318),
    .D(net391),
    .Q_N(_05675_),
    .Q(\core.fetch.data[14] ));
 sg13g2_dfrbp_1 _11313_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net317),
    .D(net523),
    .Q_N(_05674_),
    .Q(\core.fetch.data[15] ));
 sg13g2_dfrbp_1 _11314_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net316),
    .D(net478),
    .Q_N(_05673_),
    .Q(\core.fetch.data[16] ));
 sg13g2_dfrbp_1 _11315_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net315),
    .D(net516),
    .Q_N(_05672_),
    .Q(\core.fetch.data[17] ));
 sg13g2_dfrbp_1 _11316_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net314),
    .D(net602),
    .Q_N(_05671_),
    .Q(\core.fetch.data[18] ));
 sg13g2_dfrbp_1 _11317_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net313),
    .D(net453),
    .Q_N(_05670_),
    .Q(\core.fetch.data[19] ));
 sg13g2_dfrbp_1 _11318_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net312),
    .D(net501),
    .Q_N(_05669_),
    .Q(\core.fetch.data[20] ));
 sg13g2_dfrbp_1 _11319_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net311),
    .D(net422),
    .Q_N(_05668_),
    .Q(\core.fetch.data[21] ));
 sg13g2_dfrbp_1 _11320_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net310),
    .D(net430),
    .Q_N(_05667_),
    .Q(\core.fetch.data[22] ));
 sg13g2_dfrbp_1 _11321_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net309),
    .D(net412),
    .Q_N(_05666_),
    .Q(\core.fetch.data[23] ));
 sg13g2_dfrbp_1 _11322_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net308),
    .D(_00209_),
    .Q_N(_05665_),
    .Q(\core.fetch.data[24] ));
 sg13g2_dfrbp_1 _11323_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net307),
    .D(net371),
    .Q_N(_05664_),
    .Q(\core.fetch.data[25] ));
 sg13g2_dfrbp_1 _11324_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net306),
    .D(net405),
    .Q_N(_05663_),
    .Q(\core.fetch.data[26] ));
 sg13g2_dfrbp_1 _11325_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net305),
    .D(net384),
    .Q_N(_05662_),
    .Q(\core.fetch.data[27] ));
 sg13g2_dfrbp_1 _11326_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net304),
    .D(net368),
    .Q_N(_05661_),
    .Q(\core.fetch.data[28] ));
 sg13g2_dfrbp_1 _11327_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net303),
    .D(net389),
    .Q_N(_05660_),
    .Q(\core.fetch.data[29] ));
 sg13g2_dfrbp_1 _11328_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net302),
    .D(net424),
    .Q_N(_05659_),
    .Q(\core.fetch.data[30] ));
 sg13g2_dfrbp_1 _11329_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net301),
    .D(net417),
    .Q_N(_05658_),
    .Q(\core.fetch.data[31] ));
 sg13g2_dfrbp_1 _11330_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net3586),
    .D(net790),
    .Q_N(_05657_),
    .Q(\core.fetch.data_size[0] ));
 sg13g2_dfrbp_1 _11331_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3585),
    .D(_00218_),
    .Q_N(_05656_),
    .Q(\core.fetch.data_size[1] ));
 sg13g2_dfrbp_1 _11332_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net3585),
    .D(net797),
    .Q_N(_05692_),
    .Q(\core.fetch.data_size[2] ));
 sg13g2_dfrbp_1 _11333_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3583),
    .D(net868),
    .Q_N(uio_out[0]),
    .Q(\core.fetch.spi_reader.cs ));
 sg13g2_dfrbp_1 _11334_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3583),
    .D(net358),
    .Q_N(_00105_),
    .Q(\core.fetch.spi_reader.sck ));
 sg13g2_dfrbp_1 _11335_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net300),
    .D(_00221_),
    .Q_N(_00096_),
    .Q(\core.fetch.cmd_data[0] ));
 sg13g2_dfrbp_1 _11336_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net299),
    .D(_00222_),
    .Q_N(_00097_),
    .Q(\core.fetch.cmd_data[1] ));
 sg13g2_dfrbp_1 _11337_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net298),
    .D(_00223_),
    .Q_N(_00098_),
    .Q(\core.fetch.cmd_data[2] ));
 sg13g2_dfrbp_1 _11338_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net297),
    .D(_00224_),
    .Q_N(_00099_),
    .Q(\core.fetch.cmd_data[3] ));
 sg13g2_dfrbp_1 _11339_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net296),
    .D(net879),
    .Q_N(_00100_),
    .Q(\core.fetch.cmd_data[4] ));
 sg13g2_dfrbp_1 _11340_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net295),
    .D(net891),
    .Q_N(_00101_),
    .Q(\core.fetch.cmd_data[5] ));
 sg13g2_dfrbp_1 _11341_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net294),
    .D(_00227_),
    .Q_N(_00102_),
    .Q(\core.fetch.cmd_data[6] ));
 sg13g2_dfrbp_1 _11342_ (.CLK(clknet_leaf_14_clk_regs),
    .RESET_B(net293),
    .D(_00228_),
    .Q_N(_00103_),
    .Q(\core.fetch.cmd_data[7] ));
 sg13g2_dfrbp_1 _11343_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net292),
    .D(_00229_),
    .Q_N(_05655_),
    .Q(\core.fetch.spi_reader.cache_bit ));
 sg13g2_dfrbp_1 _11344_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net291),
    .D(net497),
    .Q_N(_00061_),
    .Q(\core.fetch.spi_reader.addr[0] ));
 sg13g2_dfrbp_1 _11345_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net290),
    .D(_00231_),
    .Q_N(_05654_),
    .Q(\core.fetch.spi_reader.addr[1] ));
 sg13g2_dfrbp_1 _11346_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net289),
    .D(_00232_),
    .Q_N(_00063_),
    .Q(\core.fetch.spi_reader.addr[2] ));
 sg13g2_dfrbp_1 _11347_ (.CLK(clknet_leaf_16_clk_regs),
    .RESET_B(net288),
    .D(net495),
    .Q_N(_05653_),
    .Q(\core.fetch.spi_reader.addr[3] ));
 sg13g2_dfrbp_1 _11348_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net287),
    .D(_00234_),
    .Q_N(_00070_),
    .Q(\core.fetch.spi_reader.addr[4] ));
 sg13g2_dfrbp_1 _11349_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net286),
    .D(_00235_),
    .Q_N(_00068_),
    .Q(\core.fetch.spi_reader.addr[5] ));
 sg13g2_dfrbp_1 _11350_ (.CLK(clknet_leaf_20_clk_regs),
    .RESET_B(net285),
    .D(_00236_),
    .Q_N(_00067_),
    .Q(\core.fetch.spi_reader.addr[6] ));
 sg13g2_dfrbp_1 _11351_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net284),
    .D(_00237_),
    .Q_N(_05652_),
    .Q(\core.fetch.spi_reader.addr[7] ));
 sg13g2_dfrbp_1 _11352_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net283),
    .D(_00238_),
    .Q_N(_00083_),
    .Q(\core.fetch.spi_reader.addr[8] ));
 sg13g2_dfrbp_1 _11353_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net282),
    .D(_00239_),
    .Q_N(_05651_),
    .Q(\core.fetch.spi_reader.addr[9] ));
 sg13g2_dfrbp_1 _11354_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net281),
    .D(_00240_),
    .Q_N(_00081_),
    .Q(\core.fetch.spi_reader.addr[10] ));
 sg13g2_dfrbp_1 _11355_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net280),
    .D(_00241_),
    .Q_N(_05650_),
    .Q(\core.fetch.spi_reader.addr[11] ));
 sg13g2_dfrbp_1 _11356_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net279),
    .D(_00242_),
    .Q_N(_00077_),
    .Q(\core.fetch.spi_reader.addr[12] ));
 sg13g2_dfrbp_1 _11357_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net278),
    .D(_00243_),
    .Q_N(_05649_),
    .Q(\core.fetch.spi_reader.addr[13] ));
 sg13g2_dfrbp_1 _11358_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net277),
    .D(_00244_),
    .Q_N(_00074_),
    .Q(\core.fetch.spi_reader.addr[14] ));
 sg13g2_dfrbp_1 _11359_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net276),
    .D(net548),
    .Q_N(_00071_),
    .Q(\core.fetch.spi_reader.addr[15] ));
 sg13g2_dfrbp_1 _11360_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net3584),
    .D(net782),
    .Q_N(_05648_),
    .Q(\core.fetch.spi_reader.state[0] ));
 sg13g2_dfrbp_1 _11361_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net3584),
    .D(net471),
    .Q_N(_05647_),
    .Q(\core.fetch.spi_reader.state[1] ));
 sg13g2_dfrbp_1 _11362_ (.CLK(clknet_leaf_17_clk_regs),
    .RESET_B(net3584),
    .D(_00248_),
    .Q_N(_00060_),
    .Q(\core.fetch.spi_reader.state[2] ));
 sg13g2_dfrbp_1 _11363_ (.CLK(clknet_leaf_15_clk_regs),
    .RESET_B(net3586),
    .D(_00249_),
    .Q_N(_00019_),
    .Q(\core.fetch.cmd_valid ));
 sg13g2_dfrbp_1 _11364_ (.CLK(clknet_leaf_19_clk_regs),
    .RESET_B(net3584),
    .D(net437),
    .Q_N(_05646_),
    .Q(\core.fetch.spi_reader.dirty ));
 sg13g2_dfrbp_1 _11365_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net3591),
    .D(net637),
    .Q_N(_00104_),
    .Q(\core.f2e_addr[2] ));
 sg13g2_dfrbp_1 _11366_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net3591),
    .D(net623),
    .Q_N(_05645_),
    .Q(\core.f2e_addr[3] ));
 sg13g2_dfrbp_1 _11367_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net3591),
    .D(net428),
    .Q_N(_05644_),
    .Q(\core.f2e_addr[4] ));
 sg13g2_dfrbp_1 _11368_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net3591),
    .D(_00254_),
    .Q_N(_05643_),
    .Q(\core.f2e_addr[5] ));
 sg13g2_dfrbp_1 _11369_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net3594),
    .D(_00255_),
    .Q_N(_05642_),
    .Q(\core.f2e_addr[6] ));
 sg13g2_dfrbp_1 _11370_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net3592),
    .D(_00256_),
    .Q_N(_05641_),
    .Q(\core.f2e_addr[7] ));
 sg13g2_dfrbp_1 _11371_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net3591),
    .D(_00257_),
    .Q_N(_05640_),
    .Q(\core.f2e_addr[8] ));
 sg13g2_dfrbp_1 _11372_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net3591),
    .D(_00258_),
    .Q_N(_05639_),
    .Q(\core.f2e_addr[9] ));
 sg13g2_dfrbp_1 _11373_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net3591),
    .D(_00259_),
    .Q_N(_05638_),
    .Q(\core.f2e_addr[10] ));
 sg13g2_dfrbp_1 _11374_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net3591),
    .D(net686),
    .Q_N(_00078_),
    .Q(\core.f2e_addr[11] ));
 sg13g2_dfrbp_1 _11375_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net3589),
    .D(_00261_),
    .Q_N(_05637_),
    .Q(\core.f2e_addr[12] ));
 sg13g2_dfrbp_1 _11376_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net3589),
    .D(net598),
    .Q_N(_00075_),
    .Q(\core.f2e_addr[13] ));
 sg13g2_dfrbp_1 _11377_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net3589),
    .D(_00263_),
    .Q_N(_05636_),
    .Q(\core.f2e_addr[14] ));
 sg13g2_dfrbp_1 _11378_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net3589),
    .D(net618),
    .Q_N(_05635_),
    .Q(\core.f2e_addr[15] ));
 sg13g2_dfrbp_1 _11379_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net275),
    .D(_00265_),
    .Q_N(_00143_),
    .Q(\core.work.alu.sval2[1] ));
 sg13g2_dfrbp_1 _11380_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net274),
    .D(_00266_),
    .Q_N(_00142_),
    .Q(\core.work.alu.sval2[2] ));
 sg13g2_dfrbp_1 _11381_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net273),
    .D(net758),
    .Q_N(_00109_),
    .Q(\core.work.alu.sval2[3] ));
 sg13g2_dfrbp_1 _11382_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net272),
    .D(_00268_),
    .Q_N(_00054_),
    .Q(\core.work.alu.sval2[4] ));
 sg13g2_dfrbp_1 _11383_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net271),
    .D(_00269_),
    .Q_N(_00112_),
    .Q(\core.work.alu.sval2[5] ));
 sg13g2_dfrbp_1 _11384_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net270),
    .D(_00270_),
    .Q_N(_00113_),
    .Q(\core.work.alu.sval2[6] ));
 sg13g2_dfrbp_1 _11385_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net269),
    .D(_00271_),
    .Q_N(_00114_),
    .Q(\core.work.alu.sval2[7] ));
 sg13g2_dfrbp_1 _11386_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net268),
    .D(net703),
    .Q_N(_00115_),
    .Q(\core.work.alu.sval2[8] ));
 sg13g2_dfrbp_1 _11387_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net267),
    .D(_00273_),
    .Q_N(_00116_),
    .Q(\core.work.alu.sval2[9] ));
 sg13g2_dfrbp_1 _11388_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net266),
    .D(_00274_),
    .Q_N(_00117_),
    .Q(\core.work.alu.sval2[10] ));
 sg13g2_dfrbp_1 _11389_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net265),
    .D(_00275_),
    .Q_N(_00118_),
    .Q(\core.work.alu.sval2[11] ));
 sg13g2_dfrbp_1 _11390_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net264),
    .D(net827),
    .Q_N(_00119_),
    .Q(\core.work.alu.sval2[12] ));
 sg13g2_dfrbp_1 _11391_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net263),
    .D(net741),
    .Q_N(_00121_),
    .Q(\core.work.alu.sval2[13] ));
 sg13g2_dfrbp_1 _11392_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net262),
    .D(_00278_),
    .Q_N(_00123_),
    .Q(\core.work.alu.sval2[14] ));
 sg13g2_dfrbp_1 _11393_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net261),
    .D(net773),
    .Q_N(_00125_),
    .Q(\core.work.alu.sval2[15] ));
 sg13g2_dfrbp_1 _11394_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3588),
    .D(_00280_),
    .Q_N(_00055_),
    .Q(\core.work.alu.is_mem ));
 sg13g2_dfrbp_1 _11395_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net260),
    .D(_00281_),
    .Q_N(_00051_),
    .Q(\core.work.alu.sval2[29] ));
 sg13g2_dfrbp_1 _11396_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net258),
    .D(net665),
    .Q_N(_00053_),
    .Q(\core.work.alu.sval2[31] ));
 sg13g2_dfrbp_1 _11397_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net256),
    .D(_00283_),
    .Q_N(_00144_),
    .Q(\core.work.alu.sval2[0] ));
 sg13g2_dfrbp_1 _11398_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net254),
    .D(net681),
    .Q_N(_00050_),
    .Q(\core.work.alu.sval2[30] ));
 sg13g2_dfrbp_1 _11399_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net252),
    .D(net833),
    .Q_N(_00047_),
    .Q(\core.work.alu.sval2[28] ));
 sg13g2_dfrbp_1 _11400_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net250),
    .D(net812),
    .Q_N(_00045_),
    .Q(\core.work.alu.sval2[27] ));
 sg13g2_dfrbp_1 _11401_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net248),
    .D(net792),
    .Q_N(_00042_),
    .Q(\core.work.alu.sval2[26] ));
 sg13g2_dfrbp_1 _11402_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net246),
    .D(_00288_),
    .Q_N(_00043_),
    .Q(\core.work.alu.sval2[25] ));
 sg13g2_dfrbp_1 _11403_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net244),
    .D(_00289_),
    .Q_N(_00022_),
    .Q(\core.work.alu.sval2[16] ));
 sg13g2_dfrbp_1 _11404_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net242),
    .D(_00290_),
    .Q_N(_00035_),
    .Q(\core.work.alu.sval2[21] ));
 sg13g2_dfrbp_1 _11405_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net240),
    .D(net684),
    .Q_N(_00034_),
    .Q(\core.work.alu.sval2[22] ));
 sg13g2_dfrbp_1 _11406_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net238),
    .D(net861),
    .Q_N(_00037_),
    .Q(\core.work.alu.sval2[23] ));
 sg13g2_dfrbp_1 _11407_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net236),
    .D(net854),
    .Q_N(_00039_),
    .Q(\core.work.alu.sval2[24] ));
 sg13g2_dfrbp_1 _11408_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net234),
    .D(net785),
    .Q_N(_00027_),
    .Q(\core.work.alu.sval2[17] ));
 sg13g2_dfrbp_1 _11409_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net232),
    .D(net711),
    .Q_N(_00026_),
    .Q(\core.work.alu.sval2[18] ));
 sg13g2_dfrbp_1 _11410_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net230),
    .D(_00296_),
    .Q_N(_00029_),
    .Q(\core.work.alu.sval2[19] ));
 sg13g2_dfrbp_1 _11411_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net228),
    .D(net460),
    .Q_N(_00031_),
    .Q(\core.work.alu.sval2[20] ));
 sg13g2_dfrbp_1 _11412_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net3585),
    .D(_00298_),
    .Q_N(_00062_),
    .Q(\core.fetch.inst_size[0] ));
 sg13g2_dfrbp_1 _11413_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net226),
    .D(net527),
    .Q_N(_05634_),
    .Q(\core.work.registers.wr_reg[0] ));
 sg13g2_dfrbp_1 _11414_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net225),
    .D(_00300_),
    .Q_N(_05633_),
    .Q(\core.work.registers.wr_reg[1] ));
 sg13g2_dfrbp_1 _11415_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net224),
    .D(_00301_),
    .Q_N(_05632_),
    .Q(\core.work.registers.wr_reg[2] ));
 sg13g2_dfrbp_1 _11416_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net223),
    .D(_00302_),
    .Q_N(_05631_),
    .Q(\core.work.registers.wr_reg[3] ));
 sg13g2_dfrbp_1 _11417_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3588),
    .D(_00303_),
    .Q_N(_05630_),
    .Q(\core.work.op[4] ));
 sg13g2_dfrbp_1 _11418_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3585),
    .D(_00304_),
    .Q_N(_05629_),
    .Q(\core.fetch.inst_size[1] ));
 sg13g2_dfrbp_1 _11419_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net3585),
    .D(_00305_),
    .Q_N(_05628_),
    .Q(\core.fetch.inst_size[2] ));
 sg13g2_dfrbp_1 _11420_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3583),
    .D(_00306_),
    .Q_N(_05627_),
    .Q(\core.fetch.spi_reader.counter[0] ));
 sg13g2_dfrbp_1 _11421_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3583),
    .D(net366),
    .Q_N(_00163_),
    .Q(\core.fetch.spi_reader.counter[1] ));
 sg13g2_dfrbp_1 _11422_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3583),
    .D(net432),
    .Q_N(_00164_),
    .Q(\core.fetch.spi_reader.counter[2] ));
 sg13g2_dfrbp_1 _11423_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3583),
    .D(net434),
    .Q_N(_00165_),
    .Q(\core.fetch.spi_reader.counter[3] ));
 sg13g2_dfrbp_1 _11424_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3583),
    .D(net377),
    .Q_N(_00166_),
    .Q(\core.fetch.spi_reader.counter[4] ));
 sg13g2_dfrbp_1 _11425_ (.CLK(clknet_leaf_18_clk_regs),
    .RESET_B(net3583),
    .D(net426),
    .Q_N(_00167_),
    .Q(\core.fetch.spi_reader.counter[5] ));
 sg13g2_dfrbp_1 _11426_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net222),
    .D(_00312_),
    .Q_N(_05626_),
    .Q(\core.fetch.rd_addr_i[0] ));
 sg13g2_dfrbp_1 _11427_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net221),
    .D(net396),
    .Q_N(_05625_),
    .Q(\core.fetch.rd_addr_i[1] ));
 sg13g2_dfrbp_1 _11428_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net220),
    .D(_00314_),
    .Q_N(_05624_),
    .Q(\core.fetch.rd_addr_i[2] ));
 sg13g2_dfrbp_1 _11429_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net219),
    .D(net835),
    .Q_N(_00066_),
    .Q(\core.fetch.rd_addr_i[3] ));
 sg13g2_dfrbp_1 _11430_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net218),
    .D(_00316_),
    .Q_N(_05623_),
    .Q(\core.fetch.rd_addr_i[4] ));
 sg13g2_dfrbp_1 _11431_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net217),
    .D(_00317_),
    .Q_N(_00069_),
    .Q(\core.fetch.rd_addr_i[5] ));
 sg13g2_dfrbp_1 _11432_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net216),
    .D(net382),
    .Q_N(_00065_),
    .Q(\core.fetch.rd_addr_i[6] ));
 sg13g2_dfrbp_1 _11433_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net215),
    .D(_00319_),
    .Q_N(_00064_),
    .Q(\core.fetch.rd_addr_i[7] ));
 sg13g2_dfrbp_1 _11434_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net214),
    .D(_00320_),
    .Q_N(_05622_),
    .Q(\core.fetch.rd_addr_i[8] ));
 sg13g2_dfrbp_1 _11435_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net213),
    .D(_00321_),
    .Q_N(_00082_),
    .Q(\core.fetch.rd_addr_i[9] ));
 sg13g2_dfrbp_1 _11436_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net212),
    .D(net386),
    .Q_N(_00080_),
    .Q(\core.fetch.rd_addr_i[10] ));
 sg13g2_dfrbp_1 _11437_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net211),
    .D(net633),
    .Q_N(_00079_),
    .Q(\core.fetch.rd_addr_i[11] ));
 sg13g2_dfrbp_1 _11438_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net210),
    .D(_00324_),
    .Q_N(_05621_),
    .Q(\core.fetch.rd_addr_i[12] ));
 sg13g2_dfrbp_1 _11439_ (.CLK(clknet_leaf_38_clk_regs),
    .RESET_B(net209),
    .D(net631),
    .Q_N(_00076_),
    .Q(\core.fetch.rd_addr_i[13] ));
 sg13g2_dfrbp_1 _11440_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net208),
    .D(_00326_),
    .Q_N(_00073_),
    .Q(\core.fetch.rd_addr_i[14] ));
 sg13g2_dfrbp_1 _11441_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net177),
    .D(_00327_),
    .Q_N(_00072_),
    .Q(\core.fetch.rd_addr_i[15] ));
 sg13g2_dfrbp_1 _11442_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3588),
    .D(net732),
    .Q_N(_05620_),
    .Q(\core.lsu.accept ));
 sg13g2_dfrbp_1 _11443_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3590),
    .D(_00328_),
    .Q_N(_05619_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _11444_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net3587),
    .D(_00329_),
    .Q_N(_05618_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _11445_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3587),
    .D(_00330_),
    .Q_N(_05617_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _11446_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3590),
    .D(_00331_),
    .Q_N(_05616_),
    .Q(uo_out[3]));
 sg13g2_dfrbp_1 _11447_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net3587),
    .D(_00332_),
    .Q_N(_05615_),
    .Q(uo_out[4]));
 sg13g2_dfrbp_1 _11448_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net3587),
    .D(_00333_),
    .Q_N(_05614_),
    .Q(uo_out[5]));
 sg13g2_dfrbp_1 _11449_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net3587),
    .D(_00334_),
    .Q_N(_05613_),
    .Q(uo_out[6]));
 sg13g2_dfrbp_1 _11450_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net3587),
    .D(_00335_),
    .Q_N(_05612_),
    .Q(uo_out[7]));
 sg13g2_dfrbp_1 _11451_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net3586),
    .D(net737),
    .Q_N(_05611_),
    .Q(\core.lsu.state[0] ));
 sg13g2_dfrbp_1 _11452_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net3588),
    .D(net692),
    .Q_N(_05610_),
    .Q(\core.lsu.state[1] ));
 sg13g2_dfrbp_1 _11453_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net3588),
    .D(net591),
    .Q_N(_00021_),
    .Q(\core.lsu.state[2] ));
 sg13g2_dfrbp_1 _11454_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net207),
    .D(_00339_),
    .Q_N(_00059_),
    .Q(\core.gpio.stray_wr_i ));
 sg13g2_dfrbp_1 _11455_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net206),
    .D(net400),
    .Q_N(_05609_),
    .Q(\core.lsu.is_signed ));
 sg13g2_dfrbp_1 _11456_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net205),
    .D(net439),
    .Q_N(_05608_),
    .Q(\core.lsu.is_half ));
 sg13g2_dfrbp_1 _11457_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net204),
    .D(net580),
    .Q_N(_00018_),
    .Q(\core.lsu.spi_valid ));
 sg13g2_dfrbp_1 _11458_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net202),
    .D(_00343_),
    .Q_N(_05607_),
    .Q(\core.lsu.is_byte ));
 sg13g2_dfrbp_1 _11459_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net201),
    .D(_00344_),
    .Q_N(_05606_),
    .Q(\core.gpio.stray_data_i[0] ));
 sg13g2_dfrbp_1 _11460_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net200),
    .D(_00345_),
    .Q_N(_05605_),
    .Q(\core.gpio.stray_data_i[1] ));
 sg13g2_dfrbp_1 _11461_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net199),
    .D(net697),
    .Q_N(_05604_),
    .Q(\core.gpio.stray_data_i[2] ));
 sg13g2_dfrbp_1 _11462_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net198),
    .D(_00347_),
    .Q_N(_05603_),
    .Q(\core.gpio.stray_data_i[3] ));
 sg13g2_dfrbp_1 _11463_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net197),
    .D(_00348_),
    .Q_N(_05602_),
    .Q(\core.gpio.stray_data_i[4] ));
 sg13g2_dfrbp_1 _11464_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net196),
    .D(net688),
    .Q_N(_05601_),
    .Q(\core.gpio.stray_data_i[5] ));
 sg13g2_dfrbp_1 _11465_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net195),
    .D(_00350_),
    .Q_N(_05600_),
    .Q(\core.gpio.stray_data_i[6] ));
 sg13g2_dfrbp_1 _11466_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net194),
    .D(_00351_),
    .Q_N(_05599_),
    .Q(\core.gpio.stray_data_i[7] ));
 sg13g2_dfrbp_1 _11467_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net193),
    .D(_00352_),
    .Q_N(_05598_),
    .Q(\core.gpio.stray_data_i[8] ));
 sg13g2_dfrbp_1 _11468_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net192),
    .D(net727),
    .Q_N(_05597_),
    .Q(\core.gpio.stray_data_i[9] ));
 sg13g2_dfrbp_1 _11469_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net191),
    .D(_00354_),
    .Q_N(_05596_),
    .Q(\core.gpio.stray_data_i[10] ));
 sg13g2_dfrbp_1 _11470_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net190),
    .D(net720),
    .Q_N(_05595_),
    .Q(\core.gpio.stray_data_i[11] ));
 sg13g2_dfrbp_1 _11471_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net189),
    .D(net714),
    .Q_N(_05594_),
    .Q(\core.gpio.stray_data_i[12] ));
 sg13g2_dfrbp_1 _11472_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net188),
    .D(_00357_),
    .Q_N(_05593_),
    .Q(\core.gpio.stray_data_i[13] ));
 sg13g2_dfrbp_1 _11473_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net187),
    .D(net724),
    .Q_N(_05592_),
    .Q(\core.gpio.stray_data_i[14] ));
 sg13g2_dfrbp_1 _11474_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net186),
    .D(_00359_),
    .Q_N(_05591_),
    .Q(\core.gpio.stray_data_i[15] ));
 sg13g2_dfrbp_1 _11475_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net185),
    .D(net652),
    .Q_N(_05590_),
    .Q(\core.gpio.stray_data_i[16] ));
 sg13g2_dfrbp_1 _11476_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net184),
    .D(_00361_),
    .Q_N(_05589_),
    .Q(\core.gpio.stray_data_i[17] ));
 sg13g2_dfrbp_1 _11477_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net183),
    .D(_00362_),
    .Q_N(_05588_),
    .Q(\core.gpio.stray_data_i[18] ));
 sg13g2_dfrbp_1 _11478_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net182),
    .D(_00363_),
    .Q_N(_05587_),
    .Q(\core.gpio.stray_data_i[19] ));
 sg13g2_dfrbp_1 _11479_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net181),
    .D(_00364_),
    .Q_N(_05586_),
    .Q(\core.gpio.stray_data_i[20] ));
 sg13g2_dfrbp_1 _11480_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net180),
    .D(net748),
    .Q_N(_05585_),
    .Q(\core.gpio.stray_data_i[21] ));
 sg13g2_dfrbp_1 _11481_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net179),
    .D(net755),
    .Q_N(_05584_),
    .Q(\core.gpio.stray_data_i[22] ));
 sg13g2_dfrbp_1 _11482_ (.CLK(clknet_leaf_25_clk_regs),
    .RESET_B(net178),
    .D(_00367_),
    .Q_N(_05583_),
    .Q(\core.gpio.stray_data_i[23] ));
 sg13g2_dfrbp_1 _11483_ (.CLK(clknet_leaf_24_clk_regs),
    .RESET_B(net176),
    .D(_00368_),
    .Q_N(_05582_),
    .Q(\core.gpio.stray_data_i[24] ));
 sg13g2_dfrbp_1 _11484_ (.CLK(clknet_leaf_23_clk_regs),
    .RESET_B(net175),
    .D(_00369_),
    .Q_N(_05581_),
    .Q(\core.gpio.stray_data_i[25] ));
 sg13g2_dfrbp_1 _11485_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net174),
    .D(_00370_),
    .Q_N(_05580_),
    .Q(\core.gpio.stray_data_i[26] ));
 sg13g2_dfrbp_1 _11486_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net173),
    .D(_00371_),
    .Q_N(_05579_),
    .Q(\core.gpio.stray_data_i[27] ));
 sg13g2_dfrbp_1 _11487_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net172),
    .D(_00372_),
    .Q_N(_05578_),
    .Q(\core.gpio.stray_data_i[28] ));
 sg13g2_dfrbp_1 _11488_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net171),
    .D(_00373_),
    .Q_N(_05577_),
    .Q(\core.gpio.stray_data_i[29] ));
 sg13g2_dfrbp_1 _11489_ (.CLK(clknet_leaf_22_clk_regs),
    .RESET_B(net170),
    .D(_00374_),
    .Q_N(_05576_),
    .Q(\core.gpio.stray_data_i[30] ));
 sg13g2_dfrbp_1 _11490_ (.CLK(clknet_leaf_21_clk_regs),
    .RESET_B(net169),
    .D(_00375_),
    .Q_N(_05575_),
    .Q(\core.gpio.stray_data_i[31] ));
 sg13g2_dfrbp_1 _11491_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net168),
    .D(_00376_),
    .Q_N(_05574_),
    .Q(\core.lsu.dreg[0] ));
 sg13g2_dfrbp_1 _11492_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net167),
    .D(_00377_),
    .Q_N(_05573_),
    .Q(\core.lsu.dreg[1] ));
 sg13g2_dfrbp_1 _11493_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net166),
    .D(net393),
    .Q_N(_05572_),
    .Q(\core.lsu.dreg[2] ));
 sg13g2_dfrbp_1 _11494_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net165),
    .D(net415),
    .Q_N(_05571_),
    .Q(\core.lsu.dreg[3] ));
 sg13g2_dfrbp_1 _11495_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net3593),
    .D(net361),
    .Q_N(_00128_),
    .Q(\core.lsu.spi.sck ));
 sg13g2_dfrbp_1 _11496_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net84),
    .D(_00381_),
    .Q_N(_05693_),
    .Q(\core.lsu.spi.cache_bit ));
 sg13g2_dfrbp_1 _11497_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net3592),
    .D(_00002_),
    .Q_N(uio_out[4]),
    .Q(\core.lsu.spi.cs ));
 sg13g2_dfrbp_1 _11498_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net3593),
    .D(net462),
    .Q_N(_05570_),
    .Q(\core.lsu.spi.dirty ));
 sg13g2_dfrbp_1 _11499_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net164),
    .D(_00383_),
    .Q_N(_00133_),
    .Q(\core.lsu.spi.buffer[0] ));
 sg13g2_dfrbp_1 _11500_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net163),
    .D(_00384_),
    .Q_N(_00134_),
    .Q(\core.lsu.spi.buffer[1] ));
 sg13g2_dfrbp_1 _11501_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net162),
    .D(_00385_),
    .Q_N(_00135_),
    .Q(\core.lsu.spi.buffer[2] ));
 sg13g2_dfrbp_1 _11502_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net161),
    .D(_00386_),
    .Q_N(_00136_),
    .Q(\core.lsu.spi.buffer[3] ));
 sg13g2_dfrbp_1 _11503_ (.CLK(clknet_leaf_31_clk_regs),
    .RESET_B(net160),
    .D(_00387_),
    .Q_N(_00137_),
    .Q(\core.lsu.spi.buffer[4] ));
 sg13g2_dfrbp_1 _11504_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net159),
    .D(net808),
    .Q_N(_00138_),
    .Q(\core.lsu.spi.buffer[5] ));
 sg13g2_dfrbp_1 _11505_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net158),
    .D(_00389_),
    .Q_N(_00139_),
    .Q(\core.lsu.spi.buffer[6] ));
 sg13g2_dfrbp_1 _11506_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net157),
    .D(_00390_),
    .Q_N(_00140_),
    .Q(\core.lsu.spi.buffer[7] ));
 sg13g2_dfrbp_1 _11507_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net156),
    .D(net482),
    .Q_N(_00085_),
    .Q(\core.lsu.spi.addr[0] ));
 sg13g2_dfrbp_1 _11508_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net155),
    .D(_00392_),
    .Q_N(_05569_),
    .Q(\core.lsu.spi.addr[1] ));
 sg13g2_dfrbp_1 _11509_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net154),
    .D(net552),
    .Q_N(_00086_),
    .Q(\core.lsu.spi.addr[2] ));
 sg13g2_dfrbp_1 _11510_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net153),
    .D(_00394_),
    .Q_N(_05568_),
    .Q(\core.lsu.spi.addr[3] ));
 sg13g2_dfrbp_1 _11511_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net152),
    .D(net510),
    .Q_N(_00089_),
    .Q(\core.lsu.spi.addr[4] ));
 sg13g2_dfrbp_1 _11512_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net151),
    .D(net557),
    .Q_N(_00088_),
    .Q(\core.lsu.spi.addr[5] ));
 sg13g2_dfrbp_1 _11513_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net150),
    .D(_00397_),
    .Q_N(_00087_),
    .Q(\core.lsu.spi.addr[6] ));
 sg13g2_dfrbp_1 _11514_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net149),
    .D(_00398_),
    .Q_N(_05567_),
    .Q(\core.lsu.spi.addr[7] ));
 sg13g2_dfrbp_1 _11515_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net148),
    .D(_00399_),
    .Q_N(_00095_),
    .Q(\core.lsu.spi.addr[8] ));
 sg13g2_dfrbp_1 _11516_ (.CLK(clknet_leaf_36_clk_regs),
    .RESET_B(net147),
    .D(_00400_),
    .Q_N(_00094_),
    .Q(\core.lsu.spi.addr[9] ));
 sg13g2_dfrbp_1 _11517_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net146),
    .D(_00401_),
    .Q_N(_00093_),
    .Q(\core.lsu.spi.addr[10] ));
 sg13g2_dfrbp_1 _11518_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net145),
    .D(net780),
    .Q_N(_05566_),
    .Q(\core.lsu.spi.addr[11] ));
 sg13g2_dfrbp_1 _11519_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net144),
    .D(_00403_),
    .Q_N(_00092_),
    .Q(\core.lsu.spi.addr[12] ));
 sg13g2_dfrbp_1 _11520_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net143),
    .D(net820),
    .Q_N(_05565_),
    .Q(\core.lsu.spi.addr[13] ));
 sg13g2_dfrbp_1 _11521_ (.CLK(clknet_leaf_37_clk_regs),
    .RESET_B(net142),
    .D(_00405_),
    .Q_N(_00091_),
    .Q(\core.lsu.spi.addr[14] ));
 sg13g2_dfrbp_1 _11522_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net141),
    .D(net373),
    .Q_N(_00090_),
    .Q(\core.lsu.spi.addr[15] ));
 sg13g2_dfrbp_1 _11523_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net3592),
    .D(_00407_),
    .Q_N(_05564_),
    .Q(\core.lsu.spi.state[0] ));
 sg13g2_dfrbp_1 _11524_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net3592),
    .D(net718),
    .Q_N(_05563_),
    .Q(\core.lsu.spi.state[1] ));
 sg13g2_dfrbp_1 _11525_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net3592),
    .D(_00409_),
    .Q_N(_00084_),
    .Q(\core.lsu.spi.state[2] ));
 sg13g2_dfrbp_1 _11526_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net3590),
    .D(_00410_),
    .Q_N(_05562_),
    .Q(\core.lsu.write_index[0] ));
 sg13g2_dfrbp_1 _11527_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net3590),
    .D(_00411_),
    .Q_N(_00056_),
    .Q(\core.lsu.write_index[1] ));
 sg13g2_dfrbp_1 _11528_ (.CLK(clknet_leaf_30_clk_regs),
    .RESET_B(net3590),
    .D(net881),
    .Q_N(_00057_),
    .Q(\core.lsu.write_index[2] ));
 sg13g2_dfrbp_1 _11529_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net3593),
    .D(net654),
    .Q_N(_05561_),
    .Q(\core.lsu.spi.counter[0] ));
 sg13g2_dfrbp_1 _11530_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net3593),
    .D(net408),
    .Q_N(_00127_),
    .Q(\core.lsu.spi.counter[1] ));
 sg13g2_dfrbp_1 _11531_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net3593),
    .D(net380),
    .Q_N(_00129_),
    .Q(\core.lsu.spi.counter[2] ));
 sg13g2_dfrbp_1 _11532_ (.CLK(clknet_leaf_35_clk_regs),
    .RESET_B(net3592),
    .D(net485),
    .Q_N(_00130_),
    .Q(\core.lsu.spi.counter[3] ));
 sg13g2_dfrbp_1 _11533_ (.CLK(clknet_leaf_33_clk_regs),
    .RESET_B(net3592),
    .D(net446),
    .Q_N(_00131_),
    .Q(\core.lsu.spi.counter[4] ));
 sg13g2_dfrbp_1 _11534_ (.CLK(clknet_leaf_32_clk_regs),
    .RESET_B(net3593),
    .D(net363),
    .Q_N(_00132_),
    .Q(\core.lsu.spi.counter[5] ));
 sg13g2_dfrbp_1 _11535_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net140),
    .D(net858),
    .Q_N(_05560_),
    .Q(\core.f2e_inst[0] ));
 sg13g2_dfrbp_1 _11536_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net139),
    .D(net845),
    .Q_N(_05559_),
    .Q(\core.f2e_inst[1] ));
 sg13g2_dfrbp_1 _11537_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net138),
    .D(net657),
    .Q_N(_00159_),
    .Q(\core.f2e_inst[2] ));
 sg13g2_dfrbp_1 _11538_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net137),
    .D(net659),
    .Q_N(_00160_),
    .Q(\core.f2e_inst[3] ));
 sg13g2_dfrbp_1 _11539_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net136),
    .D(_00423_),
    .Q_N(_00161_),
    .Q(\core.f2e_inst[4] ));
 sg13g2_dfrbp_1 _11540_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net135),
    .D(_00424_),
    .Q_N(_00162_),
    .Q(\core.f2e_inst[5] ));
 sg13g2_dfrbp_1 _11541_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net134),
    .D(net805),
    .Q_N(_00150_),
    .Q(\core.f2e_inst[6] ));
 sg13g2_dfrbp_1 _11542_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net133),
    .D(net707),
    .Q_N(_00155_),
    .Q(\core.f2e_inst[7] ));
 sg13g2_dfrbp_1 _11543_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net132),
    .D(_00427_),
    .Q_N(_00156_),
    .Q(\core.f2e_inst[8] ));
 sg13g2_dfrbp_1 _11544_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net131),
    .D(_00428_),
    .Q_N(_00157_),
    .Q(\core.f2e_inst[9] ));
 sg13g2_dfrbp_1 _11545_ (.CLK(clknet_leaf_5_clk_regs),
    .RESET_B(net130),
    .D(_00429_),
    .Q_N(_00158_),
    .Q(\core.f2e_inst[10] ));
 sg13g2_dfrbp_1 _11546_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net129),
    .D(_00430_),
    .Q_N(_00152_),
    .Q(\core.f2e_inst[11] ));
 sg13g2_dfrbp_1 _11547_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net128),
    .D(_00431_),
    .Q_N(_00149_),
    .Q(\core.f2e_inst[12] ));
 sg13g2_dfrbp_1 _11548_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net127),
    .D(_00432_),
    .Q_N(_05558_),
    .Q(\core.f2e_inst[13] ));
 sg13g2_dfrbp_1 _11549_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net126),
    .D(_00433_),
    .Q_N(_05557_),
    .Q(\core.f2e_inst[14] ));
 sg13g2_dfrbp_1 _11550_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net125),
    .D(_00434_),
    .Q_N(_00151_),
    .Q(\core.f2e_inst[15] ));
 sg13g2_dfrbp_1 _11551_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net124),
    .D(net474),
    .Q_N(_05556_),
    .Q(\core.f2e_inst[16] ));
 sg13g2_dfrbp_1 _11552_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net123),
    .D(net508),
    .Q_N(_05555_),
    .Q(\core.f2e_inst[17] ));
 sg13g2_dfrbp_1 _11553_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net122),
    .D(net451),
    .Q_N(_05554_),
    .Q(\core.f2e_inst[18] ));
 sg13g2_dfrbp_1 _11554_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net121),
    .D(net533),
    .Q_N(_05553_),
    .Q(\core.f2e_inst[19] ));
 sg13g2_dfrbp_1 _11555_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net120),
    .D(_00439_),
    .Q_N(_05552_),
    .Q(\core.f2e_inst[20] ));
 sg13g2_dfrbp_1 _11556_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net119),
    .D(net420),
    .Q_N(_05551_),
    .Q(\core.f2e_inst[21] ));
 sg13g2_dfrbp_1 _11557_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net118),
    .D(net538),
    .Q_N(_05550_),
    .Q(\core.f2e_inst[22] ));
 sg13g2_dfrbp_1 _11558_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net117),
    .D(net540),
    .Q_N(_05549_),
    .Q(\core.f2e_inst[23] ));
 sg13g2_dfrbp_1 _11559_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net116),
    .D(_00443_),
    .Q_N(_05548_),
    .Q(\core.f2e_inst[24] ));
 sg13g2_dfrbp_1 _11560_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net115),
    .D(net606),
    .Q_N(_05547_),
    .Q(\core.f2e_inst[25] ));
 sg13g2_dfrbp_1 _11561_ (.CLK(clknet_leaf_11_clk_regs),
    .RESET_B(net114),
    .D(net519),
    .Q_N(_05546_),
    .Q(\core.f2e_inst[26] ));
 sg13g2_dfrbp_1 _11562_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net113),
    .D(_00446_),
    .Q_N(_05545_),
    .Q(\core.f2e_inst[27] ));
 sg13g2_dfrbp_1 _11563_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net112),
    .D(net499),
    .Q_N(_05544_),
    .Q(\core.f2e_inst[28] ));
 sg13g2_dfrbp_1 _11564_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net111),
    .D(_00448_),
    .Q_N(_05543_),
    .Q(\core.f2e_inst[29] ));
 sg13g2_dfrbp_1 _11565_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net110),
    .D(net487),
    .Q_N(_05542_),
    .Q(\core.f2e_inst[30] ));
 sg13g2_dfrbp_1 _11566_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net109),
    .D(net449),
    .Q_N(_05541_),
    .Q(\core.f2e_inst[31] ));
 sg13g2_dfrbp_1 _11567_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net3586),
    .D(_00451_),
    .Q_N(_05540_),
    .Q(\core.f2e_addr[1] ));
 sg13g2_dfrbp_1 _11568_ (.CLK(clknet_leaf_34_clk_regs),
    .RESET_B(net108),
    .D(net503),
    .Q_N(_05539_),
    .Q(\core.lsu.spi.iswr ));
 sg13g2_dfrbp_1 _11569_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3595),
    .D(_00453_),
    .Q_N(_05538_),
    .Q(\core.work.state[0] ));
 sg13g2_dfrbp_1 _11570_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3582),
    .D(_00454_),
    .Q_N(_05537_),
    .Q(\core.work.state[1] ));
 sg13g2_dfrbp_1 _11571_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3582),
    .D(_00455_),
    .Q_N(_05536_),
    .Q(\core.work.dreg[0] ));
 sg13g2_dfrbp_1 _11572_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3582),
    .D(_00456_),
    .Q_N(_05535_),
    .Q(\core.work.dreg[1] ));
 sg13g2_dfrbp_1 _11573_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3582),
    .D(_00457_),
    .Q_N(_05534_),
    .Q(\core.work.dreg[2] ));
 sg13g2_dfrbp_1 _11574_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net3582),
    .D(_00458_),
    .Q_N(_05533_),
    .Q(\core.work.dreg[3] ));
 sg13g2_dfrbp_1 _11575_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net107),
    .D(_00459_),
    .Q_N(_05532_),
    .Q(\core.e2m_data[0] ));
 sg13g2_dfrbp_1 _11576_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net105),
    .D(_00460_),
    .Q_N(_05531_),
    .Q(\core.e2m_data[1] ));
 sg13g2_dfrbp_1 _11577_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net103),
    .D(_00461_),
    .Q_N(_05530_),
    .Q(\core.e2m_data[2] ));
 sg13g2_dfrbp_1 _11578_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net101),
    .D(_00462_),
    .Q_N(_05529_),
    .Q(\core.e2m_data[3] ));
 sg13g2_dfrbp_1 _11579_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net99),
    .D(_00463_),
    .Q_N(_05528_),
    .Q(\core.e2m_data[4] ));
 sg13g2_dfrbp_1 _11580_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net97),
    .D(_00464_),
    .Q_N(_05527_),
    .Q(\core.e2m_data[5] ));
 sg13g2_dfrbp_1 _11581_ (.CLK(clknet_leaf_42_clk_regs),
    .RESET_B(net95),
    .D(_00465_),
    .Q_N(_05526_),
    .Q(\core.e2m_data[6] ));
 sg13g2_dfrbp_1 _11582_ (.CLK(clknet_leaf_29_clk_regs),
    .RESET_B(net93),
    .D(_00466_),
    .Q_N(_05525_),
    .Q(\core.e2m_data[7] ));
 sg13g2_dfrbp_1 _11583_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net91),
    .D(_00467_),
    .Q_N(_05524_),
    .Q(\core.e2m_data[8] ));
 sg13g2_dfrbp_1 _11584_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net89),
    .D(_00468_),
    .Q_N(_05523_),
    .Q(\core.e2m_data[9] ));
 sg13g2_dfrbp_1 _11585_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net87),
    .D(_00469_),
    .Q_N(_05522_),
    .Q(\core.e2m_data[10] ));
 sg13g2_dfrbp_1 _11586_ (.CLK(clknet_leaf_28_clk_regs),
    .RESET_B(net85),
    .D(_00470_),
    .Q_N(_05521_),
    .Q(\core.e2m_data[11] ));
 sg13g2_dfrbp_1 _11587_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net83),
    .D(_00471_),
    .Q_N(_05520_),
    .Q(\core.e2m_data[12] ));
 sg13g2_dfrbp_1 _11588_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net82),
    .D(_00472_),
    .Q_N(_05519_),
    .Q(\core.e2m_data[13] ));
 sg13g2_dfrbp_1 _11589_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net81),
    .D(_00473_),
    .Q_N(_05518_),
    .Q(\core.e2m_data[14] ));
 sg13g2_dfrbp_1 _11590_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net80),
    .D(_00474_),
    .Q_N(_05517_),
    .Q(\core.e2m_data[15] ));
 sg13g2_dfrbp_1 _11591_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net78),
    .D(_00475_),
    .Q_N(_05516_),
    .Q(\core.e2m_data[16] ));
 sg13g2_dfrbp_1 _11592_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net76),
    .D(_00476_),
    .Q_N(_05515_),
    .Q(\core.e2m_data[17] ));
 sg13g2_dfrbp_1 _11593_ (.CLK(clknet_leaf_26_clk_regs),
    .RESET_B(net74),
    .D(_00477_),
    .Q_N(_05514_),
    .Q(\core.e2m_data[18] ));
 sg13g2_dfrbp_1 _11594_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net72),
    .D(_00478_),
    .Q_N(_05513_),
    .Q(\core.e2m_data[19] ));
 sg13g2_dfrbp_1 _11595_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net70),
    .D(_00479_),
    .Q_N(_05512_),
    .Q(\core.e2m_data[20] ));
 sg13g2_dfrbp_1 _11596_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net68),
    .D(_00480_),
    .Q_N(_05511_),
    .Q(\core.e2m_data[21] ));
 sg13g2_dfrbp_1 _11597_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net66),
    .D(_00481_),
    .Q_N(_05510_),
    .Q(\core.e2m_data[22] ));
 sg13g2_dfrbp_1 _11598_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net64),
    .D(_00482_),
    .Q_N(_05509_),
    .Q(\core.e2m_data[23] ));
 sg13g2_dfrbp_1 _11599_ (.CLK(clknet_leaf_27_clk_regs),
    .RESET_B(net62),
    .D(_00483_),
    .Q_N(_05508_),
    .Q(\core.e2m_data[24] ));
 sg13g2_dfrbp_1 _11600_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net60),
    .D(_00484_),
    .Q_N(_05507_),
    .Q(\core.e2m_data[25] ));
 sg13g2_dfrbp_1 _11601_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net58),
    .D(_00485_),
    .Q_N(_05506_),
    .Q(\core.e2m_data[26] ));
 sg13g2_dfrbp_1 _11602_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net56),
    .D(_00486_),
    .Q_N(_05505_),
    .Q(\core.e2m_data[27] ));
 sg13g2_dfrbp_1 _11603_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net54),
    .D(_00487_),
    .Q_N(_05504_),
    .Q(\core.e2m_data[28] ));
 sg13g2_dfrbp_1 _11604_ (.CLK(clknet_leaf_10_clk_regs),
    .RESET_B(net52),
    .D(_00488_),
    .Q_N(_05503_),
    .Q(\core.e2m_data[29] ));
 sg13g2_dfrbp_1 _11605_ (.CLK(clknet_leaf_9_clk_regs),
    .RESET_B(net50),
    .D(_00489_),
    .Q_N(_05502_),
    .Q(\core.e2m_data[30] ));
 sg13g2_dfrbp_1 _11606_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net48),
    .D(_00490_),
    .Q_N(_05501_),
    .Q(\core.e2m_data[31] ));
 sg13g2_dfrbp_1 _11607_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net3595),
    .D(_00491_),
    .Q_N(_00107_),
    .Q(\core.work.inst_was_short ));
 sg13g2_dfrbp_1 _11608_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net46),
    .D(_00492_),
    .Q_N(_00141_),
    .Q(\core.e2m_addr[0] ));
 sg13g2_dfrbp_1 _11609_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net45),
    .D(_00493_),
    .Q_N(_00145_),
    .Q(\core.e2m_addr[1] ));
 sg13g2_dfrbp_1 _11610_ (.CLK(clknet_leaf_39_clk_regs),
    .RESET_B(net44),
    .D(_00494_),
    .Q_N(_00147_),
    .Q(\core.e2m_addr[2] ));
 sg13g2_dfrbp_1 _11611_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net43),
    .D(_00495_),
    .Q_N(_00146_),
    .Q(\core.e2m_addr[3] ));
 sg13g2_dfrbp_1 _11612_ (.CLK(clknet_leaf_40_clk_regs),
    .RESET_B(net42),
    .D(_00496_),
    .Q_N(_00148_),
    .Q(\core.e2m_addr[4] ));
 sg13g2_dfrbp_1 _11613_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net41),
    .D(_00497_),
    .Q_N(_00153_),
    .Q(\core.e2m_addr[5] ));
 sg13g2_dfrbp_1 _11614_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net40),
    .D(net856),
    .Q_N(_00020_),
    .Q(\core.e2m_addr[6] ));
 sg13g2_dfrbp_1 _11615_ (.CLK(clknet_leaf_41_clk_regs),
    .RESET_B(net39),
    .D(_00499_),
    .Q_N(_00154_),
    .Q(\core.e2m_addr[7] ));
 sg13g2_dfrbp_1 _11616_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net38),
    .D(_00500_),
    .Q_N(_00106_),
    .Q(\core.e2m_addr[8] ));
 sg13g2_dfrbp_1 _11617_ (.CLK(clknet_leaf_43_clk_regs),
    .RESET_B(net37),
    .D(_00501_),
    .Q_N(_00108_),
    .Q(\core.e2m_addr[9] ));
 sg13g2_dfrbp_1 _11618_ (.CLK(clknet_4_11_0_clk_regs),
    .RESET_B(net36),
    .D(_00502_),
    .Q_N(_00110_),
    .Q(\core.e2m_addr[10] ));
 sg13g2_dfrbp_1 _11619_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net35),
    .D(_00503_),
    .Q_N(_00111_),
    .Q(\core.e2m_addr[11] ));
 sg13g2_dfrbp_1 _11620_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net34),
    .D(_00504_),
    .Q_N(_00120_),
    .Q(\core.e2m_addr[12] ));
 sg13g2_dfrbp_1 _11621_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net33),
    .D(_00505_),
    .Q_N(_00122_),
    .Q(\core.e2m_addr[13] ));
 sg13g2_dfrbp_1 _11622_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net32),
    .D(_00506_),
    .Q_N(_00124_),
    .Q(\core.e2m_addr[14] ));
 sg13g2_dfrbp_1 _11623_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net31),
    .D(_00507_),
    .Q_N(_00126_),
    .Q(\core.e2m_addr[15] ));
 sg13g2_dfrbp_1 _11624_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net30),
    .D(_00508_),
    .Q_N(_00023_),
    .Q(\core.e2m_addr[16] ));
 sg13g2_dfrbp_1 _11625_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net29),
    .D(_00509_),
    .Q_N(_00025_),
    .Q(\core.e2m_addr[17] ));
 sg13g2_dfrbp_1 _11626_ (.CLK(clknet_leaf_46_clk_regs),
    .RESET_B(net28),
    .D(_00510_),
    .Q_N(_00028_),
    .Q(\core.e2m_addr[18] ));
 sg13g2_dfrbp_1 _11627_ (.CLK(clknet_leaf_45_clk_regs),
    .RESET_B(net27),
    .D(_00511_),
    .Q_N(_00030_),
    .Q(\core.e2m_addr[19] ));
 sg13g2_dfrbp_1 _11628_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net26),
    .D(_00512_),
    .Q_N(_00032_),
    .Q(\core.e2m_addr[20] ));
 sg13g2_dfrbp_1 _11629_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net25),
    .D(_00513_),
    .Q_N(_00033_),
    .Q(\core.e2m_addr[21] ));
 sg13g2_dfrbp_1 _11630_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net24),
    .D(_00514_),
    .Q_N(_00036_),
    .Q(\core.e2m_addr[22] ));
 sg13g2_dfrbp_1 _11631_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net23),
    .D(_00515_),
    .Q_N(_00038_),
    .Q(\core.e2m_addr[23] ));
 sg13g2_dfrbp_1 _11632_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net22),
    .D(_00516_),
    .Q_N(_00040_),
    .Q(\core.e2m_addr[24] ));
 sg13g2_dfrbp_1 _11633_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net21),
    .D(_00517_),
    .Q_N(_00041_),
    .Q(\core.e2m_addr[25] ));
 sg13g2_dfrbp_1 _11634_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net20),
    .D(_00518_),
    .Q_N(_00044_),
    .Q(\core.e2m_addr[26] ));
 sg13g2_dfrbp_1 _11635_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net19),
    .D(_00519_),
    .Q_N(_00046_),
    .Q(\core.e2m_addr[27] ));
 sg13g2_dfrbp_1 _11636_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net18),
    .D(_00520_),
    .Q_N(_00048_),
    .Q(\core.e2m_addr[28] ));
 sg13g2_dfrbp_1 _11637_ (.CLK(clknet_leaf_52_clk_regs),
    .RESET_B(net17),
    .D(_00521_),
    .Q_N(_00049_),
    .Q(\core.e2m_addr[29] ));
 sg13g2_dfrbp_1 _11638_ (.CLK(clknet_leaf_51_clk_regs),
    .RESET_B(net16),
    .D(_00522_),
    .Q_N(_00052_),
    .Q(\core.e2m_addr[30] ));
 sg13g2_dfrbp_1 _11639_ (.CLK(clknet_leaf_6_clk_regs),
    .RESET_B(net15),
    .D(_00523_),
    .Q_N(_00024_),
    .Q(\core.e2m_addr[31] ));
 sg13g2_dfrbp_1 _11640_ (.CLK(net341),
    .RESET_B(net3579),
    .D(_00007_),
    .Q_N(_05500_),
    .Q(\core.work.registers.genblk1[14].we ));
 sg13g2_dfrbp_1 _11641_ (.CLK(net342),
    .RESET_B(net3579),
    .D(_00006_),
    .Q_N(_05499_),
    .Q(\core.work.registers.genblk1[13].we ));
 sg13g2_dlhq_1 _11642_ (.D(net3438),
    .GATE(net3253),
    .Q(\core.work.registers.genblk1[8].latch[0] ));
 sg13g2_dlhq_1 _11643_ (.D(net3436),
    .GATE(net3253),
    .Q(\core.work.registers.genblk1[8].latch[1] ));
 sg13g2_dlhq_1 _11644_ (.D(net3434),
    .GATE(net3253),
    .Q(\core.work.registers.genblk1[8].latch[2] ));
 sg13g2_dlhq_1 _11645_ (.D(net3432),
    .GATE(net3253),
    .Q(\core.work.registers.genblk1[8].latch[3] ));
 sg13g2_dlhq_1 _11646_ (.D(net3429),
    .GATE(net3253),
    .Q(\core.work.registers.genblk1[8].latch[4] ));
 sg13g2_dlhq_1 _11647_ (.D(net3428),
    .GATE(net3254),
    .Q(\core.work.registers.genblk1[8].latch[5] ));
 sg13g2_dlhq_1 _11648_ (.D(net3426),
    .GATE(net3253),
    .Q(\core.work.registers.genblk1[8].latch[6] ));
 sg13g2_dlhq_1 _11649_ (.D(net3423),
    .GATE(net3253),
    .Q(\core.work.registers.genblk1[8].latch[7] ));
 sg13g2_dlhq_1 _11650_ (.D(net3422),
    .GATE(net3254),
    .Q(\core.work.registers.genblk1[8].latch[8] ));
 sg13g2_dlhq_1 _11651_ (.D(net3419),
    .GATE(net3254),
    .Q(\core.work.registers.genblk1[8].latch[9] ));
 sg13g2_dlhq_1 _11652_ (.D(\core.work.registers.tmp[10] ),
    .GATE(net3252),
    .Q(\core.work.registers.genblk1[8].latch[10] ));
 sg13g2_dlhq_1 _11653_ (.D(net3414),
    .GATE(net3252),
    .Q(\core.work.registers.genblk1[8].latch[11] ));
 sg13g2_dlhq_1 _11654_ (.D(net3413),
    .GATE(net3254),
    .Q(\core.work.registers.genblk1[8].latch[12] ));
 sg13g2_dlhq_1 _11655_ (.D(net3411),
    .GATE(net3252),
    .Q(\core.work.registers.genblk1[8].latch[13] ));
 sg13g2_dlhq_1 _11656_ (.D(net3409),
    .GATE(net3252),
    .Q(\core.work.registers.genblk1[8].latch[14] ));
 sg13g2_dlhq_1 _11657_ (.D(net3405),
    .GATE(net3251),
    .Q(\core.work.registers.genblk1[8].latch[15] ));
 sg13g2_dlhq_1 _11658_ (.D(net3402),
    .GATE(net3254),
    .Q(\core.work.registers.genblk1[8].latch[16] ));
 sg13g2_dlhq_1 _11659_ (.D(net3401),
    .GATE(net3253),
    .Q(\core.work.registers.genblk1[8].latch[17] ));
 sg13g2_dlhq_1 _11660_ (.D(net3399),
    .GATE(net3254),
    .Q(\core.work.registers.genblk1[8].latch[18] ));
 sg13g2_dlhq_1 _11661_ (.D(net3395),
    .GATE(net3255),
    .Q(\core.work.registers.genblk1[8].latch[19] ));
 sg13g2_dlhq_1 _11662_ (.D(net3393),
    .GATE(net3254),
    .Q(\core.work.registers.genblk1[8].latch[20] ));
 sg13g2_dlhq_1 _11663_ (.D(net3390),
    .GATE(net3252),
    .Q(\core.work.registers.genblk1[8].latch[21] ));
 sg13g2_dlhq_1 _11664_ (.D(net3388),
    .GATE(net3252),
    .Q(\core.work.registers.genblk1[8].latch[22] ));
 sg13g2_dlhq_1 _11665_ (.D(net3385),
    .GATE(net3251),
    .Q(\core.work.registers.genblk1[8].latch[23] ));
 sg13g2_dlhq_1 _11666_ (.D(net3382),
    .GATE(net3254),
    .Q(\core.work.registers.genblk1[8].latch[24] ));
 sg13g2_dlhq_1 _11667_ (.D(net3379),
    .GATE(net3252),
    .Q(\core.work.registers.genblk1[8].latch[25] ));
 sg13g2_dlhq_1 _11668_ (.D(net3377),
    .GATE(net3251),
    .Q(\core.work.registers.genblk1[8].latch[26] ));
 sg13g2_dlhq_1 _11669_ (.D(net3376),
    .GATE(net3251),
    .Q(\core.work.registers.genblk1[8].latch[27] ));
 sg13g2_dlhq_1 _11670_ (.D(net3372),
    .GATE(net3251),
    .Q(\core.work.registers.genblk1[8].latch[28] ));
 sg13g2_dlhq_1 _11671_ (.D(net3369),
    .GATE(net3251),
    .Q(\core.work.registers.genblk1[8].latch[29] ));
 sg13g2_dlhq_1 _11672_ (.D(net3367),
    .GATE(net3251),
    .Q(\core.work.registers.genblk1[8].latch[30] ));
 sg13g2_dlhq_1 _11673_ (.D(net3363),
    .GATE(net3251),
    .Q(\core.work.registers.genblk1[8].latch[31] ));
 sg13g2_dlhq_1 _11674_ (.D(net3438),
    .GATE(net3228),
    .Q(\core.work.registers.genblk1[3].latch[0] ));
 sg13g2_dlhq_1 _11675_ (.D(net3436),
    .GATE(net3229),
    .Q(\core.work.registers.genblk1[3].latch[1] ));
 sg13g2_dlhq_1 _11676_ (.D(net3434),
    .GATE(net3228),
    .Q(\core.work.registers.genblk1[3].latch[2] ));
 sg13g2_dlhq_1 _11677_ (.D(net3433),
    .GATE(net3228),
    .Q(\core.work.registers.genblk1[3].latch[3] ));
 sg13g2_dlhq_1 _11678_ (.D(net3429),
    .GATE(net3228),
    .Q(\core.work.registers.genblk1[3].latch[4] ));
 sg13g2_dlhq_1 _11679_ (.D(net3428),
    .GATE(net3227),
    .Q(\core.work.registers.genblk1[3].latch[5] ));
 sg13g2_dlhq_1 _11680_ (.D(net3425),
    .GATE(net3228),
    .Q(\core.work.registers.genblk1[3].latch[6] ));
 sg13g2_dlhq_1 _11681_ (.D(net3424),
    .GATE(net3229),
    .Q(\core.work.registers.genblk1[3].latch[7] ));
 sg13g2_dlhq_1 _11682_ (.D(net3422),
    .GATE(net3230),
    .Q(\core.work.registers.genblk1[3].latch[8] ));
 sg13g2_dlhq_1 _11683_ (.D(net3420),
    .GATE(net3229),
    .Q(\core.work.registers.genblk1[3].latch[9] ));
 sg13g2_dlhq_1 _11684_ (.D(net3418),
    .GATE(net3230),
    .Q(\core.work.registers.genblk1[3].latch[10] ));
 sg13g2_dlhq_1 _11685_ (.D(net3415),
    .GATE(net3227),
    .Q(\core.work.registers.genblk1[3].latch[11] ));
 sg13g2_dlhq_1 _11686_ (.D(net3412),
    .GATE(net3227),
    .Q(\core.work.registers.genblk1[3].latch[12] ));
 sg13g2_dlhq_1 _11687_ (.D(net3410),
    .GATE(net3227),
    .Q(\core.work.registers.genblk1[3].latch[13] ));
 sg13g2_dlhq_1 _11688_ (.D(net3408),
    .GATE(net3230),
    .Q(\core.work.registers.genblk1[3].latch[14] ));
 sg13g2_dlhq_1 _11689_ (.D(net3405),
    .GATE(net3226),
    .Q(\core.work.registers.genblk1[3].latch[15] ));
 sg13g2_dlhq_1 _11690_ (.D(net3402),
    .GATE(net3229),
    .Q(\core.work.registers.genblk1[3].latch[16] ));
 sg13g2_dlhq_1 _11691_ (.D(net3401),
    .GATE(net3228),
    .Q(\core.work.registers.genblk1[3].latch[17] ));
 sg13g2_dlhq_1 _11692_ (.D(net3398),
    .GATE(net3229),
    .Q(\core.work.registers.genblk1[3].latch[18] ));
 sg13g2_dlhq_1 _11693_ (.D(net3395),
    .GATE(net3228),
    .Q(\core.work.registers.genblk1[3].latch[19] ));
 sg13g2_dlhq_1 _11694_ (.D(net3394),
    .GATE(net3228),
    .Q(\core.work.registers.genblk1[3].latch[20] ));
 sg13g2_dlhq_1 _11695_ (.D(net3391),
    .GATE(net3227),
    .Q(\core.work.registers.genblk1[3].latch[21] ));
 sg13g2_dlhq_1 _11696_ (.D(net3388),
    .GATE(net3227),
    .Q(\core.work.registers.genblk1[3].latch[22] ));
 sg13g2_dlhq_1 _11697_ (.D(net3387),
    .GATE(net3226),
    .Q(\core.work.registers.genblk1[3].latch[23] ));
 sg13g2_dlhq_1 _11698_ (.D(net3383),
    .GATE(net3229),
    .Q(\core.work.registers.genblk1[3].latch[24] ));
 sg13g2_dlhq_1 _11699_ (.D(net3379),
    .GATE(net3227),
    .Q(\core.work.registers.genblk1[3].latch[25] ));
 sg13g2_dlhq_1 _11700_ (.D(net3377),
    .GATE(net3226),
    .Q(\core.work.registers.genblk1[3].latch[26] ));
 sg13g2_dlhq_1 _11701_ (.D(net3375),
    .GATE(net3226),
    .Q(\core.work.registers.genblk1[3].latch[27] ));
 sg13g2_dlhq_1 _11702_ (.D(net3374),
    .GATE(net3226),
    .Q(\core.work.registers.genblk1[3].latch[28] ));
 sg13g2_dlhq_1 _11703_ (.D(net3371),
    .GATE(net3226),
    .Q(\core.work.registers.genblk1[3].latch[29] ));
 sg13g2_dlhq_1 _11704_ (.D(net3368),
    .GATE(net3226),
    .Q(\core.work.registers.genblk1[3].latch[30] ));
 sg13g2_dlhq_1 _11705_ (.D(net3364),
    .GATE(net3226),
    .Q(\core.work.registers.genblk1[3].latch[31] ));
 sg13g2_dfrbp_1 _11706_ (.CLK(net343),
    .RESET_B(net3579),
    .D(_00005_),
    .Q_N(_05498_),
    .Q(\core.work.registers.genblk1[12].we ));
 sg13g2_dlhq_1 _11707_ (.D(net3439),
    .GATE(net3259),
    .Q(\core.work.registers.genblk1[9].latch[0] ));
 sg13g2_dlhq_1 _11708_ (.D(net3437),
    .GATE(net3259),
    .Q(\core.work.registers.genblk1[9].latch[1] ));
 sg13g2_dlhq_1 _11709_ (.D(\core.work.registers.tmp[2] ),
    .GATE(net3259),
    .Q(\core.work.registers.genblk1[9].latch[2] ));
 sg13g2_dlhq_1 _11710_ (.D(net3433),
    .GATE(net3258),
    .Q(\core.work.registers.genblk1[9].latch[3] ));
 sg13g2_dlhq_1 _11711_ (.D(net3431),
    .GATE(net3259),
    .Q(\core.work.registers.genblk1[9].latch[4] ));
 sg13g2_dlhq_1 _11712_ (.D(net3428),
    .GATE(net3257),
    .Q(\core.work.registers.genblk1[9].latch[5] ));
 sg13g2_dlhq_1 _11713_ (.D(net3426),
    .GATE(net3259),
    .Q(\core.work.registers.genblk1[9].latch[6] ));
 sg13g2_dlhq_1 _11714_ (.D(net3423),
    .GATE(net3258),
    .Q(\core.work.registers.genblk1[9].latch[7] ));
 sg13g2_dlhq_1 _11715_ (.D(\core.work.registers.tmp[8] ),
    .GATE(net3257),
    .Q(\core.work.registers.genblk1[9].latch[8] ));
 sg13g2_dlhq_1 _11716_ (.D(net3419),
    .GATE(net3258),
    .Q(\core.work.registers.genblk1[9].latch[9] ));
 sg13g2_dlhq_1 _11717_ (.D(net3418),
    .GATE(net3260),
    .Q(\core.work.registers.genblk1[9].latch[10] ));
 sg13g2_dlhq_1 _11718_ (.D(net3414),
    .GATE(net3257),
    .Q(\core.work.registers.genblk1[9].latch[11] ));
 sg13g2_dlhq_1 _11719_ (.D(net3412),
    .GATE(net3257),
    .Q(\core.work.registers.genblk1[9].latch[12] ));
 sg13g2_dlhq_1 _11720_ (.D(net3410),
    .GATE(net3257),
    .Q(\core.work.registers.genblk1[9].latch[13] ));
 sg13g2_dlhq_1 _11721_ (.D(net3409),
    .GATE(net3260),
    .Q(\core.work.registers.genblk1[9].latch[14] ));
 sg13g2_dlhq_1 _11722_ (.D(net3406),
    .GATE(net3256),
    .Q(\core.work.registers.genblk1[9].latch[15] ));
 sg13g2_dlhq_1 _11723_ (.D(net3403),
    .GATE(net3258),
    .Q(\core.work.registers.genblk1[9].latch[16] ));
 sg13g2_dlhq_1 _11724_ (.D(net3400),
    .GATE(net3258),
    .Q(\core.work.registers.genblk1[9].latch[17] ));
 sg13g2_dlhq_1 _11725_ (.D(net3399),
    .GATE(net3258),
    .Q(\core.work.registers.genblk1[9].latch[18] ));
 sg13g2_dlhq_1 _11726_ (.D(net3397),
    .GATE(net3259),
    .Q(\core.work.registers.genblk1[9].latch[19] ));
 sg13g2_dlhq_1 _11727_ (.D(net3393),
    .GATE(net3258),
    .Q(\core.work.registers.genblk1[9].latch[20] ));
 sg13g2_dlhq_1 _11728_ (.D(net3392),
    .GATE(net3257),
    .Q(\core.work.registers.genblk1[9].latch[21] ));
 sg13g2_dlhq_1 _11729_ (.D(net3388),
    .GATE(net3257),
    .Q(\core.work.registers.genblk1[9].latch[22] ));
 sg13g2_dlhq_1 _11730_ (.D(net3385),
    .GATE(net3256),
    .Q(\core.work.registers.genblk1[9].latch[23] ));
 sg13g2_dlhq_1 _11731_ (.D(net3382),
    .GATE(net3258),
    .Q(\core.work.registers.genblk1[9].latch[24] ));
 sg13g2_dlhq_1 _11732_ (.D(net3379),
    .GATE(net3260),
    .Q(\core.work.registers.genblk1[9].latch[25] ));
 sg13g2_dlhq_1 _11733_ (.D(net3377),
    .GATE(net3256),
    .Q(\core.work.registers.genblk1[9].latch[26] ));
 sg13g2_dlhq_1 _11734_ (.D(net3376),
    .GATE(net3256),
    .Q(\core.work.registers.genblk1[9].latch[27] ));
 sg13g2_dlhq_1 _11735_ (.D(net3372),
    .GATE(net3256),
    .Q(\core.work.registers.genblk1[9].latch[28] ));
 sg13g2_dlhq_1 _11736_ (.D(net3369),
    .GATE(net3256),
    .Q(\core.work.registers.genblk1[9].latch[29] ));
 sg13g2_dlhq_1 _11737_ (.D(net3366),
    .GATE(net3256),
    .Q(\core.work.registers.genblk1[9].latch[30] ));
 sg13g2_dlhq_1 _11738_ (.D(net3363),
    .GATE(net3256),
    .Q(\core.work.registers.genblk1[9].latch[31] ));
 sg13g2_dfrbp_1 _11739_ (.CLK(net344),
    .RESET_B(net3579),
    .D(_00004_),
    .Q_N(_05497_),
    .Q(\core.work.registers.genblk1[11].we ));
 sg13g2_dlhq_1 _11740_ (.D(net3438),
    .GATE(net3239),
    .Q(\core.work.registers.genblk1[5].latch[0] ));
 sg13g2_dlhq_1 _11741_ (.D(net3436),
    .GATE(net3239),
    .Q(\core.work.registers.genblk1[5].latch[1] ));
 sg13g2_dlhq_1 _11742_ (.D(net3434),
    .GATE(net3239),
    .Q(\core.work.registers.genblk1[5].latch[2] ));
 sg13g2_dlhq_1 _11743_ (.D(net3432),
    .GATE(net3239),
    .Q(\core.work.registers.genblk1[5].latch[3] ));
 sg13g2_dlhq_1 _11744_ (.D(net3430),
    .GATE(net3239),
    .Q(\core.work.registers.genblk1[5].latch[4] ));
 sg13g2_dlhq_1 _11745_ (.D(net3427),
    .GATE(net3237),
    .Q(\core.work.registers.genblk1[5].latch[5] ));
 sg13g2_dlhq_1 _11746_ (.D(net3425),
    .GATE(net3239),
    .Q(\core.work.registers.genblk1[5].latch[6] ));
 sg13g2_dlhq_1 _11747_ (.D(net3424),
    .GATE(net3238),
    .Q(\core.work.registers.genblk1[5].latch[7] ));
 sg13g2_dlhq_1 _11748_ (.D(net3421),
    .GATE(net3237),
    .Q(\core.work.registers.genblk1[5].latch[8] ));
 sg13g2_dlhq_1 _11749_ (.D(net3420),
    .GATE(net3238),
    .Q(\core.work.registers.genblk1[5].latch[9] ));
 sg13g2_dlhq_1 _11750_ (.D(net3417),
    .GATE(net3240),
    .Q(\core.work.registers.genblk1[5].latch[10] ));
 sg13g2_dlhq_1 _11751_ (.D(net3414),
    .GATE(net3237),
    .Q(\core.work.registers.genblk1[5].latch[11] ));
 sg13g2_dlhq_1 _11752_ (.D(net3413),
    .GATE(net3238),
    .Q(\core.work.registers.genblk1[5].latch[12] ));
 sg13g2_dlhq_1 _11753_ (.D(net3410),
    .GATE(net3237),
    .Q(\core.work.registers.genblk1[5].latch[13] ));
 sg13g2_dlhq_1 _11754_ (.D(net3409),
    .GATE(net3240),
    .Q(\core.work.registers.genblk1[5].latch[14] ));
 sg13g2_dlhq_1 _11755_ (.D(net3405),
    .GATE(net3236),
    .Q(\core.work.registers.genblk1[5].latch[15] ));
 sg13g2_dlhq_1 _11756_ (.D(net3403),
    .GATE(net3238),
    .Q(\core.work.registers.genblk1[5].latch[16] ));
 sg13g2_dlhq_1 _11757_ (.D(net3400),
    .GATE(net3238),
    .Q(\core.work.registers.genblk1[5].latch[17] ));
 sg13g2_dlhq_1 _11758_ (.D(net3398),
    .GATE(net3238),
    .Q(\core.work.registers.genblk1[5].latch[18] ));
 sg13g2_dlhq_1 _11759_ (.D(net3395),
    .GATE(net3239),
    .Q(\core.work.registers.genblk1[5].latch[19] ));
 sg13g2_dlhq_1 _11760_ (.D(net3393),
    .GATE(net3238),
    .Q(\core.work.registers.genblk1[5].latch[20] ));
 sg13g2_dlhq_1 _11761_ (.D(net3390),
    .GATE(net3237),
    .Q(\core.work.registers.genblk1[5].latch[21] ));
 sg13g2_dlhq_1 _11762_ (.D(net3388),
    .GATE(net3237),
    .Q(\core.work.registers.genblk1[5].latch[22] ));
 sg13g2_dlhq_1 _11763_ (.D(net3385),
    .GATE(net3236),
    .Q(\core.work.registers.genblk1[5].latch[23] ));
 sg13g2_dlhq_1 _11764_ (.D(net3384),
    .GATE(net3238),
    .Q(\core.work.registers.genblk1[5].latch[24] ));
 sg13g2_dlhq_1 _11765_ (.D(net3379),
    .GATE(net3237),
    .Q(\core.work.registers.genblk1[5].latch[25] ));
 sg13g2_dlhq_1 _11766_ (.D(net3378),
    .GATE(net3236),
    .Q(\core.work.registers.genblk1[5].latch[26] ));
 sg13g2_dlhq_1 _11767_ (.D(net3375),
    .GATE(net3236),
    .Q(\core.work.registers.genblk1[5].latch[27] ));
 sg13g2_dlhq_1 _11768_ (.D(net3372),
    .GATE(net3236),
    .Q(\core.work.registers.genblk1[5].latch[28] ));
 sg13g2_dlhq_1 _11769_ (.D(net3370),
    .GATE(net3236),
    .Q(\core.work.registers.genblk1[5].latch[29] ));
 sg13g2_dlhq_1 _11770_ (.D(net3367),
    .GATE(net3236),
    .Q(\core.work.registers.genblk1[5].latch[30] ));
 sg13g2_dlhq_1 _11771_ (.D(net3364),
    .GATE(net3236),
    .Q(\core.work.registers.genblk1[5].latch[31] ));
 sg13g2_dlhq_1 _11772_ (.D(net3439),
    .GATE(net3264),
    .Q(\core.work.registers.genblk1[10].latch[0] ));
 sg13g2_dlhq_1 _11773_ (.D(net3437),
    .GATE(net3264),
    .Q(\core.work.registers.genblk1[10].latch[1] ));
 sg13g2_dlhq_1 _11774_ (.D(net3435),
    .GATE(net3264),
    .Q(\core.work.registers.genblk1[10].latch[2] ));
 sg13g2_dlhq_1 _11775_ (.D(net3432),
    .GATE(net3263),
    .Q(\core.work.registers.genblk1[10].latch[3] ));
 sg13g2_dlhq_1 _11776_ (.D(net3431),
    .GATE(net3264),
    .Q(\core.work.registers.genblk1[10].latch[4] ));
 sg13g2_dlhq_1 _11777_ (.D(net3428),
    .GATE(net3262),
    .Q(\core.work.registers.genblk1[10].latch[5] ));
 sg13g2_dlhq_1 _11778_ (.D(net3426),
    .GATE(net3264),
    .Q(\core.work.registers.genblk1[10].latch[6] ));
 sg13g2_dlhq_1 _11779_ (.D(net3424),
    .GATE(net3263),
    .Q(\core.work.registers.genblk1[10].latch[7] ));
 sg13g2_dlhq_1 _11780_ (.D(net3422),
    .GATE(net3265),
    .Q(\core.work.registers.genblk1[10].latch[8] ));
 sg13g2_dlhq_1 _11781_ (.D(net3420),
    .GATE(net3263),
    .Q(\core.work.registers.genblk1[10].latch[9] ));
 sg13g2_dlhq_1 _11782_ (.D(net3417),
    .GATE(net3265),
    .Q(\core.work.registers.genblk1[10].latch[10] ));
 sg13g2_dlhq_1 _11783_ (.D(net3414),
    .GATE(net3262),
    .Q(\core.work.registers.genblk1[10].latch[11] ));
 sg13g2_dlhq_1 _11784_ (.D(net3412),
    .GATE(net3262),
    .Q(\core.work.registers.genblk1[10].latch[12] ));
 sg13g2_dlhq_1 _11785_ (.D(net3410),
    .GATE(net3262),
    .Q(\core.work.registers.genblk1[10].latch[13] ));
 sg13g2_dlhq_1 _11786_ (.D(net3408),
    .GATE(net3265),
    .Q(\core.work.registers.genblk1[10].latch[14] ));
 sg13g2_dlhq_1 _11787_ (.D(net3406),
    .GATE(net3261),
    .Q(\core.work.registers.genblk1[10].latch[15] ));
 sg13g2_dlhq_1 _11788_ (.D(net3403),
    .GATE(net3263),
    .Q(\core.work.registers.genblk1[10].latch[16] ));
 sg13g2_dlhq_1 _11789_ (.D(net3401),
    .GATE(net3263),
    .Q(\core.work.registers.genblk1[10].latch[17] ));
 sg13g2_dlhq_1 _11790_ (.D(net3399),
    .GATE(net3263),
    .Q(\core.work.registers.genblk1[10].latch[18] ));
 sg13g2_dlhq_1 _11791_ (.D(net3397),
    .GATE(net3264),
    .Q(\core.work.registers.genblk1[10].latch[19] ));
 sg13g2_dlhq_1 _11792_ (.D(net3393),
    .GATE(net3263),
    .Q(\core.work.registers.genblk1[10].latch[20] ));
 sg13g2_dlhq_1 _11793_ (.D(net3390),
    .GATE(net3262),
    .Q(\core.work.registers.genblk1[10].latch[21] ));
 sg13g2_dlhq_1 _11794_ (.D(net3389),
    .GATE(net3262),
    .Q(\core.work.registers.genblk1[10].latch[22] ));
 sg13g2_dlhq_1 _11795_ (.D(net3386),
    .GATE(net3261),
    .Q(\core.work.registers.genblk1[10].latch[23] ));
 sg13g2_dlhq_1 _11796_ (.D(net3383),
    .GATE(net3263),
    .Q(\core.work.registers.genblk1[10].latch[24] ));
 sg13g2_dlhq_1 _11797_ (.D(net3380),
    .GATE(net3262),
    .Q(\core.work.registers.genblk1[10].latch[25] ));
 sg13g2_dlhq_1 _11798_ (.D(net3378),
    .GATE(net3261),
    .Q(\core.work.registers.genblk1[10].latch[26] ));
 sg13g2_dlhq_1 _11799_ (.D(net3376),
    .GATE(net3261),
    .Q(\core.work.registers.genblk1[10].latch[27] ));
 sg13g2_dlhq_1 _11800_ (.D(net3372),
    .GATE(net3261),
    .Q(\core.work.registers.genblk1[10].latch[28] ));
 sg13g2_dlhq_1 _11801_ (.D(net3369),
    .GATE(net3261),
    .Q(\core.work.registers.genblk1[10].latch[29] ));
 sg13g2_dlhq_1 _11802_ (.D(net3366),
    .GATE(net3261),
    .Q(\core.work.registers.genblk1[10].latch[30] ));
 sg13g2_dlhq_1 _11803_ (.D(net3363),
    .GATE(net3261),
    .Q(\core.work.registers.genblk1[10].latch[31] ));
 sg13g2_dfrbp_1 _11804_ (.CLK(net345),
    .RESET_B(net3579),
    .D(_00003_),
    .Q_N(_05496_),
    .Q(\core.work.registers.genblk1[10].we ));
 sg13g2_dfrbp_1 _11805_ (.CLK(net346),
    .RESET_B(net3580),
    .D(_00017_),
    .Q_N(_05495_),
    .Q(\core.work.registers.genblk1[9].we ));
 sg13g2_dlhq_1 _11806_ (.D(net3438),
    .GATE(net3268),
    .Q(\core.work.registers.genblk1[11].latch[0] ));
 sg13g2_dlhq_1 _11807_ (.D(net3437),
    .GATE(net3268),
    .Q(\core.work.registers.genblk1[11].latch[1] ));
 sg13g2_dlhq_1 _11808_ (.D(net3434),
    .GATE(net3268),
    .Q(\core.work.registers.genblk1[11].latch[2] ));
 sg13g2_dlhq_1 _11809_ (.D(net3433),
    .GATE(net3268),
    .Q(\core.work.registers.genblk1[11].latch[3] ));
 sg13g2_dlhq_1 _11810_ (.D(net3429),
    .GATE(net3268),
    .Q(\core.work.registers.genblk1[11].latch[4] ));
 sg13g2_dlhq_1 _11811_ (.D(net3427),
    .GATE(net3267),
    .Q(\core.work.registers.genblk1[11].latch[5] ));
 sg13g2_dlhq_1 _11812_ (.D(net3425),
    .GATE(net3269),
    .Q(\core.work.registers.genblk1[11].latch[6] ));
 sg13g2_dlhq_1 _11813_ (.D(net3423),
    .GATE(net3268),
    .Q(\core.work.registers.genblk1[11].latch[7] ));
 sg13g2_dlhq_1 _11814_ (.D(net3421),
    .GATE(net3270),
    .Q(\core.work.registers.genblk1[11].latch[8] ));
 sg13g2_dlhq_1 _11815_ (.D(net3420),
    .GATE(net3269),
    .Q(\core.work.registers.genblk1[11].latch[9] ));
 sg13g2_dlhq_1 _11816_ (.D(net3417),
    .GATE(net3270),
    .Q(\core.work.registers.genblk1[11].latch[10] ));
 sg13g2_dlhq_1 _11817_ (.D(net3415),
    .GATE(net3267),
    .Q(\core.work.registers.genblk1[11].latch[11] ));
 sg13g2_dlhq_1 _11818_ (.D(net3412),
    .GATE(net3267),
    .Q(\core.work.registers.genblk1[11].latch[12] ));
 sg13g2_dlhq_1 _11819_ (.D(net3411),
    .GATE(net3267),
    .Q(\core.work.registers.genblk1[11].latch[13] ));
 sg13g2_dlhq_1 _11820_ (.D(\core.work.registers.tmp[14] ),
    .GATE(net3270),
    .Q(\core.work.registers.genblk1[11].latch[14] ));
 sg13g2_dlhq_1 _11821_ (.D(net3405),
    .GATE(net3266),
    .Q(\core.work.registers.genblk1[11].latch[15] ));
 sg13g2_dlhq_1 _11822_ (.D(net3402),
    .GATE(net3269),
    .Q(\core.work.registers.genblk1[11].latch[16] ));
 sg13g2_dlhq_1 _11823_ (.D(net3400),
    .GATE(net3268),
    .Q(\core.work.registers.genblk1[11].latch[17] ));
 sg13g2_dlhq_1 _11824_ (.D(net3398),
    .GATE(net3269),
    .Q(\core.work.registers.genblk1[11].latch[18] ));
 sg13g2_dlhq_1 _11825_ (.D(net3395),
    .GATE(net3268),
    .Q(\core.work.registers.genblk1[11].latch[19] ));
 sg13g2_dlhq_1 _11826_ (.D(net3394),
    .GATE(net3269),
    .Q(\core.work.registers.genblk1[11].latch[20] ));
 sg13g2_dlhq_1 _11827_ (.D(net3391),
    .GATE(net3267),
    .Q(\core.work.registers.genblk1[11].latch[21] ));
 sg13g2_dlhq_1 _11828_ (.D(net3389),
    .GATE(net3267),
    .Q(\core.work.registers.genblk1[11].latch[22] ));
 sg13g2_dlhq_1 _11829_ (.D(net3385),
    .GATE(net3266),
    .Q(\core.work.registers.genblk1[11].latch[23] ));
 sg13g2_dlhq_1 _11830_ (.D(net3382),
    .GATE(net3269),
    .Q(\core.work.registers.genblk1[11].latch[24] ));
 sg13g2_dlhq_1 _11831_ (.D(net3380),
    .GATE(net3267),
    .Q(\core.work.registers.genblk1[11].latch[25] ));
 sg13g2_dlhq_1 _11832_ (.D(net3377),
    .GATE(net3266),
    .Q(\core.work.registers.genblk1[11].latch[26] ));
 sg13g2_dlhq_1 _11833_ (.D(net3375),
    .GATE(net3266),
    .Q(\core.work.registers.genblk1[11].latch[27] ));
 sg13g2_dlhq_1 _11834_ (.D(net3373),
    .GATE(net3266),
    .Q(\core.work.registers.genblk1[11].latch[28] ));
 sg13g2_dlhq_1 _11835_ (.D(net3369),
    .GATE(net3266),
    .Q(\core.work.registers.genblk1[11].latch[29] ));
 sg13g2_dlhq_1 _11836_ (.D(net3366),
    .GATE(net3266),
    .Q(\core.work.registers.genblk1[11].latch[30] ));
 sg13g2_dlhq_1 _11837_ (.D(net3363),
    .GATE(net3266),
    .Q(\core.work.registers.genblk1[11].latch[31] ));
 sg13g2_dlhq_1 _11838_ (.D(net3439),
    .GATE(net3234),
    .Q(\core.work.registers.genblk1[4].latch[0] ));
 sg13g2_dlhq_1 _11839_ (.D(net3436),
    .GATE(net3234),
    .Q(\core.work.registers.genblk1[4].latch[1] ));
 sg13g2_dlhq_1 _11840_ (.D(net3435),
    .GATE(net3234),
    .Q(\core.work.registers.genblk1[4].latch[2] ));
 sg13g2_dlhq_1 _11841_ (.D(net3432),
    .GATE(net3234),
    .Q(\core.work.registers.genblk1[4].latch[3] ));
 sg13g2_dlhq_1 _11842_ (.D(net3429),
    .GATE(net3233),
    .Q(\core.work.registers.genblk1[4].latch[4] ));
 sg13g2_dlhq_1 _11843_ (.D(net3427),
    .GATE(net3232),
    .Q(\core.work.registers.genblk1[4].latch[5] ));
 sg13g2_dlhq_1 _11844_ (.D(net3425),
    .GATE(net3234),
    .Q(\core.work.registers.genblk1[4].latch[6] ));
 sg13g2_dlhq_1 _11845_ (.D(net3424),
    .GATE(net3233),
    .Q(\core.work.registers.genblk1[4].latch[7] ));
 sg13g2_dlhq_1 _11846_ (.D(net3421),
    .GATE(net3235),
    .Q(\core.work.registers.genblk1[4].latch[8] ));
 sg13g2_dlhq_1 _11847_ (.D(net3419),
    .GATE(net3233),
    .Q(\core.work.registers.genblk1[4].latch[9] ));
 sg13g2_dlhq_1 _11848_ (.D(net3418),
    .GATE(net3235),
    .Q(\core.work.registers.genblk1[4].latch[10] ));
 sg13g2_dlhq_1 _11849_ (.D(net3414),
    .GATE(net3231),
    .Q(\core.work.registers.genblk1[4].latch[11] ));
 sg13g2_dlhq_1 _11850_ (.D(net3413),
    .GATE(net3232),
    .Q(\core.work.registers.genblk1[4].latch[12] ));
 sg13g2_dlhq_1 _11851_ (.D(net3411),
    .GATE(net3232),
    .Q(\core.work.registers.genblk1[4].latch[13] ));
 sg13g2_dlhq_1 _11852_ (.D(net3408),
    .GATE(net3235),
    .Q(\core.work.registers.genblk1[4].latch[14] ));
 sg13g2_dlhq_1 _11853_ (.D(net3406),
    .GATE(net3231),
    .Q(\core.work.registers.genblk1[4].latch[15] ));
 sg13g2_dlhq_1 _11854_ (.D(net3402),
    .GATE(net3233),
    .Q(\core.work.registers.genblk1[4].latch[16] ));
 sg13g2_dlhq_1 _11855_ (.D(net3401),
    .GATE(net3233),
    .Q(\core.work.registers.genblk1[4].latch[17] ));
 sg13g2_dlhq_1 _11856_ (.D(net3399),
    .GATE(net3233),
    .Q(\core.work.registers.genblk1[4].latch[18] ));
 sg13g2_dlhq_1 _11857_ (.D(net3396),
    .GATE(net3234),
    .Q(\core.work.registers.genblk1[4].latch[19] ));
 sg13g2_dlhq_1 _11858_ (.D(net3394),
    .GATE(net3233),
    .Q(\core.work.registers.genblk1[4].latch[20] ));
 sg13g2_dlhq_1 _11859_ (.D(net3390),
    .GATE(net3232),
    .Q(\core.work.registers.genblk1[4].latch[21] ));
 sg13g2_dlhq_1 _11860_ (.D(net3389),
    .GATE(net3232),
    .Q(\core.work.registers.genblk1[4].latch[22] ));
 sg13g2_dlhq_1 _11861_ (.D(net3387),
    .GATE(net3231),
    .Q(\core.work.registers.genblk1[4].latch[23] ));
 sg13g2_dlhq_1 _11862_ (.D(net3382),
    .GATE(net3233),
    .Q(\core.work.registers.genblk1[4].latch[24] ));
 sg13g2_dlhq_1 _11863_ (.D(net3381),
    .GATE(net3232),
    .Q(\core.work.registers.genblk1[4].latch[25] ));
 sg13g2_dlhq_1 _11864_ (.D(net3378),
    .GATE(net3231),
    .Q(\core.work.registers.genblk1[4].latch[26] ));
 sg13g2_dlhq_1 _11865_ (.D(net3376),
    .GATE(net3232),
    .Q(\core.work.registers.genblk1[4].latch[27] ));
 sg13g2_dlhq_1 _11866_ (.D(net3374),
    .GATE(net3231),
    .Q(\core.work.registers.genblk1[4].latch[28] ));
 sg13g2_dlhq_1 _11867_ (.D(net3371),
    .GATE(net3231),
    .Q(\core.work.registers.genblk1[4].latch[29] ));
 sg13g2_dlhq_1 _11868_ (.D(net3368),
    .GATE(net3231),
    .Q(\core.work.registers.genblk1[4].latch[30] ));
 sg13g2_dlhq_1 _11869_ (.D(net3364),
    .GATE(net3231),
    .Q(\core.work.registers.genblk1[4].latch[31] ));
 sg13g2_dfrbp_1 _11870_ (.CLK(net347),
    .RESET_B(net3579),
    .D(_00016_),
    .Q_N(_05494_),
    .Q(\core.work.registers.genblk1[8].we ));
 sg13g2_dlhq_1 _11871_ (.D(net3438),
    .GATE(net3273),
    .Q(\core.work.registers.genblk1[12].latch[0] ));
 sg13g2_dlhq_1 _11872_ (.D(net3436),
    .GATE(net3273),
    .Q(\core.work.registers.genblk1[12].latch[1] ));
 sg13g2_dlhq_1 _11873_ (.D(net3434),
    .GATE(net3273),
    .Q(\core.work.registers.genblk1[12].latch[2] ));
 sg13g2_dlhq_1 _11874_ (.D(net3433),
    .GATE(net3273),
    .Q(\core.work.registers.genblk1[12].latch[3] ));
 sg13g2_dlhq_1 _11875_ (.D(net3429),
    .GATE(net3273),
    .Q(\core.work.registers.genblk1[12].latch[4] ));
 sg13g2_dlhq_1 _11876_ (.D(net3427),
    .GATE(net3272),
    .Q(\core.work.registers.genblk1[12].latch[5] ));
 sg13g2_dlhq_1 _11877_ (.D(net3426),
    .GATE(net3275),
    .Q(\core.work.registers.genblk1[12].latch[6] ));
 sg13g2_dlhq_1 _11878_ (.D(net3424),
    .GATE(net3274),
    .Q(\core.work.registers.genblk1[12].latch[7] ));
 sg13g2_dlhq_1 _11879_ (.D(net3421),
    .GATE(net3274),
    .Q(\core.work.registers.genblk1[12].latch[8] ));
 sg13g2_dlhq_1 _11880_ (.D(net3420),
    .GATE(net3274),
    .Q(\core.work.registers.genblk1[12].latch[9] ));
 sg13g2_dlhq_1 _11881_ (.D(net3417),
    .GATE(net3272),
    .Q(\core.work.registers.genblk1[12].latch[10] ));
 sg13g2_dlhq_1 _11882_ (.D(net3415),
    .GATE(net3271),
    .Q(\core.work.registers.genblk1[12].latch[11] ));
 sg13g2_dlhq_1 _11883_ (.D(net3413),
    .GATE(net3274),
    .Q(\core.work.registers.genblk1[12].latch[12] ));
 sg13g2_dlhq_1 _11884_ (.D(net3411),
    .GATE(net3272),
    .Q(\core.work.registers.genblk1[12].latch[13] ));
 sg13g2_dlhq_1 _11885_ (.D(net3408),
    .GATE(net3275),
    .Q(\core.work.registers.genblk1[12].latch[14] ));
 sg13g2_dlhq_1 _11886_ (.D(net3405),
    .GATE(net3271),
    .Q(\core.work.registers.genblk1[12].latch[15] ));
 sg13g2_dlhq_1 _11887_ (.D(net3403),
    .GATE(net3274),
    .Q(\core.work.registers.genblk1[12].latch[16] ));
 sg13g2_dlhq_1 _11888_ (.D(net3401),
    .GATE(net3273),
    .Q(\core.work.registers.genblk1[12].latch[17] ));
 sg13g2_dlhq_1 _11889_ (.D(net3399),
    .GATE(net3274),
    .Q(\core.work.registers.genblk1[12].latch[18] ));
 sg13g2_dlhq_1 _11890_ (.D(net3396),
    .GATE(net3273),
    .Q(\core.work.registers.genblk1[12].latch[19] ));
 sg13g2_dlhq_1 _11891_ (.D(net3393),
    .GATE(net3273),
    .Q(\core.work.registers.genblk1[12].latch[20] ));
 sg13g2_dlhq_1 _11892_ (.D(net3391),
    .GATE(net3272),
    .Q(\core.work.registers.genblk1[12].latch[21] ));
 sg13g2_dlhq_1 _11893_ (.D(net3388),
    .GATE(net3272),
    .Q(\core.work.registers.genblk1[12].latch[22] ));
 sg13g2_dlhq_1 _11894_ (.D(net3385),
    .GATE(net3271),
    .Q(\core.work.registers.genblk1[12].latch[23] ));
 sg13g2_dlhq_1 _11895_ (.D(net3382),
    .GATE(net3274),
    .Q(\core.work.registers.genblk1[12].latch[24] ));
 sg13g2_dlhq_1 _11896_ (.D(net3379),
    .GATE(net3272),
    .Q(\core.work.registers.genblk1[12].latch[25] ));
 sg13g2_dlhq_1 _11897_ (.D(net3378),
    .GATE(net3271),
    .Q(\core.work.registers.genblk1[12].latch[26] ));
 sg13g2_dlhq_1 _11898_ (.D(net3376),
    .GATE(net3272),
    .Q(\core.work.registers.genblk1[12].latch[27] ));
 sg13g2_dlhq_1 _11899_ (.D(net3372),
    .GATE(net3271),
    .Q(\core.work.registers.genblk1[12].latch[28] ));
 sg13g2_dlhq_1 _11900_ (.D(net3369),
    .GATE(net3271),
    .Q(\core.work.registers.genblk1[12].latch[29] ));
 sg13g2_dlhq_1 _11901_ (.D(net3366),
    .GATE(net3271),
    .Q(\core.work.registers.genblk1[12].latch[30] ));
 sg13g2_dlhq_1 _11902_ (.D(net3364),
    .GATE(net3271),
    .Q(\core.work.registers.genblk1[12].latch[31] ));
 sg13g2_dlhq_1 _11903_ (.D(net3438),
    .GATE(net3213),
    .Q(\core.work.registers.genblk1[1].latch[0] ));
 sg13g2_dlhq_1 _11904_ (.D(net3436),
    .GATE(net3213),
    .Q(\core.work.registers.genblk1[1].latch[1] ));
 sg13g2_dlhq_1 _11905_ (.D(net3434),
    .GATE(net3213),
    .Q(\core.work.registers.genblk1[1].latch[2] ));
 sg13g2_dlhq_1 _11906_ (.D(\core.work.registers.tmp[3] ),
    .GATE(net3213),
    .Q(\core.work.registers.genblk1[1].latch[3] ));
 sg13g2_dlhq_1 _11907_ (.D(net3431),
    .GATE(net3213),
    .Q(\core.work.registers.genblk1[1].latch[4] ));
 sg13g2_dlhq_1 _11908_ (.D(\core.work.registers.tmp[5] ),
    .GATE(net3212),
    .Q(\core.work.registers.genblk1[1].latch[5] ));
 sg13g2_dlhq_1 _11909_ (.D(net3425),
    .GATE(net3214),
    .Q(\core.work.registers.genblk1[1].latch[6] ));
 sg13g2_dlhq_1 _11910_ (.D(net3423),
    .GATE(net3213),
    .Q(\core.work.registers.genblk1[1].latch[7] ));
 sg13g2_dlhq_1 _11911_ (.D(net3422),
    .GATE(net3212),
    .Q(\core.work.registers.genblk1[1].latch[8] ));
 sg13g2_dlhq_1 _11912_ (.D(net3420),
    .GATE(net3214),
    .Q(\core.work.registers.genblk1[1].latch[9] ));
 sg13g2_dlhq_1 _11913_ (.D(net3418),
    .GATE(net3215),
    .Q(\core.work.registers.genblk1[1].latch[10] ));
 sg13g2_dlhq_1 _11914_ (.D(net3416),
    .GATE(net3211),
    .Q(\core.work.registers.genblk1[1].latch[11] ));
 sg13g2_dlhq_1 _11915_ (.D(\core.work.registers.tmp[12] ),
    .GATE(net3212),
    .Q(\core.work.registers.genblk1[1].latch[12] ));
 sg13g2_dlhq_1 _11916_ (.D(\core.work.registers.tmp[13] ),
    .GATE(net3215),
    .Q(\core.work.registers.genblk1[1].latch[13] ));
 sg13g2_dlhq_1 _11917_ (.D(net3409),
    .GATE(net3215),
    .Q(\core.work.registers.genblk1[1].latch[14] ));
 sg13g2_dlhq_1 _11918_ (.D(net3407),
    .GATE(net3212),
    .Q(\core.work.registers.genblk1[1].latch[15] ));
 sg13g2_dlhq_1 _11919_ (.D(net3404),
    .GATE(net3214),
    .Q(\core.work.registers.genblk1[1].latch[16] ));
 sg13g2_dlhq_1 _11920_ (.D(\core.work.registers.tmp[17] ),
    .GATE(net3213),
    .Q(\core.work.registers.genblk1[1].latch[17] ));
 sg13g2_dlhq_1 _11921_ (.D(\core.work.registers.tmp[18] ),
    .GATE(net3214),
    .Q(\core.work.registers.genblk1[1].latch[18] ));
 sg13g2_dlhq_1 _11922_ (.D(net3395),
    .GATE(net3213),
    .Q(\core.work.registers.genblk1[1].latch[19] ));
 sg13g2_dlhq_1 _11923_ (.D(net3393),
    .GATE(net3214),
    .Q(\core.work.registers.genblk1[1].latch[20] ));
 sg13g2_dlhq_1 _11924_ (.D(net3392),
    .GATE(net3212),
    .Q(\core.work.registers.genblk1[1].latch[21] ));
 sg13g2_dlhq_1 _11925_ (.D(\core.work.registers.tmp[22] ),
    .GATE(net3212),
    .Q(\core.work.registers.genblk1[1].latch[22] ));
 sg13g2_dlhq_1 _11926_ (.D(net3387),
    .GATE(net3211),
    .Q(\core.work.registers.genblk1[1].latch[23] ));
 sg13g2_dlhq_1 _11927_ (.D(net3384),
    .GATE(net3214),
    .Q(\core.work.registers.genblk1[1].latch[24] ));
 sg13g2_dlhq_1 _11928_ (.D(net3380),
    .GATE(net3212),
    .Q(\core.work.registers.genblk1[1].latch[25] ));
 sg13g2_dlhq_1 _11929_ (.D(\core.work.registers.tmp[26] ),
    .GATE(net3211),
    .Q(\core.work.registers.genblk1[1].latch[26] ));
 sg13g2_dlhq_1 _11930_ (.D(\core.work.registers.tmp[27] ),
    .GATE(net3211),
    .Q(\core.work.registers.genblk1[1].latch[27] ));
 sg13g2_dlhq_1 _11931_ (.D(\core.work.registers.tmp[28] ),
    .GATE(net3211),
    .Q(\core.work.registers.genblk1[1].latch[28] ));
 sg13g2_dlhq_1 _11932_ (.D(\core.work.registers.tmp[29] ),
    .GATE(net3211),
    .Q(\core.work.registers.genblk1[1].latch[29] ));
 sg13g2_dlhq_1 _11933_ (.D(net3368),
    .GATE(net3211),
    .Q(\core.work.registers.genblk1[1].latch[30] ));
 sg13g2_dlhq_1 _11934_ (.D(net3365),
    .GATE(net3211),
    .Q(\core.work.registers.genblk1[1].latch[31] ));
 sg13g2_dfrbp_1 _11935_ (.CLK(net348),
    .RESET_B(net3579),
    .D(_00015_),
    .Q_N(_05493_),
    .Q(\core.work.registers.genblk1[7].we ));
 sg13g2_dlhq_1 _11936_ (.D(net3439),
    .GATE(net3279),
    .Q(\core.work.registers.genblk1[13].latch[0] ));
 sg13g2_dlhq_1 _11937_ (.D(\core.work.registers.tmp[1] ),
    .GATE(net3279),
    .Q(\core.work.registers.genblk1[13].latch[1] ));
 sg13g2_dlhq_1 _11938_ (.D(net3435),
    .GATE(net3279),
    .Q(\core.work.registers.genblk1[13].latch[2] ));
 sg13g2_dlhq_1 _11939_ (.D(net3432),
    .GATE(net3279),
    .Q(\core.work.registers.genblk1[13].latch[3] ));
 sg13g2_dlhq_1 _11940_ (.D(net3430),
    .GATE(net3278),
    .Q(\core.work.registers.genblk1[13].latch[4] ));
 sg13g2_dlhq_1 _11941_ (.D(net3427),
    .GATE(net3277),
    .Q(\core.work.registers.genblk1[13].latch[5] ));
 sg13g2_dlhq_1 _11942_ (.D(net3426),
    .GATE(net3279),
    .Q(\core.work.registers.genblk1[13].latch[6] ));
 sg13g2_dlhq_1 _11943_ (.D(net3423),
    .GATE(net3278),
    .Q(\core.work.registers.genblk1[13].latch[7] ));
 sg13g2_dlhq_1 _11944_ (.D(net3421),
    .GATE(net3277),
    .Q(\core.work.registers.genblk1[13].latch[8] ));
 sg13g2_dlhq_1 _11945_ (.D(net3419),
    .GATE(net3278),
    .Q(\core.work.registers.genblk1[13].latch[9] ));
 sg13g2_dlhq_1 _11946_ (.D(net3418),
    .GATE(net3280),
    .Q(\core.work.registers.genblk1[13].latch[10] ));
 sg13g2_dlhq_1 _11947_ (.D(net3414),
    .GATE(net3277),
    .Q(\core.work.registers.genblk1[13].latch[11] ));
 sg13g2_dlhq_1 _11948_ (.D(net3413),
    .GATE(net3277),
    .Q(\core.work.registers.genblk1[13].latch[12] ));
 sg13g2_dlhq_1 _11949_ (.D(net3410),
    .GATE(net3277),
    .Q(\core.work.registers.genblk1[13].latch[13] ));
 sg13g2_dlhq_1 _11950_ (.D(net3409),
    .GATE(net3280),
    .Q(\core.work.registers.genblk1[13].latch[14] ));
 sg13g2_dlhq_1 _11951_ (.D(net3406),
    .GATE(net3276),
    .Q(\core.work.registers.genblk1[13].latch[15] ));
 sg13g2_dlhq_1 _11952_ (.D(net3402),
    .GATE(net3278),
    .Q(\core.work.registers.genblk1[13].latch[16] ));
 sg13g2_dlhq_1 _11953_ (.D(net3400),
    .GATE(net3278),
    .Q(\core.work.registers.genblk1[13].latch[17] ));
 sg13g2_dlhq_1 _11954_ (.D(net3399),
    .GATE(net3278),
    .Q(\core.work.registers.genblk1[13].latch[18] ));
 sg13g2_dlhq_1 _11955_ (.D(net3397),
    .GATE(net3279),
    .Q(\core.work.registers.genblk1[13].latch[19] ));
 sg13g2_dlhq_1 _11956_ (.D(net3394),
    .GATE(net3278),
    .Q(\core.work.registers.genblk1[13].latch[20] ));
 sg13g2_dlhq_1 _11957_ (.D(net3390),
    .GATE(net3277),
    .Q(\core.work.registers.genblk1[13].latch[21] ));
 sg13g2_dlhq_1 _11958_ (.D(net3389),
    .GATE(net3277),
    .Q(\core.work.registers.genblk1[13].latch[22] ));
 sg13g2_dlhq_1 _11959_ (.D(net3385),
    .GATE(net3276),
    .Q(\core.work.registers.genblk1[13].latch[23] ));
 sg13g2_dlhq_1 _11960_ (.D(net3382),
    .GATE(net3278),
    .Q(\core.work.registers.genblk1[13].latch[24] ));
 sg13g2_dlhq_1 _11961_ (.D(net3379),
    .GATE(net3280),
    .Q(\core.work.registers.genblk1[13].latch[25] ));
 sg13g2_dlhq_1 _11962_ (.D(net3377),
    .GATE(net3276),
    .Q(\core.work.registers.genblk1[13].latch[26] ));
 sg13g2_dlhq_1 _11963_ (.D(net3375),
    .GATE(net3276),
    .Q(\core.work.registers.genblk1[13].latch[27] ));
 sg13g2_dlhq_1 _11964_ (.D(net3372),
    .GATE(net3276),
    .Q(\core.work.registers.genblk1[13].latch[28] ));
 sg13g2_dlhq_1 _11965_ (.D(net3369),
    .GATE(net3276),
    .Q(\core.work.registers.genblk1[13].latch[29] ));
 sg13g2_dlhq_1 _11966_ (.D(net3366),
    .GATE(net3276),
    .Q(\core.work.registers.genblk1[13].latch[30] ));
 sg13g2_dlhq_1 _11967_ (.D(net3363),
    .GATE(net3276),
    .Q(\core.work.registers.genblk1[13].latch[31] ));
 sg13g2_dfrbp_1 _11968_ (.CLK(net349),
    .RESET_B(net3580),
    .D(_00014_),
    .Q_N(_05492_),
    .Q(\core.work.registers.genblk1[6].we ));
 sg13g2_dfrbp_1 _11969_ (.CLK(net350),
    .RESET_B(net3580),
    .D(_00013_),
    .Q_N(_05491_),
    .Q(\core.work.registers.genblk1[5].we ));
 sg13g2_dlhq_1 _11970_ (.D(net3438),
    .GATE(net3284),
    .Q(\core.work.registers.genblk1[14].latch[0] ));
 sg13g2_dlhq_1 _11971_ (.D(net3436),
    .GATE(net3284),
    .Q(\core.work.registers.genblk1[14].latch[1] ));
 sg13g2_dlhq_1 _11972_ (.D(net3434),
    .GATE(net3283),
    .Q(\core.work.registers.genblk1[14].latch[2] ));
 sg13g2_dlhq_1 _11973_ (.D(net3433),
    .GATE(net3284),
    .Q(\core.work.registers.genblk1[14].latch[3] ));
 sg13g2_dlhq_1 _11974_ (.D(net3430),
    .GATE(net3284),
    .Q(\core.work.registers.genblk1[14].latch[4] ));
 sg13g2_dlhq_1 _11975_ (.D(net3428),
    .GATE(net3282),
    .Q(\core.work.registers.genblk1[14].latch[5] ));
 sg13g2_dlhq_1 _11976_ (.D(net3425),
    .GATE(net3284),
    .Q(\core.work.registers.genblk1[14].latch[6] ));
 sg13g2_dlhq_1 _11977_ (.D(net3424),
    .GATE(net3283),
    .Q(\core.work.registers.genblk1[14].latch[7] ));
 sg13g2_dlhq_1 _11978_ (.D(net3422),
    .GATE(net3283),
    .Q(\core.work.registers.genblk1[14].latch[8] ));
 sg13g2_dlhq_1 _11979_ (.D(net3419),
    .GATE(net3283),
    .Q(\core.work.registers.genblk1[14].latch[9] ));
 sg13g2_dlhq_1 _11980_ (.D(net3417),
    .GATE(net3285),
    .Q(\core.work.registers.genblk1[14].latch[10] ));
 sg13g2_dlhq_1 _11981_ (.D(net3415),
    .GATE(net3282),
    .Q(\core.work.registers.genblk1[14].latch[11] ));
 sg13g2_dlhq_1 _11982_ (.D(net3412),
    .GATE(net3282),
    .Q(\core.work.registers.genblk1[14].latch[12] ));
 sg13g2_dlhq_1 _11983_ (.D(net3410),
    .GATE(net3282),
    .Q(\core.work.registers.genblk1[14].latch[13] ));
 sg13g2_dlhq_1 _11984_ (.D(net3408),
    .GATE(net3285),
    .Q(\core.work.registers.genblk1[14].latch[14] ));
 sg13g2_dlhq_1 _11985_ (.D(net3406),
    .GATE(net3281),
    .Q(\core.work.registers.genblk1[14].latch[15] ));
 sg13g2_dlhq_1 _11986_ (.D(net3402),
    .GATE(net3283),
    .Q(\core.work.registers.genblk1[14].latch[16] ));
 sg13g2_dlhq_1 _11987_ (.D(net3400),
    .GATE(net3284),
    .Q(\core.work.registers.genblk1[14].latch[17] ));
 sg13g2_dlhq_1 _11988_ (.D(net3398),
    .GATE(net3283),
    .Q(\core.work.registers.genblk1[14].latch[18] ));
 sg13g2_dlhq_1 _11989_ (.D(net3395),
    .GATE(net3284),
    .Q(\core.work.registers.genblk1[14].latch[19] ));
 sg13g2_dlhq_1 _11990_ (.D(net3394),
    .GATE(net3283),
    .Q(\core.work.registers.genblk1[14].latch[20] ));
 sg13g2_dlhq_1 _11991_ (.D(net3390),
    .GATE(net3282),
    .Q(\core.work.registers.genblk1[14].latch[21] ));
 sg13g2_dlhq_1 _11992_ (.D(net3389),
    .GATE(net3282),
    .Q(\core.work.registers.genblk1[14].latch[22] ));
 sg13g2_dlhq_1 _11993_ (.D(net3386),
    .GATE(net3281),
    .Q(\core.work.registers.genblk1[14].latch[23] ));
 sg13g2_dlhq_1 _11994_ (.D(net3382),
    .GATE(net3283),
    .Q(\core.work.registers.genblk1[14].latch[24] ));
 sg13g2_dlhq_1 _11995_ (.D(net3380),
    .GATE(net3282),
    .Q(\core.work.registers.genblk1[14].latch[25] ));
 sg13g2_dlhq_1 _11996_ (.D(net3378),
    .GATE(net3281),
    .Q(\core.work.registers.genblk1[14].latch[26] ));
 sg13g2_dlhq_1 _11997_ (.D(net3375),
    .GATE(net3281),
    .Q(\core.work.registers.genblk1[14].latch[27] ));
 sg13g2_dlhq_1 _11998_ (.D(net3373),
    .GATE(net3281),
    .Q(\core.work.registers.genblk1[14].latch[28] ));
 sg13g2_dlhq_1 _11999_ (.D(net3369),
    .GATE(net3281),
    .Q(\core.work.registers.genblk1[14].latch[29] ));
 sg13g2_dlhq_1 _12000_ (.D(net3367),
    .GATE(net3281),
    .Q(\core.work.registers.genblk1[14].latch[30] ));
 sg13g2_dlhq_1 _12001_ (.D(net3364),
    .GATE(net3281),
    .Q(\core.work.registers.genblk1[14].latch[31] ));
 sg13g2_dlhq_1 _12002_ (.D(net3439),
    .GATE(net3244),
    .Q(\core.work.registers.genblk1[6].latch[0] ));
 sg13g2_dlhq_1 _12003_ (.D(net3437),
    .GATE(net3244),
    .Q(\core.work.registers.genblk1[6].latch[1] ));
 sg13g2_dlhq_1 _12004_ (.D(net3435),
    .GATE(net3243),
    .Q(\core.work.registers.genblk1[6].latch[2] ));
 sg13g2_dlhq_1 _12005_ (.D(net3432),
    .GATE(net3244),
    .Q(\core.work.registers.genblk1[6].latch[3] ));
 sg13g2_dlhq_1 _12006_ (.D(net3430),
    .GATE(net3244),
    .Q(\core.work.registers.genblk1[6].latch[4] ));
 sg13g2_dlhq_1 _12007_ (.D(net3428),
    .GATE(net3242),
    .Q(\core.work.registers.genblk1[6].latch[5] ));
 sg13g2_dlhq_1 _12008_ (.D(net3425),
    .GATE(net3244),
    .Q(\core.work.registers.genblk1[6].latch[6] ));
 sg13g2_dlhq_1 _12009_ (.D(net3424),
    .GATE(net3243),
    .Q(\core.work.registers.genblk1[6].latch[7] ));
 sg13g2_dlhq_1 _12010_ (.D(net3421),
    .GATE(net3242),
    .Q(\core.work.registers.genblk1[6].latch[8] ));
 sg13g2_dlhq_1 _12011_ (.D(net3420),
    .GATE(net3243),
    .Q(\core.work.registers.genblk1[6].latch[9] ));
 sg13g2_dlhq_1 _12012_ (.D(net3417),
    .GATE(net3245),
    .Q(\core.work.registers.genblk1[6].latch[10] ));
 sg13g2_dlhq_1 _12013_ (.D(net3415),
    .GATE(net3242),
    .Q(\core.work.registers.genblk1[6].latch[11] ));
 sg13g2_dlhq_1 _12014_ (.D(net3412),
    .GATE(net3242),
    .Q(\core.work.registers.genblk1[6].latch[12] ));
 sg13g2_dlhq_1 _12015_ (.D(net3411),
    .GATE(net3242),
    .Q(\core.work.registers.genblk1[6].latch[13] ));
 sg13g2_dlhq_1 _12016_ (.D(net3408),
    .GATE(net3245),
    .Q(\core.work.registers.genblk1[6].latch[14] ));
 sg13g2_dlhq_1 _12017_ (.D(net3405),
    .GATE(net3241),
    .Q(\core.work.registers.genblk1[6].latch[15] ));
 sg13g2_dlhq_1 _12018_ (.D(net3403),
    .GATE(net3243),
    .Q(\core.work.registers.genblk1[6].latch[16] ));
 sg13g2_dlhq_1 _12019_ (.D(net3400),
    .GATE(net3243),
    .Q(\core.work.registers.genblk1[6].latch[17] ));
 sg13g2_dlhq_1 _12020_ (.D(net3398),
    .GATE(net3243),
    .Q(\core.work.registers.genblk1[6].latch[18] ));
 sg13g2_dlhq_1 _12021_ (.D(net3395),
    .GATE(net3244),
    .Q(\core.work.registers.genblk1[6].latch[19] ));
 sg13g2_dlhq_1 _12022_ (.D(net3393),
    .GATE(net3243),
    .Q(\core.work.registers.genblk1[6].latch[20] ));
 sg13g2_dlhq_1 _12023_ (.D(net3390),
    .GATE(net3242),
    .Q(\core.work.registers.genblk1[6].latch[21] ));
 sg13g2_dlhq_1 _12024_ (.D(net3388),
    .GATE(net3242),
    .Q(\core.work.registers.genblk1[6].latch[22] ));
 sg13g2_dlhq_1 _12025_ (.D(net3386),
    .GATE(net3241),
    .Q(\core.work.registers.genblk1[6].latch[23] ));
 sg13g2_dlhq_1 _12026_ (.D(net3383),
    .GATE(net3243),
    .Q(\core.work.registers.genblk1[6].latch[24] ));
 sg13g2_dlhq_1 _12027_ (.D(net3379),
    .GATE(net3245),
    .Q(\core.work.registers.genblk1[6].latch[25] ));
 sg13g2_dlhq_1 _12028_ (.D(net3377),
    .GATE(net3241),
    .Q(\core.work.registers.genblk1[6].latch[26] ));
 sg13g2_dlhq_1 _12029_ (.D(net3375),
    .GATE(net3241),
    .Q(\core.work.registers.genblk1[6].latch[27] ));
 sg13g2_dlhq_1 _12030_ (.D(net3374),
    .GATE(net3241),
    .Q(\core.work.registers.genblk1[6].latch[28] ));
 sg13g2_dlhq_1 _12031_ (.D(net3371),
    .GATE(net3241),
    .Q(\core.work.registers.genblk1[6].latch[29] ));
 sg13g2_dlhq_1 _12032_ (.D(net3368),
    .GATE(net3241),
    .Q(\core.work.registers.genblk1[6].latch[30] ));
 sg13g2_dlhq_1 _12033_ (.D(net3364),
    .GATE(net3241),
    .Q(\core.work.registers.genblk1[6].latch[31] ));
 sg13g2_dfrbp_1 _12034_ (.CLK(net351),
    .RESET_B(net3580),
    .D(_00012_),
    .Q_N(_05490_),
    .Q(\core.work.registers.genblk1[4].we ));
 sg13g2_dlhq_1 _12035_ (.D(net3438),
    .GATE(net3224),
    .Q(\core.work.registers.genblk1[15].latch[0] ));
 sg13g2_dlhq_1 _12036_ (.D(net3436),
    .GATE(net3224),
    .Q(\core.work.registers.genblk1[15].latch[1] ));
 sg13g2_dlhq_1 _12037_ (.D(net3434),
    .GATE(net3224),
    .Q(\core.work.registers.genblk1[15].latch[2] ));
 sg13g2_dlhq_1 _12038_ (.D(net3433),
    .GATE(net3223),
    .Q(\core.work.registers.genblk1[15].latch[3] ));
 sg13g2_dlhq_1 _12039_ (.D(net3429),
    .GATE(net3223),
    .Q(\core.work.registers.genblk1[15].latch[4] ));
 sg13g2_dlhq_1 _12040_ (.D(net3427),
    .GATE(net3222),
    .Q(\core.work.registers.genblk1[15].latch[5] ));
 sg13g2_dlhq_1 _12041_ (.D(net3426),
    .GATE(net3224),
    .Q(\core.work.registers.genblk1[15].latch[6] ));
 sg13g2_dlhq_1 _12042_ (.D(net3423),
    .GATE(net3224),
    .Q(\core.work.registers.genblk1[15].latch[7] ));
 sg13g2_dlhq_1 _12043_ (.D(net3421),
    .GATE(net3225),
    .Q(\core.work.registers.genblk1[15].latch[8] ));
 sg13g2_dlhq_1 _12044_ (.D(net3419),
    .GATE(net3223),
    .Q(\core.work.registers.genblk1[15].latch[9] ));
 sg13g2_dlhq_1 _12045_ (.D(net3417),
    .GATE(net3225),
    .Q(\core.work.registers.genblk1[15].latch[10] ));
 sg13g2_dlhq_1 _12046_ (.D(net3414),
    .GATE(net3222),
    .Q(\core.work.registers.genblk1[15].latch[11] ));
 sg13g2_dlhq_1 _12047_ (.D(net3413),
    .GATE(net3222),
    .Q(\core.work.registers.genblk1[15].latch[12] ));
 sg13g2_dlhq_1 _12048_ (.D(net3411),
    .GATE(net3222),
    .Q(\core.work.registers.genblk1[15].latch[13] ));
 sg13g2_dlhq_1 _12049_ (.D(net3408),
    .GATE(net3225),
    .Q(\core.work.registers.genblk1[15].latch[14] ));
 sg13g2_dlhq_1 _12050_ (.D(net3405),
    .GATE(net3221),
    .Q(\core.work.registers.genblk1[15].latch[15] ));
 sg13g2_dlhq_1 _12051_ (.D(net3403),
    .GATE(net3223),
    .Q(\core.work.registers.genblk1[15].latch[16] ));
 sg13g2_dlhq_1 _12052_ (.D(net3401),
    .GATE(net3223),
    .Q(\core.work.registers.genblk1[15].latch[17] ));
 sg13g2_dlhq_1 _12053_ (.D(net3398),
    .GATE(net3223),
    .Q(\core.work.registers.genblk1[15].latch[18] ));
 sg13g2_dlhq_1 _12054_ (.D(net3395),
    .GATE(net3224),
    .Q(\core.work.registers.genblk1[15].latch[19] ));
 sg13g2_dlhq_1 _12055_ (.D(net3394),
    .GATE(net3223),
    .Q(\core.work.registers.genblk1[15].latch[20] ));
 sg13g2_dlhq_1 _12056_ (.D(net3391),
    .GATE(net3222),
    .Q(\core.work.registers.genblk1[15].latch[21] ));
 sg13g2_dlhq_1 _12057_ (.D(net3388),
    .GATE(net3222),
    .Q(\core.work.registers.genblk1[15].latch[22] ));
 sg13g2_dlhq_1 _12058_ (.D(net3385),
    .GATE(net3221),
    .Q(\core.work.registers.genblk1[15].latch[23] ));
 sg13g2_dlhq_1 _12059_ (.D(net3383),
    .GATE(net3223),
    .Q(\core.work.registers.genblk1[15].latch[24] ));
 sg13g2_dlhq_1 _12060_ (.D(net3380),
    .GATE(net3222),
    .Q(\core.work.registers.genblk1[15].latch[25] ));
 sg13g2_dlhq_1 _12061_ (.D(net3377),
    .GATE(net3221),
    .Q(\core.work.registers.genblk1[15].latch[26] ));
 sg13g2_dlhq_1 _12062_ (.D(net3376),
    .GATE(net3221),
    .Q(\core.work.registers.genblk1[15].latch[27] ));
 sg13g2_dlhq_1 _12063_ (.D(net3372),
    .GATE(net3221),
    .Q(\core.work.registers.genblk1[15].latch[28] ));
 sg13g2_dlhq_1 _12064_ (.D(net3369),
    .GATE(net3221),
    .Q(\core.work.registers.genblk1[15].latch[29] ));
 sg13g2_dlhq_1 _12065_ (.D(net3366),
    .GATE(net3221),
    .Q(\core.work.registers.genblk1[15].latch[30] ));
 sg13g2_dlhq_1 _12066_ (.D(net3363),
    .GATE(net3221),
    .Q(\core.work.registers.genblk1[15].latch[31] ));
 sg13g2_dlhq_1 _12067_ (.D(net3439),
    .GATE(net3219),
    .Q(\core.work.registers.genblk1[2].latch[0] ));
 sg13g2_dlhq_1 _12068_ (.D(net3437),
    .GATE(net3219),
    .Q(\core.work.registers.genblk1[2].latch[1] ));
 sg13g2_dlhq_1 _12069_ (.D(net3435),
    .GATE(net3219),
    .Q(\core.work.registers.genblk1[2].latch[2] ));
 sg13g2_dlhq_1 _12070_ (.D(net3432),
    .GATE(net3218),
    .Q(\core.work.registers.genblk1[2].latch[3] ));
 sg13g2_dlhq_1 _12071_ (.D(net3429),
    .GATE(net3219),
    .Q(\core.work.registers.genblk1[2].latch[4] ));
 sg13g2_dlhq_1 _12072_ (.D(net3427),
    .GATE(net3217),
    .Q(\core.work.registers.genblk1[2].latch[5] ));
 sg13g2_dlhq_1 _12073_ (.D(net3426),
    .GATE(net3219),
    .Q(\core.work.registers.genblk1[2].latch[6] ));
 sg13g2_dlhq_1 _12074_ (.D(net3423),
    .GATE(net3218),
    .Q(\core.work.registers.genblk1[2].latch[7] ));
 sg13g2_dlhq_1 _12075_ (.D(net3422),
    .GATE(net3220),
    .Q(\core.work.registers.genblk1[2].latch[8] ));
 sg13g2_dlhq_1 _12076_ (.D(net3419),
    .GATE(net3218),
    .Q(\core.work.registers.genblk1[2].latch[9] ));
 sg13g2_dlhq_1 _12077_ (.D(net3418),
    .GATE(net3220),
    .Q(\core.work.registers.genblk1[2].latch[10] ));
 sg13g2_dlhq_1 _12078_ (.D(net3415),
    .GATE(net3217),
    .Q(\core.work.registers.genblk1[2].latch[11] ));
 sg13g2_dlhq_1 _12079_ (.D(net3412),
    .GATE(net3217),
    .Q(\core.work.registers.genblk1[2].latch[12] ));
 sg13g2_dlhq_1 _12080_ (.D(net3410),
    .GATE(net3217),
    .Q(\core.work.registers.genblk1[2].latch[13] ));
 sg13g2_dlhq_1 _12081_ (.D(net3409),
    .GATE(net3220),
    .Q(\core.work.registers.genblk1[2].latch[14] ));
 sg13g2_dlhq_1 _12082_ (.D(net3406),
    .GATE(net3216),
    .Q(\core.work.registers.genblk1[2].latch[15] ));
 sg13g2_dlhq_1 _12083_ (.D(net3402),
    .GATE(net3218),
    .Q(\core.work.registers.genblk1[2].latch[16] ));
 sg13g2_dlhq_1 _12084_ (.D(net3400),
    .GATE(net3218),
    .Q(\core.work.registers.genblk1[2].latch[17] ));
 sg13g2_dlhq_1 _12085_ (.D(net3398),
    .GATE(net3218),
    .Q(\core.work.registers.genblk1[2].latch[18] ));
 sg13g2_dlhq_1 _12086_ (.D(net3397),
    .GATE(net3219),
    .Q(\core.work.registers.genblk1[2].latch[19] ));
 sg13g2_dlhq_1 _12087_ (.D(\core.work.registers.tmp[20] ),
    .GATE(net3218),
    .Q(\core.work.registers.genblk1[2].latch[20] ));
 sg13g2_dlhq_1 _12088_ (.D(net3390),
    .GATE(net3217),
    .Q(\core.work.registers.genblk1[2].latch[21] ));
 sg13g2_dlhq_1 _12089_ (.D(net3389),
    .GATE(net3217),
    .Q(\core.work.registers.genblk1[2].latch[22] ));
 sg13g2_dlhq_1 _12090_ (.D(net3387),
    .GATE(net3216),
    .Q(\core.work.registers.genblk1[2].latch[23] ));
 sg13g2_dlhq_1 _12091_ (.D(net3383),
    .GATE(net3218),
    .Q(\core.work.registers.genblk1[2].latch[24] ));
 sg13g2_dlhq_1 _12092_ (.D(net3379),
    .GATE(net3217),
    .Q(\core.work.registers.genblk1[2].latch[25] ));
 sg13g2_dlhq_1 _12093_ (.D(net3377),
    .GATE(net3216),
    .Q(\core.work.registers.genblk1[2].latch[26] ));
 sg13g2_dlhq_1 _12094_ (.D(net3375),
    .GATE(net3216),
    .Q(\core.work.registers.genblk1[2].latch[27] ));
 sg13g2_dlhq_1 _12095_ (.D(net3373),
    .GATE(net3216),
    .Q(\core.work.registers.genblk1[2].latch[28] ));
 sg13g2_dlhq_1 _12096_ (.D(net3370),
    .GATE(net3216),
    .Q(\core.work.registers.genblk1[2].latch[29] ));
 sg13g2_dlhq_1 _12097_ (.D(net3366),
    .GATE(net3216),
    .Q(\core.work.registers.genblk1[2].latch[30] ));
 sg13g2_dlhq_1 _12098_ (.D(net3363),
    .GATE(net3216),
    .Q(\core.work.registers.genblk1[2].latch[31] ));
 sg13g2_dfrbp_1 _12099_ (.CLK(net352),
    .RESET_B(net3580),
    .D(_00011_),
    .Q_N(_05489_),
    .Q(\core.work.registers.genblk1[3].we ));
 sg13g2_dfrbp_1 _12100_ (.CLK(net353),
    .RESET_B(net3579),
    .D(_00008_),
    .Q_N(_05488_),
    .Q(\core.work.registers.genblk1[15].we ));
 sg13g2_dfrbp_1 _12101_ (.CLK(net354),
    .RESET_B(net3580),
    .D(_00010_),
    .Q_N(_05487_),
    .Q(\core.work.registers.genblk1[2].we ));
 sg13g2_dfrbp_1 _12102_ (.CLK(net355),
    .RESET_B(net3580),
    .D(_00009_),
    .Q_N(_05486_),
    .Q(\core.work.registers.genblk1[1].we ));
 sg13g2_dfrbp_1 _12103_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3589),
    .D(_00524_),
    .Q_N(_05485_),
    .Q(\core.work.alu.ls_size_b ));
 sg13g2_dfrbp_1 _12104_ (.CLK(clknet_leaf_8_clk_regs),
    .RESET_B(net3589),
    .D(_00525_),
    .Q_N(_05484_),
    .Q(\core.work.alu.ls_size_h ));
 sg13g2_dfrbp_1 _12105_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3595),
    .D(_00526_),
    .Q_N(_05483_),
    .Q(\core.work.alu.is_sign ));
 sg13g2_dfrbp_1 _12106_ (.CLK(clknet_leaf_7_clk_regs),
    .RESET_B(net3588),
    .D(_00527_),
    .Q_N(_05482_),
    .Q(\core.work.alu.is_wr ));
 sg13g2_dfrbp_1 _12107_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net334),
    .D(_00528_),
    .Q_N(_05481_),
    .Q(\core.fetch.inst[32] ));
 sg13g2_dfrbp_1 _12108_ (.CLK(clknet_leaf_57_clk_regs),
    .RESET_B(net259),
    .D(_00529_),
    .Q_N(_05480_),
    .Q(\core.fetch.inst[33] ));
 sg13g2_dfrbp_1 _12109_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net255),
    .D(net586),
    .Q_N(_05479_),
    .Q(\core.fetch.inst[34] ));
 sg13g2_dfrbp_1 _12110_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net251),
    .D(_00531_),
    .Q_N(_05478_),
    .Q(\core.fetch.inst[35] ));
 sg13g2_dfrbp_1 _12111_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net247),
    .D(_00532_),
    .Q_N(_05477_),
    .Q(\core.fetch.inst[36] ));
 sg13g2_dfrbp_1 _12112_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net243),
    .D(_00533_),
    .Q_N(_05476_),
    .Q(\core.fetch.inst[37] ));
 sg13g2_dfrbp_1 _12113_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net239),
    .D(_00534_),
    .Q_N(_05475_),
    .Q(\core.fetch.inst[38] ));
 sg13g2_dfrbp_1 _12114_ (.CLK(clknet_leaf_13_clk_regs),
    .RESET_B(net235),
    .D(_00535_),
    .Q_N(_05474_),
    .Q(\core.fetch.inst[39] ));
 sg13g2_dfrbp_1 _12115_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net231),
    .D(_00536_),
    .Q_N(_05473_),
    .Q(\core.fetch.inst[40] ));
 sg13g2_dfrbp_1 _12116_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net227),
    .D(_00537_),
    .Q_N(_05472_),
    .Q(\core.fetch.inst[41] ));
 sg13g2_dfrbp_1 _12117_ (.CLK(clknet_leaf_12_clk_regs),
    .RESET_B(net106),
    .D(net554),
    .Q_N(_05471_),
    .Q(\core.fetch.inst[42] ));
 sg13g2_dfrbp_1 _12118_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net102),
    .D(_00539_),
    .Q_N(_05470_),
    .Q(\core.fetch.inst[43] ));
 sg13g2_dfrbp_1 _12119_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net98),
    .D(_00540_),
    .Q_N(_05469_),
    .Q(\core.fetch.inst[44] ));
 sg13g2_dfrbp_1 _12120_ (.CLK(clknet_leaf_2_clk_regs),
    .RESET_B(net94),
    .D(_00541_),
    .Q_N(_05468_),
    .Q(\core.fetch.inst[45] ));
 sg13g2_dfrbp_1 _12121_ (.CLK(clknet_leaf_4_clk_regs),
    .RESET_B(net90),
    .D(net575),
    .Q_N(_05467_),
    .Q(\core.fetch.inst[46] ));
 sg13g2_dfrbp_1 _12122_ (.CLK(clknet_leaf_3_clk_regs),
    .RESET_B(net86),
    .D(net535),
    .Q_N(_05466_),
    .Q(\core.fetch.inst[47] ));
 sg13g2_dfrbp_1 _12123_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net3581),
    .D(net763),
    .Q_N(_05465_),
    .Q(\core.work.registers.state[0] ));
 sg13g2_dfrbp_1 _12124_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net3581),
    .D(net743),
    .Q_N(_05464_),
    .Q(\core.work.registers.state[1] ));
 sg13g2_dfrbp_1 _12125_ (.CLK(clknet_leaf_0_clk_regs),
    .RESET_B(net3581),
    .D(_00546_),
    .Q_N(_00058_),
    .Q(\core.work.registers.state[2] ));
 sg13g2_dlhq_1 _12126_ (.D(net3439),
    .GATE(net3249),
    .Q(\core.work.registers.genblk1[7].latch[0] ));
 sg13g2_dlhq_1 _12127_ (.D(net3437),
    .GATE(net3249),
    .Q(\core.work.registers.genblk1[7].latch[1] ));
 sg13g2_dlhq_1 _12128_ (.D(net3435),
    .GATE(net3249),
    .Q(\core.work.registers.genblk1[7].latch[2] ));
 sg13g2_dlhq_1 _12129_ (.D(net3432),
    .GATE(net3248),
    .Q(\core.work.registers.genblk1[7].latch[3] ));
 sg13g2_dlhq_1 _12130_ (.D(net3429),
    .GATE(net3249),
    .Q(\core.work.registers.genblk1[7].latch[4] ));
 sg13g2_dlhq_1 _12131_ (.D(net3427),
    .GATE(net3247),
    .Q(\core.work.registers.genblk1[7].latch[5] ));
 sg13g2_dlhq_1 _12132_ (.D(net3425),
    .GATE(net3249),
    .Q(\core.work.registers.genblk1[7].latch[6] ));
 sg13g2_dlhq_1 _12133_ (.D(net3423),
    .GATE(net3248),
    .Q(\core.work.registers.genblk1[7].latch[7] ));
 sg13g2_dlhq_1 _12134_ (.D(net3421),
    .GATE(net3250),
    .Q(\core.work.registers.genblk1[7].latch[8] ));
 sg13g2_dlhq_1 _12135_ (.D(net3420),
    .GATE(net3248),
    .Q(\core.work.registers.genblk1[7].latch[9] ));
 sg13g2_dlhq_1 _12136_ (.D(net3417),
    .GATE(net3250),
    .Q(\core.work.registers.genblk1[7].latch[10] ));
 sg13g2_dlhq_1 _12137_ (.D(net3414),
    .GATE(net3247),
    .Q(\core.work.registers.genblk1[7].latch[11] ));
 sg13g2_dlhq_1 _12138_ (.D(net3412),
    .GATE(net3247),
    .Q(\core.work.registers.genblk1[7].latch[12] ));
 sg13g2_dlhq_1 _12139_ (.D(net3410),
    .GATE(net3247),
    .Q(\core.work.registers.genblk1[7].latch[13] ));
 sg13g2_dlhq_1 _12140_ (.D(net3408),
    .GATE(net3250),
    .Q(\core.work.registers.genblk1[7].latch[14] ));
 sg13g2_dlhq_1 _12141_ (.D(net3405),
    .GATE(net3246),
    .Q(\core.work.registers.genblk1[7].latch[15] ));
 sg13g2_dlhq_1 _12142_ (.D(net3402),
    .GATE(net3248),
    .Q(\core.work.registers.genblk1[7].latch[16] ));
 sg13g2_dlhq_1 _12143_ (.D(net3400),
    .GATE(net3248),
    .Q(\core.work.registers.genblk1[7].latch[17] ));
 sg13g2_dlhq_1 _12144_ (.D(net3398),
    .GATE(net3248),
    .Q(\core.work.registers.genblk1[7].latch[18] ));
 sg13g2_dlhq_1 _12145_ (.D(net3396),
    .GATE(net3249),
    .Q(\core.work.registers.genblk1[7].latch[19] ));
 sg13g2_dlhq_1 _12146_ (.D(net3393),
    .GATE(net3248),
    .Q(\core.work.registers.genblk1[7].latch[20] ));
 sg13g2_dlhq_1 _12147_ (.D(net3391),
    .GATE(net3247),
    .Q(\core.work.registers.genblk1[7].latch[21] ));
 sg13g2_dlhq_1 _12148_ (.D(net3388),
    .GATE(net3247),
    .Q(\core.work.registers.genblk1[7].latch[22] ));
 sg13g2_dlhq_1 _12149_ (.D(net3385),
    .GATE(net3246),
    .Q(\core.work.registers.genblk1[7].latch[23] ));
 sg13g2_dlhq_1 _12150_ (.D(net3382),
    .GATE(net3248),
    .Q(\core.work.registers.genblk1[7].latch[24] ));
 sg13g2_dlhq_1 _12151_ (.D(net3380),
    .GATE(net3247),
    .Q(\core.work.registers.genblk1[7].latch[25] ));
 sg13g2_dlhq_1 _12152_ (.D(net3378),
    .GATE(net3246),
    .Q(\core.work.registers.genblk1[7].latch[26] ));
 sg13g2_dlhq_1 _12153_ (.D(net3375),
    .GATE(net3246),
    .Q(\core.work.registers.genblk1[7].latch[27] ));
 sg13g2_dlhq_1 _12154_ (.D(net3372),
    .GATE(net3246),
    .Q(\core.work.registers.genblk1[7].latch[28] ));
 sg13g2_dlhq_1 _12155_ (.D(net3370),
    .GATE(net3246),
    .Q(\core.work.registers.genblk1[7].latch[29] ));
 sg13g2_dlhq_1 _12156_ (.D(net3366),
    .GATE(net3246),
    .Q(\core.work.registers.genblk1[7].latch[30] ));
 sg13g2_dlhq_1 _12157_ (.D(net3363),
    .GATE(net3246),
    .Q(\core.work.registers.genblk1[7].latch[31] ));
 sg13g2_dfrbp_1 _12158_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net79),
    .D(_00547_),
    .Q_N(_05463_),
    .Q(\core.work.registers.tmp[0] ));
 sg13g2_dfrbp_1 _12159_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net77),
    .D(net745),
    .Q_N(_05462_),
    .Q(\core.work.registers.tmp[1] ));
 sg13g2_dfrbp_1 _12160_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net75),
    .D(_00549_),
    .Q_N(_05461_),
    .Q(\core.work.registers.tmp[2] ));
 sg13g2_dfrbp_1 _12161_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net73),
    .D(_00550_),
    .Q_N(_05460_),
    .Q(\core.work.registers.tmp[3] ));
 sg13g2_dfrbp_1 _12162_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net71),
    .D(_00551_),
    .Q_N(_05459_),
    .Q(\core.work.registers.tmp[4] ));
 sg13g2_dfrbp_1 _12163_ (.CLK(clknet_leaf_53_clk_regs),
    .RESET_B(net69),
    .D(net577),
    .Q_N(_05458_),
    .Q(\core.work.registers.tmp[5] ));
 sg13g2_dfrbp_1 _12164_ (.CLK(clknet_leaf_48_clk_regs),
    .RESET_B(net67),
    .D(_00553_),
    .Q_N(_05457_),
    .Q(\core.work.registers.tmp[6] ));
 sg13g2_dfrbp_1 _12165_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net65),
    .D(_00554_),
    .Q_N(_05456_),
    .Q(\core.work.registers.tmp[7] ));
 sg13g2_dfrbp_1 _12166_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net63),
    .D(net852),
    .Q_N(_05455_),
    .Q(\core.work.registers.tmp[8] ));
 sg13g2_dfrbp_1 _12167_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net61),
    .D(_00556_),
    .Q_N(_05454_),
    .Q(\core.work.registers.tmp[9] ));
 sg13g2_dfrbp_1 _12168_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net59),
    .D(_00557_),
    .Q_N(_05453_),
    .Q(\core.work.registers.tmp[10] ));
 sg13g2_dfrbp_1 _12169_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net57),
    .D(_00558_),
    .Q_N(_05452_),
    .Q(\core.work.registers.tmp[11] ));
 sg13g2_dfrbp_1 _12170_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net55),
    .D(_00559_),
    .Q_N(_05451_),
    .Q(\core.work.registers.tmp[12] ));
 sg13g2_dfrbp_1 _12171_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net53),
    .D(_00560_),
    .Q_N(_05450_),
    .Q(\core.work.registers.tmp[13] ));
 sg13g2_dfrbp_1 _12172_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net51),
    .D(_00561_),
    .Q_N(_05449_),
    .Q(\core.work.registers.tmp[14] ));
 sg13g2_dfrbp_1 _12173_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net49),
    .D(_00562_),
    .Q_N(_05448_),
    .Q(\core.work.registers.tmp[15] ));
 sg13g2_dfrbp_1 _12174_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net47),
    .D(net752),
    .Q_N(_05447_),
    .Q(\core.work.registers.tmp[16] ));
 sg13g2_dfrbp_1 _12175_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net333),
    .D(net600),
    .Q_N(_05446_),
    .Q(\core.work.registers.tmp[17] ));
 sg13g2_dfrbp_1 _12176_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net257),
    .D(_00565_),
    .Q_N(_05445_),
    .Q(\core.work.registers.tmp[18] ));
 sg13g2_dfrbp_1 _12177_ (.CLK(clknet_leaf_47_clk_regs),
    .RESET_B(net253),
    .D(net410),
    .Q_N(_05444_),
    .Q(\core.work.registers.tmp[19] ));
 sg13g2_dfrbp_1 _12178_ (.CLK(clknet_leaf_49_clk_regs),
    .RESET_B(net249),
    .D(_00567_),
    .Q_N(_05443_),
    .Q(\core.work.registers.tmp[20] ));
 sg13g2_dfrbp_1 _12179_ (.CLK(clknet_leaf_55_clk_regs),
    .RESET_B(net245),
    .D(_00568_),
    .Q_N(_05442_),
    .Q(\core.work.registers.tmp[21] ));
 sg13g2_dfrbp_1 _12180_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net241),
    .D(net441),
    .Q_N(_05441_),
    .Q(\core.work.registers.tmp[22] ));
 sg13g2_dfrbp_1 _12181_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net237),
    .D(_00570_),
    .Q_N(_05440_),
    .Q(\core.work.registers.tmp[23] ));
 sg13g2_dfrbp_1 _12182_ (.CLK(clknet_leaf_50_clk_regs),
    .RESET_B(net233),
    .D(_00571_),
    .Q_N(_05439_),
    .Q(\core.work.registers.tmp[24] ));
 sg13g2_dfrbp_1 _12183_ (.CLK(clknet_leaf_54_clk_regs),
    .RESET_B(net229),
    .D(_00572_),
    .Q_N(_05438_),
    .Q(\core.work.registers.tmp[25] ));
 sg13g2_dfrbp_1 _12184_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net203),
    .D(_00573_),
    .Q_N(_05437_),
    .Q(\core.work.registers.tmp[26] ));
 sg13g2_dfrbp_1 _12185_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net104),
    .D(_00574_),
    .Q_N(_05436_),
    .Q(\core.work.registers.tmp[27] ));
 sg13g2_dfrbp_1 _12186_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net100),
    .D(_00575_),
    .Q_N(_05435_),
    .Q(\core.work.registers.tmp[28] ));
 sg13g2_dfrbp_1 _12187_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net96),
    .D(net627),
    .Q_N(_05434_),
    .Q(\core.work.registers.tmp[29] ));
 sg13g2_dfrbp_1 _12188_ (.CLK(clknet_leaf_1_clk_regs),
    .RESET_B(net92),
    .D(_00577_),
    .Q_N(_05433_),
    .Q(\core.work.registers.tmp[30] ));
 sg13g2_dfrbp_1 _12189_ (.CLK(clknet_leaf_56_clk_regs),
    .RESET_B(net88),
    .D(_00578_),
    .Q_N(_05432_),
    .Q(\core.work.registers.tmp[31] ));
 sg13g2_tiehi _11638__16 (.L_HI(net16));
 sg13g2_tiehi _11637__17 (.L_HI(net17));
 sg13g2_tiehi _11636__18 (.L_HI(net18));
 sg13g2_tiehi _11635__19 (.L_HI(net19));
 sg13g2_tiehi _11634__20 (.L_HI(net20));
 sg13g2_tiehi _11633__21 (.L_HI(net21));
 sg13g2_tiehi _11632__22 (.L_HI(net22));
 sg13g2_tiehi _11631__23 (.L_HI(net23));
 sg13g2_tiehi _11630__24 (.L_HI(net24));
 sg13g2_tiehi _11629__25 (.L_HI(net25));
 sg13g2_tiehi _11628__26 (.L_HI(net26));
 sg13g2_tiehi _11627__27 (.L_HI(net27));
 sg13g2_tiehi _11626__28 (.L_HI(net28));
 sg13g2_tiehi _11625__29 (.L_HI(net29));
 sg13g2_tiehi _11624__30 (.L_HI(net30));
 sg13g2_tiehi _11623__31 (.L_HI(net31));
 sg13g2_tiehi _11622__32 (.L_HI(net32));
 sg13g2_tiehi _11621__33 (.L_HI(net33));
 sg13g2_tiehi _11620__34 (.L_HI(net34));
 sg13g2_tiehi _11619__35 (.L_HI(net35));
 sg13g2_tiehi _11618__36 (.L_HI(net36));
 sg13g2_tiehi _11617__37 (.L_HI(net37));
 sg13g2_tiehi _11616__38 (.L_HI(net38));
 sg13g2_tiehi _11615__39 (.L_HI(net39));
 sg13g2_tiehi _11614__40 (.L_HI(net40));
 sg13g2_tiehi _11613__41 (.L_HI(net41));
 sg13g2_tiehi _11612__42 (.L_HI(net42));
 sg13g2_tiehi _11611__43 (.L_HI(net43));
 sg13g2_tiehi _11610__44 (.L_HI(net44));
 sg13g2_tiehi _11609__45 (.L_HI(net45));
 sg13g2_tiehi _11608__46 (.L_HI(net46));
 sg13g2_tiehi _12174__47 (.L_HI(net47));
 sg13g2_tiehi _11606__48 (.L_HI(net48));
 sg13g2_tiehi _12173__49 (.L_HI(net49));
 sg13g2_tiehi _11605__50 (.L_HI(net50));
 sg13g2_tiehi _12172__51 (.L_HI(net51));
 sg13g2_tiehi _11604__52 (.L_HI(net52));
 sg13g2_tiehi _12171__53 (.L_HI(net53));
 sg13g2_tiehi _11603__54 (.L_HI(net54));
 sg13g2_tiehi _12170__55 (.L_HI(net55));
 sg13g2_tiehi _11602__56 (.L_HI(net56));
 sg13g2_tiehi _12169__57 (.L_HI(net57));
 sg13g2_tiehi _11601__58 (.L_HI(net58));
 sg13g2_tiehi _12168__59 (.L_HI(net59));
 sg13g2_tiehi _11600__60 (.L_HI(net60));
 sg13g2_tiehi _12167__61 (.L_HI(net61));
 sg13g2_tiehi _11599__62 (.L_HI(net62));
 sg13g2_tiehi _12166__63 (.L_HI(net63));
 sg13g2_tiehi _11598__64 (.L_HI(net64));
 sg13g2_tiehi _12165__65 (.L_HI(net65));
 sg13g2_tiehi _11597__66 (.L_HI(net66));
 sg13g2_tiehi _12164__67 (.L_HI(net67));
 sg13g2_tiehi _11596__68 (.L_HI(net68));
 sg13g2_tiehi _12163__69 (.L_HI(net69));
 sg13g2_tiehi _11595__70 (.L_HI(net70));
 sg13g2_tiehi _12162__71 (.L_HI(net71));
 sg13g2_tiehi _11594__72 (.L_HI(net72));
 sg13g2_tiehi _12161__73 (.L_HI(net73));
 sg13g2_tiehi _11593__74 (.L_HI(net74));
 sg13g2_tiehi _12160__75 (.L_HI(net75));
 sg13g2_tiehi _11592__76 (.L_HI(net76));
 sg13g2_tiehi _12159__77 (.L_HI(net77));
 sg13g2_tiehi _11591__78 (.L_HI(net78));
 sg13g2_tiehi _12158__79 (.L_HI(net79));
 sg13g2_tiehi _11590__80 (.L_HI(net80));
 sg13g2_tiehi _11589__81 (.L_HI(net81));
 sg13g2_tiehi _11588__82 (.L_HI(net82));
 sg13g2_tiehi _11587__83 (.L_HI(net83));
 sg13g2_tiehi _11496__84 (.L_HI(net84));
 sg13g2_tiehi _11586__85 (.L_HI(net85));
 sg13g2_tiehi _12122__86 (.L_HI(net86));
 sg13g2_tiehi _11585__87 (.L_HI(net87));
 sg13g2_tiehi _12189__88 (.L_HI(net88));
 sg13g2_tiehi _11584__89 (.L_HI(net89));
 sg13g2_tiehi _12121__90 (.L_HI(net90));
 sg13g2_tiehi _11583__91 (.L_HI(net91));
 sg13g2_tiehi _12188__92 (.L_HI(net92));
 sg13g2_tiehi _11582__93 (.L_HI(net93));
 sg13g2_tiehi _12120__94 (.L_HI(net94));
 sg13g2_tiehi _11581__95 (.L_HI(net95));
 sg13g2_tiehi _12187__96 (.L_HI(net96));
 sg13g2_tiehi _11580__97 (.L_HI(net97));
 sg13g2_tiehi _12119__98 (.L_HI(net98));
 sg13g2_tiehi _11579__99 (.L_HI(net99));
 sg13g2_tiehi _12186__100 (.L_HI(net100));
 sg13g2_tiehi _11578__101 (.L_HI(net101));
 sg13g2_tiehi _12118__102 (.L_HI(net102));
 sg13g2_tiehi _11577__103 (.L_HI(net103));
 sg13g2_tiehi _12185__104 (.L_HI(net104));
 sg13g2_tiehi _11576__105 (.L_HI(net105));
 sg13g2_tiehi _12117__106 (.L_HI(net106));
 sg13g2_tiehi _11575__107 (.L_HI(net107));
 sg13g2_tiehi _11568__108 (.L_HI(net108));
 sg13g2_tiehi _11566__109 (.L_HI(net109));
 sg13g2_tiehi _11565__110 (.L_HI(net110));
 sg13g2_tiehi _11564__111 (.L_HI(net111));
 sg13g2_tiehi _11563__112 (.L_HI(net112));
 sg13g2_tiehi _11562__113 (.L_HI(net113));
 sg13g2_tiehi _11561__114 (.L_HI(net114));
 sg13g2_tiehi _11560__115 (.L_HI(net115));
 sg13g2_tiehi _11559__116 (.L_HI(net116));
 sg13g2_tiehi _11558__117 (.L_HI(net117));
 sg13g2_tiehi _11557__118 (.L_HI(net118));
 sg13g2_tiehi _11556__119 (.L_HI(net119));
 sg13g2_tiehi _11555__120 (.L_HI(net120));
 sg13g2_tiehi _11554__121 (.L_HI(net121));
 sg13g2_tiehi _11553__122 (.L_HI(net122));
 sg13g2_tiehi _11552__123 (.L_HI(net123));
 sg13g2_tiehi _11551__124 (.L_HI(net124));
 sg13g2_tiehi _11550__125 (.L_HI(net125));
 sg13g2_tiehi _11549__126 (.L_HI(net126));
 sg13g2_tiehi _11548__127 (.L_HI(net127));
 sg13g2_tiehi _11547__128 (.L_HI(net128));
 sg13g2_tiehi _11546__129 (.L_HI(net129));
 sg13g2_tiehi _11545__130 (.L_HI(net130));
 sg13g2_tiehi _11544__131 (.L_HI(net131));
 sg13g2_tiehi _11543__132 (.L_HI(net132));
 sg13g2_tiehi _11542__133 (.L_HI(net133));
 sg13g2_tiehi _11541__134 (.L_HI(net134));
 sg13g2_tiehi _11540__135 (.L_HI(net135));
 sg13g2_tiehi _11539__136 (.L_HI(net136));
 sg13g2_tiehi _11538__137 (.L_HI(net137));
 sg13g2_tiehi _11537__138 (.L_HI(net138));
 sg13g2_tiehi _11536__139 (.L_HI(net139));
 sg13g2_tiehi _11535__140 (.L_HI(net140));
 sg13g2_tiehi _11522__141 (.L_HI(net141));
 sg13g2_tiehi _11521__142 (.L_HI(net142));
 sg13g2_tiehi _11520__143 (.L_HI(net143));
 sg13g2_tiehi _11519__144 (.L_HI(net144));
 sg13g2_tiehi _11518__145 (.L_HI(net145));
 sg13g2_tiehi _11517__146 (.L_HI(net146));
 sg13g2_tiehi _11516__147 (.L_HI(net147));
 sg13g2_tiehi _11515__148 (.L_HI(net148));
 sg13g2_tiehi _11514__149 (.L_HI(net149));
 sg13g2_tiehi _11513__150 (.L_HI(net150));
 sg13g2_tiehi _11512__151 (.L_HI(net151));
 sg13g2_tiehi _11511__152 (.L_HI(net152));
 sg13g2_tiehi _11510__153 (.L_HI(net153));
 sg13g2_tiehi _11509__154 (.L_HI(net154));
 sg13g2_tiehi _11508__155 (.L_HI(net155));
 sg13g2_tiehi _11507__156 (.L_HI(net156));
 sg13g2_tiehi _11506__157 (.L_HI(net157));
 sg13g2_tiehi _11505__158 (.L_HI(net158));
 sg13g2_tiehi _11504__159 (.L_HI(net159));
 sg13g2_tiehi _11503__160 (.L_HI(net160));
 sg13g2_tiehi _11502__161 (.L_HI(net161));
 sg13g2_tiehi _11501__162 (.L_HI(net162));
 sg13g2_tiehi _11500__163 (.L_HI(net163));
 sg13g2_tiehi _11499__164 (.L_HI(net164));
 sg13g2_tiehi _11494__165 (.L_HI(net165));
 sg13g2_tiehi _11493__166 (.L_HI(net166));
 sg13g2_tiehi _11492__167 (.L_HI(net167));
 sg13g2_tiehi _11491__168 (.L_HI(net168));
 sg13g2_tiehi _11490__169 (.L_HI(net169));
 sg13g2_tiehi _11489__170 (.L_HI(net170));
 sg13g2_tiehi _11488__171 (.L_HI(net171));
 sg13g2_tiehi _11487__172 (.L_HI(net172));
 sg13g2_tiehi _11486__173 (.L_HI(net173));
 sg13g2_tiehi _11485__174 (.L_HI(net174));
 sg13g2_tiehi _11484__175 (.L_HI(net175));
 sg13g2_tiehi _11483__176 (.L_HI(net176));
 sg13g2_tiehi _11441__177 (.L_HI(net177));
 sg13g2_tiehi _11482__178 (.L_HI(net178));
 sg13g2_tiehi _11481__179 (.L_HI(net179));
 sg13g2_tiehi _11480__180 (.L_HI(net180));
 sg13g2_tiehi _11479__181 (.L_HI(net181));
 sg13g2_tiehi _11478__182 (.L_HI(net182));
 sg13g2_tiehi _11477__183 (.L_HI(net183));
 sg13g2_tiehi _11476__184 (.L_HI(net184));
 sg13g2_tiehi _11475__185 (.L_HI(net185));
 sg13g2_tiehi _11474__186 (.L_HI(net186));
 sg13g2_tiehi _11473__187 (.L_HI(net187));
 sg13g2_tiehi _11472__188 (.L_HI(net188));
 sg13g2_tiehi _11471__189 (.L_HI(net189));
 sg13g2_tiehi _11470__190 (.L_HI(net190));
 sg13g2_tiehi _11469__191 (.L_HI(net191));
 sg13g2_tiehi _11468__192 (.L_HI(net192));
 sg13g2_tiehi _11467__193 (.L_HI(net193));
 sg13g2_tiehi _11466__194 (.L_HI(net194));
 sg13g2_tiehi _11465__195 (.L_HI(net195));
 sg13g2_tiehi _11464__196 (.L_HI(net196));
 sg13g2_tiehi _11463__197 (.L_HI(net197));
 sg13g2_tiehi _11462__198 (.L_HI(net198));
 sg13g2_tiehi _11461__199 (.L_HI(net199));
 sg13g2_tiehi _11460__200 (.L_HI(net200));
 sg13g2_tiehi _11459__201 (.L_HI(net201));
 sg13g2_tiehi _11458__202 (.L_HI(net202));
 sg13g2_tiehi _12184__203 (.L_HI(net203));
 sg13g2_tiehi _11457__204 (.L_HI(net204));
 sg13g2_tiehi _11456__205 (.L_HI(net205));
 sg13g2_tiehi _11455__206 (.L_HI(net206));
 sg13g2_tiehi _11454__207 (.L_HI(net207));
 sg13g2_tiehi _11440__208 (.L_HI(net208));
 sg13g2_tiehi _11439__209 (.L_HI(net209));
 sg13g2_tiehi _11438__210 (.L_HI(net210));
 sg13g2_tiehi _11437__211 (.L_HI(net211));
 sg13g2_tiehi _11436__212 (.L_HI(net212));
 sg13g2_tiehi _11435__213 (.L_HI(net213));
 sg13g2_tiehi _11434__214 (.L_HI(net214));
 sg13g2_tiehi _11433__215 (.L_HI(net215));
 sg13g2_tiehi _11432__216 (.L_HI(net216));
 sg13g2_tiehi _11431__217 (.L_HI(net217));
 sg13g2_tiehi _11430__218 (.L_HI(net218));
 sg13g2_tiehi _11429__219 (.L_HI(net219));
 sg13g2_tiehi _11428__220 (.L_HI(net220));
 sg13g2_tiehi _11427__221 (.L_HI(net221));
 sg13g2_tiehi _11426__222 (.L_HI(net222));
 sg13g2_tiehi _11416__223 (.L_HI(net223));
 sg13g2_tiehi _11415__224 (.L_HI(net224));
 sg13g2_tiehi _11414__225 (.L_HI(net225));
 sg13g2_tiehi _11413__226 (.L_HI(net226));
 sg13g2_tiehi _12116__227 (.L_HI(net227));
 sg13g2_tiehi _11411__228 (.L_HI(net228));
 sg13g2_tiehi _12183__229 (.L_HI(net229));
 sg13g2_tiehi _11410__230 (.L_HI(net230));
 sg13g2_tiehi _12115__231 (.L_HI(net231));
 sg13g2_tiehi _11409__232 (.L_HI(net232));
 sg13g2_tiehi _12182__233 (.L_HI(net233));
 sg13g2_tiehi _11408__234 (.L_HI(net234));
 sg13g2_tiehi _12114__235 (.L_HI(net235));
 sg13g2_tiehi _11407__236 (.L_HI(net236));
 sg13g2_tiehi _12181__237 (.L_HI(net237));
 sg13g2_tiehi _11406__238 (.L_HI(net238));
 sg13g2_tiehi _12113__239 (.L_HI(net239));
 sg13g2_tiehi _11405__240 (.L_HI(net240));
 sg13g2_tiehi _12180__241 (.L_HI(net241));
 sg13g2_tiehi _11404__242 (.L_HI(net242));
 sg13g2_tiehi _12112__243 (.L_HI(net243));
 sg13g2_tiehi _11403__244 (.L_HI(net244));
 sg13g2_tiehi _12179__245 (.L_HI(net245));
 sg13g2_tiehi _11402__246 (.L_HI(net246));
 sg13g2_tiehi _12111__247 (.L_HI(net247));
 sg13g2_tiehi _11401__248 (.L_HI(net248));
 sg13g2_tiehi _12178__249 (.L_HI(net249));
 sg13g2_tiehi _11400__250 (.L_HI(net250));
 sg13g2_tiehi _12110__251 (.L_HI(net251));
 sg13g2_tiehi _11399__252 (.L_HI(net252));
 sg13g2_tiehi _12177__253 (.L_HI(net253));
 sg13g2_tiehi _11398__254 (.L_HI(net254));
 sg13g2_tiehi _12109__255 (.L_HI(net255));
 sg13g2_tiehi _11397__256 (.L_HI(net256));
 sg13g2_tiehi _12176__257 (.L_HI(net257));
 sg13g2_tiehi _11396__258 (.L_HI(net258));
 sg13g2_tiehi _12108__259 (.L_HI(net259));
 sg13g2_tiehi _11395__260 (.L_HI(net260));
 sg13g2_tiehi _11393__261 (.L_HI(net261));
 sg13g2_tiehi _11392__262 (.L_HI(net262));
 sg13g2_tiehi _11391__263 (.L_HI(net263));
 sg13g2_tiehi _11390__264 (.L_HI(net264));
 sg13g2_tiehi _11389__265 (.L_HI(net265));
 sg13g2_tiehi _11388__266 (.L_HI(net266));
 sg13g2_tiehi _11387__267 (.L_HI(net267));
 sg13g2_tiehi _11386__268 (.L_HI(net268));
 sg13g2_tiehi _11385__269 (.L_HI(net269));
 sg13g2_tiehi _11384__270 (.L_HI(net270));
 sg13g2_tiehi _11383__271 (.L_HI(net271));
 sg13g2_tiehi _11382__272 (.L_HI(net272));
 sg13g2_tiehi _11381__273 (.L_HI(net273));
 sg13g2_tiehi _11380__274 (.L_HI(net274));
 sg13g2_tiehi _11379__275 (.L_HI(net275));
 sg13g2_tiehi _11359__276 (.L_HI(net276));
 sg13g2_tiehi _11358__277 (.L_HI(net277));
 sg13g2_tiehi _11357__278 (.L_HI(net278));
 sg13g2_tiehi _11356__279 (.L_HI(net279));
 sg13g2_tiehi _11355__280 (.L_HI(net280));
 sg13g2_tiehi _11354__281 (.L_HI(net281));
 sg13g2_tiehi _11353__282 (.L_HI(net282));
 sg13g2_tiehi _11352__283 (.L_HI(net283));
 sg13g2_tiehi _11351__284 (.L_HI(net284));
 sg13g2_tiehi _11350__285 (.L_HI(net285));
 sg13g2_tiehi _11349__286 (.L_HI(net286));
 sg13g2_tiehi _11348__287 (.L_HI(net287));
 sg13g2_tiehi _11347__288 (.L_HI(net288));
 sg13g2_tiehi _11346__289 (.L_HI(net289));
 sg13g2_tiehi _11345__290 (.L_HI(net290));
 sg13g2_tiehi _11344__291 (.L_HI(net291));
 sg13g2_tiehi _11343__292 (.L_HI(net292));
 sg13g2_tiehi _11342__293 (.L_HI(net293));
 sg13g2_tiehi _11341__294 (.L_HI(net294));
 sg13g2_tiehi _11340__295 (.L_HI(net295));
 sg13g2_tiehi _11339__296 (.L_HI(net296));
 sg13g2_tiehi _11338__297 (.L_HI(net297));
 sg13g2_tiehi _11337__298 (.L_HI(net298));
 sg13g2_tiehi _11336__299 (.L_HI(net299));
 sg13g2_tiehi _11335__300 (.L_HI(net300));
 sg13g2_tiehi _11329__301 (.L_HI(net301));
 sg13g2_tiehi _11328__302 (.L_HI(net302));
 sg13g2_tiehi _11327__303 (.L_HI(net303));
 sg13g2_tiehi _11326__304 (.L_HI(net304));
 sg13g2_tiehi _11325__305 (.L_HI(net305));
 sg13g2_tiehi _11324__306 (.L_HI(net306));
 sg13g2_tiehi _11323__307 (.L_HI(net307));
 sg13g2_tiehi _11322__308 (.L_HI(net308));
 sg13g2_tiehi _11321__309 (.L_HI(net309));
 sg13g2_tiehi _11320__310 (.L_HI(net310));
 sg13g2_tiehi _11319__311 (.L_HI(net311));
 sg13g2_tiehi _11318__312 (.L_HI(net312));
 sg13g2_tiehi _11317__313 (.L_HI(net313));
 sg13g2_tiehi _11316__314 (.L_HI(net314));
 sg13g2_tiehi _11315__315 (.L_HI(net315));
 sg13g2_tiehi _11314__316 (.L_HI(net316));
 sg13g2_tiehi _11313__317 (.L_HI(net317));
 sg13g2_tiehi _11312__318 (.L_HI(net318));
 sg13g2_tiehi _11311__319 (.L_HI(net319));
 sg13g2_tiehi _11310__320 (.L_HI(net320));
 sg13g2_tiehi _11309__321 (.L_HI(net321));
 sg13g2_tiehi _11308__322 (.L_HI(net322));
 sg13g2_tiehi _11307__323 (.L_HI(net323));
 sg13g2_tiehi _11306__324 (.L_HI(net324));
 sg13g2_tiehi _11305__325 (.L_HI(net325));
 sg13g2_tiehi _11304__326 (.L_HI(net326));
 sg13g2_tiehi _11303__327 (.L_HI(net327));
 sg13g2_tiehi _11302__328 (.L_HI(net328));
 sg13g2_tiehi _11301__329 (.L_HI(net329));
 sg13g2_tiehi _11300__330 (.L_HI(net330));
 sg13g2_tiehi _11299__331 (.L_HI(net331));
 sg13g2_tiehi _11298__332 (.L_HI(net332));
 sg13g2_tiehi _12175__333 (.L_HI(net333));
 sg13g2_tiehi _12107__334 (.L_HI(net334));
 sg13g2_tiehi tt_um_dumbrv_yliu_hashed_335 (.L_HI(net335));
 sg13g2_tiehi tt_um_dumbrv_yliu_hashed_336 (.L_HI(net336));
 sg13g2_tiehi tt_um_dumbrv_yliu_hashed_337 (.L_HI(net337));
 sg13g2_tiehi tt_um_dumbrv_yliu_hashed_338 (.L_HI(net338));
 sg13g2_tiehi tt_um_dumbrv_yliu_hashed_339 (.L_HI(net339));
 sg13g2_tiehi tt_um_dumbrv_yliu_hashed_340 (.L_HI(net340));
 sg13g2_inv_1 _06169__1 (.Y(net341),
    .A(clknet_2_1__leaf_clk));
 sg13g2_tielo tt_um_dumbrv_yliu_hashed_12 (.L_LO(net12));
 sg13g2_tielo tt_um_dumbrv_yliu_hashed_13 (.L_LO(net13));
 sg13g2_tielo tt_um_dumbrv_yliu_hashed_14 (.L_LO(net14));
 sg13g2_tiehi _11639__15 (.L_HI(net15));
 sg13g2_buf_2 _12520_ (.A(\core.fetch.cmd_data[7] ),
    .X(uio_out[1]));
 sg13g2_buf_2 _12521_ (.A(net3573),
    .X(uio_out[3]));
 sg13g2_buf_2 _12522_ (.A(\core.lsu.spi.buffer[7] ),
    .X(uio_out[5]));
 sg13g2_buf_2 _12523_ (.A(net3522),
    .X(uio_out[7]));
 sg13g2_buf_2 fanout2714 (.A(net2715),
    .X(net2714));
 sg13g2_buf_2 fanout2715 (.A(net2716),
    .X(net2715));
 sg13g2_buf_2 fanout2716 (.A(net2718),
    .X(net2716));
 sg13g2_buf_2 fanout2717 (.A(net2718),
    .X(net2717));
 sg13g2_buf_1 fanout2718 (.A(net2730),
    .X(net2718));
 sg13g2_buf_2 fanout2719 (.A(net2720),
    .X(net2719));
 sg13g2_buf_2 fanout2720 (.A(net2723),
    .X(net2720));
 sg13g2_buf_2 fanout2721 (.A(net2723),
    .X(net2721));
 sg13g2_buf_1 fanout2722 (.A(net2723),
    .X(net2722));
 sg13g2_buf_2 fanout2723 (.A(net2730),
    .X(net2723));
 sg13g2_buf_2 fanout2724 (.A(net2725),
    .X(net2724));
 sg13g2_buf_2 fanout2725 (.A(net2726),
    .X(net2725));
 sg13g2_buf_1 fanout2726 (.A(net2730),
    .X(net2726));
 sg13g2_buf_2 fanout2727 (.A(net2729),
    .X(net2727));
 sg13g2_buf_2 fanout2728 (.A(net2729),
    .X(net2728));
 sg13g2_buf_2 fanout2729 (.A(net2730),
    .X(net2729));
 sg13g2_buf_2 fanout2730 (.A(_03019_),
    .X(net2730));
 sg13g2_buf_2 fanout2731 (.A(net2735),
    .X(net2731));
 sg13g2_buf_2 fanout2732 (.A(net2735),
    .X(net2732));
 sg13g2_buf_2 fanout2733 (.A(net2735),
    .X(net2733));
 sg13g2_buf_1 fanout2734 (.A(net2735),
    .X(net2734));
 sg13g2_buf_1 fanout2735 (.A(_01564_),
    .X(net2735));
 sg13g2_buf_4 fanout2736 (.X(net2736),
    .A(_01322_));
 sg13g2_buf_2 fanout2737 (.A(_01321_),
    .X(net2737));
 sg13g2_buf_2 fanout2738 (.A(net2741),
    .X(net2738));
 sg13g2_buf_2 fanout2739 (.A(net2741),
    .X(net2739));
 sg13g2_buf_1 fanout2740 (.A(net2741),
    .X(net2740));
 sg13g2_buf_1 fanout2741 (.A(_01321_),
    .X(net2741));
 sg13g2_buf_2 fanout2742 (.A(net2743),
    .X(net2742));
 sg13g2_buf_2 fanout2743 (.A(net2744),
    .X(net2743));
 sg13g2_buf_4 fanout2744 (.X(net2744),
    .A(net2751));
 sg13g2_buf_2 fanout2745 (.A(net2746),
    .X(net2745));
 sg13g2_buf_2 fanout2746 (.A(net2747),
    .X(net2746));
 sg13g2_buf_2 fanout2747 (.A(net2751),
    .X(net2747));
 sg13g2_buf_2 fanout2748 (.A(net2750),
    .X(net2748));
 sg13g2_buf_2 fanout2749 (.A(net2750),
    .X(net2749));
 sg13g2_buf_4 fanout2750 (.X(net2750),
    .A(net2751));
 sg13g2_buf_4 fanout2751 (.X(net2751),
    .A(_03965_));
 sg13g2_buf_2 fanout2752 (.A(net2756),
    .X(net2752));
 sg13g2_buf_2 fanout2753 (.A(net2756),
    .X(net2753));
 sg13g2_buf_4 fanout2754 (.X(net2754),
    .A(net2756));
 sg13g2_buf_2 fanout2755 (.A(net2756),
    .X(net2755));
 sg13g2_buf_2 fanout2756 (.A(_01464_),
    .X(net2756));
 sg13g2_buf_2 fanout2757 (.A(net2758),
    .X(net2757));
 sg13g2_buf_2 fanout2758 (.A(_02894_),
    .X(net2758));
 sg13g2_buf_2 fanout2759 (.A(net2761),
    .X(net2759));
 sg13g2_buf_2 fanout2760 (.A(net2761),
    .X(net2760));
 sg13g2_buf_2 fanout2761 (.A(_02894_),
    .X(net2761));
 sg13g2_buf_2 fanout2762 (.A(net2764),
    .X(net2762));
 sg13g2_buf_2 fanout2763 (.A(net2764),
    .X(net2763));
 sg13g2_buf_2 fanout2764 (.A(net2765),
    .X(net2764));
 sg13g2_buf_2 fanout2765 (.A(net2766),
    .X(net2765));
 sg13g2_buf_2 fanout2766 (.A(_03196_),
    .X(net2766));
 sg13g2_buf_2 fanout2767 (.A(net2768),
    .X(net2767));
 sg13g2_buf_2 fanout2768 (.A(_02777_),
    .X(net2768));
 sg13g2_buf_2 fanout2769 (.A(net2772),
    .X(net2769));
 sg13g2_buf_2 fanout2770 (.A(net2772),
    .X(net2770));
 sg13g2_buf_1 fanout2771 (.A(net2772),
    .X(net2771));
 sg13g2_buf_1 fanout2772 (.A(net2773),
    .X(net2772));
 sg13g2_buf_2 fanout2773 (.A(net2780),
    .X(net2773));
 sg13g2_buf_2 fanout2774 (.A(net2780),
    .X(net2774));
 sg13g2_buf_4 fanout2775 (.X(net2775),
    .A(net2779));
 sg13g2_buf_1 fanout2776 (.A(net2779),
    .X(net2776));
 sg13g2_buf_2 fanout2777 (.A(net2779),
    .X(net2777));
 sg13g2_buf_1 fanout2778 (.A(net2779),
    .X(net2778));
 sg13g2_buf_4 fanout2779 (.X(net2779),
    .A(net2780));
 sg13g2_buf_2 fanout2780 (.A(_01724_),
    .X(net2780));
 sg13g2_buf_2 fanout2781 (.A(net2784),
    .X(net2781));
 sg13g2_buf_1 fanout2782 (.A(net2784),
    .X(net2782));
 sg13g2_buf_2 fanout2783 (.A(net2784),
    .X(net2783));
 sg13g2_buf_4 fanout2784 (.X(net2784),
    .A(net2785));
 sg13g2_buf_2 fanout2785 (.A(_03194_),
    .X(net2785));
 sg13g2_buf_2 fanout2786 (.A(net2787),
    .X(net2786));
 sg13g2_buf_2 fanout2787 (.A(_02064_),
    .X(net2787));
 sg13g2_buf_4 fanout2788 (.X(net2788),
    .A(net2791));
 sg13g2_buf_2 fanout2789 (.A(net2791),
    .X(net2789));
 sg13g2_buf_4 fanout2790 (.X(net2790),
    .A(net2791));
 sg13g2_buf_2 fanout2791 (.A(_04006_),
    .X(net2791));
 sg13g2_buf_4 fanout2792 (.X(net2792),
    .A(net2793));
 sg13g2_buf_4 fanout2793 (.X(net2793),
    .A(_04005_));
 sg13g2_buf_2 fanout2794 (.A(net2797),
    .X(net2794));
 sg13g2_buf_2 fanout2795 (.A(net2796),
    .X(net2795));
 sg13g2_buf_2 fanout2796 (.A(net2797),
    .X(net2796));
 sg13g2_buf_2 fanout2797 (.A(_04005_),
    .X(net2797));
 sg13g2_buf_2 fanout2798 (.A(net2800),
    .X(net2798));
 sg13g2_buf_2 fanout2799 (.A(net2800),
    .X(net2799));
 sg13g2_buf_1 fanout2800 (.A(net2801),
    .X(net2800));
 sg13g2_buf_1 fanout2801 (.A(net2807),
    .X(net2801));
 sg13g2_buf_2 fanout2802 (.A(net2807),
    .X(net2802));
 sg13g2_buf_2 fanout2803 (.A(net2806),
    .X(net2803));
 sg13g2_buf_2 fanout2804 (.A(net2806),
    .X(net2804));
 sg13g2_buf_1 fanout2805 (.A(net2806),
    .X(net2805));
 sg13g2_buf_2 fanout2806 (.A(net2807),
    .X(net2806));
 sg13g2_buf_2 fanout2807 (.A(_02609_),
    .X(net2807));
 sg13g2_buf_2 fanout2808 (.A(net2812),
    .X(net2808));
 sg13g2_buf_1 fanout2809 (.A(net2812),
    .X(net2809));
 sg13g2_buf_2 fanout2810 (.A(net2812),
    .X(net2810));
 sg13g2_buf_2 fanout2811 (.A(net2812),
    .X(net2811));
 sg13g2_buf_1 fanout2812 (.A(net2815),
    .X(net2812));
 sg13g2_buf_2 fanout2813 (.A(net2815),
    .X(net2813));
 sg13g2_buf_2 fanout2814 (.A(net2815),
    .X(net2814));
 sg13g2_buf_2 fanout2815 (.A(_02440_),
    .X(net2815));
 sg13g2_buf_2 fanout2816 (.A(net2820),
    .X(net2816));
 sg13g2_buf_1 fanout2817 (.A(net2820),
    .X(net2817));
 sg13g2_buf_2 fanout2818 (.A(net2820),
    .X(net2818));
 sg13g2_buf_1 fanout2819 (.A(net2820),
    .X(net2819));
 sg13g2_buf_2 fanout2820 (.A(_02440_),
    .X(net2820));
 sg13g2_buf_2 fanout2821 (.A(net2822),
    .X(net2821));
 sg13g2_buf_2 fanout2822 (.A(_04092_),
    .X(net2822));
 sg13g2_buf_2 fanout2823 (.A(_04092_),
    .X(net2823));
 sg13g2_buf_2 fanout2824 (.A(_04092_),
    .X(net2824));
 sg13g2_buf_4 fanout2825 (.X(net2825),
    .A(net2828));
 sg13g2_buf_4 fanout2826 (.X(net2826),
    .A(net2828));
 sg13g2_buf_1 fanout2827 (.A(net2828),
    .X(net2827));
 sg13g2_buf_2 fanout2828 (.A(_04016_),
    .X(net2828));
 sg13g2_buf_2 fanout2829 (.A(_04009_),
    .X(net2829));
 sg13g2_buf_1 fanout2830 (.A(_04009_),
    .X(net2830));
 sg13g2_buf_2 fanout2831 (.A(net2832),
    .X(net2831));
 sg13g2_buf_4 fanout2832 (.X(net2832),
    .A(_04009_));
 sg13g2_buf_2 fanout2833 (.A(net2834),
    .X(net2833));
 sg13g2_buf_2 fanout2834 (.A(_03991_),
    .X(net2834));
 sg13g2_buf_2 fanout2835 (.A(_03991_),
    .X(net2835));
 sg13g2_buf_2 fanout2836 (.A(_03464_),
    .X(net2836));
 sg13g2_buf_4 fanout2837 (.X(net2837),
    .A(net2839));
 sg13g2_buf_1 fanout2838 (.A(net2839),
    .X(net2838));
 sg13g2_buf_2 fanout2839 (.A(_02450_),
    .X(net2839));
 sg13g2_buf_4 fanout2840 (.X(net2840),
    .A(_02134_));
 sg13g2_buf_2 fanout2841 (.A(net2844),
    .X(net2841));
 sg13g2_buf_1 fanout2842 (.A(net2844),
    .X(net2842));
 sg13g2_buf_4 fanout2843 (.X(net2843),
    .A(net2844));
 sg13g2_buf_4 fanout2844 (.X(net2844),
    .A(_02133_));
 sg13g2_buf_2 fanout2845 (.A(_01361_),
    .X(net2845));
 sg13g2_buf_2 fanout2846 (.A(_01361_),
    .X(net2846));
 sg13g2_buf_2 fanout2847 (.A(net2848),
    .X(net2847));
 sg13g2_buf_2 fanout2848 (.A(_01351_),
    .X(net2848));
 sg13g2_buf_2 fanout2849 (.A(_01343_),
    .X(net2849));
 sg13g2_buf_2 fanout2850 (.A(_01343_),
    .X(net2850));
 sg13g2_buf_2 fanout2851 (.A(_04205_),
    .X(net2851));
 sg13g2_buf_2 fanout2852 (.A(_04127_),
    .X(net2852));
 sg13g2_buf_4 fanout2853 (.X(net2853),
    .A(_03989_));
 sg13g2_buf_4 fanout2854 (.X(net2854),
    .A(net2856));
 sg13g2_buf_2 fanout2855 (.A(net2856),
    .X(net2855));
 sg13g2_buf_2 fanout2856 (.A(net2858),
    .X(net2856));
 sg13g2_buf_4 fanout2857 (.X(net2857),
    .A(net2858));
 sg13g2_buf_2 fanout2858 (.A(_03971_),
    .X(net2858));
 sg13g2_buf_4 fanout2859 (.X(net2859),
    .A(net2860));
 sg13g2_buf_4 fanout2860 (.X(net2860),
    .A(_03970_));
 sg13g2_buf_2 fanout2861 (.A(_03463_),
    .X(net2861));
 sg13g2_buf_4 fanout2862 (.X(net2862),
    .A(_02518_));
 sg13g2_buf_4 fanout2863 (.X(net2863),
    .A(_02494_));
 sg13g2_buf_2 fanout2864 (.A(net2867),
    .X(net2864));
 sg13g2_buf_2 fanout2865 (.A(net2866),
    .X(net2865));
 sg13g2_buf_2 fanout2866 (.A(net2867),
    .X(net2866));
 sg13g2_buf_1 fanout2867 (.A(net2868),
    .X(net2867));
 sg13g2_buf_1 fanout2868 (.A(_02494_),
    .X(net2868));
 sg13g2_buf_2 fanout2869 (.A(net2871),
    .X(net2869));
 sg13g2_buf_1 fanout2870 (.A(net2871),
    .X(net2870));
 sg13g2_buf_2 fanout2871 (.A(net2872),
    .X(net2871));
 sg13g2_buf_4 fanout2872 (.X(net2872),
    .A(net2875));
 sg13g2_buf_4 fanout2873 (.X(net2873),
    .A(net2874));
 sg13g2_buf_4 fanout2874 (.X(net2874),
    .A(net2875));
 sg13g2_buf_4 fanout2875 (.X(net2875),
    .A(_02432_));
 sg13g2_buf_4 fanout2876 (.X(net2876),
    .A(net2877));
 sg13g2_buf_4 fanout2877 (.X(net2877),
    .A(_02432_));
 sg13g2_buf_4 fanout2878 (.X(net2878),
    .A(net2879));
 sg13g2_buf_2 fanout2879 (.A(_02432_),
    .X(net2879));
 sg13g2_buf_2 fanout2880 (.A(net2882),
    .X(net2880));
 sg13g2_buf_1 fanout2881 (.A(net2882),
    .X(net2881));
 sg13g2_buf_2 fanout2882 (.A(net2885),
    .X(net2882));
 sg13g2_buf_2 fanout2883 (.A(net2884),
    .X(net2883));
 sg13g2_buf_2 fanout2884 (.A(net2885),
    .X(net2884));
 sg13g2_buf_1 fanout2885 (.A(_02420_),
    .X(net2885));
 sg13g2_buf_2 fanout2886 (.A(net2887),
    .X(net2886));
 sg13g2_buf_2 fanout2887 (.A(net2888),
    .X(net2887));
 sg13g2_buf_2 fanout2888 (.A(_02420_),
    .X(net2888));
 sg13g2_buf_2 fanout2889 (.A(_02132_),
    .X(net2889));
 sg13g2_buf_1 fanout2890 (.A(_02132_),
    .X(net2890));
 sg13g2_buf_2 fanout2891 (.A(net2892),
    .X(net2891));
 sg13g2_buf_2 fanout2892 (.A(net2893),
    .X(net2892));
 sg13g2_buf_2 fanout2893 (.A(_01995_),
    .X(net2893));
 sg13g2_buf_2 fanout2894 (.A(net2895),
    .X(net2894));
 sg13g2_buf_2 fanout2895 (.A(net2896),
    .X(net2895));
 sg13g2_buf_2 fanout2896 (.A(_01978_),
    .X(net2896));
 sg13g2_buf_2 fanout2897 (.A(net2898),
    .X(net2897));
 sg13g2_buf_2 fanout2898 (.A(net2899),
    .X(net2898));
 sg13g2_buf_2 fanout2899 (.A(net2902),
    .X(net2899));
 sg13g2_buf_2 fanout2900 (.A(net2901),
    .X(net2900));
 sg13g2_buf_2 fanout2901 (.A(net2902),
    .X(net2901));
 sg13g2_buf_2 fanout2902 (.A(net2904),
    .X(net2902));
 sg13g2_buf_2 fanout2903 (.A(net2904),
    .X(net2903));
 sg13g2_buf_2 fanout2904 (.A(_01728_),
    .X(net2904));
 sg13g2_buf_2 fanout2905 (.A(net2907),
    .X(net2905));
 sg13g2_buf_1 fanout2906 (.A(net2907),
    .X(net2906));
 sg13g2_buf_2 fanout2907 (.A(_01728_),
    .X(net2907));
 sg13g2_buf_4 fanout2908 (.X(net2908),
    .A(_01727_));
 sg13g2_buf_4 fanout2909 (.X(net2909),
    .A(net2911));
 sg13g2_buf_2 fanout2910 (.A(net2911),
    .X(net2910));
 sg13g2_buf_2 fanout2911 (.A(_01726_),
    .X(net2911));
 sg13g2_buf_8 fanout2912 (.A(_01688_),
    .X(net2912));
 sg13g2_buf_2 fanout2913 (.A(net2914),
    .X(net2913));
 sg13g2_buf_2 fanout2914 (.A(net2915),
    .X(net2914));
 sg13g2_buf_2 fanout2915 (.A(net2921),
    .X(net2915));
 sg13g2_buf_2 fanout2916 (.A(net2918),
    .X(net2916));
 sg13g2_buf_1 fanout2917 (.A(net2918),
    .X(net2917));
 sg13g2_buf_2 fanout2918 (.A(net2921),
    .X(net2918));
 sg13g2_buf_2 fanout2919 (.A(net2920),
    .X(net2919));
 sg13g2_buf_2 fanout2920 (.A(net2921),
    .X(net2920));
 sg13g2_buf_2 fanout2921 (.A(_01687_),
    .X(net2921));
 sg13g2_buf_4 fanout2922 (.X(net2922),
    .A(_01683_));
 sg13g2_buf_1 fanout2923 (.A(_01683_),
    .X(net2923));
 sg13g2_buf_4 fanout2924 (.X(net2924),
    .A(_04012_));
 sg13g2_buf_4 fanout2925 (.X(net2925),
    .A(net2926));
 sg13g2_buf_2 fanout2926 (.A(_04011_),
    .X(net2926));
 sg13g2_buf_4 fanout2927 (.X(net2927),
    .A(_04011_));
 sg13g2_buf_4 fanout2928 (.X(net2928),
    .A(net2929));
 sg13g2_buf_2 fanout2929 (.A(_03994_),
    .X(net2929));
 sg13g2_buf_2 fanout2930 (.A(net2931),
    .X(net2930));
 sg13g2_buf_2 fanout2931 (.A(net2932),
    .X(net2931));
 sg13g2_buf_2 fanout2932 (.A(_03993_),
    .X(net2932));
 sg13g2_buf_2 fanout2933 (.A(net2934),
    .X(net2933));
 sg13g2_buf_2 fanout2934 (.A(net2936),
    .X(net2934));
 sg13g2_buf_2 fanout2935 (.A(net2936),
    .X(net2935));
 sg13g2_buf_2 fanout2936 (.A(_03993_),
    .X(net2936));
 sg13g2_buf_2 fanout2937 (.A(net2938),
    .X(net2937));
 sg13g2_buf_4 fanout2938 (.X(net2938),
    .A(net2941));
 sg13g2_buf_4 fanout2939 (.X(net2939),
    .A(net2941));
 sg13g2_buf_4 fanout2940 (.X(net2940),
    .A(net2941));
 sg13g2_buf_2 fanout2941 (.A(_03981_),
    .X(net2941));
 sg13g2_buf_2 fanout2942 (.A(net2944),
    .X(net2942));
 sg13g2_buf_2 fanout2943 (.A(net2944),
    .X(net2943));
 sg13g2_buf_2 fanout2944 (.A(net2948),
    .X(net2944));
 sg13g2_buf_2 fanout2945 (.A(net2946),
    .X(net2945));
 sg13g2_buf_2 fanout2946 (.A(net2948),
    .X(net2946));
 sg13g2_buf_2 fanout2947 (.A(net2948),
    .X(net2947));
 sg13g2_buf_2 fanout2948 (.A(_03980_),
    .X(net2948));
 sg13g2_buf_4 fanout2949 (.X(net2949),
    .A(net2950));
 sg13g2_buf_2 fanout2950 (.A(net2951),
    .X(net2950));
 sg13g2_buf_4 fanout2951 (.X(net2951),
    .A(_03979_));
 sg13g2_buf_4 fanout2952 (.X(net2952),
    .A(net2953));
 sg13g2_buf_4 fanout2953 (.X(net2953),
    .A(_03978_));
 sg13g2_buf_4 fanout2954 (.X(net2954),
    .A(_03977_));
 sg13g2_buf_4 fanout2955 (.X(net2955),
    .A(_03977_));
 sg13g2_buf_2 fanout2956 (.A(net2957),
    .X(net2956));
 sg13g2_buf_2 fanout2957 (.A(net2958),
    .X(net2957));
 sg13g2_buf_2 fanout2958 (.A(net2961),
    .X(net2958));
 sg13g2_buf_2 fanout2959 (.A(net2960),
    .X(net2959));
 sg13g2_buf_2 fanout2960 (.A(net2961),
    .X(net2960));
 sg13g2_buf_2 fanout2961 (.A(net2966),
    .X(net2961));
 sg13g2_buf_2 fanout2962 (.A(net2963),
    .X(net2962));
 sg13g2_buf_2 fanout2963 (.A(net2966),
    .X(net2963));
 sg13g2_buf_2 fanout2964 (.A(net2965),
    .X(net2964));
 sg13g2_buf_2 fanout2965 (.A(net2966),
    .X(net2965));
 sg13g2_buf_2 fanout2966 (.A(_03969_),
    .X(net2966));
 sg13g2_buf_2 fanout2967 (.A(net2972),
    .X(net2967));
 sg13g2_buf_2 fanout2968 (.A(net2972),
    .X(net2968));
 sg13g2_buf_2 fanout2969 (.A(net2971),
    .X(net2969));
 sg13g2_buf_2 fanout2970 (.A(net2971),
    .X(net2970));
 sg13g2_buf_2 fanout2971 (.A(net2972),
    .X(net2971));
 sg13g2_buf_2 fanout2972 (.A(_02613_),
    .X(net2972));
 sg13g2_buf_2 fanout2973 (.A(net2975),
    .X(net2973));
 sg13g2_buf_2 fanout2974 (.A(net2975),
    .X(net2974));
 sg13g2_buf_2 fanout2975 (.A(_02578_),
    .X(net2975));
 sg13g2_buf_2 fanout2976 (.A(_02523_),
    .X(net2976));
 sg13g2_buf_2 fanout2977 (.A(net2978),
    .X(net2977));
 sg13g2_buf_2 fanout2978 (.A(_02521_),
    .X(net2978));
 sg13g2_buf_2 fanout2979 (.A(net2980),
    .X(net2979));
 sg13g2_buf_2 fanout2980 (.A(_02517_),
    .X(net2980));
 sg13g2_buf_2 fanout2981 (.A(_02511_),
    .X(net2981));
 sg13g2_buf_2 fanout2982 (.A(_02511_),
    .X(net2982));
 sg13g2_buf_4 fanout2983 (.X(net2983),
    .A(net2984));
 sg13g2_buf_4 fanout2984 (.X(net2984),
    .A(net2987));
 sg13g2_buf_4 fanout2985 (.X(net2985),
    .A(net2987));
 sg13g2_buf_4 fanout2986 (.X(net2986),
    .A(net2987));
 sg13g2_buf_4 fanout2987 (.X(net2987),
    .A(_01751_));
 sg13g2_buf_4 fanout2988 (.X(net2988),
    .A(net2989));
 sg13g2_buf_4 fanout2989 (.X(net2989),
    .A(net2992));
 sg13g2_buf_4 fanout2990 (.X(net2990),
    .A(net2992));
 sg13g2_buf_4 fanout2991 (.X(net2991),
    .A(net2992));
 sg13g2_buf_4 fanout2992 (.X(net2992),
    .A(_01749_));
 sg13g2_buf_4 fanout2993 (.X(net2993),
    .A(net2994));
 sg13g2_buf_4 fanout2994 (.X(net2994),
    .A(net2997));
 sg13g2_buf_4 fanout2995 (.X(net2995),
    .A(net2997));
 sg13g2_buf_4 fanout2996 (.X(net2996),
    .A(net2997));
 sg13g2_buf_4 fanout2997 (.X(net2997),
    .A(_01748_));
 sg13g2_buf_4 fanout2998 (.X(net2998),
    .A(net2999));
 sg13g2_buf_4 fanout2999 (.X(net2999),
    .A(net3002));
 sg13g2_buf_4 fanout3000 (.X(net3000),
    .A(net3002));
 sg13g2_buf_4 fanout3001 (.X(net3001),
    .A(net3002));
 sg13g2_buf_4 fanout3002 (.X(net3002),
    .A(_01745_));
 sg13g2_buf_4 fanout3003 (.X(net3003),
    .A(net3004));
 sg13g2_buf_4 fanout3004 (.X(net3004),
    .A(net3007));
 sg13g2_buf_4 fanout3005 (.X(net3005),
    .A(net3007));
 sg13g2_buf_4 fanout3006 (.X(net3006),
    .A(net3007));
 sg13g2_buf_4 fanout3007 (.X(net3007),
    .A(_01744_));
 sg13g2_buf_4 fanout3008 (.X(net3008),
    .A(net3009));
 sg13g2_buf_4 fanout3009 (.X(net3009),
    .A(net3012));
 sg13g2_buf_4 fanout3010 (.X(net3010),
    .A(net3012));
 sg13g2_buf_4 fanout3011 (.X(net3011),
    .A(net3012));
 sg13g2_buf_4 fanout3012 (.X(net3012),
    .A(_01741_));
 sg13g2_buf_4 fanout3013 (.X(net3013),
    .A(net3014));
 sg13g2_buf_4 fanout3014 (.X(net3014),
    .A(net3017));
 sg13g2_buf_4 fanout3015 (.X(net3015),
    .A(net3017));
 sg13g2_buf_4 fanout3016 (.X(net3016),
    .A(net3017));
 sg13g2_buf_4 fanout3017 (.X(net3017),
    .A(_01738_));
 sg13g2_buf_4 fanout3018 (.X(net3018),
    .A(net3019));
 sg13g2_buf_4 fanout3019 (.X(net3019),
    .A(net3022));
 sg13g2_buf_4 fanout3020 (.X(net3020),
    .A(net3022));
 sg13g2_buf_4 fanout3021 (.X(net3021),
    .A(net3022));
 sg13g2_buf_2 fanout3022 (.A(_01737_),
    .X(net3022));
 sg13g2_buf_4 fanout3023 (.X(net3023),
    .A(net3024));
 sg13g2_buf_4 fanout3024 (.X(net3024),
    .A(net3027));
 sg13g2_buf_4 fanout3025 (.X(net3025),
    .A(net3027));
 sg13g2_buf_4 fanout3026 (.X(net3026),
    .A(net3027));
 sg13g2_buf_4 fanout3027 (.X(net3027),
    .A(_01734_));
 sg13g2_buf_2 fanout3028 (.A(net3030),
    .X(net3028));
 sg13g2_buf_2 fanout3029 (.A(net3030),
    .X(net3029));
 sg13g2_buf_4 fanout3030 (.X(net3030),
    .A(_01725_));
 sg13g2_buf_4 fanout3031 (.X(net3031),
    .A(_01669_));
 sg13g2_buf_2 fanout3032 (.A(net3033),
    .X(net3032));
 sg13g2_buf_2 fanout3033 (.A(net3034),
    .X(net3033));
 sg13g2_buf_4 fanout3034 (.X(net3034),
    .A(_01668_));
 sg13g2_buf_4 fanout3035 (.X(net3035),
    .A(net3036));
 sg13g2_buf_4 fanout3036 (.X(net3036),
    .A(_01668_));
 sg13g2_buf_2 fanout3037 (.A(net3038),
    .X(net3037));
 sg13g2_buf_2 fanout3038 (.A(_01667_),
    .X(net3038));
 sg13g2_buf_2 fanout3039 (.A(_01392_),
    .X(net3039));
 sg13g2_buf_2 fanout3040 (.A(net3041),
    .X(net3040));
 sg13g2_buf_2 fanout3041 (.A(net3042),
    .X(net3041));
 sg13g2_buf_1 fanout3042 (.A(_01372_),
    .X(net3042));
 sg13g2_buf_2 fanout3043 (.A(net3045),
    .X(net3043));
 sg13g2_buf_2 fanout3044 (.A(net3045),
    .X(net3044));
 sg13g2_buf_2 fanout3045 (.A(_01328_),
    .X(net3045));
 sg13g2_buf_4 fanout3046 (.X(net3046),
    .A(net3047));
 sg13g2_buf_4 fanout3047 (.X(net3047),
    .A(_05367_));
 sg13g2_buf_2 fanout3048 (.A(net3050),
    .X(net3048));
 sg13g2_buf_2 fanout3049 (.A(net3050),
    .X(net3049));
 sg13g2_buf_2 fanout3050 (.A(_05276_),
    .X(net3050));
 sg13g2_buf_2 fanout3051 (.A(net3052),
    .X(net3051));
 sg13g2_buf_4 fanout3052 (.X(net3052),
    .A(_05251_));
 sg13g2_buf_4 fanout3053 (.X(net3053),
    .A(_04022_));
 sg13g2_buf_2 fanout3054 (.A(_04022_),
    .X(net3054));
 sg13g2_buf_2 fanout3055 (.A(net3056),
    .X(net3055));
 sg13g2_buf_2 fanout3056 (.A(net3057),
    .X(net3056));
 sg13g2_buf_2 fanout3057 (.A(_03987_),
    .X(net3057));
 sg13g2_buf_2 fanout3058 (.A(net3059),
    .X(net3058));
 sg13g2_buf_1 fanout3059 (.A(net3060),
    .X(net3059));
 sg13g2_buf_4 fanout3060 (.X(net3060),
    .A(_03987_));
 sg13g2_buf_2 fanout3061 (.A(net3062),
    .X(net3061));
 sg13g2_buf_2 fanout3062 (.A(net3063),
    .X(net3062));
 sg13g2_buf_2 fanout3063 (.A(_03986_),
    .X(net3063));
 sg13g2_buf_2 fanout3064 (.A(_03986_),
    .X(net3064));
 sg13g2_buf_2 fanout3065 (.A(_03986_),
    .X(net3065));
 sg13g2_buf_4 fanout3066 (.X(net3066),
    .A(net3067));
 sg13g2_buf_4 fanout3067 (.X(net3067),
    .A(net3070));
 sg13g2_buf_4 fanout3068 (.X(net3068),
    .A(net3069));
 sg13g2_buf_4 fanout3069 (.X(net3069),
    .A(net3070));
 sg13g2_buf_4 fanout3070 (.X(net3070),
    .A(_03221_));
 sg13g2_buf_4 fanout3071 (.X(net3071),
    .A(net3072));
 sg13g2_buf_4 fanout3072 (.X(net3072),
    .A(net3075));
 sg13g2_buf_4 fanout3073 (.X(net3073),
    .A(net3075));
 sg13g2_buf_4 fanout3074 (.X(net3074),
    .A(net3075));
 sg13g2_buf_4 fanout3075 (.X(net3075),
    .A(_03220_));
 sg13g2_buf_4 fanout3076 (.X(net3076),
    .A(net3077));
 sg13g2_buf_4 fanout3077 (.X(net3077),
    .A(net3080));
 sg13g2_buf_4 fanout3078 (.X(net3078),
    .A(net3080));
 sg13g2_buf_4 fanout3079 (.X(net3079),
    .A(net3080));
 sg13g2_buf_4 fanout3080 (.X(net3080),
    .A(_03219_));
 sg13g2_buf_4 fanout3081 (.X(net3081),
    .A(net3082));
 sg13g2_buf_4 fanout3082 (.X(net3082),
    .A(net3085));
 sg13g2_buf_4 fanout3083 (.X(net3083),
    .A(net3085));
 sg13g2_buf_4 fanout3084 (.X(net3084),
    .A(net3085));
 sg13g2_buf_4 fanout3085 (.X(net3085),
    .A(_03218_));
 sg13g2_buf_4 fanout3086 (.X(net3086),
    .A(net3087));
 sg13g2_buf_4 fanout3087 (.X(net3087),
    .A(net3090));
 sg13g2_buf_4 fanout3088 (.X(net3088),
    .A(net3090));
 sg13g2_buf_4 fanout3089 (.X(net3089),
    .A(net3090));
 sg13g2_buf_4 fanout3090 (.X(net3090),
    .A(_03216_));
 sg13g2_buf_4 fanout3091 (.X(net3091),
    .A(net3092));
 sg13g2_buf_4 fanout3092 (.X(net3092),
    .A(net3095));
 sg13g2_buf_4 fanout3093 (.X(net3093),
    .A(net3095));
 sg13g2_buf_4 fanout3094 (.X(net3094),
    .A(net3095));
 sg13g2_buf_4 fanout3095 (.X(net3095),
    .A(_03214_));
 sg13g2_buf_4 fanout3096 (.X(net3096),
    .A(net3097));
 sg13g2_buf_4 fanout3097 (.X(net3097),
    .A(net3100));
 sg13g2_buf_4 fanout3098 (.X(net3098),
    .A(net3100));
 sg13g2_buf_2 fanout3099 (.A(net3100),
    .X(net3099));
 sg13g2_buf_4 fanout3100 (.X(net3100),
    .A(_03213_));
 sg13g2_buf_4 fanout3101 (.X(net3101),
    .A(net3102));
 sg13g2_buf_4 fanout3102 (.X(net3102),
    .A(net3105));
 sg13g2_buf_4 fanout3103 (.X(net3103),
    .A(net3105));
 sg13g2_buf_4 fanout3104 (.X(net3104),
    .A(net3105));
 sg13g2_buf_4 fanout3105 (.X(net3105),
    .A(_03212_));
 sg13g2_buf_4 fanout3106 (.X(net3106),
    .A(net3107));
 sg13g2_buf_4 fanout3107 (.X(net3107),
    .A(net3110));
 sg13g2_buf_4 fanout3108 (.X(net3108),
    .A(net3110));
 sg13g2_buf_4 fanout3109 (.X(net3109),
    .A(net3110));
 sg13g2_buf_4 fanout3110 (.X(net3110),
    .A(_03210_));
 sg13g2_buf_4 fanout3111 (.X(net3111),
    .A(net3112));
 sg13g2_buf_4 fanout3112 (.X(net3112),
    .A(net3115));
 sg13g2_buf_4 fanout3113 (.X(net3113),
    .A(net3115));
 sg13g2_buf_2 fanout3114 (.A(net3115),
    .X(net3114));
 sg13g2_buf_4 fanout3115 (.X(net3115),
    .A(_03208_));
 sg13g2_buf_4 fanout3116 (.X(net3116),
    .A(net3117));
 sg13g2_buf_4 fanout3117 (.X(net3117),
    .A(net3120));
 sg13g2_buf_4 fanout3118 (.X(net3118),
    .A(net3120));
 sg13g2_buf_4 fanout3119 (.X(net3119),
    .A(net3120));
 sg13g2_buf_4 fanout3120 (.X(net3120),
    .A(_03207_));
 sg13g2_buf_4 fanout3121 (.X(net3121),
    .A(net3122));
 sg13g2_buf_4 fanout3122 (.X(net3122),
    .A(net3125));
 sg13g2_buf_4 fanout3123 (.X(net3123),
    .A(net3124));
 sg13g2_buf_4 fanout3124 (.X(net3124),
    .A(net3125));
 sg13g2_buf_4 fanout3125 (.X(net3125),
    .A(_03206_));
 sg13g2_buf_4 fanout3126 (.X(net3126),
    .A(net3127));
 sg13g2_buf_4 fanout3127 (.X(net3127),
    .A(net3130));
 sg13g2_buf_4 fanout3128 (.X(net3128),
    .A(net3129));
 sg13g2_buf_4 fanout3129 (.X(net3129),
    .A(net3130));
 sg13g2_buf_4 fanout3130 (.X(net3130),
    .A(_03203_));
 sg13g2_buf_4 fanout3131 (.X(net3131),
    .A(net3132));
 sg13g2_buf_4 fanout3132 (.X(net3132),
    .A(net3135));
 sg13g2_buf_4 fanout3133 (.X(net3133),
    .A(net3135));
 sg13g2_buf_4 fanout3134 (.X(net3134),
    .A(net3135));
 sg13g2_buf_4 fanout3135 (.X(net3135),
    .A(_03201_));
 sg13g2_buf_4 fanout3136 (.X(net3136),
    .A(net3137));
 sg13g2_buf_2 fanout3137 (.A(_03115_),
    .X(net3137));
 sg13g2_buf_2 fanout3138 (.A(_03070_),
    .X(net3138));
 sg13g2_buf_2 fanout3139 (.A(_03070_),
    .X(net3139));
 sg13g2_buf_2 fanout3140 (.A(net3141),
    .X(net3140));
 sg13g2_buf_2 fanout3141 (.A(_03021_),
    .X(net3141));
 sg13g2_buf_2 fanout3142 (.A(_02793_),
    .X(net3142));
 sg13g2_buf_2 fanout3143 (.A(_02793_),
    .X(net3143));
 sg13g2_buf_2 fanout3144 (.A(_02782_),
    .X(net3144));
 sg13g2_buf_2 fanout3145 (.A(_02723_),
    .X(net3145));
 sg13g2_buf_2 fanout3146 (.A(_02723_),
    .X(net3146));
 sg13g2_buf_2 fanout3147 (.A(net3149),
    .X(net3147));
 sg13g2_buf_1 fanout3148 (.A(net3149),
    .X(net3148));
 sg13g2_buf_2 fanout3149 (.A(net3150),
    .X(net3149));
 sg13g2_buf_2 fanout3150 (.A(_02579_),
    .X(net3150));
 sg13g2_buf_2 fanout3151 (.A(_02573_),
    .X(net3151));
 sg13g2_buf_1 fanout3152 (.A(_02573_),
    .X(net3152));
 sg13g2_buf_2 fanout3153 (.A(net3154),
    .X(net3153));
 sg13g2_buf_2 fanout3154 (.A(net3155),
    .X(net3154));
 sg13g2_buf_2 fanout3155 (.A(net3156),
    .X(net3155));
 sg13g2_buf_4 fanout3156 (.X(net3156),
    .A(_02572_));
 sg13g2_buf_2 fanout3157 (.A(_02525_),
    .X(net3157));
 sg13g2_buf_4 fanout3158 (.X(net3158),
    .A(net3159));
 sg13g2_buf_2 fanout3159 (.A(_02455_),
    .X(net3159));
 sg13g2_buf_4 fanout3160 (.X(net3160),
    .A(net3161));
 sg13g2_buf_4 fanout3161 (.X(net3161),
    .A(_01768_));
 sg13g2_buf_4 fanout3162 (.X(net3162),
    .A(net3163));
 sg13g2_buf_2 fanout3163 (.A(net3164),
    .X(net3163));
 sg13g2_buf_4 fanout3164 (.X(net3164),
    .A(_01767_));
 sg13g2_buf_4 fanout3165 (.X(net3165),
    .A(net3168));
 sg13g2_buf_1 fanout3166 (.A(net3168),
    .X(net3166));
 sg13g2_buf_2 fanout3167 (.A(net3168),
    .X(net3167));
 sg13g2_buf_2 fanout3168 (.A(_01767_),
    .X(net3168));
 sg13g2_buf_4 fanout3169 (.X(net3169),
    .A(net3170));
 sg13g2_buf_4 fanout3170 (.X(net3170),
    .A(net3173));
 sg13g2_buf_4 fanout3171 (.X(net3171),
    .A(net3173));
 sg13g2_buf_4 fanout3172 (.X(net3172),
    .A(net3173));
 sg13g2_buf_4 fanout3173 (.X(net3173),
    .A(_01752_));
 sg13g2_buf_4 fanout3174 (.X(net3174),
    .A(net3175));
 sg13g2_buf_4 fanout3175 (.X(net3175),
    .A(net3178));
 sg13g2_buf_4 fanout3176 (.X(net3176),
    .A(net3177));
 sg13g2_buf_4 fanout3177 (.X(net3177),
    .A(net3178));
 sg13g2_buf_4 fanout3178 (.X(net3178),
    .A(_01747_));
 sg13g2_buf_4 fanout3179 (.X(net3179),
    .A(net3180));
 sg13g2_buf_4 fanout3180 (.X(net3180),
    .A(net3183));
 sg13g2_buf_4 fanout3181 (.X(net3181),
    .A(net3183));
 sg13g2_buf_4 fanout3182 (.X(net3182),
    .A(net3183));
 sg13g2_buf_4 fanout3183 (.X(net3183),
    .A(_01746_));
 sg13g2_buf_4 fanout3184 (.X(net3184),
    .A(net3185));
 sg13g2_buf_4 fanout3185 (.X(net3185),
    .A(net3188));
 sg13g2_buf_4 fanout3186 (.X(net3186),
    .A(net3188));
 sg13g2_buf_2 fanout3187 (.A(net3188),
    .X(net3187));
 sg13g2_buf_4 fanout3188 (.X(net3188),
    .A(_01743_));
 sg13g2_buf_4 fanout3189 (.X(net3189),
    .A(net3190));
 sg13g2_buf_4 fanout3190 (.X(net3190),
    .A(net3193));
 sg13g2_buf_4 fanout3191 (.X(net3191),
    .A(net3193));
 sg13g2_buf_4 fanout3192 (.X(net3192),
    .A(net3193));
 sg13g2_buf_4 fanout3193 (.X(net3193),
    .A(_01739_));
 sg13g2_buf_2 fanout3194 (.A(net3195),
    .X(net3194));
 sg13g2_buf_4 fanout3195 (.X(net3195),
    .A(net3196));
 sg13g2_buf_4 fanout3196 (.X(net3196),
    .A(_01692_));
 sg13g2_buf_2 fanout3197 (.A(net3198),
    .X(net3197));
 sg13g2_buf_2 fanout3198 (.A(_01657_),
    .X(net3198));
 sg13g2_buf_4 fanout3199 (.X(net3199),
    .A(_01657_));
 sg13g2_buf_2 fanout3200 (.A(_01394_),
    .X(net3200));
 sg13g2_buf_2 fanout3201 (.A(net3203),
    .X(net3201));
 sg13g2_buf_2 fanout3202 (.A(net3203),
    .X(net3202));
 sg13g2_buf_2 fanout3203 (.A(_01142_),
    .X(net3203));
 sg13g2_buf_2 fanout3204 (.A(net3205),
    .X(net3204));
 sg13g2_buf_2 fanout3205 (.A(_01142_),
    .X(net3205));
 sg13g2_buf_2 fanout3206 (.A(_00981_),
    .X(net3206));
 sg13g2_buf_4 fanout3207 (.X(net3207),
    .A(_00981_));
 sg13g2_buf_2 fanout3208 (.A(_00980_),
    .X(net3208));
 sg13g2_buf_1 fanout3209 (.A(_00980_),
    .X(net3209));
 sg13g2_buf_2 fanout3210 (.A(_00980_),
    .X(net3210));
 sg13g2_buf_2 fanout3211 (.A(net3212),
    .X(net3211));
 sg13g2_buf_2 fanout3212 (.A(net3215),
    .X(net3212));
 sg13g2_buf_4 fanout3213 (.X(net3213),
    .A(net3214));
 sg13g2_buf_2 fanout3214 (.A(net3215),
    .X(net3214));
 sg13g2_buf_2 fanout3215 (.A(\core.work.registers.genblk1[1].we ),
    .X(net3215));
 sg13g2_buf_4 fanout3216 (.X(net3216),
    .A(net3217));
 sg13g2_buf_4 fanout3217 (.X(net3217),
    .A(net3220));
 sg13g2_buf_4 fanout3218 (.X(net3218),
    .A(net3220));
 sg13g2_buf_2 fanout3219 (.A(net3220),
    .X(net3219));
 sg13g2_buf_4 fanout3220 (.X(net3220),
    .A(\core.work.registers.genblk1[2].we ));
 sg13g2_buf_4 fanout3221 (.X(net3221),
    .A(net3222));
 sg13g2_buf_4 fanout3222 (.X(net3222),
    .A(net3225));
 sg13g2_buf_4 fanout3223 (.X(net3223),
    .A(net3225));
 sg13g2_buf_4 fanout3224 (.X(net3224),
    .A(net3225));
 sg13g2_buf_4 fanout3225 (.X(net3225),
    .A(\core.work.registers.genblk1[15].we ));
 sg13g2_buf_4 fanout3226 (.X(net3226),
    .A(net3227));
 sg13g2_buf_4 fanout3227 (.X(net3227),
    .A(net3230));
 sg13g2_buf_4 fanout3228 (.X(net3228),
    .A(net3229));
 sg13g2_buf_4 fanout3229 (.X(net3229),
    .A(net3230));
 sg13g2_buf_4 fanout3230 (.X(net3230),
    .A(\core.work.registers.genblk1[3].we ));
 sg13g2_buf_4 fanout3231 (.X(net3231),
    .A(net3232));
 sg13g2_buf_4 fanout3232 (.X(net3232),
    .A(net3235));
 sg13g2_buf_4 fanout3233 (.X(net3233),
    .A(net3235));
 sg13g2_buf_4 fanout3234 (.X(net3234),
    .A(net3235));
 sg13g2_buf_4 fanout3235 (.X(net3235),
    .A(\core.work.registers.genblk1[4].we ));
 sg13g2_buf_4 fanout3236 (.X(net3236),
    .A(net3237));
 sg13g2_buf_4 fanout3237 (.X(net3237),
    .A(net3240));
 sg13g2_buf_4 fanout3238 (.X(net3238),
    .A(net3240));
 sg13g2_buf_4 fanout3239 (.X(net3239),
    .A(net3240));
 sg13g2_buf_4 fanout3240 (.X(net3240),
    .A(\core.work.registers.genblk1[5].we ));
 sg13g2_buf_4 fanout3241 (.X(net3241),
    .A(net3242));
 sg13g2_buf_4 fanout3242 (.X(net3242),
    .A(net3245));
 sg13g2_buf_4 fanout3243 (.X(net3243),
    .A(net3245));
 sg13g2_buf_4 fanout3244 (.X(net3244),
    .A(net3245));
 sg13g2_buf_4 fanout3245 (.X(net3245),
    .A(\core.work.registers.genblk1[6].we ));
 sg13g2_buf_4 fanout3246 (.X(net3246),
    .A(net3247));
 sg13g2_buf_4 fanout3247 (.X(net3247),
    .A(net3250));
 sg13g2_buf_4 fanout3248 (.X(net3248),
    .A(net3250));
 sg13g2_buf_2 fanout3249 (.A(net3250),
    .X(net3249));
 sg13g2_buf_4 fanout3250 (.X(net3250),
    .A(\core.work.registers.genblk1[7].we ));
 sg13g2_buf_4 fanout3251 (.X(net3251),
    .A(net3252));
 sg13g2_buf_4 fanout3252 (.X(net3252),
    .A(net3255));
 sg13g2_buf_4 fanout3253 (.X(net3253),
    .A(net3255));
 sg13g2_buf_4 fanout3254 (.X(net3254),
    .A(net3255));
 sg13g2_buf_4 fanout3255 (.X(net3255),
    .A(\core.work.registers.genblk1[8].we ));
 sg13g2_buf_4 fanout3256 (.X(net3256),
    .A(net3257));
 sg13g2_buf_4 fanout3257 (.X(net3257),
    .A(net3260));
 sg13g2_buf_4 fanout3258 (.X(net3258),
    .A(net3260));
 sg13g2_buf_4 fanout3259 (.X(net3259),
    .A(net3260));
 sg13g2_buf_4 fanout3260 (.X(net3260),
    .A(\core.work.registers.genblk1[9].we ));
 sg13g2_buf_4 fanout3261 (.X(net3261),
    .A(net3262));
 sg13g2_buf_4 fanout3262 (.X(net3262),
    .A(net3265));
 sg13g2_buf_4 fanout3263 (.X(net3263),
    .A(net3265));
 sg13g2_buf_4 fanout3264 (.X(net3264),
    .A(net3265));
 sg13g2_buf_4 fanout3265 (.X(net3265),
    .A(\core.work.registers.genblk1[10].we ));
 sg13g2_buf_4 fanout3266 (.X(net3266),
    .A(net3267));
 sg13g2_buf_4 fanout3267 (.X(net3267),
    .A(net3270));
 sg13g2_buf_4 fanout3268 (.X(net3268),
    .A(net3269));
 sg13g2_buf_4 fanout3269 (.X(net3269),
    .A(net3270));
 sg13g2_buf_4 fanout3270 (.X(net3270),
    .A(\core.work.registers.genblk1[11].we ));
 sg13g2_buf_4 fanout3271 (.X(net3271),
    .A(net3272));
 sg13g2_buf_4 fanout3272 (.X(net3272),
    .A(net3275));
 sg13g2_buf_4 fanout3273 (.X(net3273),
    .A(net3274));
 sg13g2_buf_4 fanout3274 (.X(net3274),
    .A(net3275));
 sg13g2_buf_4 fanout3275 (.X(net3275),
    .A(\core.work.registers.genblk1[12].we ));
 sg13g2_buf_4 fanout3276 (.X(net3276),
    .A(net3277));
 sg13g2_buf_4 fanout3277 (.X(net3277),
    .A(net3280));
 sg13g2_buf_4 fanout3278 (.X(net3278),
    .A(net3280));
 sg13g2_buf_4 fanout3279 (.X(net3279),
    .A(net3280));
 sg13g2_buf_4 fanout3280 (.X(net3280),
    .A(\core.work.registers.genblk1[13].we ));
 sg13g2_buf_4 fanout3281 (.X(net3281),
    .A(net3282));
 sg13g2_buf_4 fanout3282 (.X(net3282),
    .A(net3285));
 sg13g2_buf_4 fanout3283 (.X(net3283),
    .A(net3285));
 sg13g2_buf_4 fanout3284 (.X(net3284),
    .A(net3285));
 sg13g2_buf_4 fanout3285 (.X(net3285),
    .A(\core.work.registers.genblk1[14].we ));
 sg13g2_buf_4 fanout3286 (.X(net3286),
    .A(_05333_));
 sg13g2_buf_4 fanout3287 (.X(net3287),
    .A(net3288));
 sg13g2_buf_4 fanout3288 (.X(net3288),
    .A(_03984_));
 sg13g2_buf_4 fanout3289 (.X(net3289),
    .A(_03972_));
 sg13g2_buf_2 fanout3290 (.A(_03972_),
    .X(net3290));
 sg13g2_buf_4 fanout3291 (.X(net3291),
    .A(net3292));
 sg13g2_buf_4 fanout3292 (.X(net3292),
    .A(_03180_));
 sg13g2_buf_2 fanout3293 (.A(_02764_),
    .X(net3293));
 sg13g2_buf_1 fanout3294 (.A(_02764_),
    .X(net3294));
 sg13g2_buf_2 fanout3295 (.A(_01833_),
    .X(net3295));
 sg13g2_buf_2 fanout3296 (.A(_01812_),
    .X(net3296));
 sg13g2_buf_4 fanout3297 (.X(net3297),
    .A(net3298));
 sg13g2_buf_4 fanout3298 (.X(net3298),
    .A(_01710_));
 sg13g2_buf_2 fanout3299 (.A(net3302),
    .X(net3299));
 sg13g2_buf_1 fanout3300 (.A(net3302),
    .X(net3300));
 sg13g2_buf_4 fanout3301 (.X(net3301),
    .A(net3302));
 sg13g2_buf_4 fanout3302 (.X(net3302),
    .A(_01710_));
 sg13g2_buf_4 fanout3303 (.X(net3303),
    .A(net3307));
 sg13g2_buf_2 fanout3304 (.A(net3307),
    .X(net3304));
 sg13g2_buf_4 fanout3305 (.X(net3305),
    .A(net3307));
 sg13g2_buf_2 fanout3306 (.A(net3307),
    .X(net3306));
 sg13g2_buf_2 fanout3307 (.A(_01709_),
    .X(net3307));
 sg13g2_buf_4 fanout3308 (.X(net3308),
    .A(net3309));
 sg13g2_buf_4 fanout3309 (.X(net3309),
    .A(_01709_));
 sg13g2_buf_4 fanout3310 (.X(net3310),
    .A(net3312));
 sg13g2_buf_4 fanout3311 (.X(net3311),
    .A(net3312));
 sg13g2_buf_2 fanout3312 (.A(net3320),
    .X(net3312));
 sg13g2_buf_4 fanout3313 (.X(net3313),
    .A(net3314));
 sg13g2_buf_4 fanout3314 (.X(net3314),
    .A(net3320));
 sg13g2_buf_4 fanout3315 (.X(net3315),
    .A(net3320));
 sg13g2_buf_2 fanout3316 (.A(net3320),
    .X(net3316));
 sg13g2_buf_4 fanout3317 (.X(net3317),
    .A(net3319));
 sg13g2_buf_2 fanout3318 (.A(net3319),
    .X(net3318));
 sg13g2_buf_2 fanout3319 (.A(net3320),
    .X(net3319));
 sg13g2_buf_4 fanout3320 (.X(net3320),
    .A(_01675_));
 sg13g2_buf_4 fanout3321 (.X(net3321),
    .A(net3324));
 sg13g2_buf_4 fanout3322 (.X(net3322),
    .A(net3323));
 sg13g2_buf_2 fanout3323 (.A(net3324),
    .X(net3323));
 sg13g2_buf_2 fanout3324 (.A(_01656_),
    .X(net3324));
 sg13g2_buf_2 fanout3325 (.A(net3327),
    .X(net3325));
 sg13g2_buf_2 fanout3326 (.A(net3327),
    .X(net3326));
 sg13g2_buf_2 fanout3327 (.A(net3328),
    .X(net3327));
 sg13g2_buf_2 fanout3328 (.A(_01656_),
    .X(net3328));
 sg13g2_buf_2 fanout3329 (.A(net3330),
    .X(net3329));
 sg13g2_buf_4 fanout3330 (.X(net3330),
    .A(_01646_));
 sg13g2_buf_4 fanout3331 (.X(net3331),
    .A(net3332));
 sg13g2_buf_2 fanout3332 (.A(_01645_),
    .X(net3332));
 sg13g2_buf_2 fanout3333 (.A(_01385_),
    .X(net3333));
 sg13g2_buf_2 fanout3334 (.A(_01385_),
    .X(net3334));
 sg13g2_buf_2 fanout3335 (.A(net3339),
    .X(net3335));
 sg13g2_buf_4 fanout3336 (.X(net3336),
    .A(net3338));
 sg13g2_buf_2 fanout3337 (.A(net3338),
    .X(net3337));
 sg13g2_buf_2 fanout3338 (.A(net3339),
    .X(net3338));
 sg13g2_buf_2 fanout3339 (.A(_01325_),
    .X(net3339));
 sg13g2_buf_2 fanout3340 (.A(net3342),
    .X(net3340));
 sg13g2_buf_1 fanout3341 (.A(net3342),
    .X(net3341));
 sg13g2_buf_2 fanout3342 (.A(net3343),
    .X(net3342));
 sg13g2_buf_2 fanout3343 (.A(net3344),
    .X(net3343));
 sg13g2_buf_2 fanout3344 (.A(net3349),
    .X(net3344));
 sg13g2_buf_2 fanout3345 (.A(net3347),
    .X(net3345));
 sg13g2_buf_2 fanout3346 (.A(net3347),
    .X(net3346));
 sg13g2_buf_2 fanout3347 (.A(net3348),
    .X(net3347));
 sg13g2_buf_2 fanout3348 (.A(net3349),
    .X(net3348));
 sg13g2_buf_4 fanout3349 (.X(net3349),
    .A(_01324_));
 sg13g2_buf_4 fanout3350 (.X(net3350),
    .A(net3351));
 sg13g2_buf_4 fanout3351 (.X(net3351),
    .A(_01132_));
 sg13g2_buf_2 fanout3352 (.A(net3354),
    .X(net3352));
 sg13g2_buf_1 fanout3353 (.A(net3354),
    .X(net3353));
 sg13g2_buf_4 fanout3354 (.X(net3354),
    .A(_00766_));
 sg13g2_buf_2 fanout3355 (.A(net3358),
    .X(net3355));
 sg13g2_buf_2 fanout3356 (.A(net3358),
    .X(net3356));
 sg13g2_buf_1 fanout3357 (.A(net3358),
    .X(net3357));
 sg13g2_buf_2 fanout3358 (.A(_00765_),
    .X(net3358));
 sg13g2_buf_4 fanout3359 (.X(net3359),
    .A(net3360));
 sg13g2_buf_2 fanout3360 (.A(net3361),
    .X(net3360));
 sg13g2_buf_4 fanout3361 (.X(net3361),
    .A(_00636_));
 sg13g2_buf_2 fanout3362 (.A(_00631_),
    .X(net3362));
 sg13g2_buf_2 fanout3363 (.A(net3365),
    .X(net3363));
 sg13g2_buf_1 fanout3364 (.A(net3365),
    .X(net3364));
 sg13g2_buf_1 fanout3365 (.A(net771),
    .X(net3365));
 sg13g2_buf_2 fanout3366 (.A(net3367),
    .X(net3366));
 sg13g2_buf_1 fanout3367 (.A(net3368),
    .X(net3367));
 sg13g2_buf_2 fanout3368 (.A(net783),
    .X(net3368));
 sg13g2_buf_2 fanout3369 (.A(net3370),
    .X(net3369));
 sg13g2_buf_1 fanout3370 (.A(net3371),
    .X(net3370));
 sg13g2_buf_1 fanout3371 (.A(\core.work.registers.tmp[29] ),
    .X(net3371));
 sg13g2_buf_2 fanout3372 (.A(net3373),
    .X(net3372));
 sg13g2_buf_1 fanout3373 (.A(net3374),
    .X(net3373));
 sg13g2_buf_1 fanout3374 (.A(\core.work.registers.tmp[28] ),
    .X(net3374));
 sg13g2_buf_2 fanout3375 (.A(net3376),
    .X(net3375));
 sg13g2_buf_2 fanout3376 (.A(\core.work.registers.tmp[27] ),
    .X(net3376));
 sg13g2_buf_2 fanout3377 (.A(net3378),
    .X(net3377));
 sg13g2_buf_2 fanout3378 (.A(\core.work.registers.tmp[26] ),
    .X(net3378));
 sg13g2_buf_2 fanout3379 (.A(net3381),
    .X(net3379));
 sg13g2_buf_1 fanout3380 (.A(net3381),
    .X(net3380));
 sg13g2_buf_1 fanout3381 (.A(net775),
    .X(net3381));
 sg13g2_buf_2 fanout3382 (.A(net3384),
    .X(net3382));
 sg13g2_buf_1 fanout3383 (.A(net3384),
    .X(net3383));
 sg13g2_buf_2 fanout3384 (.A(net770),
    .X(net3384));
 sg13g2_buf_2 fanout3385 (.A(net3386),
    .X(net3385));
 sg13g2_buf_1 fanout3386 (.A(net3387),
    .X(net3386));
 sg13g2_buf_2 fanout3387 (.A(\core.work.registers.tmp[23] ),
    .X(net3387));
 sg13g2_buf_2 fanout3388 (.A(net3389),
    .X(net3388));
 sg13g2_buf_2 fanout3389 (.A(\core.work.registers.tmp[22] ),
    .X(net3389));
 sg13g2_buf_2 fanout3390 (.A(net3392),
    .X(net3390));
 sg13g2_buf_1 fanout3391 (.A(net3392),
    .X(net3391));
 sg13g2_buf_2 fanout3392 (.A(net800),
    .X(net3392));
 sg13g2_buf_2 fanout3393 (.A(net3394),
    .X(net3393));
 sg13g2_buf_2 fanout3394 (.A(net830),
    .X(net3394));
 sg13g2_buf_2 fanout3395 (.A(net3396),
    .X(net3395));
 sg13g2_buf_1 fanout3396 (.A(net3397),
    .X(net3396));
 sg13g2_buf_2 fanout3397 (.A(\core.work.registers.tmp[19] ),
    .X(net3397));
 sg13g2_buf_2 fanout3398 (.A(net3399),
    .X(net3398));
 sg13g2_buf_2 fanout3399 (.A(\core.work.registers.tmp[18] ),
    .X(net3399));
 sg13g2_buf_2 fanout3400 (.A(net3401),
    .X(net3400));
 sg13g2_buf_2 fanout3401 (.A(\core.work.registers.tmp[17] ),
    .X(net3401));
 sg13g2_buf_2 fanout3402 (.A(net3404),
    .X(net3402));
 sg13g2_buf_1 fanout3403 (.A(net3404),
    .X(net3403));
 sg13g2_buf_2 fanout3404 (.A(net751),
    .X(net3404));
 sg13g2_buf_2 fanout3405 (.A(net3407),
    .X(net3405));
 sg13g2_buf_2 fanout3406 (.A(net3407),
    .X(net3406));
 sg13g2_buf_2 fanout3407 (.A(net761),
    .X(net3407));
 sg13g2_buf_2 fanout3408 (.A(net3409),
    .X(net3408));
 sg13g2_buf_2 fanout3409 (.A(net818),
    .X(net3409));
 sg13g2_buf_2 fanout3410 (.A(net3411),
    .X(net3410));
 sg13g2_buf_2 fanout3411 (.A(\core.work.registers.tmp[13] ),
    .X(net3411));
 sg13g2_buf_2 fanout3412 (.A(net3413),
    .X(net3412));
 sg13g2_buf_2 fanout3413 (.A(\core.work.registers.tmp[12] ),
    .X(net3413));
 sg13g2_buf_2 fanout3414 (.A(net3416),
    .X(net3414));
 sg13g2_buf_1 fanout3415 (.A(net3416),
    .X(net3415));
 sg13g2_buf_1 fanout3416 (.A(net769),
    .X(net3416));
 sg13g2_buf_2 fanout3417 (.A(net3418),
    .X(net3417));
 sg13g2_buf_2 fanout3418 (.A(net624),
    .X(net3418));
 sg13g2_buf_2 fanout3419 (.A(net821),
    .X(net3419));
 sg13g2_buf_2 fanout3420 (.A(\core.work.registers.tmp[9] ),
    .X(net3420));
 sg13g2_buf_2 fanout3421 (.A(net3422),
    .X(net3421));
 sg13g2_buf_2 fanout3422 (.A(net851),
    .X(net3422));
 sg13g2_buf_2 fanout3423 (.A(net3424),
    .X(net3423));
 sg13g2_buf_2 fanout3424 (.A(\core.work.registers.tmp[7] ),
    .X(net3424));
 sg13g2_buf_2 fanout3425 (.A(net3426),
    .X(net3425));
 sg13g2_buf_2 fanout3426 (.A(\core.work.registers.tmp[6] ),
    .X(net3426));
 sg13g2_buf_2 fanout3427 (.A(net3428),
    .X(net3427));
 sg13g2_buf_2 fanout3428 (.A(\core.work.registers.tmp[5] ),
    .X(net3428));
 sg13g2_buf_2 fanout3429 (.A(net3431),
    .X(net3429));
 sg13g2_buf_1 fanout3430 (.A(net3431),
    .X(net3430));
 sg13g2_buf_2 fanout3431 (.A(net764),
    .X(net3431));
 sg13g2_buf_2 fanout3432 (.A(net3433),
    .X(net3432));
 sg13g2_buf_2 fanout3433 (.A(\core.work.registers.tmp[3] ),
    .X(net3433));
 sg13g2_buf_2 fanout3434 (.A(net3435),
    .X(net3434));
 sg13g2_buf_2 fanout3435 (.A(net837),
    .X(net3435));
 sg13g2_buf_2 fanout3436 (.A(net3437),
    .X(net3436));
 sg13g2_buf_2 fanout3437 (.A(\core.work.registers.tmp[1] ),
    .X(net3437));
 sg13g2_buf_2 fanout3438 (.A(\core.work.registers.tmp[0] ),
    .X(net3438));
 sg13g2_buf_1 fanout3439 (.A(\core.work.registers.tmp[0] ),
    .X(net3439));
 sg13g2_buf_4 fanout3440 (.X(net3440),
    .A(net883));
 sg13g2_buf_4 fanout3441 (.X(net3441),
    .A(net438));
 sg13g2_buf_4 fanout3442 (.X(net3442),
    .A(_00024_));
 sg13g2_buf_4 fanout3443 (.X(net3443),
    .A(\core.e2m_addr[31] ));
 sg13g2_buf_4 fanout3444 (.X(net3444),
    .A(\core.e2m_addr[30] ));
 sg13g2_buf_4 fanout3445 (.X(net3445),
    .A(net3446));
 sg13g2_buf_4 fanout3446 (.X(net3446),
    .A(\core.e2m_addr[29] ));
 sg13g2_buf_4 fanout3447 (.X(net3447),
    .A(\core.e2m_addr[28] ));
 sg13g2_buf_4 fanout3448 (.X(net3448),
    .A(net885));
 sg13g2_buf_4 fanout3449 (.X(net3449),
    .A(net873));
 sg13g2_buf_4 fanout3450 (.X(net3450),
    .A(\core.e2m_addr[25] ));
 sg13g2_buf_4 fanout3451 (.X(net3451),
    .A(net863));
 sg13g2_buf_4 fanout3452 (.X(net3452),
    .A(_00038_));
 sg13g2_buf_2 fanout3453 (.A(net3454),
    .X(net3453));
 sg13g2_buf_4 fanout3454 (.X(net3454),
    .A(net828));
 sg13g2_buf_2 fanout3455 (.A(net3456),
    .X(net3455));
 sg13g2_buf_4 fanout3456 (.X(net3456),
    .A(net815));
 sg13g2_buf_2 fanout3457 (.A(net3458),
    .X(net3457));
 sg13g2_buf_2 fanout3458 (.A(net3459),
    .X(net3458));
 sg13g2_buf_2 fanout3459 (.A(\core.e2m_addr[21] ),
    .X(net3459));
 sg13g2_buf_4 fanout3460 (.X(net3460),
    .A(_00032_));
 sg13g2_buf_2 fanout3461 (.A(net3463),
    .X(net3461));
 sg13g2_buf_4 fanout3462 (.X(net3462),
    .A(net3463));
 sg13g2_buf_2 fanout3463 (.A(\core.e2m_addr[20] ),
    .X(net3463));
 sg13g2_buf_4 fanout3464 (.X(net3464),
    .A(net3466));
 sg13g2_buf_4 fanout3465 (.X(net3465),
    .A(net3466));
 sg13g2_buf_2 fanout3466 (.A(net3467),
    .X(net3466));
 sg13g2_buf_2 fanout3467 (.A(\core.e2m_addr[20] ),
    .X(net3467));
 sg13g2_buf_4 fanout3468 (.X(net3468),
    .A(\core.e2m_addr[18] ));
 sg13g2_buf_4 fanout3469 (.X(net3469),
    .A(net3470));
 sg13g2_buf_4 fanout3470 (.X(net3470),
    .A(net864));
 sg13g2_buf_4 fanout3471 (.X(net3471),
    .A(net3472));
 sg13g2_buf_4 fanout3472 (.X(net3472),
    .A(net793));
 sg13g2_buf_2 fanout3473 (.A(net3475),
    .X(net3473));
 sg13g2_buf_4 fanout3474 (.X(net3474),
    .A(net3475));
 sg13g2_buf_4 fanout3475 (.X(net3475),
    .A(\core.e2m_addr[15] ));
 sg13g2_buf_2 fanout3476 (.A(net3477),
    .X(net3476));
 sg13g2_buf_2 fanout3477 (.A(net3478),
    .X(net3477));
 sg13g2_buf_4 fanout3478 (.X(net3478),
    .A(net3479));
 sg13g2_buf_2 fanout3479 (.A(\core.e2m_addr[15] ),
    .X(net3479));
 sg13g2_buf_4 fanout3480 (.X(net3480),
    .A(net3481));
 sg13g2_buf_4 fanout3481 (.X(net3481),
    .A(\core.e2m_addr[14] ));
 sg13g2_buf_2 fanout3482 (.A(net3483),
    .X(net3482));
 sg13g2_buf_4 fanout3483 (.X(net3483),
    .A(\core.e2m_addr[13] ));
 sg13g2_buf_4 fanout3484 (.X(net3484),
    .A(\core.e2m_addr[12] ));
 sg13g2_buf_1 fanout3485 (.A(\core.e2m_addr[12] ),
    .X(net3485));
 sg13g2_buf_4 fanout3486 (.X(net3486),
    .A(net385));
 sg13g2_buf_2 fanout3487 (.A(net385),
    .X(net3487));
 sg13g2_buf_4 fanout3488 (.X(net3488),
    .A(net573));
 sg13g2_buf_2 fanout3489 (.A(net3491),
    .X(net3489));
 sg13g2_buf_2 fanout3490 (.A(net3491),
    .X(net3490));
 sg13g2_buf_2 fanout3491 (.A(net3492),
    .X(net3491));
 sg13g2_buf_4 fanout3492 (.X(net3492),
    .A(\core.e2m_addr[5] ));
 sg13g2_buf_4 fanout3493 (.X(net3493),
    .A(net3494));
 sg13g2_buf_4 fanout3494 (.X(net3494),
    .A(\core.e2m_addr[5] ));
 sg13g2_buf_4 fanout3495 (.X(net3495),
    .A(net704));
 sg13g2_buf_4 fanout3496 (.X(net3496),
    .A(net869));
 sg13g2_buf_4 fanout3497 (.X(net3497),
    .A(net774));
 sg13g2_buf_2 fanout3498 (.A(net774),
    .X(net3498));
 sg13g2_buf_4 fanout3499 (.X(net3499),
    .A(net744));
 sg13g2_buf_4 fanout3500 (.X(net3500),
    .A(net900));
 sg13g2_buf_4 fanout3501 (.X(net3501),
    .A(net887));
 sg13g2_buf_4 fanout3502 (.X(net3502),
    .A(\core.work.state[0] ));
 sg13g2_buf_4 fanout3503 (.X(net3503),
    .A(net886));
 sg13g2_buf_2 fanout3504 (.A(net3505),
    .X(net3504));
 sg13g2_buf_2 fanout3505 (.A(net756),
    .X(net3505));
 sg13g2_buf_2 fanout3506 (.A(_00149_),
    .X(net3506));
 sg13g2_buf_4 fanout3507 (.X(net3507),
    .A(net825));
 sg13g2_buf_2 fanout3508 (.A(net3509),
    .X(net3508));
 sg13g2_buf_2 fanout3509 (.A(net813),
    .X(net3509));
 sg13g2_buf_4 fanout3510 (.X(net3510),
    .A(net804));
 sg13g2_buf_4 fanout3511 (.X(net3511),
    .A(net822));
 sg13g2_buf_4 fanout3512 (.X(net3512),
    .A(net844));
 sg13g2_buf_4 fanout3513 (.X(net3513),
    .A(net857));
 sg13g2_buf_4 fanout3514 (.X(net3514),
    .A(_00057_));
 sg13g2_buf_4 fanout3515 (.X(net3515),
    .A(net3516));
 sg13g2_buf_2 fanout3516 (.A(\core.lsu.write_index[1] ),
    .X(net3516));
 sg13g2_buf_4 fanout3517 (.X(net3517),
    .A(net3519));
 sg13g2_buf_1 fanout3518 (.A(net3519),
    .X(net3518));
 sg13g2_buf_4 fanout3519 (.X(net3519),
    .A(\core.lsu.write_index[0] ));
 sg13g2_buf_2 fanout3520 (.A(net866),
    .X(net3520));
 sg13g2_buf_4 fanout3521 (.X(net3521),
    .A(net3522));
 sg13g2_buf_2 fanout3522 (.A(\core.lsu.spi.sck ),
    .X(net3522));
 sg13g2_buf_2 fanout3523 (.A(net843),
    .X(net3523));
 sg13g2_buf_4 fanout3524 (.X(net3524),
    .A(\core.lsu.is_byte ));
 sg13g2_buf_2 fanout3525 (.A(net788),
    .X(net3525));
 sg13g2_buf_4 fanout3526 (.X(net3526),
    .A(\core.fetch.rd_addr_i[1] ));
 sg13g2_buf_2 fanout3527 (.A(\core.fetch.inst_size[2] ),
    .X(net3527));
 sg13g2_buf_4 fanout3528 (.X(net3528),
    .A(net898));
 sg13g2_buf_2 fanout3529 (.A(\core.fetch.inst_size[0] ),
    .X(net3529));
 sg13g2_buf_4 fanout3530 (.X(net3530),
    .A(\core.work.alu.sval2[20] ));
 sg13g2_buf_2 fanout3531 (.A(\core.work.alu.sval2[19] ),
    .X(net3531));
 sg13g2_buf_2 fanout3532 (.A(\core.work.alu.sval2[17] ),
    .X(net3532));
 sg13g2_buf_2 fanout3533 (.A(net853),
    .X(net3533));
 sg13g2_buf_2 fanout3534 (.A(\core.work.alu.sval2[23] ),
    .X(net3534));
 sg13g2_buf_4 fanout3535 (.X(net3535),
    .A(net784));
 sg13g2_buf_2 fanout3536 (.A(net838),
    .X(net3536));
 sg13g2_buf_2 fanout3537 (.A(\core.work.alu.sval2[27] ),
    .X(net3537));
 sg13g2_buf_4 fanout3538 (.X(net3538),
    .A(net3539));
 sg13g2_buf_4 fanout3539 (.X(net3539),
    .A(\core.work.alu.sval2[0] ));
 sg13g2_buf_2 fanout3540 (.A(net848),
    .X(net3540));
 sg13g2_buf_4 fanout3541 (.X(net3541),
    .A(net826));
 sg13g2_buf_2 fanout3542 (.A(net875),
    .X(net3542));
 sg13g2_buf_2 fanout3543 (.A(net846),
    .X(net3543));
 sg13g2_buf_4 fanout3544 (.X(net3544),
    .A(_00054_));
 sg13g2_buf_2 fanout3545 (.A(net3546),
    .X(net3545));
 sg13g2_buf_2 fanout3546 (.A(_00054_),
    .X(net3546));
 sg13g2_buf_2 fanout3547 (.A(net3550),
    .X(net3547));
 sg13g2_buf_4 fanout3548 (.X(net3548),
    .A(net3550));
 sg13g2_buf_2 fanout3549 (.A(net3550),
    .X(net3549));
 sg13g2_buf_2 fanout3550 (.A(\core.work.alu.sval2[4] ),
    .X(net3550));
 sg13g2_buf_4 fanout3551 (.X(net3551),
    .A(_00109_));
 sg13g2_buf_4 fanout3552 (.X(net3552),
    .A(net3554));
 sg13g2_buf_2 fanout3553 (.A(net3554),
    .X(net3553));
 sg13g2_buf_4 fanout3554 (.X(net3554),
    .A(net757));
 sg13g2_buf_4 fanout3555 (.X(net3555),
    .A(net3556));
 sg13g2_buf_2 fanout3556 (.A(_00142_),
    .X(net3556));
 sg13g2_buf_2 fanout3557 (.A(net3558),
    .X(net3557));
 sg13g2_buf_2 fanout3558 (.A(net3559),
    .X(net3558));
 sg13g2_buf_4 fanout3559 (.X(net3559),
    .A(\core.work.alu.sval2[2] ));
 sg13g2_buf_4 fanout3560 (.X(net3560),
    .A(\core.work.alu.sval2[1] ));
 sg13g2_buf_2 fanout3561 (.A(net831),
    .X(net3561));
 sg13g2_buf_4 fanout3562 (.X(net3562),
    .A(\core.work.alu.sval2[1] ));
 sg13g2_buf_2 fanout3563 (.A(net874),
    .X(net3563));
 sg13g2_buf_2 fanout3564 (.A(\core.f2e_addr[4] ),
    .X(net3564));
 sg13g2_buf_4 fanout3565 (.X(net3565),
    .A(\core.fetch.cmd_valid ));
 sg13g2_buf_2 fanout3566 (.A(net862),
    .X(net3566));
 sg13g2_buf_2 fanout3567 (.A(\core.fetch.spi_reader.state[1] ),
    .X(net3567));
 sg13g2_buf_4 fanout3568 (.X(net3568),
    .A(net795));
 sg13g2_buf_4 fanout3569 (.X(net3569),
    .A(net587));
 sg13g2_buf_4 fanout3570 (.X(net3570),
    .A(net418));
 sg13g2_buf_4 fanout3571 (.X(net3571),
    .A(net3573));
 sg13g2_buf_2 fanout3572 (.A(net3573),
    .X(net3572));
 sg13g2_buf_2 fanout3573 (.A(\core.fetch.spi_reader.sck ),
    .X(net3573));
 sg13g2_buf_2 fanout3574 (.A(net3575),
    .X(net3574));
 sg13g2_buf_2 fanout3575 (.A(\core.fetch.spi_reader.cs ),
    .X(net3575));
 sg13g2_buf_2 fanout3576 (.A(net799),
    .X(net3576));
 sg13g2_buf_2 fanout3577 (.A(net789),
    .X(net3577));
 sg13g2_buf_2 fanout3578 (.A(net847),
    .X(net3578));
 sg13g2_buf_4 fanout3579 (.X(net3579),
    .A(net3580));
 sg13g2_buf_4 fanout3580 (.X(net3580),
    .A(net3581));
 sg13g2_buf_2 fanout3581 (.A(net3582),
    .X(net3581));
 sg13g2_buf_4 fanout3582 (.X(net3582),
    .A(net3596));
 sg13g2_buf_4 fanout3583 (.X(net3583),
    .A(net3584));
 sg13g2_buf_4 fanout3584 (.X(net3584),
    .A(net3596));
 sg13g2_buf_4 fanout3585 (.X(net3585),
    .A(net3586));
 sg13g2_buf_4 fanout3586 (.X(net3586),
    .A(net3587));
 sg13g2_buf_4 fanout3587 (.X(net3587),
    .A(net3596));
 sg13g2_buf_4 fanout3588 (.X(net3588),
    .A(net3589));
 sg13g2_buf_4 fanout3589 (.X(net3589),
    .A(net3590));
 sg13g2_buf_4 fanout3590 (.X(net3590),
    .A(net3594));
 sg13g2_buf_4 fanout3591 (.X(net3591),
    .A(net3594));
 sg13g2_buf_4 fanout3592 (.X(net3592),
    .A(net3593));
 sg13g2_buf_4 fanout3593 (.X(net3593),
    .A(net3594));
 sg13g2_buf_2 fanout3594 (.A(net3595),
    .X(net3594));
 sg13g2_buf_4 fanout3595 (.X(net3595),
    .A(net3596));
 sg13g2_buf_4 fanout3596 (.X(net3596),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[2]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[6]),
    .X(net10));
 sg13g2_tielo tt_um_dumbrv_yliu_hashed_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_3__leaf_clk));
 sg13g2_buf_2 clkbuf_leaf_0_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_1_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_2_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_3_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_4_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_5_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_6_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_7_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_8_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_9_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_10_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_11_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_12_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_13_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_14_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_15_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_16_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_17_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_18_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_19_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_20_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_21_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_22_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_23_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_23_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_24_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_25_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_26_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_27_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_28_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_29_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_29_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_30_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_30_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_31_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_31_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_32_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_32_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_33_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_33_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_34_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_34_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_35_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_35_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_36_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_36_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_37_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_37_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_38_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_38_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_39_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_39_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_40_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_40_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_41_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_41_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_42_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_42_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_43_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_43_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_45_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_45_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_46_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_46_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_47_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_47_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_48_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_48_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_49_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_49_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_50_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_50_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_51_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_51_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_52_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_52_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_53_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_53_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_54_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_54_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_55_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_55_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_56_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_56_clk_regs));
 sg13g2_buf_2 clkbuf_leaf_57_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_57_clk_regs));
 sg13g2_buf_2 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_2 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_2 clkload1 (.A(clknet_4_3_0_clk_regs));
 sg13g2_buf_2 clkload2 (.A(clknet_4_5_0_clk_regs));
 sg13g2_buf_2 clkload3 (.A(clknet_4_7_0_clk_regs));
 sg13g2_buf_1 clkload4 (.A(clknet_4_11_0_clk_regs));
 sg13g2_buf_2 clkload5 (.A(clknet_4_13_0_clk_regs));
 sg13g2_buf_2 clkload6 (.A(clknet_4_15_0_clk_regs));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_1_clk_regs));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_56_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_57_clk_regs));
 sg13g2_inv_8 clkload10 (.A(clknet_leaf_5_clk_regs));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_53_clk_regs));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_55_clk_regs));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_12_clk_regs));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_17_clk_regs));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_19_clk_regs));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_21_clk_regs));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_7_clk_regs));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_50_clk_regs));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_8_clk_regs));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_45_clk_regs));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_46_clk_regs));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_48_clk_regs));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_42_clk_regs));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_34_clk_regs));
 sg13g2_inv_4 clkload25 (.A(clknet_leaf_40_clk_regs));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_41_clk_regs));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_36_clk_regs));
 sg13g2_inv_1 clkload28 (.A(clknet_leaf_37_clk_regs));
 sg13g2_buf_2 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(delaynet_1_clk));
 sg13g2_buf_2 delaybuf_1_clk (.A(delaynet_1_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_00105_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold2 (.A(_01383_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold3 (.A(_00220_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold4 (.A(_00128_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold5 (.A(_02761_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold6 (.A(_00380_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold7 (.A(\core.lsu.spi.counter[5] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold8 (.A(_00418_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold9 (.A(\core.fetch.inst_size[0] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold10 (.A(_00163_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold11 (.A(_00307_),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold12 (.A(\core.fetch.data[28] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold13 (.A(_00213_),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold14 (.A(\core.fetch.rd_addr_i[7] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold15 (.A(\core.fetch.data[25] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold16 (.A(_00210_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold17 (.A(\core.lsu.spi.addr[15] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold18 (.A(_00406_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold19 (.A(\core.e2m_data[1] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold20 (.A(\core.fetch.rd_addr_i[15] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold21 (.A(\core.fetch.spi_reader.counter[4] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold22 (.A(_00310_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold23 (.A(\core.fetch.rd_addr_i[14] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold24 (.A(\core.lsu.spi.counter[2] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold25 (.A(_00415_),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold26 (.A(\core.fetch.rd_addr_i[6] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold27 (.A(_00318_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold28 (.A(\core.fetch.data[27] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold29 (.A(_00212_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold30 (.A(\core.e2m_addr[10] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold31 (.A(_00322_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold32 (.A(\core.fetch.spi_reader.cache_bit ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold33 (.A(\core.fetch.data[29] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold34 (.A(_00214_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold35 (.A(\core.fetch.data[14] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold36 (.A(_00199_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold37 (.A(\core.work.dreg[2] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold38 (.A(_00378_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold39 (.A(\core.work.registers.tmp[7] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold40 (.A(\core.fetch.rd_addr_i[1] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold41 (.A(_00313_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold42 (.A(\core.fetch.data[13] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold43 (.A(_00198_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold44 (.A(\core.lsu.is_signed ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold45 (.A(_00340_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold46 (.A(\core.fetch.data[5] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold47 (.A(_00190_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold48 (.A(\core.work.registers.tmp[23] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold49 (.A(\core.fetch.data[26] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold50 (.A(_00211_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold51 (.A(_00127_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold52 (.A(_03000_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold53 (.A(_00414_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold54 (.A(\core.work.registers.tmp[19] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold55 (.A(_00566_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold56 (.A(_00103_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold57 (.A(_00208_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold58 (.A(\core.e2m_data[24] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold59 (.A(\core.work.dreg[3] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold60 (.A(_00379_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold61 (.A(\core.fetch.data[31] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold62 (.A(_00216_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold63 (.A(\core.fetch.cmd_data[0] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold64 (.A(\core.f2e_inst[21] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold65 (.A(_00440_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold66 (.A(_00101_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold67 (.A(_00206_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold68 (.A(\core.fetch.data[30] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold69 (.A(_00215_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold70 (.A(\core.fetch.spi_reader.counter[5] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold71 (.A(_00311_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold72 (.A(\core.f2e_addr[4] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold73 (.A(_00253_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold74 (.A(_00102_),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold75 (.A(_00207_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold76 (.A(_00164_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold77 (.A(_00308_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold78 (.A(\core.fetch.spi_reader.counter[3] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold79 (.A(_00309_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold80 (.A(\core.lsu.spi.cache_bit ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold81 (.A(\core.fetch.spi_reader.dirty ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold82 (.A(_00250_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold83 (.A(\core.work.alu.ls_size_h ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold84 (.A(_00341_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold85 (.A(\core.work.registers.tmp[22] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold86 (.A(_00569_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold87 (.A(\core.fetch.data[6] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold88 (.A(_00191_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold89 (.A(\core.e2m_data[16] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold90 (.A(\core.lsu.spi.counter[4] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold91 (.A(_00417_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold92 (.A(\core.fetch.rd_addr_i[5] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold93 (.A(\core.f2e_inst[31] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold94 (.A(_00450_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold95 (.A(\core.f2e_inst[18] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold96 (.A(_00437_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold97 (.A(_00099_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold98 (.A(_00204_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold99 (.A(\core.e2m_data[7] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold100 (.A(\core.fetch.data[7] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold101 (.A(_00192_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold102 (.A(\core.e2m_data[3] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold103 (.A(\core.work.inst_was_short ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold104 (.A(\core.work.alu.sval2[20] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold105 (.A(_00297_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold106 (.A(\core.lsu.spi.dirty ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold107 (.A(_00382_),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold108 (.A(\core.e2m_data[4] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold109 (.A(\core.fetch.data[24] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold110 (.A(\core.fetch.data[3] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold111 (.A(_00188_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold112 (.A(\core.e2m_data[19] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold113 (.A(\core.e2m_data[0] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold114 (.A(\core.fetch.spi_reader.addr[14] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold115 (.A(\core.fetch.spi_reader.state[1] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold116 (.A(_00247_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold117 (.A(\core.fetch.inst[32] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold118 (.A(_03117_),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold119 (.A(_00435_),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold120 (.A(\core.e2m_data[18] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold121 (.A(\core.e2m_data[25] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold122 (.A(_00096_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold123 (.A(_00201_),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold124 (.A(\core.fetch.data[9] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold125 (.A(_00194_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold126 (.A(\core.lsu.spi.addr[0] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold127 (.A(_00391_),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold128 (.A(\core.e2m_data[22] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold129 (.A(\core.lsu.spi.counter[3] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold130 (.A(_00416_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold131 (.A(\core.f2e_inst[30] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold132 (.A(_00449_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold133 (.A(\core.e2m_data[20] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold134 (.A(\core.e2m_data[17] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold135 (.A(\core.fetch.data[8] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold136 (.A(\core.e2m_data[21] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold137 (.A(\core.fetch.data[0] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold138 (.A(\core.e2m_data[26] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold139 (.A(\core.fetch.spi_reader.addr[3] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold140 (.A(_00233_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold141 (.A(\core.fetch.spi_reader.addr[0] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold142 (.A(_00230_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold143 (.A(\core.f2e_inst[28] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold144 (.A(_00447_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold145 (.A(_00100_),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold146 (.A(_00205_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold147 (.A(\core.lsu.spi.iswr ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold148 (.A(_00452_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold149 (.A(\core.fetch.data[10] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold150 (.A(_00195_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold151 (.A(\core.fetch.inst[33] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold152 (.A(_03121_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold153 (.A(_00436_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold154 (.A(\core.lsu.spi.addr[4] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold155 (.A(_00395_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold156 (.A(\core.work.registers.tmp[13] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold157 (.A(\core.e2m_data[29] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold158 (.A(\core.work.op[4] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold159 (.A(\core.work.registers.tmp[0] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold160 (.A(_00097_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold161 (.A(_00202_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold162 (.A(\core.e2m_data[6] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold163 (.A(\core.f2e_inst[26] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold164 (.A(_00445_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold165 (.A(\core.fetch.inst[36] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold166 (.A(\core.e2m_data[12] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold167 (.A(\core.fetch.data[15] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold168 (.A(_00200_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold169 (.A(\core.fetch.inst[41] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold170 (.A(\core.work.registers.tmp[6] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold171 (.A(\core.work.registers.wr_reg[0] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold172 (.A(_00299_),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold173 (.A(\core.fetch.inst[40] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold174 (.A(\core.e2m_data[27] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold175 (.A(\core.fetch.inst[45] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold176 (.A(\core.fetch.inst[35] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold177 (.A(_03127_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold178 (.A(_00438_),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold179 (.A(\core.fetch.inst[47] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold180 (.A(_00543_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold181 (.A(\core.fetch.inst[38] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold182 (.A(_03140_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold183 (.A(_00441_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold184 (.A(\core.fetch.inst[39] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold185 (.A(_00442_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold186 (.A(\core.work.dreg[0] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold187 (.A(\core.e2m_data[10] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold188 (.A(\core.f2e_inst[20] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold189 (.A(\core.work.registers.state[2] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold190 (.A(\core.f2e_inst[29] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold191 (.A(\core.e2m_data[5] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold192 (.A(\core.fetch.spi_reader.addr[15] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold193 (.A(_00245_),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold194 (.A(\core.lsu.spi.addr[14] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold195 (.A(\core.lsu.spi.addr[6] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold196 (.A(\core.lsu.spi.addr[2] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold197 (.A(_00393_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold198 (.A(\core.fetch.inst[42] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold199 (.A(_00538_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold200 (.A(\core.f2e_inst[24] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold201 (.A(\core.lsu.spi.addr[5] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold202 (.A(_00396_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold203 (.A(\core.lsu.spi.addr[8] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold204 (.A(\core.lsu.dreg[0] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold205 (.A(\core.e2m_data[8] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold206 (.A(\core.lsu.spi.addr[12] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold207 (.A(\core.work.dreg[1] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold208 (.A(\core.fetch.inst[44] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold209 (.A(\core.fetch.inst[43] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold210 (.A(\core.fetch.cmd_data[6] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold211 (.A(_05270_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold212 (.A(uo_out[1]),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold213 (.A(\core.work.registers.wr_reg[1] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold214 (.A(\core.fetch.data[2] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold215 (.A(_00187_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold216 (.A(\core.fetch.cmd_data[3] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold217 (.A(\core.lsu.dreg[1] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold218 (.A(\core.e2m_addr[9] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold219 (.A(\core.fetch.inst[46] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold220 (.A(_00542_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold221 (.A(\core.work.registers.tmp[5] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold222 (.A(_00552_),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold223 (.A(\core.lsu.spi.addr[9] ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold224 (.A(\core.lsu.spi_valid ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold225 (.A(_00342_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold226 (.A(\core.fetch.inst[37] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold227 (.A(\core.f2e_inst[8] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold228 (.A(\core.work.registers.tmp[12] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold229 (.A(\core.e2m_data[23] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold230 (.A(\core.fetch.inst[34] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold231 (.A(_00530_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold232 (.A(\core.fetch.cmd_data[1] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold233 (.A(\core.fetch.spi_reader.addr[4] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold234 (.A(uo_out[7]),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold235 (.A(\core.lsu.state[2] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold236 (.A(_00338_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold237 (.A(\core.e2m_data[30] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold238 (.A(\core.fetch.data[4] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold239 (.A(_00189_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold240 (.A(\core.work.registers.tmp[27] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold241 (.A(\core.fetch.spi_reader.addr[12] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold242 (.A(\core.e2m_data[13] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold243 (.A(_00262_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold244 (.A(\core.work.registers.tmp[17] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold245 (.A(_00564_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold246 (.A(_00098_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold247 (.A(_00203_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold248 (.A(\core.f2e_inst[27] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold249 (.A(\core.e2m_data[13] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold250 (.A(\core.f2e_inst[25] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold251 (.A(_00444_),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold252 (.A(\core.fetch.cmd_data[7] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold253 (.A(uo_out[5]),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold254 (.A(\core.lsu.spi.addr[10] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold255 (.A(\core.fetch.data[1] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold256 (.A(uo_out[2]),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold257 (.A(\core.f2e_addr[12] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold258 (.A(\core.f2e_addr[6] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold259 (.A(\core.gpio.stray_data_i[24] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold260 (.A(_00018_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold261 (.A(_01002_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold262 (.A(\core.e2m_data[15] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold263 (.A(_00264_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold264 (.A(\core.e2m_data[11] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold265 (.A(\core.work.registers.tmp[28] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold266 (.A(\core.e2m_data[31] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold267 (.A(\core.f2e_addr[3] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold268 (.A(_00252_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold269 (.A(\core.work.registers.tmp[10] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold270 (.A(\core.gpio.stray_data_i[20] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold271 (.A(\core.work.registers.tmp[29] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold272 (.A(_00576_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold273 (.A(\core.fetch.spi_reader.addr[2] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold274 (.A(\core.e2m_data[2] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold275 (.A(\core.fetch.rd_addr_i[13] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold276 (.A(_00325_),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold277 (.A(\core.fetch.rd_addr_i[11] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold278 (.A(_00323_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold279 (.A(\core.lsu.spi.buffer[1] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold280 (.A(\core.e2m_data[9] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold281 (.A(_00104_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold282 (.A(_00251_),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold283 (.A(uo_out[6]),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold284 (.A(uo_out[4]),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold285 (.A(\core.fetch.data[11] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold286 (.A(\core.lsu.spi.buffer[2] ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold287 (.A(\core.fetch.data[12] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold288 (.A(_00197_),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold289 (.A(\core.e2m_data[14] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold290 (.A(\core.fetch.spi_reader.addr[5] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold291 (.A(\core.lsu.spi.buffer[4] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold292 (.A(\core.work.registers.tmp[26] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold293 (.A(\core.work.registers.tmp[18] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold294 (.A(\core.gpio.stray_data_i[18] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold295 (.A(\core.gpio.stray_data_i[6] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold296 (.A(\core.gpio.stray_data_i[16] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold297 (.A(_00360_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold298 (.A(\core.lsu.spi.counter[0] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold299 (.A(_00413_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold300 (.A(\core.fetch.spi_reader.addr[10] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold301 (.A(\core.f2e_inst[2] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold302 (.A(_00421_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold303 (.A(\core.f2e_inst[3] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold304 (.A(_00422_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold305 (.A(uo_out[3]),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold306 (.A(uo_out[0]),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold307 (.A(\core.e2m_data[28] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold308 (.A(_00053_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold309 (.A(_02098_),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold310 (.A(_00282_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold311 (.A(\core.work.alu.is_mem ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold312 (.A(\core.gpio.stray_data_i[31] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold313 (.A(\core.gpio.stray_data_i[3] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold314 (.A(\core.f2e_addr[14] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold315 (.A(\core.f2e_addr[9] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold316 (.A(\core.work.registers.wr_reg[2] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold317 (.A(\core.lsu.spi.addr[1] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold318 (.A(\core.gpio.stray_data_i[19] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold319 (.A(\core.fetch.spi_reader.addr[6] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold320 (.A(\core.gpio.stray_data_i[23] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold321 (.A(\core.fetch.spi_reader.addr[8] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold322 (.A(\core.lsu.spi.buffer[7] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold323 (.A(\core.fetch.spi_reader.counter[0] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold324 (.A(_00050_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold325 (.A(_02141_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold326 (.A(_00284_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold327 (.A(_00034_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold328 (.A(_02286_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold329 (.A(_00291_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold330 (.A(\core.f2e_addr[11] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold331 (.A(_00260_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold332 (.A(\core.gpio.stray_data_i[5] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold333 (.A(_00349_),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold334 (.A(\core.f2e_inst[11] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold335 (.A(\core.work.registers.wr_reg[3] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold336 (.A(\core.lsu.state[1] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold337 (.A(_00337_),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold338 (.A(\core.gpio.stray_data_i[7] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold339 (.A(\core.work.registers.tmp[3] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold340 (.A(\core.fetch.spi_reader.addr[7] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold341 (.A(\core.gpio.stray_data_i[2] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold342 (.A(_00346_),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold343 (.A(\core.f2e_addr[5] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold344 (.A(\core.work.alu.sval2[7] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold345 (.A(\core.gpio.stray_data_i[15] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold346 (.A(\core.gpio.stray_data_i[26] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold347 (.A(\core.work.alu.sval2[8] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold348 (.A(_00272_),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold349 (.A(\core.e2m_addr[4] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold350 (.A(\core.fetch.spi_reader.addr[13] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold351 (.A(\core.f2e_inst[7] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold352 (.A(_00426_),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold353 (.A(\core.e2m_addr[18] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold354 (.A(_00026_),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold355 (.A(_02363_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold356 (.A(_00295_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold357 (.A(\core.f2e_inst[4] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold358 (.A(\core.gpio.stray_data_i[12] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold359 (.A(_00356_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold360 (.A(\core.f2e_inst[14] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold361 (.A(\core.lsu.spi.addr[3] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold362 (.A(\core.lsu.spi.state[1] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold363 (.A(_00408_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold364 (.A(\core.gpio.stray_data_i[11] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold365 (.A(_00355_),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold366 (.A(_00029_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold367 (.A(\core.f2e_inst[9] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold368 (.A(\core.gpio.stray_data_i[14] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold369 (.A(_00358_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold370 (.A(\core.gpio.stray_data_i[0] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold371 (.A(\core.gpio.stray_data_i[9] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold372 (.A(_00353_),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold373 (.A(\core.gpio.stray_data_i[10] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold374 (.A(\core.lsu.spi.buffer[0] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold375 (.A(_00055_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold376 (.A(_01128_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold377 (.A(_00001_),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold378 (.A(\core.gpio.stray_data_i[8] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold379 (.A(\core.fetch.rd_addr_i[9] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold380 (.A(\core.gpio.stray_data_i[4] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold381 (.A(\core.lsu.state[0] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold382 (.A(_00336_),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold383 (.A(\core.lsu.spi.buffer[3] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold384 (.A(\core.fetch.spi_reader.addr[1] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold385 (.A(\core.work.alu.sval2[13] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold386 (.A(_00277_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold387 (.A(\core.work.registers.state[1] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold388 (.A(_00545_),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold389 (.A(\core.e2m_addr[1] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold390 (.A(_00548_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold391 (.A(\core.lsu.spi.state[2] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold392 (.A(\core.gpio.stray_data_i[21] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold393 (.A(_00365_),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold394 (.A(\core.work.alu.sval2[11] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold395 (.A(\core.lsu.spi.buffer[6] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold396 (.A(\core.work.registers.tmp[16] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold397 (.A(_00563_),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold398 (.A(\core.gpio.stray_data_i[13] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold399 (.A(\core.gpio.stray_data_i[22] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold400 (.A(_00366_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold401 (.A(\core.f2e_inst[13] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold402 (.A(\core.work.alu.sval2[3] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold403 (.A(_00267_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold404 (.A(\core.f2e_addr[10] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold405 (.A(\core.gpio.stray_data_i[17] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold406 (.A(\core.work.registers.tmp[15] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold407 (.A(\core.work.registers.state[0] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold408 (.A(_00544_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold409 (.A(\core.work.registers.tmp[4] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold410 (.A(_00119_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold411 (.A(\core.gpio.stray_data_i[29] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold412 (.A(\core.gpio.stray_data_i[27] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold413 (.A(\core.gpio.stray_data_i[30] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold414 (.A(\core.work.registers.tmp[11] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold415 (.A(\core.work.registers.tmp[24] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold416 (.A(\core.work.registers.tmp[31] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold417 (.A(\core.work.alu.sval2[15] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold418 (.A(_00279_),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold419 (.A(\core.e2m_addr[2] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold420 (.A(\core.work.registers.tmp[25] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold421 (.A(\core.work.alu.sval2[14] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold422 (.A(\core.f2e_addr[8] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold423 (.A(\core.work.alu.sval2[21] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold424 (.A(\core.lsu.spi.addr[11] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold425 (.A(_00402_),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold426 (.A(\core.fetch.spi_reader.state[0] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold427 (.A(_00246_),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold428 (.A(\core.work.registers.tmp[30] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold429 (.A(\core.work.alu.sval2[16] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold430 (.A(_00294_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold431 (.A(\core.gpio.stray_data_i[25] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold432 (.A(\core.gpio.stray_data_i[1] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold433 (.A(\core.fetch.rd_addr_i[12] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold434 (.A(\core.fetch.data_size[0] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold435 (.A(_00217_),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold436 (.A(\core.work.alu.sval2[26] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold437 (.A(_00287_),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold438 (.A(\core.e2m_addr[16] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold439 (.A(\core.f2e_inst[15] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold440 (.A(\core.fetch.spi_reader.addr[11] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold441 (.A(\core.fetch.data_size[2] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold442 (.A(_00219_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold443 (.A(_00022_),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold444 (.A(\core.fetch.data_size[1] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold445 (.A(\core.work.registers.tmp[21] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold446 (.A(\core.fetch.spi_reader.addr[9] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold447 (.A(\core.gpio.stray_data_i[28] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold448 (.A(_00114_),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold449 (.A(\core.f2e_inst[6] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold450 (.A(_00425_),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold451 (.A(\core.fetch.inst_size[1] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold452 (.A(\core.lsu.spi.buffer[5] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold453 (.A(_00388_),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold454 (.A(\core.fetch.rd_addr_i[8] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold455 (.A(_00045_),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold456 (.A(_02196_),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold457 (.A(_00286_),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold458 (.A(\core.f2e_inst[10] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold459 (.A(\core.fetch.rd_addr_i[2] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold460 (.A(\core.e2m_addr[22] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold461 (.A(\core.work.alu.sval2[0] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold462 (.A(_02115_),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold463 (.A(\core.work.registers.tmp[14] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold464 (.A(\core.lsu.spi.addr[13] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold465 (.A(_00404_),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold466 (.A(\core.work.registers.tmp[9] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold467 (.A(\core.f2e_inst[5] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold468 (.A(\core.e2m_addr[0] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold469 (.A(\core.e2m_addr[19] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold470 (.A(\core.f2e_inst[12] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold471 (.A(\core.work.alu.sval2[12] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold472 (.A(_00276_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold473 (.A(\core.e2m_addr[23] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold474 (.A(\core.fetch.spi_reader.state[2] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold475 (.A(\core.work.registers.tmp[20] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold476 (.A(\core.work.alu.sval2[1] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold477 (.A(\core.work.alu.sval2[28] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold478 (.A(_00285_),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold479 (.A(\core.fetch.rd_addr_i[3] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold480 (.A(_00315_),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold481 (.A(\core.lsu.spi.state[0] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold482 (.A(\core.work.registers.tmp[2] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold483 (.A(\core.work.alu.sval2[25] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold484 (.A(_02222_),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold485 (.A(\core.work.alu.ls_size_b ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold486 (.A(\core.fetch.rd_addr_i[4] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold487 (.A(\core.work.alu.sval2[6] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold488 (.A(\core.lsu.is_byte ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold489 (.A(\core.f2e_inst[1] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold490 (.A(_00420_),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold491 (.A(\core.work.alu.sval2[5] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold492 (.A(\core.fetch.state[1] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold493 (.A(\core.work.alu.sval2[29] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold494 (.A(\core.gpio.stray_wr_i ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold495 (.A(_00123_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold496 (.A(\core.work.registers.tmp[8] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold497 (.A(_00555_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold498 (.A(\core.work.alu.sval2[24] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold499 (.A(_00293_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold500 (.A(_00113_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold501 (.A(_00498_),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold502 (.A(\core.f2e_inst[0] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold503 (.A(_00419_),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold504 (.A(\core.work.state[0] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold505 (.A(_02322_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold506 (.A(_00292_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold507 (.A(\core.fetch.cmd_valid ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold508 (.A(\core.e2m_addr[24] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold509 (.A(\core.e2m_addr[17] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold510 (.A(\core.work.alu.is_sign ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold511 (.A(\core.lsu.spi.addr[7] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold512 (.A(uio_out[0]),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold513 (.A(_00000_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold514 (.A(\core.e2m_addr[3] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold515 (.A(_00096_),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold516 (.A(_00098_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold517 (.A(_01422_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold518 (.A(\core.e2m_addr[25] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold519 (.A(\core.f2e_addr[7] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold520 (.A(\core.work.alu.sval2[9] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold521 (.A(\core.e2m_addr[11] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold522 (.A(_00099_),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold523 (.A(_01426_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold524 (.A(_00225_),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold525 (.A(\core.lsu.write_index[2] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold526 (.A(_00412_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold527 (.A(_00112_),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold528 (.A(\core.work.alu.is_wr ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold529 (.A(\core.fetch.cmd_data[2] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold530 (.A(\core.e2m_addr[27] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold531 (.A(\core.f2e_addr[1] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold532 (.A(\core.work.state[1] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold533 (.A(_00101_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold534 (.A(_01442_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold535 (.A(_00100_),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold536 (.A(_00226_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold537 (.A(\core.e2m_addr[8] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold538 (.A(_00103_),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold539 (.A(_01450_),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold540 (.A(\core.e2m_addr[0] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold541 (.A(_00123_),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold542 (.A(\core.f2e_inst[9] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold543 (.A(\core.fetch.inst_size[1] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold544 (.A(\core.gpio.stray_data_i[3] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold545 (.A(\core.e2m_addr[0] ),
    .X(net900));
 sg13g2_antennanp ANTENNA_1 (.A(_00283_));
 sg13g2_antennanp ANTENNA_2 (.A(_01383_));
 sg13g2_antennanp ANTENNA_3 (.A(_04230_));
 sg13g2_antennanp ANTENNA_4 (.A(_04262_));
 sg13g2_antennanp ANTENNA_5 (.A(_04718_));
 sg13g2_antennanp ANTENNA_6 (.A(_04781_));
 sg13g2_antennanp ANTENNA_7 (.A(_04882_));
 sg13g2_antennanp ANTENNA_8 (.A(clk));
 sg13g2_antennanp ANTENNA_9 (.A(clk));
 sg13g2_antennanp ANTENNA_10 (.A(uio_out[4]));
 sg13g2_antennanp ANTENNA_11 (.A(uo_out[0]));
 sg13g2_antennanp ANTENNA_12 (.A(uo_out[0]));
 sg13g2_antennanp ANTENNA_13 (.A(uo_out[3]));
 sg13g2_antennanp ANTENNA_14 (.A(uo_out[3]));
 sg13g2_antennanp ANTENNA_15 (.A(uo_out[4]));
 sg13g2_antennanp ANTENNA_16 (.A(uo_out[4]));
 sg13g2_antennanp ANTENNA_17 (.A(uo_out[6]));
 sg13g2_antennanp ANTENNA_18 (.A(uo_out[6]));
 sg13g2_antennanp ANTENNA_19 (.A(_00283_));
 sg13g2_antennanp ANTENNA_20 (.A(_04230_));
 sg13g2_antennanp ANTENNA_21 (.A(_04262_));
 sg13g2_antennanp ANTENNA_22 (.A(_04718_));
 sg13g2_antennanp ANTENNA_23 (.A(_04781_));
 sg13g2_antennanp ANTENNA_24 (.A(_04882_));
 sg13g2_antennanp ANTENNA_25 (.A(clk));
 sg13g2_antennanp ANTENNA_26 (.A(clk));
 sg13g2_antennanp ANTENNA_27 (.A(uio_out[4]));
 sg13g2_antennanp ANTENNA_28 (.A(uio_out[4]));
 sg13g2_antennanp ANTENNA_29 (.A(uo_out[0]));
 sg13g2_antennanp ANTENNA_30 (.A(uo_out[0]));
 sg13g2_antennanp ANTENNA_31 (.A(uo_out[3]));
 sg13g2_antennanp ANTENNA_32 (.A(uo_out[3]));
 sg13g2_antennanp ANTENNA_33 (.A(uo_out[4]));
 sg13g2_antennanp ANTENNA_34 (.A(uo_out[4]));
 sg13g2_antennanp ANTENNA_35 (.A(uo_out[6]));
 sg13g2_antennanp ANTENNA_36 (.A(uo_out[6]));
 sg13g2_antennanp ANTENNA_37 (.A(_00283_));
 sg13g2_antennanp ANTENNA_38 (.A(_04230_));
 sg13g2_antennanp ANTENNA_39 (.A(_04262_));
 sg13g2_antennanp ANTENNA_40 (.A(_04718_));
 sg13g2_antennanp ANTENNA_41 (.A(_04781_));
 sg13g2_antennanp ANTENNA_42 (.A(clk));
 sg13g2_antennanp ANTENNA_43 (.A(clk));
 sg13g2_antennanp ANTENNA_44 (.A(uio_out[4]));
 sg13g2_antennanp ANTENNA_45 (.A(uio_out[4]));
 sg13g2_antennanp ANTENNA_46 (.A(uo_out[0]));
 sg13g2_antennanp ANTENNA_47 (.A(uo_out[0]));
 sg13g2_antennanp ANTENNA_48 (.A(uo_out[3]));
 sg13g2_antennanp ANTENNA_49 (.A(uo_out[3]));
 sg13g2_antennanp ANTENNA_50 (.A(uo_out[4]));
 sg13g2_antennanp ANTENNA_51 (.A(uo_out[4]));
 sg13g2_antennanp ANTENNA_52 (.A(uo_out[6]));
 sg13g2_antennanp ANTENNA_53 (.A(uo_out[6]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_fill_1 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_67 ();
 sg13g2_decap_8 FILLER_0_74 ();
 sg13g2_decap_8 FILLER_0_81 ();
 sg13g2_decap_4 FILLER_0_88 ();
 sg13g2_fill_1 FILLER_0_92 ();
 sg13g2_fill_2 FILLER_0_98 ();
 sg13g2_fill_1 FILLER_0_100 ();
 sg13g2_fill_1 FILLER_0_118 ();
 sg13g2_decap_8 FILLER_0_136 ();
 sg13g2_decap_4 FILLER_0_143 ();
 sg13g2_fill_1 FILLER_0_164 ();
 sg13g2_decap_4 FILLER_0_182 ();
 sg13g2_fill_2 FILLER_0_186 ();
 sg13g2_decap_4 FILLER_0_205 ();
 sg13g2_fill_1 FILLER_0_209 ();
 sg13g2_fill_1 FILLER_0_218 ();
 sg13g2_decap_8 FILLER_0_227 ();
 sg13g2_decap_8 FILLER_0_251 ();
 sg13g2_fill_2 FILLER_0_258 ();
 sg13g2_fill_1 FILLER_0_260 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_fill_2 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_321 ();
 sg13g2_fill_2 FILLER_0_328 ();
 sg13g2_decap_4 FILLER_0_347 ();
 sg13g2_fill_2 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_4 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_4 FILLER_0_480 ();
 sg13g2_fill_2 FILLER_0_484 ();
 sg13g2_decap_8 FILLER_0_503 ();
 sg13g2_decap_8 FILLER_0_510 ();
 sg13g2_fill_2 FILLER_0_534 ();
 sg13g2_fill_1 FILLER_0_536 ();
 sg13g2_decap_8 FILLER_0_554 ();
 sg13g2_decap_4 FILLER_0_578 ();
 sg13g2_decap_8 FILLER_0_599 ();
 sg13g2_decap_8 FILLER_0_606 ();
 sg13g2_decap_4 FILLER_0_613 ();
 sg13g2_decap_8 FILLER_0_702 ();
 sg13g2_decap_4 FILLER_0_709 ();
 sg13g2_fill_2 FILLER_0_713 ();
 sg13g2_decap_8 FILLER_0_740 ();
 sg13g2_decap_8 FILLER_0_764 ();
 sg13g2_decap_8 FILLER_0_771 ();
 sg13g2_decap_8 FILLER_0_778 ();
 sg13g2_decap_8 FILLER_0_785 ();
 sg13g2_decap_8 FILLER_0_792 ();
 sg13g2_decap_8 FILLER_0_799 ();
 sg13g2_decap_8 FILLER_0_806 ();
 sg13g2_decap_8 FILLER_0_813 ();
 sg13g2_decap_8 FILLER_0_820 ();
 sg13g2_decap_8 FILLER_0_827 ();
 sg13g2_decap_8 FILLER_0_834 ();
 sg13g2_decap_8 FILLER_0_841 ();
 sg13g2_decap_8 FILLER_0_848 ();
 sg13g2_decap_8 FILLER_0_855 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_4 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_46 ();
 sg13g2_fill_1 FILLER_1_51 ();
 sg13g2_decap_8 FILLER_1_69 ();
 sg13g2_decap_8 FILLER_1_76 ();
 sg13g2_decap_4 FILLER_1_83 ();
 sg13g2_decap_4 FILLER_1_121 ();
 sg13g2_fill_1 FILLER_1_125 ();
 sg13g2_fill_2 FILLER_1_143 ();
 sg13g2_fill_2 FILLER_1_170 ();
 sg13g2_decap_4 FILLER_1_206 ();
 sg13g2_fill_1 FILLER_1_210 ();
 sg13g2_fill_1 FILLER_1_279 ();
 sg13g2_fill_1 FILLER_1_348 ();
 sg13g2_fill_2 FILLER_1_400 ();
 sg13g2_decap_4 FILLER_1_419 ();
 sg13g2_fill_2 FILLER_1_423 ();
 sg13g2_fill_1 FILLER_1_430 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_4 FILLER_1_462 ();
 sg13g2_fill_1 FILLER_1_466 ();
 sg13g2_fill_2 FILLER_1_484 ();
 sg13g2_fill_2 FILLER_1_509 ();
 sg13g2_decap_4 FILLER_1_528 ();
 sg13g2_fill_2 FILLER_1_532 ();
 sg13g2_fill_1 FILLER_1_551 ();
 sg13g2_fill_2 FILLER_1_556 ();
 sg13g2_fill_1 FILLER_1_558 ();
 sg13g2_decap_8 FILLER_1_576 ();
 sg13g2_decap_8 FILLER_1_583 ();
 sg13g2_decap_8 FILLER_1_646 ();
 sg13g2_fill_1 FILLER_1_653 ();
 sg13g2_decap_8 FILLER_1_676 ();
 sg13g2_decap_8 FILLER_1_683 ();
 sg13g2_decap_4 FILLER_1_707 ();
 sg13g2_fill_1 FILLER_1_711 ();
 sg13g2_fill_1 FILLER_1_746 ();
 sg13g2_decap_8 FILLER_1_781 ();
 sg13g2_decap_8 FILLER_1_788 ();
 sg13g2_decap_8 FILLER_1_795 ();
 sg13g2_decap_8 FILLER_1_802 ();
 sg13g2_decap_8 FILLER_1_809 ();
 sg13g2_decap_8 FILLER_1_816 ();
 sg13g2_decap_8 FILLER_1_823 ();
 sg13g2_decap_8 FILLER_1_830 ();
 sg13g2_decap_8 FILLER_1_837 ();
 sg13g2_decap_8 FILLER_1_844 ();
 sg13g2_decap_8 FILLER_1_851 ();
 sg13g2_decap_4 FILLER_1_858 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_4 FILLER_2_7 ();
 sg13g2_fill_1 FILLER_2_11 ();
 sg13g2_fill_2 FILLER_2_46 ();
 sg13g2_fill_1 FILLER_2_48 ();
 sg13g2_fill_2 FILLER_2_66 ();
 sg13g2_fill_1 FILLER_2_68 ();
 sg13g2_decap_4 FILLER_2_86 ();
 sg13g2_fill_2 FILLER_2_90 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_fill_2 FILLER_2_116 ();
 sg13g2_fill_1 FILLER_2_118 ();
 sg13g2_decap_4 FILLER_2_136 ();
 sg13g2_decap_4 FILLER_2_162 ();
 sg13g2_fill_2 FILLER_2_166 ();
 sg13g2_fill_1 FILLER_2_193 ();
 sg13g2_fill_2 FILLER_2_211 ();
 sg13g2_fill_2 FILLER_2_229 ();
 sg13g2_decap_4 FILLER_2_253 ();
 sg13g2_fill_2 FILLER_2_274 ();
 sg13g2_fill_1 FILLER_2_276 ();
 sg13g2_decap_4 FILLER_2_299 ();
 sg13g2_fill_1 FILLER_2_303 ();
 sg13g2_decap_8 FILLER_2_321 ();
 sg13g2_decap_4 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_337 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_419 ();
 sg13g2_fill_2 FILLER_2_426 ();
 sg13g2_decap_8 FILLER_2_445 ();
 sg13g2_fill_2 FILLER_2_452 ();
 sg13g2_decap_4 FILLER_2_471 ();
 sg13g2_fill_2 FILLER_2_475 ();
 sg13g2_fill_1 FILLER_2_515 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_fill_1 FILLER_2_546 ();
 sg13g2_fill_2 FILLER_2_570 ();
 sg13g2_fill_1 FILLER_2_585 ();
 sg13g2_fill_1 FILLER_2_603 ();
 sg13g2_fill_2 FILLER_2_609 ();
 sg13g2_fill_1 FILLER_2_611 ();
 sg13g2_decap_8 FILLER_2_618 ();
 sg13g2_decap_8 FILLER_2_625 ();
 sg13g2_decap_4 FILLER_2_649 ();
 sg13g2_fill_2 FILLER_2_653 ();
 sg13g2_fill_2 FILLER_2_672 ();
 sg13g2_fill_1 FILLER_2_674 ();
 sg13g2_decap_4 FILLER_2_709 ();
 sg13g2_fill_2 FILLER_2_713 ();
 sg13g2_decap_8 FILLER_2_723 ();
 sg13g2_decap_8 FILLER_2_730 ();
 sg13g2_decap_8 FILLER_2_737 ();
 sg13g2_decap_8 FILLER_2_744 ();
 sg13g2_decap_4 FILLER_2_768 ();
 sg13g2_fill_2 FILLER_2_789 ();
 sg13g2_decap_8 FILLER_2_808 ();
 sg13g2_decap_8 FILLER_2_815 ();
 sg13g2_decap_8 FILLER_2_822 ();
 sg13g2_decap_8 FILLER_2_829 ();
 sg13g2_decap_8 FILLER_2_836 ();
 sg13g2_decap_8 FILLER_2_843 ();
 sg13g2_decap_8 FILLER_2_850 ();
 sg13g2_decap_4 FILLER_2_857 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_7 ();
 sg13g2_decap_4 FILLER_3_25 ();
 sg13g2_fill_1 FILLER_3_29 ();
 sg13g2_decap_4 FILLER_3_64 ();
 sg13g2_decap_8 FILLER_3_80 ();
 sg13g2_decap_4 FILLER_3_87 ();
 sg13g2_fill_2 FILLER_3_91 ();
 sg13g2_decap_4 FILLER_3_110 ();
 sg13g2_fill_1 FILLER_3_114 ();
 sg13g2_decap_8 FILLER_3_132 ();
 sg13g2_decap_8 FILLER_3_139 ();
 sg13g2_fill_2 FILLER_3_146 ();
 sg13g2_decap_4 FILLER_3_165 ();
 sg13g2_fill_1 FILLER_3_169 ();
 sg13g2_fill_2 FILLER_3_184 ();
 sg13g2_fill_2 FILLER_3_196 ();
 sg13g2_fill_1 FILLER_3_198 ();
 sg13g2_fill_2 FILLER_3_205 ();
 sg13g2_fill_2 FILLER_3_215 ();
 sg13g2_fill_1 FILLER_3_217 ();
 sg13g2_fill_1 FILLER_3_234 ();
 sg13g2_decap_4 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_279 ();
 sg13g2_decap_4 FILLER_3_286 ();
 sg13g2_decap_8 FILLER_3_307 ();
 sg13g2_fill_2 FILLER_3_320 ();
 sg13g2_fill_1 FILLER_3_322 ();
 sg13g2_fill_1 FILLER_3_361 ();
 sg13g2_fill_2 FILLER_3_384 ();
 sg13g2_fill_1 FILLER_3_386 ();
 sg13g2_fill_1 FILLER_3_426 ();
 sg13g2_decap_8 FILLER_3_444 ();
 sg13g2_fill_2 FILLER_3_451 ();
 sg13g2_fill_1 FILLER_3_453 ();
 sg13g2_decap_4 FILLER_3_471 ();
 sg13g2_fill_1 FILLER_3_475 ();
 sg13g2_fill_1 FILLER_3_529 ();
 sg13g2_fill_2 FILLER_3_548 ();
 sg13g2_fill_2 FILLER_3_562 ();
 sg13g2_fill_1 FILLER_3_564 ();
 sg13g2_fill_1 FILLER_3_594 ();
 sg13g2_fill_2 FILLER_3_630 ();
 sg13g2_fill_2 FILLER_3_653 ();
 sg13g2_decap_4 FILLER_3_678 ();
 sg13g2_decap_4 FILLER_3_764 ();
 sg13g2_fill_2 FILLER_3_768 ();
 sg13g2_decap_8 FILLER_3_821 ();
 sg13g2_decap_8 FILLER_3_828 ();
 sg13g2_decap_8 FILLER_3_835 ();
 sg13g2_decap_8 FILLER_3_842 ();
 sg13g2_decap_8 FILLER_3_849 ();
 sg13g2_decap_4 FILLER_3_856 ();
 sg13g2_fill_2 FILLER_3_860 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_24 ();
 sg13g2_decap_4 FILLER_4_31 ();
 sg13g2_fill_2 FILLER_4_35 ();
 sg13g2_decap_4 FILLER_4_42 ();
 sg13g2_fill_2 FILLER_4_46 ();
 sg13g2_fill_2 FILLER_4_90 ();
 sg13g2_fill_2 FILLER_4_109 ();
 sg13g2_fill_1 FILLER_4_123 ();
 sg13g2_fill_1 FILLER_4_142 ();
 sg13g2_fill_2 FILLER_4_190 ();
 sg13g2_fill_1 FILLER_4_192 ();
 sg13g2_decap_4 FILLER_4_205 ();
 sg13g2_fill_1 FILLER_4_209 ();
 sg13g2_fill_2 FILLER_4_234 ();
 sg13g2_fill_1 FILLER_4_236 ();
 sg13g2_decap_4 FILLER_4_255 ();
 sg13g2_decap_4 FILLER_4_277 ();
 sg13g2_fill_2 FILLER_4_281 ();
 sg13g2_decap_4 FILLER_4_327 ();
 sg13g2_fill_1 FILLER_4_331 ();
 sg13g2_fill_1 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_421 ();
 sg13g2_fill_1 FILLER_4_425 ();
 sg13g2_decap_8 FILLER_4_431 ();
 sg13g2_fill_2 FILLER_4_438 ();
 sg13g2_fill_1 FILLER_4_474 ();
 sg13g2_decap_4 FILLER_4_527 ();
 sg13g2_fill_2 FILLER_4_567 ();
 sg13g2_fill_1 FILLER_4_569 ();
 sg13g2_fill_2 FILLER_4_582 ();
 sg13g2_fill_1 FILLER_4_584 ();
 sg13g2_decap_4 FILLER_4_602 ();
 sg13g2_fill_1 FILLER_4_632 ();
 sg13g2_decap_8 FILLER_4_656 ();
 sg13g2_decap_8 FILLER_4_720 ();
 sg13g2_decap_8 FILLER_4_727 ();
 sg13g2_decap_8 FILLER_4_746 ();
 sg13g2_decap_8 FILLER_4_753 ();
 sg13g2_decap_8 FILLER_4_760 ();
 sg13g2_decap_8 FILLER_4_767 ();
 sg13g2_decap_4 FILLER_4_774 ();
 sg13g2_decap_4 FILLER_4_786 ();
 sg13g2_decap_8 FILLER_4_801 ();
 sg13g2_fill_2 FILLER_4_830 ();
 sg13g2_decap_8 FILLER_4_849 ();
 sg13g2_decap_4 FILLER_4_856 ();
 sg13g2_fill_2 FILLER_4_860 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_9 ();
 sg13g2_decap_4 FILLER_5_27 ();
 sg13g2_fill_2 FILLER_5_31 ();
 sg13g2_decap_4 FILLER_5_50 ();
 sg13g2_fill_1 FILLER_5_54 ();
 sg13g2_fill_1 FILLER_5_73 ();
 sg13g2_decap_8 FILLER_5_90 ();
 sg13g2_fill_2 FILLER_5_97 ();
 sg13g2_fill_1 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_145 ();
 sg13g2_decap_8 FILLER_5_152 ();
 sg13g2_decap_4 FILLER_5_159 ();
 sg13g2_fill_1 FILLER_5_181 ();
 sg13g2_fill_2 FILLER_5_230 ();
 sg13g2_fill_1 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_4 FILLER_5_291 ();
 sg13g2_fill_2 FILLER_5_355 ();
 sg13g2_fill_2 FILLER_5_363 ();
 sg13g2_fill_2 FILLER_5_383 ();
 sg13g2_fill_1 FILLER_5_385 ();
 sg13g2_fill_1 FILLER_5_392 ();
 sg13g2_fill_1 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_424 ();
 sg13g2_fill_2 FILLER_5_431 ();
 sg13g2_fill_1 FILLER_5_433 ();
 sg13g2_decap_4 FILLER_5_451 ();
 sg13g2_decap_4 FILLER_5_472 ();
 sg13g2_fill_2 FILLER_5_505 ();
 sg13g2_fill_1 FILLER_5_524 ();
 sg13g2_fill_1 FILLER_5_553 ();
 sg13g2_decap_4 FILLER_5_558 ();
 sg13g2_decap_4 FILLER_5_579 ();
 sg13g2_fill_2 FILLER_5_611 ();
 sg13g2_fill_1 FILLER_5_613 ();
 sg13g2_decap_8 FILLER_5_622 ();
 sg13g2_fill_1 FILLER_5_629 ();
 sg13g2_fill_1 FILLER_5_638 ();
 sg13g2_fill_1 FILLER_5_657 ();
 sg13g2_decap_8 FILLER_5_675 ();
 sg13g2_fill_2 FILLER_5_699 ();
 sg13g2_fill_1 FILLER_5_701 ();
 sg13g2_fill_1 FILLER_5_727 ();
 sg13g2_fill_1 FILLER_5_734 ();
 sg13g2_decap_8 FILLER_5_753 ();
 sg13g2_fill_2 FILLER_5_760 ();
 sg13g2_fill_1 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_851 ();
 sg13g2_decap_4 FILLER_5_858 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_2 ();
 sg13g2_decap_8 FILLER_6_20 ();
 sg13g2_decap_4 FILLER_6_27 ();
 sg13g2_fill_2 FILLER_6_31 ();
 sg13g2_fill_2 FILLER_6_50 ();
 sg13g2_fill_1 FILLER_6_52 ();
 sg13g2_fill_2 FILLER_6_115 ();
 sg13g2_fill_2 FILLER_6_145 ();
 sg13g2_fill_1 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_decap_4 FILLER_6_172 ();
 sg13g2_fill_1 FILLER_6_176 ();
 sg13g2_decap_4 FILLER_6_188 ();
 sg13g2_fill_2 FILLER_6_197 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_fill_1 FILLER_6_210 ();
 sg13g2_fill_1 FILLER_6_219 ();
 sg13g2_fill_2 FILLER_6_228 ();
 sg13g2_fill_1 FILLER_6_230 ();
 sg13g2_fill_2 FILLER_6_248 ();
 sg13g2_fill_1 FILLER_6_256 ();
 sg13g2_decap_4 FILLER_6_263 ();
 sg13g2_fill_1 FILLER_6_267 ();
 sg13g2_fill_2 FILLER_6_278 ();
 sg13g2_fill_1 FILLER_6_280 ();
 sg13g2_fill_1 FILLER_6_298 ();
 sg13g2_fill_2 FILLER_6_329 ();
 sg13g2_decap_4 FILLER_6_358 ();
 sg13g2_fill_2 FILLER_6_368 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_414 ();
 sg13g2_decap_8 FILLER_6_419 ();
 sg13g2_decap_8 FILLER_6_426 ();
 sg13g2_fill_1 FILLER_6_433 ();
 sg13g2_decap_4 FILLER_6_530 ();
 sg13g2_decap_8 FILLER_6_538 ();
 sg13g2_fill_1 FILLER_6_545 ();
 sg13g2_decap_4 FILLER_6_579 ();
 sg13g2_decap_4 FILLER_6_600 ();
 sg13g2_decap_4 FILLER_6_621 ();
 sg13g2_fill_2 FILLER_6_625 ();
 sg13g2_fill_2 FILLER_6_633 ();
 sg13g2_fill_1 FILLER_6_635 ();
 sg13g2_decap_8 FILLER_6_653 ();
 sg13g2_decap_8 FILLER_6_660 ();
 sg13g2_fill_1 FILLER_6_667 ();
 sg13g2_fill_2 FILLER_6_692 ();
 sg13g2_fill_1 FILLER_6_694 ();
 sg13g2_fill_2 FILLER_6_720 ();
 sg13g2_fill_1 FILLER_6_728 ();
 sg13g2_fill_2 FILLER_6_779 ();
 sg13g2_fill_2 FILLER_6_793 ();
 sg13g2_fill_1 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_830 ();
 sg13g2_fill_2 FILLER_6_837 ();
 sg13g2_fill_1 FILLER_6_839 ();
 sg13g2_decap_4 FILLER_6_857 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_24 ();
 sg13g2_fill_1 FILLER_7_26 ();
 sg13g2_fill_2 FILLER_7_35 ();
 sg13g2_fill_1 FILLER_7_37 ();
 sg13g2_decap_4 FILLER_7_88 ();
 sg13g2_fill_1 FILLER_7_92 ();
 sg13g2_decap_4 FILLER_7_110 ();
 sg13g2_decap_4 FILLER_7_120 ();
 sg13g2_fill_2 FILLER_7_135 ();
 sg13g2_fill_2 FILLER_7_153 ();
 sg13g2_fill_1 FILLER_7_155 ();
 sg13g2_decap_8 FILLER_7_198 ();
 sg13g2_fill_1 FILLER_7_205 ();
 sg13g2_fill_2 FILLER_7_214 ();
 sg13g2_fill_1 FILLER_7_216 ();
 sg13g2_decap_4 FILLER_7_225 ();
 sg13g2_fill_2 FILLER_7_229 ();
 sg13g2_fill_1 FILLER_7_248 ();
 sg13g2_fill_2 FILLER_7_261 ();
 sg13g2_fill_2 FILLER_7_279 ();
 sg13g2_decap_8 FILLER_7_326 ();
 sg13g2_fill_2 FILLER_7_373 ();
 sg13g2_fill_1 FILLER_7_375 ();
 sg13g2_fill_2 FILLER_7_382 ();
 sg13g2_fill_1 FILLER_7_384 ();
 sg13g2_fill_1 FILLER_7_393 ();
 sg13g2_fill_2 FILLER_7_418 ();
 sg13g2_fill_1 FILLER_7_420 ();
 sg13g2_decap_4 FILLER_7_429 ();
 sg13g2_fill_2 FILLER_7_433 ();
 sg13g2_decap_4 FILLER_7_452 ();
 sg13g2_fill_1 FILLER_7_456 ();
 sg13g2_decap_4 FILLER_7_474 ();
 sg13g2_fill_1 FILLER_7_478 ();
 sg13g2_decap_8 FILLER_7_502 ();
 sg13g2_decap_8 FILLER_7_509 ();
 sg13g2_decap_8 FILLER_7_516 ();
 sg13g2_decap_8 FILLER_7_523 ();
 sg13g2_decap_8 FILLER_7_530 ();
 sg13g2_fill_2 FILLER_7_561 ();
 sg13g2_fill_2 FILLER_7_580 ();
 sg13g2_decap_4 FILLER_7_599 ();
 sg13g2_decap_4 FILLER_7_608 ();
 sg13g2_fill_1 FILLER_7_612 ();
 sg13g2_decap_8 FILLER_7_621 ();
 sg13g2_fill_2 FILLER_7_628 ();
 sg13g2_decap_4 FILLER_7_688 ();
 sg13g2_decap_4 FILLER_7_717 ();
 sg13g2_fill_2 FILLER_7_727 ();
 sg13g2_decap_4 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_765 ();
 sg13g2_fill_2 FILLER_7_772 ();
 sg13g2_fill_1 FILLER_7_774 ();
 sg13g2_fill_2 FILLER_7_804 ();
 sg13g2_fill_1 FILLER_7_806 ();
 sg13g2_decap_4 FILLER_7_858 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_9 ();
 sg13g2_decap_4 FILLER_8_27 ();
 sg13g2_fill_2 FILLER_8_31 ();
 sg13g2_fill_1 FILLER_8_67 ();
 sg13g2_decap_8 FILLER_8_131 ();
 sg13g2_fill_1 FILLER_8_138 ();
 sg13g2_decap_8 FILLER_8_164 ();
 sg13g2_fill_1 FILLER_8_171 ();
 sg13g2_decap_4 FILLER_8_193 ();
 sg13g2_fill_1 FILLER_8_197 ();
 sg13g2_fill_2 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_4 FILLER_8_231 ();
 sg13g2_fill_1 FILLER_8_235 ();
 sg13g2_decap_8 FILLER_8_253 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_decap_8 FILLER_8_291 ();
 sg13g2_fill_2 FILLER_8_298 ();
 sg13g2_decap_4 FILLER_8_327 ();
 sg13g2_fill_1 FILLER_8_331 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_fill_1 FILLER_8_356 ();
 sg13g2_fill_2 FILLER_8_373 ();
 sg13g2_fill_1 FILLER_8_375 ();
 sg13g2_decap_4 FILLER_8_407 ();
 sg13g2_fill_2 FILLER_8_411 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_fill_2 FILLER_8_434 ();
 sg13g2_fill_1 FILLER_8_436 ();
 sg13g2_decap_8 FILLER_8_454 ();
 sg13g2_fill_1 FILLER_8_461 ();
 sg13g2_decap_4 FILLER_8_479 ();
 sg13g2_fill_2 FILLER_8_483 ();
 sg13g2_decap_4 FILLER_8_507 ();
 sg13g2_fill_1 FILLER_8_511 ();
 sg13g2_decap_4 FILLER_8_537 ();
 sg13g2_fill_2 FILLER_8_541 ();
 sg13g2_fill_2 FILLER_8_551 ();
 sg13g2_fill_1 FILLER_8_553 ();
 sg13g2_fill_1 FILLER_8_562 ();
 sg13g2_decap_8 FILLER_8_580 ();
 sg13g2_fill_2 FILLER_8_587 ();
 sg13g2_fill_1 FILLER_8_638 ();
 sg13g2_fill_1 FILLER_8_649 ();
 sg13g2_decap_8 FILLER_8_655 ();
 sg13g2_fill_2 FILLER_8_662 ();
 sg13g2_fill_1 FILLER_8_664 ();
 sg13g2_decap_4 FILLER_8_689 ();
 sg13g2_fill_2 FILLER_8_701 ();
 sg13g2_fill_1 FILLER_8_703 ();
 sg13g2_fill_1 FILLER_8_721 ();
 sg13g2_fill_1 FILLER_8_786 ();
 sg13g2_fill_2 FILLER_8_793 ();
 sg13g2_fill_1 FILLER_8_795 ();
 sg13g2_fill_1 FILLER_8_814 ();
 sg13g2_decap_8 FILLER_8_849 ();
 sg13g2_decap_4 FILLER_8_856 ();
 sg13g2_fill_2 FILLER_8_860 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_32 ();
 sg13g2_decap_8 FILLER_9_51 ();
 sg13g2_fill_1 FILLER_9_58 ();
 sg13g2_decap_8 FILLER_9_87 ();
 sg13g2_decap_4 FILLER_9_94 ();
 sg13g2_fill_2 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_104 ();
 sg13g2_decap_8 FILLER_9_111 ();
 sg13g2_fill_2 FILLER_9_118 ();
 sg13g2_fill_1 FILLER_9_120 ();
 sg13g2_fill_1 FILLER_9_143 ();
 sg13g2_decap_4 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_9_206 ();
 sg13g2_fill_2 FILLER_9_213 ();
 sg13g2_fill_1 FILLER_9_215 ();
 sg13g2_fill_2 FILLER_9_238 ();
 sg13g2_fill_1 FILLER_9_240 ();
 sg13g2_decap_4 FILLER_9_258 ();
 sg13g2_decap_8 FILLER_9_267 ();
 sg13g2_fill_2 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_318 ();
 sg13g2_decap_8 FILLER_9_325 ();
 sg13g2_fill_2 FILLER_9_349 ();
 sg13g2_fill_1 FILLER_9_351 ();
 sg13g2_fill_1 FILLER_9_377 ();
 sg13g2_fill_1 FILLER_9_406 ();
 sg13g2_fill_2 FILLER_9_432 ();
 sg13g2_fill_1 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_443 ();
 sg13g2_fill_2 FILLER_9_450 ();
 sg13g2_fill_1 FILLER_9_457 ();
 sg13g2_fill_1 FILLER_9_479 ();
 sg13g2_fill_2 FILLER_9_506 ();
 sg13g2_decap_8 FILLER_9_533 ();
 sg13g2_decap_4 FILLER_9_557 ();
 sg13g2_fill_1 FILLER_9_561 ();
 sg13g2_fill_1 FILLER_9_602 ();
 sg13g2_fill_2 FILLER_9_640 ();
 sg13g2_decap_4 FILLER_9_665 ();
 sg13g2_fill_2 FILLER_9_691 ();
 sg13g2_decap_8 FILLER_9_710 ();
 sg13g2_fill_1 FILLER_9_717 ();
 sg13g2_decap_4 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_748 ();
 sg13g2_decap_8 FILLER_9_755 ();
 sg13g2_fill_1 FILLER_9_776 ();
 sg13g2_fill_2 FILLER_9_783 ();
 sg13g2_fill_1 FILLER_9_785 ();
 sg13g2_decap_8 FILLER_9_804 ();
 sg13g2_fill_2 FILLER_9_811 ();
 sg13g2_fill_1 FILLER_9_813 ();
 sg13g2_decap_8 FILLER_9_831 ();
 sg13g2_fill_1 FILLER_9_838 ();
 sg13g2_decap_4 FILLER_9_856 ();
 sg13g2_fill_2 FILLER_9_860 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_fill_2 FILLER_10_20 ();
 sg13g2_fill_1 FILLER_10_22 ();
 sg13g2_decap_8 FILLER_10_45 ();
 sg13g2_decap_8 FILLER_10_52 ();
 sg13g2_fill_2 FILLER_10_59 ();
 sg13g2_fill_2 FILLER_10_119 ();
 sg13g2_fill_1 FILLER_10_121 ();
 sg13g2_fill_1 FILLER_10_139 ();
 sg13g2_fill_1 FILLER_10_162 ();
 sg13g2_decap_4 FILLER_10_167 ();
 sg13g2_fill_2 FILLER_10_171 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_4 FILLER_10_196 ();
 sg13g2_fill_2 FILLER_10_200 ();
 sg13g2_fill_2 FILLER_10_278 ();
 sg13g2_fill_1 FILLER_10_280 ();
 sg13g2_decap_4 FILLER_10_298 ();
 sg13g2_fill_1 FILLER_10_302 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_fill_1 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_fill_2 FILLER_10_385 ();
 sg13g2_decap_4 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_fill_2 FILLER_10_459 ();
 sg13g2_fill_1 FILLER_10_461 ();
 sg13g2_decap_4 FILLER_10_479 ();
 sg13g2_fill_1 FILLER_10_493 ();
 sg13g2_fill_2 FILLER_10_506 ();
 sg13g2_fill_1 FILLER_10_508 ();
 sg13g2_fill_2 FILLER_10_517 ();
 sg13g2_fill_1 FILLER_10_519 ();
 sg13g2_fill_2 FILLER_10_537 ();
 sg13g2_decap_8 FILLER_10_556 ();
 sg13g2_decap_8 FILLER_10_563 ();
 sg13g2_decap_8 FILLER_10_578 ();
 sg13g2_decap_8 FILLER_10_585 ();
 sg13g2_fill_2 FILLER_10_592 ();
 sg13g2_decap_4 FILLER_10_619 ();
 sg13g2_fill_1 FILLER_10_623 ();
 sg13g2_fill_1 FILLER_10_635 ();
 sg13g2_decap_4 FILLER_10_670 ();
 sg13g2_fill_2 FILLER_10_674 ();
 sg13g2_decap_8 FILLER_10_688 ();
 sg13g2_decap_8 FILLER_10_695 ();
 sg13g2_decap_4 FILLER_10_702 ();
 sg13g2_fill_2 FILLER_10_706 ();
 sg13g2_decap_8 FILLER_10_713 ();
 sg13g2_fill_1 FILLER_10_720 ();
 sg13g2_fill_2 FILLER_10_745 ();
 sg13g2_fill_1 FILLER_10_747 ();
 sg13g2_fill_1 FILLER_10_810 ();
 sg13g2_fill_2 FILLER_10_828 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_88 ();
 sg13g2_decap_8 FILLER_11_95 ();
 sg13g2_fill_2 FILLER_11_102 ();
 sg13g2_fill_1 FILLER_11_104 ();
 sg13g2_decap_4 FILLER_11_122 ();
 sg13g2_fill_2 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_174 ();
 sg13g2_fill_2 FILLER_11_189 ();
 sg13g2_fill_1 FILLER_11_191 ();
 sg13g2_fill_1 FILLER_11_200 ();
 sg13g2_decap_4 FILLER_11_218 ();
 sg13g2_fill_2 FILLER_11_222 ();
 sg13g2_decap_8 FILLER_11_242 ();
 sg13g2_fill_2 FILLER_11_249 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_decap_8 FILLER_11_274 ();
 sg13g2_decap_8 FILLER_11_281 ();
 sg13g2_fill_2 FILLER_11_375 ();
 sg13g2_decap_4 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_fill_1 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_11_435 ();
 sg13g2_fill_1 FILLER_11_459 ();
 sg13g2_decap_4 FILLER_11_477 ();
 sg13g2_fill_1 FILLER_11_481 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_4 FILLER_11_535 ();
 sg13g2_fill_2 FILLER_11_539 ();
 sg13g2_decap_4 FILLER_11_569 ();
 sg13g2_fill_2 FILLER_11_573 ();
 sg13g2_fill_2 FILLER_11_596 ();
 sg13g2_fill_2 FILLER_11_603 ();
 sg13g2_fill_1 FILLER_11_605 ();
 sg13g2_decap_8 FILLER_11_612 ();
 sg13g2_fill_1 FILLER_11_619 ();
 sg13g2_decap_4 FILLER_11_655 ();
 sg13g2_fill_1 FILLER_11_696 ();
 sg13g2_decap_8 FILLER_11_720 ();
 sg13g2_fill_2 FILLER_11_727 ();
 sg13g2_fill_1 FILLER_11_729 ();
 sg13g2_fill_2 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_754 ();
 sg13g2_decap_4 FILLER_11_761 ();
 sg13g2_decap_8 FILLER_11_769 ();
 sg13g2_fill_2 FILLER_11_776 ();
 sg13g2_decap_4 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_806 ();
 sg13g2_fill_2 FILLER_11_813 ();
 sg13g2_fill_1 FILLER_11_815 ();
 sg13g2_decap_8 FILLER_11_820 ();
 sg13g2_decap_8 FILLER_11_827 ();
 sg13g2_decap_4 FILLER_11_834 ();
 sg13g2_decap_8 FILLER_11_855 ();
 sg13g2_fill_2 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_48 ();
 sg13g2_decap_4 FILLER_12_55 ();
 sg13g2_fill_1 FILLER_12_59 ();
 sg13g2_decap_8 FILLER_12_82 ();
 sg13g2_fill_1 FILLER_12_89 ();
 sg13g2_decap_4 FILLER_12_111 ();
 sg13g2_fill_1 FILLER_12_115 ();
 sg13g2_fill_1 FILLER_12_133 ();
 sg13g2_fill_1 FILLER_12_146 ();
 sg13g2_decap_8 FILLER_12_159 ();
 sg13g2_decap_8 FILLER_12_166 ();
 sg13g2_fill_1 FILLER_12_173 ();
 sg13g2_decap_8 FILLER_12_199 ();
 sg13g2_decap_4 FILLER_12_206 ();
 sg13g2_fill_2 FILLER_12_210 ();
 sg13g2_fill_1 FILLER_12_251 ();
 sg13g2_fill_2 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_327 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_fill_1 FILLER_12_371 ();
 sg13g2_fill_2 FILLER_12_395 ();
 sg13g2_fill_1 FILLER_12_397 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_425 ();
 sg13g2_fill_2 FILLER_12_460 ();
 sg13g2_fill_1 FILLER_12_462 ();
 sg13g2_fill_2 FILLER_12_480 ();
 sg13g2_decap_4 FILLER_12_509 ();
 sg13g2_decap_8 FILLER_12_530 ();
 sg13g2_decap_4 FILLER_12_537 ();
 sg13g2_decap_4 FILLER_12_561 ();
 sg13g2_fill_2 FILLER_12_573 ();
 sg13g2_fill_1 FILLER_12_575 ();
 sg13g2_decap_4 FILLER_12_584 ();
 sg13g2_decap_4 FILLER_12_622 ();
 sg13g2_fill_2 FILLER_12_626 ();
 sg13g2_decap_4 FILLER_12_649 ();
 sg13g2_fill_1 FILLER_12_653 ();
 sg13g2_fill_2 FILLER_12_679 ();
 sg13g2_fill_1 FILLER_12_681 ();
 sg13g2_fill_2 FILLER_12_705 ();
 sg13g2_fill_1 FILLER_12_755 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_fill_1 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_830 ();
 sg13g2_fill_2 FILLER_12_837 ();
 sg13g2_decap_4 FILLER_12_856 ();
 sg13g2_fill_2 FILLER_12_860 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_24 ();
 sg13g2_fill_1 FILLER_13_70 ();
 sg13g2_decap_4 FILLER_13_83 ();
 sg13g2_fill_1 FILLER_13_87 ();
 sg13g2_fill_1 FILLER_13_93 ();
 sg13g2_decap_4 FILLER_13_128 ();
 sg13g2_decap_4 FILLER_13_144 ();
 sg13g2_fill_1 FILLER_13_148 ();
 sg13g2_decap_4 FILLER_13_155 ();
 sg13g2_fill_1 FILLER_13_159 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_fill_2 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_268 ();
 sg13g2_fill_1 FILLER_13_275 ();
 sg13g2_decap_4 FILLER_13_329 ();
 sg13g2_fill_2 FILLER_13_333 ();
 sg13g2_fill_1 FILLER_13_369 ();
 sg13g2_fill_1 FILLER_13_382 ();
 sg13g2_fill_2 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_415 ();
 sg13g2_fill_1 FILLER_13_417 ();
 sg13g2_decap_8 FILLER_13_432 ();
 sg13g2_fill_1 FILLER_13_439 ();
 sg13g2_decap_8 FILLER_13_457 ();
 sg13g2_fill_1 FILLER_13_464 ();
 sg13g2_fill_1 FILLER_13_482 ();
 sg13g2_decap_4 FILLER_13_507 ();
 sg13g2_fill_2 FILLER_13_511 ();
 sg13g2_fill_2 FILLER_13_521 ();
 sg13g2_fill_2 FILLER_13_577 ();
 sg13g2_fill_1 FILLER_13_587 ();
 sg13g2_decap_8 FILLER_13_604 ();
 sg13g2_decap_4 FILLER_13_611 ();
 sg13g2_decap_4 FILLER_13_631 ();
 sg13g2_fill_2 FILLER_13_635 ();
 sg13g2_decap_8 FILLER_13_675 ();
 sg13g2_fill_2 FILLER_13_682 ();
 sg13g2_decap_8 FILLER_13_689 ();
 sg13g2_decap_4 FILLER_13_696 ();
 sg13g2_fill_1 FILLER_13_700 ();
 sg13g2_fill_2 FILLER_13_718 ();
 sg13g2_fill_1 FILLER_13_720 ();
 sg13g2_decap_4 FILLER_13_739 ();
 sg13g2_fill_2 FILLER_13_760 ();
 sg13g2_fill_2 FILLER_13_775 ();
 sg13g2_fill_1 FILLER_13_777 ();
 sg13g2_decap_4 FILLER_13_782 ();
 sg13g2_fill_2 FILLER_13_860 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_4 ();
 sg13g2_decap_8 FILLER_14_45 ();
 sg13g2_fill_2 FILLER_14_52 ();
 sg13g2_fill_2 FILLER_14_83 ();
 sg13g2_fill_1 FILLER_14_85 ();
 sg13g2_decap_8 FILLER_14_103 ();
 sg13g2_fill_2 FILLER_14_110 ();
 sg13g2_fill_2 FILLER_14_134 ();
 sg13g2_fill_2 FILLER_14_148 ();
 sg13g2_fill_1 FILLER_14_150 ();
 sg13g2_decap_4 FILLER_14_157 ();
 sg13g2_fill_1 FILLER_14_161 ();
 sg13g2_decap_4 FILLER_14_185 ();
 sg13g2_decap_4 FILLER_14_195 ();
 sg13g2_fill_1 FILLER_14_199 ();
 sg13g2_fill_1 FILLER_14_223 ();
 sg13g2_fill_2 FILLER_14_236 ();
 sg13g2_fill_1 FILLER_14_238 ();
 sg13g2_fill_2 FILLER_14_257 ();
 sg13g2_fill_1 FILLER_14_259 ();
 sg13g2_fill_2 FILLER_14_285 ();
 sg13g2_fill_2 FILLER_14_295 ();
 sg13g2_fill_1 FILLER_14_297 ();
 sg13g2_fill_1 FILLER_14_308 ();
 sg13g2_decap_4 FILLER_14_326 ();
 sg13g2_fill_2 FILLER_14_330 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_fill_1 FILLER_14_347 ();
 sg13g2_fill_1 FILLER_14_365 ();
 sg13g2_fill_2 FILLER_14_384 ();
 sg13g2_fill_1 FILLER_14_386 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_1 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_14_429 ();
 sg13g2_decap_4 FILLER_14_436 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_4 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_fill_2 FILLER_14_483 ();
 sg13g2_decap_4 FILLER_14_505 ();
 sg13g2_fill_1 FILLER_14_509 ();
 sg13g2_decap_4 FILLER_14_535 ();
 sg13g2_fill_1 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_570 ();
 sg13g2_decap_4 FILLER_14_603 ();
 sg13g2_fill_2 FILLER_14_607 ();
 sg13g2_fill_2 FILLER_14_654 ();
 sg13g2_decap_8 FILLER_14_662 ();
 sg13g2_fill_2 FILLER_14_669 ();
 sg13g2_decap_4 FILLER_14_690 ();
 sg13g2_decap_8 FILLER_14_716 ();
 sg13g2_fill_2 FILLER_14_765 ();
 sg13g2_fill_1 FILLER_14_767 ();
 sg13g2_fill_2 FILLER_14_785 ();
 sg13g2_fill_1 FILLER_14_811 ();
 sg13g2_decap_4 FILLER_14_829 ();
 sg13g2_fill_1 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_851 ();
 sg13g2_decap_4 FILLER_14_858 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_4 ();
 sg13g2_decap_4 FILLER_15_23 ();
 sg13g2_fill_2 FILLER_15_27 ();
 sg13g2_decap_4 FILLER_15_46 ();
 sg13g2_fill_1 FILLER_15_50 ();
 sg13g2_decap_4 FILLER_15_55 ();
 sg13g2_fill_1 FILLER_15_83 ();
 sg13g2_fill_1 FILLER_15_90 ();
 sg13g2_decap_8 FILLER_15_103 ();
 sg13g2_fill_2 FILLER_15_155 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_1 FILLER_15_176 ();
 sg13g2_fill_1 FILLER_15_183 ();
 sg13g2_fill_2 FILLER_15_196 ();
 sg13g2_fill_1 FILLER_15_250 ();
 sg13g2_fill_1 FILLER_15_276 ();
 sg13g2_fill_2 FILLER_15_293 ();
 sg13g2_fill_1 FILLER_15_295 ();
 sg13g2_fill_2 FILLER_15_316 ();
 sg13g2_decap_4 FILLER_15_348 ();
 sg13g2_fill_2 FILLER_15_352 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_fill_2 FILLER_15_434 ();
 sg13g2_fill_1 FILLER_15_460 ();
 sg13g2_decap_8 FILLER_15_478 ();
 sg13g2_fill_2 FILLER_15_485 ();
 sg13g2_fill_1 FILLER_15_493 ();
 sg13g2_decap_4 FILLER_15_508 ();
 sg13g2_fill_1 FILLER_15_512 ();
 sg13g2_fill_1 FILLER_15_521 ();
 sg13g2_fill_1 FILLER_15_539 ();
 sg13g2_decap_4 FILLER_15_546 ();
 sg13g2_fill_2 FILLER_15_602 ();
 sg13g2_fill_1 FILLER_15_604 ();
 sg13g2_decap_8 FILLER_15_622 ();
 sg13g2_decap_4 FILLER_15_629 ();
 sg13g2_decap_4 FILLER_15_655 ();
 sg13g2_fill_1 FILLER_15_664 ();
 sg13g2_decap_8 FILLER_15_696 ();
 sg13g2_fill_1 FILLER_15_703 ();
 sg13g2_fill_1 FILLER_15_729 ();
 sg13g2_fill_2 FILLER_15_744 ();
 sg13g2_fill_1 FILLER_15_746 ();
 sg13g2_fill_2 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_fill_1 FILLER_15_777 ();
 sg13g2_fill_2 FILLER_15_808 ();
 sg13g2_fill_1 FILLER_15_810 ();
 sg13g2_decap_4 FILLER_15_828 ();
 sg13g2_fill_1 FILLER_15_832 ();
 sg13g2_decap_8 FILLER_15_850 ();
 sg13g2_decap_4 FILLER_15_857 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_23 ();
 sg13g2_fill_1 FILLER_16_30 ();
 sg13g2_fill_1 FILLER_16_82 ();
 sg13g2_decap_4 FILLER_16_109 ();
 sg13g2_fill_2 FILLER_16_113 ();
 sg13g2_decap_8 FILLER_16_132 ();
 sg13g2_decap_4 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_143 ();
 sg13g2_decap_4 FILLER_16_149 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_decap_4 FILLER_16_194 ();
 sg13g2_fill_1 FILLER_16_202 ();
 sg13g2_fill_2 FILLER_16_220 ();
 sg13g2_fill_1 FILLER_16_222 ();
 sg13g2_fill_2 FILLER_16_239 ();
 sg13g2_fill_2 FILLER_16_258 ();
 sg13g2_decap_4 FILLER_16_294 ();
 sg13g2_decap_4 FILLER_16_376 ();
 sg13g2_fill_2 FILLER_16_384 ();
 sg13g2_fill_1 FILLER_16_386 ();
 sg13g2_fill_1 FILLER_16_412 ();
 sg13g2_decap_8 FILLER_16_426 ();
 sg13g2_decap_8 FILLER_16_433 ();
 sg13g2_decap_4 FILLER_16_440 ();
 sg13g2_fill_2 FILLER_16_444 ();
 sg13g2_decap_4 FILLER_16_462 ();
 sg13g2_fill_1 FILLER_16_466 ();
 sg13g2_decap_8 FILLER_16_506 ();
 sg13g2_fill_1 FILLER_16_521 ();
 sg13g2_decap_8 FILLER_16_573 ();
 sg13g2_fill_1 FILLER_16_580 ();
 sg13g2_decap_4 FILLER_16_597 ();
 sg13g2_fill_2 FILLER_16_618 ();
 sg13g2_fill_1 FILLER_16_620 ();
 sg13g2_fill_1 FILLER_16_638 ();
 sg13g2_fill_2 FILLER_16_645 ();
 sg13g2_decap_4 FILLER_16_694 ();
 sg13g2_fill_1 FILLER_16_698 ();
 sg13g2_fill_1 FILLER_16_712 ();
 sg13g2_fill_2 FILLER_16_719 ();
 sg13g2_fill_1 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_726 ();
 sg13g2_fill_1 FILLER_16_733 ();
 sg13g2_decap_4 FILLER_16_755 ();
 sg13g2_fill_2 FILLER_16_776 ();
 sg13g2_fill_2 FILLER_16_807 ();
 sg13g2_decap_8 FILLER_16_843 ();
 sg13g2_decap_8 FILLER_16_850 ();
 sg13g2_decap_4 FILLER_16_857 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_4 ();
 sg13g2_decap_8 FILLER_17_23 ();
 sg13g2_fill_1 FILLER_17_30 ();
 sg13g2_decap_8 FILLER_17_48 ();
 sg13g2_decap_4 FILLER_17_55 ();
 sg13g2_fill_1 FILLER_17_76 ();
 sg13g2_decap_8 FILLER_17_102 ();
 sg13g2_decap_4 FILLER_17_126 ();
 sg13g2_fill_2 FILLER_17_130 ();
 sg13g2_fill_1 FILLER_17_138 ();
 sg13g2_fill_2 FILLER_17_156 ();
 sg13g2_fill_1 FILLER_17_158 ();
 sg13g2_decap_4 FILLER_17_185 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_208 ();
 sg13g2_decap_4 FILLER_17_215 ();
 sg13g2_decap_4 FILLER_17_236 ();
 sg13g2_fill_2 FILLER_17_257 ();
 sg13g2_decap_8 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_fill_2 FILLER_17_290 ();
 sg13g2_fill_1 FILLER_17_292 ();
 sg13g2_decap_4 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_341 ();
 sg13g2_decap_4 FILLER_17_348 ();
 sg13g2_fill_2 FILLER_17_352 ();
 sg13g2_fill_2 FILLER_17_371 ();
 sg13g2_fill_1 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_fill_2 FILLER_17_387 ();
 sg13g2_fill_1 FILLER_17_406 ();
 sg13g2_fill_2 FILLER_17_412 ();
 sg13g2_fill_1 FILLER_17_414 ();
 sg13g2_decap_4 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_442 ();
 sg13g2_decap_4 FILLER_17_461 ();
 sg13g2_fill_2 FILLER_17_465 ();
 sg13g2_decap_8 FILLER_17_475 ();
 sg13g2_decap_8 FILLER_17_510 ();
 sg13g2_decap_8 FILLER_17_530 ();
 sg13g2_decap_4 FILLER_17_537 ();
 sg13g2_fill_2 FILLER_17_541 ();
 sg13g2_decap_8 FILLER_17_559 ();
 sg13g2_decap_8 FILLER_17_566 ();
 sg13g2_fill_2 FILLER_17_573 ();
 sg13g2_fill_2 FILLER_17_599 ();
 sg13g2_fill_1 FILLER_17_617 ();
 sg13g2_fill_2 FILLER_17_635 ();
 sg13g2_decap_4 FILLER_17_654 ();
 sg13g2_decap_4 FILLER_17_663 ();
 sg13g2_fill_2 FILLER_17_667 ();
 sg13g2_fill_2 FILLER_17_700 ();
 sg13g2_fill_1 FILLER_17_702 ();
 sg13g2_fill_1 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_745 ();
 sg13g2_decap_8 FILLER_17_752 ();
 sg13g2_fill_1 FILLER_17_759 ();
 sg13g2_fill_2 FILLER_17_777 ();
 sg13g2_fill_1 FILLER_17_783 ();
 sg13g2_fill_2 FILLER_17_792 ();
 sg13g2_fill_2 FILLER_17_800 ();
 sg13g2_fill_1 FILLER_17_802 ();
 sg13g2_decap_8 FILLER_17_820 ();
 sg13g2_decap_8 FILLER_17_827 ();
 sg13g2_decap_8 FILLER_17_834 ();
 sg13g2_decap_8 FILLER_17_841 ();
 sg13g2_decap_8 FILLER_17_848 ();
 sg13g2_decap_8 FILLER_17_855 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_24 ();
 sg13g2_fill_1 FILLER_18_31 ();
 sg13g2_fill_2 FILLER_18_49 ();
 sg13g2_decap_4 FILLER_18_85 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_decap_8 FILLER_18_99 ();
 sg13g2_decap_4 FILLER_18_106 ();
 sg13g2_fill_2 FILLER_18_139 ();
 sg13g2_decap_4 FILLER_18_159 ();
 sg13g2_fill_2 FILLER_18_163 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_fill_1 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_238 ();
 sg13g2_fill_1 FILLER_18_240 ();
 sg13g2_fill_2 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_285 ();
 sg13g2_fill_2 FILLER_18_306 ();
 sg13g2_fill_1 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_317 ();
 sg13g2_decap_4 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_352 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_decap_4 FILLER_18_372 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_decap_4 FILLER_18_394 ();
 sg13g2_fill_2 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_418 ();
 sg13g2_decap_4 FILLER_18_439 ();
 sg13g2_fill_1 FILLER_18_443 ();
 sg13g2_fill_2 FILLER_18_461 ();
 sg13g2_fill_2 FILLER_18_480 ();
 sg13g2_fill_2 FILLER_18_496 ();
 sg13g2_fill_1 FILLER_18_498 ();
 sg13g2_decap_4 FILLER_18_513 ();
 sg13g2_fill_2 FILLER_18_517 ();
 sg13g2_fill_2 FILLER_18_524 ();
 sg13g2_fill_1 FILLER_18_526 ();
 sg13g2_fill_2 FILLER_18_606 ();
 sg13g2_decap_8 FILLER_18_624 ();
 sg13g2_fill_2 FILLER_18_681 ();
 sg13g2_fill_1 FILLER_18_683 ();
 sg13g2_decap_8 FILLER_18_701 ();
 sg13g2_decap_8 FILLER_18_708 ();
 sg13g2_fill_1 FILLER_18_732 ();
 sg13g2_decap_8 FILLER_18_745 ();
 sg13g2_fill_2 FILLER_18_752 ();
 sg13g2_fill_1 FILLER_18_754 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_fill_2 FILLER_18_799 ();
 sg13g2_fill_1 FILLER_18_805 ();
 sg13g2_decap_4 FILLER_18_815 ();
 sg13g2_fill_1 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_2 ();
 sg13g2_decap_8 FILLER_19_20 ();
 sg13g2_decap_4 FILLER_19_27 ();
 sg13g2_decap_8 FILLER_19_48 ();
 sg13g2_fill_2 FILLER_19_85 ();
 sg13g2_decap_8 FILLER_19_104 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_fill_1 FILLER_19_129 ();
 sg13g2_decap_4 FILLER_19_152 ();
 sg13g2_fill_2 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_fill_2 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_219 ();
 sg13g2_decap_4 FILLER_19_228 ();
 sg13g2_fill_2 FILLER_19_240 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_fill_2 FILLER_19_262 ();
 sg13g2_fill_2 FILLER_19_269 ();
 sg13g2_fill_2 FILLER_19_275 ();
 sg13g2_fill_1 FILLER_19_277 ();
 sg13g2_fill_2 FILLER_19_295 ();
 sg13g2_fill_1 FILLER_19_305 ();
 sg13g2_fill_2 FILLER_19_324 ();
 sg13g2_decap_4 FILLER_19_343 ();
 sg13g2_fill_1 FILLER_19_347 ();
 sg13g2_fill_2 FILLER_19_365 ();
 sg13g2_fill_1 FILLER_19_367 ();
 sg13g2_fill_1 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_fill_1 FILLER_19_409 ();
 sg13g2_fill_2 FILLER_19_415 ();
 sg13g2_fill_1 FILLER_19_417 ();
 sg13g2_fill_1 FILLER_19_452 ();
 sg13g2_decap_8 FILLER_19_463 ();
 sg13g2_fill_2 FILLER_19_470 ();
 sg13g2_fill_1 FILLER_19_472 ();
 sg13g2_decap_4 FILLER_19_478 ();
 sg13g2_fill_1 FILLER_19_482 ();
 sg13g2_fill_2 FILLER_19_512 ();
 sg13g2_fill_1 FILLER_19_514 ();
 sg13g2_fill_1 FILLER_19_542 ();
 sg13g2_fill_2 FILLER_19_551 ();
 sg13g2_decap_8 FILLER_19_559 ();
 sg13g2_decap_4 FILLER_19_566 ();
 sg13g2_decap_4 FILLER_19_588 ();
 sg13g2_fill_2 FILLER_19_592 ();
 sg13g2_fill_1 FILLER_19_598 ();
 sg13g2_fill_2 FILLER_19_607 ();
 sg13g2_decap_4 FILLER_19_631 ();
 sg13g2_fill_1 FILLER_19_635 ();
 sg13g2_fill_2 FILLER_19_647 ();
 sg13g2_decap_8 FILLER_19_657 ();
 sg13g2_decap_8 FILLER_19_664 ();
 sg13g2_decap_4 FILLER_19_671 ();
 sg13g2_decap_8 FILLER_19_690 ();
 sg13g2_decap_8 FILLER_19_720 ();
 sg13g2_fill_2 FILLER_19_727 ();
 sg13g2_fill_1 FILLER_19_741 ();
 sg13g2_fill_1 FILLER_19_775 ();
 sg13g2_fill_1 FILLER_19_797 ();
 sg13g2_decap_8 FILLER_19_829 ();
 sg13g2_decap_8 FILLER_19_836 ();
 sg13g2_decap_8 FILLER_19_843 ();
 sg13g2_decap_8 FILLER_19_850 ();
 sg13g2_decap_4 FILLER_19_857 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_decap_4 FILLER_20_23 ();
 sg13g2_fill_1 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_50 ();
 sg13g2_decap_4 FILLER_20_57 ();
 sg13g2_fill_1 FILLER_20_61 ();
 sg13g2_fill_2 FILLER_20_88 ();
 sg13g2_fill_1 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_108 ();
 sg13g2_decap_8 FILLER_20_115 ();
 sg13g2_fill_1 FILLER_20_156 ();
 sg13g2_fill_1 FILLER_20_179 ();
 sg13g2_decap_4 FILLER_20_197 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_223 ();
 sg13g2_fill_2 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_233 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_decap_8 FILLER_20_268 ();
 sg13g2_fill_2 FILLER_20_283 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_decap_4 FILLER_20_325 ();
 sg13g2_fill_1 FILLER_20_329 ();
 sg13g2_decap_4 FILLER_20_347 ();
 sg13g2_fill_1 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_1 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_423 ();
 sg13g2_fill_1 FILLER_20_428 ();
 sg13g2_fill_2 FILLER_20_441 ();
 sg13g2_fill_1 FILLER_20_443 ();
 sg13g2_fill_2 FILLER_20_450 ();
 sg13g2_fill_1 FILLER_20_463 ();
 sg13g2_fill_2 FILLER_20_468 ();
 sg13g2_decap_8 FILLER_20_513 ();
 sg13g2_decap_4 FILLER_20_520 ();
 sg13g2_fill_2 FILLER_20_524 ();
 sg13g2_decap_4 FILLER_20_535 ();
 sg13g2_fill_2 FILLER_20_539 ();
 sg13g2_fill_1 FILLER_20_569 ();
 sg13g2_decap_8 FILLER_20_578 ();
 sg13g2_fill_2 FILLER_20_615 ();
 sg13g2_fill_2 FILLER_20_646 ();
 sg13g2_fill_1 FILLER_20_648 ();
 sg13g2_fill_1 FILLER_20_661 ();
 sg13g2_fill_2 FILLER_20_670 ();
 sg13g2_fill_1 FILLER_20_698 ();
 sg13g2_fill_1 FILLER_20_707 ();
 sg13g2_fill_1 FILLER_20_750 ();
 sg13g2_fill_2 FILLER_20_765 ();
 sg13g2_fill_1 FILLER_20_767 ();
 sg13g2_fill_2 FILLER_20_780 ();
 sg13g2_fill_2 FILLER_20_796 ();
 sg13g2_fill_1 FILLER_20_798 ();
 sg13g2_fill_1 FILLER_20_830 ();
 sg13g2_decap_8 FILLER_20_836 ();
 sg13g2_decap_8 FILLER_20_843 ();
 sg13g2_decap_8 FILLER_20_850 ();
 sg13g2_decap_4 FILLER_20_857 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_12 ();
 sg13g2_decap_4 FILLER_21_19 ();
 sg13g2_fill_1 FILLER_21_23 ();
 sg13g2_decap_4 FILLER_21_40 ();
 sg13g2_fill_2 FILLER_21_68 ();
 sg13g2_decap_4 FILLER_21_104 ();
 sg13g2_fill_2 FILLER_21_108 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_fill_2 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_162 ();
 sg13g2_fill_2 FILLER_21_170 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_201 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_fill_2 FILLER_21_224 ();
 sg13g2_fill_2 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_fill_2 FILLER_21_279 ();
 sg13g2_fill_2 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_322 ();
 sg13g2_decap_4 FILLER_21_362 ();
 sg13g2_fill_1 FILLER_21_366 ();
 sg13g2_fill_1 FILLER_21_385 ();
 sg13g2_fill_2 FILLER_21_418 ();
 sg13g2_fill_2 FILLER_21_432 ();
 sg13g2_fill_1 FILLER_21_434 ();
 sg13g2_fill_1 FILLER_21_466 ();
 sg13g2_fill_2 FILLER_21_493 ();
 sg13g2_fill_2 FILLER_21_504 ();
 sg13g2_fill_1 FILLER_21_550 ();
 sg13g2_fill_1 FILLER_21_586 ();
 sg13g2_fill_1 FILLER_21_611 ();
 sg13g2_fill_2 FILLER_21_625 ();
 sg13g2_fill_2 FILLER_21_645 ();
 sg13g2_fill_1 FILLER_21_647 ();
 sg13g2_fill_1 FILLER_21_656 ();
 sg13g2_decap_4 FILLER_21_669 ();
 sg13g2_fill_2 FILLER_21_673 ();
 sg13g2_decap_4 FILLER_21_680 ();
 sg13g2_fill_1 FILLER_21_692 ();
 sg13g2_fill_2 FILLER_21_708 ();
 sg13g2_fill_1 FILLER_21_710 ();
 sg13g2_decap_4 FILLER_21_769 ();
 sg13g2_fill_2 FILLER_21_808 ();
 sg13g2_decap_8 FILLER_21_845 ();
 sg13g2_decap_8 FILLER_21_852 ();
 sg13g2_fill_2 FILLER_21_859 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_69 ();
 sg13g2_fill_1 FILLER_22_75 ();
 sg13g2_decap_4 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_114 ();
 sg13g2_decap_8 FILLER_22_123 ();
 sg13g2_decap_8 FILLER_22_130 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_fill_2 FILLER_22_155 ();
 sg13g2_fill_1 FILLER_22_157 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_4 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_192 ();
 sg13g2_fill_1 FILLER_22_194 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_fill_2 FILLER_22_272 ();
 sg13g2_fill_1 FILLER_22_285 ();
 sg13g2_fill_2 FILLER_22_298 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_307 ();
 sg13g2_fill_2 FILLER_22_326 ();
 sg13g2_fill_1 FILLER_22_328 ();
 sg13g2_decap_4 FILLER_22_346 ();
 sg13g2_decap_4 FILLER_22_367 ();
 sg13g2_fill_1 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_4 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_410 ();
 sg13g2_fill_2 FILLER_22_421 ();
 sg13g2_fill_1 FILLER_22_423 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_fill_2 FILLER_22_453 ();
 sg13g2_fill_1 FILLER_22_455 ();
 sg13g2_fill_2 FILLER_22_466 ();
 sg13g2_fill_1 FILLER_22_468 ();
 sg13g2_fill_2 FILLER_22_474 ();
 sg13g2_fill_1 FILLER_22_476 ();
 sg13g2_fill_2 FILLER_22_572 ();
 sg13g2_fill_2 FILLER_22_583 ();
 sg13g2_fill_1 FILLER_22_585 ();
 sg13g2_decap_4 FILLER_22_590 ();
 sg13g2_fill_2 FILLER_22_594 ();
 sg13g2_decap_8 FILLER_22_600 ();
 sg13g2_decap_4 FILLER_22_607 ();
 sg13g2_fill_2 FILLER_22_611 ();
 sg13g2_fill_2 FILLER_22_659 ();
 sg13g2_fill_1 FILLER_22_661 ();
 sg13g2_fill_1 FILLER_22_697 ();
 sg13g2_decap_8 FILLER_22_724 ();
 sg13g2_fill_1 FILLER_22_731 ();
 sg13g2_decap_8 FILLER_22_740 ();
 sg13g2_decap_4 FILLER_22_747 ();
 sg13g2_fill_1 FILLER_22_751 ();
 sg13g2_decap_8 FILLER_22_757 ();
 sg13g2_fill_2 FILLER_22_764 ();
 sg13g2_fill_2 FILLER_22_775 ();
 sg13g2_fill_1 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_822 ();
 sg13g2_decap_8 FILLER_22_829 ();
 sg13g2_decap_8 FILLER_22_836 ();
 sg13g2_decap_8 FILLER_22_843 ();
 sg13g2_decap_8 FILLER_22_850 ();
 sg13g2_decap_4 FILLER_22_857 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_27 ();
 sg13g2_decap_4 FILLER_23_34 ();
 sg13g2_fill_1 FILLER_23_38 ();
 sg13g2_fill_1 FILLER_23_48 ();
 sg13g2_fill_2 FILLER_23_79 ();
 sg13g2_decap_8 FILLER_23_114 ();
 sg13g2_fill_1 FILLER_23_137 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_1 FILLER_23_221 ();
 sg13g2_fill_1 FILLER_23_236 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_317 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_fill_2 FILLER_23_335 ();
 sg13g2_fill_1 FILLER_23_337 ();
 sg13g2_fill_2 FILLER_23_364 ();
 sg13g2_fill_2 FILLER_23_388 ();
 sg13g2_fill_1 FILLER_23_390 ();
 sg13g2_fill_2 FILLER_23_416 ();
 sg13g2_fill_1 FILLER_23_418 ();
 sg13g2_fill_2 FILLER_23_458 ();
 sg13g2_fill_2 FILLER_23_501 ();
 sg13g2_decap_4 FILLER_23_507 ();
 sg13g2_fill_1 FILLER_23_567 ();
 sg13g2_fill_2 FILLER_23_573 ();
 sg13g2_fill_1 FILLER_23_605 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_fill_2 FILLER_23_639 ();
 sg13g2_fill_2 FILLER_23_658 ();
 sg13g2_fill_2 FILLER_23_685 ();
 sg13g2_fill_1 FILLER_23_687 ();
 sg13g2_fill_2 FILLER_23_693 ();
 sg13g2_fill_1 FILLER_23_695 ();
 sg13g2_fill_1 FILLER_23_707 ();
 sg13g2_fill_2 FILLER_23_747 ();
 sg13g2_fill_1 FILLER_23_775 ();
 sg13g2_decap_8 FILLER_23_829 ();
 sg13g2_decap_8 FILLER_23_836 ();
 sg13g2_decap_8 FILLER_23_843 ();
 sg13g2_decap_8 FILLER_23_850 ();
 sg13g2_decap_4 FILLER_23_857 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_fill_2 FILLER_24_17 ();
 sg13g2_fill_1 FILLER_24_44 ();
 sg13g2_fill_2 FILLER_24_76 ();
 sg13g2_fill_2 FILLER_24_85 ();
 sg13g2_decap_8 FILLER_24_113 ();
 sg13g2_fill_2 FILLER_24_120 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_fill_1 FILLER_24_156 ();
 sg13g2_fill_2 FILLER_24_179 ();
 sg13g2_fill_1 FILLER_24_181 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_321 ();
 sg13g2_decap_8 FILLER_24_344 ();
 sg13g2_fill_2 FILLER_24_351 ();
 sg13g2_fill_2 FILLER_24_370 ();
 sg13g2_fill_2 FILLER_24_388 ();
 sg13g2_fill_2 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_430 ();
 sg13g2_decap_8 FILLER_24_437 ();
 sg13g2_decap_4 FILLER_24_444 ();
 sg13g2_fill_2 FILLER_24_448 ();
 sg13g2_fill_2 FILLER_24_460 ();
 sg13g2_decap_4 FILLER_24_475 ();
 sg13g2_fill_2 FILLER_24_479 ();
 sg13g2_decap_4 FILLER_24_495 ();
 sg13g2_fill_2 FILLER_24_573 ();
 sg13g2_fill_1 FILLER_24_575 ();
 sg13g2_fill_1 FILLER_24_633 ();
 sg13g2_fill_1 FILLER_24_673 ();
 sg13g2_fill_1 FILLER_24_690 ();
 sg13g2_fill_1 FILLER_24_718 ();
 sg13g2_fill_1 FILLER_24_727 ();
 sg13g2_decap_8 FILLER_24_736 ();
 sg13g2_fill_2 FILLER_24_743 ();
 sg13g2_fill_1 FILLER_24_745 ();
 sg13g2_fill_1 FILLER_24_826 ();
 sg13g2_decap_4 FILLER_24_857 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_66 ();
 sg13g2_fill_1 FILLER_25_120 ();
 sg13g2_fill_2 FILLER_25_137 ();
 sg13g2_fill_2 FILLER_25_165 ();
 sg13g2_decap_8 FILLER_25_192 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_243 ();
 sg13g2_fill_2 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_fill_2 FILLER_25_306 ();
 sg13g2_fill_1 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_318 ();
 sg13g2_fill_2 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_331 ();
 sg13g2_fill_1 FILLER_25_364 ();
 sg13g2_fill_1 FILLER_25_391 ();
 sg13g2_fill_1 FILLER_25_418 ();
 sg13g2_decap_8 FILLER_25_426 ();
 sg13g2_fill_2 FILLER_25_433 ();
 sg13g2_fill_1 FILLER_25_435 ();
 sg13g2_decap_4 FILLER_25_472 ();
 sg13g2_fill_2 FILLER_25_476 ();
 sg13g2_fill_1 FILLER_25_508 ();
 sg13g2_fill_2 FILLER_25_533 ();
 sg13g2_fill_2 FILLER_25_541 ();
 sg13g2_fill_2 FILLER_25_561 ();
 sg13g2_fill_1 FILLER_25_563 ();
 sg13g2_fill_2 FILLER_25_577 ();
 sg13g2_fill_1 FILLER_25_704 ();
 sg13g2_fill_2 FILLER_25_715 ();
 sg13g2_fill_2 FILLER_25_766 ();
 sg13g2_fill_1 FILLER_25_786 ();
 sg13g2_fill_2 FILLER_25_804 ();
 sg13g2_fill_1 FILLER_25_821 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_fill_2 FILLER_26_41 ();
 sg13g2_fill_2 FILLER_26_59 ();
 sg13g2_fill_1 FILLER_26_67 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_79 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_decap_4 FILLER_26_109 ();
 sg13g2_fill_2 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_162 ();
 sg13g2_decap_8 FILLER_26_185 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_fill_2 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_271 ();
 sg13g2_fill_1 FILLER_26_273 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_decap_4 FILLER_26_355 ();
 sg13g2_fill_1 FILLER_26_391 ();
 sg13g2_fill_2 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_432 ();
 sg13g2_fill_2 FILLER_26_466 ();
 sg13g2_fill_1 FILLER_26_468 ();
 sg13g2_fill_2 FILLER_26_509 ();
 sg13g2_fill_1 FILLER_26_528 ();
 sg13g2_fill_2 FILLER_26_563 ();
 sg13g2_fill_1 FILLER_26_565 ();
 sg13g2_fill_1 FILLER_26_614 ();
 sg13g2_decap_4 FILLER_26_667 ();
 sg13g2_fill_2 FILLER_26_696 ();
 sg13g2_decap_4 FILLER_26_724 ();
 sg13g2_fill_2 FILLER_26_728 ();
 sg13g2_fill_1 FILLER_26_782 ();
 sg13g2_fill_2 FILLER_26_808 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_10 ();
 sg13g2_fill_2 FILLER_27_83 ();
 sg13g2_fill_2 FILLER_27_111 ();
 sg13g2_fill_1 FILLER_27_172 ();
 sg13g2_fill_1 FILLER_27_204 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_268 ();
 sg13g2_decap_8 FILLER_27_274 ();
 sg13g2_decap_4 FILLER_27_281 ();
 sg13g2_fill_2 FILLER_27_349 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_fill_2 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_411 ();
 sg13g2_fill_1 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_419 ();
 sg13g2_decap_8 FILLER_27_426 ();
 sg13g2_fill_1 FILLER_27_453 ();
 sg13g2_fill_2 FILLER_27_530 ();
 sg13g2_fill_1 FILLER_27_564 ();
 sg13g2_fill_2 FILLER_27_594 ();
 sg13g2_fill_2 FILLER_27_633 ();
 sg13g2_fill_1 FILLER_27_635 ();
 sg13g2_fill_2 FILLER_27_641 ();
 sg13g2_fill_1 FILLER_27_643 ();
 sg13g2_fill_2 FILLER_27_689 ();
 sg13g2_fill_1 FILLER_27_691 ();
 sg13g2_decap_4 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_720 ();
 sg13g2_fill_2 FILLER_27_727 ();
 sg13g2_decap_4 FILLER_27_742 ();
 sg13g2_fill_2 FILLER_27_746 ();
 sg13g2_fill_2 FILLER_27_761 ();
 sg13g2_fill_2 FILLER_27_777 ();
 sg13g2_fill_1 FILLER_27_779 ();
 sg13g2_fill_2 FILLER_27_803 ();
 sg13g2_fill_2 FILLER_27_829 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_36 ();
 sg13g2_fill_1 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_fill_2 FILLER_28_108 ();
 sg13g2_fill_2 FILLER_28_135 ();
 sg13g2_fill_2 FILLER_28_155 ();
 sg13g2_fill_1 FILLER_28_182 ();
 sg13g2_fill_2 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_decap_4 FILLER_28_270 ();
 sg13g2_fill_2 FILLER_28_274 ();
 sg13g2_fill_2 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_289 ();
 sg13g2_fill_1 FILLER_28_296 ();
 sg13g2_fill_1 FILLER_28_305 ();
 sg13g2_fill_2 FILLER_28_314 ();
 sg13g2_decap_4 FILLER_28_352 ();
 sg13g2_fill_2 FILLER_28_365 ();
 sg13g2_decap_4 FILLER_28_410 ();
 sg13g2_decap_8 FILLER_28_424 ();
 sg13g2_fill_2 FILLER_28_431 ();
 sg13g2_fill_1 FILLER_28_433 ();
 sg13g2_fill_1 FILLER_28_479 ();
 sg13g2_fill_1 FILLER_28_499 ();
 sg13g2_fill_2 FILLER_28_545 ();
 sg13g2_fill_1 FILLER_28_547 ();
 sg13g2_fill_1 FILLER_28_569 ();
 sg13g2_fill_2 FILLER_28_586 ();
 sg13g2_decap_4 FILLER_28_616 ();
 sg13g2_fill_1 FILLER_28_620 ();
 sg13g2_decap_8 FILLER_28_629 ();
 sg13g2_fill_2 FILLER_28_667 ();
 sg13g2_fill_1 FILLER_28_669 ();
 sg13g2_fill_2 FILLER_28_675 ();
 sg13g2_fill_1 FILLER_28_677 ();
 sg13g2_decap_4 FILLER_28_687 ();
 sg13g2_fill_2 FILLER_28_691 ();
 sg13g2_fill_2 FILLER_28_744 ();
 sg13g2_fill_1 FILLER_28_746 ();
 sg13g2_fill_2 FILLER_28_777 ();
 sg13g2_decap_4 FILLER_28_836 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_34 ();
 sg13g2_fill_1 FILLER_29_62 ();
 sg13g2_fill_2 FILLER_29_144 ();
 sg13g2_fill_1 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_152 ();
 sg13g2_fill_1 FILLER_29_154 ();
 sg13g2_decap_4 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_fill_2 FILLER_29_191 ();
 sg13g2_fill_1 FILLER_29_193 ();
 sg13g2_fill_2 FILLER_29_218 ();
 sg13g2_fill_2 FILLER_29_245 ();
 sg13g2_fill_2 FILLER_29_255 ();
 sg13g2_decap_4 FILLER_29_288 ();
 sg13g2_fill_2 FILLER_29_292 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_fill_2 FILLER_29_388 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_fill_2 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_407 ();
 sg13g2_fill_2 FILLER_29_419 ();
 sg13g2_decap_4 FILLER_29_429 ();
 sg13g2_fill_2 FILLER_29_433 ();
 sg13g2_fill_2 FILLER_29_445 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_fill_2 FILLER_29_469 ();
 sg13g2_fill_2 FILLER_29_482 ();
 sg13g2_fill_1 FILLER_29_484 ();
 sg13g2_fill_2 FILLER_29_559 ();
 sg13g2_fill_1 FILLER_29_569 ();
 sg13g2_fill_1 FILLER_29_575 ();
 sg13g2_decap_8 FILLER_29_591 ();
 sg13g2_fill_2 FILLER_29_598 ();
 sg13g2_fill_1 FILLER_29_609 ();
 sg13g2_fill_2 FILLER_29_614 ();
 sg13g2_fill_2 FILLER_29_621 ();
 sg13g2_decap_8 FILLER_29_636 ();
 sg13g2_fill_1 FILLER_29_648 ();
 sg13g2_fill_2 FILLER_29_659 ();
 sg13g2_decap_8 FILLER_29_698 ();
 sg13g2_decap_8 FILLER_29_705 ();
 sg13g2_fill_2 FILLER_29_721 ();
 sg13g2_fill_1 FILLER_29_723 ();
 sg13g2_fill_2 FILLER_29_740 ();
 sg13g2_fill_1 FILLER_29_742 ();
 sg13g2_fill_2 FILLER_29_751 ();
 sg13g2_fill_1 FILLER_29_753 ();
 sg13g2_fill_1 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_768 ();
 sg13g2_decap_4 FILLER_29_775 ();
 sg13g2_fill_1 FILLER_29_779 ();
 sg13g2_fill_2 FILLER_29_796 ();
 sg13g2_fill_1 FILLER_29_828 ();
 sg13g2_fill_2 FILLER_29_833 ();
 sg13g2_fill_1 FILLER_29_835 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_fill_1 FILLER_30_53 ();
 sg13g2_fill_1 FILLER_30_113 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_145 ();
 sg13g2_fill_2 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_182 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_decap_4 FILLER_30_257 ();
 sg13g2_decap_8 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_276 ();
 sg13g2_fill_2 FILLER_30_282 ();
 sg13g2_decap_4 FILLER_30_289 ();
 sg13g2_fill_2 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_30_323 ();
 sg13g2_fill_2 FILLER_30_357 ();
 sg13g2_fill_2 FILLER_30_371 ();
 sg13g2_fill_2 FILLER_30_378 ();
 sg13g2_fill_1 FILLER_30_380 ();
 sg13g2_fill_2 FILLER_30_404 ();
 sg13g2_decap_4 FILLER_30_437 ();
 sg13g2_fill_2 FILLER_30_441 ();
 sg13g2_decap_4 FILLER_30_453 ();
 sg13g2_decap_4 FILLER_30_465 ();
 sg13g2_fill_2 FILLER_30_519 ();
 sg13g2_fill_1 FILLER_30_521 ();
 sg13g2_decap_8 FILLER_30_555 ();
 sg13g2_fill_2 FILLER_30_589 ();
 sg13g2_fill_1 FILLER_30_615 ();
 sg13g2_fill_2 FILLER_30_621 ();
 sg13g2_fill_2 FILLER_30_647 ();
 sg13g2_fill_1 FILLER_30_649 ();
 sg13g2_fill_2 FILLER_30_667 ();
 sg13g2_fill_1 FILLER_30_669 ();
 sg13g2_fill_1 FILLER_30_723 ();
 sg13g2_fill_2 FILLER_30_730 ();
 sg13g2_fill_2 FILLER_30_743 ();
 sg13g2_decap_8 FILLER_30_769 ();
 sg13g2_fill_1 FILLER_30_796 ();
 sg13g2_fill_1 FILLER_30_834 ();
 sg13g2_fill_2 FILLER_30_840 ();
 sg13g2_fill_1 FILLER_30_842 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_150 ();
 sg13g2_fill_2 FILLER_31_183 ();
 sg13g2_fill_1 FILLER_31_185 ();
 sg13g2_decap_4 FILLER_31_255 ();
 sg13g2_fill_2 FILLER_31_267 ();
 sg13g2_fill_2 FILLER_31_295 ();
 sg13g2_fill_1 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_302 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_4 FILLER_31_331 ();
 sg13g2_fill_1 FILLER_31_335 ();
 sg13g2_fill_2 FILLER_31_361 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_31_412 ();
 sg13g2_decap_8 FILLER_31_427 ();
 sg13g2_fill_2 FILLER_31_462 ();
 sg13g2_fill_1 FILLER_31_482 ();
 sg13g2_fill_1 FILLER_31_509 ();
 sg13g2_fill_2 FILLER_31_519 ();
 sg13g2_fill_1 FILLER_31_545 ();
 sg13g2_decap_8 FILLER_31_551 ();
 sg13g2_decap_8 FILLER_31_558 ();
 sg13g2_decap_8 FILLER_31_588 ();
 sg13g2_fill_1 FILLER_31_595 ();
 sg13g2_fill_1 FILLER_31_601 ();
 sg13g2_fill_1 FILLER_31_613 ();
 sg13g2_fill_2 FILLER_31_618 ();
 sg13g2_fill_2 FILLER_31_639 ();
 sg13g2_fill_2 FILLER_31_669 ();
 sg13g2_fill_1 FILLER_31_671 ();
 sg13g2_decap_8 FILLER_31_688 ();
 sg13g2_fill_2 FILLER_31_695 ();
 sg13g2_fill_1 FILLER_31_697 ();
 sg13g2_decap_8 FILLER_31_708 ();
 sg13g2_decap_8 FILLER_31_715 ();
 sg13g2_fill_2 FILLER_31_722 ();
 sg13g2_decap_4 FILLER_31_745 ();
 sg13g2_decap_4 FILLER_31_774 ();
 sg13g2_fill_2 FILLER_31_778 ();
 sg13g2_fill_2 FILLER_31_796 ();
 sg13g2_fill_1 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_821 ();
 sg13g2_decap_4 FILLER_31_828 ();
 sg13g2_fill_1 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_94 ();
 sg13g2_fill_1 FILLER_32_96 ();
 sg13g2_fill_1 FILLER_32_123 ();
 sg13g2_fill_2 FILLER_32_168 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_206 ();
 sg13g2_decap_4 FILLER_32_221 ();
 sg13g2_fill_2 FILLER_32_225 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_fill_1 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_267 ();
 sg13g2_fill_1 FILLER_32_269 ();
 sg13g2_decap_8 FILLER_32_286 ();
 sg13g2_fill_2 FILLER_32_293 ();
 sg13g2_fill_1 FILLER_32_304 ();
 sg13g2_decap_4 FILLER_32_333 ();
 sg13g2_fill_2 FILLER_32_337 ();
 sg13g2_decap_4 FILLER_32_355 ();
 sg13g2_fill_2 FILLER_32_359 ();
 sg13g2_fill_2 FILLER_32_369 ();
 sg13g2_fill_1 FILLER_32_381 ();
 sg13g2_fill_1 FILLER_32_398 ();
 sg13g2_fill_1 FILLER_32_431 ();
 sg13g2_decap_8 FILLER_32_460 ();
 sg13g2_fill_2 FILLER_32_467 ();
 sg13g2_fill_1 FILLER_32_469 ();
 sg13g2_fill_2 FILLER_32_478 ();
 sg13g2_decap_4 FILLER_32_531 ();
 sg13g2_fill_2 FILLER_32_547 ();
 sg13g2_fill_1 FILLER_32_549 ();
 sg13g2_fill_1 FILLER_32_558 ();
 sg13g2_fill_2 FILLER_32_579 ();
 sg13g2_fill_2 FILLER_32_593 ();
 sg13g2_fill_1 FILLER_32_595 ();
 sg13g2_fill_2 FILLER_32_600 ();
 sg13g2_fill_1 FILLER_32_602 ();
 sg13g2_fill_2 FILLER_32_609 ();
 sg13g2_fill_1 FILLER_32_632 ();
 sg13g2_fill_2 FILLER_32_650 ();
 sg13g2_fill_2 FILLER_32_657 ();
 sg13g2_fill_1 FILLER_32_659 ();
 sg13g2_fill_2 FILLER_32_665 ();
 sg13g2_fill_1 FILLER_32_667 ();
 sg13g2_fill_2 FILLER_32_699 ();
 sg13g2_fill_2 FILLER_32_741 ();
 sg13g2_fill_1 FILLER_32_743 ();
 sg13g2_fill_1 FILLER_32_753 ();
 sg13g2_fill_2 FILLER_32_768 ();
 sg13g2_fill_1 FILLER_32_806 ();
 sg13g2_fill_2 FILLER_32_827 ();
 sg13g2_fill_1 FILLER_32_843 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_32 ();
 sg13g2_fill_2 FILLER_33_72 ();
 sg13g2_fill_1 FILLER_33_87 ();
 sg13g2_fill_1 FILLER_33_114 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_fill_2 FILLER_33_214 ();
 sg13g2_fill_1 FILLER_33_216 ();
 sg13g2_decap_8 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_244 ();
 sg13g2_fill_1 FILLER_33_246 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_fill_1 FILLER_33_311 ();
 sg13g2_decap_4 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_354 ();
 sg13g2_fill_1 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_382 ();
 sg13g2_fill_1 FILLER_33_384 ();
 sg13g2_fill_2 FILLER_33_400 ();
 sg13g2_decap_4 FILLER_33_407 ();
 sg13g2_fill_2 FILLER_33_411 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_decap_4 FILLER_33_429 ();
 sg13g2_fill_1 FILLER_33_433 ();
 sg13g2_fill_1 FILLER_33_444 ();
 sg13g2_fill_2 FILLER_33_460 ();
 sg13g2_fill_2 FILLER_33_472 ();
 sg13g2_fill_1 FILLER_33_474 ();
 sg13g2_fill_1 FILLER_33_493 ();
 sg13g2_fill_2 FILLER_33_503 ();
 sg13g2_fill_2 FILLER_33_561 ();
 sg13g2_fill_2 FILLER_33_567 ();
 sg13g2_decap_8 FILLER_33_580 ();
 sg13g2_fill_1 FILLER_33_587 ();
 sg13g2_fill_2 FILLER_33_598 ();
 sg13g2_fill_1 FILLER_33_604 ();
 sg13g2_fill_2 FILLER_33_648 ();
 sg13g2_fill_1 FILLER_33_650 ();
 sg13g2_fill_2 FILLER_33_670 ();
 sg13g2_fill_1 FILLER_33_672 ();
 sg13g2_decap_4 FILLER_33_697 ();
 sg13g2_fill_2 FILLER_33_701 ();
 sg13g2_fill_2 FILLER_33_716 ();
 sg13g2_fill_1 FILLER_33_718 ();
 sg13g2_fill_1 FILLER_33_724 ();
 sg13g2_fill_2 FILLER_33_741 ();
 sg13g2_fill_1 FILLER_33_743 ();
 sg13g2_fill_1 FILLER_33_753 ();
 sg13g2_fill_2 FILLER_33_769 ();
 sg13g2_fill_2 FILLER_33_790 ();
 sg13g2_decap_4 FILLER_33_805 ();
 sg13g2_decap_4 FILLER_33_822 ();
 sg13g2_fill_1 FILLER_33_826 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_27 ();
 sg13g2_fill_1 FILLER_34_37 ();
 sg13g2_fill_2 FILLER_34_174 ();
 sg13g2_fill_2 FILLER_34_181 ();
 sg13g2_decap_8 FILLER_34_193 ();
 sg13g2_decap_4 FILLER_34_200 ();
 sg13g2_decap_4 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_decap_4 FILLER_34_238 ();
 sg13g2_fill_1 FILLER_34_242 ();
 sg13g2_fill_2 FILLER_34_269 ();
 sg13g2_fill_2 FILLER_34_331 ();
 sg13g2_fill_2 FILLER_34_338 ();
 sg13g2_fill_1 FILLER_34_340 ();
 sg13g2_decap_4 FILLER_34_375 ();
 sg13g2_fill_2 FILLER_34_395 ();
 sg13g2_fill_1 FILLER_34_397 ();
 sg13g2_fill_2 FILLER_34_403 ();
 sg13g2_fill_1 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_34_424 ();
 sg13g2_fill_2 FILLER_34_431 ();
 sg13g2_fill_2 FILLER_34_443 ();
 sg13g2_fill_1 FILLER_34_537 ();
 sg13g2_decap_8 FILLER_34_554 ();
 sg13g2_fill_1 FILLER_34_570 ();
 sg13g2_fill_2 FILLER_34_581 ();
 sg13g2_decap_8 FILLER_34_587 ();
 sg13g2_fill_2 FILLER_34_594 ();
 sg13g2_fill_1 FILLER_34_624 ();
 sg13g2_fill_2 FILLER_34_629 ();
 sg13g2_fill_1 FILLER_34_644 ();
 sg13g2_fill_1 FILLER_34_650 ();
 sg13g2_fill_2 FILLER_34_658 ();
 sg13g2_decap_4 FILLER_34_668 ();
 sg13g2_fill_1 FILLER_34_672 ();
 sg13g2_decap_4 FILLER_34_699 ();
 sg13g2_fill_2 FILLER_34_703 ();
 sg13g2_fill_2 FILLER_34_717 ();
 sg13g2_fill_2 FILLER_34_724 ();
 sg13g2_fill_1 FILLER_34_726 ();
 sg13g2_fill_1 FILLER_34_731 ();
 sg13g2_fill_2 FILLER_34_752 ();
 sg13g2_decap_8 FILLER_34_787 ();
 sg13g2_decap_4 FILLER_34_794 ();
 sg13g2_decap_4 FILLER_34_829 ();
 sg13g2_decap_4 FILLER_34_844 ();
 sg13g2_decap_4 FILLER_34_858 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_48 ();
 sg13g2_fill_2 FILLER_35_92 ();
 sg13g2_fill_1 FILLER_35_146 ();
 sg13g2_fill_2 FILLER_35_202 ();
 sg13g2_fill_1 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_248 ();
 sg13g2_fill_2 FILLER_35_254 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_fill_1 FILLER_35_281 ();
 sg13g2_fill_2 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_305 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_fill_2 FILLER_35_349 ();
 sg13g2_fill_2 FILLER_35_381 ();
 sg13g2_fill_2 FILLER_35_416 ();
 sg13g2_decap_8 FILLER_35_423 ();
 sg13g2_decap_4 FILLER_35_434 ();
 sg13g2_fill_2 FILLER_35_443 ();
 sg13g2_fill_1 FILLER_35_445 ();
 sg13g2_fill_1 FILLER_35_456 ();
 sg13g2_fill_2 FILLER_35_475 ();
 sg13g2_fill_2 FILLER_35_518 ();
 sg13g2_fill_2 FILLER_35_525 ();
 sg13g2_fill_1 FILLER_35_537 ();
 sg13g2_fill_2 FILLER_35_555 ();
 sg13g2_fill_1 FILLER_35_595 ();
 sg13g2_fill_1 FILLER_35_614 ();
 sg13g2_fill_1 FILLER_35_639 ();
 sg13g2_fill_2 FILLER_35_645 ();
 sg13g2_fill_1 FILLER_35_647 ();
 sg13g2_fill_1 FILLER_35_656 ();
 sg13g2_decap_4 FILLER_35_677 ();
 sg13g2_fill_1 FILLER_35_681 ();
 sg13g2_fill_2 FILLER_35_687 ();
 sg13g2_fill_1 FILLER_35_689 ();
 sg13g2_decap_8 FILLER_35_696 ();
 sg13g2_fill_1 FILLER_35_703 ();
 sg13g2_fill_2 FILLER_35_732 ();
 sg13g2_decap_8 FILLER_35_744 ();
 sg13g2_fill_2 FILLER_35_755 ();
 sg13g2_fill_1 FILLER_35_757 ();
 sg13g2_fill_2 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_796 ();
 sg13g2_fill_2 FILLER_35_803 ();
 sg13g2_fill_1 FILLER_35_829 ();
 sg13g2_fill_2 FILLER_36_25 ();
 sg13g2_fill_1 FILLER_36_46 ();
 sg13g2_fill_2 FILLER_36_52 ();
 sg13g2_fill_2 FILLER_36_66 ();
 sg13g2_fill_1 FILLER_36_82 ();
 sg13g2_fill_1 FILLER_36_115 ();
 sg13g2_fill_2 FILLER_36_129 ();
 sg13g2_fill_1 FILLER_36_143 ();
 sg13g2_fill_2 FILLER_36_174 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_decap_4 FILLER_36_234 ();
 sg13g2_fill_2 FILLER_36_316 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_fill_2 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_decap_8 FILLER_36_361 ();
 sg13g2_decap_4 FILLER_36_368 ();
 sg13g2_fill_1 FILLER_36_372 ();
 sg13g2_fill_1 FILLER_36_413 ();
 sg13g2_fill_1 FILLER_36_419 ();
 sg13g2_fill_2 FILLER_36_446 ();
 sg13g2_fill_1 FILLER_36_448 ();
 sg13g2_fill_1 FILLER_36_528 ();
 sg13g2_decap_8 FILLER_36_550 ();
 sg13g2_fill_2 FILLER_36_562 ();
 sg13g2_decap_4 FILLER_36_587 ();
 sg13g2_fill_1 FILLER_36_596 ();
 sg13g2_decap_8 FILLER_36_611 ();
 sg13g2_decap_8 FILLER_36_618 ();
 sg13g2_decap_4 FILLER_36_625 ();
 sg13g2_fill_2 FILLER_36_629 ();
 sg13g2_fill_2 FILLER_36_637 ();
 sg13g2_fill_1 FILLER_36_639 ();
 sg13g2_decap_4 FILLER_36_671 ();
 sg13g2_fill_2 FILLER_36_675 ();
 sg13g2_decap_4 FILLER_36_685 ();
 sg13g2_fill_2 FILLER_36_689 ();
 sg13g2_fill_2 FILLER_36_697 ();
 sg13g2_fill_1 FILLER_36_699 ();
 sg13g2_fill_2 FILLER_36_715 ();
 sg13g2_decap_4 FILLER_36_737 ();
 sg13g2_fill_2 FILLER_36_754 ();
 sg13g2_fill_1 FILLER_36_756 ();
 sg13g2_decap_4 FILLER_36_771 ();
 sg13g2_fill_1 FILLER_36_775 ();
 sg13g2_fill_1 FILLER_36_784 ();
 sg13g2_fill_2 FILLER_36_817 ();
 sg13g2_decap_4 FILLER_36_829 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_65 ();
 sg13g2_fill_2 FILLER_37_86 ();
 sg13g2_fill_1 FILLER_37_123 ();
 sg13g2_fill_1 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_160 ();
 sg13g2_fill_1 FILLER_37_179 ();
 sg13g2_fill_2 FILLER_37_207 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_fill_2 FILLER_37_215 ();
 sg13g2_fill_1 FILLER_37_222 ();
 sg13g2_decap_4 FILLER_37_236 ();
 sg13g2_fill_2 FILLER_37_245 ();
 sg13g2_fill_1 FILLER_37_247 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_decap_8 FILLER_37_288 ();
 sg13g2_fill_2 FILLER_37_295 ();
 sg13g2_fill_1 FILLER_37_297 ();
 sg13g2_decap_4 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_306 ();
 sg13g2_fill_2 FILLER_37_321 ();
 sg13g2_fill_1 FILLER_37_329 ();
 sg13g2_fill_2 FILLER_37_335 ();
 sg13g2_fill_1 FILLER_37_337 ();
 sg13g2_decap_4 FILLER_37_387 ();
 sg13g2_fill_2 FILLER_37_412 ();
 sg13g2_fill_2 FILLER_37_418 ();
 sg13g2_decap_4 FILLER_37_436 ();
 sg13g2_decap_4 FILLER_37_445 ();
 sg13g2_fill_2 FILLER_37_514 ();
 sg13g2_fill_2 FILLER_37_524 ();
 sg13g2_fill_1 FILLER_37_551 ();
 sg13g2_fill_2 FILLER_37_565 ();
 sg13g2_fill_1 FILLER_37_567 ();
 sg13g2_decap_4 FILLER_37_584 ();
 sg13g2_fill_1 FILLER_37_588 ();
 sg13g2_decap_4 FILLER_37_615 ();
 sg13g2_fill_2 FILLER_37_619 ();
 sg13g2_fill_2 FILLER_37_634 ();
 sg13g2_fill_2 FILLER_37_640 ();
 sg13g2_fill_1 FILLER_37_642 ();
 sg13g2_fill_2 FILLER_37_648 ();
 sg13g2_fill_1 FILLER_37_650 ();
 sg13g2_fill_1 FILLER_37_733 ();
 sg13g2_fill_2 FILLER_37_740 ();
 sg13g2_fill_2 FILLER_37_747 ();
 sg13g2_fill_1 FILLER_37_776 ();
 sg13g2_fill_2 FILLER_37_806 ();
 sg13g2_fill_2 FILLER_37_834 ();
 sg13g2_decap_4 FILLER_37_858 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_62 ();
 sg13g2_fill_1 FILLER_38_68 ();
 sg13g2_fill_2 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_117 ();
 sg13g2_fill_2 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_134 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_fill_1 FILLER_38_162 ();
 sg13g2_fill_2 FILLER_38_185 ();
 sg13g2_fill_1 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_198 ();
 sg13g2_fill_1 FILLER_38_200 ();
 sg13g2_fill_1 FILLER_38_205 ();
 sg13g2_fill_2 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_246 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_254 ();
 sg13g2_fill_2 FILLER_38_277 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_2 FILLER_38_284 ();
 sg13g2_fill_1 FILLER_38_290 ();
 sg13g2_decap_8 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_fill_1 FILLER_38_371 ();
 sg13g2_fill_1 FILLER_38_376 ();
 sg13g2_decap_4 FILLER_38_398 ();
 sg13g2_fill_1 FILLER_38_402 ();
 sg13g2_fill_1 FILLER_38_449 ();
 sg13g2_fill_1 FILLER_38_473 ();
 sg13g2_fill_1 FILLER_38_503 ();
 sg13g2_fill_1 FILLER_38_535 ();
 sg13g2_decap_8 FILLER_38_544 ();
 sg13g2_fill_2 FILLER_38_551 ();
 sg13g2_decap_8 FILLER_38_561 ();
 sg13g2_decap_4 FILLER_38_568 ();
 sg13g2_fill_2 FILLER_38_572 ();
 sg13g2_decap_4 FILLER_38_579 ();
 sg13g2_fill_2 FILLER_38_588 ();
 sg13g2_fill_1 FILLER_38_590 ();
 sg13g2_fill_2 FILLER_38_620 ();
 sg13g2_decap_4 FILLER_38_643 ();
 sg13g2_fill_1 FILLER_38_647 ();
 sg13g2_fill_1 FILLER_38_657 ();
 sg13g2_decap_4 FILLER_38_674 ();
 sg13g2_fill_2 FILLER_38_678 ();
 sg13g2_decap_8 FILLER_38_684 ();
 sg13g2_decap_4 FILLER_38_691 ();
 sg13g2_fill_1 FILLER_38_707 ();
 sg13g2_decap_8 FILLER_38_726 ();
 sg13g2_fill_2 FILLER_38_733 ();
 sg13g2_fill_2 FILLER_38_740 ();
 sg13g2_fill_1 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_747 ();
 sg13g2_fill_2 FILLER_38_754 ();
 sg13g2_fill_1 FILLER_38_761 ();
 sg13g2_fill_2 FILLER_38_784 ();
 sg13g2_fill_2 FILLER_38_805 ();
 sg13g2_fill_1 FILLER_38_807 ();
 sg13g2_fill_1 FILLER_38_827 ();
 sg13g2_fill_1 FILLER_38_836 ();
 sg13g2_fill_2 FILLER_38_845 ();
 sg13g2_fill_1 FILLER_38_847 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_fill_2 FILLER_39_52 ();
 sg13g2_fill_1 FILLER_39_88 ();
 sg13g2_fill_2 FILLER_39_191 ();
 sg13g2_decap_8 FILLER_39_212 ();
 sg13g2_fill_2 FILLER_39_219 ();
 sg13g2_decap_8 FILLER_39_234 ();
 sg13g2_fill_2 FILLER_39_241 ();
 sg13g2_fill_1 FILLER_39_243 ();
 sg13g2_decap_4 FILLER_39_312 ();
 sg13g2_fill_2 FILLER_39_316 ();
 sg13g2_fill_2 FILLER_39_344 ();
 sg13g2_decap_4 FILLER_39_365 ();
 sg13g2_fill_1 FILLER_39_369 ();
 sg13g2_fill_1 FILLER_39_374 ();
 sg13g2_fill_2 FILLER_39_386 ();
 sg13g2_fill_2 FILLER_39_405 ();
 sg13g2_fill_1 FILLER_39_407 ();
 sg13g2_fill_1 FILLER_39_430 ();
 sg13g2_decap_4 FILLER_39_539 ();
 sg13g2_fill_2 FILLER_39_543 ();
 sg13g2_fill_2 FILLER_39_550 ();
 sg13g2_fill_1 FILLER_39_591 ();
 sg13g2_fill_2 FILLER_39_615 ();
 sg13g2_fill_1 FILLER_39_617 ();
 sg13g2_decap_4 FILLER_39_626 ();
 sg13g2_decap_4 FILLER_39_673 ();
 sg13g2_fill_2 FILLER_39_677 ();
 sg13g2_decap_4 FILLER_39_684 ();
 sg13g2_fill_2 FILLER_39_712 ();
 sg13g2_decap_4 FILLER_39_733 ();
 sg13g2_fill_1 FILLER_39_737 ();
 sg13g2_fill_2 FILLER_39_763 ();
 sg13g2_fill_1 FILLER_39_765 ();
 sg13g2_decap_4 FILLER_39_776 ();
 sg13g2_decap_4 FILLER_39_793 ();
 sg13g2_fill_2 FILLER_39_797 ();
 sg13g2_fill_1 FILLER_39_823 ();
 sg13g2_fill_2 FILLER_39_832 ();
 sg13g2_fill_2 FILLER_39_848 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_37 ();
 sg13g2_fill_2 FILLER_40_69 ();
 sg13g2_fill_1 FILLER_40_149 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_fill_2 FILLER_40_175 ();
 sg13g2_fill_2 FILLER_40_182 ();
 sg13g2_fill_1 FILLER_40_194 ();
 sg13g2_fill_2 FILLER_40_216 ();
 sg13g2_fill_1 FILLER_40_218 ();
 sg13g2_decap_8 FILLER_40_242 ();
 sg13g2_fill_2 FILLER_40_249 ();
 sg13g2_fill_1 FILLER_40_279 ();
 sg13g2_fill_2 FILLER_40_285 ();
 sg13g2_fill_1 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_305 ();
 sg13g2_fill_2 FILLER_40_312 ();
 sg13g2_decap_8 FILLER_40_325 ();
 sg13g2_decap_4 FILLER_40_332 ();
 sg13g2_fill_2 FILLER_40_336 ();
 sg13g2_fill_2 FILLER_40_343 ();
 sg13g2_fill_1 FILLER_40_360 ();
 sg13g2_fill_2 FILLER_40_373 ();
 sg13g2_fill_1 FILLER_40_375 ();
 sg13g2_decap_4 FILLER_40_394 ();
 sg13g2_fill_1 FILLER_40_398 ();
 sg13g2_fill_2 FILLER_40_436 ();
 sg13g2_fill_2 FILLER_40_450 ();
 sg13g2_fill_1 FILLER_40_452 ();
 sg13g2_decap_8 FILLER_40_558 ();
 sg13g2_fill_1 FILLER_40_565 ();
 sg13g2_decap_4 FILLER_40_574 ();
 sg13g2_fill_1 FILLER_40_586 ();
 sg13g2_decap_4 FILLER_40_591 ();
 sg13g2_fill_2 FILLER_40_595 ();
 sg13g2_decap_4 FILLER_40_601 ();
 sg13g2_fill_1 FILLER_40_605 ();
 sg13g2_fill_1 FILLER_40_622 ();
 sg13g2_decap_4 FILLER_40_645 ();
 sg13g2_fill_2 FILLER_40_649 ();
 sg13g2_fill_1 FILLER_40_674 ();
 sg13g2_decap_4 FILLER_40_679 ();
 sg13g2_fill_1 FILLER_40_700 ();
 sg13g2_decap_8 FILLER_40_723 ();
 sg13g2_decap_8 FILLER_40_730 ();
 sg13g2_fill_1 FILLER_40_737 ();
 sg13g2_fill_2 FILLER_40_781 ();
 sg13g2_decap_4 FILLER_40_796 ();
 sg13g2_fill_1 FILLER_40_800 ();
 sg13g2_fill_2 FILLER_40_807 ();
 sg13g2_decap_8 FILLER_40_813 ();
 sg13g2_fill_2 FILLER_40_850 ();
 sg13g2_fill_1 FILLER_40_852 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_42 ();
 sg13g2_fill_1 FILLER_41_52 ();
 sg13g2_fill_1 FILLER_41_93 ();
 sg13g2_fill_2 FILLER_41_157 ();
 sg13g2_fill_1 FILLER_41_171 ();
 sg13g2_fill_1 FILLER_41_190 ();
 sg13g2_fill_2 FILLER_41_196 ();
 sg13g2_fill_1 FILLER_41_198 ();
 sg13g2_decap_4 FILLER_41_250 ();
 sg13g2_fill_1 FILLER_41_254 ();
 sg13g2_fill_2 FILLER_41_298 ();
 sg13g2_fill_1 FILLER_41_300 ();
 sg13g2_fill_1 FILLER_41_309 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_fill_1 FILLER_41_362 ();
 sg13g2_fill_1 FILLER_41_369 ();
 sg13g2_decap_4 FILLER_41_398 ();
 sg13g2_fill_2 FILLER_41_402 ();
 sg13g2_fill_1 FILLER_41_409 ();
 sg13g2_fill_1 FILLER_41_424 ();
 sg13g2_fill_1 FILLER_41_434 ();
 sg13g2_fill_1 FILLER_41_453 ();
 sg13g2_fill_1 FILLER_41_500 ();
 sg13g2_decap_8 FILLER_41_517 ();
 sg13g2_fill_1 FILLER_41_536 ();
 sg13g2_fill_1 FILLER_41_550 ();
 sg13g2_decap_8 FILLER_41_556 ();
 sg13g2_decap_8 FILLER_41_563 ();
 sg13g2_fill_2 FILLER_41_584 ();
 sg13g2_fill_1 FILLER_41_592 ();
 sg13g2_decap_8 FILLER_41_598 ();
 sg13g2_decap_4 FILLER_41_621 ();
 sg13g2_decap_8 FILLER_41_649 ();
 sg13g2_fill_2 FILLER_41_656 ();
 sg13g2_fill_1 FILLER_41_658 ();
 sg13g2_fill_2 FILLER_41_671 ();
 sg13g2_fill_1 FILLER_41_702 ();
 sg13g2_fill_2 FILLER_41_716 ();
 sg13g2_decap_8 FILLER_41_752 ();
 sg13g2_fill_1 FILLER_41_759 ();
 sg13g2_fill_2 FILLER_41_764 ();
 sg13g2_fill_1 FILLER_41_766 ();
 sg13g2_fill_2 FILLER_41_780 ();
 sg13g2_fill_1 FILLER_41_792 ();
 sg13g2_fill_2 FILLER_41_827 ();
 sg13g2_fill_1 FILLER_41_834 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_fill_1 FILLER_42_35 ();
 sg13g2_fill_2 FILLER_42_95 ();
 sg13g2_decap_4 FILLER_42_127 ();
 sg13g2_fill_2 FILLER_42_149 ();
 sg13g2_fill_2 FILLER_42_162 ();
 sg13g2_fill_1 FILLER_42_174 ();
 sg13g2_decap_4 FILLER_42_179 ();
 sg13g2_fill_1 FILLER_42_183 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_fill_1 FILLER_42_214 ();
 sg13g2_fill_1 FILLER_42_230 ();
 sg13g2_decap_4 FILLER_42_241 ();
 sg13g2_fill_2 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_270 ();
 sg13g2_fill_1 FILLER_42_277 ();
 sg13g2_fill_1 FILLER_42_292 ();
 sg13g2_decap_8 FILLER_42_325 ();
 sg13g2_decap_8 FILLER_42_332 ();
 sg13g2_fill_2 FILLER_42_339 ();
 sg13g2_fill_1 FILLER_42_341 ();
 sg13g2_decap_4 FILLER_42_402 ();
 sg13g2_fill_1 FILLER_42_406 ();
 sg13g2_fill_2 FILLER_42_419 ();
 sg13g2_decap_8 FILLER_42_437 ();
 sg13g2_decap_8 FILLER_42_444 ();
 sg13g2_decap_4 FILLER_42_451 ();
 sg13g2_fill_1 FILLER_42_490 ();
 sg13g2_decap_8 FILLER_42_508 ();
 sg13g2_decap_4 FILLER_42_542 ();
 sg13g2_fill_2 FILLER_42_546 ();
 sg13g2_fill_2 FILLER_42_558 ();
 sg13g2_fill_1 FILLER_42_560 ();
 sg13g2_fill_2 FILLER_42_569 ();
 sg13g2_fill_1 FILLER_42_585 ();
 sg13g2_decap_8 FILLER_42_600 ();
 sg13g2_fill_2 FILLER_42_607 ();
 sg13g2_decap_4 FILLER_42_626 ();
 sg13g2_fill_2 FILLER_42_630 ();
 sg13g2_fill_1 FILLER_42_637 ();
 sg13g2_decap_4 FILLER_42_643 ();
 sg13g2_fill_2 FILLER_42_647 ();
 sg13g2_fill_1 FILLER_42_680 ();
 sg13g2_fill_2 FILLER_42_695 ();
 sg13g2_decap_8 FILLER_42_703 ();
 sg13g2_fill_2 FILLER_42_710 ();
 sg13g2_fill_2 FILLER_42_716 ();
 sg13g2_decap_8 FILLER_42_728 ();
 sg13g2_decap_8 FILLER_42_739 ();
 sg13g2_fill_2 FILLER_42_746 ();
 sg13g2_decap_4 FILLER_42_759 ();
 sg13g2_fill_2 FILLER_42_763 ();
 sg13g2_fill_2 FILLER_42_795 ();
 sg13g2_fill_1 FILLER_42_797 ();
 sg13g2_decap_4 FILLER_42_808 ();
 sg13g2_fill_2 FILLER_42_812 ();
 sg13g2_decap_8 FILLER_42_850 ();
 sg13g2_decap_4 FILLER_42_857 ();
 sg13g2_fill_1 FILLER_42_861 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_72 ();
 sg13g2_fill_1 FILLER_43_74 ();
 sg13g2_fill_1 FILLER_43_80 ();
 sg13g2_fill_2 FILLER_43_115 ();
 sg13g2_fill_2 FILLER_43_151 ();
 sg13g2_fill_2 FILLER_43_171 ();
 sg13g2_fill_1 FILLER_43_173 ();
 sg13g2_fill_2 FILLER_43_179 ();
 sg13g2_fill_1 FILLER_43_181 ();
 sg13g2_fill_1 FILLER_43_194 ();
 sg13g2_fill_1 FILLER_43_222 ();
 sg13g2_decap_4 FILLER_43_235 ();
 sg13g2_fill_1 FILLER_43_239 ();
 sg13g2_decap_8 FILLER_43_254 ();
 sg13g2_decap_4 FILLER_43_261 ();
 sg13g2_fill_1 FILLER_43_279 ();
 sg13g2_decap_4 FILLER_43_311 ();
 sg13g2_decap_4 FILLER_43_321 ();
 sg13g2_fill_2 FILLER_43_325 ();
 sg13g2_fill_1 FILLER_43_344 ();
 sg13g2_fill_2 FILLER_43_349 ();
 sg13g2_fill_1 FILLER_43_351 ();
 sg13g2_fill_1 FILLER_43_373 ();
 sg13g2_fill_2 FILLER_43_379 ();
 sg13g2_fill_1 FILLER_43_381 ();
 sg13g2_fill_2 FILLER_43_388 ();
 sg13g2_decap_4 FILLER_43_395 ();
 sg13g2_fill_1 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_404 ();
 sg13g2_fill_2 FILLER_43_411 ();
 sg13g2_fill_2 FILLER_43_426 ();
 sg13g2_fill_2 FILLER_43_436 ();
 sg13g2_fill_1 FILLER_43_447 ();
 sg13g2_decap_8 FILLER_43_452 ();
 sg13g2_fill_1 FILLER_43_459 ();
 sg13g2_fill_2 FILLER_43_465 ();
 sg13g2_fill_2 FILLER_43_485 ();
 sg13g2_fill_1 FILLER_43_487 ();
 sg13g2_fill_2 FILLER_43_551 ();
 sg13g2_fill_1 FILLER_43_553 ();
 sg13g2_fill_1 FILLER_43_573 ();
 sg13g2_decap_4 FILLER_43_590 ();
 sg13g2_decap_4 FILLER_43_602 ();
 sg13g2_decap_4 FILLER_43_653 ();
 sg13g2_fill_1 FILLER_43_657 ();
 sg13g2_decap_4 FILLER_43_668 ();
 sg13g2_fill_2 FILLER_43_672 ();
 sg13g2_decap_4 FILLER_43_691 ();
 sg13g2_fill_2 FILLER_43_695 ();
 sg13g2_fill_2 FILLER_43_722 ();
 sg13g2_decap_4 FILLER_43_737 ();
 sg13g2_fill_2 FILLER_43_763 ();
 sg13g2_fill_1 FILLER_43_773 ();
 sg13g2_decap_4 FILLER_43_780 ();
 sg13g2_fill_1 FILLER_43_800 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_58 ();
 sg13g2_fill_2 FILLER_44_116 ();
 sg13g2_fill_1 FILLER_44_172 ();
 sg13g2_fill_1 FILLER_44_178 ();
 sg13g2_fill_2 FILLER_44_191 ();
 sg13g2_fill_1 FILLER_44_193 ();
 sg13g2_fill_2 FILLER_44_204 ();
 sg13g2_fill_1 FILLER_44_206 ();
 sg13g2_fill_2 FILLER_44_212 ();
 sg13g2_fill_2 FILLER_44_229 ();
 sg13g2_fill_1 FILLER_44_241 ();
 sg13g2_fill_2 FILLER_44_268 ();
 sg13g2_fill_1 FILLER_44_270 ();
 sg13g2_fill_2 FILLER_44_281 ();
 sg13g2_fill_1 FILLER_44_283 ();
 sg13g2_fill_1 FILLER_44_327 ();
 sg13g2_fill_2 FILLER_44_344 ();
 sg13g2_fill_1 FILLER_44_346 ();
 sg13g2_fill_2 FILLER_44_357 ();
 sg13g2_fill_1 FILLER_44_359 ();
 sg13g2_decap_4 FILLER_44_371 ();
 sg13g2_decap_4 FILLER_44_380 ();
 sg13g2_fill_1 FILLER_44_389 ();
 sg13g2_decap_4 FILLER_44_399 ();
 sg13g2_fill_1 FILLER_44_403 ();
 sg13g2_fill_1 FILLER_44_409 ();
 sg13g2_decap_8 FILLER_44_436 ();
 sg13g2_fill_1 FILLER_44_443 ();
 sg13g2_fill_2 FILLER_44_449 ();
 sg13g2_fill_2 FILLER_44_468 ();
 sg13g2_decap_8 FILLER_44_475 ();
 sg13g2_fill_2 FILLER_44_482 ();
 sg13g2_fill_1 FILLER_44_484 ();
 sg13g2_fill_2 FILLER_44_529 ();
 sg13g2_fill_1 FILLER_44_531 ();
 sg13g2_fill_2 FILLER_44_544 ();
 sg13g2_fill_2 FILLER_44_553 ();
 sg13g2_fill_1 FILLER_44_570 ();
 sg13g2_fill_2 FILLER_44_577 ();
 sg13g2_fill_1 FILLER_44_579 ();
 sg13g2_fill_1 FILLER_44_584 ();
 sg13g2_decap_4 FILLER_44_595 ();
 sg13g2_fill_2 FILLER_44_599 ();
 sg13g2_fill_2 FILLER_44_606 ();
 sg13g2_fill_2 FILLER_44_618 ();
 sg13g2_decap_4 FILLER_44_625 ();
 sg13g2_fill_2 FILLER_44_629 ();
 sg13g2_decap_8 FILLER_44_647 ();
 sg13g2_decap_4 FILLER_44_654 ();
 sg13g2_fill_1 FILLER_44_658 ();
 sg13g2_fill_2 FILLER_44_663 ();
 sg13g2_fill_1 FILLER_44_665 ();
 sg13g2_decap_8 FILLER_44_674 ();
 sg13g2_fill_1 FILLER_44_690 ();
 sg13g2_fill_1 FILLER_44_707 ();
 sg13g2_fill_1 FILLER_44_721 ();
 sg13g2_fill_2 FILLER_44_730 ();
 sg13g2_fill_1 FILLER_44_732 ();
 sg13g2_fill_1 FILLER_44_743 ();
 sg13g2_decap_8 FILLER_44_758 ();
 sg13g2_decap_8 FILLER_44_765 ();
 sg13g2_fill_2 FILLER_44_772 ();
 sg13g2_decap_4 FILLER_44_780 ();
 sg13g2_fill_2 FILLER_44_788 ();
 sg13g2_fill_1 FILLER_44_790 ();
 sg13g2_decap_4 FILLER_44_799 ();
 sg13g2_fill_2 FILLER_44_803 ();
 sg13g2_decap_8 FILLER_44_810 ();
 sg13g2_fill_2 FILLER_44_827 ();
 sg13g2_fill_1 FILLER_44_829 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_fill_1 FILLER_45_29 ();
 sg13g2_fill_2 FILLER_45_71 ();
 sg13g2_fill_1 FILLER_45_73 ();
 sg13g2_fill_2 FILLER_45_96 ();
 sg13g2_fill_2 FILLER_45_102 ();
 sg13g2_fill_1 FILLER_45_108 ();
 sg13g2_fill_2 FILLER_45_123 ();
 sg13g2_fill_1 FILLER_45_129 ();
 sg13g2_fill_2 FILLER_45_167 ();
 sg13g2_fill_1 FILLER_45_169 ();
 sg13g2_fill_1 FILLER_45_192 ();
 sg13g2_fill_2 FILLER_45_198 ();
 sg13g2_fill_2 FILLER_45_205 ();
 sg13g2_fill_1 FILLER_45_207 ();
 sg13g2_fill_1 FILLER_45_226 ();
 sg13g2_fill_2 FILLER_45_240 ();
 sg13g2_fill_2 FILLER_45_275 ();
 sg13g2_decap_8 FILLER_45_330 ();
 sg13g2_fill_1 FILLER_45_337 ();
 sg13g2_fill_2 FILLER_45_352 ();
 sg13g2_fill_1 FILLER_45_354 ();
 sg13g2_fill_2 FILLER_45_366 ();
 sg13g2_fill_1 FILLER_45_368 ();
 sg13g2_fill_2 FILLER_45_384 ();
 sg13g2_fill_1 FILLER_45_391 ();
 sg13g2_decap_8 FILLER_45_398 ();
 sg13g2_decap_4 FILLER_45_405 ();
 sg13g2_fill_1 FILLER_45_409 ();
 sg13g2_fill_1 FILLER_45_431 ();
 sg13g2_decap_4 FILLER_45_457 ();
 sg13g2_fill_1 FILLER_45_461 ();
 sg13g2_fill_2 FILLER_45_467 ();
 sg13g2_fill_1 FILLER_45_469 ();
 sg13g2_decap_4 FILLER_45_488 ();
 sg13g2_fill_1 FILLER_45_492 ();
 sg13g2_decap_8 FILLER_45_509 ();
 sg13g2_fill_1 FILLER_45_516 ();
 sg13g2_fill_2 FILLER_45_528 ();
 sg13g2_fill_2 FILLER_45_535 ();
 sg13g2_decap_4 FILLER_45_582 ();
 sg13g2_fill_1 FILLER_45_586 ();
 sg13g2_fill_1 FILLER_45_604 ();
 sg13g2_decap_8 FILLER_45_623 ();
 sg13g2_fill_1 FILLER_45_630 ();
 sg13g2_fill_1 FILLER_45_649 ();
 sg13g2_fill_2 FILLER_45_672 ();
 sg13g2_fill_1 FILLER_45_674 ();
 sg13g2_fill_2 FILLER_45_684 ();
 sg13g2_fill_2 FILLER_45_727 ();
 sg13g2_fill_2 FILLER_45_740 ();
 sg13g2_fill_1 FILLER_45_742 ();
 sg13g2_decap_4 FILLER_45_755 ();
 sg13g2_fill_1 FILLER_45_759 ();
 sg13g2_fill_2 FILLER_45_765 ();
 sg13g2_fill_1 FILLER_45_767 ();
 sg13g2_decap_4 FILLER_45_789 ();
 sg13g2_fill_1 FILLER_45_793 ();
 sg13g2_decap_4 FILLER_45_823 ();
 sg13g2_fill_1 FILLER_45_827 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_fill_2 FILLER_46_85 ();
 sg13g2_fill_1 FILLER_46_87 ();
 sg13g2_fill_2 FILLER_46_96 ();
 sg13g2_fill_1 FILLER_46_107 ();
 sg13g2_fill_2 FILLER_46_123 ();
 sg13g2_fill_1 FILLER_46_138 ();
 sg13g2_fill_2 FILLER_46_156 ();
 sg13g2_fill_1 FILLER_46_169 ();
 sg13g2_fill_2 FILLER_46_190 ();
 sg13g2_fill_1 FILLER_46_197 ();
 sg13g2_fill_1 FILLER_46_206 ();
 sg13g2_fill_2 FILLER_46_226 ();
 sg13g2_fill_1 FILLER_46_228 ();
 sg13g2_fill_2 FILLER_46_313 ();
 sg13g2_fill_2 FILLER_46_336 ();
 sg13g2_fill_2 FILLER_46_346 ();
 sg13g2_fill_2 FILLER_46_364 ();
 sg13g2_fill_2 FILLER_46_374 ();
 sg13g2_fill_1 FILLER_46_376 ();
 sg13g2_fill_2 FILLER_46_449 ();
 sg13g2_fill_2 FILLER_46_476 ();
 sg13g2_fill_2 FILLER_46_492 ();
 sg13g2_decap_4 FILLER_46_500 ();
 sg13g2_fill_2 FILLER_46_504 ();
 sg13g2_fill_2 FILLER_46_562 ();
 sg13g2_fill_1 FILLER_46_564 ();
 sg13g2_decap_4 FILLER_46_596 ();
 sg13g2_decap_4 FILLER_46_623 ();
 sg13g2_fill_2 FILLER_46_627 ();
 sg13g2_fill_2 FILLER_46_645 ();
 sg13g2_fill_1 FILLER_46_647 ();
 sg13g2_fill_2 FILLER_46_653 ();
 sg13g2_decap_8 FILLER_46_702 ();
 sg13g2_fill_1 FILLER_46_709 ();
 sg13g2_decap_8 FILLER_46_715 ();
 sg13g2_fill_2 FILLER_46_722 ();
 sg13g2_fill_1 FILLER_46_724 ();
 sg13g2_decap_4 FILLER_46_735 ();
 sg13g2_fill_2 FILLER_46_749 ();
 sg13g2_fill_2 FILLER_46_768 ();
 sg13g2_fill_2 FILLER_46_781 ();
 sg13g2_fill_1 FILLER_46_783 ();
 sg13g2_fill_1 FILLER_46_806 ();
 sg13g2_fill_2 FILLER_46_827 ();
 sg13g2_fill_2 FILLER_46_834 ();
 sg13g2_fill_1 FILLER_46_836 ();
 sg13g2_decap_8 FILLER_46_853 ();
 sg13g2_fill_2 FILLER_46_860 ();
 sg13g2_fill_1 FILLER_47_31 ();
 sg13g2_fill_1 FILLER_47_55 ();
 sg13g2_fill_1 FILLER_47_70 ();
 sg13g2_fill_2 FILLER_47_110 ();
 sg13g2_fill_2 FILLER_47_116 ();
 sg13g2_fill_1 FILLER_47_118 ();
 sg13g2_fill_2 FILLER_47_150 ();
 sg13g2_fill_1 FILLER_47_183 ();
 sg13g2_fill_1 FILLER_47_190 ();
 sg13g2_fill_1 FILLER_47_202 ();
 sg13g2_fill_2 FILLER_47_240 ();
 sg13g2_fill_1 FILLER_47_276 ();
 sg13g2_fill_1 FILLER_47_287 ();
 sg13g2_decap_4 FILLER_47_314 ();
 sg13g2_fill_1 FILLER_47_324 ();
 sg13g2_fill_2 FILLER_47_330 ();
 sg13g2_fill_1 FILLER_47_340 ();
 sg13g2_fill_1 FILLER_47_371 ();
 sg13g2_fill_2 FILLER_47_383 ();
 sg13g2_fill_2 FILLER_47_411 ();
 sg13g2_fill_1 FILLER_47_413 ();
 sg13g2_fill_2 FILLER_47_423 ();
 sg13g2_fill_2 FILLER_47_457 ();
 sg13g2_fill_1 FILLER_47_459 ();
 sg13g2_fill_2 FILLER_47_471 ();
 sg13g2_fill_1 FILLER_47_473 ();
 sg13g2_fill_2 FILLER_47_510 ();
 sg13g2_fill_1 FILLER_47_512 ();
 sg13g2_decap_4 FILLER_47_526 ();
 sg13g2_fill_1 FILLER_47_530 ();
 sg13g2_fill_1 FILLER_47_543 ();
 sg13g2_fill_1 FILLER_47_552 ();
 sg13g2_fill_2 FILLER_47_582 ();
 sg13g2_fill_1 FILLER_47_584 ();
 sg13g2_decap_8 FILLER_47_590 ();
 sg13g2_fill_1 FILLER_47_597 ();
 sg13g2_fill_1 FILLER_47_613 ();
 sg13g2_decap_4 FILLER_47_641 ();
 sg13g2_fill_2 FILLER_47_668 ();
 sg13g2_fill_2 FILLER_47_703 ();
 sg13g2_fill_1 FILLER_47_753 ();
 sg13g2_fill_2 FILLER_47_766 ();
 sg13g2_fill_2 FILLER_47_777 ();
 sg13g2_fill_1 FILLER_47_779 ();
 sg13g2_fill_1 FILLER_47_791 ();
 sg13g2_fill_1 FILLER_47_811 ();
 sg13g2_fill_1 FILLER_47_832 ();
 sg13g2_fill_1 FILLER_48_40 ();
 sg13g2_fill_1 FILLER_48_81 ();
 sg13g2_fill_1 FILLER_48_96 ();
 sg13g2_fill_1 FILLER_48_123 ();
 sg13g2_fill_2 FILLER_48_206 ();
 sg13g2_fill_2 FILLER_48_221 ();
 sg13g2_fill_1 FILLER_48_223 ();
 sg13g2_fill_2 FILLER_48_237 ();
 sg13g2_fill_1 FILLER_48_239 ();
 sg13g2_decap_4 FILLER_48_246 ();
 sg13g2_fill_2 FILLER_48_276 ();
 sg13g2_fill_1 FILLER_48_278 ();
 sg13g2_fill_2 FILLER_48_309 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_fill_2 FILLER_48_328 ();
 sg13g2_fill_2 FILLER_48_352 ();
 sg13g2_fill_2 FILLER_48_359 ();
 sg13g2_decap_4 FILLER_48_367 ();
 sg13g2_fill_2 FILLER_48_371 ();
 sg13g2_fill_2 FILLER_48_401 ();
 sg13g2_fill_2 FILLER_48_431 ();
 sg13g2_fill_1 FILLER_48_456 ();
 sg13g2_decap_8 FILLER_48_461 ();
 sg13g2_fill_2 FILLER_48_468 ();
 sg13g2_fill_2 FILLER_48_478 ();
 sg13g2_fill_2 FILLER_48_569 ();
 sg13g2_fill_1 FILLER_48_571 ();
 sg13g2_fill_2 FILLER_48_577 ();
 sg13g2_fill_1 FILLER_48_579 ();
 sg13g2_fill_2 FILLER_48_611 ();
 sg13g2_fill_1 FILLER_48_613 ();
 sg13g2_fill_1 FILLER_48_647 ();
 sg13g2_fill_2 FILLER_48_658 ();
 sg13g2_fill_2 FILLER_48_696 ();
 sg13g2_fill_1 FILLER_48_698 ();
 sg13g2_fill_2 FILLER_48_703 ();
 sg13g2_fill_2 FILLER_48_714 ();
 sg13g2_fill_1 FILLER_48_725 ();
 sg13g2_fill_2 FILLER_48_735 ();
 sg13g2_fill_2 FILLER_48_772 ();
 sg13g2_fill_1 FILLER_48_774 ();
 sg13g2_fill_2 FILLER_48_792 ();
 sg13g2_decap_4 FILLER_48_824 ();
 sg13g2_fill_1 FILLER_48_828 ();
 sg13g2_fill_2 FILLER_48_841 ();
 sg13g2_decap_4 FILLER_48_858 ();
 sg13g2_fill_2 FILLER_49_26 ();
 sg13g2_fill_2 FILLER_49_45 ();
 sg13g2_fill_1 FILLER_49_88 ();
 sg13g2_fill_1 FILLER_49_94 ();
 sg13g2_fill_1 FILLER_49_104 ();
 sg13g2_fill_2 FILLER_49_118 ();
 sg13g2_fill_1 FILLER_49_137 ();
 sg13g2_fill_1 FILLER_49_147 ();
 sg13g2_fill_2 FILLER_49_165 ();
 sg13g2_fill_1 FILLER_49_233 ();
 sg13g2_fill_1 FILLER_49_278 ();
 sg13g2_fill_2 FILLER_49_288 ();
 sg13g2_fill_1 FILLER_49_290 ();
 sg13g2_fill_2 FILLER_49_352 ();
 sg13g2_fill_2 FILLER_49_415 ();
 sg13g2_fill_2 FILLER_49_445 ();
 sg13g2_fill_1 FILLER_49_478 ();
 sg13g2_fill_1 FILLER_49_496 ();
 sg13g2_decap_8 FILLER_49_519 ();
 sg13g2_decap_8 FILLER_49_526 ();
 sg13g2_fill_2 FILLER_49_533 ();
 sg13g2_fill_1 FILLER_49_553 ();
 sg13g2_fill_2 FILLER_49_562 ();
 sg13g2_fill_1 FILLER_49_564 ();
 sg13g2_fill_1 FILLER_49_578 ();
 sg13g2_decap_8 FILLER_49_596 ();
 sg13g2_fill_2 FILLER_49_603 ();
 sg13g2_decap_4 FILLER_49_623 ();
 sg13g2_fill_2 FILLER_49_627 ();
 sg13g2_decap_4 FILLER_49_645 ();
 sg13g2_fill_2 FILLER_49_664 ();
 sg13g2_fill_2 FILLER_49_674 ();
 sg13g2_fill_1 FILLER_49_676 ();
 sg13g2_decap_4 FILLER_49_683 ();
 sg13g2_fill_2 FILLER_49_687 ();
 sg13g2_decap_8 FILLER_49_716 ();
 sg13g2_fill_2 FILLER_49_723 ();
 sg13g2_decap_4 FILLER_49_745 ();
 sg13g2_fill_1 FILLER_49_749 ();
 sg13g2_fill_1 FILLER_49_759 ();
 sg13g2_fill_1 FILLER_49_765 ();
 sg13g2_fill_2 FILLER_49_774 ();
 sg13g2_fill_1 FILLER_49_776 ();
 sg13g2_decap_8 FILLER_49_792 ();
 sg13g2_fill_2 FILLER_49_799 ();
 sg13g2_fill_2 FILLER_49_818 ();
 sg13g2_decap_4 FILLER_49_833 ();
 sg13g2_fill_2 FILLER_49_837 ();
 sg13g2_decap_8 FILLER_49_849 ();
 sg13g2_decap_4 FILLER_49_856 ();
 sg13g2_fill_2 FILLER_49_860 ();
 sg13g2_fill_2 FILLER_50_40 ();
 sg13g2_fill_1 FILLER_50_62 ();
 sg13g2_fill_1 FILLER_50_72 ();
 sg13g2_fill_1 FILLER_50_100 ();
 sg13g2_fill_2 FILLER_50_139 ();
 sg13g2_fill_1 FILLER_50_141 ();
 sg13g2_fill_2 FILLER_50_147 ();
 sg13g2_fill_1 FILLER_50_149 ();
 sg13g2_fill_1 FILLER_50_160 ();
 sg13g2_fill_2 FILLER_50_176 ();
 sg13g2_fill_1 FILLER_50_204 ();
 sg13g2_fill_2 FILLER_50_213 ();
 sg13g2_fill_2 FILLER_50_229 ();
 sg13g2_fill_1 FILLER_50_240 ();
 sg13g2_fill_2 FILLER_50_249 ();
 sg13g2_fill_1 FILLER_50_251 ();
 sg13g2_fill_2 FILLER_50_263 ();
 sg13g2_fill_1 FILLER_50_265 ();
 sg13g2_fill_2 FILLER_50_282 ();
 sg13g2_fill_2 FILLER_50_289 ();
 sg13g2_fill_1 FILLER_50_291 ();
 sg13g2_fill_1 FILLER_50_314 ();
 sg13g2_fill_2 FILLER_50_361 ();
 sg13g2_fill_1 FILLER_50_514 ();
 sg13g2_decap_4 FILLER_50_561 ();
 sg13g2_fill_1 FILLER_50_565 ();
 sg13g2_decap_4 FILLER_50_610 ();
 sg13g2_fill_1 FILLER_50_618 ();
 sg13g2_decap_8 FILLER_50_636 ();
 sg13g2_decap_4 FILLER_50_643 ();
 sg13g2_decap_4 FILLER_50_670 ();
 sg13g2_fill_1 FILLER_50_674 ();
 sg13g2_fill_2 FILLER_50_679 ();
 sg13g2_fill_1 FILLER_50_681 ();
 sg13g2_fill_1 FILLER_50_686 ();
 sg13g2_fill_1 FILLER_50_690 ();
 sg13g2_fill_1 FILLER_50_703 ();
 sg13g2_decap_4 FILLER_50_714 ();
 sg13g2_fill_1 FILLER_50_718 ();
 sg13g2_fill_2 FILLER_50_731 ();
 sg13g2_fill_2 FILLER_50_773 ();
 sg13g2_fill_2 FILLER_50_803 ();
 sg13g2_fill_1 FILLER_50_825 ();
 sg13g2_fill_2 FILLER_50_859 ();
 sg13g2_fill_1 FILLER_50_861 ();
 sg13g2_fill_2 FILLER_51_56 ();
 sg13g2_fill_2 FILLER_51_62 ();
 sg13g2_fill_2 FILLER_51_112 ();
 sg13g2_fill_1 FILLER_51_133 ();
 sg13g2_fill_2 FILLER_51_180 ();
 sg13g2_fill_2 FILLER_51_191 ();
 sg13g2_fill_2 FILLER_51_324 ();
 sg13g2_fill_1 FILLER_51_349 ();
 sg13g2_fill_2 FILLER_51_390 ();
 sg13g2_fill_1 FILLER_51_432 ();
 sg13g2_fill_1 FILLER_51_438 ();
 sg13g2_decap_4 FILLER_51_453 ();
 sg13g2_fill_1 FILLER_51_461 ();
 sg13g2_fill_2 FILLER_51_471 ();
 sg13g2_fill_1 FILLER_51_473 ();
 sg13g2_decap_8 FILLER_51_478 ();
 sg13g2_fill_2 FILLER_51_485 ();
 sg13g2_fill_1 FILLER_51_505 ();
 sg13g2_fill_2 FILLER_51_536 ();
 sg13g2_fill_2 FILLER_51_552 ();
 sg13g2_decap_8 FILLER_51_568 ();
 sg13g2_fill_2 FILLER_51_575 ();
 sg13g2_decap_4 FILLER_51_629 ();
 sg13g2_fill_2 FILLER_51_633 ();
 sg13g2_fill_2 FILLER_51_647 ();
 sg13g2_fill_2 FILLER_51_658 ();
 sg13g2_fill_1 FILLER_51_660 ();
 sg13g2_fill_1 FILLER_51_674 ();
 sg13g2_fill_1 FILLER_51_694 ();
 sg13g2_fill_2 FILLER_51_726 ();
 sg13g2_fill_1 FILLER_51_728 ();
 sg13g2_fill_2 FILLER_51_757 ();
 sg13g2_fill_2 FILLER_51_791 ();
 sg13g2_fill_1 FILLER_51_793 ();
 sg13g2_fill_1 FILLER_51_810 ();
 sg13g2_decap_4 FILLER_51_819 ();
 sg13g2_fill_2 FILLER_51_823 ();
 sg13g2_fill_1 FILLER_51_830 ();
 sg13g2_fill_1 FILLER_51_842 ();
 sg13g2_fill_1 FILLER_51_861 ();
 sg13g2_fill_2 FILLER_52_33 ();
 sg13g2_fill_2 FILLER_52_127 ();
 sg13g2_fill_1 FILLER_52_129 ();
 sg13g2_fill_2 FILLER_52_191 ();
 sg13g2_fill_1 FILLER_52_238 ();
 sg13g2_fill_2 FILLER_52_272 ();
 sg13g2_fill_2 FILLER_52_284 ();
 sg13g2_fill_2 FILLER_52_291 ();
 sg13g2_fill_1 FILLER_52_358 ();
 sg13g2_fill_1 FILLER_52_371 ();
 sg13g2_fill_2 FILLER_52_405 ();
 sg13g2_fill_2 FILLER_52_419 ();
 sg13g2_decap_4 FILLER_52_472 ();
 sg13g2_fill_2 FILLER_52_476 ();
 sg13g2_fill_2 FILLER_52_486 ();
 sg13g2_fill_1 FILLER_52_488 ();
 sg13g2_decap_4 FILLER_52_505 ();
 sg13g2_decap_4 FILLER_52_565 ();
 sg13g2_fill_1 FILLER_52_569 ();
 sg13g2_fill_1 FILLER_52_580 ();
 sg13g2_decap_4 FILLER_52_603 ();
 sg13g2_fill_2 FILLER_52_607 ();
 sg13g2_fill_2 FILLER_52_629 ();
 sg13g2_fill_1 FILLER_52_659 ();
 sg13g2_decap_8 FILLER_52_676 ();
 sg13g2_fill_2 FILLER_52_683 ();
 sg13g2_fill_2 FILLER_52_689 ();
 sg13g2_fill_1 FILLER_52_691 ();
 sg13g2_decap_4 FILLER_52_749 ();
 sg13g2_fill_2 FILLER_52_753 ();
 sg13g2_fill_2 FILLER_52_771 ();
 sg13g2_decap_8 FILLER_52_796 ();
 sg13g2_fill_2 FILLER_52_803 ();
 sg13g2_fill_1 FILLER_52_805 ();
 sg13g2_fill_1 FILLER_52_817 ();
 sg13g2_fill_2 FILLER_52_823 ();
 sg13g2_fill_2 FILLER_52_859 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_fill_2 FILLER_53_39 ();
 sg13g2_fill_2 FILLER_53_51 ();
 sg13g2_fill_1 FILLER_53_66 ();
 sg13g2_fill_1 FILLER_53_91 ();
 sg13g2_fill_2 FILLER_53_197 ();
 sg13g2_fill_1 FILLER_53_235 ();
 sg13g2_fill_2 FILLER_53_282 ();
 sg13g2_fill_1 FILLER_53_318 ();
 sg13g2_fill_1 FILLER_53_380 ();
 sg13g2_fill_2 FILLER_53_459 ();
 sg13g2_fill_1 FILLER_53_461 ();
 sg13g2_fill_1 FILLER_53_474 ();
 sg13g2_fill_1 FILLER_53_540 ();
 sg13g2_fill_1 FILLER_53_568 ();
 sg13g2_decap_4 FILLER_53_594 ();
 sg13g2_fill_1 FILLER_53_598 ();
 sg13g2_fill_2 FILLER_53_607 ();
 sg13g2_fill_1 FILLER_53_609 ();
 sg13g2_fill_2 FILLER_53_618 ();
 sg13g2_fill_1 FILLER_53_620 ();
 sg13g2_decap_4 FILLER_53_627 ();
 sg13g2_fill_2 FILLER_53_636 ();
 sg13g2_fill_1 FILLER_53_638 ();
 sg13g2_fill_2 FILLER_53_655 ();
 sg13g2_fill_1 FILLER_53_657 ();
 sg13g2_fill_2 FILLER_53_688 ();
 sg13g2_fill_1 FILLER_53_690 ();
 sg13g2_fill_1 FILLER_53_696 ();
 sg13g2_decap_4 FILLER_53_727 ();
 sg13g2_fill_2 FILLER_53_747 ();
 sg13g2_fill_1 FILLER_53_749 ();
 sg13g2_fill_2 FILLER_53_755 ();
 sg13g2_decap_8 FILLER_53_762 ();
 sg13g2_decap_8 FILLER_53_769 ();
 sg13g2_fill_2 FILLER_53_776 ();
 sg13g2_fill_1 FILLER_53_778 ();
 sg13g2_decap_8 FILLER_53_802 ();
 sg13g2_fill_2 FILLER_53_809 ();
 sg13g2_fill_1 FILLER_53_814 ();
 sg13g2_fill_2 FILLER_53_825 ();
 sg13g2_fill_2 FILLER_53_837 ();
 sg13g2_fill_2 FILLER_53_860 ();
 sg13g2_fill_2 FILLER_54_34 ();
 sg13g2_fill_2 FILLER_54_70 ();
 sg13g2_fill_2 FILLER_54_121 ();
 sg13g2_fill_2 FILLER_54_170 ();
 sg13g2_fill_1 FILLER_54_204 ();
 sg13g2_fill_2 FILLER_54_240 ();
 sg13g2_fill_1 FILLER_54_242 ();
 sg13g2_fill_1 FILLER_54_258 ();
 sg13g2_fill_1 FILLER_54_299 ();
 sg13g2_fill_1 FILLER_54_307 ();
 sg13g2_fill_2 FILLER_54_362 ();
 sg13g2_fill_2 FILLER_54_390 ();
 sg13g2_fill_1 FILLER_54_392 ();
 sg13g2_fill_1 FILLER_54_428 ();
 sg13g2_fill_2 FILLER_54_468 ();
 sg13g2_fill_1 FILLER_54_470 ();
 sg13g2_fill_2 FILLER_54_474 ();
 sg13g2_decap_4 FILLER_54_502 ();
 sg13g2_fill_2 FILLER_54_558 ();
 sg13g2_fill_1 FILLER_54_560 ();
 sg13g2_fill_2 FILLER_54_579 ();
 sg13g2_fill_1 FILLER_54_581 ();
 sg13g2_fill_2 FILLER_54_588 ();
 sg13g2_fill_1 FILLER_54_590 ();
 sg13g2_fill_2 FILLER_54_662 ();
 sg13g2_decap_8 FILLER_54_669 ();
 sg13g2_fill_2 FILLER_54_676 ();
 sg13g2_fill_1 FILLER_54_698 ();
 sg13g2_fill_1 FILLER_54_720 ();
 sg13g2_fill_2 FILLER_54_770 ();
 sg13g2_fill_1 FILLER_54_808 ();
 sg13g2_fill_1 FILLER_54_853 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_60 ();
 sg13g2_fill_2 FILLER_55_97 ();
 sg13g2_fill_2 FILLER_55_125 ();
 sg13g2_fill_1 FILLER_55_127 ();
 sg13g2_fill_2 FILLER_55_136 ();
 sg13g2_fill_1 FILLER_55_138 ();
 sg13g2_fill_1 FILLER_55_170 ();
 sg13g2_fill_2 FILLER_55_221 ();
 sg13g2_fill_1 FILLER_55_268 ();
 sg13g2_fill_1 FILLER_55_321 ();
 sg13g2_fill_1 FILLER_55_416 ();
 sg13g2_fill_1 FILLER_55_510 ();
 sg13g2_fill_2 FILLER_55_541 ();
 sg13g2_fill_1 FILLER_55_543 ();
 sg13g2_fill_2 FILLER_55_573 ();
 sg13g2_fill_1 FILLER_55_597 ();
 sg13g2_fill_2 FILLER_55_616 ();
 sg13g2_fill_1 FILLER_55_618 ();
 sg13g2_decap_4 FILLER_55_624 ();
 sg13g2_fill_1 FILLER_55_628 ();
 sg13g2_fill_2 FILLER_55_652 ();
 sg13g2_decap_8 FILLER_55_676 ();
 sg13g2_decap_4 FILLER_55_683 ();
 sg13g2_fill_2 FILLER_55_687 ();
 sg13g2_fill_2 FILLER_55_734 ();
 sg13g2_fill_2 FILLER_55_741 ();
 sg13g2_fill_1 FILLER_55_748 ();
 sg13g2_fill_1 FILLER_55_757 ();
 sg13g2_fill_1 FILLER_55_773 ();
 sg13g2_decap_4 FILLER_55_791 ();
 sg13g2_fill_2 FILLER_55_795 ();
 sg13g2_decap_4 FILLER_55_800 ();
 sg13g2_fill_2 FILLER_55_829 ();
 sg13g2_fill_1 FILLER_55_861 ();
 sg13g2_fill_1 FILLER_56_21 ();
 sg13g2_fill_1 FILLER_56_36 ();
 sg13g2_fill_2 FILLER_56_80 ();
 sg13g2_fill_1 FILLER_56_98 ();
 sg13g2_fill_2 FILLER_56_191 ();
 sg13g2_fill_1 FILLER_56_193 ();
 sg13g2_fill_1 FILLER_56_220 ();
 sg13g2_fill_2 FILLER_56_247 ();
 sg13g2_fill_1 FILLER_56_249 ();
 sg13g2_fill_2 FILLER_56_280 ();
 sg13g2_fill_1 FILLER_56_282 ();
 sg13g2_fill_1 FILLER_56_310 ();
 sg13g2_fill_2 FILLER_56_324 ();
 sg13g2_fill_1 FILLER_56_398 ();
 sg13g2_fill_1 FILLER_56_432 ();
 sg13g2_fill_2 FILLER_56_446 ();
 sg13g2_fill_2 FILLER_56_465 ();
 sg13g2_fill_1 FILLER_56_467 ();
 sg13g2_fill_2 FILLER_56_477 ();
 sg13g2_decap_8 FILLER_56_501 ();
 sg13g2_decap_8 FILLER_56_586 ();
 sg13g2_decap_8 FILLER_56_593 ();
 sg13g2_fill_1 FILLER_56_600 ();
 sg13g2_fill_2 FILLER_56_638 ();
 sg13g2_fill_1 FILLER_56_640 ();
 sg13g2_fill_2 FILLER_56_651 ();
 sg13g2_fill_1 FILLER_56_653 ();
 sg13g2_decap_4 FILLER_56_678 ();
 sg13g2_fill_2 FILLER_56_728 ();
 sg13g2_fill_1 FILLER_56_730 ();
 sg13g2_fill_2 FILLER_56_748 ();
 sg13g2_fill_1 FILLER_56_750 ();
 sg13g2_decap_4 FILLER_56_759 ();
 sg13g2_decap_4 FILLER_56_779 ();
 sg13g2_fill_2 FILLER_56_783 ();
 sg13g2_fill_2 FILLER_56_797 ();
 sg13g2_fill_1 FILLER_56_817 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_fill_1 FILLER_57_35 ();
 sg13g2_fill_1 FILLER_57_63 ();
 sg13g2_fill_2 FILLER_57_112 ();
 sg13g2_fill_1 FILLER_57_114 ();
 sg13g2_fill_2 FILLER_57_165 ();
 sg13g2_fill_1 FILLER_57_180 ();
 sg13g2_fill_2 FILLER_57_186 ();
 sg13g2_fill_2 FILLER_57_209 ();
 sg13g2_fill_2 FILLER_57_256 ();
 sg13g2_fill_2 FILLER_57_281 ();
 sg13g2_fill_1 FILLER_57_293 ();
 sg13g2_fill_1 FILLER_57_332 ();
 sg13g2_fill_2 FILLER_57_396 ();
 sg13g2_fill_1 FILLER_57_459 ();
 sg13g2_fill_1 FILLER_57_465 ();
 sg13g2_decap_8 FILLER_57_514 ();
 sg13g2_decap_8 FILLER_57_521 ();
 sg13g2_fill_2 FILLER_57_528 ();
 sg13g2_fill_1 FILLER_57_530 ();
 sg13g2_fill_2 FILLER_57_538 ();
 sg13g2_fill_1 FILLER_57_540 ();
 sg13g2_decap_4 FILLER_57_545 ();
 sg13g2_fill_2 FILLER_57_549 ();
 sg13g2_decap_8 FILLER_57_558 ();
 sg13g2_fill_2 FILLER_57_565 ();
 sg13g2_fill_1 FILLER_57_567 ();
 sg13g2_decap_4 FILLER_57_572 ();
 sg13g2_decap_8 FILLER_57_599 ();
 sg13g2_fill_1 FILLER_57_606 ();
 sg13g2_fill_2 FILLER_57_640 ();
 sg13g2_decap_4 FILLER_57_657 ();
 sg13g2_fill_2 FILLER_57_661 ();
 sg13g2_fill_2 FILLER_57_668 ();
 sg13g2_fill_1 FILLER_57_670 ();
 sg13g2_fill_2 FILLER_57_676 ();
 sg13g2_fill_1 FILLER_57_678 ();
 sg13g2_fill_1 FILLER_57_696 ();
 sg13g2_fill_1 FILLER_57_773 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_49 ();
 sg13g2_fill_1 FILLER_58_86 ();
 sg13g2_fill_1 FILLER_58_97 ();
 sg13g2_fill_1 FILLER_58_141 ();
 sg13g2_fill_1 FILLER_58_185 ();
 sg13g2_fill_2 FILLER_58_360 ();
 sg13g2_fill_1 FILLER_58_362 ();
 sg13g2_fill_1 FILLER_58_439 ();
 sg13g2_fill_1 FILLER_58_462 ();
 sg13g2_fill_2 FILLER_58_520 ();
 sg13g2_fill_1 FILLER_58_522 ();
 sg13g2_fill_2 FILLER_58_577 ();
 sg13g2_fill_2 FILLER_58_605 ();
 sg13g2_fill_2 FILLER_58_615 ();
 sg13g2_fill_1 FILLER_58_617 ();
 sg13g2_fill_2 FILLER_58_627 ();
 sg13g2_fill_2 FILLER_58_645 ();
 sg13g2_fill_2 FILLER_58_710 ();
 sg13g2_fill_1 FILLER_58_712 ();
 sg13g2_fill_2 FILLER_58_727 ();
 sg13g2_fill_2 FILLER_58_749 ();
 sg13g2_fill_1 FILLER_58_861 ();
 sg13g2_fill_1 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_133 ();
 sg13g2_fill_1 FILLER_59_135 ();
 sg13g2_fill_1 FILLER_59_172 ();
 sg13g2_fill_1 FILLER_59_223 ();
 sg13g2_fill_1 FILLER_59_457 ();
 sg13g2_fill_2 FILLER_59_467 ();
 sg13g2_fill_1 FILLER_59_482 ();
 sg13g2_fill_2 FILLER_59_492 ();
 sg13g2_fill_2 FILLER_59_515 ();
 sg13g2_fill_2 FILLER_59_550 ();
 sg13g2_fill_1 FILLER_59_552 ();
 sg13g2_fill_1 FILLER_59_557 ();
 sg13g2_fill_2 FILLER_59_619 ();
 sg13g2_fill_1 FILLER_59_621 ();
 sg13g2_decap_8 FILLER_59_645 ();
 sg13g2_fill_2 FILLER_59_668 ();
 sg13g2_fill_1 FILLER_59_670 ();
 sg13g2_fill_1 FILLER_59_680 ();
 sg13g2_fill_2 FILLER_59_710 ();
 sg13g2_fill_1 FILLER_59_821 ();
 sg13g2_fill_1 FILLER_60_56 ();
 sg13g2_fill_2 FILLER_60_97 ();
 sg13g2_fill_2 FILLER_60_140 ();
 sg13g2_fill_1 FILLER_60_142 ();
 sg13g2_fill_1 FILLER_60_153 ();
 sg13g2_fill_2 FILLER_60_191 ();
 sg13g2_fill_2 FILLER_60_224 ();
 sg13g2_fill_1 FILLER_60_226 ();
 sg13g2_fill_1 FILLER_60_316 ();
 sg13g2_fill_1 FILLER_60_362 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_fill_1 FILLER_60_409 ();
 sg13g2_fill_2 FILLER_60_436 ();
 sg13g2_fill_2 FILLER_60_510 ();
 sg13g2_fill_1 FILLER_60_521 ();
 sg13g2_fill_2 FILLER_60_526 ();
 sg13g2_fill_1 FILLER_60_528 ();
 sg13g2_fill_2 FILLER_60_542 ();
 sg13g2_fill_1 FILLER_60_544 ();
 sg13g2_fill_2 FILLER_60_600 ();
 sg13g2_fill_2 FILLER_60_663 ();
 sg13g2_fill_2 FILLER_60_814 ();
 sg13g2_fill_2 FILLER_60_859 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_fill_2 FILLER_61_18 ();
 sg13g2_fill_1 FILLER_61_20 ();
 sg13g2_fill_2 FILLER_61_51 ();
 sg13g2_fill_1 FILLER_61_94 ();
 sg13g2_fill_1 FILLER_61_104 ();
 sg13g2_fill_2 FILLER_61_174 ();
 sg13g2_fill_1 FILLER_61_191 ();
 sg13g2_fill_2 FILLER_61_218 ();
 sg13g2_fill_1 FILLER_61_249 ();
 sg13g2_fill_1 FILLER_61_263 ();
 sg13g2_fill_2 FILLER_61_313 ();
 sg13g2_fill_1 FILLER_61_323 ();
 sg13g2_fill_1 FILLER_61_333 ();
 sg13g2_fill_2 FILLER_61_364 ();
 sg13g2_fill_2 FILLER_61_374 ();
 sg13g2_fill_2 FILLER_61_398 ();
 sg13g2_fill_2 FILLER_61_409 ();
 sg13g2_fill_1 FILLER_61_411 ();
 sg13g2_fill_1 FILLER_61_437 ();
 sg13g2_decap_8 FILLER_61_459 ();
 sg13g2_fill_2 FILLER_61_466 ();
 sg13g2_fill_1 FILLER_61_468 ();
 sg13g2_fill_2 FILLER_61_479 ();
 sg13g2_decap_4 FILLER_61_532 ();
 sg13g2_fill_1 FILLER_61_545 ();
 sg13g2_fill_2 FILLER_61_598 ();
 sg13g2_fill_2 FILLER_61_605 ();
 sg13g2_fill_2 FILLER_61_658 ();
 sg13g2_fill_1 FILLER_61_660 ();
 sg13g2_fill_2 FILLER_61_678 ();
 sg13g2_fill_2 FILLER_61_694 ();
 sg13g2_fill_1 FILLER_61_708 ();
 sg13g2_fill_2 FILLER_61_722 ();
 sg13g2_fill_1 FILLER_61_724 ();
 sg13g2_fill_2 FILLER_61_742 ();
 sg13g2_fill_1 FILLER_61_744 ();
 sg13g2_fill_2 FILLER_61_785 ();
 sg13g2_fill_1 FILLER_61_787 ();
 sg13g2_fill_2 FILLER_61_831 ();
 sg13g2_fill_1 FILLER_61_842 ();
 sg13g2_fill_2 FILLER_61_860 ();
 sg13g2_fill_2 FILLER_62_50 ();
 sg13g2_fill_1 FILLER_62_52 ();
 sg13g2_fill_1 FILLER_62_62 ();
 sg13g2_fill_2 FILLER_62_176 ();
 sg13g2_fill_1 FILLER_62_198 ();
 sg13g2_fill_2 FILLER_62_208 ();
 sg13g2_fill_1 FILLER_62_245 ();
 sg13g2_fill_2 FILLER_62_263 ();
 sg13g2_fill_1 FILLER_62_287 ();
 sg13g2_fill_2 FILLER_62_311 ();
 sg13g2_fill_1 FILLER_62_313 ();
 sg13g2_fill_2 FILLER_62_331 ();
 sg13g2_fill_1 FILLER_62_333 ();
 sg13g2_fill_1 FILLER_62_365 ();
 sg13g2_fill_1 FILLER_62_439 ();
 sg13g2_decap_8 FILLER_62_462 ();
 sg13g2_fill_2 FILLER_62_469 ();
 sg13g2_fill_1 FILLER_62_471 ();
 sg13g2_fill_1 FILLER_62_493 ();
 sg13g2_fill_2 FILLER_62_512 ();
 sg13g2_fill_1 FILLER_62_541 ();
 sg13g2_fill_2 FILLER_62_581 ();
 sg13g2_fill_1 FILLER_62_583 ();
 sg13g2_fill_2 FILLER_62_604 ();
 sg13g2_fill_2 FILLER_62_623 ();
 sg13g2_fill_2 FILLER_62_681 ();
 sg13g2_fill_1 FILLER_62_687 ();
 sg13g2_fill_2 FILLER_62_697 ();
 sg13g2_fill_1 FILLER_62_748 ();
 sg13g2_fill_2 FILLER_62_788 ();
 sg13g2_fill_1 FILLER_62_790 ();
 sg13g2_fill_2 FILLER_62_805 ();
 sg13g2_fill_1 FILLER_62_812 ();
 sg13g2_fill_2 FILLER_62_823 ();
 sg13g2_fill_1 FILLER_62_825 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_2 ();
 sg13g2_fill_1 FILLER_63_38 ();
 sg13g2_fill_2 FILLER_63_84 ();
 sg13g2_fill_1 FILLER_63_86 ();
 sg13g2_fill_1 FILLER_63_113 ();
 sg13g2_fill_1 FILLER_63_123 ();
 sg13g2_fill_1 FILLER_63_138 ();
 sg13g2_fill_1 FILLER_63_181 ();
 sg13g2_fill_1 FILLER_63_224 ();
 sg13g2_fill_1 FILLER_63_246 ();
 sg13g2_fill_1 FILLER_63_300 ();
 sg13g2_fill_2 FILLER_63_325 ();
 sg13g2_fill_2 FILLER_63_353 ();
 sg13g2_fill_2 FILLER_63_374 ();
 sg13g2_fill_2 FILLER_63_411 ();
 sg13g2_decap_8 FILLER_63_465 ();
 sg13g2_fill_1 FILLER_63_480 ();
 sg13g2_fill_2 FILLER_63_578 ();
 sg13g2_fill_1 FILLER_63_595 ();
 sg13g2_fill_2 FILLER_63_671 ();
 sg13g2_fill_1 FILLER_63_673 ();
 sg13g2_fill_2 FILLER_63_705 ();
 sg13g2_fill_1 FILLER_63_793 ();
 sg13g2_fill_2 FILLER_63_834 ();
 sg13g2_fill_2 FILLER_64_43 ();
 sg13g2_fill_1 FILLER_64_55 ();
 sg13g2_fill_1 FILLER_64_121 ();
 sg13g2_fill_2 FILLER_64_157 ();
 sg13g2_fill_1 FILLER_64_159 ();
 sg13g2_fill_1 FILLER_64_199 ();
 sg13g2_fill_2 FILLER_64_237 ();
 sg13g2_fill_1 FILLER_64_239 ();
 sg13g2_fill_2 FILLER_64_307 ();
 sg13g2_fill_2 FILLER_64_317 ();
 sg13g2_fill_1 FILLER_64_362 ();
 sg13g2_fill_1 FILLER_64_395 ();
 sg13g2_fill_2 FILLER_64_438 ();
 sg13g2_fill_1 FILLER_64_440 ();
 sg13g2_decap_4 FILLER_64_474 ();
 sg13g2_fill_1 FILLER_64_478 ();
 sg13g2_fill_1 FILLER_64_521 ();
 sg13g2_fill_1 FILLER_64_555 ();
 sg13g2_fill_1 FILLER_64_565 ();
 sg13g2_fill_2 FILLER_64_614 ();
 sg13g2_fill_2 FILLER_64_621 ();
 sg13g2_fill_1 FILLER_64_632 ();
 sg13g2_fill_1 FILLER_64_642 ();
 sg13g2_fill_1 FILLER_64_656 ();
 sg13g2_decap_4 FILLER_64_683 ();
 sg13g2_fill_2 FILLER_64_687 ();
 sg13g2_fill_2 FILLER_64_743 ();
 sg13g2_fill_2 FILLER_64_758 ();
 sg13g2_fill_1 FILLER_64_770 ();
 sg13g2_fill_2 FILLER_64_816 ();
 sg13g2_fill_1 FILLER_64_818 ();
 sg13g2_fill_1 FILLER_64_845 ();
 sg13g2_fill_2 FILLER_64_859 ();
 sg13g2_fill_1 FILLER_64_861 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_2 ();
 sg13g2_fill_1 FILLER_65_31 ();
 sg13g2_fill_2 FILLER_65_136 ();
 sg13g2_fill_1 FILLER_65_231 ();
 sg13g2_fill_1 FILLER_65_285 ();
 sg13g2_fill_1 FILLER_65_316 ();
 sg13g2_fill_1 FILLER_65_404 ();
 sg13g2_fill_2 FILLER_65_410 ();
 sg13g2_fill_1 FILLER_65_412 ();
 sg13g2_fill_1 FILLER_65_430 ();
 sg13g2_decap_8 FILLER_65_483 ();
 sg13g2_decap_4 FILLER_65_490 ();
 sg13g2_fill_1 FILLER_65_494 ();
 sg13g2_fill_2 FILLER_65_527 ();
 sg13g2_fill_1 FILLER_65_529 ();
 sg13g2_fill_1 FILLER_65_571 ();
 sg13g2_fill_2 FILLER_65_580 ();
 sg13g2_fill_1 FILLER_65_646 ();
 sg13g2_fill_2 FILLER_65_663 ();
 sg13g2_fill_1 FILLER_65_665 ();
 sg13g2_fill_1 FILLER_65_678 ();
 sg13g2_fill_2 FILLER_65_698 ();
 sg13g2_fill_1 FILLER_65_720 ();
 sg13g2_fill_2 FILLER_65_798 ();
 sg13g2_fill_2 FILLER_65_826 ();
 sg13g2_fill_1 FILLER_65_828 ();
 sg13g2_fill_2 FILLER_65_834 ();
 sg13g2_fill_2 FILLER_66_65 ();
 sg13g2_fill_2 FILLER_66_75 ();
 sg13g2_fill_1 FILLER_66_77 ();
 sg13g2_fill_1 FILLER_66_109 ();
 sg13g2_fill_2 FILLER_66_119 ();
 sg13g2_fill_1 FILLER_66_130 ();
 sg13g2_fill_1 FILLER_66_183 ();
 sg13g2_fill_2 FILLER_66_245 ();
 sg13g2_fill_1 FILLER_66_321 ();
 sg13g2_fill_2 FILLER_66_327 ();
 sg13g2_fill_1 FILLER_66_350 ();
 sg13g2_fill_2 FILLER_66_361 ();
 sg13g2_fill_2 FILLER_66_368 ();
 sg13g2_fill_1 FILLER_66_370 ();
 sg13g2_fill_1 FILLER_66_386 ();
 sg13g2_fill_1 FILLER_66_415 ();
 sg13g2_fill_1 FILLER_66_488 ();
 sg13g2_fill_2 FILLER_66_515 ();
 sg13g2_fill_1 FILLER_66_522 ();
 sg13g2_fill_2 FILLER_66_548 ();
 sg13g2_fill_1 FILLER_66_550 ();
 sg13g2_fill_1 FILLER_66_557 ();
 sg13g2_fill_2 FILLER_66_566 ();
 sg13g2_fill_2 FILLER_66_577 ();
 sg13g2_fill_1 FILLER_66_579 ();
 sg13g2_fill_1 FILLER_66_600 ();
 sg13g2_fill_2 FILLER_66_605 ();
 sg13g2_fill_1 FILLER_66_641 ();
 sg13g2_fill_2 FILLER_66_666 ();
 sg13g2_fill_1 FILLER_66_668 ();
 sg13g2_fill_2 FILLER_66_687 ();
 sg13g2_decap_4 FILLER_66_698 ();
 sg13g2_fill_2 FILLER_66_702 ();
 sg13g2_fill_2 FILLER_66_718 ();
 sg13g2_fill_1 FILLER_66_720 ();
 sg13g2_fill_2 FILLER_66_744 ();
 sg13g2_fill_1 FILLER_66_746 ();
 sg13g2_fill_1 FILLER_66_752 ();
 sg13g2_fill_1 FILLER_66_757 ();
 sg13g2_fill_1 FILLER_66_797 ();
 sg13g2_fill_2 FILLER_66_818 ();
 sg13g2_fill_1 FILLER_66_850 ();
 sg13g2_fill_2 FILLER_66_860 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_2 ();
 sg13g2_fill_1 FILLER_67_59 ();
 sg13g2_fill_2 FILLER_67_65 ();
 sg13g2_fill_2 FILLER_67_80 ();
 sg13g2_fill_1 FILLER_67_109 ();
 sg13g2_fill_1 FILLER_67_205 ();
 sg13g2_fill_2 FILLER_67_274 ();
 sg13g2_fill_2 FILLER_67_291 ();
 sg13g2_fill_1 FILLER_67_293 ();
 sg13g2_fill_1 FILLER_67_371 ();
 sg13g2_fill_1 FILLER_67_404 ();
 sg13g2_fill_2 FILLER_67_418 ();
 sg13g2_fill_2 FILLER_67_425 ();
 sg13g2_fill_1 FILLER_67_427 ();
 sg13g2_fill_1 FILLER_67_466 ();
 sg13g2_fill_1 FILLER_67_614 ();
 sg13g2_fill_2 FILLER_67_632 ();
 sg13g2_fill_1 FILLER_67_634 ();
 sg13g2_fill_1 FILLER_67_643 ();
 sg13g2_fill_1 FILLER_67_666 ();
 sg13g2_fill_1 FILLER_67_695 ();
 sg13g2_fill_1 FILLER_67_741 ();
 sg13g2_fill_2 FILLER_67_794 ();
 sg13g2_fill_1 FILLER_68_26 ();
 sg13g2_fill_1 FILLER_68_69 ();
 sg13g2_fill_1 FILLER_68_86 ();
 sg13g2_fill_2 FILLER_68_157 ();
 sg13g2_fill_2 FILLER_68_185 ();
 sg13g2_fill_2 FILLER_68_285 ();
 sg13g2_fill_1 FILLER_68_287 ();
 sg13g2_fill_2 FILLER_68_297 ();
 sg13g2_fill_2 FILLER_68_371 ();
 sg13g2_fill_2 FILLER_68_408 ();
 sg13g2_fill_1 FILLER_68_410 ();
 sg13g2_fill_1 FILLER_68_444 ();
 sg13g2_fill_1 FILLER_68_497 ();
 sg13g2_decap_4 FILLER_68_535 ();
 sg13g2_fill_1 FILLER_68_578 ();
 sg13g2_fill_1 FILLER_68_618 ();
 sg13g2_fill_2 FILLER_68_640 ();
 sg13g2_fill_2 FILLER_68_668 ();
 sg13g2_fill_1 FILLER_68_679 ();
 sg13g2_fill_1 FILLER_68_715 ();
 sg13g2_fill_2 FILLER_68_814 ();
 sg13g2_fill_1 FILLER_68_829 ();
 sg13g2_fill_2 FILLER_68_834 ();
 sg13g2_fill_1 FILLER_68_861 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_27 ();
 sg13g2_fill_1 FILLER_69_49 ();
 sg13g2_fill_2 FILLER_69_108 ();
 sg13g2_fill_2 FILLER_69_115 ();
 sg13g2_fill_1 FILLER_69_125 ();
 sg13g2_fill_2 FILLER_69_283 ();
 sg13g2_fill_1 FILLER_69_311 ();
 sg13g2_fill_2 FILLER_69_399 ();
 sg13g2_fill_1 FILLER_69_401 ();
 sg13g2_fill_2 FILLER_69_442 ();
 sg13g2_fill_1 FILLER_69_444 ();
 sg13g2_fill_2 FILLER_69_461 ();
 sg13g2_fill_2 FILLER_69_509 ();
 sg13g2_fill_1 FILLER_69_563 ();
 sg13g2_fill_1 FILLER_69_601 ();
 sg13g2_decap_8 FILLER_69_609 ();
 sg13g2_decap_4 FILLER_69_616 ();
 sg13g2_fill_1 FILLER_69_620 ();
 sg13g2_decap_8 FILLER_69_626 ();
 sg13g2_decap_8 FILLER_69_633 ();
 sg13g2_fill_1 FILLER_69_640 ();
 sg13g2_fill_2 FILLER_69_650 ();
 sg13g2_fill_2 FILLER_69_656 ();
 sg13g2_fill_2 FILLER_69_734 ();
 sg13g2_fill_1 FILLER_69_753 ();
 sg13g2_fill_2 FILLER_69_775 ();
 sg13g2_fill_1 FILLER_69_777 ();
 sg13g2_fill_1 FILLER_69_791 ();
 sg13g2_fill_2 FILLER_69_826 ();
 sg13g2_fill_1 FILLER_70_37 ();
 sg13g2_fill_2 FILLER_70_102 ();
 sg13g2_fill_2 FILLER_70_109 ();
 sg13g2_fill_1 FILLER_70_116 ();
 sg13g2_fill_2 FILLER_70_211 ();
 sg13g2_fill_2 FILLER_70_365 ();
 sg13g2_fill_1 FILLER_70_383 ();
 sg13g2_fill_2 FILLER_70_394 ();
 sg13g2_fill_1 FILLER_70_410 ();
 sg13g2_fill_2 FILLER_70_415 ();
 sg13g2_fill_2 FILLER_70_422 ();
 sg13g2_fill_1 FILLER_70_424 ();
 sg13g2_fill_2 FILLER_70_436 ();
 sg13g2_fill_2 FILLER_70_539 ();
 sg13g2_fill_1 FILLER_70_562 ();
 sg13g2_fill_2 FILLER_70_589 ();
 sg13g2_fill_1 FILLER_70_677 ();
 sg13g2_fill_1 FILLER_70_686 ();
 sg13g2_fill_1 FILLER_70_720 ();
 sg13g2_fill_1 FILLER_70_747 ();
 sg13g2_fill_1 FILLER_70_769 ();
 sg13g2_fill_1 FILLER_70_778 ();
 sg13g2_fill_1 FILLER_70_791 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_30 ();
 sg13g2_fill_1 FILLER_71_37 ();
 sg13g2_fill_1 FILLER_71_69 ();
 sg13g2_fill_2 FILLER_71_77 ();
 sg13g2_fill_1 FILLER_71_79 ();
 sg13g2_fill_1 FILLER_71_101 ();
 sg13g2_fill_2 FILLER_71_112 ();
 sg13g2_fill_1 FILLER_71_114 ();
 sg13g2_fill_1 FILLER_71_123 ();
 sg13g2_fill_1 FILLER_71_146 ();
 sg13g2_fill_1 FILLER_71_166 ();
 sg13g2_fill_2 FILLER_71_257 ();
 sg13g2_fill_1 FILLER_71_259 ();
 sg13g2_fill_2 FILLER_71_277 ();
 sg13g2_fill_1 FILLER_71_279 ();
 sg13g2_fill_1 FILLER_71_332 ();
 sg13g2_fill_2 FILLER_71_369 ();
 sg13g2_fill_1 FILLER_71_381 ();
 sg13g2_fill_2 FILLER_71_405 ();
 sg13g2_fill_2 FILLER_71_454 ();
 sg13g2_fill_2 FILLER_71_474 ();
 sg13g2_fill_1 FILLER_71_497 ();
 sg13g2_fill_1 FILLER_71_575 ();
 sg13g2_fill_1 FILLER_71_599 ();
 sg13g2_fill_2 FILLER_71_741 ();
 sg13g2_fill_1 FILLER_71_743 ();
 sg13g2_fill_2 FILLER_71_766 ();
 sg13g2_fill_1 FILLER_71_795 ();
 sg13g2_fill_1 FILLER_71_809 ();
 sg13g2_fill_2 FILLER_71_827 ();
 sg13g2_fill_1 FILLER_71_846 ();
 sg13g2_fill_2 FILLER_71_851 ();
 sg13g2_fill_1 FILLER_72_91 ();
 sg13g2_fill_1 FILLER_72_97 ();
 sg13g2_fill_2 FILLER_72_103 ();
 sg13g2_fill_2 FILLER_72_114 ();
 sg13g2_fill_2 FILLER_72_126 ();
 sg13g2_fill_1 FILLER_72_128 ();
 sg13g2_fill_2 FILLER_72_134 ();
 sg13g2_fill_1 FILLER_72_136 ();
 sg13g2_fill_2 FILLER_72_223 ();
 sg13g2_fill_1 FILLER_72_225 ();
 sg13g2_fill_1 FILLER_72_235 ();
 sg13g2_fill_2 FILLER_72_244 ();
 sg13g2_fill_1 FILLER_72_246 ();
 sg13g2_fill_2 FILLER_72_252 ();
 sg13g2_fill_1 FILLER_72_254 ();
 sg13g2_fill_2 FILLER_72_272 ();
 sg13g2_fill_1 FILLER_72_274 ();
 sg13g2_fill_2 FILLER_72_280 ();
 sg13g2_fill_2 FILLER_72_298 ();
 sg13g2_fill_2 FILLER_72_309 ();
 sg13g2_fill_1 FILLER_72_311 ();
 sg13g2_fill_2 FILLER_72_334 ();
 sg13g2_fill_1 FILLER_72_336 ();
 sg13g2_fill_2 FILLER_72_353 ();
 sg13g2_fill_1 FILLER_72_355 ();
 sg13g2_fill_2 FILLER_72_361 ();
 sg13g2_fill_1 FILLER_72_363 ();
 sg13g2_fill_2 FILLER_72_379 ();
 sg13g2_fill_2 FILLER_72_424 ();
 sg13g2_fill_1 FILLER_72_426 ();
 sg13g2_fill_2 FILLER_72_442 ();
 sg13g2_fill_1 FILLER_72_507 ();
 sg13g2_fill_2 FILLER_72_512 ();
 sg13g2_fill_2 FILLER_72_542 ();
 sg13g2_fill_1 FILLER_72_553 ();
 sg13g2_fill_1 FILLER_72_568 ();
 sg13g2_fill_1 FILLER_72_635 ();
 sg13g2_fill_2 FILLER_72_701 ();
 sg13g2_fill_1 FILLER_72_716 ();
 sg13g2_fill_2 FILLER_72_771 ();
 sg13g2_fill_1 FILLER_72_783 ();
 sg13g2_fill_1 FILLER_72_789 ();
 sg13g2_fill_2 FILLER_72_798 ();
 sg13g2_fill_1 FILLER_72_800 ();
 sg13g2_fill_1 FILLER_72_806 ();
 sg13g2_fill_1 FILLER_72_835 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_2 ();
 sg13g2_fill_1 FILLER_73_25 ();
 sg13g2_fill_1 FILLER_73_61 ();
 sg13g2_fill_1 FILLER_73_67 ();
 sg13g2_fill_1 FILLER_73_107 ();
 sg13g2_fill_2 FILLER_73_120 ();
 sg13g2_fill_1 FILLER_73_122 ();
 sg13g2_fill_1 FILLER_73_162 ();
 sg13g2_fill_1 FILLER_73_177 ();
 sg13g2_fill_1 FILLER_73_199 ();
 sg13g2_fill_1 FILLER_73_220 ();
 sg13g2_fill_2 FILLER_73_228 ();
 sg13g2_fill_1 FILLER_73_338 ();
 sg13g2_fill_2 FILLER_73_360 ();
 sg13g2_fill_1 FILLER_73_362 ();
 sg13g2_fill_2 FILLER_73_369 ();
 sg13g2_fill_2 FILLER_73_422 ();
 sg13g2_fill_1 FILLER_73_430 ();
 sg13g2_fill_1 FILLER_73_440 ();
 sg13g2_fill_2 FILLER_73_527 ();
 sg13g2_fill_1 FILLER_73_538 ();
 sg13g2_fill_2 FILLER_73_635 ();
 sg13g2_fill_1 FILLER_73_673 ();
 sg13g2_fill_2 FILLER_73_694 ();
 sg13g2_fill_2 FILLER_73_710 ();
 sg13g2_fill_1 FILLER_73_734 ();
 sg13g2_fill_1 FILLER_73_744 ();
 sg13g2_fill_2 FILLER_73_750 ();
 sg13g2_fill_1 FILLER_73_752 ();
 sg13g2_fill_1 FILLER_73_768 ();
 sg13g2_fill_1 FILLER_73_795 ();
 sg13g2_fill_1 FILLER_73_818 ();
 sg13g2_fill_1 FILLER_73_832 ();
 sg13g2_fill_2 FILLER_73_837 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_63 ();
 sg13g2_fill_1 FILLER_74_70 ();
 sg13g2_fill_1 FILLER_74_87 ();
 sg13g2_fill_2 FILLER_74_150 ();
 sg13g2_fill_1 FILLER_74_152 ();
 sg13g2_fill_2 FILLER_74_189 ();
 sg13g2_fill_1 FILLER_74_197 ();
 sg13g2_fill_1 FILLER_74_206 ();
 sg13g2_fill_1 FILLER_74_217 ();
 sg13g2_fill_2 FILLER_74_226 ();
 sg13g2_fill_1 FILLER_74_228 ();
 sg13g2_fill_1 FILLER_74_244 ();
 sg13g2_fill_2 FILLER_74_256 ();
 sg13g2_fill_2 FILLER_74_292 ();
 sg13g2_fill_1 FILLER_74_308 ();
 sg13g2_fill_2 FILLER_74_326 ();
 sg13g2_fill_1 FILLER_74_328 ();
 sg13g2_fill_1 FILLER_74_362 ();
 sg13g2_fill_2 FILLER_74_429 ();
 sg13g2_fill_2 FILLER_74_451 ();
 sg13g2_fill_1 FILLER_74_495 ();
 sg13g2_fill_1 FILLER_74_583 ();
 sg13g2_fill_1 FILLER_74_601 ();
 sg13g2_fill_1 FILLER_74_650 ();
 sg13g2_fill_1 FILLER_74_736 ();
 sg13g2_fill_1 FILLER_74_776 ();
 sg13g2_fill_2 FILLER_74_803 ();
 sg13g2_fill_1 FILLER_74_805 ();
 sg13g2_fill_1 FILLER_74_829 ();
 sg13g2_fill_2 FILLER_74_860 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_51 ();
 sg13g2_fill_1 FILLER_75_72 ();
 sg13g2_fill_2 FILLER_75_105 ();
 sg13g2_fill_1 FILLER_75_111 ();
 sg13g2_fill_2 FILLER_75_169 ();
 sg13g2_fill_1 FILLER_75_241 ();
 sg13g2_fill_1 FILLER_75_333 ();
 sg13g2_fill_2 FILLER_75_344 ();
 sg13g2_fill_2 FILLER_75_361 ();
 sg13g2_fill_1 FILLER_75_363 ();
 sg13g2_fill_2 FILLER_75_375 ();
 sg13g2_fill_1 FILLER_75_406 ();
 sg13g2_fill_2 FILLER_75_424 ();
 sg13g2_fill_1 FILLER_75_470 ();
 sg13g2_fill_2 FILLER_75_506 ();
 sg13g2_fill_1 FILLER_75_517 ();
 sg13g2_fill_1 FILLER_75_533 ();
 sg13g2_fill_1 FILLER_75_602 ();
 sg13g2_fill_2 FILLER_75_613 ();
 sg13g2_fill_2 FILLER_75_620 ();
 sg13g2_fill_2 FILLER_75_637 ();
 sg13g2_fill_1 FILLER_75_644 ();
 sg13g2_fill_2 FILLER_75_740 ();
 sg13g2_fill_1 FILLER_75_742 ();
 sg13g2_fill_2 FILLER_75_748 ();
 sg13g2_fill_1 FILLER_75_750 ();
 sg13g2_fill_2 FILLER_75_756 ();
 sg13g2_fill_2 FILLER_75_812 ();
 sg13g2_fill_1 FILLER_76_48 ();
 sg13g2_fill_1 FILLER_76_131 ();
 sg13g2_fill_1 FILLER_76_150 ();
 sg13g2_fill_1 FILLER_76_160 ();
 sg13g2_fill_1 FILLER_76_186 ();
 sg13g2_fill_2 FILLER_76_221 ();
 sg13g2_fill_1 FILLER_76_223 ();
 sg13g2_fill_1 FILLER_76_239 ();
 sg13g2_fill_1 FILLER_76_269 ();
 sg13g2_fill_2 FILLER_76_306 ();
 sg13g2_fill_1 FILLER_76_334 ();
 sg13g2_fill_2 FILLER_76_346 ();
 sg13g2_fill_1 FILLER_76_348 ();
 sg13g2_fill_2 FILLER_76_422 ();
 sg13g2_fill_1 FILLER_76_459 ();
 sg13g2_fill_2 FILLER_76_546 ();
 sg13g2_fill_2 FILLER_76_635 ();
 sg13g2_fill_2 FILLER_76_679 ();
 sg13g2_fill_1 FILLER_76_716 ();
 sg13g2_fill_1 FILLER_76_722 ();
 sg13g2_fill_2 FILLER_76_735 ();
 sg13g2_fill_2 FILLER_76_757 ();
 sg13g2_fill_1 FILLER_76_759 ();
 sg13g2_fill_1 FILLER_76_765 ();
 sg13g2_fill_1 FILLER_76_785 ();
 sg13g2_fill_2 FILLER_76_815 ();
 sg13g2_fill_1 FILLER_76_827 ();
 sg13g2_fill_2 FILLER_76_833 ();
 sg13g2_fill_2 FILLER_76_848 ();
 sg13g2_fill_1 FILLER_76_850 ();
 sg13g2_fill_2 FILLER_76_860 ();
 sg13g2_fill_2 FILLER_77_108 ();
 sg13g2_fill_2 FILLER_77_255 ();
 sg13g2_fill_2 FILLER_77_266 ();
 sg13g2_fill_1 FILLER_77_268 ();
 sg13g2_fill_2 FILLER_77_274 ();
 sg13g2_fill_1 FILLER_77_280 ();
 sg13g2_fill_1 FILLER_77_304 ();
 sg13g2_fill_1 FILLER_77_338 ();
 sg13g2_fill_1 FILLER_77_347 ();
 sg13g2_fill_2 FILLER_77_381 ();
 sg13g2_fill_2 FILLER_77_440 ();
 sg13g2_fill_1 FILLER_77_510 ();
 sg13g2_fill_2 FILLER_77_624 ();
 sg13g2_fill_1 FILLER_77_657 ();
 sg13g2_fill_1 FILLER_77_736 ();
 sg13g2_fill_1 FILLER_77_742 ();
 sg13g2_fill_2 FILLER_77_851 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_27 ();
 sg13g2_fill_2 FILLER_78_65 ();
 sg13g2_fill_2 FILLER_78_140 ();
 sg13g2_fill_1 FILLER_78_142 ();
 sg13g2_fill_2 FILLER_78_148 ();
 sg13g2_fill_1 FILLER_78_150 ();
 sg13g2_fill_2 FILLER_78_181 ();
 sg13g2_fill_2 FILLER_78_199 ();
 sg13g2_fill_1 FILLER_78_224 ();
 sg13g2_fill_2 FILLER_78_238 ();
 sg13g2_fill_1 FILLER_78_240 ();
 sg13g2_fill_1 FILLER_78_263 ();
 sg13g2_fill_2 FILLER_78_274 ();
 sg13g2_fill_2 FILLER_78_306 ();
 sg13g2_fill_1 FILLER_78_395 ();
 sg13g2_fill_2 FILLER_78_579 ();
 sg13g2_fill_1 FILLER_78_604 ();
 sg13g2_fill_1 FILLER_78_628 ();
 sg13g2_fill_1 FILLER_78_645 ();
 sg13g2_fill_1 FILLER_78_660 ();
 sg13g2_fill_1 FILLER_78_707 ();
 sg13g2_fill_1 FILLER_78_731 ();
 sg13g2_fill_1 FILLER_78_741 ();
 sg13g2_fill_1 FILLER_78_784 ();
 sg13g2_fill_1 FILLER_78_815 ();
 sg13g2_fill_2 FILLER_78_826 ();
 sg13g2_fill_1 FILLER_78_828 ();
 sg13g2_fill_2 FILLER_78_834 ();
 sg13g2_fill_1 FILLER_79_81 ();
 sg13g2_fill_2 FILLER_79_91 ();
 sg13g2_fill_2 FILLER_79_128 ();
 sg13g2_fill_2 FILLER_79_147 ();
 sg13g2_fill_1 FILLER_79_187 ();
 sg13g2_fill_1 FILLER_79_206 ();
 sg13g2_fill_1 FILLER_79_271 ();
 sg13g2_fill_2 FILLER_79_285 ();
 sg13g2_fill_1 FILLER_79_287 ();
 sg13g2_fill_1 FILLER_79_314 ();
 sg13g2_fill_2 FILLER_79_341 ();
 sg13g2_fill_1 FILLER_79_402 ();
 sg13g2_fill_1 FILLER_79_436 ();
 sg13g2_fill_1 FILLER_79_463 ();
 sg13g2_fill_2 FILLER_79_482 ();
 sg13g2_fill_1 FILLER_79_487 ();
 sg13g2_fill_2 FILLER_79_508 ();
 sg13g2_fill_1 FILLER_79_568 ();
 sg13g2_fill_2 FILLER_79_764 ();
 sg13g2_fill_2 FILLER_79_854 ();
 sg13g2_fill_2 FILLER_79_860 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_121 ();
 sg13g2_fill_1 FILLER_80_183 ();
 sg13g2_fill_1 FILLER_80_236 ();
 sg13g2_fill_1 FILLER_80_250 ();
 sg13g2_fill_2 FILLER_80_300 ();
 sg13g2_fill_1 FILLER_80_302 ();
 sg13g2_fill_1 FILLER_80_319 ();
 sg13g2_fill_1 FILLER_80_361 ();
 sg13g2_fill_1 FILLER_80_372 ();
 sg13g2_fill_2 FILLER_80_429 ();
 sg13g2_fill_2 FILLER_80_503 ();
 sg13g2_fill_2 FILLER_80_536 ();
 sg13g2_fill_1 FILLER_80_564 ();
 sg13g2_fill_2 FILLER_80_609 ();
 sg13g2_fill_2 FILLER_80_624 ();
 sg13g2_fill_2 FILLER_80_665 ();
 sg13g2_fill_1 FILLER_80_681 ();
 sg13g2_fill_2 FILLER_80_712 ();
 sg13g2_fill_2 FILLER_80_771 ();
 sg13g2_fill_2 FILLER_80_799 ();
 sg13g2_fill_1 FILLER_80_810 ();
 sg13g2_fill_1 FILLER_80_841 ();
 assign uio_oe[0] = net335;
 assign uio_oe[1] = net336;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net337;
 assign uio_oe[4] = net338;
 assign uio_oe[5] = net339;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net340;
 assign uio_out[2] = net13;
 assign uio_out[6] = net14;
endmodule
