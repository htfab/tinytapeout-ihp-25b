module tt_um_izh_neuron_lite (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire params_ready_internal;
 wire spike_out_internal;
 wire \system_inst.internal_param_a[0] ;
 wire \system_inst.internal_param_a[1] ;
 wire \system_inst.internal_param_a[2] ;
 wire \system_inst.internal_param_a[3] ;
 wire \system_inst.internal_param_a[4] ;
 wire \system_inst.internal_param_a[5] ;
 wire \system_inst.internal_param_b[0] ;
 wire \system_inst.internal_param_b[1] ;
 wire \system_inst.internal_param_b[2] ;
 wire \system_inst.internal_param_b[3] ;
 wire \system_inst.internal_param_b[4] ;
 wire \system_inst.internal_param_b[5] ;
 wire \system_inst.internal_param_c[0] ;
 wire \system_inst.internal_param_c[1] ;
 wire \system_inst.internal_param_c[2] ;
 wire \system_inst.internal_param_c[3] ;
 wire \system_inst.internal_param_c[4] ;
 wire \system_inst.internal_param_c[5] ;
 wire \system_inst.internal_param_d[0] ;
 wire \system_inst.internal_param_d[1] ;
 wire \system_inst.internal_param_d[2] ;
 wire \system_inst.internal_param_d[3] ;
 wire \system_inst.internal_param_d[4] ;
 wire \system_inst.internal_param_d[5] ;
 wire \system_inst.loader.bit_count[0] ;
 wire \system_inst.loader.bit_count[1] ;
 wire \system_inst.loader.bit_count[2] ;
 wire \system_inst.loader.load_enable_prev ;
 wire \system_inst.loader.shift_reg[0] ;
 wire \system_inst.loader.shift_reg[1] ;
 wire \system_inst.loader.shift_reg[2] ;
 wire \system_inst.loader.shift_reg[3] ;
 wire \system_inst.loader.shift_reg[4] ;
 wire \system_inst.loader.state[0] ;
 wire \system_inst.loader.state[1] ;
 wire \system_inst.loader.state[2] ;
 wire \system_inst.loader.state[3] ;
 wire \system_inst.loader.state[4] ;
 wire \system_inst.loader.state[5] ;
 wire \system_inst.neuron.u[0] ;
 wire \system_inst.neuron.u[1] ;
 wire \system_inst.neuron.u[2] ;
 wire \system_inst.neuron.u[3] ;
 wire \system_inst.neuron.u[4] ;
 wire \system_inst.neuron.u[5] ;
 wire \system_inst.neuron.u[6] ;
 wire \system_inst.neuron.u[7] ;
 wire \system_inst.neuron.u[8] ;
 wire \system_inst.neuron.u[9] ;
 wire \system_inst.neuron.v[0] ;
 wire \system_inst.neuron.v[1] ;
 wire \system_inst.neuron.v[2] ;
 wire \system_inst.neuron.v[3] ;
 wire \system_inst.neuron.v[4] ;
 wire \system_inst.neuron.v[5] ;
 wire \system_inst.neuron.v[6] ;
 wire \system_inst.neuron.v[7] ;
 wire \system_inst.neuron.v[8] ;
 wire \system_inst.neuron.v[9] ;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire clknet_0_clk;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;

 sg13g2_xnor2_1 _1900_ (.Y(_0351_),
    .A(_0023_),
    .B(_0350_));
 sg13g2_nand2_1 _1901_ (.Y(_0352_),
    .A(_0345_),
    .B(_0351_));
 sg13g2_nand2_1 _1902_ (.Y(_0353_),
    .A(net365),
    .B(net377));
 sg13g2_inv_1 _1903_ (.Y(_0354_),
    .A(_0353_));
 sg13g2_xnor2_1 _1904_ (.Y(_0355_),
    .A(_0301_),
    .B(_0303_));
 sg13g2_and2_1 _1905_ (.A(_0343_),
    .B(_0355_),
    .X(_0356_));
 sg13g2_xor2_1 _1906_ (.B(_0355_),
    .A(_0343_),
    .X(_0357_));
 sg13g2_xnor2_1 _1907_ (.Y(_0358_),
    .A(_0353_),
    .B(_0357_));
 sg13g2_nor2b_1 _1908_ (.A(_0352_),
    .B_N(_0358_),
    .Y(_0359_));
 sg13g2_xnor2_1 _1909_ (.Y(_0360_),
    .A(_0352_),
    .B(_0358_));
 sg13g2_xor2_1 _1910_ (.B(_0347_),
    .A(_0346_),
    .X(_0361_));
 sg13g2_a21oi_1 _1911_ (.A1(_0360_),
    .A2(_0361_),
    .Y(_0362_),
    .B1(_0359_));
 sg13g2_a21oi_1 _1912_ (.A1(_0354_),
    .A2(_0357_),
    .Y(_0363_),
    .B1(_0356_));
 sg13g2_xnor2_1 _1913_ (.Y(_0364_),
    .A(_0993_),
    .B(_0307_));
 sg13g2_nand2b_1 _1914_ (.Y(_0365_),
    .B(_0364_),
    .A_N(_0363_));
 sg13g2_xor2_1 _1915_ (.B(_0364_),
    .A(_0363_),
    .X(_0366_));
 sg13g2_o21ai_1 _1916_ (.B1(_0331_),
    .Y(_0367_),
    .A1(_0301_),
    .A2(_0332_));
 sg13g2_and2_1 _1917_ (.A(net370),
    .B(net373),
    .X(_0368_));
 sg13g2_nand2_1 _1918_ (.Y(_0369_),
    .A(net368),
    .B(net373));
 sg13g2_xor2_1 _1919_ (.B(_0271_),
    .A(_0152_),
    .X(_0370_));
 sg13g2_nand2_1 _1920_ (.Y(_0371_),
    .A(_0368_),
    .B(_0370_));
 sg13g2_xnor2_1 _1921_ (.Y(_0372_),
    .A(_0369_),
    .B(_0370_));
 sg13g2_nand2_1 _1922_ (.Y(_0373_),
    .A(_0367_),
    .B(_0372_));
 sg13g2_xnor2_1 _1923_ (.Y(_0374_),
    .A(_0367_),
    .B(_0372_));
 sg13g2_xnor2_1 _1924_ (.Y(_0375_),
    .A(_0366_),
    .B(_0374_));
 sg13g2_nor2_1 _1925_ (.A(_0362_),
    .B(_0375_),
    .Y(_0376_));
 sg13g2_xnor2_1 _1926_ (.Y(_0377_),
    .A(_0273_),
    .B(_0348_));
 sg13g2_xor2_1 _1927_ (.B(_0375_),
    .A(_0362_),
    .X(_0378_));
 sg13g2_a21oi_1 _1928_ (.A1(_0377_),
    .A2(_0378_),
    .Y(_0379_),
    .B1(_0376_));
 sg13g2_a21oi_2 _1929_ (.B1(_0235_),
    .Y(_0380_),
    .A2(_0373_),
    .A1(_0371_));
 sg13g2_nand3_1 _1930_ (.B(_0371_),
    .C(_0373_),
    .A(_0235_),
    .Y(_0381_));
 sg13g2_nand2b_1 _1931_ (.Y(_0382_),
    .B(_0381_),
    .A_N(_0380_));
 sg13g2_o21ai_1 _1932_ (.B1(_0365_),
    .Y(_0383_),
    .A1(_0366_),
    .A2(_0374_));
 sg13g2_xnor2_1 _1933_ (.Y(_0384_),
    .A(_0311_),
    .B(_0316_));
 sg13g2_nand2b_1 _1934_ (.Y(_0385_),
    .B(_0383_),
    .A_N(_0384_));
 sg13g2_xor2_1 _1935_ (.B(_0384_),
    .A(_0383_),
    .X(_0386_));
 sg13g2_xor2_1 _1936_ (.B(_0386_),
    .A(_0382_),
    .X(_0387_));
 sg13g2_nand2b_1 _1937_ (.Y(_0388_),
    .B(_0387_),
    .A_N(_0379_));
 sg13g2_xnor2_1 _1938_ (.Y(_0389_),
    .A(_0379_),
    .B(_0387_));
 sg13g2_nand2b_1 _1939_ (.Y(_0390_),
    .B(_0389_),
    .A_N(_0349_));
 sg13g2_xnor2_1 _1940_ (.Y(_0391_),
    .A(_0349_),
    .B(_0389_));
 sg13g2_and2_1 _1941_ (.A(net372),
    .B(net375),
    .X(_0392_));
 sg13g2_nand2_1 _1942_ (.Y(_0393_),
    .A(net372),
    .B(net375));
 sg13g2_and4_1 _1943_ (.A(net366),
    .B(net367),
    .C(net379),
    .D(net384),
    .X(_0394_));
 sg13g2_a22oi_1 _1944_ (.Y(_0395_),
    .B1(net385),
    .B2(net366),
    .A2(net379),
    .A1(net367));
 sg13g2_nor2_2 _1945_ (.A(_0394_),
    .B(_0395_),
    .Y(_0396_));
 sg13g2_xnor2_1 _1946_ (.Y(_0397_),
    .A(_0393_),
    .B(_0396_));
 sg13g2_nand3_1 _1947_ (.B(net390),
    .C(_0397_),
    .A(net360),
    .Y(_0398_));
 sg13g2_xnor2_1 _1948_ (.Y(_0399_),
    .A(_0345_),
    .B(_0351_));
 sg13g2_nor2_1 _1949_ (.A(_0398_),
    .B(_0399_),
    .Y(_0400_));
 sg13g2_xor2_1 _1950_ (.B(_0399_),
    .A(_0398_),
    .X(_0401_));
 sg13g2_a21oi_1 _1951_ (.A1(_0392_),
    .A2(_0396_),
    .Y(_0402_),
    .B1(_0394_));
 sg13g2_xor2_1 _1952_ (.B(_0345_),
    .A(_0338_),
    .X(_0403_));
 sg13g2_nor2b_1 _1953_ (.A(_0402_),
    .B_N(_0403_),
    .Y(_0404_));
 sg13g2_xnor2_1 _1954_ (.Y(_0405_),
    .A(_0402_),
    .B(_0403_));
 sg13g2_a21oi_1 _1955_ (.A1(net360),
    .A2(net390),
    .Y(_0406_),
    .B1(_0394_));
 sg13g2_nor2_1 _1956_ (.A(_0395_),
    .B(_0406_),
    .Y(_0407_));
 sg13g2_xnor2_1 _1957_ (.Y(_0408_),
    .A(_0405_),
    .B(_0407_));
 sg13g2_inv_1 _1958_ (.Y(_0409_),
    .A(_0408_));
 sg13g2_a21oi_1 _1959_ (.A1(_0401_),
    .A2(_0409_),
    .Y(_0410_),
    .B1(_0400_));
 sg13g2_xnor2_1 _1960_ (.Y(_0411_),
    .A(_0360_),
    .B(_0361_));
 sg13g2_or2_1 _1961_ (.X(_0412_),
    .B(_0411_),
    .A(_0410_));
 sg13g2_xnor2_1 _1962_ (.Y(_0413_),
    .A(_0410_),
    .B(_0411_));
 sg13g2_a21o_1 _1963_ (.A2(_0407_),
    .A1(_0405_),
    .B1(_0404_),
    .X(_0414_));
 sg13g2_xnor2_1 _1964_ (.Y(_0415_),
    .A(net349),
    .B(_0414_));
 sg13g2_xnor2_1 _1965_ (.Y(_0416_),
    .A(_0354_),
    .B(_0415_));
 sg13g2_o21ai_1 _1966_ (.B1(_0412_),
    .Y(_0417_),
    .A1(_0413_),
    .A2(_0416_));
 sg13g2_xor2_1 _1967_ (.B(_0378_),
    .A(_0377_),
    .X(_0418_));
 sg13g2_nand2_1 _1968_ (.Y(_0419_),
    .A(_0417_),
    .B(_0418_));
 sg13g2_a22oi_1 _1969_ (.Y(_0420_),
    .B1(_0415_),
    .B2(_0354_),
    .A2(_0414_),
    .A1(_1004_));
 sg13g2_nor2_1 _1970_ (.A(_0417_),
    .B(_0418_),
    .Y(_0421_));
 sg13g2_xor2_1 _1971_ (.B(_0418_),
    .A(_0417_),
    .X(_0422_));
 sg13g2_o21ai_1 _1972_ (.B1(_0419_),
    .Y(_0423_),
    .A1(_0420_),
    .A2(_0421_));
 sg13g2_and2_1 _1973_ (.A(_0391_),
    .B(_0423_),
    .X(_0424_));
 sg13g2_xor2_1 _1974_ (.B(_0423_),
    .A(_0391_),
    .X(_0425_));
 sg13g2_xnor2_1 _1975_ (.Y(_0426_),
    .A(_0391_),
    .B(_0423_));
 sg13g2_a22oi_1 _1976_ (.Y(_0427_),
    .B1(net390),
    .B2(net368),
    .A2(net385),
    .A1(net371));
 sg13g2_a21oi_2 _1977_ (.B1(_0427_),
    .Y(_0428_),
    .A2(_0368_),
    .A1(_1172_));
 sg13g2_inv_1 _1978_ (.Y(_0429_),
    .A(_0428_));
 sg13g2_nand2_1 _1979_ (.Y(_0430_),
    .A(_0335_),
    .B(_0428_));
 sg13g2_nand2_1 _1980_ (.Y(_0431_),
    .A(net371),
    .B(net379));
 sg13g2_nand2_1 _1981_ (.Y(_0432_),
    .A(_1172_),
    .B(_0130_));
 sg13g2_a22oi_1 _1982_ (.Y(_0433_),
    .B1(net390),
    .B2(net363),
    .A2(net385),
    .A1(net368));
 sg13g2_a21oi_1 _1983_ (.A1(_1172_),
    .A2(_0130_),
    .Y(_0434_),
    .B1(_0433_));
 sg13g2_nand2b_1 _1984_ (.Y(_0435_),
    .B(_0434_),
    .A_N(_0431_));
 sg13g2_xnor2_1 _1985_ (.Y(_0436_),
    .A(_0431_),
    .B(_0434_));
 sg13g2_nand2_1 _1986_ (.Y(_0437_),
    .A(_0430_),
    .B(_0436_));
 sg13g2_nand2b_1 _1987_ (.Y(_0438_),
    .B(_0436_),
    .A_N(_0430_));
 sg13g2_o21ai_1 _1988_ (.B1(_0438_),
    .Y(_0439_),
    .A1(_1173_),
    .A2(_0369_));
 sg13g2_and2_1 _1989_ (.A(_0392_),
    .B(_0439_),
    .X(_0440_));
 sg13g2_mux2_1 _1990_ (.A0(_0393_),
    .A1(_0437_),
    .S(_0439_),
    .X(_0441_));
 sg13g2_a21oi_2 _1991_ (.B1(_0337_),
    .Y(_0442_),
    .A2(_0435_),
    .A1(_0432_));
 sg13g2_nand3_1 _1992_ (.B(_0432_),
    .C(_0435_),
    .A(_0337_),
    .Y(_0443_));
 sg13g2_nor2b_1 _1993_ (.A(_0442_),
    .B_N(_0443_),
    .Y(_0444_));
 sg13g2_a21oi_1 _1994_ (.A1(net359),
    .A2(net391),
    .Y(_0445_),
    .B1(_0396_));
 sg13g2_a21oi_1 _1995_ (.A1(_0392_),
    .A2(_0396_),
    .Y(_0446_),
    .B1(_0445_));
 sg13g2_and2_1 _1996_ (.A(_0398_),
    .B(_0446_),
    .X(_0447_));
 sg13g2_inv_1 _1997_ (.Y(_0448_),
    .A(_0447_));
 sg13g2_xor2_1 _1998_ (.B(_0408_),
    .A(_0401_),
    .X(_0449_));
 sg13g2_nor2_1 _1999_ (.A(_0448_),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_xnor2_1 _2000_ (.Y(_0451_),
    .A(_0447_),
    .B(_0449_));
 sg13g2_xnor2_1 _2001_ (.Y(_0452_),
    .A(_0444_),
    .B(_0451_));
 sg13g2_xor2_1 _2002_ (.B(_0452_),
    .A(_0441_),
    .X(_0453_));
 sg13g2_nand2_1 _2003_ (.Y(_0454_),
    .A(_0440_),
    .B(_0453_));
 sg13g2_o21ai_1 _2004_ (.B1(_0454_),
    .Y(_0455_),
    .A1(_0441_),
    .A2(_0452_));
 sg13g2_a21oi_1 _2005_ (.A1(_0444_),
    .A2(_0451_),
    .Y(_0456_),
    .B1(_0450_));
 sg13g2_xnor2_1 _2006_ (.Y(_0457_),
    .A(_0413_),
    .B(_0416_));
 sg13g2_nor2_1 _2007_ (.A(_0456_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_xor2_1 _2008_ (.B(_0457_),
    .A(_0456_),
    .X(_0459_));
 sg13g2_xor2_1 _2009_ (.B(_0459_),
    .A(_0442_),
    .X(_0460_));
 sg13g2_nor2_1 _2010_ (.A(_0455_),
    .B(_0460_),
    .Y(_0461_));
 sg13g2_nand2_1 _2011_ (.Y(_0462_),
    .A(net371),
    .B(net391));
 sg13g2_and4_1 _2012_ (.A(net371),
    .B(net376),
    .C(net384),
    .D(net391),
    .X(_0463_));
 sg13g2_a22oi_1 _2013_ (.Y(_0464_),
    .B1(net391),
    .B2(net372),
    .A2(net384),
    .A1(net376));
 sg13g2_nor2_1 _2014_ (.A(net380),
    .B(_0463_),
    .Y(_0465_));
 sg13g2_nor2_1 _2015_ (.A(_0464_),
    .B(_0465_),
    .Y(_0466_));
 sg13g2_nor2_1 _2016_ (.A(_0429_),
    .B(_0466_),
    .Y(_0467_));
 sg13g2_a22oi_1 _2017_ (.Y(_0468_),
    .B1(_0467_),
    .B2(net376),
    .A2(_0428_),
    .A1(_0335_));
 sg13g2_xor2_1 _2018_ (.B(_0439_),
    .A(_0437_),
    .X(_0469_));
 sg13g2_nor2_1 _2019_ (.A(_0468_),
    .B(_0469_),
    .Y(_0470_));
 sg13g2_or2_1 _2020_ (.X(_0471_),
    .B(_0428_),
    .A(_0335_));
 sg13g2_nand3_1 _2021_ (.B(_0466_),
    .C(_0471_),
    .A(_0430_),
    .Y(_0472_));
 sg13g2_nor2_1 _2022_ (.A(_0025_),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_xor2_1 _2023_ (.B(_0469_),
    .A(_0468_),
    .X(_0474_));
 sg13g2_a21oi_1 _2024_ (.A1(_0473_),
    .A2(_0474_),
    .Y(_0475_),
    .B1(_0470_));
 sg13g2_xnor2_1 _2025_ (.Y(_0476_),
    .A(_0440_),
    .B(_0453_));
 sg13g2_nor2_1 _2026_ (.A(_0475_),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_o21ai_1 _2027_ (.B1(_0026_),
    .Y(_0478_),
    .A1(_0463_),
    .A2(_0464_));
 sg13g2_or3_1 _2028_ (.A(_0026_),
    .B(_0463_),
    .C(_0464_),
    .X(_0479_));
 sg13g2_a22oi_1 _2029_ (.Y(_0480_),
    .B1(_0478_),
    .B2(_0479_),
    .A2(net384),
    .A1(net380));
 sg13g2_and4_1 _2030_ (.A(net379),
    .B(net384),
    .C(_0478_),
    .D(_0479_),
    .X(_0481_));
 sg13g2_nor3_1 _2031_ (.A(_0462_),
    .B(_0480_),
    .C(_0481_),
    .Y(_0482_));
 sg13g2_xnor2_1 _2032_ (.Y(_0483_),
    .A(_0336_),
    .B(_0466_));
 sg13g2_nand2_1 _2033_ (.Y(_0484_),
    .A(_0482_),
    .B(_0483_));
 sg13g2_xnor2_1 _2034_ (.Y(_0485_),
    .A(_0482_),
    .B(_0483_));
 sg13g2_nand2_1 _2035_ (.Y(_0486_),
    .A(net375),
    .B(_0481_));
 sg13g2_o21ai_1 _2036_ (.B1(_0486_),
    .Y(_0487_),
    .A1(_0335_),
    .A2(_0481_));
 sg13g2_o21ai_1 _2037_ (.B1(_0484_),
    .Y(_0488_),
    .A1(_0485_),
    .A2(_0487_));
 sg13g2_nand2b_1 _2038_ (.Y(_0489_),
    .B(_0472_),
    .A_N(_0467_));
 sg13g2_xnor2_1 _2039_ (.Y(_0490_),
    .A(_0757_),
    .B(_0489_));
 sg13g2_nand2_1 _2040_ (.Y(_0491_),
    .A(_0488_),
    .B(_0490_));
 sg13g2_xnor2_1 _2041_ (.Y(_0492_),
    .A(_0488_),
    .B(_0490_));
 sg13g2_o21ai_1 _2042_ (.B1(_0491_),
    .Y(_0493_),
    .A1(_0486_),
    .A2(_0492_));
 sg13g2_xor2_1 _2043_ (.B(_0474_),
    .A(_0473_),
    .X(_0494_));
 sg13g2_nand2_1 _2044_ (.Y(_0495_),
    .A(_0493_),
    .B(_0494_));
 sg13g2_nand2_1 _2045_ (.Y(_0496_),
    .A(net378),
    .B(net392));
 sg13g2_nand2_2 _2046_ (.Y(_0497_),
    .A(_1172_),
    .B(_0335_));
 sg13g2_o21ai_1 _2047_ (.B1(net382),
    .Y(_0498_),
    .A1(net387),
    .A2(_0027_));
 sg13g2_or2_1 _2048_ (.X(_0499_),
    .B(_0498_),
    .A(_0496_));
 sg13g2_o21ai_1 _2049_ (.B1(_0499_),
    .Y(_0500_),
    .A1(_0757_),
    .A2(_0779_));
 sg13g2_nand2_2 _2050_ (.Y(_0501_),
    .A(_0497_),
    .B(_0500_));
 sg13g2_mux2_1 _2051_ (.A0(_0026_),
    .A1(_0025_),
    .S(net387),
    .X(_0502_));
 sg13g2_nor2_1 _2052_ (.A(_0501_),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_xor2_1 _2053_ (.B(_0487_),
    .A(_0485_),
    .X(_0504_));
 sg13g2_inv_1 _2054_ (.Y(_0505_),
    .A(_0504_));
 sg13g2_nand2_1 _2055_ (.Y(_0506_),
    .A(_0503_),
    .B(_0504_));
 sg13g2_xor2_1 _2056_ (.B(_0504_),
    .A(_0503_),
    .X(_0507_));
 sg13g2_o21ai_1 _2057_ (.B1(_0506_),
    .Y(_0508_),
    .A1(_0497_),
    .A2(_0505_));
 sg13g2_xor2_1 _2058_ (.B(_0492_),
    .A(_0486_),
    .X(_0509_));
 sg13g2_and2_1 _2059_ (.A(_0508_),
    .B(_0509_),
    .X(_0510_));
 sg13g2_xnor2_1 _2060_ (.Y(_0511_),
    .A(_0497_),
    .B(_0507_));
 sg13g2_xor2_1 _2061_ (.B(_0502_),
    .A(_0501_),
    .X(_0512_));
 sg13g2_xnor2_1 _2062_ (.Y(_0513_),
    .A(_0501_),
    .B(_0502_));
 sg13g2_nand3_1 _2063_ (.B(net387),
    .C(net392),
    .A(net376),
    .Y(_0514_));
 sg13g2_nand2_1 _2064_ (.Y(_0515_),
    .A(_1173_),
    .B(_0496_));
 sg13g2_nand2_1 _2065_ (.Y(_0516_),
    .A(_0514_),
    .B(_0515_));
 sg13g2_nand2_1 _2066_ (.Y(_0517_),
    .A(_0757_),
    .B(_0498_));
 sg13g2_nand3_1 _2067_ (.B(_0499_),
    .C(_0517_),
    .A(net393),
    .Y(_0518_));
 sg13g2_nor2_1 _2068_ (.A(_0516_),
    .B(_0518_),
    .Y(_0519_));
 sg13g2_xnor2_1 _2069_ (.Y(_0520_),
    .A(_0512_),
    .B(_0519_));
 sg13g2_nor2_1 _2070_ (.A(_0514_),
    .B(_0520_),
    .Y(_0521_));
 sg13g2_a21oi_1 _2071_ (.A1(_0512_),
    .A2(_0519_),
    .Y(_0522_),
    .B1(_0521_));
 sg13g2_nor2b_1 _2072_ (.A(_0522_),
    .B_N(_0511_),
    .Y(_0523_));
 sg13g2_xor2_1 _2073_ (.B(_0509_),
    .A(_0508_),
    .X(_0524_));
 sg13g2_a21oi_1 _2074_ (.A1(_0523_),
    .A2(_0524_),
    .Y(_0525_),
    .B1(_0510_));
 sg13g2_xnor2_1 _2075_ (.Y(_0526_),
    .A(_0493_),
    .B(_0494_));
 sg13g2_o21ai_1 _2076_ (.B1(_0495_),
    .Y(_0527_),
    .A1(_0525_),
    .A2(_0526_));
 sg13g2_xor2_1 _2077_ (.B(_0476_),
    .A(_0475_),
    .X(_0528_));
 sg13g2_a21oi_1 _2078_ (.A1(_0527_),
    .A2(_0528_),
    .Y(_0529_),
    .B1(_0477_));
 sg13g2_a221oi_1 _2079_ (.B2(_0528_),
    .C1(_0477_),
    .B1(_0527_),
    .A1(_0455_),
    .Y(_0530_),
    .A2(_0460_));
 sg13g2_nor2_1 _2080_ (.A(_0461_),
    .B(_0530_),
    .Y(_0531_));
 sg13g2_xnor2_1 _2081_ (.Y(_0532_),
    .A(_0420_),
    .B(_0422_));
 sg13g2_a21oi_1 _2082_ (.A1(_0442_),
    .A2(_0459_),
    .Y(_0533_),
    .B1(_0458_));
 sg13g2_nor2b_1 _2083_ (.A(_0533_),
    .B_N(_0532_),
    .Y(_0534_));
 sg13g2_xor2_1 _2084_ (.B(_0533_),
    .A(_0532_),
    .X(_0535_));
 sg13g2_or3_1 _2085_ (.A(_0461_),
    .B(_0530_),
    .C(_0535_),
    .X(_0536_));
 sg13g2_nor2_1 _2086_ (.A(_0426_),
    .B(_0535_),
    .Y(_0537_));
 sg13g2_or4_2 _2087_ (.A(_0426_),
    .B(_0461_),
    .C(_0530_),
    .D(_0535_),
    .X(_0538_));
 sg13g2_and2_1 _2088_ (.A(_0425_),
    .B(_0534_),
    .X(_0539_));
 sg13g2_nand2_1 _2089_ (.Y(_0540_),
    .A(_0425_),
    .B(_0534_));
 sg13g2_a21oi_1 _2090_ (.A1(_0425_),
    .A2(_0534_),
    .Y(_0541_),
    .B1(_0424_));
 sg13g2_o21ai_1 _2091_ (.B1(_0385_),
    .Y(_0542_),
    .A1(_0382_),
    .A2(_0386_));
 sg13g2_xor2_1 _2092_ (.B(_0323_),
    .A(_0322_),
    .X(_0543_));
 sg13g2_nand2_1 _2093_ (.Y(_0544_),
    .A(_0542_),
    .B(_0543_));
 sg13g2_xor2_1 _2094_ (.B(_0543_),
    .A(_0542_),
    .X(_0545_));
 sg13g2_nand2_1 _2095_ (.Y(_0546_),
    .A(_0380_),
    .B(_0545_));
 sg13g2_xnor2_1 _2096_ (.Y(_0547_),
    .A(_0380_),
    .B(_0545_));
 sg13g2_a21oi_1 _2097_ (.A1(_0388_),
    .A2(_0390_),
    .Y(_0548_),
    .B1(_0547_));
 sg13g2_inv_1 _2098_ (.Y(_0549_),
    .A(_0548_));
 sg13g2_nand3_1 _2099_ (.B(_0390_),
    .C(_0547_),
    .A(_0388_),
    .Y(_0550_));
 sg13g2_nand2b_1 _2100_ (.Y(_0551_),
    .B(_0550_),
    .A_N(_0548_));
 sg13g2_a21o_1 _2101_ (.A2(_0541_),
    .A1(_0538_),
    .B1(_0551_),
    .X(_0552_));
 sg13g2_and2_1 _2102_ (.A(_0544_),
    .B(_0546_),
    .X(_0553_));
 sg13g2_xnor2_1 _2103_ (.Y(_0554_),
    .A(_0321_),
    .B(_0327_));
 sg13g2_or2_1 _2104_ (.X(_0555_),
    .B(_0554_),
    .A(_0553_));
 sg13g2_and2_1 _2105_ (.A(_0553_),
    .B(_0554_),
    .X(_0556_));
 sg13g2_nand2b_1 _2106_ (.Y(_0557_),
    .B(_0554_),
    .A_N(_0553_));
 sg13g2_nand3b_1 _2107_ (.B(_0546_),
    .C(_0544_),
    .Y(_0558_),
    .A_N(_0554_));
 sg13g2_a221oi_1 _2108_ (.B2(_0558_),
    .C1(_0551_),
    .B1(_0557_),
    .A1(_0538_),
    .Y(_0559_),
    .A2(_0541_));
 sg13g2_o21ai_1 _2109_ (.B1(_0555_),
    .Y(_0560_),
    .A1(_0549_),
    .A2(_0556_));
 sg13g2_xor2_1 _2110_ (.B(_0329_),
    .A(_0328_),
    .X(_0561_));
 sg13g2_o21ai_1 _2111_ (.B1(_0561_),
    .Y(_0562_),
    .A1(_0559_),
    .A2(_0560_));
 sg13g2_nand2_1 _2112_ (.Y(_0563_),
    .A(_0330_),
    .B(_0562_));
 sg13g2_nand3_1 _2113_ (.B(_0330_),
    .C(_0562_),
    .A(_0296_),
    .Y(_0564_));
 sg13g2_nand3_1 _2114_ (.B(_0297_),
    .C(_0564_),
    .A(_0268_),
    .Y(_0565_));
 sg13g2_xnor2_1 _2115_ (.Y(_0566_),
    .A(_0214_),
    .B(_0233_));
 sg13g2_a21oi_1 _2116_ (.A1(_0267_),
    .A2(_0565_),
    .Y(_0567_),
    .B1(_0566_));
 sg13g2_a21oi_1 _2117_ (.A1(_0214_),
    .A2(_0233_),
    .Y(_0568_),
    .B1(_0567_));
 sg13g2_inv_1 _2118_ (.Y(_0569_),
    .A(_0568_));
 sg13g2_o21ai_1 _2119_ (.B1(_0230_),
    .Y(_0570_),
    .A1(_0190_),
    .A2(_0232_));
 sg13g2_a21oi_1 _2120_ (.A1(_0219_),
    .A2(_0226_),
    .Y(_0571_),
    .B1(_0228_));
 sg13g2_or2_1 _2121_ (.X(_0572_),
    .B(_0223_),
    .A(_0198_));
 sg13g2_a22oi_1 _2122_ (.Y(_0573_),
    .B1(_0224_),
    .B2(_0572_),
    .A2(_0222_),
    .A1(_0199_));
 sg13g2_a22oi_1 _2123_ (.Y(_0574_),
    .B1(_0174_),
    .B2(_0221_),
    .A2(_1060_),
    .A1(\system_inst.neuron.v[8] ));
 sg13g2_xor2_1 _2124_ (.B(_0174_),
    .A(_0137_),
    .X(_0575_));
 sg13g2_xnor2_1 _2125_ (.Y(_0576_),
    .A(_0574_),
    .B(_0575_));
 sg13g2_xnor2_1 _2126_ (.Y(_0577_),
    .A(_0217_),
    .B(_0576_));
 sg13g2_xnor2_1 _2127_ (.Y(_0578_),
    .A(_0573_),
    .B(_0577_));
 sg13g2_xnor2_1 _2128_ (.Y(_0579_),
    .A(_0571_),
    .B(_0578_));
 sg13g2_xnor2_1 _2129_ (.Y(_0580_),
    .A(_0570_),
    .B(_0579_));
 sg13g2_nor2_2 _2130_ (.A(_0569_),
    .B(_0580_),
    .Y(_0581_));
 sg13g2_nand2_1 _2131_ (.Y(_0582_),
    .A(_0944_),
    .B(net8));
 sg13g2_xnor2_1 _2132_ (.Y(_0583_),
    .A(\system_inst.neuron.u[9] ),
    .B(net8));
 sg13g2_nand2_1 _2133_ (.Y(_0584_),
    .A(_0581_),
    .B(_0583_));
 sg13g2_xnor2_1 _2134_ (.Y(_0585_),
    .A(_0581_),
    .B(_0583_));
 sg13g2_nor2b_1 _2135_ (.A(net415),
    .B_N(net7),
    .Y(_0586_));
 sg13g2_xnor2_1 _2136_ (.Y(_0587_),
    .A(net415),
    .B(net7));
 sg13g2_a21oi_2 _2137_ (.B1(_0586_),
    .Y(_0588_),
    .A2(_0587_),
    .A1(net358));
 sg13g2_nor2_1 _2138_ (.A(_0585_),
    .B(_0588_),
    .Y(_0589_));
 sg13g2_xnor2_1 _2139_ (.Y(_0590_),
    .A(net415),
    .B(net9));
 sg13g2_xnor2_1 _2140_ (.Y(_0591_),
    .A(net355),
    .B(_0590_));
 sg13g2_a21oi_1 _2141_ (.A1(_0582_),
    .A2(_0584_),
    .Y(_0592_),
    .B1(_0591_));
 sg13g2_nand3_1 _2142_ (.B(_0584_),
    .C(_0591_),
    .A(_0582_),
    .Y(_0593_));
 sg13g2_nand2b_1 _2143_ (.Y(_0594_),
    .B(_0593_),
    .A_N(_0592_));
 sg13g2_xor2_1 _2144_ (.B(_0594_),
    .A(_0581_),
    .X(_0595_));
 sg13g2_or3_1 _2145_ (.A(_0585_),
    .B(_0588_),
    .C(_0595_),
    .X(_0596_));
 sg13g2_a21oi_1 _2146_ (.A1(_0581_),
    .A2(_0593_),
    .Y(_0597_),
    .B1(_0592_));
 sg13g2_or3_1 _2147_ (.A(net355),
    .B(_0944_),
    .C(net9),
    .X(_0598_));
 sg13g2_nand3_1 _2148_ (.B(_0944_),
    .C(net9),
    .A(net355),
    .Y(_0599_));
 sg13g2_nand2_1 _2149_ (.Y(_0600_),
    .A(_0598_),
    .B(_0599_));
 sg13g2_mux2_1 _2150_ (.A0(_0600_),
    .A1(_0599_),
    .S(_0581_),
    .X(_0601_));
 sg13g2_xnor2_1 _2151_ (.Y(_0602_),
    .A(_0597_),
    .B(_0601_));
 sg13g2_nand2_1 _2152_ (.Y(_0603_),
    .A(_0596_),
    .B(_0602_));
 sg13g2_xor2_1 _2153_ (.B(_0595_),
    .A(_0589_),
    .X(_0604_));
 sg13g2_nor2b_1 _2154_ (.A(net415),
    .B_N(net6),
    .Y(_0605_));
 sg13g2_xnor2_1 _2155_ (.Y(_0606_),
    .A(net415),
    .B(net6));
 sg13g2_a21oi_1 _2156_ (.A1(net362),
    .A2(_0606_),
    .Y(_0607_),
    .B1(_0605_));
 sg13g2_xnor2_1 _2157_ (.Y(_0608_),
    .A(net358),
    .B(_0587_));
 sg13g2_nor2_1 _2158_ (.A(_0607_),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_xor2_1 _2159_ (.B(_0608_),
    .A(_0607_),
    .X(_0610_));
 sg13g2_xor2_1 _2160_ (.B(_0580_),
    .A(_0568_),
    .X(_0611_));
 sg13g2_inv_1 _2161_ (.Y(_0612_),
    .A(_0611_));
 sg13g2_nand3_1 _2162_ (.B(_0565_),
    .C(_0566_),
    .A(_0267_),
    .Y(_0613_));
 sg13g2_nand2b_2 _2163_ (.Y(_0614_),
    .B(_0613_),
    .A_N(_0567_));
 sg13g2_a21o_1 _2164_ (.A2(_0564_),
    .A1(_0297_),
    .B1(_0268_),
    .X(_0615_));
 sg13g2_nand2_1 _2165_ (.Y(_0616_),
    .A(_0565_),
    .B(_0615_));
 sg13g2_xor2_1 _2166_ (.B(_0616_),
    .A(_0611_),
    .X(_0617_));
 sg13g2_and2_1 _2167_ (.A(_0296_),
    .B(_0297_),
    .X(_0618_));
 sg13g2_xnor2_1 _2168_ (.Y(_0619_),
    .A(_0563_),
    .B(_0618_));
 sg13g2_nor2_1 _2169_ (.A(_0614_),
    .B(_0619_),
    .Y(_0620_));
 sg13g2_nor4_1 _2170_ (.A(_0581_),
    .B(_0614_),
    .C(_0617_),
    .D(_0619_),
    .Y(_0621_));
 sg13g2_and4_1 _2171_ (.A(_0549_),
    .B(_0552_),
    .C(_0557_),
    .D(_0558_),
    .X(_0622_));
 sg13g2_a22oi_1 _2172_ (.Y(_0623_),
    .B1(_0557_),
    .B2(_0558_),
    .A2(_0552_),
    .A1(_0549_));
 sg13g2_or2_1 _2173_ (.X(_0624_),
    .B(_0623_),
    .A(_0622_));
 sg13g2_or2_1 _2174_ (.X(_0625_),
    .B(_0624_),
    .A(_0619_));
 sg13g2_or3_1 _2175_ (.A(_0559_),
    .B(_0560_),
    .C(_0561_),
    .X(_0626_));
 sg13g2_and2_2 _2176_ (.A(_0562_),
    .B(_0626_),
    .X(_0627_));
 sg13g2_and3_2 _2177_ (.X(_0628_),
    .A(_0565_),
    .B(_0615_),
    .C(_0627_));
 sg13g2_a21oi_2 _2178_ (.B1(_0627_),
    .Y(_0629_),
    .A2(_0615_),
    .A1(_0565_));
 sg13g2_or2_1 _2179_ (.X(_0630_),
    .B(_0629_),
    .A(_0628_));
 sg13g2_nor3_2 _2180_ (.A(_0625_),
    .B(_0628_),
    .C(_0629_),
    .Y(_0631_));
 sg13g2_xor2_1 _2181_ (.B(_0619_),
    .A(_0614_),
    .X(_0632_));
 sg13g2_nand2_1 _2182_ (.Y(_0633_),
    .A(_0631_),
    .B(_0632_));
 sg13g2_nand3_1 _2183_ (.B(_0541_),
    .C(_0551_),
    .A(_0538_),
    .Y(_0634_));
 sg13g2_nand2_2 _2184_ (.Y(_0635_),
    .A(_0552_),
    .B(_0634_));
 sg13g2_and3_1 _2185_ (.X(_0636_),
    .A(_0552_),
    .B(_0627_),
    .C(_0634_));
 sg13g2_nand2_1 _2186_ (.Y(_0637_),
    .A(_0619_),
    .B(_0624_));
 sg13g2_xnor2_1 _2187_ (.Y(_0638_),
    .A(_0619_),
    .B(_0624_));
 sg13g2_nand3_1 _2188_ (.B(_0636_),
    .C(_0637_),
    .A(_0625_),
    .Y(_0639_));
 sg13g2_o21ai_1 _2189_ (.B1(_0625_),
    .Y(_0640_),
    .A1(_0628_),
    .A2(_0629_));
 sg13g2_nand2b_1 _2190_ (.Y(_0641_),
    .B(_0640_),
    .A_N(_0631_));
 sg13g2_nor2_1 _2191_ (.A(_0639_),
    .B(_0641_),
    .Y(_0642_));
 sg13g2_nor2_1 _2192_ (.A(_0425_),
    .B(_0534_),
    .Y(_0643_));
 sg13g2_nand2_1 _2193_ (.Y(_0644_),
    .A(_0536_),
    .B(_0643_));
 sg13g2_a221oi_1 _2194_ (.B2(_0536_),
    .C1(_0539_),
    .B1(_0643_),
    .A1(_0531_),
    .Y(_0645_),
    .A2(_0537_));
 sg13g2_nand3_1 _2195_ (.B(_0540_),
    .C(_0644_),
    .A(_0538_),
    .Y(_0646_));
 sg13g2_nor2_1 _2196_ (.A(_0624_),
    .B(_0646_),
    .Y(_0647_));
 sg13g2_or3_1 _2197_ (.A(_0622_),
    .B(_0623_),
    .C(_0646_),
    .X(_0648_));
 sg13g2_xnor2_1 _2198_ (.Y(_0649_),
    .A(_0627_),
    .B(_0635_));
 sg13g2_and2_1 _2199_ (.A(_0647_),
    .B(_0649_),
    .X(_0650_));
 sg13g2_xnor2_1 _2200_ (.Y(_0651_),
    .A(_0636_),
    .B(_0638_));
 sg13g2_nor2_1 _2201_ (.A(_0650_),
    .B(_0651_),
    .Y(_0652_));
 sg13g2_xor2_1 _2202_ (.B(_0460_),
    .A(_0455_),
    .X(_0653_));
 sg13g2_xnor2_1 _2203_ (.Y(_0654_),
    .A(_0529_),
    .B(_0653_));
 sg13g2_nand2_1 _2204_ (.Y(_0655_),
    .A(_0645_),
    .B(_0654_));
 sg13g2_xor2_1 _2205_ (.B(_0535_),
    .A(_0531_),
    .X(_0656_));
 sg13g2_nor2_1 _2206_ (.A(_0635_),
    .B(_0656_),
    .Y(_0657_));
 sg13g2_xor2_1 _2207_ (.B(_0656_),
    .A(_0635_),
    .X(_0658_));
 sg13g2_nor2b_1 _2208_ (.A(_0655_),
    .B_N(_0658_),
    .Y(_0659_));
 sg13g2_nand2b_1 _2209_ (.Y(_0660_),
    .B(_0658_),
    .A_N(_0655_));
 sg13g2_xor2_1 _2210_ (.B(_0658_),
    .A(_0655_),
    .X(_0661_));
 sg13g2_xnor2_1 _2211_ (.Y(_0662_),
    .A(_0527_),
    .B(_0528_));
 sg13g2_nor2_1 _2212_ (.A(_0656_),
    .B(_0662_),
    .Y(_0663_));
 sg13g2_xnor2_1 _2213_ (.Y(_0664_),
    .A(_0645_),
    .B(_0654_));
 sg13g2_or3_2 _2214_ (.A(_0656_),
    .B(_0662_),
    .C(_0664_),
    .X(_0665_));
 sg13g2_nor2_1 _2215_ (.A(_0661_),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_o21ai_1 _2216_ (.B1(_0660_),
    .Y(_0667_),
    .A1(_0661_),
    .A2(_0665_));
 sg13g2_o21ai_1 _2217_ (.B1(_0646_),
    .Y(_0668_),
    .A1(_0622_),
    .A2(_0623_));
 sg13g2_nand3_1 _2218_ (.B(_0657_),
    .C(_0668_),
    .A(_0648_),
    .Y(_0669_));
 sg13g2_a21o_1 _2219_ (.A2(_0668_),
    .A1(_0648_),
    .B1(_0657_),
    .X(_0670_));
 sg13g2_and3_1 _2220_ (.X(_0671_),
    .A(_0667_),
    .B(_0669_),
    .C(_0670_));
 sg13g2_xor2_1 _2221_ (.B(_0665_),
    .A(_0661_),
    .X(_0672_));
 sg13g2_xnor2_1 _2222_ (.Y(_0673_),
    .A(_0661_),
    .B(_0665_));
 sg13g2_xnor2_1 _2223_ (.Y(_0674_),
    .A(_0656_),
    .B(_0662_));
 sg13g2_xnor2_1 _2224_ (.Y(_0675_),
    .A(_0525_),
    .B(_0526_));
 sg13g2_nand2b_1 _2225_ (.Y(_0676_),
    .B(_0654_),
    .A_N(_0675_));
 sg13g2_or2_1 _2226_ (.X(_0677_),
    .B(_0676_),
    .A(_0674_));
 sg13g2_xor2_1 _2227_ (.B(_0664_),
    .A(_0663_),
    .X(_0678_));
 sg13g2_nor2_1 _2228_ (.A(_0677_),
    .B(_0678_),
    .Y(_0679_));
 sg13g2_xnor2_1 _2229_ (.Y(_0680_),
    .A(_0514_),
    .B(_0520_));
 sg13g2_xor2_1 _2230_ (.B(_0522_),
    .A(_0511_),
    .X(_0681_));
 sg13g2_and2_1 _2231_ (.A(_0680_),
    .B(_0681_),
    .X(_0682_));
 sg13g2_xor2_1 _2232_ (.B(_0524_),
    .A(_0523_),
    .X(_0683_));
 sg13g2_inv_1 _2233_ (.Y(_0684_),
    .A(_0683_));
 sg13g2_o21ai_1 _2234_ (.B1(_0684_),
    .Y(_0685_),
    .A1(_0662_),
    .A2(_0682_));
 sg13g2_nand2b_1 _2235_ (.Y(_0686_),
    .B(_0675_),
    .A_N(_0654_));
 sg13g2_xor2_1 _2236_ (.B(_0518_),
    .A(_0516_),
    .X(_0687_));
 sg13g2_nor3_1 _2237_ (.A(_0779_),
    .B(net393),
    .C(_0513_),
    .Y(_0688_));
 sg13g2_nor2_1 _2238_ (.A(_0687_),
    .B(_0688_),
    .Y(_0689_));
 sg13g2_a21oi_1 _2239_ (.A1(_0675_),
    .A2(_0689_),
    .Y(_0690_),
    .B1(_0681_));
 sg13g2_nor2_1 _2240_ (.A(_0680_),
    .B(_0684_),
    .Y(_0691_));
 sg13g2_nor2b_1 _2241_ (.A(_0524_),
    .B_N(_0680_),
    .Y(_0692_));
 sg13g2_o21ai_1 _2242_ (.B1(_0675_),
    .Y(_0693_),
    .A1(_0681_),
    .A2(_0692_));
 sg13g2_o21ai_1 _2243_ (.B1(_0693_),
    .Y(_0694_),
    .A1(_0690_),
    .A2(_0691_));
 sg13g2_o21ai_1 _2244_ (.B1(_0694_),
    .Y(_0695_),
    .A1(_0662_),
    .A2(_0684_));
 sg13g2_nand4_1 _2245_ (.B(_0685_),
    .C(_0686_),
    .A(_0676_),
    .Y(_0696_),
    .D(_0695_));
 sg13g2_nor2_1 _2246_ (.A(_0674_),
    .B(_0696_),
    .Y(_0697_));
 sg13g2_or2_1 _2247_ (.X(_0698_),
    .B(_0696_),
    .A(_0674_));
 sg13g2_xor2_1 _2248_ (.B(_0678_),
    .A(_0677_),
    .X(_0699_));
 sg13g2_a21oi_1 _2249_ (.A1(_0697_),
    .A2(_0699_),
    .Y(_0700_),
    .B1(_0679_));
 sg13g2_a21o_1 _2250_ (.A2(_0699_),
    .A1(_0697_),
    .B1(_0679_),
    .X(_0701_));
 sg13g2_a21oi_1 _2251_ (.A1(_0669_),
    .A2(_0670_),
    .Y(_0702_),
    .B1(_0659_));
 sg13g2_and3_1 _2252_ (.X(_0703_),
    .A(_0648_),
    .B(_0659_),
    .C(_0668_));
 sg13g2_or2_1 _2253_ (.X(_0704_),
    .B(_0703_),
    .A(_0702_));
 sg13g2_nor4_1 _2254_ (.A(_0673_),
    .B(_0700_),
    .C(_0702_),
    .D(_0703_),
    .Y(_0705_));
 sg13g2_or2_1 _2255_ (.X(_0706_),
    .B(_0705_),
    .A(_0671_));
 sg13g2_xnor2_1 _2256_ (.Y(_0707_),
    .A(_0647_),
    .B(_0649_));
 sg13g2_nor2_1 _2257_ (.A(_0669_),
    .B(_0707_),
    .Y(_0708_));
 sg13g2_xor2_1 _2258_ (.B(_0707_),
    .A(_0669_),
    .X(_0709_));
 sg13g2_o21ai_1 _2259_ (.B1(_0709_),
    .Y(_0710_),
    .A1(_0671_),
    .A2(_0705_));
 sg13g2_a21oi_1 _2260_ (.A1(_0650_),
    .A2(_0651_),
    .Y(_0711_),
    .B1(_0708_));
 sg13g2_a21oi_1 _2261_ (.A1(_0710_),
    .A2(_0711_),
    .Y(_0712_),
    .B1(_0652_));
 sg13g2_nand3b_1 _2262_ (.B(_0639_),
    .C(_0640_),
    .Y(_0714_),
    .A_N(_0631_));
 sg13g2_nand4_1 _2263_ (.B(_0630_),
    .C(_0636_),
    .A(_0625_),
    .Y(_0715_),
    .D(_0637_));
 sg13g2_nand2_1 _2264_ (.Y(_0716_),
    .A(_0714_),
    .B(_0715_));
 sg13g2_a221oi_1 _2265_ (.B2(_0715_),
    .C1(_0652_),
    .B1(_0714_),
    .A1(_0710_),
    .Y(_0717_),
    .A2(_0711_));
 sg13g2_nor2_1 _2266_ (.A(_0628_),
    .B(_0631_),
    .Y(_0718_));
 sg13g2_xnor2_1 _2267_ (.Y(_0719_),
    .A(_0632_),
    .B(_0718_));
 sg13g2_o21ai_1 _2268_ (.B1(_0719_),
    .Y(_0720_),
    .A1(_0642_),
    .A2(_0717_));
 sg13g2_a21oi_1 _2269_ (.A1(_0628_),
    .A2(_0632_),
    .Y(_0721_),
    .B1(_0620_));
 sg13g2_xnor2_1 _2270_ (.Y(_0722_),
    .A(_0617_),
    .B(_0721_));
 sg13g2_a21oi_1 _2271_ (.A1(_0633_),
    .A2(_0720_),
    .Y(_0723_),
    .B1(_0722_));
 sg13g2_and3_1 _2272_ (.X(_0725_),
    .A(_0612_),
    .B(_0628_),
    .C(_0632_));
 sg13g2_nor2_1 _2273_ (.A(_0723_),
    .B(_0725_),
    .Y(_0726_));
 sg13g2_nor3_1 _2274_ (.A(_0621_),
    .B(_0723_),
    .C(_0725_),
    .Y(_0727_));
 sg13g2_o21ai_1 _2275_ (.B1(_0612_),
    .Y(_0728_),
    .A1(_0614_),
    .A2(_0727_));
 sg13g2_xnor2_1 _2276_ (.Y(_0729_),
    .A(_0024_),
    .B(_0728_));
 sg13g2_a21oi_1 _2277_ (.A1(_0610_),
    .A2(_0729_),
    .Y(_0730_),
    .B1(_0609_));
 sg13g2_xnor2_1 _2278_ (.Y(_0731_),
    .A(_0585_),
    .B(_0588_));
 sg13g2_nand2_1 _2279_ (.Y(_0732_),
    .A(net355),
    .B(_0728_));
 sg13g2_xor2_1 _2280_ (.B(_0731_),
    .A(_0730_),
    .X(_0733_));
 sg13g2_nand2b_1 _2281_ (.Y(_0734_),
    .B(_0733_),
    .A_N(_0732_));
 sg13g2_o21ai_1 _2282_ (.B1(_0734_),
    .Y(_0736_),
    .A1(_0730_),
    .A2(_0731_));
 sg13g2_nor2b_1 _2283_ (.A(_0604_),
    .B_N(_0736_),
    .Y(_0737_));
 sg13g2_xor2_1 _2284_ (.B(_0736_),
    .A(_0604_),
    .X(_0738_));
 sg13g2_nor2b_1 _2285_ (.A(\system_inst.neuron.u[6] ),
    .B_N(net3),
    .Y(_0739_));
 sg13g2_xnor2_1 _2286_ (.Y(_0740_),
    .A(\system_inst.neuron.u[6] ),
    .B(net3));
 sg13g2_a21oi_1 _2287_ (.A1(net374),
    .A2(_0740_),
    .Y(_0741_),
    .B1(_0739_));
 sg13g2_nor2_1 _2288_ (.A(_0954_),
    .B(net4),
    .Y(_0742_));
 sg13g2_xnor2_1 _2289_ (.Y(_0743_),
    .A(\system_inst.neuron.u[7] ),
    .B(net4));
 sg13g2_nor2_1 _2290_ (.A(_0741_),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_nand2_1 _2291_ (.Y(_0745_),
    .A(_0741_),
    .B(_0743_));
 sg13g2_nand2b_1 _2292_ (.Y(_0747_),
    .B(_0745_),
    .A_N(_0744_));
 sg13g2_nor2_1 _2293_ (.A(net361),
    .B(net370),
    .Y(_0748_));
 sg13g2_nor2_1 _2294_ (.A(_0120_),
    .B(_0748_),
    .Y(_0749_));
 sg13g2_or3_1 _2295_ (.A(_0642_),
    .B(_0717_),
    .C(_0719_),
    .X(_0750_));
 sg13g2_nand2_1 _2296_ (.Y(_0751_),
    .A(_0720_),
    .B(_0750_));
 sg13g2_xnor2_1 _2297_ (.Y(_0752_),
    .A(_0749_),
    .B(_0751_));
 sg13g2_a21oi_1 _2298_ (.A1(_0745_),
    .A2(_0752_),
    .Y(_0753_),
    .B1(_0744_));
 sg13g2_nor2b_1 _2299_ (.A(net5),
    .B_N(\system_inst.neuron.u[8] ),
    .Y(_0754_));
 sg13g2_xnor2_1 _2300_ (.Y(_0755_),
    .A(\system_inst.neuron.u[8] ),
    .B(net5));
 sg13g2_nor2_1 _2301_ (.A(_0742_),
    .B(_0755_),
    .Y(_0756_));
 sg13g2_xor2_1 _2302_ (.B(_0755_),
    .A(_0742_),
    .X(_0758_));
 sg13g2_nand3_1 _2303_ (.B(_0720_),
    .C(_0722_),
    .A(_0633_),
    .Y(_0759_));
 sg13g2_nor2b_1 _2304_ (.A(_0723_),
    .B_N(_0759_),
    .Y(_0760_));
 sg13g2_nand2_1 _2305_ (.Y(_0761_),
    .A(_1067_),
    .B(_0760_));
 sg13g2_xor2_1 _2306_ (.B(_0760_),
    .A(_1067_),
    .X(_0762_));
 sg13g2_xnor2_1 _2307_ (.Y(_0763_),
    .A(_0758_),
    .B(_0762_));
 sg13g2_nor2_1 _2308_ (.A(_0753_),
    .B(_0763_),
    .Y(_0764_));
 sg13g2_o21ai_1 _2309_ (.B1(_0119_),
    .Y(_0765_),
    .A1(_0748_),
    .A2(_0751_));
 sg13g2_xor2_1 _2310_ (.B(_0763_),
    .A(_0753_),
    .X(_0766_));
 sg13g2_a21oi_1 _2311_ (.A1(_0765_),
    .A2(_0766_),
    .Y(_0767_),
    .B1(_0764_));
 sg13g2_nand2_1 _2312_ (.Y(_0769_),
    .A(_1061_),
    .B(_0761_));
 sg13g2_a21oi_1 _2313_ (.A1(_0758_),
    .A2(_0762_),
    .Y(_0770_),
    .B1(_0756_));
 sg13g2_xnor2_1 _2314_ (.Y(_0771_),
    .A(net362),
    .B(_0606_));
 sg13g2_nor2_1 _2315_ (.A(_0754_),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_xor2_1 _2316_ (.B(_0771_),
    .A(_0754_),
    .X(_0773_));
 sg13g2_nor2_1 _2317_ (.A(_0614_),
    .B(_0621_),
    .Y(_0774_));
 sg13g2_xnor2_1 _2318_ (.Y(_0775_),
    .A(_0726_),
    .B(_0774_));
 sg13g2_xnor2_1 _2319_ (.Y(_0776_),
    .A(_0024_),
    .B(_0775_));
 sg13g2_xnor2_1 _2320_ (.Y(_0777_),
    .A(_0773_),
    .B(_0776_));
 sg13g2_nor2_1 _2321_ (.A(_0770_),
    .B(_0777_),
    .Y(_0778_));
 sg13g2_xor2_1 _2322_ (.B(_0777_),
    .A(_0770_),
    .X(_0780_));
 sg13g2_xnor2_1 _2323_ (.Y(_0781_),
    .A(_0769_),
    .B(_0780_));
 sg13g2_nor2_1 _2324_ (.A(_0767_),
    .B(_0781_),
    .Y(_0782_));
 sg13g2_nor2b_1 _2325_ (.A(net416),
    .B_N(net2),
    .Y(_0783_));
 sg13g2_xnor2_1 _2326_ (.Y(_0784_),
    .A(net416),
    .B(net2));
 sg13g2_a21oi_1 _2327_ (.A1(\system_inst.neuron.v[3] ),
    .A2(_0784_),
    .Y(_0785_),
    .B1(_0783_));
 sg13g2_xnor2_1 _2328_ (.Y(_0786_),
    .A(net374),
    .B(_0740_));
 sg13g2_nor2_1 _2329_ (.A(_0785_),
    .B(_0786_),
    .Y(_0787_));
 sg13g2_xor2_1 _2330_ (.B(_0786_),
    .A(_0785_),
    .X(_0788_));
 sg13g2_xor2_1 _2331_ (.B(_0716_),
    .A(_0712_),
    .X(_0789_));
 sg13g2_xnor2_1 _2332_ (.Y(_0791_),
    .A(_0021_),
    .B(_0789_));
 sg13g2_a21oi_1 _2333_ (.A1(_0788_),
    .A2(_0791_),
    .Y(_0792_),
    .B1(_0787_));
 sg13g2_xnor2_1 _2334_ (.Y(_0793_),
    .A(_0747_),
    .B(_0752_));
 sg13g2_nand2b_1 _2335_ (.Y(_0794_),
    .B(_0793_),
    .A_N(_0792_));
 sg13g2_nand2_1 _2336_ (.Y(_0795_),
    .A(net364),
    .B(_0789_));
 sg13g2_xnor2_1 _2337_ (.Y(_0796_),
    .A(_0792_),
    .B(_0793_));
 sg13g2_nand2b_1 _2338_ (.Y(_0797_),
    .B(_0796_),
    .A_N(_0795_));
 sg13g2_nand2_1 _2339_ (.Y(_0798_),
    .A(_0794_),
    .B(_0797_));
 sg13g2_xnor2_1 _2340_ (.Y(_0799_),
    .A(_0765_),
    .B(_0766_));
 sg13g2_nand2b_1 _2341_ (.Y(_0800_),
    .B(_0798_),
    .A_N(_0799_));
 sg13g2_nor2_1 _2342_ (.A(_0768_),
    .B(\system_inst.neuron.u[4] ),
    .Y(_0802_));
 sg13g2_xnor2_1 _2343_ (.Y(_0803_),
    .A(net382),
    .B(\system_inst.neuron.u[4] ));
 sg13g2_a21oi_1 _2344_ (.A1(\system_inst.neuron.v[4] ),
    .A2(_0803_),
    .Y(_0804_),
    .B1(_0802_));
 sg13g2_xnor2_1 _2345_ (.Y(_0805_),
    .A(net378),
    .B(_0784_));
 sg13g2_nor2_1 _2346_ (.A(_0804_),
    .B(_0805_),
    .Y(_0806_));
 sg13g2_nand2_1 _2347_ (.Y(_0807_),
    .A(_0804_),
    .B(_0805_));
 sg13g2_nand2b_1 _2348_ (.Y(_0808_),
    .B(_0807_),
    .A_N(_0806_));
 sg13g2_xor2_1 _2349_ (.B(_0651_),
    .A(_0650_),
    .X(_0809_));
 sg13g2_nor2b_1 _2350_ (.A(_0708_),
    .B_N(_0710_),
    .Y(_0810_));
 sg13g2_xnor2_1 _2351_ (.Y(_0811_),
    .A(_0809_),
    .B(_0810_));
 sg13g2_xnor2_1 _2352_ (.Y(_0813_),
    .A(_0022_),
    .B(_0811_));
 sg13g2_a21oi_1 _2353_ (.A1(_0807_),
    .A2(_0813_),
    .Y(_0814_),
    .B1(_0806_));
 sg13g2_xnor2_1 _2354_ (.Y(_0815_),
    .A(_0788_),
    .B(_0791_));
 sg13g2_nand2_1 _2355_ (.Y(_0816_),
    .A(net370),
    .B(_0811_));
 sg13g2_xor2_1 _2356_ (.B(_0815_),
    .A(_0814_),
    .X(_0817_));
 sg13g2_nand2b_1 _2357_ (.Y(_0818_),
    .B(_0817_),
    .A_N(_0816_));
 sg13g2_o21ai_1 _2358_ (.B1(_0818_),
    .Y(_0819_),
    .A1(_0814_),
    .A2(_0815_));
 sg13g2_xnor2_1 _2359_ (.Y(_0820_),
    .A(_0795_),
    .B(_0796_));
 sg13g2_and2_1 _2360_ (.A(_0819_),
    .B(_0820_),
    .X(_0821_));
 sg13g2_xnor2_1 _2361_ (.Y(_0822_),
    .A(_0808_),
    .B(_0813_));
 sg13g2_nor2_1 _2362_ (.A(_0779_),
    .B(\system_inst.neuron.u[3] ),
    .Y(_0824_));
 sg13g2_xnor2_1 _2363_ (.Y(_0825_),
    .A(net388),
    .B(\system_inst.neuron.u[3] ));
 sg13g2_a21oi_2 _2364_ (.B1(_0824_),
    .Y(_0826_),
    .A2(_0825_),
    .A1(net378));
 sg13g2_xnor2_1 _2365_ (.Y(_0827_),
    .A(net374),
    .B(_0803_));
 sg13g2_xnor2_1 _2366_ (.Y(_0828_),
    .A(_0706_),
    .B(_0709_));
 sg13g2_xor2_1 _2367_ (.B(_0827_),
    .A(_0826_),
    .X(_0829_));
 sg13g2_nand2b_1 _2368_ (.Y(_0830_),
    .B(_0829_),
    .A_N(_0828_));
 sg13g2_o21ai_1 _2369_ (.B1(_0830_),
    .Y(_0831_),
    .A1(_0826_),
    .A2(_0827_));
 sg13g2_nand2_1 _2370_ (.Y(_0832_),
    .A(_0822_),
    .B(_0831_));
 sg13g2_xnor2_1 _2371_ (.Y(_0833_),
    .A(_0816_),
    .B(_0817_));
 sg13g2_nor2b_1 _2372_ (.A(_0832_),
    .B_N(_0833_),
    .Y(_0835_));
 sg13g2_xnor2_1 _2373_ (.Y(_0836_),
    .A(_0828_),
    .B(_0829_));
 sg13g2_nor2b_1 _2374_ (.A(\system_inst.neuron.u[2] ),
    .B_N(net393),
    .Y(_0837_));
 sg13g2_xnor2_1 _2375_ (.Y(_0838_),
    .A(net393),
    .B(\system_inst.neuron.u[2] ));
 sg13g2_a21oi_1 _2376_ (.A1(net382),
    .A2(_0838_),
    .Y(_0839_),
    .B1(_0837_));
 sg13g2_xnor2_1 _2377_ (.Y(_0840_),
    .A(net378),
    .B(_0825_));
 sg13g2_nor2_1 _2378_ (.A(_0839_),
    .B(_0840_),
    .Y(_0841_));
 sg13g2_xor2_1 _2379_ (.B(_0840_),
    .A(_0839_),
    .X(_0842_));
 sg13g2_a21oi_1 _2380_ (.A1(_0672_),
    .A2(_0701_),
    .Y(_0843_),
    .B1(_0666_));
 sg13g2_xor2_1 _2381_ (.B(_0843_),
    .A(_0704_),
    .X(_0844_));
 sg13g2_a21oi_1 _2382_ (.A1(_0842_),
    .A2(_0844_),
    .Y(_0846_),
    .B1(_0841_));
 sg13g2_nor2b_1 _2383_ (.A(_0846_),
    .B_N(_0836_),
    .Y(_0847_));
 sg13g2_xor2_1 _2384_ (.B(_0831_),
    .A(_0822_),
    .X(_0848_));
 sg13g2_and2_1 _2385_ (.A(_0847_),
    .B(_0848_),
    .X(_0849_));
 sg13g2_xnor2_1 _2386_ (.Y(_0850_),
    .A(_0842_),
    .B(_0844_));
 sg13g2_nor2_1 _2387_ (.A(_0779_),
    .B(\system_inst.neuron.u[1] ),
    .Y(_0851_));
 sg13g2_xnor2_1 _2388_ (.Y(_0852_),
    .A(net388),
    .B(\system_inst.neuron.u[1] ));
 sg13g2_xnor2_1 _2389_ (.Y(_0853_),
    .A(_0698_),
    .B(_0699_));
 sg13g2_a21oi_1 _2390_ (.A1(_0852_),
    .A2(_0853_),
    .Y(_0854_),
    .B1(_0851_));
 sg13g2_xnor2_1 _2391_ (.Y(_0855_),
    .A(net382),
    .B(_0838_));
 sg13g2_nor2_1 _2392_ (.A(_0854_),
    .B(_0855_),
    .Y(_0857_));
 sg13g2_xnor2_1 _2393_ (.Y(_0858_),
    .A(_0672_),
    .B(_0700_));
 sg13g2_xor2_1 _2394_ (.B(_0855_),
    .A(_0854_),
    .X(_0859_));
 sg13g2_a21oi_1 _2395_ (.A1(_0858_),
    .A2(_0859_),
    .Y(_0860_),
    .B1(_0857_));
 sg13g2_nor2_1 _2396_ (.A(_0850_),
    .B(_0860_),
    .Y(_0861_));
 sg13g2_inv_1 _2397_ (.Y(_0862_),
    .A(_0861_));
 sg13g2_xor2_1 _2398_ (.B(_0846_),
    .A(_0836_),
    .X(_0863_));
 sg13g2_or2_1 _2399_ (.X(_0864_),
    .B(_0863_),
    .A(_0862_));
 sg13g2_xnor2_1 _2400_ (.Y(_0865_),
    .A(_0850_),
    .B(_0860_));
 sg13g2_xnor2_1 _2401_ (.Y(_0866_),
    .A(_0852_),
    .B(_0853_));
 sg13g2_nor2b_1 _2402_ (.A(net393),
    .B_N(\system_inst.neuron.u[0] ),
    .Y(_0868_));
 sg13g2_nor2_1 _2403_ (.A(_0866_),
    .B(_0868_),
    .Y(_0869_));
 sg13g2_xnor2_1 _2404_ (.Y(_0870_),
    .A(_0858_),
    .B(_0859_));
 sg13g2_or3_1 _2405_ (.A(_0866_),
    .B(_0868_),
    .C(_0870_),
    .X(_0871_));
 sg13g2_nor2_1 _2406_ (.A(_0865_),
    .B(_0871_),
    .Y(_0872_));
 sg13g2_xor2_1 _2407_ (.B(_0868_),
    .A(_0866_),
    .X(_0873_));
 sg13g2_xor2_1 _2408_ (.B(\system_inst.neuron.u[0] ),
    .A(net392),
    .X(_0874_));
 sg13g2_nand3_1 _2409_ (.B(_0676_),
    .C(_0696_),
    .A(_0674_),
    .Y(_0875_));
 sg13g2_and4_1 _2410_ (.A(_0677_),
    .B(_0698_),
    .C(_0874_),
    .D(_0875_),
    .X(_0876_));
 sg13g2_nand2_1 _2411_ (.Y(_0877_),
    .A(_0873_),
    .B(_0876_));
 sg13g2_nor2_1 _2412_ (.A(_0870_),
    .B(_0877_),
    .Y(_0879_));
 sg13g2_xor2_1 _2413_ (.B(_0871_),
    .A(_0865_),
    .X(_0880_));
 sg13g2_a21oi_1 _2414_ (.A1(_0879_),
    .A2(_0880_),
    .Y(_0881_),
    .B1(_0872_));
 sg13g2_xnor2_1 _2415_ (.Y(_0882_),
    .A(_0862_),
    .B(_0863_));
 sg13g2_o21ai_1 _2416_ (.B1(_0864_),
    .Y(_0883_),
    .A1(_0881_),
    .A2(_0882_));
 sg13g2_xor2_1 _2417_ (.B(_0848_),
    .A(_0847_),
    .X(_0884_));
 sg13g2_a21o_1 _2418_ (.A2(_0884_),
    .A1(_0883_),
    .B1(_0849_),
    .X(_0885_));
 sg13g2_xnor2_1 _2419_ (.Y(_0886_),
    .A(_0832_),
    .B(_0833_));
 sg13g2_a21o_1 _2420_ (.A2(_0886_),
    .A1(_0885_),
    .B1(_0835_),
    .X(_0887_));
 sg13g2_xor2_1 _2421_ (.B(_0820_),
    .A(_0819_),
    .X(_0888_));
 sg13g2_a21oi_1 _2422_ (.A1(_0887_),
    .A2(_0888_),
    .Y(_0890_),
    .B1(_0821_));
 sg13g2_xor2_1 _2423_ (.B(_0799_),
    .A(_0798_),
    .X(_0891_));
 sg13g2_nor2_1 _2424_ (.A(_0890_),
    .B(_0891_),
    .Y(_0892_));
 sg13g2_o21ai_1 _2425_ (.B1(_0800_),
    .Y(_0893_),
    .A1(_0890_),
    .A2(_0891_));
 sg13g2_xor2_1 _2426_ (.B(_0781_),
    .A(_0767_),
    .X(_0894_));
 sg13g2_a21o_1 _2427_ (.A2(_0894_),
    .A1(_0893_),
    .B1(_0782_),
    .X(_0895_));
 sg13g2_nand2_1 _2428_ (.Y(_0896_),
    .A(net354),
    .B(_0775_));
 sg13g2_a21oi_1 _2429_ (.A1(_0773_),
    .A2(_0776_),
    .Y(_0897_),
    .B1(_0772_));
 sg13g2_xor2_1 _2430_ (.B(_0729_),
    .A(_0610_),
    .X(_0898_));
 sg13g2_nand2b_1 _2431_ (.Y(_0899_),
    .B(_0898_),
    .A_N(_0897_));
 sg13g2_xnor2_1 _2432_ (.Y(_0901_),
    .A(_0897_),
    .B(_0898_));
 sg13g2_nand2b_1 _2433_ (.Y(_0902_),
    .B(_0901_),
    .A_N(_0896_));
 sg13g2_xnor2_1 _2434_ (.Y(_0903_),
    .A(_0896_),
    .B(_0901_));
 sg13g2_a21oi_1 _2435_ (.A1(_0769_),
    .A2(_0780_),
    .Y(_0904_),
    .B1(_0778_));
 sg13g2_nand2b_1 _2436_ (.Y(_0905_),
    .B(_0903_),
    .A_N(_0904_));
 sg13g2_inv_1 _2437_ (.Y(_0906_),
    .A(_0905_));
 sg13g2_xnor2_1 _2438_ (.Y(_0907_),
    .A(_0903_),
    .B(_0904_));
 sg13g2_xor2_1 _2439_ (.B(_0733_),
    .A(_0732_),
    .X(_0908_));
 sg13g2_a21o_1 _2440_ (.A2(_0902_),
    .A1(_0899_),
    .B1(_0908_),
    .X(_0909_));
 sg13g2_nand3_1 _2441_ (.B(_0902_),
    .C(_0908_),
    .A(_0899_),
    .Y(_0910_));
 sg13g2_and2_1 _2442_ (.A(_0909_),
    .B(_0910_),
    .X(_0912_));
 sg13g2_nand3_1 _2443_ (.B(_0907_),
    .C(_0912_),
    .A(_0895_),
    .Y(_0913_));
 sg13g2_nand2_1 _2444_ (.Y(_0914_),
    .A(_0905_),
    .B(_0909_));
 sg13g2_nand2_1 _2445_ (.Y(_0915_),
    .A(_0910_),
    .B(_0914_));
 sg13g2_a21oi_2 _2446_ (.B1(_0738_),
    .Y(_0916_),
    .A2(_0915_),
    .A1(_0913_));
 sg13g2_or2_1 _2447_ (.X(_0917_),
    .B(_0916_),
    .A(_0737_));
 sg13g2_or2_1 _2448_ (.X(_0918_),
    .B(_0602_),
    .A(_0596_));
 sg13g2_and2_1 _2449_ (.A(_0603_),
    .B(_0918_),
    .X(_0919_));
 sg13g2_o21ai_1 _2450_ (.B1(_0919_),
    .Y(_0920_),
    .A1(_0737_),
    .A2(_0916_));
 sg13g2_or3_1 _2451_ (.A(_0581_),
    .B(_0597_),
    .C(_0600_),
    .X(_0921_));
 sg13g2_nand3_1 _2452_ (.B(_0918_),
    .C(_0921_),
    .A(_0598_),
    .Y(_0923_));
 sg13g2_nor2b_1 _2453_ (.A(_0923_),
    .B_N(_0920_),
    .Y(_0924_));
 sg13g2_nand2b_1 _2454_ (.Y(_0925_),
    .B(_0920_),
    .A_N(_0923_));
 sg13g2_or3_1 _2455_ (.A(_0737_),
    .B(_0916_),
    .C(_0919_),
    .X(_0926_));
 sg13g2_and3_1 _2456_ (.X(_0927_),
    .A(_0738_),
    .B(_0913_),
    .C(_0915_));
 sg13g2_nor2_1 _2457_ (.A(_0916_),
    .B(_0927_),
    .Y(_0928_));
 sg13g2_a21oi_1 _2458_ (.A1(_0895_),
    .A2(_0907_),
    .Y(_0929_),
    .B1(_0906_));
 sg13g2_xor2_1 _2459_ (.B(_0929_),
    .A(_0912_),
    .X(_0930_));
 sg13g2_xor2_1 _2460_ (.B(_0907_),
    .A(_0895_),
    .X(_0931_));
 sg13g2_xor2_1 _2461_ (.B(_0894_),
    .A(_0893_),
    .X(_0932_));
 sg13g2_nor2_1 _2462_ (.A(_0931_),
    .B(_0932_),
    .Y(_0934_));
 sg13g2_nand2_1 _2463_ (.Y(_0935_),
    .A(_0930_),
    .B(_0934_));
 sg13g2_a21o_1 _2464_ (.A2(_0926_),
    .A1(_0920_),
    .B1(_0935_),
    .X(_0936_));
 sg13g2_o21ai_1 _2465_ (.B1(_0925_),
    .Y(_0937_),
    .A1(_0928_),
    .A2(_0936_));
 sg13g2_nand2_1 _2466_ (.Y(_0938_),
    .A(_0931_),
    .B(_0932_));
 sg13g2_nor4_1 _2467_ (.A(_0916_),
    .B(_0927_),
    .C(_0930_),
    .D(_0938_),
    .Y(_0939_));
 sg13g2_a221oi_1 _2468_ (.B2(_0939_),
    .C1(_0923_),
    .B1(_0926_),
    .A1(_0603_),
    .Y(_0940_),
    .A2(_0917_));
 sg13g2_xnor2_1 _2469_ (.Y(_0941_),
    .A(_0873_),
    .B(_0876_));
 sg13g2_or2_1 _2470_ (.X(_0942_),
    .B(_0941_),
    .A(_0940_));
 sg13g2_a21oi_1 _2471_ (.A1(net324),
    .A2(_0942_),
    .Y(_0943_),
    .B1(net344));
 sg13g2_xnor2_1 _2472_ (.Y(_0945_),
    .A(net394),
    .B(_0943_));
 sg13g2_nor3_1 _2473_ (.A(net417),
    .B(_1684_),
    .C(_0945_),
    .Y(_0072_));
 sg13g2_nand2_1 _2474_ (.Y(_0946_),
    .A(net388),
    .B(net344));
 sg13g2_a21oi_1 _2475_ (.A1(net324),
    .A2(_0942_),
    .Y(_0947_),
    .B1(net136));
 sg13g2_a21oi_1 _2476_ (.A1(_0873_),
    .A2(_0876_),
    .Y(_0948_),
    .B1(_0869_));
 sg13g2_xnor2_1 _2477_ (.Y(_0949_),
    .A(_0870_),
    .B(_0948_));
 sg13g2_or2_1 _2478_ (.X(_0950_),
    .B(_0949_),
    .A(_0940_));
 sg13g2_nand3_1 _2479_ (.B(net324),
    .C(_0950_),
    .A(_0027_),
    .Y(_0951_));
 sg13g2_a21o_1 _2480_ (.A2(_0950_),
    .A1(net324),
    .B1(_0027_),
    .X(_0952_));
 sg13g2_nand3_1 _2481_ (.B(_0951_),
    .C(_0952_),
    .A(_0947_),
    .Y(_0953_));
 sg13g2_a21oi_1 _2482_ (.A1(_0951_),
    .A2(_0952_),
    .Y(_0955_),
    .B1(_0947_));
 sg13g2_nand3b_1 _2483_ (.B(_1682_),
    .C(_0953_),
    .Y(_0956_),
    .A_N(_0955_));
 sg13g2_a21oi_1 _2484_ (.A1(_0946_),
    .A2(_0956_),
    .Y(_0073_),
    .B1(net417));
 sg13g2_a21o_1 _2485_ (.A2(_0950_),
    .A1(net324),
    .B1(_0779_),
    .X(_0957_));
 sg13g2_xnor2_1 _2486_ (.Y(_0958_),
    .A(_0879_),
    .B(_0880_));
 sg13g2_o21ai_1 _2487_ (.B1(net324),
    .Y(_0959_),
    .A1(_0940_),
    .A2(_0958_));
 sg13g2_xnor2_1 _2488_ (.Y(_0960_),
    .A(net383),
    .B(_0959_));
 sg13g2_nand3_1 _2489_ (.B(_0957_),
    .C(_0960_),
    .A(_0953_),
    .Y(_0961_));
 sg13g2_a21oi_1 _2490_ (.A1(_0953_),
    .A2(_0957_),
    .Y(_0962_),
    .B1(_0960_));
 sg13g2_nand3b_1 _2491_ (.B(_1682_),
    .C(_0961_),
    .Y(_0963_),
    .A_N(_0962_));
 sg13g2_a22oi_1 _2492_ (.Y(_0965_),
    .B1(_1684_),
    .B2(net96),
    .A2(net345),
    .A1(net382));
 sg13g2_a21oi_1 _2493_ (.A1(_0963_),
    .A2(_0965_),
    .Y(_0074_),
    .B1(net417));
 sg13g2_nor2b_1 _2494_ (.A(_0026_),
    .B_N(_0959_),
    .Y(_0966_));
 sg13g2_xnor2_1 _2495_ (.Y(_0967_),
    .A(_0881_),
    .B(_0882_));
 sg13g2_o21ai_1 _2496_ (.B1(net324),
    .Y(_0968_),
    .A1(_0940_),
    .A2(_0967_));
 sg13g2_xnor2_1 _2497_ (.Y(_0969_),
    .A(_0757_),
    .B(_0968_));
 sg13g2_nor3_1 _2498_ (.A(_0962_),
    .B(_0966_),
    .C(_0969_),
    .Y(_0970_));
 sg13g2_o21ai_1 _2499_ (.B1(_0969_),
    .Y(_0971_),
    .A1(_0962_),
    .A2(_0966_));
 sg13g2_nand3b_1 _2500_ (.B(_0971_),
    .C(_1682_),
    .Y(_0972_),
    .A_N(_0970_));
 sg13g2_a22oi_1 _2501_ (.Y(_0973_),
    .B1(_1684_),
    .B2(net98),
    .A2(net344),
    .A1(net378));
 sg13g2_a21oi_1 _2502_ (.A1(_0972_),
    .A2(net99),
    .Y(_0075_),
    .B1(net417));
 sg13g2_nand2b_1 _2503_ (.Y(_0975_),
    .B(_0968_),
    .A_N(_0025_));
 sg13g2_nand2_1 _2504_ (.Y(_0976_),
    .A(_0971_),
    .B(_0975_));
 sg13g2_xnor2_1 _2505_ (.Y(_0977_),
    .A(_0883_),
    .B(_0884_));
 sg13g2_o21ai_1 _2506_ (.B1(net324),
    .Y(_0978_),
    .A1(_0940_),
    .A2(_0977_));
 sg13g2_xor2_1 _2507_ (.B(_0978_),
    .A(net374),
    .X(_0979_));
 sg13g2_xnor2_1 _2508_ (.Y(_0980_),
    .A(_0976_),
    .B(_0979_));
 sg13g2_a22oi_1 _2509_ (.Y(_0981_),
    .B1(_1684_),
    .B2(net113),
    .A2(net345),
    .A1(net374));
 sg13g2_o21ai_1 _2510_ (.B1(_0981_),
    .Y(_0982_),
    .A1(_1683_),
    .A2(_0980_));
 sg13g2_and2_1 _2511_ (.A(net426),
    .B(_0982_),
    .X(_0076_));
 sg13g2_nor2b_1 _2512_ (.A(_0023_),
    .B_N(_0978_),
    .Y(_0984_));
 sg13g2_a21oi_1 _2513_ (.A1(_0976_),
    .A2(_0979_),
    .Y(_0985_),
    .B1(_0984_));
 sg13g2_xnor2_1 _2514_ (.Y(_0986_),
    .A(_0885_),
    .B(_0886_));
 sg13g2_o21ai_1 _2515_ (.B1(net325),
    .Y(_0987_),
    .A1(_0940_),
    .A2(_0986_));
 sg13g2_xor2_1 _2516_ (.B(_0987_),
    .A(\system_inst.neuron.v[5] ),
    .X(_0988_));
 sg13g2_xor2_1 _2517_ (.B(_0988_),
    .A(_0985_),
    .X(_0989_));
 sg13g2_nand2b_1 _2518_ (.Y(_0990_),
    .B(_1682_),
    .A_N(_0989_));
 sg13g2_a22oi_1 _2519_ (.Y(_0991_),
    .B1(_1684_),
    .B2(net89),
    .A2(net344),
    .A1(net95));
 sg13g2_a21oi_1 _2520_ (.A1(_0990_),
    .A2(_0991_),
    .Y(_0077_),
    .B1(net417));
 sg13g2_nand2_1 _2521_ (.Y(_0992_),
    .A(_0979_),
    .B(_0988_));
 sg13g2_a21oi_1 _2522_ (.A1(_0971_),
    .A2(_0975_),
    .Y(_0994_),
    .B1(_0992_));
 sg13g2_a22oi_1 _2523_ (.Y(_0995_),
    .B1(_0988_),
    .B2(_0984_),
    .A2(_0987_),
    .A1(_0993_));
 sg13g2_inv_1 _2524_ (.Y(_0996_),
    .A(_0995_));
 sg13g2_xnor2_1 _2525_ (.Y(_0997_),
    .A(_0887_),
    .B(_0888_));
 sg13g2_o21ai_1 _2526_ (.B1(net325),
    .Y(_0998_),
    .A1(_0940_),
    .A2(_0997_));
 sg13g2_xnor2_1 _2527_ (.Y(_0999_),
    .A(_0746_),
    .B(_0998_));
 sg13g2_nor3_1 _2528_ (.A(_0994_),
    .B(_0996_),
    .C(_0999_),
    .Y(_1000_));
 sg13g2_o21ai_1 _2529_ (.B1(_0999_),
    .Y(_1001_),
    .A1(_0994_),
    .A2(_0996_));
 sg13g2_nor2b_1 _2530_ (.A(_1000_),
    .B_N(_1001_),
    .Y(_1002_));
 sg13g2_a21oi_1 _2531_ (.A1(net364),
    .A2(net346),
    .Y(_1003_),
    .B1(net418));
 sg13g2_a22oi_1 _2532_ (.Y(_1005_),
    .B1(_1002_),
    .B2(_1682_),
    .A2(_1684_),
    .A1(net88));
 sg13g2_nand2_1 _2533_ (.Y(_0078_),
    .A(_1003_),
    .B(_1005_));
 sg13g2_a21oi_1 _2534_ (.A1(\system_inst.internal_param_c[5] ),
    .A2(\system_inst.internal_param_c[4] ),
    .Y(_1006_),
    .B1(_1063_));
 sg13g2_nand2b_1 _2535_ (.Y(_1007_),
    .B(net348),
    .A_N(_1006_));
 sg13g2_or2_1 _2536_ (.X(_1008_),
    .B(\system_inst.internal_param_c[4] ),
    .A(\system_inst.internal_param_c[5] ));
 sg13g2_a21oi_1 _2537_ (.A1(_1006_),
    .A2(_1008_),
    .Y(_1009_),
    .B1(net346));
 sg13g2_and2_1 _2538_ (.A(_0890_),
    .B(_0891_),
    .X(_1010_));
 sg13g2_or3_1 _2539_ (.A(_0892_),
    .B(_0940_),
    .C(_1010_),
    .X(_1011_));
 sg13g2_nand2_1 _2540_ (.Y(_1012_),
    .A(net325),
    .B(_1011_));
 sg13g2_a21oi_1 _2541_ (.A1(net325),
    .A2(_1011_),
    .Y(_1013_),
    .B1(_0735_));
 sg13g2_xnor2_1 _2542_ (.Y(_1015_),
    .A(net362),
    .B(_1012_));
 sg13g2_nand2b_1 _2543_ (.Y(_1016_),
    .B(_0998_),
    .A_N(_0021_));
 sg13g2_a21oi_1 _2544_ (.A1(_1001_),
    .A2(_1016_),
    .Y(_1017_),
    .B1(_1015_));
 sg13g2_nand3_1 _2545_ (.B(_1015_),
    .C(_1016_),
    .A(_1001_),
    .Y(_1018_));
 sg13g2_nand2_1 _2546_ (.Y(_1019_),
    .A(net336),
    .B(_1018_));
 sg13g2_o21ai_1 _2547_ (.B1(_1009_),
    .Y(_1020_),
    .A1(_1017_),
    .A2(_1019_));
 sg13g2_o21ai_1 _2548_ (.B1(_1020_),
    .Y(_1021_),
    .A1(net362),
    .A2(net348));
 sg13g2_nor2_1 _2549_ (.A(net418),
    .B(_1021_),
    .Y(_0079_));
 sg13g2_nor2_1 _2550_ (.A(net358),
    .B(net348),
    .Y(_1022_));
 sg13g2_xnor2_1 _2551_ (.Y(_1023_),
    .A(_0009_),
    .B(_0924_));
 sg13g2_o21ai_1 _2552_ (.B1(_1023_),
    .Y(_1025_),
    .A1(_1013_),
    .A2(_1017_));
 sg13g2_nor3_1 _2553_ (.A(_1013_),
    .B(_1017_),
    .C(_1023_),
    .Y(_1026_));
 sg13g2_nor2_1 _2554_ (.A(_1062_),
    .B(_1026_),
    .Y(_1027_));
 sg13g2_a21oi_1 _2555_ (.A1(_1025_),
    .A2(_1027_),
    .Y(_1028_),
    .B1(_1007_));
 sg13g2_o21ai_1 _2556_ (.B1(net426),
    .Y(_0080_),
    .A1(_1022_),
    .A2(_1028_));
 sg13g2_o21ai_1 _2557_ (.B1(_1025_),
    .Y(_1029_),
    .A1(_0724_),
    .A2(_0925_));
 sg13g2_xnor2_1 _2558_ (.Y(_1030_),
    .A(_0024_),
    .B(_0924_));
 sg13g2_xnor2_1 _2559_ (.Y(_1031_),
    .A(_1029_),
    .B(_1030_));
 sg13g2_nand2_1 _2560_ (.Y(_1032_),
    .A(net349),
    .B(net346));
 sg13g2_a21oi_1 _2561_ (.A1(_1007_),
    .A2(_1032_),
    .Y(_1033_),
    .B1(net418));
 sg13g2_o21ai_1 _2562_ (.B1(_1033_),
    .Y(_0081_),
    .A1(_1683_),
    .A2(_1031_));
 sg13g2_inv_2 _2563_ (.Y(_0713_),
    .A(net350));
 sg13g2_inv_1 _2564_ (.Y(_0724_),
    .A(net358));
 sg13g2_inv_2 _2565_ (.Y(_0735_),
    .A(net362));
 sg13g2_inv_2 _2566_ (.Y(_0746_),
    .A(net364));
 sg13g2_inv_2 _2567_ (.Y(_0757_),
    .A(net378));
 sg13g2_inv_2 _2568_ (.Y(_0768_),
    .A(net383));
 sg13g2_inv_2 _2569_ (.Y(_0779_),
    .A(net387));
 sg13g2_inv_1 _2570_ (.Y(_0790_),
    .A(net106));
 sg13g2_inv_1 _2571_ (.Y(_0801_),
    .A(net138));
 sg13g2_inv_2 _2572_ (.Y(_0812_),
    .A(net109));
 sg13g2_inv_2 _2573_ (.Y(_0823_),
    .A(net120));
 sg13g2_inv_1 _2574_ (.Y(_0834_),
    .A(\system_inst.loader.shift_reg[1] ));
 sg13g2_inv_2 _2575_ (.Y(_0845_),
    .A(net104));
 sg13g2_inv_1 _2576_ (.Y(_0856_),
    .A(net100));
 sg13g2_inv_1 _2577_ (.Y(_0867_),
    .A(net12));
 sg13g2_inv_1 _2578_ (.Y(_0878_),
    .A(net89));
 sg13g2_inv_1 _2579_ (.Y(_0889_),
    .A(net400));
 sg13g2_inv_1 _2580_ (.Y(_0900_),
    .A(net408));
 sg13g2_inv_2 _2581_ (.Y(_0911_),
    .A(net146));
 sg13g2_inv_1 _2582_ (.Y(_0922_),
    .A(net410));
 sg13g2_inv_1 _2583_ (.Y(_0933_),
    .A(net412));
 sg13g2_inv_1 _2584_ (.Y(_0944_),
    .A(net415));
 sg13g2_inv_2 _2585_ (.Y(_0954_),
    .A(\system_inst.neuron.u[7] ));
 sg13g2_inv_1 _2586_ (.Y(_0964_),
    .A(\system_inst.neuron.u[4] ));
 sg13g2_inv_1 _2587_ (.Y(_0974_),
    .A(net425));
 sg13g2_inv_1 _2588_ (.Y(_0983_),
    .A(net102));
 sg13g2_inv_2 _2589_ (.Y(_0993_),
    .A(_0022_));
 sg13g2_inv_1 _2590_ (.Y(_1004_),
    .A(_0024_));
 sg13g2_inv_1 _2591_ (.Y(_1014_),
    .A(_0011_));
 sg13g2_inv_2 _2592_ (.Y(_1024_),
    .A(_0016_));
 sg13g2_inv_2 _2593_ (.Y(_1034_),
    .A(_0017_));
 sg13g2_inv_1 _2594_ (.Y(_1035_),
    .A(_0018_));
 sg13g2_nand3b_1 _2595_ (.B(\system_inst.loader.bit_count[0] ),
    .C(\system_inst.loader.bit_count[2] ),
    .Y(_1036_),
    .A_N(\system_inst.loader.bit_count[1] ));
 sg13g2_nand2_1 _2596_ (.Y(_1037_),
    .A(net1),
    .B(net11));
 sg13g2_nor2_2 _2597_ (.A(_1036_),
    .B(_1037_),
    .Y(_1038_));
 sg13g2_or2_2 _2598_ (.X(_1039_),
    .B(_1037_),
    .A(_1036_));
 sg13g2_and2_1 _2599_ (.A(net111),
    .B(_1038_),
    .X(_1040_));
 sg13g2_nand2_2 _2600_ (.Y(_1041_),
    .A(net111),
    .B(_1038_));
 sg13g2_a21oi_1 _2601_ (.A1(net108),
    .A2(_1039_),
    .Y(_1042_),
    .B1(_1040_));
 sg13g2_nor2_1 _2602_ (.A(net420),
    .B(_1042_),
    .Y(_0005_));
 sg13g2_and2_2 _2603_ (.A(net108),
    .B(_1038_),
    .X(_1043_));
 sg13g2_nand2_2 _2604_ (.Y(_1044_),
    .A(net108),
    .B(_1038_));
 sg13g2_a21oi_1 _2605_ (.A1(net102),
    .A2(_1039_),
    .Y(_1045_),
    .B1(_1043_));
 sg13g2_nor2_1 _2606_ (.A(net419),
    .B(net103),
    .Y(_0001_));
 sg13g2_nor2_2 _2607_ (.A(\system_inst.loader.state[4] ),
    .B(\system_inst.loader.state[0] ),
    .Y(_1046_));
 sg13g2_or2_1 _2608_ (.X(_1047_),
    .B(net129),
    .A(net116));
 sg13g2_nand2b_1 _2609_ (.Y(_1048_),
    .B(net11),
    .A_N(\system_inst.loader.load_enable_prev ));
 sg13g2_nor2_1 _2610_ (.A(\system_inst.loader.load_enable_prev ),
    .B(_1037_),
    .Y(_1049_));
 sg13g2_a22oi_1 _2611_ (.Y(_1050_),
    .B1(_1047_),
    .B2(_1049_),
    .A2(_1039_),
    .A1(net93));
 sg13g2_nor2_1 _2612_ (.A(net419),
    .B(net94),
    .Y(_0003_));
 sg13g2_and2_1 _2613_ (.A(net426),
    .B(net11),
    .X(_0082_));
 sg13g2_nor2_1 _2614_ (.A(net1),
    .B(net419),
    .Y(_1051_));
 sg13g2_a21o_1 _2615_ (.A2(_0082_),
    .A1(\system_inst.loader.load_enable_prev ),
    .B1(_1051_),
    .X(_1052_));
 sg13g2_and2_1 _2616_ (.A(net11),
    .B(\system_inst.loader.state[1] ),
    .X(_1053_));
 sg13g2_nor2_2 _2617_ (.A(_0983_),
    .B(_1039_),
    .Y(_1054_));
 sg13g2_a22oi_1 _2618_ (.Y(_1055_),
    .B1(_1054_),
    .B2(net426),
    .A2(_1052_),
    .A1(net116));
 sg13g2_inv_1 _2619_ (.Y(_0004_),
    .A(net117));
 sg13g2_o21ai_1 _2620_ (.B1(net129),
    .Y(_1056_),
    .A1(_1048_),
    .A2(_1051_));
 sg13g2_nand3b_1 _2621_ (.B(net1),
    .C(net116),
    .Y(_1057_),
    .A_N(net11));
 sg13g2_nand3_1 _2622_ (.B(net130),
    .C(_1057_),
    .A(net426),
    .Y(_0000_));
 sg13g2_and2_1 _2623_ (.A(net93),
    .B(_1038_),
    .X(_1058_));
 sg13g2_a21oi_1 _2624_ (.A1(net111),
    .A2(_1039_),
    .Y(_1059_),
    .B1(net338));
 sg13g2_nor2_1 _2625_ (.A(net419),
    .B(_1059_),
    .Y(_0002_));
 sg13g2_nor2_1 _2626_ (.A(_0713_),
    .B(net361),
    .Y(_1060_));
 sg13g2_nand2_2 _2627_ (.Y(_1061_),
    .A(net358),
    .B(net366));
 sg13g2_o21ai_1 _2628_ (.B1(net354),
    .Y(_1062_),
    .A1(_0735_),
    .A2(_1061_));
 sg13g2_a21o_1 _2629_ (.A2(_1061_),
    .A1(net354),
    .B1(_1060_),
    .X(_1063_));
 sg13g2_nand2_2 _2630_ (.Y(uo_out[0]),
    .A(_0026_),
    .B(net334));
 sg13g2_nand2_2 _2631_ (.Y(uo_out[1]),
    .A(_0025_),
    .B(net334));
 sg13g2_nand2_2 _2632_ (.Y(uo_out[2]),
    .A(_0023_),
    .B(net336));
 sg13g2_nand2_2 _2633_ (.Y(uo_out[3]),
    .A(_0022_),
    .B(net336));
 sg13g2_nand2_2 _2634_ (.Y(_1064_),
    .A(\system_inst.neuron.v[8] ),
    .B(net361));
 sg13g2_nand3_1 _2635_ (.B(net364),
    .C(_1064_),
    .A(net354),
    .Y(uo_out[4]));
 sg13g2_nand2_2 _2636_ (.Y(_1065_),
    .A(net361),
    .B(net364));
 sg13g2_o21ai_1 _2637_ (.B1(net354),
    .Y(_1066_),
    .A1(net361),
    .A2(net364));
 sg13g2_nand2b_1 _2638_ (.Y(uo_out[5]),
    .B(_1065_),
    .A_N(_1066_));
 sg13g2_xor2_1 _2639_ (.B(net364),
    .A(net358),
    .X(_1067_));
 sg13g2_o21ai_1 _2640_ (.B1(_1064_),
    .Y(_1068_),
    .A1(net361),
    .A2(_1067_));
 sg13g2_nand2_2 _2641_ (.Y(uo_out[6]),
    .A(net336),
    .B(_1068_));
 sg13g2_nand3_1 _2642_ (.B(_1061_),
    .C(_1064_),
    .A(net354),
    .Y(uo_out[7]));
 sg13g2_nand2_1 _2643_ (.Y(_1069_),
    .A(net392),
    .B(net400));
 sg13g2_and4_1 _2644_ (.A(net387),
    .B(net392),
    .C(net398),
    .D(net400),
    .X(_1070_));
 sg13g2_nand2_1 _2645_ (.Y(_1071_),
    .A(net380),
    .B(net400));
 sg13g2_and4_1 _2646_ (.A(net389),
    .B(net391),
    .C(net396),
    .D(net398),
    .X(_1072_));
 sg13g2_a22oi_1 _2647_ (.Y(_1073_),
    .B1(net398),
    .B2(net387),
    .A2(net396),
    .A1(net391));
 sg13g2_or3_1 _2648_ (.A(_1071_),
    .B(_1072_),
    .C(_1073_),
    .X(_1074_));
 sg13g2_o21ai_1 _2649_ (.B1(_1071_),
    .Y(_1075_),
    .A1(_1072_),
    .A2(_1073_));
 sg13g2_nand3_1 _2650_ (.B(_1074_),
    .C(_1075_),
    .A(_1070_),
    .Y(_1076_));
 sg13g2_a21o_1 _2651_ (.A2(_1075_),
    .A1(_1074_),
    .B1(_1070_),
    .X(_1077_));
 sg13g2_nand2_1 _2652_ (.Y(_1078_),
    .A(net368),
    .B(\system_inst.internal_param_b[0] ));
 sg13g2_nand2_1 _2653_ (.Y(_1079_),
    .A(net371),
    .B(net401));
 sg13g2_nand2_1 _2654_ (.Y(_1080_),
    .A(net372),
    .B(net404));
 sg13g2_nand2_1 _2655_ (.Y(_1081_),
    .A(net376),
    .B(net402));
 sg13g2_xor2_1 _2656_ (.B(_1081_),
    .A(_1080_),
    .X(_1082_));
 sg13g2_nand2b_1 _2657_ (.Y(_1083_),
    .B(_1082_),
    .A_N(_1078_));
 sg13g2_xnor2_1 _2658_ (.Y(_1084_),
    .A(_1078_),
    .B(_1082_));
 sg13g2_nand3_1 _2659_ (.B(_1077_),
    .C(_1084_),
    .A(_1076_),
    .Y(_1085_));
 sg13g2_nand2_1 _2660_ (.Y(_1086_),
    .A(_1076_),
    .B(_1085_));
 sg13g2_nand2b_1 _2661_ (.Y(_1087_),
    .B(_1074_),
    .A_N(_1072_));
 sg13g2_nand2_1 _2662_ (.Y(_1088_),
    .A(net375),
    .B(net399));
 sg13g2_nand2_1 _2663_ (.Y(_1089_),
    .A(net379),
    .B(net395));
 sg13g2_and4_1 _2664_ (.A(net379),
    .B(net384),
    .C(net395),
    .D(net397),
    .X(_1090_));
 sg13g2_a22oi_1 _2665_ (.Y(_1091_),
    .B1(net397),
    .B2(net379),
    .A2(net395),
    .A1(net384));
 sg13g2_nor3_1 _2666_ (.A(_1088_),
    .B(_1090_),
    .C(_1091_),
    .Y(_1092_));
 sg13g2_o21ai_1 _2667_ (.B1(_1088_),
    .Y(_1093_),
    .A1(_1090_),
    .A2(_1091_));
 sg13g2_nor2b_1 _2668_ (.A(_1092_),
    .B_N(_1093_),
    .Y(_1094_));
 sg13g2_xnor2_1 _2669_ (.Y(_1095_),
    .A(_1087_),
    .B(_1094_));
 sg13g2_nand2_1 _2670_ (.Y(_1096_),
    .A(net363),
    .B(net405));
 sg13g2_nand2_1 _2671_ (.Y(_1097_),
    .A(net367),
    .B(net401));
 sg13g2_nand2_1 _2672_ (.Y(_1098_),
    .A(net367),
    .B(net403));
 sg13g2_xor2_1 _2673_ (.B(_1098_),
    .A(_1079_),
    .X(_1099_));
 sg13g2_nand2b_1 _2674_ (.Y(_1100_),
    .B(_1099_),
    .A_N(_1096_));
 sg13g2_xnor2_1 _2675_ (.Y(_1101_),
    .A(_1096_),
    .B(_1099_));
 sg13g2_nor2b_1 _2676_ (.A(_1095_),
    .B_N(_1101_),
    .Y(_1102_));
 sg13g2_xnor2_1 _2677_ (.Y(_1103_),
    .A(_1095_),
    .B(_1101_));
 sg13g2_o21ai_1 _2678_ (.B1(_1083_),
    .Y(_1104_),
    .A1(_1080_),
    .A2(_1081_));
 sg13g2_xnor2_1 _2679_ (.Y(_1105_),
    .A(_1086_),
    .B(_1103_));
 sg13g2_nor2b_1 _2680_ (.A(_1105_),
    .B_N(_1104_),
    .Y(_1106_));
 sg13g2_a21o_1 _2681_ (.A2(_1103_),
    .A1(_1086_),
    .B1(_1106_),
    .X(_1107_));
 sg13g2_o21ai_1 _2682_ (.B1(_1100_),
    .Y(_1108_),
    .A1(_1079_),
    .A2(_1098_));
 sg13g2_a21o_1 _2683_ (.A2(_1094_),
    .A1(_1087_),
    .B1(_1102_),
    .X(_1109_));
 sg13g2_or2_1 _2684_ (.X(_1110_),
    .B(_1092_),
    .A(_1090_));
 sg13g2_nand2_1 _2685_ (.Y(_1111_),
    .A(net371),
    .B(net399));
 sg13g2_nand2_1 _2686_ (.Y(_1112_),
    .A(net375),
    .B(net395));
 sg13g2_nand2_1 _2687_ (.Y(_1113_),
    .A(net375),
    .B(net397));
 sg13g2_xor2_1 _2688_ (.B(_1113_),
    .A(_1089_),
    .X(_1114_));
 sg13g2_nand2b_1 _2689_ (.Y(_1115_),
    .B(_1114_),
    .A_N(_1111_));
 sg13g2_xnor2_1 _2690_ (.Y(_1116_),
    .A(_1111_),
    .B(_1114_));
 sg13g2_xnor2_1 _2691_ (.Y(_1117_),
    .A(_1110_),
    .B(_1116_));
 sg13g2_nand2_1 _2692_ (.Y(_1118_),
    .A(net359),
    .B(net405));
 sg13g2_nand2_1 _2693_ (.Y(_1119_),
    .A(net363),
    .B(net401));
 sg13g2_nand2_1 _2694_ (.Y(_1120_),
    .A(net363),
    .B(net403));
 sg13g2_xor2_1 _2695_ (.B(_1120_),
    .A(_1097_),
    .X(_1121_));
 sg13g2_nand2b_1 _2696_ (.Y(_1122_),
    .B(_1121_),
    .A_N(_1118_));
 sg13g2_xnor2_1 _2697_ (.Y(_1123_),
    .A(_1118_),
    .B(_1121_));
 sg13g2_nor2b_1 _2698_ (.A(_1117_),
    .B_N(_1123_),
    .Y(_1124_));
 sg13g2_xnor2_1 _2699_ (.Y(_1125_),
    .A(_1117_),
    .B(_1123_));
 sg13g2_xnor2_1 _2700_ (.Y(_1126_),
    .A(_1109_),
    .B(_1125_));
 sg13g2_nor2b_1 _2701_ (.A(_1126_),
    .B_N(_1108_),
    .Y(_1127_));
 sg13g2_xor2_1 _2702_ (.B(_1126_),
    .A(_1108_),
    .X(_1128_));
 sg13g2_nor2b_1 _2703_ (.A(_1128_),
    .B_N(_1107_),
    .Y(_1129_));
 sg13g2_a22oi_1 _2704_ (.Y(_1130_),
    .B1(net399),
    .B2(net387),
    .A2(net398),
    .A1(net392));
 sg13g2_nor2_1 _2705_ (.A(_1070_),
    .B(_1130_),
    .Y(_1131_));
 sg13g2_nand2_1 _2706_ (.Y(_1132_),
    .A(net372),
    .B(\system_inst.internal_param_b[0] ));
 sg13g2_nand2_1 _2707_ (.Y(_1133_),
    .A(net382),
    .B(net404));
 sg13g2_and4_1 _2708_ (.A(net376),
    .B(net380),
    .C(net402),
    .D(net403),
    .X(_1134_));
 sg13g2_a22oi_1 _2709_ (.Y(_1135_),
    .B1(net403),
    .B2(net378),
    .A2(net402),
    .A1(net382));
 sg13g2_o21ai_1 _2710_ (.B1(_1132_),
    .Y(_1136_),
    .A1(_1134_),
    .A2(_1135_));
 sg13g2_or3_1 _2711_ (.A(_1132_),
    .B(_1134_),
    .C(_1135_),
    .X(_1137_));
 sg13g2_nand3_1 _2712_ (.B(_1136_),
    .C(_1137_),
    .A(_1131_),
    .Y(_1138_));
 sg13g2_inv_1 _2713_ (.Y(_1139_),
    .A(_1138_));
 sg13g2_a21o_1 _2714_ (.A2(_1077_),
    .A1(_1076_),
    .B1(_1084_),
    .X(_1140_));
 sg13g2_and2_1 _2715_ (.A(_1085_),
    .B(_1140_),
    .X(_1141_));
 sg13g2_nand3_1 _2716_ (.B(_1139_),
    .C(_1140_),
    .A(_1085_),
    .Y(_1142_));
 sg13g2_nand2b_1 _2717_ (.Y(_1143_),
    .B(_1137_),
    .A_N(_1134_));
 sg13g2_a21o_1 _2718_ (.A2(_1140_),
    .A1(_1085_),
    .B1(_1139_),
    .X(_1144_));
 sg13g2_and3_1 _2719_ (.X(_1145_),
    .A(_1142_),
    .B(_1143_),
    .C(_1144_));
 sg13g2_a21oi_2 _2720_ (.B1(_1145_),
    .Y(_1146_),
    .A2(_1141_),
    .A1(_1139_));
 sg13g2_xor2_1 _2721_ (.B(_1105_),
    .A(_1104_),
    .X(_1147_));
 sg13g2_or2_1 _2722_ (.X(_1148_),
    .B(_1147_),
    .A(_1146_));
 sg13g2_nand2_1 _2723_ (.Y(_1149_),
    .A(net378),
    .B(net405));
 sg13g2_nand2_1 _2724_ (.Y(_1150_),
    .A(net387),
    .B(net402));
 sg13g2_xor2_1 _2725_ (.B(_1150_),
    .A(_1133_),
    .X(_1151_));
 sg13g2_nand2b_1 _2726_ (.Y(_1152_),
    .B(_1151_),
    .A_N(_1149_));
 sg13g2_xnor2_1 _2727_ (.Y(_1153_),
    .A(_1149_),
    .B(_1151_));
 sg13g2_nand2b_1 _2728_ (.Y(_1154_),
    .B(_1153_),
    .A_N(_1069_));
 sg13g2_a21o_1 _2729_ (.A2(_1137_),
    .A1(_1136_),
    .B1(_1131_),
    .X(_1155_));
 sg13g2_nand2_1 _2730_ (.Y(_1156_),
    .A(_1138_),
    .B(_1155_));
 sg13g2_nor2_1 _2731_ (.A(_1154_),
    .B(_1156_),
    .Y(_1157_));
 sg13g2_o21ai_1 _2732_ (.B1(_1152_),
    .Y(_1158_),
    .A1(_1133_),
    .A2(_1150_));
 sg13g2_xor2_1 _2733_ (.B(_1156_),
    .A(_1154_),
    .X(_1159_));
 sg13g2_a21oi_1 _2734_ (.A1(_1158_),
    .A2(_1159_),
    .Y(_1160_),
    .B1(_1157_));
 sg13g2_a21oi_1 _2735_ (.A1(_1142_),
    .A2(_1144_),
    .Y(_1161_),
    .B1(_1143_));
 sg13g2_nor3_1 _2736_ (.A(_1145_),
    .B(_1160_),
    .C(_1161_),
    .Y(_1162_));
 sg13g2_xnor2_1 _2737_ (.Y(_1163_),
    .A(_1069_),
    .B(_1153_));
 sg13g2_a22oi_1 _2738_ (.Y(_1164_),
    .B1(net404),
    .B2(net388),
    .A2(net401),
    .A1(net392));
 sg13g2_nand2_1 _2739_ (.Y(_1165_),
    .A(net382),
    .B(net405));
 sg13g2_nand4_1 _2740_ (.B(net392),
    .C(net402),
    .A(net388),
    .Y(_1166_),
    .D(net404));
 sg13g2_a21oi_1 _2741_ (.A1(_1165_),
    .A2(_1166_),
    .Y(_1167_),
    .B1(_1164_));
 sg13g2_nand2_1 _2742_ (.Y(_1168_),
    .A(_1163_),
    .B(_1167_));
 sg13g2_xnor2_1 _2743_ (.Y(_1169_),
    .A(_1158_),
    .B(_1159_));
 sg13g2_nor2_1 _2744_ (.A(_1168_),
    .B(_1169_),
    .Y(_1170_));
 sg13g2_xnor2_1 _2745_ (.Y(_1171_),
    .A(_1163_),
    .B(_1167_));
 sg13g2_and2_2 _2746_ (.A(net385),
    .B(net390),
    .X(_1172_));
 sg13g2_nand2_2 _2747_ (.Y(_1173_),
    .A(net384),
    .B(net391));
 sg13g2_nand2_1 _2748_ (.Y(_1174_),
    .A(net403),
    .B(net405));
 sg13g2_nor3_1 _2749_ (.A(_1151_),
    .B(_1173_),
    .C(_1174_),
    .Y(_1175_));
 sg13g2_nand2b_1 _2750_ (.Y(_1176_),
    .B(_1175_),
    .A_N(_1171_));
 sg13g2_a21oi_1 _2751_ (.A1(_1168_),
    .A2(_1176_),
    .Y(_1177_),
    .B1(_1169_));
 sg13g2_o21ai_1 _2752_ (.B1(_1160_),
    .Y(_1178_),
    .A1(_1145_),
    .A2(_1161_));
 sg13g2_nor2b_1 _2753_ (.A(_1162_),
    .B_N(_1178_),
    .Y(_1179_));
 sg13g2_a21oi_1 _2754_ (.A1(_1177_),
    .A2(_1178_),
    .Y(_1180_),
    .B1(_1162_));
 sg13g2_and2_1 _2755_ (.A(_1146_),
    .B(_1147_),
    .X(_1181_));
 sg13g2_xor2_1 _2756_ (.B(_1147_),
    .A(_1146_),
    .X(_1182_));
 sg13g2_o21ai_1 _2757_ (.B1(_1148_),
    .Y(_1183_),
    .A1(_1180_),
    .A2(_1181_));
 sg13g2_xnor2_1 _2758_ (.Y(_1184_),
    .A(_1107_),
    .B(_1128_));
 sg13g2_a21o_1 _2759_ (.A2(_1184_),
    .A1(_1183_),
    .B1(_1129_),
    .X(_1185_));
 sg13g2_a21o_1 _2760_ (.A2(_1125_),
    .A1(_1109_),
    .B1(_1127_),
    .X(_1186_));
 sg13g2_o21ai_1 _2761_ (.B1(_1122_),
    .Y(_1187_),
    .A1(_1097_),
    .A2(_1120_));
 sg13g2_inv_1 _2762_ (.Y(_1188_),
    .A(_1187_));
 sg13g2_a21o_1 _2763_ (.A2(_1116_),
    .A1(_1110_),
    .B1(_1124_),
    .X(_1189_));
 sg13g2_o21ai_1 _2764_ (.B1(_1115_),
    .Y(_1190_),
    .A1(_1089_),
    .A2(_1113_));
 sg13g2_nand2_1 _2765_ (.Y(_1191_),
    .A(net367),
    .B(net399));
 sg13g2_nand2_1 _2766_ (.Y(_1192_),
    .A(net371),
    .B(net395));
 sg13g2_nand2_1 _2767_ (.Y(_1193_),
    .A(net371),
    .B(net397));
 sg13g2_xor2_1 _2768_ (.B(_1193_),
    .A(_1112_),
    .X(_1194_));
 sg13g2_nand2b_1 _2769_ (.Y(_1195_),
    .B(_1194_),
    .A_N(_1191_));
 sg13g2_xnor2_1 _2770_ (.Y(_1196_),
    .A(_1191_),
    .B(_1194_));
 sg13g2_xnor2_1 _2771_ (.Y(_1197_),
    .A(_1190_),
    .B(_1196_));
 sg13g2_nand2_1 _2772_ (.Y(_1198_),
    .A(net356),
    .B(net405));
 sg13g2_nand2_1 _2773_ (.Y(_1199_),
    .A(net359),
    .B(net401));
 sg13g2_nand2_1 _2774_ (.Y(_1200_),
    .A(net359),
    .B(net403));
 sg13g2_xor2_1 _2775_ (.B(_1200_),
    .A(_1119_),
    .X(_1201_));
 sg13g2_nand2b_1 _2776_ (.Y(_1202_),
    .B(_1201_),
    .A_N(_1198_));
 sg13g2_xnor2_1 _2777_ (.Y(_1203_),
    .A(_1198_),
    .B(_1201_));
 sg13g2_nor2b_1 _2778_ (.A(_1197_),
    .B_N(_1203_),
    .Y(_1204_));
 sg13g2_xnor2_1 _2779_ (.Y(_1205_),
    .A(_1197_),
    .B(_1203_));
 sg13g2_nand2_1 _2780_ (.Y(_1206_),
    .A(_1189_),
    .B(_1205_));
 sg13g2_xnor2_1 _2781_ (.Y(_1207_),
    .A(_1189_),
    .B(_1205_));
 sg13g2_xnor2_1 _2782_ (.Y(_1208_),
    .A(_1188_),
    .B(_1207_));
 sg13g2_nor2b_1 _2783_ (.A(_1208_),
    .B_N(_1186_),
    .Y(_1209_));
 sg13g2_nand2b_1 _2784_ (.Y(_1210_),
    .B(_1208_),
    .A_N(_1186_));
 sg13g2_xor2_1 _2785_ (.B(_1208_),
    .A(_1186_),
    .X(_1211_));
 sg13g2_xnor2_1 _2786_ (.Y(_1212_),
    .A(_1185_),
    .B(_1211_));
 sg13g2_and2_1 _2787_ (.A(_0012_),
    .B(_1212_),
    .X(_1213_));
 sg13g2_xor2_1 _2788_ (.B(_1179_),
    .A(_1177_),
    .X(_1214_));
 sg13g2_nand2b_1 _2789_ (.Y(_1215_),
    .B(\system_inst.neuron.u[0] ),
    .A_N(_1214_));
 sg13g2_xnor2_1 _2790_ (.Y(_1216_),
    .A(_1180_),
    .B(_1182_));
 sg13g2_xnor2_1 _2791_ (.Y(_1217_),
    .A(\system_inst.neuron.u[1] ),
    .B(_1216_));
 sg13g2_a22oi_1 _2792_ (.Y(_1218_),
    .B1(_1217_),
    .B2(_1215_),
    .A2(_1216_),
    .A1(_0013_));
 sg13g2_xnor2_1 _2793_ (.Y(_1219_),
    .A(_1183_),
    .B(_1184_));
 sg13g2_xor2_1 _2794_ (.B(_1219_),
    .A(_0014_),
    .X(_1220_));
 sg13g2_or2_1 _2795_ (.X(_1221_),
    .B(_1219_),
    .A(\system_inst.neuron.u[2] ));
 sg13g2_o21ai_1 _2796_ (.B1(_1221_),
    .Y(_1222_),
    .A1(_1218_),
    .A2(_1220_));
 sg13g2_or2_1 _2797_ (.X(_1223_),
    .B(_1212_),
    .A(_0012_));
 sg13g2_xnor2_1 _2798_ (.Y(_1224_),
    .A(_0012_),
    .B(_1212_));
 sg13g2_a21o_1 _2799_ (.A2(_1223_),
    .A1(_1222_),
    .B1(_1213_),
    .X(_1225_));
 sg13g2_a21oi_1 _2800_ (.A1(_1185_),
    .A2(_1210_),
    .Y(_1226_),
    .B1(_1209_));
 sg13g2_o21ai_1 _2801_ (.B1(_1206_),
    .Y(_1227_),
    .A1(_1188_),
    .A2(_1207_));
 sg13g2_o21ai_1 _2802_ (.B1(_1202_),
    .Y(_1228_),
    .A1(_1119_),
    .A2(_1200_));
 sg13g2_inv_1 _2803_ (.Y(_1229_),
    .A(_1228_));
 sg13g2_a21o_1 _2804_ (.A2(_1196_),
    .A1(_1190_),
    .B1(_1204_),
    .X(_1230_));
 sg13g2_o21ai_1 _2805_ (.B1(_1195_),
    .Y(_1231_),
    .A1(_1112_),
    .A2(_1193_));
 sg13g2_nand2_1 _2806_ (.Y(_1232_),
    .A(net363),
    .B(net399));
 sg13g2_nand2_1 _2807_ (.Y(_1233_),
    .A(net367),
    .B(net395));
 sg13g2_nand2_1 _2808_ (.Y(_1234_),
    .A(net367),
    .B(net397));
 sg13g2_xor2_1 _2809_ (.B(_1234_),
    .A(_1192_),
    .X(_1235_));
 sg13g2_nand2b_1 _2810_ (.Y(_1236_),
    .B(_1235_),
    .A_N(_1232_));
 sg13g2_xnor2_1 _2811_ (.Y(_1237_),
    .A(_1232_),
    .B(_1235_));
 sg13g2_xnor2_1 _2812_ (.Y(_1238_),
    .A(_1231_),
    .B(_1237_));
 sg13g2_nand2_1 _2813_ (.Y(_1239_),
    .A(net353),
    .B(net405));
 sg13g2_nand2_1 _2814_ (.Y(_1240_),
    .A(net356),
    .B(net403));
 sg13g2_xor2_1 _2815_ (.B(_1240_),
    .A(_1199_),
    .X(_1241_));
 sg13g2_nand2b_1 _2816_ (.Y(_1242_),
    .B(_1241_),
    .A_N(_1239_));
 sg13g2_xnor2_1 _2817_ (.Y(_1243_),
    .A(_1239_),
    .B(_1241_));
 sg13g2_nor2b_1 _2818_ (.A(_1238_),
    .B_N(_1243_),
    .Y(_1244_));
 sg13g2_xnor2_1 _2819_ (.Y(_1245_),
    .A(_1238_),
    .B(_1243_));
 sg13g2_nand2_1 _2820_ (.Y(_1246_),
    .A(_1230_),
    .B(_1245_));
 sg13g2_xnor2_1 _2821_ (.Y(_1247_),
    .A(_1230_),
    .B(_1245_));
 sg13g2_xnor2_1 _2822_ (.Y(_1248_),
    .A(_1229_),
    .B(_1247_));
 sg13g2_nand2b_1 _2823_ (.Y(_1249_),
    .B(_1227_),
    .A_N(_1248_));
 sg13g2_xor2_1 _2824_ (.B(_1248_),
    .A(_1227_),
    .X(_1250_));
 sg13g2_xnor2_1 _2825_ (.Y(_1251_),
    .A(_1226_),
    .B(_1250_));
 sg13g2_xor2_1 _2826_ (.B(_1251_),
    .A(_0015_),
    .X(_1252_));
 sg13g2_xnor2_1 _2827_ (.Y(_1253_),
    .A(_0015_),
    .B(_1251_));
 sg13g2_nor2_1 _2828_ (.A(\system_inst.neuron.u[4] ),
    .B(_1251_),
    .Y(_1254_));
 sg13g2_a21o_2 _2829_ (.A2(_1253_),
    .A1(_1225_),
    .B1(_1254_),
    .X(_1255_));
 sg13g2_o21ai_1 _2830_ (.B1(_1249_),
    .Y(_1256_),
    .A1(_1226_),
    .A2(_1250_));
 sg13g2_o21ai_1 _2831_ (.B1(_1246_),
    .Y(_1257_),
    .A1(_1229_),
    .A2(_1247_));
 sg13g2_o21ai_1 _2832_ (.B1(_1242_),
    .Y(_1258_),
    .A1(_1199_),
    .A2(_1240_));
 sg13g2_a21o_1 _2833_ (.A2(_1237_),
    .A1(_1231_),
    .B1(_1244_),
    .X(_1259_));
 sg13g2_nand2_1 _2834_ (.Y(_1260_),
    .A(net353),
    .B(net401));
 sg13g2_or2_1 _2835_ (.X(_1261_),
    .B(_1260_),
    .A(_1240_));
 sg13g2_inv_1 _2836_ (.Y(_1262_),
    .A(_1261_));
 sg13g2_a22oi_1 _2837_ (.Y(_1263_),
    .B1(net403),
    .B2(net353),
    .A2(net401),
    .A1(net356));
 sg13g2_nor2_1 _2838_ (.A(_1262_),
    .B(_1263_),
    .Y(_1264_));
 sg13g2_inv_1 _2839_ (.Y(_1265_),
    .A(_1264_));
 sg13g2_o21ai_1 _2840_ (.B1(_1236_),
    .Y(_1266_),
    .A1(_1192_),
    .A2(_1234_));
 sg13g2_nand2_1 _2841_ (.Y(_1267_),
    .A(net359),
    .B(net399));
 sg13g2_nand2_1 _2842_ (.Y(_1268_),
    .A(net363),
    .B(net395));
 sg13g2_nand2_1 _2843_ (.Y(_1269_),
    .A(net363),
    .B(net397));
 sg13g2_xor2_1 _2844_ (.B(_1269_),
    .A(_1233_),
    .X(_1270_));
 sg13g2_nand2b_1 _2845_ (.Y(_1271_),
    .B(_1270_),
    .A_N(_1267_));
 sg13g2_xnor2_1 _2846_ (.Y(_1272_),
    .A(_1267_),
    .B(_1270_));
 sg13g2_nand2_1 _2847_ (.Y(_1273_),
    .A(_1266_),
    .B(_1272_));
 sg13g2_xnor2_1 _2848_ (.Y(_1274_),
    .A(_1266_),
    .B(_1272_));
 sg13g2_xnor2_1 _2849_ (.Y(_1275_),
    .A(_1265_),
    .B(_1274_));
 sg13g2_nor2b_1 _2850_ (.A(_1275_),
    .B_N(_1259_),
    .Y(_1276_));
 sg13g2_xor2_1 _2851_ (.B(_1275_),
    .A(_1259_),
    .X(_1277_));
 sg13g2_nor2b_1 _2852_ (.A(_1277_),
    .B_N(_1258_),
    .Y(_1278_));
 sg13g2_xor2_1 _2853_ (.B(_1277_),
    .A(_1258_),
    .X(_1279_));
 sg13g2_nor2b_1 _2854_ (.A(_1279_),
    .B_N(_1257_),
    .Y(_1280_));
 sg13g2_xor2_1 _2855_ (.B(_1279_),
    .A(_1257_),
    .X(_1281_));
 sg13g2_inv_1 _2856_ (.Y(_1282_),
    .A(_1281_));
 sg13g2_xnor2_1 _2857_ (.Y(_1283_),
    .A(_1256_),
    .B(_1282_));
 sg13g2_nor2_1 _2858_ (.A(net416),
    .B(_1283_),
    .Y(_1284_));
 sg13g2_xor2_1 _2859_ (.B(_1283_),
    .A(net416),
    .X(_1285_));
 sg13g2_xor2_1 _2860_ (.B(_1285_),
    .A(_1255_),
    .X(_1286_));
 sg13g2_xnor2_1 _2861_ (.Y(_1287_),
    .A(_1255_),
    .B(_1285_));
 sg13g2_nor2_1 _2862_ (.A(_0016_),
    .B(_1287_),
    .Y(_1288_));
 sg13g2_xnor2_1 _2863_ (.Y(_1289_),
    .A(_1225_),
    .B(_1252_));
 sg13g2_xnor2_1 _2864_ (.Y(_1290_),
    .A(_1225_),
    .B(_1253_));
 sg13g2_and2_1 _2865_ (.A(net407),
    .B(_1289_),
    .X(_1291_));
 sg13g2_nand2_1 _2866_ (.Y(_1292_),
    .A(net407),
    .B(_1286_));
 sg13g2_nor2_1 _2867_ (.A(_0016_),
    .B(_1290_),
    .Y(_1293_));
 sg13g2_a21oi_2 _2868_ (.B1(_1284_),
    .Y(_1294_),
    .A2(_1285_),
    .A1(_1255_));
 sg13g2_o21ai_1 _2869_ (.B1(_1273_),
    .Y(_1295_),
    .A1(_1265_),
    .A2(_1274_));
 sg13g2_o21ai_1 _2870_ (.B1(_1271_),
    .Y(_1296_),
    .A1(_1233_),
    .A2(_1269_));
 sg13g2_nand2_1 _2871_ (.Y(_1297_),
    .A(net356),
    .B(net399));
 sg13g2_nand2_1 _2872_ (.Y(_1298_),
    .A(net359),
    .B(net395));
 sg13g2_nand2_1 _2873_ (.Y(_1299_),
    .A(net359),
    .B(net397));
 sg13g2_xor2_1 _2874_ (.B(_1299_),
    .A(_1268_),
    .X(_1300_));
 sg13g2_nand2b_1 _2875_ (.Y(_1301_),
    .B(_1300_),
    .A_N(_1297_));
 sg13g2_xnor2_1 _2876_ (.Y(_1302_),
    .A(_1297_),
    .B(_1300_));
 sg13g2_nand2_1 _2877_ (.Y(_1303_),
    .A(_1296_),
    .B(_1302_));
 sg13g2_xnor2_1 _2878_ (.Y(_1304_),
    .A(_1296_),
    .B(_1302_));
 sg13g2_xor2_1 _2879_ (.B(_1304_),
    .A(_1260_),
    .X(_1305_));
 sg13g2_nand2_1 _2880_ (.Y(_1306_),
    .A(_1295_),
    .B(_1305_));
 sg13g2_xnor2_1 _2881_ (.Y(_1307_),
    .A(_1295_),
    .B(_1305_));
 sg13g2_xnor2_1 _2882_ (.Y(_1308_),
    .A(_1262_),
    .B(_1307_));
 sg13g2_nor3_1 _2883_ (.A(_1276_),
    .B(_1278_),
    .C(_1308_),
    .Y(_1309_));
 sg13g2_o21ai_1 _2884_ (.B1(_1308_),
    .Y(_1310_),
    .A1(_1276_),
    .A2(_1278_));
 sg13g2_nand2b_1 _2885_ (.Y(_1311_),
    .B(_1310_),
    .A_N(_1309_));
 sg13g2_a21oi_1 _2886_ (.A1(_1256_),
    .A2(_1282_),
    .Y(_1312_),
    .B1(_1280_));
 sg13g2_xnor2_1 _2887_ (.Y(_1313_),
    .A(_1311_),
    .B(_1312_));
 sg13g2_xnor2_1 _2888_ (.Y(_1314_),
    .A(_1014_),
    .B(_1313_));
 sg13g2_xor2_1 _2889_ (.B(_1314_),
    .A(_1294_),
    .X(_1315_));
 sg13g2_nand2_1 _2890_ (.Y(_1316_),
    .A(net409),
    .B(_1315_));
 sg13g2_xnor2_1 _2891_ (.Y(_1317_),
    .A(_1292_),
    .B(_1293_));
 sg13g2_nor2b_1 _2892_ (.A(_1316_),
    .B_N(_1317_),
    .Y(_1318_));
 sg13g2_a21oi_1 _2893_ (.A1(_1288_),
    .A2(_1291_),
    .Y(_1319_),
    .B1(_1318_));
 sg13g2_or2_1 _2894_ (.X(_1320_),
    .B(_1313_),
    .A(\system_inst.neuron.u[6] ));
 sg13g2_o21ai_1 _2895_ (.B1(_1320_),
    .Y(_1321_),
    .A1(_1294_),
    .A2(_1314_));
 sg13g2_o21ai_1 _2896_ (.B1(_1310_),
    .Y(_1322_),
    .A1(_1309_),
    .A2(_1312_));
 sg13g2_o21ai_1 _2897_ (.B1(_1306_),
    .Y(_1323_),
    .A1(_1261_),
    .A2(_1307_));
 sg13g2_o21ai_1 _2898_ (.B1(_1303_),
    .Y(_1324_),
    .A1(_1260_),
    .A2(_1304_));
 sg13g2_o21ai_1 _2899_ (.B1(_1301_),
    .Y(_1325_),
    .A1(_1268_),
    .A2(_1299_));
 sg13g2_nand2_1 _2900_ (.Y(_1326_),
    .A(net353),
    .B(net399));
 sg13g2_nand2_1 _2901_ (.Y(_1327_),
    .A(net356),
    .B(net397));
 sg13g2_xor2_1 _2902_ (.B(_1327_),
    .A(_1298_),
    .X(_1328_));
 sg13g2_xnor2_1 _2903_ (.Y(_1329_),
    .A(_1326_),
    .B(_1328_));
 sg13g2_xnor2_1 _2904_ (.Y(_1330_),
    .A(_1325_),
    .B(_1329_));
 sg13g2_xnor2_1 _2905_ (.Y(_1331_),
    .A(_1324_),
    .B(_1330_));
 sg13g2_xnor2_1 _2906_ (.Y(_1332_),
    .A(_1323_),
    .B(_1331_));
 sg13g2_xnor2_1 _2907_ (.Y(_1333_),
    .A(_1322_),
    .B(_1332_));
 sg13g2_xor2_1 _2908_ (.B(_1333_),
    .A(_0010_),
    .X(_1334_));
 sg13g2_xor2_1 _2909_ (.B(_1334_),
    .A(_1321_),
    .X(_1335_));
 sg13g2_nand2_1 _2910_ (.Y(_1336_),
    .A(net409),
    .B(_1335_));
 sg13g2_and2_1 _2911_ (.A(_1024_),
    .B(_1315_),
    .X(_1337_));
 sg13g2_nand2_1 _2912_ (.Y(_1338_),
    .A(net407),
    .B(_1315_));
 sg13g2_nor2b_1 _2913_ (.A(_1292_),
    .B_N(_1337_),
    .Y(_1339_));
 sg13g2_xor2_1 _2914_ (.B(_1338_),
    .A(_1288_),
    .X(_1340_));
 sg13g2_nor2_1 _2915_ (.A(_1336_),
    .B(_1340_),
    .Y(_1341_));
 sg13g2_xor2_1 _2916_ (.B(_1340_),
    .A(_1336_),
    .X(_1342_));
 sg13g2_nor2b_1 _2917_ (.A(_1319_),
    .B_N(_1342_),
    .Y(_1343_));
 sg13g2_a22oi_1 _2918_ (.Y(_1344_),
    .B1(_1334_),
    .B2(_1321_),
    .A2(_1333_),
    .A1(_0954_));
 sg13g2_or3_2 _2919_ (.A(net415),
    .B(\system_inst.neuron.u[8] ),
    .C(_1344_),
    .X(_1345_));
 sg13g2_nand2_2 _2920_ (.Y(_1346_),
    .A(net414),
    .B(_1345_));
 sg13g2_inv_1 _2921_ (.Y(_1347_),
    .A(_1346_));
 sg13g2_nor2b_1 _2922_ (.A(_1344_),
    .B_N(_0008_),
    .Y(_1348_));
 sg13g2_xnor2_1 _2923_ (.Y(_1349_),
    .A(_0008_),
    .B(_1344_));
 sg13g2_and2_1 _2924_ (.A(_1034_),
    .B(_1349_),
    .X(_1350_));
 sg13g2_xnor2_1 _2925_ (.Y(_1351_),
    .A(net415),
    .B(_1348_));
 sg13g2_and3_1 _2926_ (.X(_1352_),
    .A(_1035_),
    .B(_1350_),
    .C(_1351_));
 sg13g2_a21oi_1 _2927_ (.A1(_1035_),
    .A2(_1351_),
    .Y(_1353_),
    .B1(_1350_));
 sg13g2_nor2_1 _2928_ (.A(_1352_),
    .B(_1353_),
    .Y(_1354_));
 sg13g2_xnor2_1 _2929_ (.Y(_1355_),
    .A(_1346_),
    .B(_1354_));
 sg13g2_xor2_1 _2930_ (.B(_1342_),
    .A(_1319_),
    .X(_1356_));
 sg13g2_inv_1 _2931_ (.Y(_1357_),
    .A(_1356_));
 sg13g2_a21oi_1 _2932_ (.A1(_1355_),
    .A2(_1357_),
    .Y(_1358_),
    .B1(_1343_));
 sg13g2_nand3_1 _2933_ (.B(_1034_),
    .C(_1345_),
    .A(net410),
    .Y(_1359_));
 sg13g2_inv_1 _2934_ (.Y(_1360_),
    .A(_1359_));
 sg13g2_a22oi_1 _2935_ (.Y(_1361_),
    .B1(net326),
    .B2(_1034_),
    .A2(_1345_),
    .A1(net410));
 sg13g2_a21oi_1 _2936_ (.A1(net326),
    .A2(_1360_),
    .Y(_1362_),
    .B1(_1361_));
 sg13g2_xnor2_1 _2937_ (.Y(_1363_),
    .A(_1346_),
    .B(_1362_));
 sg13g2_nor2_1 _2938_ (.A(_1339_),
    .B(_1341_),
    .Y(_1364_));
 sg13g2_nand2_1 _2939_ (.Y(_1365_),
    .A(net409),
    .B(net327));
 sg13g2_and2_1 _2940_ (.A(_1024_),
    .B(_1335_),
    .X(_1366_));
 sg13g2_nor2b_1 _2941_ (.A(_1338_),
    .B_N(_1366_),
    .Y(_1367_));
 sg13g2_a21oi_1 _2942_ (.A1(net407),
    .A2(_1335_),
    .Y(_1368_),
    .B1(_1337_));
 sg13g2_or2_1 _2943_ (.X(_1369_),
    .B(_1368_),
    .A(_1367_));
 sg13g2_nor2_1 _2944_ (.A(_1365_),
    .B(_1369_),
    .Y(_1370_));
 sg13g2_xor2_1 _2945_ (.B(_1369_),
    .A(_1365_),
    .X(_1371_));
 sg13g2_nor2b_1 _2946_ (.A(_1364_),
    .B_N(_1371_),
    .Y(_1372_));
 sg13g2_xnor2_1 _2947_ (.Y(_1373_),
    .A(_1364_),
    .B(_1371_));
 sg13g2_xnor2_1 _2948_ (.Y(_1374_),
    .A(_1363_),
    .B(_1373_));
 sg13g2_nor2_1 _2949_ (.A(_1358_),
    .B(_1374_),
    .Y(_1375_));
 sg13g2_a21o_1 _2950_ (.A2(_1354_),
    .A1(_1347_),
    .B1(_1352_),
    .X(_1376_));
 sg13g2_xor2_1 _2951_ (.B(_1374_),
    .A(_1358_),
    .X(_1377_));
 sg13g2_a21oi_1 _2952_ (.A1(_1376_),
    .A2(_1377_),
    .Y(_1378_),
    .B1(_1375_));
 sg13g2_a22oi_1 _2953_ (.Y(_1379_),
    .B1(_1362_),
    .B2(_1347_),
    .A2(_1360_),
    .A1(net326));
 sg13g2_a21oi_1 _2954_ (.A1(_1363_),
    .A2(_1373_),
    .Y(_1380_),
    .B1(_1372_));
 sg13g2_o21ai_1 _2955_ (.B1(_1345_),
    .Y(_1381_),
    .A1(net410),
    .A2(_1034_));
 sg13g2_nor2_1 _2956_ (.A(_1360_),
    .B(_1381_),
    .Y(_1382_));
 sg13g2_xnor2_1 _2957_ (.Y(_1383_),
    .A(_1346_),
    .B(_1382_));
 sg13g2_nor2_1 _2958_ (.A(_1367_),
    .B(_1370_),
    .Y(_1384_));
 sg13g2_nand2_1 _2959_ (.Y(_1385_),
    .A(net409),
    .B(net326));
 sg13g2_nand3_1 _2960_ (.B(net327),
    .C(_1366_),
    .A(net407),
    .Y(_1386_));
 sg13g2_a21o_1 _2961_ (.A2(net327),
    .A1(net407),
    .B1(_1366_),
    .X(_1387_));
 sg13g2_and2_1 _2962_ (.A(_1386_),
    .B(_1387_),
    .X(_1388_));
 sg13g2_nand2b_1 _2963_ (.Y(_1389_),
    .B(_1388_),
    .A_N(_1385_));
 sg13g2_xnor2_1 _2964_ (.Y(_1390_),
    .A(_1385_),
    .B(_1388_));
 sg13g2_nor2b_1 _2965_ (.A(_1384_),
    .B_N(_1390_),
    .Y(_1391_));
 sg13g2_xnor2_1 _2966_ (.Y(_1392_),
    .A(_1384_),
    .B(_1390_));
 sg13g2_xnor2_1 _2967_ (.Y(_1393_),
    .A(_1383_),
    .B(_1392_));
 sg13g2_xor2_1 _2968_ (.B(_1393_),
    .A(_1380_),
    .X(_1394_));
 sg13g2_nand2b_1 _2969_ (.Y(_1395_),
    .B(_1394_),
    .A_N(_1379_));
 sg13g2_xnor2_1 _2970_ (.Y(_1396_),
    .A(_1379_),
    .B(_1394_));
 sg13g2_nand2b_1 _2971_ (.Y(_1397_),
    .B(_1396_),
    .A_N(_1378_));
 sg13g2_xnor2_1 _2972_ (.Y(_1398_),
    .A(_1222_),
    .B(_1224_));
 sg13g2_xor2_1 _2973_ (.B(_1224_),
    .A(_1222_),
    .X(_1399_));
 sg13g2_nor2_2 _2974_ (.A(_0016_),
    .B(_1399_),
    .Y(_1400_));
 sg13g2_nand2_1 _2975_ (.Y(_1401_),
    .A(net409),
    .B(_1286_));
 sg13g2_xor2_1 _2976_ (.B(_1400_),
    .A(_1291_),
    .X(_1402_));
 sg13g2_nor2b_1 _2977_ (.A(_1401_),
    .B_N(_1402_),
    .Y(_1403_));
 sg13g2_a21oi_1 _2978_ (.A1(_1291_),
    .A2(_1400_),
    .Y(_1404_),
    .B1(_1403_));
 sg13g2_xnor2_1 _2979_ (.Y(_1405_),
    .A(_1316_),
    .B(_1317_));
 sg13g2_nor2b_1 _2980_ (.A(_1404_),
    .B_N(_1405_),
    .Y(_1406_));
 sg13g2_and2_1 _2981_ (.A(\system_inst.internal_param_a[2] ),
    .B(_1335_),
    .X(_1407_));
 sg13g2_nand3_1 _2982_ (.B(_1349_),
    .C(_1407_),
    .A(net410),
    .Y(_1408_));
 sg13g2_a21o_1 _2983_ (.A2(net327),
    .A1(net410),
    .B1(_1407_),
    .X(_1409_));
 sg13g2_and4_1 _2984_ (.A(net413),
    .B(net326),
    .C(_1408_),
    .D(_1409_),
    .X(_1410_));
 sg13g2_nand4_1 _2985_ (.B(net326),
    .C(_1408_),
    .A(net413),
    .Y(_1411_),
    .D(_1409_));
 sg13g2_a22oi_1 _2986_ (.Y(_1412_),
    .B1(_1408_),
    .B2(_1409_),
    .A2(net326),
    .A1(net413));
 sg13g2_xnor2_1 _2987_ (.Y(_1413_),
    .A(_1404_),
    .B(_1405_));
 sg13g2_inv_1 _2988_ (.Y(_1414_),
    .A(_1413_));
 sg13g2_nor3_1 _2989_ (.A(_1410_),
    .B(_1412_),
    .C(_1414_),
    .Y(_1415_));
 sg13g2_nor2_1 _2990_ (.A(_1406_),
    .B(_1415_),
    .Y(_1416_));
 sg13g2_xnor2_1 _2991_ (.Y(_1417_),
    .A(_1355_),
    .B(_1357_));
 sg13g2_nor2_1 _2992_ (.A(_1416_),
    .B(_1417_),
    .Y(_1418_));
 sg13g2_nand2_1 _2993_ (.Y(_1419_),
    .A(_1408_),
    .B(_1411_));
 sg13g2_xor2_1 _2994_ (.B(_1417_),
    .A(_1416_),
    .X(_1420_));
 sg13g2_a21oi_1 _2995_ (.A1(_1419_),
    .A2(_1420_),
    .Y(_1421_),
    .B1(_1418_));
 sg13g2_xnor2_1 _2996_ (.Y(_1422_),
    .A(_1376_),
    .B(_1377_));
 sg13g2_or2_1 _2997_ (.X(_1423_),
    .B(_1422_),
    .A(_1421_));
 sg13g2_xor2_1 _2998_ (.B(_1220_),
    .A(_1218_),
    .X(_1424_));
 sg13g2_and2_1 _2999_ (.A(net406),
    .B(_1424_),
    .X(_1425_));
 sg13g2_nor2_1 _3000_ (.A(_0900_),
    .B(_1290_),
    .Y(_1426_));
 sg13g2_a22oi_1 _3001_ (.Y(_1427_),
    .B1(_1424_),
    .B2(_1024_),
    .A2(_1398_),
    .A1(net406));
 sg13g2_a21oi_1 _3002_ (.A1(_1400_),
    .A2(_1425_),
    .Y(_1428_),
    .B1(_1427_));
 sg13g2_a22oi_1 _3003_ (.Y(_1429_),
    .B1(_1426_),
    .B2(_1428_),
    .A2(_1425_),
    .A1(_1400_));
 sg13g2_xnor2_1 _3004_ (.Y(_1430_),
    .A(_1401_),
    .B(_1402_));
 sg13g2_nand2b_1 _3005_ (.Y(_1431_),
    .B(_1430_),
    .A_N(_1429_));
 sg13g2_and2_1 _3006_ (.A(\system_inst.internal_param_a[2] ),
    .B(_1315_),
    .X(_1432_));
 sg13g2_nand3_1 _3007_ (.B(_1335_),
    .C(_1432_),
    .A(\system_inst.internal_param_a[1] ),
    .Y(_1433_));
 sg13g2_a21o_1 _3008_ (.A2(_1335_),
    .A1(\system_inst.internal_param_a[1] ),
    .B1(_1432_),
    .X(_1434_));
 sg13g2_and4_1 _3009_ (.A(net414),
    .B(net327),
    .C(_1433_),
    .D(_1434_),
    .X(_1435_));
 sg13g2_nand4_1 _3010_ (.B(net327),
    .C(_1433_),
    .A(net413),
    .Y(_1436_),
    .D(_1434_));
 sg13g2_a22oi_1 _3011_ (.Y(_1437_),
    .B1(_1433_),
    .B2(_1434_),
    .A2(net327),
    .A1(net414));
 sg13g2_xor2_1 _3012_ (.B(_1430_),
    .A(_1429_),
    .X(_1438_));
 sg13g2_or3_1 _3013_ (.A(_1435_),
    .B(_1437_),
    .C(_1438_),
    .X(_1439_));
 sg13g2_nand2_1 _3014_ (.Y(_1440_),
    .A(_1431_),
    .B(_1439_));
 sg13g2_o21ai_1 _3015_ (.B1(_1414_),
    .Y(_1441_),
    .A1(_1410_),
    .A2(_1412_));
 sg13g2_nor2b_1 _3016_ (.A(_1415_),
    .B_N(_1441_),
    .Y(_1442_));
 sg13g2_nand2_1 _3017_ (.Y(_1443_),
    .A(_1440_),
    .B(_1442_));
 sg13g2_nand2_1 _3018_ (.Y(_1444_),
    .A(_1433_),
    .B(_1436_));
 sg13g2_xor2_1 _3019_ (.B(_1442_),
    .A(_1440_),
    .X(_1445_));
 sg13g2_nand2_1 _3020_ (.Y(_1446_),
    .A(_1444_),
    .B(_1445_));
 sg13g2_and2_1 _3021_ (.A(_1443_),
    .B(_1446_),
    .X(_1447_));
 sg13g2_xnor2_1 _3022_ (.Y(_1448_),
    .A(_1419_),
    .B(_1420_));
 sg13g2_nor2_1 _3023_ (.A(_1447_),
    .B(_1448_),
    .Y(_1449_));
 sg13g2_xor2_1 _3024_ (.B(_1217_),
    .A(_1215_),
    .X(_1450_));
 sg13g2_nand2_1 _3025_ (.Y(_1451_),
    .A(net406),
    .B(_1450_));
 sg13g2_and2_1 _3026_ (.A(_1024_),
    .B(_1450_),
    .X(_1452_));
 sg13g2_nand2_1 _3027_ (.Y(_1453_),
    .A(net409),
    .B(_1398_));
 sg13g2_xor2_1 _3028_ (.B(_1452_),
    .A(_1425_),
    .X(_1454_));
 sg13g2_nor2b_1 _3029_ (.A(_1453_),
    .B_N(_1454_),
    .Y(_1455_));
 sg13g2_a21oi_1 _3030_ (.A1(_1425_),
    .A2(_1452_),
    .Y(_1456_),
    .B1(_1455_));
 sg13g2_xor2_1 _3031_ (.B(_1428_),
    .A(_1426_),
    .X(_1457_));
 sg13g2_nand2b_1 _3032_ (.Y(_1458_),
    .B(_1457_),
    .A_N(_1456_));
 sg13g2_nor2_2 _3033_ (.A(_0922_),
    .B(_1287_),
    .Y(_1459_));
 sg13g2_nor2_1 _3034_ (.A(_0911_),
    .B(_1287_),
    .Y(_1460_));
 sg13g2_nand2_1 _3035_ (.Y(_1461_),
    .A(_1432_),
    .B(_1459_));
 sg13g2_a21o_1 _3036_ (.A2(_1315_),
    .A1(net410),
    .B1(_1460_),
    .X(_1462_));
 sg13g2_and4_1 _3037_ (.A(net413),
    .B(_1335_),
    .C(_1461_),
    .D(_1462_),
    .X(_1463_));
 sg13g2_a22oi_1 _3038_ (.Y(_1464_),
    .B1(_1461_),
    .B2(_1462_),
    .A2(_1335_),
    .A1(net413));
 sg13g2_xor2_1 _3039_ (.B(_1457_),
    .A(_1456_),
    .X(_1465_));
 sg13g2_or3_1 _3040_ (.A(_1463_),
    .B(_1464_),
    .C(_1465_),
    .X(_1466_));
 sg13g2_nand2_1 _3041_ (.Y(_1467_),
    .A(_1458_),
    .B(_1466_));
 sg13g2_o21ai_1 _3042_ (.B1(_1438_),
    .Y(_1468_),
    .A1(_1435_),
    .A2(_1437_));
 sg13g2_nand3_1 _3043_ (.B(_1467_),
    .C(_1468_),
    .A(_1439_),
    .Y(_1469_));
 sg13g2_a21o_1 _3044_ (.A2(_1459_),
    .A1(_1432_),
    .B1(_1463_),
    .X(_1470_));
 sg13g2_inv_1 _3045_ (.Y(_1471_),
    .A(_1470_));
 sg13g2_a21oi_1 _3046_ (.A1(_1439_),
    .A2(_1468_),
    .Y(_1472_),
    .B1(_1467_));
 sg13g2_a21o_1 _3047_ (.A2(_1468_),
    .A1(_1439_),
    .B1(_1467_),
    .X(_1473_));
 sg13g2_and3_1 _3048_ (.X(_1474_),
    .A(_1469_),
    .B(_1470_),
    .C(_1473_));
 sg13g2_o21ai_1 _3049_ (.B1(_1469_),
    .Y(_1475_),
    .A1(_1471_),
    .A2(_1472_));
 sg13g2_or2_1 _3050_ (.X(_1476_),
    .B(_1445_),
    .A(_1444_));
 sg13g2_and3_1 _3051_ (.X(_1477_),
    .A(_1446_),
    .B(_1475_),
    .C(_1476_));
 sg13g2_nand3_1 _3052_ (.B(_1475_),
    .C(_1476_),
    .A(_1446_),
    .Y(_1478_));
 sg13g2_xor2_1 _3053_ (.B(_1214_),
    .A(\system_inst.neuron.u[0] ),
    .X(_1479_));
 sg13g2_nand2_1 _3054_ (.Y(_1480_),
    .A(net406),
    .B(net328));
 sg13g2_nand2_1 _3055_ (.Y(_1481_),
    .A(_1024_),
    .B(net328));
 sg13g2_nor2_1 _3056_ (.A(_1451_),
    .B(_1481_),
    .Y(_1482_));
 sg13g2_nand2_1 _3057_ (.Y(_1483_),
    .A(net408),
    .B(_1424_));
 sg13g2_xor2_1 _3058_ (.B(_1481_),
    .A(_1451_),
    .X(_1484_));
 sg13g2_nor2b_1 _3059_ (.A(_1483_),
    .B_N(_1484_),
    .Y(_1485_));
 sg13g2_nor2_1 _3060_ (.A(_1482_),
    .B(_1485_),
    .Y(_1486_));
 sg13g2_xnor2_1 _3061_ (.Y(_1487_),
    .A(_1453_),
    .B(_1454_));
 sg13g2_nor2b_1 _3062_ (.A(_1486_),
    .B_N(_1487_),
    .Y(_1488_));
 sg13g2_nor2_1 _3063_ (.A(_0911_),
    .B(_1290_),
    .Y(_1489_));
 sg13g2_nand2_1 _3064_ (.Y(_1490_),
    .A(_1459_),
    .B(_1489_));
 sg13g2_or2_1 _3065_ (.X(_1491_),
    .B(_1489_),
    .A(_1459_));
 sg13g2_and4_1 _3066_ (.A(net413),
    .B(_1315_),
    .C(_1490_),
    .D(_1491_),
    .X(_1492_));
 sg13g2_a22oi_1 _3067_ (.Y(_1493_),
    .B1(_1490_),
    .B2(_1491_),
    .A2(_1315_),
    .A1(net413));
 sg13g2_xor2_1 _3068_ (.B(_1487_),
    .A(_1486_),
    .X(_1494_));
 sg13g2_or3_1 _3069_ (.A(_1492_),
    .B(_1493_),
    .C(_1494_),
    .X(_1495_));
 sg13g2_nand2b_1 _3070_ (.Y(_1496_),
    .B(_1495_),
    .A_N(_1488_));
 sg13g2_o21ai_1 _3071_ (.B1(_1465_),
    .Y(_1497_),
    .A1(_1463_),
    .A2(_1464_));
 sg13g2_nand3_1 _3072_ (.B(_1496_),
    .C(_1497_),
    .A(_1466_),
    .Y(_1498_));
 sg13g2_a21o_1 _3073_ (.A2(_1489_),
    .A1(_1459_),
    .B1(_1492_),
    .X(_1499_));
 sg13g2_a21o_1 _3074_ (.A2(_1497_),
    .A1(_1466_),
    .B1(_1496_),
    .X(_1500_));
 sg13g2_nand3_1 _3075_ (.B(_1499_),
    .C(_1500_),
    .A(_1498_),
    .Y(_1501_));
 sg13g2_and2_1 _3076_ (.A(_1498_),
    .B(_1501_),
    .X(_1502_));
 sg13g2_a21oi_1 _3077_ (.A1(_1469_),
    .A2(_1473_),
    .Y(_1503_),
    .B1(_1470_));
 sg13g2_nor3_1 _3078_ (.A(_1474_),
    .B(_1502_),
    .C(_1503_),
    .Y(_1504_));
 sg13g2_xnor2_1 _3079_ (.Y(_1505_),
    .A(_1169_),
    .B(_1176_));
 sg13g2_a21oi_1 _3080_ (.A1(_1168_),
    .A2(_1505_),
    .Y(_1506_),
    .B1(_1170_));
 sg13g2_nand2_1 _3081_ (.Y(_1507_),
    .A(\system_inst.internal_param_a[5] ),
    .B(net329));
 sg13g2_nand2_1 _3082_ (.Y(_1508_),
    .A(net408),
    .B(_1450_));
 sg13g2_xor2_1 _3083_ (.B(_1507_),
    .A(_1480_),
    .X(_1509_));
 sg13g2_nand2b_1 _3084_ (.Y(_1510_),
    .B(_1509_),
    .A_N(_1508_));
 sg13g2_o21ai_1 _3085_ (.B1(_1510_),
    .Y(_1511_),
    .A1(_1480_),
    .A2(_1507_));
 sg13g2_xnor2_1 _3086_ (.Y(_1512_),
    .A(_1483_),
    .B(_1484_));
 sg13g2_nand2_1 _3087_ (.Y(_1513_),
    .A(net411),
    .B(_1398_));
 sg13g2_nor2_1 _3088_ (.A(_0911_),
    .B(_1399_),
    .Y(_1514_));
 sg13g2_nor3_1 _3089_ (.A(_0911_),
    .B(_1290_),
    .C(_1513_),
    .Y(_1515_));
 sg13g2_nand3_1 _3090_ (.B(_1289_),
    .C(_1514_),
    .A(net411),
    .Y(_1516_));
 sg13g2_a21o_1 _3091_ (.A2(_1289_),
    .A1(net411),
    .B1(_1514_),
    .X(_1517_));
 sg13g2_and4_1 _3092_ (.A(net412),
    .B(_1286_),
    .C(_1516_),
    .D(_1517_),
    .X(_1518_));
 sg13g2_a22oi_1 _3093_ (.Y(_1519_),
    .B1(_1516_),
    .B2(_1517_),
    .A2(_1286_),
    .A1(net414));
 sg13g2_nor2_1 _3094_ (.A(_1518_),
    .B(_1519_),
    .Y(_1520_));
 sg13g2_xnor2_1 _3095_ (.Y(_1521_),
    .A(_1511_),
    .B(_1512_));
 sg13g2_nor3_1 _3096_ (.A(_1518_),
    .B(_1519_),
    .C(_1521_),
    .Y(_1522_));
 sg13g2_a21o_1 _3097_ (.A2(_1512_),
    .A1(_1511_),
    .B1(_1522_),
    .X(_1523_));
 sg13g2_o21ai_1 _3098_ (.B1(_1494_),
    .Y(_1524_),
    .A1(_1492_),
    .A2(_1493_));
 sg13g2_nand3_1 _3099_ (.B(_1523_),
    .C(_1524_),
    .A(_1495_),
    .Y(_1525_));
 sg13g2_or2_1 _3100_ (.X(_1526_),
    .B(_1518_),
    .A(_1515_));
 sg13g2_inv_1 _3101_ (.Y(_1527_),
    .A(_1526_));
 sg13g2_a21oi_1 _3102_ (.A1(_1495_),
    .A2(_1524_),
    .Y(_1528_),
    .B1(_1523_));
 sg13g2_a21o_1 _3103_ (.A2(_1524_),
    .A1(_1495_),
    .B1(_1523_),
    .X(_1529_));
 sg13g2_and3_1 _3104_ (.X(_1530_),
    .A(_1525_),
    .B(_1526_),
    .C(_1529_));
 sg13g2_o21ai_1 _3105_ (.B1(_1525_),
    .Y(_1531_),
    .A1(_1527_),
    .A2(_1528_));
 sg13g2_a21o_1 _3106_ (.A2(_1500_),
    .A1(_1498_),
    .B1(_1499_),
    .X(_1532_));
 sg13g2_and3_1 _3107_ (.X(_1533_),
    .A(_1501_),
    .B(_1531_),
    .C(_1532_));
 sg13g2_nand3_1 _3108_ (.B(_1531_),
    .C(_1532_),
    .A(_1501_),
    .Y(_1534_));
 sg13g2_xnor2_1 _3109_ (.Y(_1535_),
    .A(_1171_),
    .B(_1175_));
 sg13g2_and2_1 _3110_ (.A(_1024_),
    .B(_1535_),
    .X(_1536_));
 sg13g2_nand3_1 _3111_ (.B(net329),
    .C(_1536_),
    .A(net406),
    .Y(_1537_));
 sg13g2_a21o_1 _3112_ (.A2(_1506_),
    .A1(net406),
    .B1(_1536_),
    .X(_1538_));
 sg13g2_and2_1 _3113_ (.A(_1537_),
    .B(_1538_),
    .X(_1539_));
 sg13g2_nand3_1 _3114_ (.B(net328),
    .C(_1539_),
    .A(net408),
    .Y(_1540_));
 sg13g2_and2_1 _3115_ (.A(_1537_),
    .B(_1540_),
    .X(_1541_));
 sg13g2_xnor2_1 _3116_ (.Y(_1542_),
    .A(_1508_),
    .B(_1509_));
 sg13g2_nand2b_1 _3117_ (.Y(_1543_),
    .B(_1542_),
    .A_N(_1541_));
 sg13g2_xnor2_1 _3118_ (.Y(_1544_),
    .A(_1541_),
    .B(_1542_));
 sg13g2_inv_1 _3119_ (.Y(_1545_),
    .A(_1544_));
 sg13g2_nand2_1 _3120_ (.Y(_1546_),
    .A(\system_inst.internal_param_a[2] ),
    .B(_1424_));
 sg13g2_or2_1 _3121_ (.X(_1547_),
    .B(_1546_),
    .A(_1513_));
 sg13g2_nand2_1 _3122_ (.Y(_1548_),
    .A(_1513_),
    .B(_1546_));
 sg13g2_and4_1 _3123_ (.A(net412),
    .B(_1289_),
    .C(_1547_),
    .D(_1548_),
    .X(_1549_));
 sg13g2_nand4_1 _3124_ (.B(_1289_),
    .C(_1547_),
    .A(net412),
    .Y(_1550_),
    .D(_1548_));
 sg13g2_a22oi_1 _3125_ (.Y(_1551_),
    .B1(_1547_),
    .B2(_1548_),
    .A2(_1289_),
    .A1(net412));
 sg13g2_nand3b_1 _3126_ (.B(_1544_),
    .C(_1550_),
    .Y(_1552_),
    .A_N(_1551_));
 sg13g2_and2_1 _3127_ (.A(_1543_),
    .B(_1552_),
    .X(_1553_));
 sg13g2_nor2b_1 _3128_ (.A(_1520_),
    .B_N(_1521_),
    .Y(_1554_));
 sg13g2_nor3_1 _3129_ (.A(_1522_),
    .B(_1553_),
    .C(_1554_),
    .Y(_1555_));
 sg13g2_nand2_1 _3130_ (.Y(_1556_),
    .A(_1547_),
    .B(_1550_));
 sg13g2_o21ai_1 _3131_ (.B1(_1553_),
    .Y(_1557_),
    .A1(_1522_),
    .A2(_1554_));
 sg13g2_nor2b_1 _3132_ (.A(_1555_),
    .B_N(_1557_),
    .Y(_1558_));
 sg13g2_a21oi_1 _3133_ (.A1(_1556_),
    .A2(_1557_),
    .Y(_1559_),
    .B1(_1555_));
 sg13g2_a21oi_1 _3134_ (.A1(_1525_),
    .A2(_1529_),
    .Y(_1560_),
    .B1(_1526_));
 sg13g2_nor3_1 _3135_ (.A(_1530_),
    .B(_1559_),
    .C(_1560_),
    .Y(_1561_));
 sg13g2_nand2_1 _3136_ (.Y(_1562_),
    .A(net408),
    .B(_1535_));
 sg13g2_and2_1 _3137_ (.A(net406),
    .B(_1535_),
    .X(_1563_));
 sg13g2_nand3_1 _3138_ (.B(net329),
    .C(_1563_),
    .A(net408),
    .Y(_1564_));
 sg13g2_a21o_1 _3139_ (.A2(net328),
    .A1(net408),
    .B1(_1539_),
    .X(_1565_));
 sg13g2_and2_1 _3140_ (.A(_1540_),
    .B(_1565_),
    .X(_1566_));
 sg13g2_nor2b_1 _3141_ (.A(_1564_),
    .B_N(_1566_),
    .Y(_1567_));
 sg13g2_xnor2_1 _3142_ (.Y(_1568_),
    .A(_1564_),
    .B(_1566_));
 sg13g2_nor2_1 _3143_ (.A(_0933_),
    .B(_1399_),
    .Y(_1569_));
 sg13g2_nand2_1 _3144_ (.Y(_1570_),
    .A(net411),
    .B(_1450_));
 sg13g2_nor2_1 _3145_ (.A(_1546_),
    .B(_1570_),
    .Y(_1571_));
 sg13g2_a22oi_1 _3146_ (.Y(_1572_),
    .B1(_1450_),
    .B2(\system_inst.internal_param_a[2] ),
    .A2(_1424_),
    .A1(net411));
 sg13g2_nor2_1 _3147_ (.A(_1571_),
    .B(_1572_),
    .Y(_1573_));
 sg13g2_xor2_1 _3148_ (.B(_1573_),
    .A(_1569_),
    .X(_1574_));
 sg13g2_a21o_1 _3149_ (.A2(_1574_),
    .A1(_1568_),
    .B1(_1567_),
    .X(_1575_));
 sg13g2_o21ai_1 _3150_ (.B1(_1545_),
    .Y(_1576_),
    .A1(_1549_),
    .A2(_1551_));
 sg13g2_nand3_1 _3151_ (.B(_1575_),
    .C(_1576_),
    .A(_1552_),
    .Y(_1577_));
 sg13g2_a21oi_1 _3152_ (.A1(_1569_),
    .A2(_1573_),
    .Y(_1578_),
    .B1(_1571_));
 sg13g2_inv_1 _3153_ (.Y(_1579_),
    .A(_1578_));
 sg13g2_a21oi_1 _3154_ (.A1(_1552_),
    .A2(_1576_),
    .Y(_1580_),
    .B1(_1575_));
 sg13g2_a21o_1 _3155_ (.A2(_1576_),
    .A1(_1552_),
    .B1(_1575_),
    .X(_1581_));
 sg13g2_and3_1 _3156_ (.X(_1582_),
    .A(_1577_),
    .B(_1579_),
    .C(_1581_));
 sg13g2_o21ai_1 _3157_ (.B1(_1577_),
    .Y(_1583_),
    .A1(_1578_),
    .A2(_1580_));
 sg13g2_xor2_1 _3158_ (.B(_1558_),
    .A(_1556_),
    .X(_1584_));
 sg13g2_nand2_1 _3159_ (.Y(_1585_),
    .A(_1583_),
    .B(_1584_));
 sg13g2_xnor2_1 _3160_ (.Y(_1586_),
    .A(_1568_),
    .B(_1574_));
 sg13g2_nand2_1 _3161_ (.Y(_1587_),
    .A(net412),
    .B(_1424_));
 sg13g2_nand2_1 _3162_ (.Y(_1588_),
    .A(net411),
    .B(_1479_));
 sg13g2_nand2_1 _3163_ (.Y(_1589_),
    .A(\system_inst.internal_param_a[2] ),
    .B(net328));
 sg13g2_xor2_1 _3164_ (.B(_1589_),
    .A(_1570_),
    .X(_1590_));
 sg13g2_nand2b_1 _3165_ (.Y(_1591_),
    .B(_1590_),
    .A_N(_1587_));
 sg13g2_xnor2_1 _3166_ (.Y(_1592_),
    .A(_1587_),
    .B(_1590_));
 sg13g2_a21o_1 _3167_ (.A2(net329),
    .A1(net408),
    .B1(_1563_),
    .X(_1593_));
 sg13g2_and2_1 _3168_ (.A(_1564_),
    .B(_1593_),
    .X(_1594_));
 sg13g2_and2_1 _3169_ (.A(_1592_),
    .B(_1594_),
    .X(_1595_));
 sg13g2_nor2b_1 _3170_ (.A(_1586_),
    .B_N(_1595_),
    .Y(_1596_));
 sg13g2_o21ai_1 _3171_ (.B1(_1591_),
    .Y(_1597_),
    .A1(_1570_),
    .A2(_1589_));
 sg13g2_xnor2_1 _3172_ (.Y(_1598_),
    .A(_1586_),
    .B(_1595_));
 sg13g2_nand2_1 _3173_ (.Y(_1599_),
    .A(_1597_),
    .B(_1598_));
 sg13g2_a21oi_1 _3174_ (.A1(_1597_),
    .A2(_1598_),
    .Y(_1600_),
    .B1(_1596_));
 sg13g2_a21oi_1 _3175_ (.A1(_1577_),
    .A2(_1581_),
    .Y(_1601_),
    .B1(_1579_));
 sg13g2_nor3_1 _3176_ (.A(_1582_),
    .B(_1600_),
    .C(_1601_),
    .Y(_1602_));
 sg13g2_nand2_1 _3177_ (.Y(_1603_),
    .A(net412),
    .B(_1450_));
 sg13g2_nand2_1 _3178_ (.Y(_1604_),
    .A(\system_inst.internal_param_a[2] ),
    .B(net329));
 sg13g2_or2_1 _3179_ (.X(_1605_),
    .B(_1604_),
    .A(_1588_));
 sg13g2_xnor2_1 _3180_ (.Y(_1606_),
    .A(_1588_),
    .B(_1604_));
 sg13g2_xnor2_1 _3181_ (.Y(_1607_),
    .A(_1603_),
    .B(_1606_));
 sg13g2_nor2_1 _3182_ (.A(_1562_),
    .B(_1607_),
    .Y(_1608_));
 sg13g2_xor2_1 _3183_ (.B(_1594_),
    .A(_1592_),
    .X(_1609_));
 sg13g2_and2_1 _3184_ (.A(_1608_),
    .B(_1609_),
    .X(_1610_));
 sg13g2_o21ai_1 _3185_ (.B1(_1605_),
    .Y(_1611_),
    .A1(_1603_),
    .A2(_1606_));
 sg13g2_and4_1 _3186_ (.A(net411),
    .B(_1034_),
    .C(net329),
    .D(_1535_),
    .X(_1612_));
 sg13g2_a22oi_1 _3187_ (.Y(_1613_),
    .B1(_1535_),
    .B2(_1034_),
    .A2(net329),
    .A1(net411));
 sg13g2_nor2_1 _3188_ (.A(_1612_),
    .B(_1613_),
    .Y(_1614_));
 sg13g2_and4_1 _3189_ (.A(net412),
    .B(_1035_),
    .C(net329),
    .D(_1535_),
    .X(_1615_));
 sg13g2_o21ai_1 _3190_ (.B1(_1615_),
    .Y(_1616_),
    .A1(net328),
    .A2(_1614_));
 sg13g2_nor2_1 _3191_ (.A(_0933_),
    .B(_1613_),
    .Y(_1617_));
 sg13g2_a21oi_1 _3192_ (.A1(net328),
    .A2(_1617_),
    .Y(_1618_),
    .B1(_1612_));
 sg13g2_nand3_1 _3193_ (.B(_1612_),
    .C(_1615_),
    .A(net328),
    .Y(_1619_));
 sg13g2_a22oi_1 _3194_ (.Y(_1620_),
    .B1(_1616_),
    .B2(_1618_),
    .A2(_1607_),
    .A1(_1562_));
 sg13g2_nand2b_1 _3195_ (.Y(_1621_),
    .B(_1620_),
    .A_N(_1608_));
 sg13g2_and2_1 _3196_ (.A(_1619_),
    .B(_1621_),
    .X(_1622_));
 sg13g2_nor2b_1 _3197_ (.A(_1622_),
    .B_N(_1611_),
    .Y(_1623_));
 sg13g2_and2_1 _3198_ (.A(_1610_),
    .B(_1623_),
    .X(_1624_));
 sg13g2_nor2_1 _3199_ (.A(_1610_),
    .B(_1611_),
    .Y(_1625_));
 sg13g2_or3_1 _3200_ (.A(_1608_),
    .B(_1609_),
    .C(_1623_),
    .X(_1626_));
 sg13g2_o21ai_1 _3201_ (.B1(_1626_),
    .Y(_1627_),
    .A1(_1597_),
    .A2(_1598_));
 sg13g2_a21oi_1 _3202_ (.A1(_1622_),
    .A2(_1625_),
    .Y(_1628_),
    .B1(_1627_));
 sg13g2_a21o_1 _3203_ (.A2(_1628_),
    .A1(_1599_),
    .B1(_1624_),
    .X(_1629_));
 sg13g2_o21ai_1 _3204_ (.B1(_1600_),
    .Y(_1630_),
    .A1(_1582_),
    .A2(_1601_));
 sg13g2_nor2b_1 _3205_ (.A(_1602_),
    .B_N(_1630_),
    .Y(_1631_));
 sg13g2_a21oi_1 _3206_ (.A1(_1629_),
    .A2(_1631_),
    .Y(_1632_),
    .B1(_1602_));
 sg13g2_xnor2_1 _3207_ (.Y(_1633_),
    .A(_1583_),
    .B(_1584_));
 sg13g2_o21ai_1 _3208_ (.B1(_1585_),
    .Y(_1634_),
    .A1(_1632_),
    .A2(_1633_));
 sg13g2_o21ai_1 _3209_ (.B1(_1559_),
    .Y(_1635_),
    .A1(_1530_),
    .A2(_1560_));
 sg13g2_nor2b_1 _3210_ (.A(_1561_),
    .B_N(_1635_),
    .Y(_1636_));
 sg13g2_a21oi_1 _3211_ (.A1(_1634_),
    .A2(_1636_),
    .Y(_1637_),
    .B1(_1561_));
 sg13g2_a21oi_1 _3212_ (.A1(_1501_),
    .A2(_1532_),
    .Y(_1638_),
    .B1(_1531_));
 sg13g2_nor2_1 _3213_ (.A(_1533_),
    .B(_1638_),
    .Y(_1639_));
 sg13g2_o21ai_1 _3214_ (.B1(_1534_),
    .Y(_1640_),
    .A1(_1637_),
    .A2(_1638_));
 sg13g2_o21ai_1 _3215_ (.B1(_1502_),
    .Y(_1641_),
    .A1(_1474_),
    .A2(_1503_));
 sg13g2_nor2b_1 _3216_ (.A(_1504_),
    .B_N(_1641_),
    .Y(_1642_));
 sg13g2_a21oi_1 _3217_ (.A1(_1640_),
    .A2(_1642_),
    .Y(_1643_),
    .B1(_1504_));
 sg13g2_a21oi_1 _3218_ (.A1(_1446_),
    .A2(_1476_),
    .Y(_1644_),
    .B1(_1475_));
 sg13g2_nor2_1 _3219_ (.A(_1477_),
    .B(_1644_),
    .Y(_1645_));
 sg13g2_o21ai_1 _3220_ (.B1(_1478_),
    .Y(_1646_),
    .A1(_1643_),
    .A2(_1644_));
 sg13g2_xor2_1 _3221_ (.B(_1448_),
    .A(_1447_),
    .X(_1647_));
 sg13g2_a21oi_1 _3222_ (.A1(_1646_),
    .A2(_1647_),
    .Y(_1648_),
    .B1(_1449_));
 sg13g2_xnor2_1 _3223_ (.Y(_1649_),
    .A(_1421_),
    .B(_1422_));
 sg13g2_o21ai_1 _3224_ (.B1(_1423_),
    .Y(_1650_),
    .A1(_1648_),
    .A2(_1649_));
 sg13g2_xnor2_1 _3225_ (.Y(_1651_),
    .A(_1378_),
    .B(_1396_));
 sg13g2_nand2_1 _3226_ (.Y(_1652_),
    .A(_1650_),
    .B(_1651_));
 sg13g2_o21ai_1 _3227_ (.B1(_1395_),
    .Y(_1653_),
    .A1(_1380_),
    .A2(_1393_));
 sg13g2_nand2_1 _3228_ (.Y(_1654_),
    .A(net406),
    .B(net326));
 sg13g2_nand2_1 _3229_ (.Y(_1655_),
    .A(_1386_),
    .B(_1389_));
 sg13g2_xor2_1 _3230_ (.B(_1655_),
    .A(_1654_),
    .X(_1656_));
 sg13g2_nand2_1 _3231_ (.Y(_1657_),
    .A(\system_inst.internal_param_a[5] ),
    .B(net327));
 sg13g2_nand2_1 _3232_ (.Y(_1658_),
    .A(net409),
    .B(_1345_));
 sg13g2_xnor2_1 _3233_ (.Y(_1659_),
    .A(_1657_),
    .B(_1658_));
 sg13g2_xnor2_1 _3234_ (.Y(_1660_),
    .A(_1383_),
    .B(_1659_));
 sg13g2_xnor2_1 _3235_ (.Y(_1661_),
    .A(_1656_),
    .B(_1660_));
 sg13g2_a21oi_1 _3236_ (.A1(_1383_),
    .A2(_1392_),
    .Y(_1662_),
    .B1(_1391_));
 sg13g2_a21o_1 _3237_ (.A2(_1382_),
    .A1(_1347_),
    .B1(_1360_),
    .X(_1663_));
 sg13g2_xnor2_1 _3238_ (.Y(_1664_),
    .A(_1662_),
    .B(_1663_));
 sg13g2_xnor2_1 _3239_ (.Y(_1665_),
    .A(_1661_),
    .B(_1664_));
 sg13g2_xnor2_1 _3240_ (.Y(_1666_),
    .A(_1653_),
    .B(_1665_));
 sg13g2_a21oi_1 _3241_ (.A1(_1397_),
    .A2(_1652_),
    .Y(_1667_),
    .B1(_1666_));
 sg13g2_xnor2_1 _3242_ (.Y(_1668_),
    .A(_1648_),
    .B(_1649_));
 sg13g2_a21o_1 _3243_ (.A2(_1666_),
    .A1(_1397_),
    .B1(_1651_),
    .X(_1669_));
 sg13g2_o21ai_1 _3244_ (.B1(_1652_),
    .Y(_1670_),
    .A1(_1650_),
    .A2(_1669_));
 sg13g2_nand3b_1 _3245_ (.B(_1668_),
    .C(_1670_),
    .Y(_1671_),
    .A_N(_1667_));
 sg13g2_xor2_1 _3246_ (.B(_1631_),
    .A(_1629_),
    .X(_1672_));
 sg13g2_or2_1 _3247_ (.X(_1673_),
    .B(_1672_),
    .A(_1671_));
 sg13g2_and2_1 _3248_ (.A(\system_inst.neuron.u[0] ),
    .B(_1673_),
    .X(_1674_));
 sg13g2_xnor2_1 _3249_ (.Y(_1675_),
    .A(_1632_),
    .B(_1633_));
 sg13g2_nand2b_1 _3250_ (.Y(_1676_),
    .B(_1675_),
    .A_N(_1671_));
 sg13g2_xor2_1 _3251_ (.B(_1676_),
    .A(net141),
    .X(_1677_));
 sg13g2_nor2b_1 _3252_ (.A(_1677_),
    .B_N(_1674_),
    .Y(_1678_));
 sg13g2_xor2_1 _3253_ (.B(_1677_),
    .A(_1674_),
    .X(_1679_));
 sg13g2_and3_1 _3254_ (.X(_1680_),
    .A(params_ready_internal),
    .B(net1),
    .C(net10));
 sg13g2_nand3_1 _3255_ (.B(net1),
    .C(net10),
    .A(net131),
    .Y(_1681_));
 sg13g2_nor2_2 _3256_ (.A(_1062_),
    .B(net344),
    .Y(_1682_));
 sg13g2_nand2_1 _3257_ (.Y(_1683_),
    .A(net336),
    .B(net348));
 sg13g2_nor2_2 _3258_ (.A(net334),
    .B(net344),
    .Y(_1684_));
 sg13g2_xnor2_1 _3259_ (.Y(_1685_),
    .A(net140),
    .B(\system_inst.neuron.u[1] ));
 sg13g2_o21ai_1 _3260_ (.B1(net421),
    .Y(_1686_),
    .A1(\system_inst.neuron.u[1] ),
    .A2(net347));
 sg13g2_a221oi_1 _3261_ (.B2(_1685_),
    .C1(_1686_),
    .B1(_1684_),
    .A1(_1679_),
    .Y(_0028_),
    .A2(_1682_));
 sg13g2_and2_1 _3262_ (.A(\system_inst.neuron.u[1] ),
    .B(_1676_),
    .X(_1687_));
 sg13g2_xnor2_1 _3263_ (.Y(_1688_),
    .A(_1634_),
    .B(_1636_));
 sg13g2_nand2b_1 _3264_ (.Y(_1689_),
    .B(_1688_),
    .A_N(_1671_));
 sg13g2_xor2_1 _3265_ (.B(_1689_),
    .A(\system_inst.neuron.u[2] ),
    .X(_1690_));
 sg13g2_o21ai_1 _3266_ (.B1(_1690_),
    .Y(_1691_),
    .A1(_1678_),
    .A2(_1687_));
 sg13g2_nor3_1 _3267_ (.A(_1678_),
    .B(_1687_),
    .C(_1690_),
    .Y(_1692_));
 sg13g2_nor2_1 _3268_ (.A(_1062_),
    .B(_1692_),
    .Y(_1693_));
 sg13g2_nand2_1 _3269_ (.Y(_1694_),
    .A(\system_inst.internal_param_d[1] ),
    .B(\system_inst.neuron.u[2] ));
 sg13g2_xor2_1 _3270_ (.B(\system_inst.neuron.u[2] ),
    .A(\system_inst.internal_param_d[1] ),
    .X(_1695_));
 sg13g2_a21oi_1 _3271_ (.A1(net140),
    .A2(\system_inst.neuron.u[1] ),
    .Y(_1696_),
    .B1(_1695_));
 sg13g2_nand3_1 _3272_ (.B(\system_inst.neuron.u[1] ),
    .C(_1695_),
    .A(net140),
    .Y(_1697_));
 sg13g2_nor2_1 _3273_ (.A(net334),
    .B(_1696_),
    .Y(_1698_));
 sg13g2_a221oi_1 _3274_ (.B2(_1698_),
    .C1(net344),
    .B1(_1697_),
    .A1(_1691_),
    .Y(_1699_),
    .A2(_1693_));
 sg13g2_o21ai_1 _3275_ (.B1(net421),
    .Y(_1700_),
    .A1(net153),
    .A2(net347));
 sg13g2_nor2_1 _3276_ (.A(_1699_),
    .B(_1700_),
    .Y(_0029_));
 sg13g2_nand2b_1 _3277_ (.Y(_1701_),
    .B(_1689_),
    .A_N(_0014_));
 sg13g2_xnor2_1 _3278_ (.Y(_1702_),
    .A(_1637_),
    .B(_1639_));
 sg13g2_or2_1 _3279_ (.X(_1703_),
    .B(_1702_),
    .A(_1671_));
 sg13g2_and2_1 _3280_ (.A(\system_inst.neuron.u[3] ),
    .B(_1703_),
    .X(_1704_));
 sg13g2_xor2_1 _3281_ (.B(_1703_),
    .A(\system_inst.neuron.u[3] ),
    .X(_1705_));
 sg13g2_inv_1 _3282_ (.Y(_1706_),
    .A(_1705_));
 sg13g2_a21oi_2 _3283_ (.B1(_1706_),
    .Y(_1707_),
    .A2(_1701_),
    .A1(_1691_));
 sg13g2_nand3_1 _3284_ (.B(_1701_),
    .C(_1706_),
    .A(_1691_),
    .Y(_1708_));
 sg13g2_nor2b_1 _3285_ (.A(_1707_),
    .B_N(_1708_),
    .Y(_1709_));
 sg13g2_nand2_1 _3286_ (.Y(_1710_),
    .A(\system_inst.internal_param_d[2] ),
    .B(\system_inst.neuron.u[3] ));
 sg13g2_xnor2_1 _3287_ (.Y(_1711_),
    .A(\system_inst.internal_param_d[2] ),
    .B(\system_inst.neuron.u[3] ));
 sg13g2_nand2_1 _3288_ (.Y(_1712_),
    .A(_1694_),
    .B(_1697_));
 sg13g2_inv_1 _3289_ (.Y(_1713_),
    .A(_1712_));
 sg13g2_nand2b_1 _3290_ (.Y(_1714_),
    .B(_1712_),
    .A_N(_1711_));
 sg13g2_a21oi_1 _3291_ (.A1(_1711_),
    .A2(_1713_),
    .Y(_1715_),
    .B1(net334));
 sg13g2_a221oi_1 _3292_ (.B2(_1715_),
    .C1(net344),
    .B1(_1714_),
    .A1(net334),
    .Y(_1716_),
    .A2(_1709_));
 sg13g2_o21ai_1 _3293_ (.B1(net424),
    .Y(_1717_),
    .A1(net157),
    .A2(net347));
 sg13g2_nor2_1 _3294_ (.A(_1716_),
    .B(_1717_),
    .Y(_0030_));
 sg13g2_xor2_1 _3295_ (.B(_1642_),
    .A(_1640_),
    .X(_1718_));
 sg13g2_or2_1 _3296_ (.X(_1719_),
    .B(_1718_),
    .A(_1671_));
 sg13g2_xnor2_1 _3297_ (.Y(_1720_),
    .A(_0964_),
    .B(_1719_));
 sg13g2_o21ai_1 _3298_ (.B1(_1720_),
    .Y(_1721_),
    .A1(_1704_),
    .A2(_1707_));
 sg13g2_nor3_1 _3299_ (.A(_1704_),
    .B(_1707_),
    .C(_1720_),
    .Y(_1722_));
 sg13g2_nor2_1 _3300_ (.A(_1062_),
    .B(_1722_),
    .Y(_1723_));
 sg13g2_xnor2_1 _3301_ (.Y(_1724_),
    .A(\system_inst.internal_param_d[3] ),
    .B(\system_inst.neuron.u[4] ));
 sg13g2_nand2_1 _3302_ (.Y(_1725_),
    .A(_1710_),
    .B(_1714_));
 sg13g2_inv_1 _3303_ (.Y(_1726_),
    .A(_1725_));
 sg13g2_nand2b_1 _3304_ (.Y(_1727_),
    .B(_1725_),
    .A_N(_1724_));
 sg13g2_a21oi_1 _3305_ (.A1(_1724_),
    .A2(_1726_),
    .Y(_1728_),
    .B1(net335));
 sg13g2_a221oi_1 _3306_ (.B2(_1728_),
    .C1(net345),
    .B1(_1727_),
    .A1(_1721_),
    .Y(_1729_),
    .A2(_1723_));
 sg13g2_o21ai_1 _3307_ (.B1(net422),
    .Y(_1730_),
    .A1(net150),
    .A2(net347));
 sg13g2_nor2_1 _3308_ (.A(_1729_),
    .B(_1730_),
    .Y(_0031_));
 sg13g2_nand2b_1 _3309_ (.Y(_1731_),
    .B(_1719_),
    .A_N(_0015_));
 sg13g2_and2_1 _3310_ (.A(_1721_),
    .B(_1731_),
    .X(_1732_));
 sg13g2_xnor2_1 _3311_ (.Y(_1733_),
    .A(_1643_),
    .B(_1645_));
 sg13g2_or2_1 _3312_ (.X(_1734_),
    .B(_1733_),
    .A(_1671_));
 sg13g2_nor2_1 _3313_ (.A(net416),
    .B(_1734_),
    .Y(_1735_));
 sg13g2_nand2_1 _3314_ (.Y(_1736_),
    .A(net416),
    .B(_1734_));
 sg13g2_nor2b_1 _3315_ (.A(_1735_),
    .B_N(_1736_),
    .Y(_1737_));
 sg13g2_xnor2_1 _3316_ (.Y(_1738_),
    .A(_1732_),
    .B(_1737_));
 sg13g2_xnor2_1 _3317_ (.Y(_1739_),
    .A(\system_inst.internal_param_d[4] ),
    .B(net416));
 sg13g2_o21ai_1 _3318_ (.B1(_1727_),
    .Y(_1740_),
    .A1(_0856_),
    .A2(_0964_));
 sg13g2_inv_1 _3319_ (.Y(_1741_),
    .A(_1740_));
 sg13g2_nand2b_1 _3320_ (.Y(_1742_),
    .B(_1740_),
    .A_N(_1739_));
 sg13g2_inv_1 _3321_ (.Y(_1743_),
    .A(_1742_));
 sg13g2_a21oi_1 _3322_ (.A1(_1739_),
    .A2(_1741_),
    .Y(_1744_),
    .B1(net334));
 sg13g2_a221oi_1 _3323_ (.B2(_1744_),
    .C1(net345),
    .B1(_1742_),
    .A1(net334),
    .Y(_1745_),
    .A2(_1738_));
 sg13g2_o21ai_1 _3324_ (.B1(net423),
    .Y(_1746_),
    .A1(net416),
    .A2(net347));
 sg13g2_nor2_1 _3325_ (.A(_1745_),
    .B(_1746_),
    .Y(_0032_));
 sg13g2_o21ai_1 _3326_ (.B1(_1736_),
    .Y(_1747_),
    .A1(_1732_),
    .A2(_1735_));
 sg13g2_xnor2_1 _3327_ (.Y(_1748_),
    .A(_1646_),
    .B(_1647_));
 sg13g2_nand2b_2 _3328_ (.Y(_1749_),
    .B(_1748_),
    .A_N(_1671_));
 sg13g2_xor2_1 _3329_ (.B(_1749_),
    .A(\system_inst.neuron.u[6] ),
    .X(_1750_));
 sg13g2_and2_1 _3330_ (.A(_1747_),
    .B(_1750_),
    .X(_1751_));
 sg13g2_o21ai_1 _3331_ (.B1(net335),
    .Y(_1752_),
    .A1(_1747_),
    .A2(_1750_));
 sg13g2_nor2_1 _3332_ (.A(_1751_),
    .B(_1752_),
    .Y(_1753_));
 sg13g2_a21oi_1 _3333_ (.A1(\system_inst.internal_param_d[4] ),
    .A2(\system_inst.neuron.u[5] ),
    .Y(_1754_),
    .B1(_1743_));
 sg13g2_nor2_1 _3334_ (.A(\system_inst.internal_param_d[5] ),
    .B(\system_inst.neuron.u[6] ),
    .Y(_1755_));
 sg13g2_nand2_1 _3335_ (.Y(_1756_),
    .A(\system_inst.internal_param_d[5] ),
    .B(\system_inst.neuron.u[6] ));
 sg13g2_nor2b_1 _3336_ (.A(_1755_),
    .B_N(_1756_),
    .Y(_1757_));
 sg13g2_xnor2_1 _3337_ (.Y(_1758_),
    .A(_1754_),
    .B(_1757_));
 sg13g2_a21oi_1 _3338_ (.A1(_1062_),
    .A2(_1758_),
    .Y(_1759_),
    .B1(_1753_));
 sg13g2_o21ai_1 _3339_ (.B1(net423),
    .Y(_1760_),
    .A1(net158),
    .A2(net347));
 sg13g2_a21oi_1 _3340_ (.A1(net347),
    .A2(_1759_),
    .Y(_0033_),
    .B1(_1760_));
 sg13g2_a21oi_2 _3341_ (.B1(_1751_),
    .Y(_1761_),
    .A2(_1749_),
    .A1(_1014_));
 sg13g2_o21ai_1 _3342_ (.B1(_1756_),
    .Y(_1762_),
    .A1(_1754_),
    .A2(_1755_));
 sg13g2_nor2_1 _3343_ (.A(net335),
    .B(_1762_),
    .Y(_1763_));
 sg13g2_a21oi_1 _3344_ (.A1(net335),
    .A2(_1761_),
    .Y(_1764_),
    .B1(_1763_));
 sg13g2_or2_1 _3345_ (.X(_1765_),
    .B(_1764_),
    .A(net143));
 sg13g2_a21oi_1 _3346_ (.A1(net143),
    .A2(_1764_),
    .Y(_1766_),
    .B1(net345));
 sg13g2_a221oi_1 _3347_ (.B2(_1766_),
    .C1(net420),
    .B1(_1765_),
    .A1(_0954_),
    .Y(_0034_),
    .A2(net345));
 sg13g2_o21ai_1 _3348_ (.B1(_0008_),
    .Y(_1767_),
    .A1(net143),
    .A2(_1761_));
 sg13g2_nor3_1 _3349_ (.A(_0010_),
    .B(_0008_),
    .C(_1761_),
    .Y(_1768_));
 sg13g2_nor2_1 _3350_ (.A(_1062_),
    .B(_1768_),
    .Y(_1769_));
 sg13g2_a21o_1 _3351_ (.A2(_1762_),
    .A1(\system_inst.neuron.u[7] ),
    .B1(\system_inst.neuron.u[8] ),
    .X(_1770_));
 sg13g2_nand3_1 _3352_ (.B(\system_inst.neuron.u[7] ),
    .C(_1762_),
    .A(\system_inst.neuron.u[8] ),
    .Y(_1771_));
 sg13g2_and2_1 _3353_ (.A(_1062_),
    .B(_1771_),
    .X(_1772_));
 sg13g2_a221oi_1 _3354_ (.B2(_1772_),
    .C1(net345),
    .B1(_1770_),
    .A1(_1767_),
    .Y(_1773_),
    .A2(_1769_));
 sg13g2_o21ai_1 _3355_ (.B1(net422),
    .Y(_1774_),
    .A1(net147),
    .A2(net347));
 sg13g2_nor2_1 _3356_ (.A(_1773_),
    .B(_1774_),
    .Y(_0035_));
 sg13g2_nor2_2 _3357_ (.A(_1769_),
    .B(_1772_),
    .Y(_1775_));
 sg13g2_or2_1 _3358_ (.X(_1776_),
    .B(_1775_),
    .A(net91));
 sg13g2_a21oi_1 _3359_ (.A1(net91),
    .A2(_1775_),
    .Y(_1777_),
    .B1(net346));
 sg13g2_a221oi_1 _3360_ (.B2(_1777_),
    .C1(net419),
    .B1(_1776_),
    .A1(_0944_),
    .Y(_0036_),
    .A2(net346));
 sg13g2_a21oi_1 _3361_ (.A1(_1673_),
    .A2(_1682_),
    .Y(_1778_),
    .B1(net154));
 sg13g2_a21oi_1 _3362_ (.A1(_1674_),
    .A2(_1682_),
    .Y(_1779_),
    .B1(_1778_));
 sg13g2_and2_1 _3363_ (.A(net421),
    .B(_1779_),
    .X(_0037_));
 sg13g2_o21ai_1 _3364_ (.B1(_1046_),
    .Y(_1780_),
    .A1(net11),
    .A2(_0983_));
 sg13g2_nand2_1 _3365_ (.Y(_1781_),
    .A(_1048_),
    .B(_1780_));
 sg13g2_nand2_1 _3366_ (.Y(_1782_),
    .A(net1),
    .B(_1781_));
 sg13g2_a22oi_1 _3367_ (.Y(_1783_),
    .B1(_1053_),
    .B2(_1036_),
    .A2(_1046_),
    .A1(_0983_));
 sg13g2_nand3_1 _3368_ (.B(_1781_),
    .C(_1783_),
    .A(net1),
    .Y(_1784_));
 sg13g2_a21oi_1 _3369_ (.A1(net131),
    .A2(_1784_),
    .Y(_1785_),
    .B1(net419));
 sg13g2_o21ai_1 _3370_ (.B1(_1785_),
    .Y(_0038_),
    .A1(_1047_),
    .A2(_1784_));
 sg13g2_a21oi_1 _3371_ (.A1(net12),
    .A2(net337),
    .Y(_1786_),
    .B1(net417));
 sg13g2_o21ai_1 _3372_ (.B1(_1786_),
    .Y(_0039_),
    .A1(_0933_),
    .A2(net337));
 sg13g2_o21ai_1 _3373_ (.B1(net422),
    .Y(_1787_),
    .A1(net410),
    .A2(net338));
 sg13g2_a21oi_1 _3374_ (.A1(_0845_),
    .A2(net338),
    .Y(_0040_),
    .B1(_1787_));
 sg13g2_a21oi_1 _3375_ (.A1(net127),
    .A2(net338),
    .Y(_1788_),
    .B1(net420));
 sg13g2_o21ai_1 _3376_ (.B1(_1788_),
    .Y(_0041_),
    .A1(_0911_),
    .A2(net337));
 sg13g2_a21oi_1 _3377_ (.A1(net137),
    .A2(net337),
    .Y(_1789_),
    .B1(net417));
 sg13g2_o21ai_1 _3378_ (.B1(_1789_),
    .Y(_0042_),
    .A1(_0900_),
    .A2(net337));
 sg13g2_o21ai_1 _3379_ (.B1(net422),
    .Y(_1790_),
    .A1(net407),
    .A2(net338));
 sg13g2_a21oi_1 _3380_ (.A1(_0823_),
    .A2(net337),
    .Y(_0043_),
    .B1(_1790_));
 sg13g2_o21ai_1 _3381_ (.B1(net422),
    .Y(_1791_),
    .A1(net121),
    .A2(net337));
 sg13g2_a21oi_1 _3382_ (.A1(_0812_),
    .A2(net337),
    .Y(_0044_),
    .B1(_1791_));
 sg13g2_o21ai_1 _3383_ (.B1(net421),
    .Y(_1792_),
    .A1(_0867_),
    .A2(_1041_));
 sg13g2_a21o_1 _3384_ (.A2(_1041_),
    .A1(net405),
    .B1(_1792_),
    .X(_0045_));
 sg13g2_o21ai_1 _3385_ (.B1(net421),
    .Y(_1793_),
    .A1(net404),
    .A2(net341));
 sg13g2_a21oi_1 _3386_ (.A1(_0845_),
    .A2(net341),
    .Y(_0046_),
    .B1(_1793_));
 sg13g2_o21ai_1 _3387_ (.B1(net421),
    .Y(_1794_),
    .A1(_0834_),
    .A2(_1041_));
 sg13g2_a21o_1 _3388_ (.A2(_1041_),
    .A1(net401),
    .B1(_1794_),
    .X(_0047_));
 sg13g2_a21oi_1 _3389_ (.A1(net137),
    .A2(net341),
    .Y(_1795_),
    .B1(net417));
 sg13g2_o21ai_1 _3390_ (.B1(_1795_),
    .Y(_0048_),
    .A1(_0889_),
    .A2(net341));
 sg13g2_o21ai_1 _3391_ (.B1(net422),
    .Y(_1796_),
    .A1(net134),
    .A2(net341));
 sg13g2_a21oi_1 _3392_ (.A1(_0823_),
    .A2(net341),
    .Y(_0049_),
    .B1(_1796_));
 sg13g2_o21ai_1 _3393_ (.B1(net422),
    .Y(_1797_),
    .A1(net396),
    .A2(net341));
 sg13g2_a21oi_1 _3394_ (.A1(_0812_),
    .A2(net341),
    .Y(_0050_),
    .B1(_1797_));
 sg13g2_a21oi_1 _3395_ (.A1(net96),
    .A2(_1044_),
    .Y(_1798_),
    .B1(net418));
 sg13g2_o21ai_1 _3396_ (.B1(_1798_),
    .Y(_0051_),
    .A1(_0867_),
    .A2(_1044_));
 sg13g2_a21oi_1 _3397_ (.A1(net98),
    .A2(_1044_),
    .Y(_1799_),
    .B1(net420));
 sg13g2_o21ai_1 _3398_ (.B1(_1799_),
    .Y(_0052_),
    .A1(_0845_),
    .A2(_1044_));
 sg13g2_a21oi_1 _3399_ (.A1(net113),
    .A2(_1044_),
    .Y(_0083_),
    .B1(net418));
 sg13g2_o21ai_1 _3400_ (.B1(_0083_),
    .Y(_0053_),
    .A1(_0834_),
    .A2(_1044_));
 sg13g2_a21oi_1 _3401_ (.A1(\system_inst.loader.shift_reg[2] ),
    .A2(_1043_),
    .Y(_0084_),
    .B1(net420));
 sg13g2_o21ai_1 _3402_ (.B1(_0084_),
    .Y(_0054_),
    .A1(_0878_),
    .A2(_1043_));
 sg13g2_a21oi_1 _3403_ (.A1(net118),
    .A2(_1044_),
    .Y(_0085_),
    .B1(net419));
 sg13g2_o21ai_1 _3404_ (.B1(_0085_),
    .Y(_0055_),
    .A1(_0823_),
    .A2(_1044_));
 sg13g2_o21ai_1 _3405_ (.B1(net425),
    .Y(_0086_),
    .A1(net115),
    .A2(_1043_));
 sg13g2_a21oi_1 _3406_ (.A1(_0812_),
    .A2(_1043_),
    .Y(_0056_),
    .B1(_0086_));
 sg13g2_o21ai_1 _3407_ (.B1(net421),
    .Y(_0087_),
    .A1(net140),
    .A2(net339));
 sg13g2_a21oi_1 _3408_ (.A1(_0867_),
    .A2(net339),
    .Y(_0057_),
    .B1(_0087_));
 sg13g2_o21ai_1 _3409_ (.B1(net421),
    .Y(_0088_),
    .A1(net135),
    .A2(net339));
 sg13g2_a21oi_1 _3410_ (.A1(_0845_),
    .A2(net339),
    .Y(_0058_),
    .B1(_0088_));
 sg13g2_o21ai_1 _3411_ (.B1(net424),
    .Y(_0089_),
    .A1(net124),
    .A2(net339));
 sg13g2_a21oi_1 _3412_ (.A1(_0834_),
    .A2(net339),
    .Y(_0059_),
    .B1(_0089_));
 sg13g2_a21oi_1 _3413_ (.A1(\system_inst.loader.shift_reg[2] ),
    .A2(net340),
    .Y(_0090_),
    .B1(net420));
 sg13g2_o21ai_1 _3414_ (.B1(_0090_),
    .Y(_0060_),
    .A1(_0856_),
    .A2(net340));
 sg13g2_o21ai_1 _3415_ (.B1(net423),
    .Y(_0091_),
    .A1(net126),
    .A2(net339));
 sg13g2_a21oi_1 _3416_ (.A1(_0823_),
    .A2(net339),
    .Y(_0061_),
    .B1(_0091_));
 sg13g2_o21ai_1 _3417_ (.B1(net423),
    .Y(_0092_),
    .A1(net112),
    .A2(net340));
 sg13g2_a21oi_1 _3418_ (.A1(_0812_),
    .A2(net340),
    .Y(_0062_),
    .B1(_0092_));
 sg13g2_nor3_1 _3419_ (.A(\system_inst.loader.state[5] ),
    .B(\system_inst.loader.state[2] ),
    .C(\system_inst.loader.state[3] ),
    .Y(_0093_));
 sg13g2_nand3_1 _3420_ (.B(_1046_),
    .C(_0093_),
    .A(_0019_),
    .Y(_0094_));
 sg13g2_o21ai_1 _3421_ (.B1(_0094_),
    .Y(_0095_),
    .A1(net11),
    .A2(_0093_));
 sg13g2_or2_1 _3422_ (.X(_0096_),
    .B(_0095_),
    .A(_1782_));
 sg13g2_inv_1 _3423_ (.Y(_0097_),
    .A(net330));
 sg13g2_a21o_2 _3424_ (.A2(_1046_),
    .A1(_1036_),
    .B1(\system_inst.loader.state[1] ),
    .X(_0098_));
 sg13g2_a21oi_1 _3425_ (.A1(net12),
    .A2(_0098_),
    .Y(_0099_),
    .B1(net330));
 sg13g2_o21ai_1 _3426_ (.B1(net425),
    .Y(_0100_),
    .A1(net104),
    .A2(_0097_));
 sg13g2_nor2_1 _3427_ (.A(_0099_),
    .B(_0100_),
    .Y(_0063_));
 sg13g2_a21oi_1 _3428_ (.A1(net104),
    .A2(_0098_),
    .Y(_0101_),
    .B1(net330));
 sg13g2_o21ai_1 _3429_ (.B1(net422),
    .Y(_0102_),
    .A1(\system_inst.loader.shift_reg[1] ),
    .A2(_0097_));
 sg13g2_nor2_1 _3430_ (.A(_0101_),
    .B(_0102_),
    .Y(_0064_));
 sg13g2_a21oi_1 _3431_ (.A1(net127),
    .A2(_0098_),
    .Y(_0103_),
    .B1(net330));
 sg13g2_o21ai_1 _3432_ (.B1(net425),
    .Y(_0104_),
    .A1(\system_inst.loader.shift_reg[2] ),
    .A2(_0097_));
 sg13g2_nor2_1 _3433_ (.A(_0103_),
    .B(_0104_),
    .Y(_0065_));
 sg13g2_a21oi_1 _3434_ (.A1(net137),
    .A2(_0098_),
    .Y(_0105_),
    .B1(net330));
 sg13g2_o21ai_1 _3435_ (.B1(net425),
    .Y(_0106_),
    .A1(net120),
    .A2(_0097_));
 sg13g2_nor2_1 _3436_ (.A(_0105_),
    .B(_0106_),
    .Y(_0066_));
 sg13g2_a21oi_1 _3437_ (.A1(net120),
    .A2(_0098_),
    .Y(_0107_),
    .B1(net330));
 sg13g2_o21ai_1 _3438_ (.B1(net425),
    .Y(_0108_),
    .A1(net109),
    .A2(_0097_));
 sg13g2_nor2_1 _3439_ (.A(_0107_),
    .B(_0108_),
    .Y(_0067_));
 sg13g2_o21ai_1 _3440_ (.B1(_0801_),
    .Y(_0109_),
    .A1(_1783_),
    .A2(_0096_));
 sg13g2_nor2_1 _3441_ (.A(_0801_),
    .B(net330),
    .Y(_0110_));
 sg13g2_nand2_1 _3442_ (.Y(_0111_),
    .A(net425),
    .B(net139));
 sg13g2_nor2_1 _3443_ (.A(_0110_),
    .B(_0111_),
    .Y(_0068_));
 sg13g2_nand2_1 _3444_ (.Y(_0112_),
    .A(net122),
    .B(_0110_));
 sg13g2_o21ai_1 _3445_ (.B1(_0112_),
    .Y(_0113_),
    .A1(net330),
    .A2(_0098_));
 sg13g2_o21ai_1 _3446_ (.B1(net425),
    .Y(_0114_),
    .A1(net122),
    .A2(_0110_));
 sg13g2_nor2_1 _3447_ (.A(_0113_),
    .B(net123),
    .Y(_0069_));
 sg13g2_nand2_1 _3448_ (.Y(_0115_),
    .A(_0790_),
    .B(_0098_));
 sg13g2_a221oi_1 _3449_ (.B2(_0115_),
    .C1(net419),
    .B1(_0113_),
    .A1(_0790_),
    .Y(_0070_),
    .A2(_0112_));
 sg13g2_nor3_1 _3450_ (.A(net418),
    .B(net336),
    .C(net346),
    .Y(_0071_));
 sg13g2_nand2_2 _3451_ (.Y(_0116_),
    .A(net357),
    .B(net373));
 sg13g2_nor2b_1 _3452_ (.A(net377),
    .B_N(net350),
    .Y(_0117_));
 sg13g2_nor2b_1 _3453_ (.A(_0116_),
    .B_N(_0117_),
    .Y(_0118_));
 sg13g2_nand2_2 _3454_ (.Y(_0119_),
    .A(net361),
    .B(net370));
 sg13g2_inv_1 _3455_ (.Y(_0120_),
    .A(_0119_));
 sg13g2_xnor2_1 _3456_ (.Y(_0121_),
    .A(_0116_),
    .B(_0117_));
 sg13g2_a21oi_2 _3457_ (.B1(_0118_),
    .Y(_0122_),
    .A2(_0121_),
    .A1(_0120_));
 sg13g2_nand2b_1 _3458_ (.Y(_0123_),
    .B(net352),
    .A_N(net374));
 sg13g2_nand2_2 _3459_ (.Y(_0124_),
    .A(net356),
    .B(net369));
 sg13g2_xor2_1 _3460_ (.B(_0124_),
    .A(_0123_),
    .X(_0125_));
 sg13g2_nand2b_1 _3461_ (.Y(_0126_),
    .B(_0125_),
    .A_N(_1065_));
 sg13g2_xnor2_1 _3462_ (.Y(_0127_),
    .A(_1065_),
    .B(_0125_));
 sg13g2_nor2b_1 _3463_ (.A(_0122_),
    .B_N(_0127_),
    .Y(_0128_));
 sg13g2_nand2_2 _3464_ (.Y(_0129_),
    .A(net351),
    .B(net373));
 sg13g2_and2_2 _3465_ (.A(net365),
    .B(net369),
    .X(_0130_));
 sg13g2_nand2_2 _3466_ (.Y(_0131_),
    .A(net365),
    .B(net369));
 sg13g2_xor2_1 _3467_ (.B(_0124_),
    .A(_1065_),
    .X(_0132_));
 sg13g2_nand2b_1 _3468_ (.Y(_0133_),
    .B(_0132_),
    .A_N(_0129_));
 sg13g2_xnor2_1 _3469_ (.Y(_0134_),
    .A(_0129_),
    .B(_0132_));
 sg13g2_nand2b_1 _3470_ (.Y(_0135_),
    .B(_0122_),
    .A_N(_0127_));
 sg13g2_a21oi_1 _3471_ (.A1(_0134_),
    .A2(_0135_),
    .Y(_0136_),
    .B1(_0128_));
 sg13g2_nor2_2 _3472_ (.A(_0713_),
    .B(_0724_),
    .Y(_0137_));
 sg13g2_nand2_1 _3473_ (.Y(_0138_),
    .A(_0130_),
    .B(_0137_));
 sg13g2_a22oi_1 _3474_ (.Y(_0139_),
    .B1(net369),
    .B2(net351),
    .A2(net365),
    .A1(net357));
 sg13g2_a21oi_1 _3475_ (.A1(_0130_),
    .A2(_0137_),
    .Y(_0140_),
    .B1(_0139_));
 sg13g2_xnor2_1 _3476_ (.Y(_0141_),
    .A(_0129_),
    .B(_0140_));
 sg13g2_o21ai_1 _3477_ (.B1(_0126_),
    .Y(_0142_),
    .A1(_0123_),
    .A2(_0124_));
 sg13g2_nor2_1 _3478_ (.A(_0713_),
    .B(net370),
    .Y(_0143_));
 sg13g2_nor3_1 _3479_ (.A(net349),
    .B(net370),
    .C(_1061_),
    .Y(_0144_));
 sg13g2_xnor2_1 _3480_ (.Y(_0145_),
    .A(_1061_),
    .B(_0143_));
 sg13g2_xnor2_1 _3481_ (.Y(_0146_),
    .A(net360),
    .B(_0145_));
 sg13g2_nor2b_1 _3482_ (.A(_0146_),
    .B_N(_0142_),
    .Y(_0147_));
 sg13g2_xor2_1 _3483_ (.B(_0146_),
    .A(_0142_),
    .X(_0148_));
 sg13g2_inv_1 _3484_ (.Y(_0149_),
    .A(_0148_));
 sg13g2_xor2_1 _3485_ (.B(_0148_),
    .A(_0141_),
    .X(_0150_));
 sg13g2_nor2_1 _3486_ (.A(net349),
    .B(_1172_),
    .Y(_0151_));
 sg13g2_o21ai_1 _3487_ (.B1(_0151_),
    .Y(_0152_),
    .A1(net386),
    .A2(net394));
 sg13g2_nor2_1 _3488_ (.A(net349),
    .B(_0768_),
    .Y(_0153_));
 sg13g2_nand2_1 _3489_ (.Y(_0154_),
    .A(net350),
    .B(_1172_));
 sg13g2_o21ai_1 _3490_ (.B1(_0154_),
    .Y(_0155_),
    .A1(_0768_),
    .A2(_0152_));
 sg13g2_mux2_1 _3491_ (.A0(_0768_),
    .A1(_0153_),
    .S(_0152_),
    .X(_0156_));
 sg13g2_o21ai_1 _3492_ (.B1(_0133_),
    .Y(_0157_),
    .A1(_1064_),
    .A2(_0131_));
 sg13g2_and2_1 _3493_ (.A(net331),
    .B(_0157_),
    .X(_0158_));
 sg13g2_xor2_1 _3494_ (.B(_0157_),
    .A(net331),
    .X(_0159_));
 sg13g2_xnor2_1 _3495_ (.Y(_0160_),
    .A(net333),
    .B(_0159_));
 sg13g2_xor2_1 _3496_ (.B(_0150_),
    .A(_0136_),
    .X(_0161_));
 sg13g2_nand2b_1 _3497_ (.Y(_0162_),
    .B(_0161_),
    .A_N(_0160_));
 sg13g2_o21ai_1 _3498_ (.B1(_0162_),
    .Y(_0163_),
    .A1(_0136_),
    .A2(_0150_));
 sg13g2_o21ai_1 _3499_ (.B1(_0138_),
    .Y(_0164_),
    .A1(_0129_),
    .A2(_0139_));
 sg13g2_and2_1 _3500_ (.A(net332),
    .B(_0164_),
    .X(_0165_));
 sg13g2_xor2_1 _3501_ (.B(_0164_),
    .A(net332),
    .X(_0166_));
 sg13g2_xnor2_1 _3502_ (.Y(_0167_),
    .A(_0155_),
    .B(_0166_));
 sg13g2_inv_1 _3503_ (.Y(_0168_),
    .A(_0167_));
 sg13g2_a21oi_1 _3504_ (.A1(_0141_),
    .A2(_0149_),
    .Y(_0169_),
    .B1(_0147_));
 sg13g2_nand3_1 _3505_ (.B(net365),
    .C(net369),
    .A(net351),
    .Y(_0170_));
 sg13g2_o21ai_1 _3506_ (.B1(net351),
    .Y(_0171_),
    .A1(net365),
    .A2(net369));
 sg13g2_inv_1 _3507_ (.Y(_0172_),
    .A(_0171_));
 sg13g2_nand2_1 _3508_ (.Y(_0173_),
    .A(_0170_),
    .B(_0172_));
 sg13g2_xor2_1 _3509_ (.B(_0173_),
    .A(_0129_),
    .X(_0174_));
 sg13g2_nor4_2 _3510_ (.A(net349),
    .B(_0735_),
    .C(net364),
    .Y(_0175_),
    .D(net370));
 sg13g2_a221oi_1 _3511_ (.B2(net360),
    .C1(_0144_),
    .B1(_0145_),
    .A1(net352),
    .Y(_0176_),
    .A2(_0746_));
 sg13g2_nor2_1 _3512_ (.A(_0175_),
    .B(_0176_),
    .Y(_0177_));
 sg13g2_xnor2_1 _3513_ (.Y(_0178_),
    .A(_0174_),
    .B(_0177_));
 sg13g2_nor2_1 _3514_ (.A(_0169_),
    .B(_0178_),
    .Y(_0179_));
 sg13g2_xor2_1 _3515_ (.B(_0178_),
    .A(_0169_),
    .X(_0180_));
 sg13g2_xnor2_1 _3516_ (.Y(_0181_),
    .A(_0167_),
    .B(_0180_));
 sg13g2_nand2_1 _3517_ (.Y(_0182_),
    .A(_0163_),
    .B(_0181_));
 sg13g2_nand2_1 _3518_ (.Y(_0183_),
    .A(net350),
    .B(net377));
 sg13g2_a21o_1 _3519_ (.A2(_0159_),
    .A1(net333),
    .B1(_0158_),
    .X(_0184_));
 sg13g2_nand2b_1 _3520_ (.Y(_0185_),
    .B(_0184_),
    .A_N(net342));
 sg13g2_xor2_1 _3521_ (.B(_0184_),
    .A(net342),
    .X(_0186_));
 sg13g2_xnor2_1 _3522_ (.Y(_0187_),
    .A(_0163_),
    .B(_0181_));
 sg13g2_o21ai_1 _3523_ (.B1(_0182_),
    .Y(_0188_),
    .A1(_0186_),
    .A2(_0187_));
 sg13g2_a21o_1 _3524_ (.A2(_0166_),
    .A1(_0155_),
    .B1(_0165_),
    .X(_0189_));
 sg13g2_nand2b_1 _3525_ (.Y(_0190_),
    .B(_0189_),
    .A_N(net343));
 sg13g2_xor2_1 _3526_ (.B(_0189_),
    .A(net343),
    .X(_0191_));
 sg13g2_inv_1 _3527_ (.Y(_0192_),
    .A(_0191_));
 sg13g2_a21oi_1 _3528_ (.A1(_0168_),
    .A2(_0180_),
    .Y(_0193_),
    .B1(_0179_));
 sg13g2_o21ai_1 _3529_ (.B1(_0170_),
    .Y(_0194_),
    .A1(_0129_),
    .A2(_0171_));
 sg13g2_nand2_1 _3530_ (.Y(_0195_),
    .A(net332),
    .B(_0194_));
 sg13g2_xor2_1 _3531_ (.B(_0194_),
    .A(net332),
    .X(_0196_));
 sg13g2_nand2_1 _3532_ (.Y(_0197_),
    .A(net333),
    .B(_0196_));
 sg13g2_xnor2_1 _3533_ (.Y(_0198_),
    .A(net333),
    .B(_0196_));
 sg13g2_inv_1 _3534_ (.Y(_0199_),
    .A(_0198_));
 sg13g2_a21oi_2 _3535_ (.B1(_0175_),
    .Y(_0200_),
    .A2(_0177_),
    .A1(_0174_));
 sg13g2_nand2_1 _3536_ (.Y(_0201_),
    .A(net354),
    .B(net361));
 sg13g2_xnor2_1 _3537_ (.Y(_0202_),
    .A(net354),
    .B(_0009_));
 sg13g2_nor2b_1 _3538_ (.A(_1064_),
    .B_N(_0202_),
    .Y(_0203_));
 sg13g2_xnor2_1 _3539_ (.Y(_0204_),
    .A(_1064_),
    .B(_0202_));
 sg13g2_xnor2_1 _3540_ (.Y(_0205_),
    .A(_0174_),
    .B(_0204_));
 sg13g2_xor2_1 _3541_ (.B(_0205_),
    .A(_0200_),
    .X(_0206_));
 sg13g2_nand2_1 _3542_ (.Y(_0207_),
    .A(_0199_),
    .B(_0206_));
 sg13g2_xnor2_1 _3543_ (.Y(_0208_),
    .A(_0198_),
    .B(_0206_));
 sg13g2_nor2b_1 _3544_ (.A(_0193_),
    .B_N(_0208_),
    .Y(_0209_));
 sg13g2_xnor2_1 _3545_ (.Y(_0210_),
    .A(_0193_),
    .B(_0208_));
 sg13g2_xnor2_1 _3546_ (.Y(_0211_),
    .A(_0191_),
    .B(_0210_));
 sg13g2_nand2_1 _3547_ (.Y(_0212_),
    .A(_0188_),
    .B(_0211_));
 sg13g2_xnor2_1 _3548_ (.Y(_0213_),
    .A(_0188_),
    .B(_0211_));
 sg13g2_o21ai_1 _3549_ (.B1(_0212_),
    .Y(_0214_),
    .A1(_0185_),
    .A2(_0213_));
 sg13g2_a21oi_1 _3550_ (.A1(_0192_),
    .A2(_0210_),
    .Y(_0215_),
    .B1(_0209_));
 sg13g2_nand2_1 _3551_ (.Y(_0216_),
    .A(_0195_),
    .B(_0197_));
 sg13g2_nand3_1 _3552_ (.B(_0195_),
    .C(_0197_),
    .A(net343),
    .Y(_0217_));
 sg13g2_xor2_1 _3553_ (.B(_0216_),
    .A(net343),
    .X(_0218_));
 sg13g2_o21ai_1 _3554_ (.B1(_0207_),
    .Y(_0219_),
    .A1(_0200_),
    .A2(_0205_));
 sg13g2_nand2_1 _3555_ (.Y(_0220_),
    .A(_0724_),
    .B(_1060_));
 sg13g2_o21ai_1 _3556_ (.B1(_0220_),
    .Y(_0221_),
    .A1(_0009_),
    .A2(_0201_));
 sg13g2_xor2_1 _3557_ (.B(_0221_),
    .A(_0174_),
    .X(_0222_));
 sg13g2_a21o_1 _3558_ (.A2(_0204_),
    .A1(_0174_),
    .B1(_0203_),
    .X(_0223_));
 sg13g2_nand2_1 _3559_ (.Y(_0224_),
    .A(_0222_),
    .B(_0223_));
 sg13g2_xnor2_1 _3560_ (.Y(_0225_),
    .A(_0222_),
    .B(_0223_));
 sg13g2_xnor2_1 _3561_ (.Y(_0226_),
    .A(_0199_),
    .B(_0225_));
 sg13g2_xor2_1 _3562_ (.B(_0226_),
    .A(_0219_),
    .X(_0227_));
 sg13g2_nor2b_1 _3563_ (.A(_0218_),
    .B_N(_0227_),
    .Y(_0228_));
 sg13g2_xnor2_1 _3564_ (.Y(_0229_),
    .A(_0218_),
    .B(_0227_));
 sg13g2_nand2b_1 _3565_ (.Y(_0230_),
    .B(_0229_),
    .A_N(_0215_));
 sg13g2_xnor2_1 _3566_ (.Y(_0231_),
    .A(_0215_),
    .B(_0229_));
 sg13g2_inv_1 _3567_ (.Y(_0232_),
    .A(_0231_));
 sg13g2_xnor2_1 _3568_ (.Y(_0233_),
    .A(_0190_),
    .B(_0231_));
 sg13g2_xnor2_1 _3569_ (.Y(_0234_),
    .A(_0119_),
    .B(_0121_));
 sg13g2_nand2_2 _3570_ (.Y(_0235_),
    .A(net357),
    .B(net377));
 sg13g2_nor3_1 _3571_ (.A(net349),
    .B(net381),
    .C(_0235_),
    .Y(_0236_));
 sg13g2_o21ai_1 _3572_ (.B1(_0235_),
    .Y(_0237_),
    .A1(net349),
    .A2(net381));
 sg13g2_and2_1 _3573_ (.A(net360),
    .B(net373),
    .X(_0238_));
 sg13g2_o21ai_1 _3574_ (.B1(_0237_),
    .Y(_0239_),
    .A1(_0236_),
    .A2(_0238_));
 sg13g2_nor2b_1 _3575_ (.A(_0239_),
    .B_N(_0234_),
    .Y(_0240_));
 sg13g2_xor2_1 _3576_ (.B(_0119_),
    .A(_0021_),
    .X(_0241_));
 sg13g2_nand2b_1 _3577_ (.Y(_0242_),
    .B(_0241_),
    .A_N(_0116_));
 sg13g2_xnor2_1 _3578_ (.Y(_0243_),
    .A(_0116_),
    .B(_0241_));
 sg13g2_xnor2_1 _3579_ (.Y(_0244_),
    .A(_0234_),
    .B(_0239_));
 sg13g2_a21oi_1 _3580_ (.A1(_0243_),
    .A2(_0244_),
    .Y(_0245_),
    .B1(_0240_));
 sg13g2_xnor2_1 _3581_ (.Y(_0246_),
    .A(net350),
    .B(_0122_));
 sg13g2_nand2b_1 _3582_ (.Y(_0247_),
    .B(_0246_),
    .A_N(_0245_));
 sg13g2_o21ai_1 _3583_ (.B1(_0242_),
    .Y(_0248_),
    .A1(_0735_),
    .A2(_0131_));
 sg13g2_and2_1 _3584_ (.A(net331),
    .B(_0248_),
    .X(_0249_));
 sg13g2_xor2_1 _3585_ (.B(_0248_),
    .A(net331),
    .X(_0250_));
 sg13g2_xnor2_1 _3586_ (.Y(_0251_),
    .A(net333),
    .B(_0250_));
 sg13g2_xnor2_1 _3587_ (.Y(_0252_),
    .A(_0245_),
    .B(_0246_));
 sg13g2_inv_1 _3588_ (.Y(_0253_),
    .A(_0252_));
 sg13g2_o21ai_1 _3589_ (.B1(_0247_),
    .Y(_0254_),
    .A1(_0251_),
    .A2(_0253_));
 sg13g2_xnor2_1 _3590_ (.Y(_0255_),
    .A(_0160_),
    .B(_0161_));
 sg13g2_nand2_1 _3591_ (.Y(_0256_),
    .A(_0254_),
    .B(_0255_));
 sg13g2_a21o_1 _3592_ (.A2(_0250_),
    .A1(net333),
    .B1(_0249_),
    .X(_0257_));
 sg13g2_nand2b_1 _3593_ (.Y(_0258_),
    .B(_0257_),
    .A_N(net342));
 sg13g2_xor2_1 _3594_ (.B(_0257_),
    .A(net342),
    .X(_0259_));
 sg13g2_xnor2_1 _3595_ (.Y(_0260_),
    .A(_0254_),
    .B(_0255_));
 sg13g2_o21ai_1 _3596_ (.B1(_0256_),
    .Y(_0261_),
    .A1(_0259_),
    .A2(_0260_));
 sg13g2_xor2_1 _3597_ (.B(_0187_),
    .A(_0186_),
    .X(_0262_));
 sg13g2_xnor2_1 _3598_ (.Y(_0263_),
    .A(_0261_),
    .B(_0262_));
 sg13g2_nor2_1 _3599_ (.A(_0258_),
    .B(_0263_),
    .Y(_0264_));
 sg13g2_a21oi_2 _3600_ (.B1(_0264_),
    .Y(_0265_),
    .A2(_0262_),
    .A1(_0261_));
 sg13g2_xor2_1 _3601_ (.B(_0213_),
    .A(_0185_),
    .X(_0266_));
 sg13g2_nand2b_1 _3602_ (.Y(_0267_),
    .B(_0266_),
    .A_N(_0265_));
 sg13g2_xnor2_1 _3603_ (.Y(_0268_),
    .A(_0265_),
    .B(_0266_));
 sg13g2_nor2b_1 _3604_ (.A(_0236_),
    .B_N(_0237_),
    .Y(_0269_));
 sg13g2_nand2b_1 _3605_ (.Y(_0270_),
    .B(net350),
    .A_N(net386));
 sg13g2_nand2_2 _3606_ (.Y(_0271_),
    .A(net357),
    .B(net381));
 sg13g2_or2_1 _3607_ (.X(_0272_),
    .B(_0271_),
    .A(_0270_));
 sg13g2_nand2_2 _3608_ (.Y(_0273_),
    .A(net360),
    .B(net377));
 sg13g2_xnor2_1 _3609_ (.Y(_0274_),
    .A(_0270_),
    .B(_0271_));
 sg13g2_o21ai_1 _3610_ (.B1(_0272_),
    .Y(_0275_),
    .A1(_0273_),
    .A2(_0274_));
 sg13g2_mux2_1 _3611_ (.A0(_0238_),
    .A1(_0275_),
    .S(_0269_),
    .X(_0276_));
 sg13g2_xor2_1 _3612_ (.B(_0244_),
    .A(_0243_),
    .X(_0277_));
 sg13g2_and2_1 _3613_ (.A(_0276_),
    .B(_0277_),
    .X(_0278_));
 sg13g2_and2_1 _3614_ (.A(_0130_),
    .B(net331),
    .X(_0279_));
 sg13g2_xnor2_1 _3615_ (.Y(_0280_),
    .A(_0131_),
    .B(net331));
 sg13g2_xor2_1 _3616_ (.B(_0280_),
    .A(net333),
    .X(_0281_));
 sg13g2_xor2_1 _3617_ (.B(_0277_),
    .A(_0276_),
    .X(_0282_));
 sg13g2_a21o_1 _3618_ (.A2(_0282_),
    .A1(_0281_),
    .B1(_0278_),
    .X(_0283_));
 sg13g2_xnor2_1 _3619_ (.Y(_0284_),
    .A(_0251_),
    .B(_0252_));
 sg13g2_and2_1 _3620_ (.A(_0283_),
    .B(_0284_),
    .X(_0285_));
 sg13g2_a21oi_1 _3621_ (.A1(net333),
    .A2(_0280_),
    .Y(_0286_),
    .B1(_0279_));
 sg13g2_nor2_1 _3622_ (.A(net342),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_xor2_1 _3623_ (.B(_0286_),
    .A(net342),
    .X(_0288_));
 sg13g2_xor2_1 _3624_ (.B(_0284_),
    .A(_0283_),
    .X(_0289_));
 sg13g2_a21o_1 _3625_ (.A2(_0289_),
    .A1(_0288_),
    .B1(_0285_),
    .X(_0290_));
 sg13g2_xor2_1 _3626_ (.B(_0260_),
    .A(_0259_),
    .X(_0291_));
 sg13g2_nand2_1 _3627_ (.Y(_0292_),
    .A(_0290_),
    .B(_0291_));
 sg13g2_xor2_1 _3628_ (.B(_0291_),
    .A(_0290_),
    .X(_0293_));
 sg13g2_nand2_1 _3629_ (.Y(_0294_),
    .A(_0287_),
    .B(_0293_));
 sg13g2_xnor2_1 _3630_ (.Y(_0295_),
    .A(_0258_),
    .B(_0263_));
 sg13g2_a21o_1 _3631_ (.A2(_0294_),
    .A1(_0292_),
    .B1(_0295_),
    .X(_0296_));
 sg13g2_nand3_1 _3632_ (.B(_0294_),
    .C(_0295_),
    .A(_0292_),
    .Y(_0297_));
 sg13g2_nand2_1 _3633_ (.Y(_0298_),
    .A(net357),
    .B(net386));
 sg13g2_nor2b_1 _3634_ (.A(net391),
    .B_N(net350),
    .Y(_0299_));
 sg13g2_nand2b_1 _3635_ (.Y(_0300_),
    .B(_0299_),
    .A_N(_0298_));
 sg13g2_nand2_2 _3636_ (.Y(_0301_),
    .A(net360),
    .B(net381));
 sg13g2_a21oi_1 _3637_ (.A1(net357),
    .A2(net385),
    .Y(_0302_),
    .B1(_0299_));
 sg13g2_xnor2_1 _3638_ (.Y(_0303_),
    .A(_0298_),
    .B(_0299_));
 sg13g2_o21ai_1 _3639_ (.B1(_0300_),
    .Y(_0304_),
    .A1(_0301_),
    .A2(_0302_));
 sg13g2_xor2_1 _3640_ (.B(_0274_),
    .A(_0273_),
    .X(_0305_));
 sg13g2_nand2_1 _3641_ (.Y(_0306_),
    .A(_0304_),
    .B(_0305_));
 sg13g2_xnor2_1 _3642_ (.Y(_0307_),
    .A(_0304_),
    .B(_0305_));
 sg13g2_o21ai_1 _3643_ (.B1(_0306_),
    .Y(_0308_),
    .A1(_0022_),
    .A2(_0307_));
 sg13g2_xor2_1 _3644_ (.B(_0275_),
    .A(_0269_),
    .X(_0309_));
 sg13g2_nand2_1 _3645_ (.Y(_0310_),
    .A(_0308_),
    .B(_0309_));
 sg13g2_xnor2_1 _3646_ (.Y(_0311_),
    .A(_0308_),
    .B(_0309_));
 sg13g2_o21ai_1 _3647_ (.B1(_0154_),
    .Y(_0312_),
    .A1(_0152_),
    .A2(_0271_));
 sg13g2_nand2_1 _3648_ (.Y(_0313_),
    .A(net365),
    .B(net373));
 sg13g2_and3_1 _3649_ (.X(_0314_),
    .A(net365),
    .B(net373),
    .C(net331));
 sg13g2_xnor2_1 _3650_ (.Y(_0315_),
    .A(net331),
    .B(_0313_));
 sg13g2_xnor2_1 _3651_ (.Y(_0316_),
    .A(_0312_),
    .B(_0315_));
 sg13g2_o21ai_1 _3652_ (.B1(_0310_),
    .Y(_0317_),
    .A1(_0311_),
    .A2(_0316_));
 sg13g2_xor2_1 _3653_ (.B(_0282_),
    .A(_0281_),
    .X(_0318_));
 sg13g2_nand2_1 _3654_ (.Y(_0319_),
    .A(_0317_),
    .B(_0318_));
 sg13g2_a21oi_1 _3655_ (.A1(_0312_),
    .A2(_0315_),
    .Y(_0320_),
    .B1(_0314_));
 sg13g2_nor2_1 _3656_ (.A(net342),
    .B(_0320_),
    .Y(_0321_));
 sg13g2_xnor2_1 _3657_ (.Y(_0322_),
    .A(net342),
    .B(_0320_));
 sg13g2_xnor2_1 _3658_ (.Y(_0323_),
    .A(_0317_),
    .B(_0318_));
 sg13g2_o21ai_1 _3659_ (.B1(_0319_),
    .Y(_0324_),
    .A1(_0322_),
    .A2(_0323_));
 sg13g2_xor2_1 _3660_ (.B(_0289_),
    .A(_0288_),
    .X(_0325_));
 sg13g2_and2_1 _3661_ (.A(_0324_),
    .B(_0325_),
    .X(_0326_));
 sg13g2_xor2_1 _3662_ (.B(_0325_),
    .A(_0324_),
    .X(_0327_));
 sg13g2_a21oi_1 _3663_ (.A1(_0321_),
    .A2(_0327_),
    .Y(_0328_),
    .B1(_0326_));
 sg13g2_xnor2_1 _3664_ (.Y(_0329_),
    .A(_0287_),
    .B(_0293_));
 sg13g2_or2_1 _3665_ (.X(_0330_),
    .B(_0329_),
    .A(_0328_));
 sg13g2_nand2_1 _3666_ (.Y(_0331_),
    .A(_1172_),
    .B(_0137_));
 sg13g2_a22oi_1 _3667_ (.Y(_0332_),
    .B1(net390),
    .B2(net350),
    .A2(net385),
    .A1(net357));
 sg13g2_a21oi_1 _3668_ (.A1(_1172_),
    .A2(_0137_),
    .Y(_0333_),
    .B1(_0332_));
 sg13g2_xnor2_1 _3669_ (.Y(_0334_),
    .A(_0301_),
    .B(_0333_));
 sg13g2_and2_2 _3670_ (.A(net375),
    .B(net379),
    .X(_0335_));
 sg13g2_nand2_1 _3671_ (.Y(_0336_),
    .A(net375),
    .B(net380));
 sg13g2_nand2_1 _3672_ (.Y(_0337_),
    .A(net367),
    .B(net377));
 sg13g2_nor2_2 _3673_ (.A(_0746_),
    .B(_0768_),
    .Y(_0338_));
 sg13g2_a22oi_1 _3674_ (.Y(_0339_),
    .B1(net381),
    .B2(net363),
    .A2(net377),
    .A1(net369));
 sg13g2_a21oi_1 _3675_ (.A1(_0130_),
    .A2(_0335_),
    .Y(_0340_),
    .B1(net373));
 sg13g2_nor2_1 _3676_ (.A(_0339_),
    .B(_0340_),
    .Y(_0341_));
 sg13g2_nand2_1 _3677_ (.Y(_0342_),
    .A(_0334_),
    .B(_0341_));
 sg13g2_and4_2 _3678_ (.A(net356),
    .B(\system_inst.neuron.v[7] ),
    .C(net385),
    .D(net390),
    .X(_0343_));
 sg13g2_a22oi_1 _3679_ (.Y(_0344_),
    .B1(net390),
    .B2(net356),
    .A2(net385),
    .A1(net359));
 sg13g2_nor2_2 _3680_ (.A(_0343_),
    .B(_0344_),
    .Y(_0345_));
 sg13g2_a21oi_1 _3681_ (.A1(_0338_),
    .A2(_0345_),
    .Y(_0346_),
    .B1(_0343_));
 sg13g2_xnor2_1 _3682_ (.Y(_0347_),
    .A(_0334_),
    .B(_0341_));
 sg13g2_o21ai_1 _3683_ (.B1(_0342_),
    .Y(_0348_),
    .A1(_0346_),
    .A2(_0347_));
 sg13g2_nand2b_1 _3684_ (.Y(_0349_),
    .B(_0348_),
    .A_N(_0273_));
 sg13g2_a21oi_1 _3685_ (.A1(_0130_),
    .A2(_0335_),
    .Y(_0350_),
    .B1(_0339_));
 sg13g2_dfrbp_1 _3686_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net65),
    .D(net142),
    .Q_N(_0013_),
    .Q(\system_inst.neuron.u[1] ));
 sg13g2_dfrbp_1 _3687_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net27),
    .D(_0029_),
    .Q_N(_0014_),
    .Q(\system_inst.neuron.u[2] ));
 sg13g2_dfrbp_1 _3688_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net25),
    .D(_0030_),
    .Q_N(_0012_),
    .Q(\system_inst.neuron.u[3] ));
 sg13g2_dfrbp_1 _3689_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net23),
    .D(_0031_),
    .Q_N(_0015_),
    .Q(\system_inst.neuron.u[4] ));
 sg13g2_dfrbp_1 _3690_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net82),
    .D(_0032_),
    .Q_N(_1833_),
    .Q(\system_inst.neuron.u[5] ));
 sg13g2_dfrbp_1 _3691_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net80),
    .D(_0033_),
    .Q_N(_0011_),
    .Q(\system_inst.neuron.u[6] ));
 sg13g2_dfrbp_1 _3692_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net78),
    .D(net144),
    .Q_N(_0010_),
    .Q(\system_inst.neuron.u[7] ));
 sg13g2_dfrbp_1 _3693_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net76),
    .D(net148),
    .Q_N(_0008_),
    .Q(\system_inst.neuron.u[8] ));
 sg13g2_dfrbp_1 _3694_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net74),
    .D(net92),
    .Q_N(_0020_),
    .Q(\system_inst.neuron.u[9] ));
 sg13g2_dfrbp_1 _3695_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net72),
    .D(_0037_),
    .Q_N(_1832_),
    .Q(\system_inst.neuron.u[0] ));
 sg13g2_dfrbp_1 _3696_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net64),
    .D(_0038_),
    .Q_N(_1831_),
    .Q(params_ready_internal));
 sg13g2_dfrbp_1 _3697_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net62),
    .D(_0039_),
    .Q_N(_1830_),
    .Q(\system_inst.internal_param_a[0] ));
 sg13g2_dfrbp_1 _3698_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net60),
    .D(_0040_),
    .Q_N(_0018_),
    .Q(\system_inst.internal_param_a[1] ));
 sg13g2_dfrbp_1 _3699_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net58),
    .D(_0041_),
    .Q_N(_0017_),
    .Q(\system_inst.internal_param_a[2] ));
 sg13g2_dfrbp_1 _3700_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net56),
    .D(_0042_),
    .Q_N(_1829_),
    .Q(\system_inst.internal_param_a[3] ));
 sg13g2_dfrbp_1 _3701_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net54),
    .D(_0043_),
    .Q_N(_1828_),
    .Q(\system_inst.internal_param_a[4] ));
 sg13g2_dfrbp_1 _3702_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net52),
    .D(_0044_),
    .Q_N(_0016_),
    .Q(\system_inst.internal_param_a[5] ));
 sg13g2_dfrbp_1 _3703_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net50),
    .D(_0045_),
    .Q_N(_1827_),
    .Q(\system_inst.internal_param_b[0] ));
 sg13g2_dfrbp_1 _3704_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net48),
    .D(_0046_),
    .Q_N(_1826_),
    .Q(\system_inst.internal_param_b[1] ));
 sg13g2_dfrbp_1 _3705_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net46),
    .D(net152),
    .Q_N(_1825_),
    .Q(\system_inst.internal_param_b[2] ));
 sg13g2_dfrbp_1 _3706_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net44),
    .D(_0048_),
    .Q_N(_1824_),
    .Q(\system_inst.internal_param_b[3] ));
 sg13g2_dfrbp_1 _3707_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net42),
    .D(_0049_),
    .Q_N(_1823_),
    .Q(\system_inst.internal_param_b[4] ));
 sg13g2_dfrbp_1 _3708_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net40),
    .D(net110),
    .Q_N(_1822_),
    .Q(\system_inst.internal_param_b[5] ));
 sg13g2_dfrbp_1 _3709_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net38),
    .D(_0051_),
    .Q_N(_1821_),
    .Q(\system_inst.internal_param_c[0] ));
 sg13g2_dfrbp_1 _3710_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net36),
    .D(_0052_),
    .Q_N(_1820_),
    .Q(\system_inst.internal_param_c[1] ));
 sg13g2_dfrbp_1 _3711_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net34),
    .D(net114),
    .Q_N(_1819_),
    .Q(\system_inst.internal_param_c[2] ));
 sg13g2_dfrbp_1 _3712_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net32),
    .D(net90),
    .Q_N(_1818_),
    .Q(\system_inst.internal_param_c[3] ));
 sg13g2_dfrbp_1 _3713_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net30),
    .D(net119),
    .Q_N(_0007_),
    .Q(\system_inst.internal_param_c[4] ));
 sg13g2_dfrbp_1 _3714_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net28),
    .D(_0056_),
    .Q_N(_1817_),
    .Q(\system_inst.internal_param_c[5] ));
 sg13g2_dfrbp_1 _3715_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net24),
    .D(_0057_),
    .Q_N(_1816_),
    .Q(\system_inst.internal_param_d[0] ));
 sg13g2_dfrbp_1 _3716_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net81),
    .D(_0058_),
    .Q_N(_1815_),
    .Q(\system_inst.internal_param_d[1] ));
 sg13g2_dfrbp_1 _3717_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net77),
    .D(net125),
    .Q_N(_1814_),
    .Q(\system_inst.internal_param_d[2] ));
 sg13g2_dfrbp_1 _3718_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net73),
    .D(net101),
    .Q_N(_1813_),
    .Q(\system_inst.internal_param_d[3] ));
 sg13g2_dfrbp_1 _3719_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net63),
    .D(_0061_),
    .Q_N(_1812_),
    .Q(\system_inst.internal_param_d[4] ));
 sg13g2_dfrbp_1 _3720_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net59),
    .D(_0062_),
    .Q_N(_1811_),
    .Q(\system_inst.internal_param_d[5] ));
 sg13g2_dfrbp_1 _3721_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net55),
    .D(_0063_),
    .Q_N(_1810_),
    .Q(\system_inst.loader.shift_reg[0] ));
 sg13g2_dfrbp_1 _3722_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net51),
    .D(net105),
    .Q_N(_1809_),
    .Q(\system_inst.loader.shift_reg[1] ));
 sg13g2_dfrbp_1 _3723_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net47),
    .D(net128),
    .Q_N(_1808_),
    .Q(\system_inst.loader.shift_reg[2] ));
 sg13g2_dfrbp_1 _3724_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net43),
    .D(_0066_),
    .Q_N(_1807_),
    .Q(\system_inst.loader.shift_reg[3] ));
 sg13g2_dfrbp_1 _3725_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net39),
    .D(_0067_),
    .Q_N(_1806_),
    .Q(\system_inst.loader.shift_reg[4] ));
 sg13g2_dfrbp_1 _3726_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net35),
    .D(_0068_),
    .Q_N(_1805_),
    .Q(\system_inst.loader.bit_count[0] ));
 sg13g2_dfrbp_1 _3727_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net31),
    .D(_0069_),
    .Q_N(_1804_),
    .Q(\system_inst.loader.bit_count[1] ));
 sg13g2_dfrbp_1 _3728_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net66),
    .D(net107),
    .Q_N(_1834_),
    .Q(\system_inst.loader.bit_count[2] ));
 sg13g2_dfrbp_1 _3729_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net67),
    .D(_0000_),
    .Q_N(_1835_),
    .Q(\system_inst.loader.state[0] ));
 sg13g2_dfrbp_1 _3730_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net68),
    .D(_0001_),
    .Q_N(_0019_),
    .Q(\system_inst.loader.state[1] ));
 sg13g2_dfrbp_1 _3731_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net69),
    .D(_0002_),
    .Q_N(_1836_),
    .Q(\system_inst.loader.state[2] ));
 sg13g2_dfrbp_1 _3732_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net70),
    .D(_0003_),
    .Q_N(_1837_),
    .Q(\system_inst.loader.state[3] ));
 sg13g2_dfrbp_1 _3733_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net41),
    .D(_0004_),
    .Q_N(_1838_),
    .Q(\system_inst.loader.state[4] ));
 sg13g2_dfrbp_1 _3734_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net26),
    .D(_0005_),
    .Q_N(_1803_),
    .Q(\system_inst.loader.state[5] ));
 sg13g2_dfrbp_1 _3735_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net79),
    .D(_0071_),
    .Q_N(_1802_),
    .Q(spike_out_internal));
 sg13g2_dfrbp_1 _3736_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net75),
    .D(_0072_),
    .Q_N(_0006_),
    .Q(\system_inst.neuron.v[0] ));
 sg13g2_dfrbp_1 _3737_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net61),
    .D(_0073_),
    .Q_N(_0027_),
    .Q(\system_inst.neuron.v[1] ));
 sg13g2_dfrbp_1 _3738_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net53),
    .D(net97),
    .Q_N(_0026_),
    .Q(\system_inst.neuron.v[2] ));
 sg13g2_dfrbp_1 _3739_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net45),
    .D(_0075_),
    .Q_N(_0025_),
    .Q(\system_inst.neuron.v[3] ));
 sg13g2_dfrbp_1 _3740_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net37),
    .D(_0076_),
    .Q_N(_0023_),
    .Q(\system_inst.neuron.v[4] ));
 sg13g2_dfrbp_1 _3741_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net29),
    .D(_0077_),
    .Q_N(_0022_),
    .Q(\system_inst.neuron.v[5] ));
 sg13g2_dfrbp_1 _3742_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net71),
    .D(_0078_),
    .Q_N(_0021_),
    .Q(\system_inst.neuron.v[6] ));
 sg13g2_dfrbp_1 _3743_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net49),
    .D(_0079_),
    .Q_N(_1801_),
    .Q(\system_inst.neuron.v[7] ));
 sg13g2_dfrbp_1 _3744_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net33),
    .D(_0080_),
    .Q_N(_0009_),
    .Q(\system_inst.neuron.v[8] ));
 sg13g2_dfrbp_1 _3745_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net57),
    .D(_0081_),
    .Q_N(_0024_),
    .Q(\system_inst.neuron.v[9] ));
 sg13g2_dfrbp_1 _3746_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net22),
    .D(_0082_),
    .Q_N(_1800_),
    .Q(\system_inst.loader.load_enable_prev ));
 sg13g2_tiehi _3689__23 (.L_HI(net23));
 sg13g2_tiehi _3715__24 (.L_HI(net24));
 sg13g2_tiehi _3688__25 (.L_HI(net25));
 sg13g2_tiehi _3734__26 (.L_HI(net26));
 sg13g2_tiehi _3687__27 (.L_HI(net27));
 sg13g2_tiehi _3714__28 (.L_HI(net28));
 sg13g2_tiehi _3741__29 (.L_HI(net29));
 sg13g2_tiehi _3713__30 (.L_HI(net30));
 sg13g2_tiehi _3727__31 (.L_HI(net31));
 sg13g2_tiehi _3712__32 (.L_HI(net32));
 sg13g2_tiehi _3744__33 (.L_HI(net33));
 sg13g2_tiehi _3711__34 (.L_HI(net34));
 sg13g2_tiehi _3726__35 (.L_HI(net35));
 sg13g2_tiehi _3710__36 (.L_HI(net36));
 sg13g2_tiehi _3740__37 (.L_HI(net37));
 sg13g2_tiehi _3709__38 (.L_HI(net38));
 sg13g2_tiehi _3725__39 (.L_HI(net39));
 sg13g2_tiehi _3708__40 (.L_HI(net40));
 sg13g2_tiehi _3733__41 (.L_HI(net41));
 sg13g2_tiehi _3707__42 (.L_HI(net42));
 sg13g2_tiehi _3724__43 (.L_HI(net43));
 sg13g2_tiehi _3706__44 (.L_HI(net44));
 sg13g2_tiehi _3739__45 (.L_HI(net45));
 sg13g2_tiehi _3705__46 (.L_HI(net46));
 sg13g2_tiehi _3723__47 (.L_HI(net47));
 sg13g2_tiehi _3704__48 (.L_HI(net48));
 sg13g2_tiehi _3743__49 (.L_HI(net49));
 sg13g2_tiehi _3703__50 (.L_HI(net50));
 sg13g2_tiehi _3722__51 (.L_HI(net51));
 sg13g2_tiehi _3702__52 (.L_HI(net52));
 sg13g2_tiehi _3738__53 (.L_HI(net53));
 sg13g2_tiehi _3701__54 (.L_HI(net54));
 sg13g2_tiehi _3721__55 (.L_HI(net55));
 sg13g2_tiehi _3700__56 (.L_HI(net56));
 sg13g2_tiehi _3745__57 (.L_HI(net57));
 sg13g2_tiehi _3699__58 (.L_HI(net58));
 sg13g2_tiehi _3720__59 (.L_HI(net59));
 sg13g2_tiehi _3698__60 (.L_HI(net60));
 sg13g2_tiehi _3737__61 (.L_HI(net61));
 sg13g2_tiehi _3697__62 (.L_HI(net62));
 sg13g2_tiehi _3719__63 (.L_HI(net63));
 sg13g2_tiehi _3696__64 (.L_HI(net64));
 sg13g2_tiehi _3686__65 (.L_HI(net65));
 sg13g2_tiehi _3728__66 (.L_HI(net66));
 sg13g2_tiehi _3729__67 (.L_HI(net67));
 sg13g2_tiehi _3730__68 (.L_HI(net68));
 sg13g2_tiehi _3731__69 (.L_HI(net69));
 sg13g2_tiehi _3732__70 (.L_HI(net70));
 sg13g2_tiehi _3742__71 (.L_HI(net71));
 sg13g2_tiehi _3695__72 (.L_HI(net72));
 sg13g2_tiehi _3718__73 (.L_HI(net73));
 sg13g2_tiehi _3694__74 (.L_HI(net74));
 sg13g2_tiehi _3736__75 (.L_HI(net75));
 sg13g2_tiehi _3693__76 (.L_HI(net76));
 sg13g2_tiehi _3717__77 (.L_HI(net77));
 sg13g2_tiehi _3692__78 (.L_HI(net78));
 sg13g2_tiehi _3735__79 (.L_HI(net79));
 sg13g2_tiehi _3691__80 (.L_HI(net80));
 sg13g2_tiehi _3716__81 (.L_HI(net81));
 sg13g2_tiehi _3690__82 (.L_HI(net82));
 sg13g2_tiehi tt_um_izh_neuron_lite_83 (.L_HI(net83));
 sg13g2_tiehi tt_um_izh_neuron_lite_84 (.L_HI(net84));
 sg13g2_tiehi tt_um_izh_neuron_lite_85 (.L_HI(net85));
 sg13g2_tiehi tt_um_izh_neuron_lite_86 (.L_HI(net86));
 sg13g2_tiehi tt_um_izh_neuron_lite_87 (.L_HI(net87));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_izh_neuron_lite_14 (.L_LO(net14));
 sg13g2_tielo tt_um_izh_neuron_lite_15 (.L_LO(net15));
 sg13g2_tielo tt_um_izh_neuron_lite_16 (.L_LO(net16));
 sg13g2_tielo tt_um_izh_neuron_lite_17 (.L_LO(net17));
 sg13g2_tielo tt_um_izh_neuron_lite_18 (.L_LO(net18));
 sg13g2_tielo tt_um_izh_neuron_lite_19 (.L_LO(net19));
 sg13g2_tielo tt_um_izh_neuron_lite_20 (.L_LO(net20));
 sg13g2_tielo tt_um_izh_neuron_lite_21 (.L_LO(net21));
 sg13g2_tiehi _3746__22 (.L_HI(net22));
 sg13g2_buf_1 _3822_ (.A(spike_out_internal),
    .X(uio_out[0]));
 sg13g2_buf_2 _3823_ (.A(params_ready_internal),
    .X(uio_out[1]));
 sg13g2_buf_2 fanout324 (.A(_0937_),
    .X(net324));
 sg13g2_buf_1 fanout325 (.A(_0937_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_1351_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_1349_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_1479_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_1506_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_0096_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_0156_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_0156_),
    .X(net332));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(_0155_));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(net336));
 sg13g2_buf_1 fanout335 (.A(net336),
    .X(net335));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(_1063_));
 sg13g2_buf_2 fanout337 (.A(net338),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_1058_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_1054_),
    .X(net339));
 sg13g2_buf_1 fanout340 (.A(_1054_),
    .X(net340));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(_1040_));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(_0183_));
 sg13g2_buf_1 fanout343 (.A(_0183_),
    .X(net343));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(net345));
 sg13g2_buf_2 fanout345 (.A(net346),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_1681_),
    .X(net346));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(_1680_));
 sg13g2_buf_1 fanout348 (.A(_1680_),
    .X(net348));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(_0713_));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(net352));
 sg13g2_buf_1 fanout351 (.A(net352),
    .X(net351));
 sg13g2_buf_1 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(\system_inst.neuron.v[9] ));
 sg13g2_buf_2 fanout354 (.A(\system_inst.neuron.v[9] ),
    .X(net354));
 sg13g2_buf_1 fanout355 (.A(\system_inst.neuron.v[9] ),
    .X(net355));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(net358));
 sg13g2_buf_2 fanout357 (.A(net358),
    .X(net357));
 sg13g2_buf_4 fanout358 (.X(net358),
    .A(\system_inst.neuron.v[8] ));
 sg13g2_buf_2 fanout359 (.A(net360),
    .X(net359));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(\system_inst.neuron.v[7] ));
 sg13g2_buf_2 fanout361 (.A(net362),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(\system_inst.neuron.v[7] ),
    .X(net362));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(net366));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(net366));
 sg13g2_buf_2 fanout365 (.A(net366),
    .X(net365));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(\system_inst.neuron.v[6] ));
 sg13g2_buf_2 fanout367 (.A(net368),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(net369),
    .X(net368));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(net370));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(\system_inst.neuron.v[5] ));
 sg13g2_buf_2 fanout371 (.A(net372),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(net374),
    .X(net372));
 sg13g2_buf_4 fanout373 (.X(net373),
    .A(net374));
 sg13g2_buf_4 fanout374 (.X(net374),
    .A(\system_inst.neuron.v[4] ));
 sg13g2_buf_2 fanout375 (.A(net376),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(net377),
    .X(net376));
 sg13g2_buf_4 fanout377 (.X(net377),
    .A(\system_inst.neuron.v[3] ));
 sg13g2_buf_4 fanout378 (.X(net378),
    .A(\system_inst.neuron.v[3] ));
 sg13g2_buf_2 fanout379 (.A(net380),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(net381),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(net383),
    .X(net381));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(net383));
 sg13g2_buf_2 fanout383 (.A(\system_inst.neuron.v[2] ),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(net389),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(net386),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(net389),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(net388),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(net389),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(\system_inst.neuron.v[1] ),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(net394),
    .X(net390));
 sg13g2_buf_4 fanout391 (.X(net391),
    .A(net394));
 sg13g2_buf_2 fanout392 (.A(net393),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(net394),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(net149),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(net396),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(\system_inst.internal_param_b[5] ),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(\system_inst.internal_param_b[4] ),
    .X(net397));
 sg13g2_buf_1 fanout398 (.A(\system_inst.internal_param_b[4] ),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(net400),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(net145),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(net151),
    .X(net401));
 sg13g2_buf_1 fanout402 (.A(\system_inst.internal_param_b[2] ),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(net404),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(net133),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(net156),
    .X(net405));
 sg13g2_buf_4 fanout406 (.X(net406),
    .A(\system_inst.internal_param_a[4] ));
 sg13g2_buf_2 fanout407 (.A(net132),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(net409),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(\system_inst.internal_param_a[3] ),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(\system_inst.internal_param_a[1] ),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(\system_inst.internal_param_a[1] ),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(net414),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(\system_inst.internal_param_a[0] ),
    .X(net414));
 sg13g2_buf_4 fanout415 (.X(net415),
    .A(\system_inst.neuron.u[9] ));
 sg13g2_buf_4 fanout416 (.X(net416),
    .A(net155));
 sg13g2_buf_2 fanout417 (.A(net418),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_0974_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(net420),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_0974_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(net424),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(net424),
    .X(net422));
 sg13g2_buf_1 fanout423 (.A(net424),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(rst_n),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(net426),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(rst_n),
    .X(net426));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[2]),
    .X(net12));
 sg13g2_tielo tt_um_izh_neuron_lite_13 (.L_LO(net13));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_0007_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold2 (.A(\system_inst.internal_param_c[3] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0054_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0020_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0036_),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold6 (.A(\system_inst.loader.state[3] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold7 (.A(_1050_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold8 (.A(\system_inst.neuron.v[5] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold9 (.A(\system_inst.internal_param_c[0] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0074_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold11 (.A(\system_inst.internal_param_c[1] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0973_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold13 (.A(\system_inst.internal_param_d[3] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0060_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold15 (.A(\system_inst.loader.state[1] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold16 (.A(_1045_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold17 (.A(\system_inst.loader.shift_reg[0] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0064_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold19 (.A(\system_inst.loader.bit_count[2] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0070_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold21 (.A(\system_inst.loader.state[5] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold22 (.A(\system_inst.loader.shift_reg[4] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0050_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold24 (.A(\system_inst.loader.state[2] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold25 (.A(\system_inst.internal_param_d[5] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold26 (.A(\system_inst.internal_param_c[2] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0053_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold28 (.A(\system_inst.internal_param_c[5] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold29 (.A(\system_inst.loader.state[4] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold30 (.A(_1055_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold31 (.A(\system_inst.internal_param_c[4] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0055_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold33 (.A(\system_inst.loader.shift_reg[3] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold34 (.A(\system_inst.internal_param_a[5] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold35 (.A(\system_inst.loader.bit_count[1] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0114_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold37 (.A(\system_inst.internal_param_d[2] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0059_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold39 (.A(\system_inst.internal_param_d[4] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold40 (.A(\system_inst.loader.shift_reg[1] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0065_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold42 (.A(\system_inst.loader.state[0] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold43 (.A(_1056_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold44 (.A(params_ready_internal),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold45 (.A(\system_inst.internal_param_a[4] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold46 (.A(\system_inst.internal_param_b[1] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold47 (.A(\system_inst.internal_param_b[4] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold48 (.A(\system_inst.internal_param_d[1] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0006_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold50 (.A(\system_inst.loader.shift_reg[2] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold51 (.A(\system_inst.loader.bit_count[0] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0109_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold53 (.A(\system_inst.internal_param_d[0] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0013_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0028_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0010_),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0034_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold58 (.A(\system_inst.internal_param_b[3] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold59 (.A(\system_inst.internal_param_a[2] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold60 (.A(\system_inst.neuron.u[8] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0035_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold62 (.A(\system_inst.neuron.v[0] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold63 (.A(\system_inst.neuron.u[4] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold64 (.A(\system_inst.internal_param_b[2] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0047_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold66 (.A(\system_inst.neuron.u[2] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold67 (.A(\system_inst.neuron.u[0] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold68 (.A(\system_inst.neuron.u[5] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold69 (.A(\system_inst.internal_param_b[0] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold70 (.A(\system_inst.neuron.u[3] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold71 (.A(\system_inst.neuron.u[6] ),
    .X(net158));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_fill_1 FILLER_0_140 ();
 sg13g2_decap_4 FILLER_0_153 ();
 sg13g2_decap_8 FILLER_0_162 ();
 sg13g2_decap_4 FILLER_0_169 ();
 sg13g2_decap_4 FILLER_0_185 ();
 sg13g2_fill_1 FILLER_0_193 ();
 sg13g2_fill_2 FILLER_0_206 ();
 sg13g2_fill_1 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_226 ();
 sg13g2_decap_8 FILLER_0_233 ();
 sg13g2_decap_8 FILLER_0_240 ();
 sg13g2_decap_4 FILLER_0_247 ();
 sg13g2_fill_2 FILLER_0_256 ();
 sg13g2_fill_1 FILLER_0_258 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_4 FILLER_0_299 ();
 sg13g2_fill_2 FILLER_0_303 ();
 sg13g2_fill_2 FILLER_0_309 ();
 sg13g2_fill_1 FILLER_0_311 ();
 sg13g2_decap_4 FILLER_0_329 ();
 sg13g2_fill_2 FILLER_0_333 ();
 sg13g2_fill_2 FILLER_0_356 ();
 sg13g2_fill_1 FILLER_0_358 ();
 sg13g2_fill_2 FILLER_0_392 ();
 sg13g2_fill_2 FILLER_0_398 ();
 sg13g2_fill_1 FILLER_0_400 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_fill_2 FILLER_1_126 ();
 sg13g2_fill_1 FILLER_1_128 ();
 sg13g2_fill_2 FILLER_1_141 ();
 sg13g2_fill_1 FILLER_1_143 ();
 sg13g2_fill_1 FILLER_1_166 ();
 sg13g2_decap_8 FILLER_1_200 ();
 sg13g2_fill_1 FILLER_1_207 ();
 sg13g2_fill_1 FILLER_1_231 ();
 sg13g2_fill_1 FILLER_1_257 ();
 sg13g2_fill_2 FILLER_1_278 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_291 ();
 sg13g2_fill_1 FILLER_1_318 ();
 sg13g2_fill_2 FILLER_1_331 ();
 sg13g2_fill_1 FILLER_1_333 ();
 sg13g2_fill_2 FILLER_1_391 ();
 sg13g2_fill_1 FILLER_1_393 ();
 sg13g2_fill_1 FILLER_1_398 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_4 FILLER_2_112 ();
 sg13g2_fill_2 FILLER_2_116 ();
 sg13g2_fill_2 FILLER_2_123 ();
 sg13g2_fill_1 FILLER_2_125 ();
 sg13g2_fill_2 FILLER_2_139 ();
 sg13g2_decap_4 FILLER_2_162 ();
 sg13g2_fill_1 FILLER_2_166 ();
 sg13g2_fill_2 FILLER_2_176 ();
 sg13g2_fill_2 FILLER_2_187 ();
 sg13g2_fill_2 FILLER_2_204 ();
 sg13g2_fill_1 FILLER_2_206 ();
 sg13g2_fill_2 FILLER_2_232 ();
 sg13g2_fill_1 FILLER_2_234 ();
 sg13g2_fill_1 FILLER_2_247 ();
 sg13g2_fill_2 FILLER_2_253 ();
 sg13g2_fill_1 FILLER_2_255 ();
 sg13g2_fill_2 FILLER_2_261 ();
 sg13g2_decap_4 FILLER_2_268 ();
 sg13g2_fill_2 FILLER_2_272 ();
 sg13g2_decap_8 FILLER_2_293 ();
 sg13g2_fill_2 FILLER_2_300 ();
 sg13g2_fill_1 FILLER_2_302 ();
 sg13g2_fill_2 FILLER_2_328 ();
 sg13g2_fill_2 FILLER_2_379 ();
 sg13g2_fill_1 FILLER_2_381 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_4 FILLER_3_98 ();
 sg13g2_fill_2 FILLER_3_102 ();
 sg13g2_fill_1 FILLER_3_128 ();
 sg13g2_fill_2 FILLER_3_142 ();
 sg13g2_fill_2 FILLER_3_149 ();
 sg13g2_fill_1 FILLER_3_159 ();
 sg13g2_fill_2 FILLER_3_177 ();
 sg13g2_fill_1 FILLER_3_179 ();
 sg13g2_fill_2 FILLER_3_200 ();
 sg13g2_fill_1 FILLER_3_215 ();
 sg13g2_fill_1 FILLER_3_221 ();
 sg13g2_fill_2 FILLER_3_233 ();
 sg13g2_fill_2 FILLER_3_245 ();
 sg13g2_fill_1 FILLER_3_247 ();
 sg13g2_fill_2 FILLER_3_338 ();
 sg13g2_fill_1 FILLER_3_349 ();
 sg13g2_fill_2 FILLER_3_380 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_fill_2 FILLER_4_105 ();
 sg13g2_decap_4 FILLER_4_120 ();
 sg13g2_fill_2 FILLER_4_134 ();
 sg13g2_fill_1 FILLER_4_171 ();
 sg13g2_fill_1 FILLER_4_210 ();
 sg13g2_fill_2 FILLER_4_235 ();
 sg13g2_fill_2 FILLER_4_246 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_265 ();
 sg13g2_fill_2 FILLER_4_272 ();
 sg13g2_decap_4 FILLER_4_280 ();
 sg13g2_fill_1 FILLER_4_284 ();
 sg13g2_decap_4 FILLER_4_298 ();
 sg13g2_fill_2 FILLER_4_320 ();
 sg13g2_fill_2 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_fill_2 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_38 ();
 sg13g2_decap_8 FILLER_5_44 ();
 sg13g2_decap_4 FILLER_5_51 ();
 sg13g2_fill_2 FILLER_5_55 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_85 ();
 sg13g2_decap_4 FILLER_5_92 ();
 sg13g2_fill_1 FILLER_5_96 ();
 sg13g2_decap_4 FILLER_5_107 ();
 sg13g2_fill_2 FILLER_5_111 ();
 sg13g2_fill_2 FILLER_5_122 ();
 sg13g2_fill_1 FILLER_5_124 ();
 sg13g2_decap_4 FILLER_5_135 ();
 sg13g2_fill_1 FILLER_5_139 ();
 sg13g2_fill_2 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_165 ();
 sg13g2_fill_1 FILLER_5_167 ();
 sg13g2_fill_1 FILLER_5_173 ();
 sg13g2_fill_1 FILLER_5_187 ();
 sg13g2_fill_1 FILLER_5_192 ();
 sg13g2_decap_4 FILLER_5_200 ();
 sg13g2_fill_1 FILLER_5_204 ();
 sg13g2_fill_1 FILLER_5_218 ();
 sg13g2_fill_2 FILLER_5_232 ();
 sg13g2_fill_1 FILLER_5_234 ();
 sg13g2_fill_1 FILLER_5_248 ();
 sg13g2_fill_1 FILLER_5_280 ();
 sg13g2_fill_2 FILLER_5_296 ();
 sg13g2_decap_8 FILLER_5_320 ();
 sg13g2_fill_1 FILLER_5_327 ();
 sg13g2_fill_1 FILLER_5_343 ();
 sg13g2_fill_2 FILLER_5_360 ();
 sg13g2_fill_1 FILLER_5_385 ();
 sg13g2_fill_2 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_18 ();
 sg13g2_fill_1 FILLER_6_60 ();
 sg13g2_fill_2 FILLER_6_110 ();
 sg13g2_fill_1 FILLER_6_161 ();
 sg13g2_fill_1 FILLER_6_188 ();
 sg13g2_decap_8 FILLER_6_205 ();
 sg13g2_fill_2 FILLER_6_212 ();
 sg13g2_fill_1 FILLER_6_214 ();
 sg13g2_fill_1 FILLER_6_231 ();
 sg13g2_fill_1 FILLER_6_248 ();
 sg13g2_fill_1 FILLER_6_252 ();
 sg13g2_fill_2 FILLER_6_257 ();
 sg13g2_fill_2 FILLER_6_316 ();
 sg13g2_fill_1 FILLER_6_318 ();
 sg13g2_fill_1 FILLER_6_329 ();
 sg13g2_fill_1 FILLER_6_361 ();
 sg13g2_fill_2 FILLER_6_379 ();
 sg13g2_fill_2 FILLER_6_391 ();
 sg13g2_fill_1 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_23 ();
 sg13g2_fill_1 FILLER_7_30 ();
 sg13g2_fill_1 FILLER_7_36 ();
 sg13g2_decap_8 FILLER_7_45 ();
 sg13g2_decap_4 FILLER_7_52 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_74 ();
 sg13g2_decap_8 FILLER_7_80 ();
 sg13g2_fill_2 FILLER_7_87 ();
 sg13g2_fill_1 FILLER_7_89 ();
 sg13g2_fill_2 FILLER_7_107 ();
 sg13g2_decap_8 FILLER_7_116 ();
 sg13g2_fill_1 FILLER_7_128 ();
 sg13g2_decap_4 FILLER_7_134 ();
 sg13g2_fill_1 FILLER_7_138 ();
 sg13g2_decap_4 FILLER_7_160 ();
 sg13g2_fill_2 FILLER_7_207 ();
 sg13g2_decap_4 FILLER_7_229 ();
 sg13g2_fill_2 FILLER_7_238 ();
 sg13g2_fill_1 FILLER_7_240 ();
 sg13g2_fill_2 FILLER_7_258 ();
 sg13g2_fill_1 FILLER_7_267 ();
 sg13g2_fill_1 FILLER_7_278 ();
 sg13g2_fill_2 FILLER_7_289 ();
 sg13g2_fill_1 FILLER_7_343 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_28 ();
 sg13g2_fill_1 FILLER_8_30 ();
 sg13g2_fill_1 FILLER_8_100 ();
 sg13g2_fill_2 FILLER_8_114 ();
 sg13g2_fill_1 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_152 ();
 sg13g2_fill_1 FILLER_8_159 ();
 sg13g2_fill_2 FILLER_8_169 ();
 sg13g2_fill_1 FILLER_8_171 ();
 sg13g2_fill_1 FILLER_8_182 ();
 sg13g2_fill_2 FILLER_8_191 ();
 sg13g2_fill_1 FILLER_8_193 ();
 sg13g2_decap_8 FILLER_8_207 ();
 sg13g2_decap_4 FILLER_8_214 ();
 sg13g2_fill_1 FILLER_8_218 ();
 sg13g2_fill_2 FILLER_8_239 ();
 sg13g2_fill_1 FILLER_8_241 ();
 sg13g2_fill_2 FILLER_8_255 ();
 sg13g2_decap_4 FILLER_8_265 ();
 sg13g2_fill_2 FILLER_8_278 ();
 sg13g2_fill_2 FILLER_8_312 ();
 sg13g2_fill_2 FILLER_8_319 ();
 sg13g2_fill_2 FILLER_8_326 ();
 sg13g2_fill_2 FILLER_8_332 ();
 sg13g2_fill_1 FILLER_8_334 ();
 sg13g2_fill_2 FILLER_8_366 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_4 ();
 sg13g2_fill_2 FILLER_9_47 ();
 sg13g2_fill_1 FILLER_9_49 ();
 sg13g2_fill_1 FILLER_9_79 ();
 sg13g2_decap_8 FILLER_9_85 ();
 sg13g2_fill_2 FILLER_9_99 ();
 sg13g2_fill_1 FILLER_9_101 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_decap_4 FILLER_9_130 ();
 sg13g2_fill_2 FILLER_9_134 ();
 sg13g2_fill_1 FILLER_9_157 ();
 sg13g2_fill_2 FILLER_9_179 ();
 sg13g2_fill_1 FILLER_9_181 ();
 sg13g2_fill_2 FILLER_9_209 ();
 sg13g2_fill_1 FILLER_9_211 ();
 sg13g2_decap_4 FILLER_9_217 ();
 sg13g2_fill_2 FILLER_9_235 ();
 sg13g2_fill_2 FILLER_9_251 ();
 sg13g2_fill_1 FILLER_9_253 ();
 sg13g2_fill_1 FILLER_9_360 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_fill_2 FILLER_10_23 ();
 sg13g2_fill_2 FILLER_10_38 ();
 sg13g2_fill_1 FILLER_10_40 ();
 sg13g2_decap_4 FILLER_10_59 ();
 sg13g2_fill_1 FILLER_10_63 ();
 sg13g2_decap_4 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_124 ();
 sg13g2_decap_4 FILLER_10_149 ();
 sg13g2_fill_2 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_176 ();
 sg13g2_decap_4 FILLER_10_183 ();
 sg13g2_fill_1 FILLER_10_187 ();
 sg13g2_fill_1 FILLER_10_245 ();
 sg13g2_fill_1 FILLER_10_277 ();
 sg13g2_fill_1 FILLER_10_305 ();
 sg13g2_fill_2 FILLER_10_320 ();
 sg13g2_fill_1 FILLER_10_343 ();
 sg13g2_fill_1 FILLER_10_354 ();
 sg13g2_fill_2 FILLER_10_360 ();
 sg13g2_fill_1 FILLER_10_367 ();
 sg13g2_fill_2 FILLER_10_381 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_15 ();
 sg13g2_fill_2 FILLER_11_29 ();
 sg13g2_fill_1 FILLER_11_49 ();
 sg13g2_decap_4 FILLER_11_75 ();
 sg13g2_decap_4 FILLER_11_89 ();
 sg13g2_fill_2 FILLER_11_122 ();
 sg13g2_fill_1 FILLER_11_148 ();
 sg13g2_fill_2 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_176 ();
 sg13g2_fill_1 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_320 ();
 sg13g2_fill_2 FILLER_11_396 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_fill_2 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_23 ();
 sg13g2_fill_1 FILLER_12_27 ();
 sg13g2_fill_2 FILLER_12_50 ();
 sg13g2_fill_1 FILLER_12_52 ();
 sg13g2_fill_2 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_97 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_fill_2 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_128 ();
 sg13g2_decap_4 FILLER_12_146 ();
 sg13g2_fill_1 FILLER_12_154 ();
 sg13g2_fill_1 FILLER_12_160 ();
 sg13g2_fill_1 FILLER_12_182 ();
 sg13g2_fill_2 FILLER_12_200 ();
 sg13g2_fill_1 FILLER_12_202 ();
 sg13g2_fill_2 FILLER_12_271 ();
 sg13g2_fill_2 FILLER_12_323 ();
 sg13g2_fill_2 FILLER_12_354 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_26 ();
 sg13g2_fill_2 FILLER_13_92 ();
 sg13g2_fill_2 FILLER_13_145 ();
 sg13g2_fill_1 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_178 ();
 sg13g2_fill_2 FILLER_13_209 ();
 sg13g2_fill_2 FILLER_13_248 ();
 sg13g2_fill_1 FILLER_13_304 ();
 sg13g2_fill_2 FILLER_13_368 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_2 FILLER_14_20 ();
 sg13g2_fill_1 FILLER_14_22 ();
 sg13g2_fill_2 FILLER_14_39 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_63 ();
 sg13g2_decap_4 FILLER_14_70 ();
 sg13g2_fill_2 FILLER_14_83 ();
 sg13g2_fill_1 FILLER_14_85 ();
 sg13g2_fill_2 FILLER_14_90 ();
 sg13g2_fill_1 FILLER_14_92 ();
 sg13g2_decap_8 FILLER_14_101 ();
 sg13g2_decap_4 FILLER_14_116 ();
 sg13g2_fill_2 FILLER_14_157 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_decap_4 FILLER_14_211 ();
 sg13g2_decap_4 FILLER_14_220 ();
 sg13g2_fill_2 FILLER_14_253 ();
 sg13g2_fill_1 FILLER_14_263 ();
 sg13g2_fill_2 FILLER_14_317 ();
 sg13g2_fill_2 FILLER_14_339 ();
 sg13g2_fill_1 FILLER_14_375 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_30 ();
 sg13g2_fill_2 FILLER_15_44 ();
 sg13g2_fill_1 FILLER_15_46 ();
 sg13g2_fill_2 FILLER_15_76 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_fill_1 FILLER_15_84 ();
 sg13g2_fill_2 FILLER_15_93 ();
 sg13g2_fill_1 FILLER_15_95 ();
 sg13g2_fill_2 FILLER_15_101 ();
 sg13g2_fill_2 FILLER_15_129 ();
 sg13g2_fill_1 FILLER_15_135 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_fill_1 FILLER_15_204 ();
 sg13g2_fill_1 FILLER_15_274 ();
 sg13g2_fill_1 FILLER_15_329 ();
 sg13g2_fill_1 FILLER_15_364 ();
 sg13g2_fill_2 FILLER_15_375 ();
 sg13g2_fill_1 FILLER_15_382 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_2 FILLER_16_24 ();
 sg13g2_fill_2 FILLER_16_55 ();
 sg13g2_fill_1 FILLER_16_57 ();
 sg13g2_fill_2 FILLER_16_87 ();
 sg13g2_fill_1 FILLER_16_89 ();
 sg13g2_fill_2 FILLER_16_106 ();
 sg13g2_fill_1 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_128 ();
 sg13g2_decap_4 FILLER_16_151 ();
 sg13g2_fill_2 FILLER_16_159 ();
 sg13g2_fill_1 FILLER_16_161 ();
 sg13g2_fill_2 FILLER_16_167 ();
 sg13g2_fill_1 FILLER_16_169 ();
 sg13g2_fill_2 FILLER_16_186 ();
 sg13g2_fill_2 FILLER_16_201 ();
 sg13g2_fill_1 FILLER_16_211 ();
 sg13g2_fill_1 FILLER_16_217 ();
 sg13g2_fill_1 FILLER_16_228 ();
 sg13g2_fill_1 FILLER_16_274 ();
 sg13g2_fill_1 FILLER_16_284 ();
 sg13g2_fill_2 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_25 ();
 sg13g2_fill_1 FILLER_17_45 ();
 sg13g2_decap_4 FILLER_17_51 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_fill_2 FILLER_17_68 ();
 sg13g2_fill_2 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_100 ();
 sg13g2_fill_2 FILLER_17_106 ();
 sg13g2_fill_1 FILLER_17_116 ();
 sg13g2_fill_2 FILLER_17_125 ();
 sg13g2_fill_1 FILLER_17_127 ();
 sg13g2_fill_2 FILLER_17_133 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_fill_2 FILLER_17_180 ();
 sg13g2_fill_1 FILLER_17_182 ();
 sg13g2_fill_2 FILLER_17_191 ();
 sg13g2_fill_1 FILLER_17_218 ();
 sg13g2_fill_2 FILLER_17_281 ();
 sg13g2_fill_2 FILLER_17_355 ();
 sg13g2_fill_1 FILLER_17_366 ();
 sg13g2_fill_1 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_29 ();
 sg13g2_fill_2 FILLER_18_55 ();
 sg13g2_fill_2 FILLER_18_109 ();
 sg13g2_fill_1 FILLER_18_111 ();
 sg13g2_fill_2 FILLER_18_120 ();
 sg13g2_fill_1 FILLER_18_122 ();
 sg13g2_fill_2 FILLER_18_152 ();
 sg13g2_fill_2 FILLER_18_176 ();
 sg13g2_fill_1 FILLER_18_178 ();
 sg13g2_fill_1 FILLER_18_208 ();
 sg13g2_fill_2 FILLER_18_214 ();
 sg13g2_fill_2 FILLER_18_233 ();
 sg13g2_fill_2 FILLER_18_244 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_fill_2 FILLER_18_276 ();
 sg13g2_fill_1 FILLER_18_357 ();
 sg13g2_fill_1 FILLER_18_394 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_31 ();
 sg13g2_fill_1 FILLER_19_38 ();
 sg13g2_decap_8 FILLER_19_53 ();
 sg13g2_fill_2 FILLER_19_60 ();
 sg13g2_decap_4 FILLER_19_83 ();
 sg13g2_fill_2 FILLER_19_87 ();
 sg13g2_fill_2 FILLER_19_111 ();
 sg13g2_fill_2 FILLER_19_123 ();
 sg13g2_fill_2 FILLER_19_157 ();
 sg13g2_decap_4 FILLER_19_163 ();
 sg13g2_fill_1 FILLER_19_167 ();
 sg13g2_fill_2 FILLER_19_185 ();
 sg13g2_decap_8 FILLER_19_204 ();
 sg13g2_fill_1 FILLER_19_239 ();
 sg13g2_fill_1 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_4 ();
 sg13g2_fill_2 FILLER_20_34 ();
 sg13g2_fill_2 FILLER_20_58 ();
 sg13g2_fill_2 FILLER_20_83 ();
 sg13g2_fill_2 FILLER_20_93 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_fill_1 FILLER_20_113 ();
 sg13g2_fill_2 FILLER_20_127 ();
 sg13g2_fill_2 FILLER_20_183 ();
 sg13g2_decap_4 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_272 ();
 sg13g2_fill_1 FILLER_20_274 ();
 sg13g2_fill_1 FILLER_20_324 ();
 sg13g2_fill_1 FILLER_20_330 ();
 sg13g2_fill_1 FILLER_20_363 ();
 sg13g2_fill_1 FILLER_20_373 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_1 FILLER_21_19 ();
 sg13g2_fill_2 FILLER_21_33 ();
 sg13g2_fill_2 FILLER_21_47 ();
 sg13g2_decap_8 FILLER_21_62 ();
 sg13g2_decap_8 FILLER_21_93 ();
 sg13g2_fill_2 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_122 ();
 sg13g2_decap_8 FILLER_21_129 ();
 sg13g2_decap_4 FILLER_21_136 ();
 sg13g2_fill_2 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_152 ();
 sg13g2_fill_2 FILLER_21_161 ();
 sg13g2_fill_1 FILLER_21_163 ();
 sg13g2_decap_8 FILLER_21_188 ();
 sg13g2_fill_2 FILLER_21_208 ();
 sg13g2_fill_1 FILLER_21_210 ();
 sg13g2_fill_2 FILLER_21_223 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_235 ();
 sg13g2_fill_2 FILLER_21_248 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_fill_2 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_299 ();
 sg13g2_fill_1 FILLER_21_384 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_7 ();
 sg13g2_decap_4 FILLER_22_51 ();
 sg13g2_fill_1 FILLER_22_75 ();
 sg13g2_fill_2 FILLER_22_102 ();
 sg13g2_fill_1 FILLER_22_104 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_decap_4 FILLER_22_141 ();
 sg13g2_fill_2 FILLER_22_145 ();
 sg13g2_fill_2 FILLER_22_189 ();
 sg13g2_fill_1 FILLER_22_191 ();
 sg13g2_fill_1 FILLER_22_196 ();
 sg13g2_fill_1 FILLER_22_209 ();
 sg13g2_decap_4 FILLER_22_215 ();
 sg13g2_fill_2 FILLER_22_219 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_254 ();
 sg13g2_fill_1 FILLER_22_295 ();
 sg13g2_fill_2 FILLER_22_311 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_fill_2 FILLER_23_14 ();
 sg13g2_fill_1 FILLER_23_16 ();
 sg13g2_fill_1 FILLER_23_40 ();
 sg13g2_decap_4 FILLER_23_46 ();
 sg13g2_fill_1 FILLER_23_58 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_decap_4 FILLER_23_102 ();
 sg13g2_fill_2 FILLER_23_111 ();
 sg13g2_fill_1 FILLER_23_113 ();
 sg13g2_decap_4 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_130 ();
 sg13g2_fill_2 FILLER_23_155 ();
 sg13g2_fill_1 FILLER_23_157 ();
 sg13g2_fill_1 FILLER_23_163 ();
 sg13g2_fill_1 FILLER_23_181 ();
 sg13g2_decap_4 FILLER_23_190 ();
 sg13g2_fill_2 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_217 ();
 sg13g2_fill_1 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_fill_2 FILLER_23_341 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_23 ();
 sg13g2_fill_2 FILLER_24_41 ();
 sg13g2_fill_1 FILLER_24_72 ();
 sg13g2_fill_2 FILLER_24_86 ();
 sg13g2_fill_1 FILLER_24_88 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_fill_2 FILLER_24_114 ();
 sg13g2_fill_1 FILLER_24_116 ();
 sg13g2_fill_2 FILLER_24_133 ();
 sg13g2_fill_1 FILLER_24_135 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_224 ();
 sg13g2_fill_2 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_fill_2 FILLER_24_254 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_fill_2 FILLER_24_282 ();
 sg13g2_fill_1 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_291 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_1 FILLER_25_37 ();
 sg13g2_fill_2 FILLER_25_57 ();
 sg13g2_fill_1 FILLER_25_59 ();
 sg13g2_fill_2 FILLER_25_76 ();
 sg13g2_fill_2 FILLER_25_94 ();
 sg13g2_fill_1 FILLER_25_96 ();
 sg13g2_decap_4 FILLER_25_106 ();
 sg13g2_fill_2 FILLER_25_110 ();
 sg13g2_fill_2 FILLER_25_133 ();
 sg13g2_fill_2 FILLER_25_144 ();
 sg13g2_fill_1 FILLER_25_146 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_167 ();
 sg13g2_fill_1 FILLER_25_169 ();
 sg13g2_decap_4 FILLER_25_190 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_250 ();
 sg13g2_fill_1 FILLER_25_256 ();
 sg13g2_fill_1 FILLER_25_267 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_fill_1 FILLER_25_283 ();
 sg13g2_fill_1 FILLER_25_360 ();
 sg13g2_fill_1 FILLER_25_392 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_32 ();
 sg13g2_decap_4 FILLER_26_37 ();
 sg13g2_fill_2 FILLER_26_41 ();
 sg13g2_fill_2 FILLER_26_57 ();
 sg13g2_fill_1 FILLER_26_59 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_fill_1 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_81 ();
 sg13g2_fill_2 FILLER_26_89 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_fill_2 FILLER_26_121 ();
 sg13g2_decap_4 FILLER_26_140 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_fill_2 FILLER_26_238 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_fill_1 FILLER_26_332 ();
 sg13g2_fill_2 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_389 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_2 FILLER_27_23 ();
 sg13g2_fill_1 FILLER_27_25 ();
 sg13g2_fill_1 FILLER_27_47 ();
 sg13g2_decap_4 FILLER_27_83 ();
 sg13g2_fill_2 FILLER_27_100 ();
 sg13g2_fill_2 FILLER_27_107 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_fill_2 FILLER_27_125 ();
 sg13g2_decap_4 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_fill_1 FILLER_27_252 ();
 sg13g2_fill_2 FILLER_27_343 ();
 sg13g2_fill_1 FILLER_27_368 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_30 ();
 sg13g2_fill_1 FILLER_28_40 ();
 sg13g2_fill_2 FILLER_28_62 ();
 sg13g2_fill_2 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_116 ();
 sg13g2_fill_1 FILLER_28_118 ();
 sg13g2_fill_1 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_135 ();
 sg13g2_decap_8 FILLER_28_159 ();
 sg13g2_fill_1 FILLER_28_192 ();
 sg13g2_fill_2 FILLER_28_222 ();
 sg13g2_fill_2 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_270 ();
 sg13g2_fill_2 FILLER_28_281 ();
 sg13g2_fill_2 FILLER_28_367 ();
 sg13g2_fill_2 FILLER_28_375 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_9 ();
 sg13g2_decap_4 FILLER_29_47 ();
 sg13g2_fill_1 FILLER_29_85 ();
 sg13g2_fill_1 FILLER_29_91 ();
 sg13g2_fill_1 FILLER_29_102 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_fill_2 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_118 ();
 sg13g2_fill_2 FILLER_29_139 ();
 sg13g2_fill_1 FILLER_29_141 ();
 sg13g2_decap_4 FILLER_29_152 ();
 sg13g2_fill_1 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_209 ();
 sg13g2_fill_2 FILLER_29_223 ();
 sg13g2_fill_1 FILLER_29_225 ();
 sg13g2_fill_1 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_355 ();
 sg13g2_fill_2 FILLER_29_375 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_32 ();
 sg13g2_decap_4 FILLER_30_45 ();
 sg13g2_fill_1 FILLER_30_49 ();
 sg13g2_fill_1 FILLER_30_80 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_decap_4 FILLER_30_131 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_172 ();
 sg13g2_fill_1 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_fill_2 FILLER_30_198 ();
 sg13g2_fill_1 FILLER_30_200 ();
 sg13g2_fill_2 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_247 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_fill_2 FILLER_30_309 ();
 sg13g2_fill_1 FILLER_30_311 ();
 sg13g2_fill_2 FILLER_30_382 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_16 ();
 sg13g2_decap_4 FILLER_31_27 ();
 sg13g2_fill_1 FILLER_31_31 ();
 sg13g2_fill_2 FILLER_31_40 ();
 sg13g2_fill_1 FILLER_31_50 ();
 sg13g2_fill_2 FILLER_31_54 ();
 sg13g2_fill_1 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_67 ();
 sg13g2_decap_4 FILLER_31_86 ();
 sg13g2_fill_1 FILLER_31_90 ();
 sg13g2_fill_2 FILLER_31_103 ();
 sg13g2_fill_1 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_111 ();
 sg13g2_decap_4 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_132 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_fill_2 FILLER_31_153 ();
 sg13g2_fill_1 FILLER_31_165 ();
 sg13g2_fill_2 FILLER_31_180 ();
 sg13g2_fill_2 FILLER_31_189 ();
 sg13g2_fill_2 FILLER_31_220 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_fill_2 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_244 ();
 sg13g2_fill_1 FILLER_31_270 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_fill_1 FILLER_31_369 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_28 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_decap_4 FILLER_32_52 ();
 sg13g2_fill_1 FILLER_32_68 ();
 sg13g2_decap_4 FILLER_32_75 ();
 sg13g2_fill_2 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_112 ();
 sg13g2_fill_2 FILLER_32_138 ();
 sg13g2_fill_2 FILLER_32_152 ();
 sg13g2_fill_1 FILLER_32_154 ();
 sg13g2_fill_1 FILLER_32_172 ();
 sg13g2_fill_2 FILLER_32_185 ();
 sg13g2_fill_2 FILLER_32_197 ();
 sg13g2_fill_1 FILLER_32_218 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_fill_2 FILLER_32_360 ();
 sg13g2_fill_2 FILLER_33_13 ();
 sg13g2_fill_1 FILLER_33_27 ();
 sg13g2_fill_2 FILLER_33_41 ();
 sg13g2_fill_1 FILLER_33_62 ();
 sg13g2_fill_1 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_fill_2 FILLER_33_135 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_188 ();
 sg13g2_fill_1 FILLER_33_194 ();
 sg13g2_fill_2 FILLER_33_228 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_288 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_fill_2 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_355 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_41 ();
 sg13g2_fill_1 FILLER_34_43 ();
 sg13g2_fill_2 FILLER_34_60 ();
 sg13g2_fill_1 FILLER_34_62 ();
 sg13g2_fill_1 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_108 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_fill_2 FILLER_34_142 ();
 sg13g2_fill_1 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_208 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_311 ();
 sg13g2_fill_2 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_fill_1 FILLER_34_393 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_28 ();
 sg13g2_fill_1 FILLER_35_30 ();
 sg13g2_fill_1 FILLER_35_39 ();
 sg13g2_fill_2 FILLER_35_57 ();
 sg13g2_fill_2 FILLER_35_82 ();
 sg13g2_fill_1 FILLER_35_84 ();
 sg13g2_fill_1 FILLER_35_90 ();
 sg13g2_fill_2 FILLER_35_130 ();
 sg13g2_fill_2 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_153 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_1 FILLER_35_177 ();
 sg13g2_fill_1 FILLER_35_211 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_238 ();
 sg13g2_fill_1 FILLER_35_251 ();
 sg13g2_fill_2 FILLER_35_280 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_2 FILLER_35_363 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_26 ();
 sg13g2_fill_2 FILLER_36_32 ();
 sg13g2_fill_1 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_156 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_fill_1 FILLER_36_191 ();
 sg13g2_fill_2 FILLER_36_209 ();
 sg13g2_fill_2 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_267 ();
 sg13g2_fill_1 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_286 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_11 ();
 sg13g2_fill_1 FILLER_37_41 ();
 sg13g2_fill_2 FILLER_37_57 ();
 sg13g2_fill_1 FILLER_37_59 ();
 sg13g2_fill_1 FILLER_37_71 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_237 ();
 sg13g2_fill_1 FILLER_37_239 ();
 sg13g2_fill_1 FILLER_37_284 ();
 sg13g2_fill_2 FILLER_37_307 ();
 sg13g2_fill_1 FILLER_37_309 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_fill_2 FILLER_37_365 ();
 sg13g2_fill_2 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_4 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_57 ();
 sg13g2_fill_2 FILLER_38_111 ();
 sg13g2_fill_1 FILLER_38_134 ();
 sg13g2_fill_2 FILLER_38_153 ();
 sg13g2_fill_1 FILLER_38_155 ();
 sg13g2_fill_1 FILLER_38_178 ();
 sg13g2_fill_2 FILLER_38_198 ();
 sg13g2_fill_1 FILLER_38_200 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_fill_1 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_337 ();
 sg13g2_fill_1 FILLER_38_339 ();
 sg13g2_fill_1 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_381 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net83;
 assign uio_oe[1] = net84;
 assign uio_oe[2] = net85;
 assign uio_oe[3] = net86;
 assign uio_oe[4] = net87;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
 assign uio_out[2] = net16;
 assign uio_out[3] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
endmodule
