module tt_um_wokwi_434917506576906241 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire params_ready;
 wire spike_out;
 wire \system_inst.leak_cycles[0] ;
 wire \system_inst.leak_cycles[1] ;
 wire \system_inst.leak_cycles[2] ;
 wire \system_inst.leak_cycles[3] ;
 wire \system_inst.leak_rate[0] ;
 wire \system_inst.leak_rate[1] ;
 wire \system_inst.leak_rate[2] ;
 wire \system_inst.leak_rate[3] ;
 wire \system_inst.leak_rate[4] ;
 wire \system_inst.leak_rate[5] ;
 wire \system_inst.leak_rate[6] ;
 wire \system_inst.leak_rate[7] ;
 wire \system_inst.loader.bit_count[0] ;
 wire \system_inst.loader.bit_count[1] ;
 wire \system_inst.loader.bit_count[2] ;
 wire \system_inst.loader.current_state[0] ;
 wire \system_inst.loader.current_state[1] ;
 wire \system_inst.loader.current_state[2] ;
 wire \system_inst.loader.current_state[3] ;
 wire \system_inst.loader.current_state[5] ;
 wire \system_inst.loader.shift_reg[0] ;
 wire \system_inst.loader.shift_reg[1] ;
 wire \system_inst.loader.shift_reg[2] ;
 wire \system_inst.loader.shift_reg[3] ;
 wire \system_inst.loader.shift_reg[4] ;
 wire \system_inst.loader.shift_reg[5] ;
 wire \system_inst.loader.shift_reg[6] ;
 wire \system_inst.loader.threshold_min[0] ;
 wire \system_inst.loader.threshold_min[1] ;
 wire \system_inst.loader.threshold_min[2] ;
 wire \system_inst.loader.threshold_min[3] ;
 wire \system_inst.loader.threshold_min[4] ;
 wire \system_inst.loader.threshold_min[5] ;
 wire \system_inst.loader.threshold_min[6] ;
 wire \system_inst.loader.threshold_min[7] ;
 wire \system_inst.loader.weight_a[0] ;
 wire \system_inst.loader.weight_a[1] ;
 wire \system_inst.loader.weight_a[2] ;
 wire \system_inst.neuron.leak_counter[0] ;
 wire \system_inst.neuron.leak_counter[1] ;
 wire \system_inst.neuron.leak_counter[2] ;
 wire \system_inst.neuron.leak_counter[3] ;
 wire \system_inst.neuron.refr_cnt[0] ;
 wire \system_inst.neuron.refr_cnt[1] ;
 wire \system_inst.neuron.refr_cnt[2] ;
 wire \system_inst.neuron.refr_cnt[3] ;
 wire \system_inst.neuron.threshold[0] ;
 wire \system_inst.neuron.threshold[1] ;
 wire \system_inst.neuron.threshold[2] ;
 wire \system_inst.neuron.threshold[3] ;
 wire \system_inst.neuron.threshold[4] ;
 wire \system_inst.neuron.threshold[5] ;
 wire \system_inst.neuron.threshold[6] ;
 wire \system_inst.neuron.threshold[7] ;
 wire \system_inst.neuron.v_mem[0] ;
 wire \system_inst.neuron.v_mem[1] ;
 wire \system_inst.neuron.v_mem[2] ;
 wire \system_inst.neuron.v_mem[3] ;
 wire \system_inst.neuron.v_mem[4] ;
 wire \system_inst.neuron.v_mem[5] ;
 wire \system_inst.neuron.v_mem[6] ;
 wire \system_inst.neuron.v_mem[7] ;
 wire \system_inst.neuron.v_mem[8] ;
 wire clknet_0_clk;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;

 sg13g2_inv_1 _0673_ (.Y(_0079_),
    .A(net96));
 sg13g2_inv_1 _0674_ (.Y(_0080_),
    .A(net182));
 sg13g2_inv_1 _0675_ (.Y(_0081_),
    .A(net108));
 sg13g2_inv_1 _0676_ (.Y(_0082_),
    .A(net179));
 sg13g2_inv_1 _0677_ (.Y(_0083_),
    .A(net128));
 sg13g2_inv_2 _0678_ (.Y(_0084_),
    .A(net126));
 sg13g2_inv_1 _0679_ (.Y(_0085_),
    .A(net104));
 sg13g2_inv_1 _0680_ (.Y(_0086_),
    .A(net116));
 sg13g2_inv_1 _0681_ (.Y(_0087_),
    .A(net98));
 sg13g2_inv_1 _0682_ (.Y(_0088_),
    .A(net4));
 sg13g2_inv_1 _0683_ (.Y(_0089_),
    .A(\system_inst.loader.threshold_min[6] ));
 sg13g2_inv_1 _0684_ (.Y(_0090_),
    .A(\system_inst.loader.threshold_min[5] ));
 sg13g2_inv_1 _0685_ (.Y(_0091_),
    .A(net203));
 sg13g2_inv_1 _0686_ (.Y(_0092_),
    .A(net206));
 sg13g2_inv_1 _0687_ (.Y(_0093_),
    .A(net198));
 sg13g2_inv_1 _0688_ (.Y(_0094_),
    .A(\system_inst.loader.threshold_min[0] ));
 sg13g2_inv_1 _0689_ (.Y(_0095_),
    .A(net187));
 sg13g2_inv_1 _0690_ (.Y(_0096_),
    .A(net158));
 sg13g2_inv_1 _0691_ (.Y(_0097_),
    .A(net212));
 sg13g2_inv_1 _0692_ (.Y(_0098_),
    .A(net221));
 sg13g2_inv_1 _0693_ (.Y(_0099_),
    .A(net192));
 sg13g2_inv_1 _0694_ (.Y(_0100_),
    .A(net210));
 sg13g2_inv_1 _0695_ (.Y(_0101_),
    .A(net217));
 sg13g2_inv_1 _0696_ (.Y(_0102_),
    .A(net205));
 sg13g2_inv_1 _0697_ (.Y(_0103_),
    .A(net161));
 sg13g2_inv_1 _0698_ (.Y(_0104_),
    .A(net162));
 sg13g2_inv_1 _0699_ (.Y(_0105_),
    .A(net207));
 sg13g2_inv_1 _0700_ (.Y(_0106_),
    .A(net107));
 sg13g2_inv_1 _0701_ (.Y(_0107_),
    .A(net173));
 sg13g2_inv_1 _0702_ (.Y(_0108_),
    .A(\system_inst.loader.current_state[0] ));
 sg13g2_inv_1 _0703_ (.Y(_0109_),
    .A(_0015_));
 sg13g2_nand2b_1 _0704_ (.Y(_0110_),
    .B(net173),
    .A_N(net1));
 sg13g2_nand2_1 _0705_ (.Y(_0111_),
    .A(net113),
    .B(\system_inst.loader.bit_count[0] ));
 sg13g2_nor2_1 _0706_ (.A(_0011_),
    .B(_0111_),
    .Y(_0112_));
 sg13g2_and2_2 _0707_ (.A(net1),
    .B(net3),
    .X(_0113_));
 sg13g2_nand2_1 _0708_ (.Y(_0114_),
    .A(net173),
    .B(_0113_));
 sg13g2_o21ai_1 _0709_ (.B1(_0110_),
    .Y(_0115_),
    .A1(net155),
    .A2(_0114_));
 sg13g2_and3_1 _0710_ (.X(_0116_),
    .A(\system_inst.loader.current_state[5] ),
    .B(_0112_),
    .C(_0113_));
 sg13g2_nand3_1 _0711_ (.B(net155),
    .C(_0113_),
    .A(\system_inst.loader.current_state[5] ),
    .Y(_0117_));
 sg13g2_a22oi_1 _0712_ (.Y(_0118_),
    .B1(net154),
    .B2(net174),
    .A2(_0115_),
    .A1(net107));
 sg13g2_inv_1 _0713_ (.Y(_0001_),
    .A(_0118_));
 sg13g2_and3_1 _0714_ (.X(_0119_),
    .A(\system_inst.loader.current_state[2] ),
    .B(_0112_),
    .C(_0113_));
 sg13g2_nand3_1 _0715_ (.B(net155),
    .C(_0113_),
    .A(net132),
    .Y(_0120_));
 sg13g2_a22oi_1 _0716_ (.Y(_0121_),
    .B1(net152),
    .B2(net173),
    .A2(_0115_),
    .A1(net133));
 sg13g2_inv_1 _0717_ (.Y(_0004_),
    .A(_0121_));
 sg13g2_nor2_1 _0718_ (.A(net118),
    .B(_0110_),
    .Y(_0122_));
 sg13g2_a21oi_1 _0719_ (.A1(net173),
    .A2(_0113_),
    .Y(_0000_),
    .B1(_0122_));
 sg13g2_nand3_1 _0720_ (.B(net155),
    .C(_0113_),
    .A(net101),
    .Y(_0123_));
 sg13g2_inv_1 _0721_ (.Y(_0124_),
    .A(_0123_));
 sg13g2_a22oi_1 _0722_ (.Y(_0125_),
    .B1(_0124_),
    .B2(net173),
    .A2(_0115_),
    .A1(net132));
 sg13g2_inv_1 _0723_ (.Y(_0002_),
    .A(_0125_));
 sg13g2_nand2_1 _0724_ (.Y(_0126_),
    .A(net101),
    .B(_0115_));
 sg13g2_o21ai_1 _0725_ (.B1(_0126_),
    .Y(_0003_),
    .A1(_0108_),
    .A2(_0114_));
 sg13g2_nor2b_1 _0726_ (.A(net163),
    .B_N(\system_inst.neuron.v_mem[0] ),
    .Y(uo_out[1]));
 sg13g2_nor2b_1 _0727_ (.A(net163),
    .B_N(\system_inst.neuron.v_mem[1] ),
    .Y(uo_out[2]));
 sg13g2_nor2b_1 _0728_ (.A(net163),
    .B_N(\system_inst.neuron.v_mem[2] ),
    .Y(uo_out[3]));
 sg13g2_nor2b_1 _0729_ (.A(\system_inst.neuron.v_mem[8] ),
    .B_N(\system_inst.neuron.v_mem[3] ),
    .Y(uo_out[4]));
 sg13g2_nor2b_1 _0730_ (.A(net163),
    .B_N(\system_inst.neuron.v_mem[4] ),
    .Y(uo_out[5]));
 sg13g2_nor2b_1 _0731_ (.A(net163),
    .B_N(\system_inst.neuron.v_mem[5] ),
    .Y(uo_out[6]));
 sg13g2_nor2b_1 _0732_ (.A(net163),
    .B_N(\system_inst.neuron.v_mem[6] ),
    .Y(uo_out[7]));
 sg13g2_nor2_1 _0733_ (.A(\system_inst.neuron.refr_cnt[1] ),
    .B(net208),
    .Y(_0127_));
 sg13g2_nor4_2 _0734_ (.A(\system_inst.neuron.refr_cnt[3] ),
    .B(\system_inst.neuron.refr_cnt[2] ),
    .C(\system_inst.neuron.refr_cnt[1] ),
    .Y(_0128_),
    .D(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_and2_2 _0735_ (.A(net124),
    .B(net1),
    .X(_0129_));
 sg13g2_nand2_1 _0736_ (.Y(_0130_),
    .A(net2),
    .B(_0129_));
 sg13g2_and3_2 _0737_ (.X(_0131_),
    .A(net2),
    .B(_0128_),
    .C(_0129_));
 sg13g2_nor2_1 _0738_ (.A(net166),
    .B(_0131_),
    .Y(_0132_));
 sg13g2_nand2_1 _0739_ (.Y(_0133_),
    .A(net91),
    .B(net150));
 sg13g2_and3_1 _0740_ (.X(_0134_),
    .A(net158),
    .B(\system_inst.neuron.v_mem[3] ),
    .C(net170));
 sg13g2_nand3_1 _0741_ (.B(\system_inst.neuron.v_mem[3] ),
    .C(net170),
    .A(\system_inst.loader.weight_a[2] ),
    .Y(_0135_));
 sg13g2_nand2_1 _0742_ (.Y(_0136_),
    .A(net159),
    .B(net7));
 sg13g2_a21oi_1 _0743_ (.A1(\system_inst.loader.weight_a[2] ),
    .A2(net170),
    .Y(_0137_),
    .B1(\system_inst.neuron.v_mem[3] ));
 sg13g2_nor2_1 _0744_ (.A(_0134_),
    .B(_0137_),
    .Y(_0138_));
 sg13g2_o21ai_1 _0745_ (.B1(_0135_),
    .Y(_0139_),
    .A1(_0136_),
    .A2(_0137_));
 sg13g2_nand2_1 _0746_ (.Y(_0140_),
    .A(net159),
    .B(net8));
 sg13g2_and3_1 _0747_ (.X(_0141_),
    .A(net158),
    .B(\system_inst.neuron.v_mem[4] ),
    .C(net7));
 sg13g2_nand3_1 _0748_ (.B(\system_inst.neuron.v_mem[4] ),
    .C(net7),
    .A(net158),
    .Y(_0142_));
 sg13g2_a21oi_1 _0749_ (.A1(net158),
    .A2(net7),
    .Y(_0143_),
    .B1(\system_inst.neuron.v_mem[4] ));
 sg13g2_nor2_1 _0750_ (.A(_0141_),
    .B(_0143_),
    .Y(_0144_));
 sg13g2_xnor2_1 _0751_ (.Y(_0145_),
    .A(_0140_),
    .B(_0144_));
 sg13g2_nand2_1 _0752_ (.Y(_0146_),
    .A(_0139_),
    .B(_0145_));
 sg13g2_nand2_1 _0753_ (.Y(_0147_),
    .A(net160),
    .B(net9));
 sg13g2_xnor2_1 _0754_ (.Y(_0148_),
    .A(_0139_),
    .B(_0145_));
 sg13g2_o21ai_1 _0755_ (.B1(_0146_),
    .Y(_0149_),
    .A1(_0147_),
    .A2(_0148_));
 sg13g2_nand2_1 _0756_ (.Y(_0150_),
    .A(net160),
    .B(net10));
 sg13g2_o21ai_1 _0757_ (.B1(_0142_),
    .Y(_0151_),
    .A1(_0140_),
    .A2(_0143_));
 sg13g2_nand2_1 _0758_ (.Y(_0152_),
    .A(net159),
    .B(net9));
 sg13g2_nand3_1 _0759_ (.B(\system_inst.neuron.v_mem[5] ),
    .C(net8),
    .A(net157),
    .Y(_0153_));
 sg13g2_a21o_1 _0760_ (.A2(net8),
    .A1(net157),
    .B1(\system_inst.neuron.v_mem[5] ),
    .X(_0154_));
 sg13g2_nand2_1 _0761_ (.Y(_0155_),
    .A(_0153_),
    .B(_0154_));
 sg13g2_xor2_1 _0762_ (.B(_0155_),
    .A(_0152_),
    .X(_0156_));
 sg13g2_nand2_1 _0763_ (.Y(_0157_),
    .A(_0151_),
    .B(_0156_));
 sg13g2_xnor2_1 _0764_ (.Y(_0158_),
    .A(_0151_),
    .B(_0156_));
 sg13g2_xor2_1 _0765_ (.B(_0158_),
    .A(_0150_),
    .X(_0159_));
 sg13g2_and2_1 _0766_ (.A(_0149_),
    .B(_0159_),
    .X(_0160_));
 sg13g2_nand3_1 _0767_ (.B(\system_inst.neuron.v_mem[2] ),
    .C(net5),
    .A(\system_inst.loader.weight_a[2] ),
    .Y(_0161_));
 sg13g2_nand2_1 _0768_ (.Y(_0162_),
    .A(net159),
    .B(net170));
 sg13g2_a21oi_1 _0769_ (.A1(net158),
    .A2(net5),
    .Y(_0163_),
    .B1(\system_inst.neuron.v_mem[2] ));
 sg13g2_a21o_1 _0770_ (.A2(net5),
    .A1(net158),
    .B1(\system_inst.neuron.v_mem[2] ),
    .X(_0164_));
 sg13g2_and4_1 _0771_ (.A(net159),
    .B(net170),
    .C(_0161_),
    .D(_0164_),
    .X(_0165_));
 sg13g2_o21ai_1 _0772_ (.B1(_0161_),
    .Y(_0166_),
    .A1(_0162_),
    .A2(_0163_));
 sg13g2_xnor2_1 _0773_ (.Y(_0167_),
    .A(_0136_),
    .B(_0138_));
 sg13g2_nand2_1 _0774_ (.Y(_0168_),
    .A(_0166_),
    .B(_0167_));
 sg13g2_nand2_1 _0775_ (.Y(_0169_),
    .A(net160),
    .B(net8));
 sg13g2_xnor2_1 _0776_ (.Y(_0170_),
    .A(_0166_),
    .B(_0167_));
 sg13g2_o21ai_1 _0777_ (.B1(_0168_),
    .Y(_0171_),
    .A1(_0169_),
    .A2(_0170_));
 sg13g2_xor2_1 _0778_ (.B(_0148_),
    .A(_0147_),
    .X(_0172_));
 sg13g2_nand2_1 _0779_ (.Y(_0173_),
    .A(_0171_),
    .B(_0172_));
 sg13g2_and2_1 _0780_ (.A(net159),
    .B(net5),
    .X(_0174_));
 sg13g2_nand2_2 _0781_ (.Y(_0175_),
    .A(\system_inst.neuron.v_mem[1] ),
    .B(_0174_));
 sg13g2_a22oi_1 _0782_ (.Y(_0176_),
    .B1(_0161_),
    .B2(_0164_),
    .A2(net170),
    .A1(net159));
 sg13g2_nor3_1 _0783_ (.A(_0165_),
    .B(_0175_),
    .C(_0176_),
    .Y(_0177_));
 sg13g2_or3_1 _0784_ (.A(_0165_),
    .B(_0175_),
    .C(_0176_),
    .X(_0178_));
 sg13g2_o21ai_1 _0785_ (.B1(_0175_),
    .Y(_0179_),
    .A1(_0165_),
    .A2(_0176_));
 sg13g2_and4_1 _0786_ (.A(net160),
    .B(net7),
    .C(_0178_),
    .D(_0179_),
    .X(_0180_));
 sg13g2_or2_1 _0787_ (.X(_0181_),
    .B(_0180_),
    .A(_0177_));
 sg13g2_xor2_1 _0788_ (.B(_0170_),
    .A(_0169_),
    .X(_0182_));
 sg13g2_and2_1 _0789_ (.A(_0181_),
    .B(_0182_),
    .X(_0183_));
 sg13g2_or2_1 _0790_ (.X(_0184_),
    .B(_0174_),
    .A(\system_inst.neuron.v_mem[1] ));
 sg13g2_and4_1 _0791_ (.A(net160),
    .B(net6),
    .C(_0175_),
    .D(_0184_),
    .X(_0185_));
 sg13g2_nand4_1 _0792_ (.B(net170),
    .C(_0175_),
    .A(net160),
    .Y(_0186_),
    .D(_0184_));
 sg13g2_a22oi_1 _0793_ (.Y(_0187_),
    .B1(_0178_),
    .B2(_0179_),
    .A2(net7),
    .A1(net160));
 sg13g2_nor3_1 _0794_ (.A(_0180_),
    .B(_0186_),
    .C(_0187_),
    .Y(_0188_));
 sg13g2_or3_1 _0795_ (.A(_0180_),
    .B(_0186_),
    .C(_0187_),
    .X(_0189_));
 sg13g2_nand2_1 _0796_ (.Y(_0190_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net5));
 sg13g2_or2_1 _0797_ (.X(_0191_),
    .B(_0190_),
    .A(_0005_));
 sg13g2_a22oi_1 _0798_ (.Y(_0192_),
    .B1(_0175_),
    .B2(_0184_),
    .A2(net170),
    .A1(net160));
 sg13g2_nor2_1 _0799_ (.A(_0185_),
    .B(_0192_),
    .Y(_0193_));
 sg13g2_nor3_1 _0800_ (.A(_0185_),
    .B(_0191_),
    .C(_0192_),
    .Y(_0194_));
 sg13g2_o21ai_1 _0801_ (.B1(_0186_),
    .Y(_0195_),
    .A1(_0180_),
    .A2(_0187_));
 sg13g2_nand3_1 _0802_ (.B(_0194_),
    .C(_0195_),
    .A(_0189_),
    .Y(_0196_));
 sg13g2_a21o_1 _0803_ (.A2(_0195_),
    .A1(_0194_),
    .B1(_0188_),
    .X(_0197_));
 sg13g2_xor2_1 _0804_ (.B(_0182_),
    .A(_0181_),
    .X(_0198_));
 sg13g2_a21oi_1 _0805_ (.A1(_0197_),
    .A2(_0198_),
    .Y(_0199_),
    .B1(_0183_));
 sg13g2_xnor2_1 _0806_ (.Y(_0200_),
    .A(_0171_),
    .B(_0172_));
 sg13g2_o21ai_1 _0807_ (.B1(_0173_),
    .Y(_0201_),
    .A1(_0199_),
    .A2(_0200_));
 sg13g2_xnor2_1 _0808_ (.Y(_0202_),
    .A(_0149_),
    .B(_0159_));
 sg13g2_inv_1 _0809_ (.Y(_0203_),
    .A(_0202_));
 sg13g2_a21oi_1 _0810_ (.A1(_0201_),
    .A2(_0203_),
    .Y(_0204_),
    .B1(_0160_));
 sg13g2_o21ai_1 _0811_ (.B1(_0157_),
    .Y(_0205_),
    .A1(_0150_),
    .A2(_0158_));
 sg13g2_o21ai_1 _0812_ (.B1(_0153_),
    .Y(_0206_),
    .A1(_0152_),
    .A2(_0155_));
 sg13g2_nand2_1 _0813_ (.Y(_0207_),
    .A(net159),
    .B(net10));
 sg13g2_and3_1 _0814_ (.X(_0208_),
    .A(net157),
    .B(\system_inst.neuron.v_mem[6] ),
    .C(net9));
 sg13g2_nand3_1 _0815_ (.B(\system_inst.neuron.v_mem[6] ),
    .C(net9),
    .A(net157),
    .Y(_0209_));
 sg13g2_a21oi_1 _0816_ (.A1(net157),
    .A2(net9),
    .Y(_0210_),
    .B1(\system_inst.neuron.v_mem[6] ));
 sg13g2_nor2_1 _0817_ (.A(_0208_),
    .B(_0210_),
    .Y(_0211_));
 sg13g2_xnor2_1 _0818_ (.Y(_0212_),
    .A(_0207_),
    .B(_0211_));
 sg13g2_nand2_1 _0819_ (.Y(_0213_),
    .A(_0206_),
    .B(_0212_));
 sg13g2_xnor2_1 _0820_ (.Y(_0214_),
    .A(_0206_),
    .B(_0212_));
 sg13g2_nand2b_1 _0821_ (.Y(_0215_),
    .B(_0205_),
    .A_N(_0214_));
 sg13g2_xor2_1 _0822_ (.B(_0214_),
    .A(_0205_),
    .X(_0216_));
 sg13g2_xnor2_1 _0823_ (.Y(_0217_),
    .A(_0204_),
    .B(_0216_));
 sg13g2_or2_1 _0824_ (.X(_0218_),
    .B(_0217_),
    .A(\system_inst.leak_rate[6] ));
 sg13g2_xnor2_1 _0825_ (.Y(_0219_),
    .A(_0201_),
    .B(_0203_));
 sg13g2_nor2_1 _0826_ (.A(\system_inst.leak_rate[5] ),
    .B(_0219_),
    .Y(_0220_));
 sg13g2_xnor2_1 _0827_ (.Y(_0221_),
    .A(_0199_),
    .B(_0200_));
 sg13g2_or2_1 _0828_ (.X(_0222_),
    .B(_0221_),
    .A(\system_inst.leak_rate[4] ));
 sg13g2_and2_1 _0829_ (.A(\system_inst.leak_rate[4] ),
    .B(_0221_),
    .X(_0223_));
 sg13g2_xor2_1 _0830_ (.B(_0221_),
    .A(\system_inst.leak_rate[4] ),
    .X(_0224_));
 sg13g2_xnor2_1 _0831_ (.Y(_0225_),
    .A(_0197_),
    .B(_0198_));
 sg13g2_nor2_1 _0832_ (.A(\system_inst.leak_rate[3] ),
    .B(_0225_),
    .Y(_0226_));
 sg13g2_a21o_1 _0833_ (.A2(_0195_),
    .A1(_0189_),
    .B1(_0194_),
    .X(_0227_));
 sg13g2_nand2_1 _0834_ (.Y(_0228_),
    .A(_0196_),
    .B(_0227_));
 sg13g2_nand3_1 _0835_ (.B(_0196_),
    .C(_0227_),
    .A(_0095_),
    .Y(_0229_));
 sg13g2_a21oi_1 _0836_ (.A1(_0196_),
    .A2(_0227_),
    .Y(_0230_),
    .B1(_0095_));
 sg13g2_xnor2_1 _0837_ (.Y(_0231_),
    .A(_0095_),
    .B(_0228_));
 sg13g2_xnor2_1 _0838_ (.Y(_0232_),
    .A(_0191_),
    .B(_0193_));
 sg13g2_nor2b_1 _0839_ (.A(\system_inst.leak_rate[1] ),
    .B_N(_0232_),
    .Y(_0233_));
 sg13g2_xor2_1 _0840_ (.B(_0190_),
    .A(_0005_),
    .X(_0234_));
 sg13g2_nand2b_1 _0841_ (.Y(_0235_),
    .B(\system_inst.leak_rate[0] ),
    .A_N(_0234_));
 sg13g2_xnor2_1 _0842_ (.Y(_0236_),
    .A(\system_inst.leak_rate[1] ),
    .B(_0232_));
 sg13g2_a21oi_1 _0843_ (.A1(_0235_),
    .A2(_0236_),
    .Y(_0237_),
    .B1(_0233_));
 sg13g2_o21ai_1 _0844_ (.B1(_0229_),
    .Y(_0238_),
    .A1(_0230_),
    .A2(_0237_));
 sg13g2_xor2_1 _0845_ (.B(_0225_),
    .A(\system_inst.leak_rate[3] ),
    .X(_0239_));
 sg13g2_a21oi_1 _0846_ (.A1(_0238_),
    .A2(_0239_),
    .Y(_0240_),
    .B1(_0226_));
 sg13g2_o21ai_1 _0847_ (.B1(_0222_),
    .Y(_0241_),
    .A1(_0223_),
    .A2(_0240_));
 sg13g2_xor2_1 _0848_ (.B(_0219_),
    .A(\system_inst.leak_rate[5] ),
    .X(_0242_));
 sg13g2_a21oi_1 _0849_ (.A1(_0241_),
    .A2(_0242_),
    .Y(_0243_),
    .B1(_0220_));
 sg13g2_xnor2_1 _0850_ (.Y(_0244_),
    .A(\system_inst.leak_rate[6] ),
    .B(_0217_));
 sg13g2_o21ai_1 _0851_ (.B1(_0218_),
    .Y(_0245_),
    .A1(_0243_),
    .A2(_0244_));
 sg13g2_o21ai_1 _0852_ (.B1(_0215_),
    .Y(_0246_),
    .A1(_0204_),
    .A2(_0216_));
 sg13g2_o21ai_1 _0853_ (.B1(_0209_),
    .Y(_0247_),
    .A1(_0207_),
    .A2(_0210_));
 sg13g2_inv_1 _0854_ (.Y(_0248_),
    .A(_0247_));
 sg13g2_and3_1 _0855_ (.X(_0249_),
    .A(net157),
    .B(\system_inst.neuron.v_mem[7] ),
    .C(net10));
 sg13g2_nand3_1 _0856_ (.B(\system_inst.neuron.v_mem[7] ),
    .C(net10),
    .A(net157),
    .Y(_0250_));
 sg13g2_a21oi_1 _0857_ (.A1(net157),
    .A2(net10),
    .Y(_0251_),
    .B1(\system_inst.neuron.v_mem[7] ));
 sg13g2_nor2_1 _0858_ (.A(_0249_),
    .B(_0251_),
    .Y(_0252_));
 sg13g2_xnor2_1 _0859_ (.Y(_0253_),
    .A(_0247_),
    .B(_0252_));
 sg13g2_nor2_1 _0860_ (.A(_0213_),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_xor2_1 _0861_ (.B(_0253_),
    .A(_0213_),
    .X(_0255_));
 sg13g2_xnor2_1 _0862_ (.Y(_0256_),
    .A(_0246_),
    .B(_0255_));
 sg13g2_xor2_1 _0863_ (.B(_0256_),
    .A(\system_inst.leak_rate[7] ),
    .X(_0257_));
 sg13g2_nand2b_1 _0864_ (.Y(_0258_),
    .B(\system_inst.leak_cycles[3] ),
    .A_N(\system_inst.neuron.leak_counter[3] ));
 sg13g2_nand2_1 _0865_ (.Y(_0259_),
    .A(_0085_),
    .B(\system_inst.neuron.leak_counter[3] ));
 sg13g2_nand2b_1 _0866_ (.Y(_0260_),
    .B(\system_inst.leak_cycles[1] ),
    .A_N(\system_inst.neuron.leak_counter[1] ));
 sg13g2_nand2b_1 _0867_ (.Y(_0261_),
    .B(\system_inst.neuron.leak_counter[1] ),
    .A_N(\system_inst.leak_cycles[1] ));
 sg13g2_nand3b_1 _0868_ (.B(_0261_),
    .C(\system_inst.leak_cycles[0] ),
    .Y(_0262_),
    .A_N(\system_inst.neuron.leak_counter[0] ));
 sg13g2_a22oi_1 _0869_ (.Y(_0263_),
    .B1(_0260_),
    .B2(_0262_),
    .A2(\system_inst.neuron.leak_counter[2] ),
    .A1(_0086_));
 sg13g2_o21ai_1 _0870_ (.B1(_0258_),
    .Y(_0264_),
    .A1(_0086_),
    .A2(\system_inst.neuron.leak_counter[2] ));
 sg13g2_o21ai_1 _0871_ (.B1(_0259_),
    .Y(_0265_),
    .A1(_0263_),
    .A2(_0264_));
 sg13g2_inv_1 _0872_ (.Y(_0266_),
    .A(_0265_));
 sg13g2_o21ai_1 _0873_ (.B1(_0265_),
    .Y(_0267_),
    .A1(\system_inst.leak_rate[7] ),
    .A2(_0256_));
 sg13g2_a21oi_1 _0874_ (.A1(_0245_),
    .A2(_0257_),
    .Y(_0268_),
    .B1(_0267_));
 sg13g2_a21oi_1 _0875_ (.A1(_0246_),
    .A2(_0255_),
    .Y(_0269_),
    .B1(_0254_));
 sg13g2_a21oi_1 _0876_ (.A1(_0248_),
    .A2(_0250_),
    .Y(_0270_),
    .B1(_0251_));
 sg13g2_xnor2_1 _0877_ (.Y(_0271_),
    .A(net163),
    .B(_0270_));
 sg13g2_xnor2_1 _0878_ (.Y(_0272_),
    .A(_0269_),
    .B(_0271_));
 sg13g2_xnor2_1 _0879_ (.Y(_0273_),
    .A(_0268_),
    .B(_0272_));
 sg13g2_nand2_1 _0880_ (.Y(_0274_),
    .A(_0217_),
    .B(net148));
 sg13g2_xnor2_1 _0881_ (.Y(_0275_),
    .A(_0243_),
    .B(_0244_));
 sg13g2_nand2_1 _0882_ (.Y(_0276_),
    .A(_0265_),
    .B(_0275_));
 sg13g2_nand3b_1 _0883_ (.B(_0274_),
    .C(_0276_),
    .Y(_0277_),
    .A_N(net142));
 sg13g2_xnor2_1 _0884_ (.Y(_0278_),
    .A(\system_inst.neuron.threshold[6] ),
    .B(_0277_));
 sg13g2_xor2_1 _0885_ (.B(_0257_),
    .A(_0245_),
    .X(_0279_));
 sg13g2_nand2_1 _0886_ (.Y(_0280_),
    .A(_0256_),
    .B(net148));
 sg13g2_o21ai_1 _0887_ (.B1(_0280_),
    .Y(_0281_),
    .A1(net148),
    .A2(_0279_));
 sg13g2_nor2_2 _0888_ (.A(net142),
    .B(_0281_),
    .Y(_0282_));
 sg13g2_or2_1 _0889_ (.X(_0283_),
    .B(_0282_),
    .A(_0006_));
 sg13g2_and2_1 _0890_ (.A(_0006_),
    .B(_0282_),
    .X(_0284_));
 sg13g2_xnor2_1 _0891_ (.Y(_0285_),
    .A(_0006_),
    .B(_0282_));
 sg13g2_nor2_1 _0892_ (.A(_0278_),
    .B(_0285_),
    .Y(_0286_));
 sg13g2_nand2_1 _0893_ (.Y(_0287_),
    .A(_0219_),
    .B(net148));
 sg13g2_xor2_1 _0894_ (.B(_0242_),
    .A(_0241_),
    .X(_0288_));
 sg13g2_o21ai_1 _0895_ (.B1(_0287_),
    .Y(_0289_),
    .A1(net148),
    .A2(_0288_));
 sg13g2_nor2_1 _0896_ (.A(net142),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_xnor2_1 _0897_ (.Y(_0291_),
    .A(_0008_),
    .B(_0290_));
 sg13g2_xnor2_1 _0898_ (.Y(_0292_),
    .A(_0224_),
    .B(_0240_));
 sg13g2_nor2_1 _0899_ (.A(net149),
    .B(_0292_),
    .Y(_0293_));
 sg13g2_a21oi_2 _0900_ (.B1(_0293_),
    .Y(_0294_),
    .A2(net148),
    .A1(_0221_));
 sg13g2_nand2b_2 _0901_ (.Y(_0295_),
    .B(_0294_),
    .A_N(net142));
 sg13g2_nand2_1 _0902_ (.Y(_0296_),
    .A(\system_inst.neuron.threshold[4] ),
    .B(_0295_));
 sg13g2_xnor2_1 _0903_ (.Y(_0297_),
    .A(\system_inst.neuron.threshold[4] ),
    .B(_0295_));
 sg13g2_nor4_1 _0904_ (.A(_0278_),
    .B(_0285_),
    .C(_0291_),
    .D(_0297_),
    .Y(_0298_));
 sg13g2_nand2_1 _0905_ (.Y(_0299_),
    .A(_0225_),
    .B(net149));
 sg13g2_xor2_1 _0906_ (.B(_0239_),
    .A(_0238_),
    .X(_0300_));
 sg13g2_o21ai_1 _0907_ (.B1(_0299_),
    .Y(_0301_),
    .A1(net149),
    .A2(_0300_));
 sg13g2_nor3_1 _0908_ (.A(\system_inst.neuron.threshold[3] ),
    .B(net141),
    .C(_0301_),
    .Y(_0302_));
 sg13g2_or3_1 _0909_ (.A(\system_inst.neuron.threshold[3] ),
    .B(net141),
    .C(_0301_),
    .X(_0303_));
 sg13g2_o21ai_1 _0910_ (.B1(net161),
    .Y(_0304_),
    .A1(net141),
    .A2(_0301_));
 sg13g2_xnor2_1 _0911_ (.Y(_0305_),
    .A(_0231_),
    .B(_0237_));
 sg13g2_nor2_1 _0912_ (.A(net149),
    .B(_0305_),
    .Y(_0306_));
 sg13g2_a21oi_1 _0913_ (.A1(_0228_),
    .A2(net149),
    .Y(_0307_),
    .B1(_0306_));
 sg13g2_inv_1 _0914_ (.Y(_0308_),
    .A(_0307_));
 sg13g2_or3_1 _0915_ (.A(\system_inst.neuron.threshold[2] ),
    .B(net141),
    .C(_0308_),
    .X(_0309_));
 sg13g2_o21ai_1 _0916_ (.B1(\system_inst.neuron.threshold[2] ),
    .Y(_0310_),
    .A1(net141),
    .A2(_0308_));
 sg13g2_nand4_1 _0917_ (.B(_0304_),
    .C(_0309_),
    .A(_0303_),
    .Y(_0311_),
    .D(_0310_));
 sg13g2_or2_1 _0918_ (.X(_0312_),
    .B(_0236_),
    .A(_0235_));
 sg13g2_a21oi_1 _0919_ (.A1(_0235_),
    .A2(_0236_),
    .Y(_0313_),
    .B1(net148));
 sg13g2_a22oi_1 _0920_ (.Y(_0314_),
    .B1(_0312_),
    .B2(_0313_),
    .A2(net148),
    .A1(_0232_));
 sg13g2_nor3_1 _0921_ (.A(\system_inst.neuron.threshold[1] ),
    .B(_0273_),
    .C(_0314_),
    .Y(_0315_));
 sg13g2_o21ai_1 _0922_ (.B1(\system_inst.neuron.threshold[1] ),
    .Y(_0316_),
    .A1(net142),
    .A2(_0314_));
 sg13g2_nand2_1 _0923_ (.Y(_0317_),
    .A(\system_inst.leak_rate[0] ),
    .B(_0265_));
 sg13g2_xor2_1 _0924_ (.B(_0317_),
    .A(_0234_),
    .X(_0318_));
 sg13g2_nor2_1 _0925_ (.A(_0273_),
    .B(_0318_),
    .Y(_0319_));
 sg13g2_nor3_1 _0926_ (.A(\system_inst.neuron.threshold[0] ),
    .B(_0273_),
    .C(_0318_),
    .Y(_0320_));
 sg13g2_a21o_1 _0927_ (.A2(_0320_),
    .A1(_0316_),
    .B1(_0315_),
    .X(_0321_));
 sg13g2_o21ai_1 _0928_ (.B1(_0105_),
    .Y(_0322_),
    .A1(net141),
    .A2(_0308_));
 sg13g2_a21o_1 _0929_ (.A2(_0322_),
    .A1(_0304_),
    .B1(_0302_),
    .X(_0323_));
 sg13g2_o21ai_1 _0930_ (.B1(_0323_),
    .Y(_0324_),
    .A1(_0311_),
    .A2(_0321_));
 sg13g2_o21ai_1 _0931_ (.B1(\system_inst.neuron.threshold[5] ),
    .Y(_0325_),
    .A1(net141),
    .A2(_0289_));
 sg13g2_o21ai_1 _0932_ (.B1(_0325_),
    .Y(_0326_),
    .A1(_0291_),
    .A2(_0296_));
 sg13g2_nand2b_1 _0933_ (.Y(_0327_),
    .B(_0277_),
    .A_N(_0007_));
 sg13g2_a21oi_1 _0934_ (.A1(_0283_),
    .A2(_0327_),
    .Y(_0328_),
    .B1(_0284_));
 sg13g2_a221oi_1 _0935_ (.B2(_0286_),
    .C1(_0328_),
    .B1(_0326_),
    .A1(_0298_),
    .Y(_0329_),
    .A2(_0324_));
 sg13g2_nor2b_1 _0936_ (.A(_0315_),
    .B_N(_0316_),
    .Y(_0330_));
 sg13g2_xnor2_1 _0937_ (.Y(_0331_),
    .A(_0010_),
    .B(_0319_));
 sg13g2_nor2_1 _0938_ (.A(_0311_),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_and3_1 _0939_ (.X(_0333_),
    .A(_0298_),
    .B(_0330_),
    .C(_0332_));
 sg13g2_nor2_2 _0940_ (.A(_0329_),
    .B(_0333_),
    .Y(_0334_));
 sg13g2_and2_1 _0941_ (.A(net171),
    .B(_0131_),
    .X(_0335_));
 sg13g2_nand2_2 _0942_ (.Y(_0336_),
    .A(net176),
    .B(_0131_));
 sg13g2_nand3_1 _0943_ (.B(net138),
    .C(_0335_),
    .A(_0319_),
    .Y(_0337_));
 sg13g2_nand2_1 _0944_ (.Y(_0019_),
    .A(_0133_),
    .B(_0337_));
 sg13g2_nor3_1 _0945_ (.A(net142),
    .B(_0314_),
    .C(_0336_),
    .Y(_0338_));
 sg13g2_a22oi_1 _0946_ (.Y(_0339_),
    .B1(net139),
    .B2(_0338_),
    .A2(net150),
    .A1(net190));
 sg13g2_inv_1 _0947_ (.Y(_0020_),
    .A(_0339_));
 sg13g2_nor3_1 _0948_ (.A(net141),
    .B(_0308_),
    .C(_0336_),
    .Y(_0340_));
 sg13g2_a22oi_1 _0949_ (.Y(_0341_),
    .B1(net139),
    .B2(_0340_),
    .A2(net150),
    .A1(net196));
 sg13g2_inv_1 _0950_ (.Y(_0021_),
    .A(_0341_));
 sg13g2_nor3_1 _0951_ (.A(net142),
    .B(_0301_),
    .C(_0336_),
    .Y(_0342_));
 sg13g2_a22oi_1 _0952_ (.Y(_0343_),
    .B1(net137),
    .B2(_0342_),
    .A2(net150),
    .A1(net200));
 sg13g2_inv_1 _0953_ (.Y(_0022_),
    .A(_0343_));
 sg13g2_nor2_1 _0954_ (.A(_0295_),
    .B(_0336_),
    .Y(_0344_));
 sg13g2_a22oi_1 _0955_ (.Y(_0345_),
    .B1(net137),
    .B2(_0344_),
    .A2(_0132_),
    .A1(net191));
 sg13g2_inv_1 _0956_ (.Y(_0023_),
    .A(_0345_));
 sg13g2_nand2_1 _0957_ (.Y(_0346_),
    .A(net103),
    .B(net150));
 sg13g2_nand3_1 _0958_ (.B(net137),
    .C(_0335_),
    .A(_0290_),
    .Y(_0347_));
 sg13g2_nand2_1 _0959_ (.Y(_0024_),
    .A(_0346_),
    .B(_0347_));
 sg13g2_nor2_1 _0960_ (.A(_0277_),
    .B(_0336_),
    .Y(_0348_));
 sg13g2_a22oi_1 _0961_ (.Y(_0349_),
    .B1(net137),
    .B2(_0348_),
    .A2(net150),
    .A1(net184));
 sg13g2_inv_1 _0962_ (.Y(_0025_),
    .A(_0349_));
 sg13g2_nand2_1 _0963_ (.Y(_0350_),
    .A(net106),
    .B(net150));
 sg13g2_nand3_1 _0964_ (.B(net138),
    .C(_0335_),
    .A(_0282_),
    .Y(_0351_));
 sg13g2_nand2_1 _0965_ (.Y(_0026_),
    .A(_0350_),
    .B(_0351_));
 sg13g2_and2_1 _0966_ (.A(net163),
    .B(_0132_),
    .X(_0027_));
 sg13g2_nor2_1 _0967_ (.A(net139),
    .B(_0336_),
    .Y(_0028_));
 sg13g2_nand2b_1 _0968_ (.Y(_0352_),
    .B(_0129_),
    .A_N(_0128_));
 sg13g2_o21ai_1 _0969_ (.B1(_0352_),
    .Y(_0353_),
    .A1(_0130_),
    .A2(_0334_));
 sg13g2_o21ai_1 _0970_ (.B1(_0353_),
    .Y(_0354_),
    .A1(net208),
    .A2(_0128_));
 sg13g2_o21ai_1 _0971_ (.B1(net175),
    .Y(_0355_),
    .A1(net208),
    .A2(_0353_));
 sg13g2_nor2b_1 _0972_ (.A(_0355_),
    .B_N(_0354_),
    .Y(_0029_));
 sg13g2_xnor2_1 _0973_ (.Y(_0356_),
    .A(\system_inst.neuron.refr_cnt[1] ),
    .B(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_nand2b_1 _0974_ (.Y(_0357_),
    .B(_0356_),
    .A_N(_0352_));
 sg13g2_o21ai_1 _0975_ (.B1(_0357_),
    .Y(_0358_),
    .A1(_0098_),
    .A2(_0353_));
 sg13g2_and2_1 _0976_ (.A(net175),
    .B(net222),
    .X(_0030_));
 sg13g2_nand3_1 _0977_ (.B(_0127_),
    .C(_0353_),
    .A(_0097_),
    .Y(_0359_));
 sg13g2_a21o_1 _0978_ (.A2(_0353_),
    .A1(_0127_),
    .B1(_0097_),
    .X(_0360_));
 sg13g2_a21oi_1 _0979_ (.A1(net213),
    .A2(_0360_),
    .Y(_0031_),
    .B1(net169));
 sg13g2_and3_1 _0980_ (.X(_0032_),
    .A(net94),
    .B(net175),
    .C(_0359_));
 sg13g2_nor2_1 _0981_ (.A(net167),
    .B(_0265_),
    .Y(_0361_));
 sg13g2_a21o_1 _0982_ (.A2(_0265_),
    .A1(_0129_),
    .B1(net168),
    .X(_0362_));
 sg13g2_xnor2_1 _0983_ (.Y(_0363_),
    .A(net189),
    .B(_0129_));
 sg13g2_nor2_1 _0984_ (.A(_0362_),
    .B(_0363_),
    .Y(_0033_));
 sg13g2_a21oi_1 _0985_ (.A1(\system_inst.neuron.leak_counter[0] ),
    .A2(_0129_),
    .Y(_0364_),
    .B1(net110));
 sg13g2_and3_1 _0986_ (.X(_0365_),
    .A(net110),
    .B(\system_inst.neuron.leak_counter[0] ),
    .C(_0129_));
 sg13g2_nor3_1 _0987_ (.A(_0362_),
    .B(net111),
    .C(_0365_),
    .Y(_0034_));
 sg13g2_nand2_1 _0988_ (.Y(_0366_),
    .A(\system_inst.neuron.leak_counter[2] ),
    .B(_0365_));
 sg13g2_xnor2_1 _0989_ (.Y(_0367_),
    .A(net185),
    .B(_0365_));
 sg13g2_nor2_1 _0990_ (.A(_0362_),
    .B(net186),
    .Y(_0035_));
 sg13g2_xor2_1 _0991_ (.B(_0366_),
    .A(net177),
    .X(_0368_));
 sg13g2_nor2_1 _0992_ (.A(_0362_),
    .B(net178),
    .Y(_0036_));
 sg13g2_nand2_1 _0993_ (.Y(_0369_),
    .A(net161),
    .B(net162));
 sg13g2_nand4_1 _0994_ (.B(\system_inst.neuron.threshold[4] ),
    .C(\system_inst.neuron.threshold[3] ),
    .A(\system_inst.neuron.threshold[5] ),
    .Y(_0370_),
    .D(net162));
 sg13g2_nor2_1 _0995_ (.A(_0007_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_xnor2_1 _0996_ (.Y(_0372_),
    .A(_0006_),
    .B(_0371_));
 sg13g2_nor2_1 _0997_ (.A(_0016_),
    .B(_0369_),
    .Y(_0373_));
 sg13g2_xor2_1 _0998_ (.B(_0373_),
    .A(_0008_),
    .X(_0374_));
 sg13g2_nor2_1 _0999_ (.A(_0109_),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_xor2_1 _1000_ (.B(net162),
    .A(net161),
    .X(_0376_));
 sg13g2_xnor2_1 _1001_ (.Y(_0377_),
    .A(_0016_),
    .B(_0369_));
 sg13g2_inv_1 _1002_ (.Y(_0378_),
    .A(_0377_));
 sg13g2_xnor2_1 _1003_ (.Y(_0379_),
    .A(_0017_),
    .B(_0377_));
 sg13g2_o21ai_1 _1004_ (.B1(_0379_),
    .Y(_0380_),
    .A1(_0018_),
    .A2(_0376_));
 sg13g2_xor2_1 _1005_ (.B(net162),
    .A(net156),
    .X(_0381_));
 sg13g2_o21ai_1 _1006_ (.B1(_0381_),
    .Y(_0382_),
    .A1(_0094_),
    .A2(\system_inst.neuron.threshold[1] ));
 sg13g2_and2_1 _1007_ (.A(_0018_),
    .B(_0376_),
    .X(_0383_));
 sg13g2_o21ai_1 _1008_ (.B1(_0382_),
    .Y(_0384_),
    .A1(net156),
    .A2(net162));
 sg13g2_nor2_1 _1009_ (.A(_0383_),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_xnor2_1 _1010_ (.Y(_0386_),
    .A(_0007_),
    .B(_0370_));
 sg13g2_nor2_1 _1011_ (.A(\system_inst.loader.threshold_min[5] ),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_a21oi_1 _1012_ (.A1(_0092_),
    .A2(_0378_),
    .Y(_0388_),
    .B1(_0387_));
 sg13g2_o21ai_1 _1013_ (.B1(_0388_),
    .Y(_0389_),
    .A1(_0380_),
    .A2(_0385_));
 sg13g2_xor2_1 _1014_ (.B(_0386_),
    .A(_0014_),
    .X(_0390_));
 sg13g2_a21oi_1 _1015_ (.A1(_0109_),
    .A2(_0374_),
    .Y(_0391_),
    .B1(_0390_));
 sg13g2_nor2b_1 _1016_ (.A(\system_inst.loader.threshold_min[0] ),
    .B_N(\system_inst.neuron.threshold[1] ),
    .Y(_0392_));
 sg13g2_nor4_1 _1017_ (.A(_0380_),
    .B(_0382_),
    .C(_0383_),
    .D(_0392_),
    .Y(_0393_));
 sg13g2_nand3_1 _1018_ (.B(_0391_),
    .C(_0393_),
    .A(_0010_),
    .Y(_0394_));
 sg13g2_a21oi_1 _1019_ (.A1(_0389_),
    .A2(_0394_),
    .Y(_0395_),
    .B1(_0375_));
 sg13g2_nor2_1 _1020_ (.A(_0387_),
    .B(_0391_),
    .Y(_0396_));
 sg13g2_nor2_1 _1021_ (.A(_0013_),
    .B(_0372_),
    .Y(_0397_));
 sg13g2_nor3_1 _1022_ (.A(_0395_),
    .B(_0396_),
    .C(_0397_),
    .Y(_0398_));
 sg13g2_nor2_1 _1023_ (.A(_0372_),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_a21o_1 _1024_ (.A2(_0372_),
    .A1(_0013_),
    .B1(_0398_),
    .X(_0400_));
 sg13g2_nand2_1 _1025_ (.Y(_0401_),
    .A(net156),
    .B(net146));
 sg13g2_o21ai_1 _1026_ (.B1(_0401_),
    .Y(_0402_),
    .A1(_0105_),
    .A2(net146));
 sg13g2_nand2_1 _1027_ (.Y(_0403_),
    .A(net156),
    .B(\system_inst.loader.threshold_min[0] ));
 sg13g2_nand4_1 _1028_ (.B(\system_inst.loader.threshold_min[2] ),
    .C(net156),
    .A(\system_inst.loader.threshold_min[3] ),
    .Y(_0404_),
    .D(\system_inst.loader.threshold_min[0] ));
 sg13g2_nor3_2 _1029_ (.A(_0090_),
    .B(_0091_),
    .C(_0404_),
    .Y(_0405_));
 sg13g2_nand2_1 _1030_ (.Y(_0406_),
    .A(\system_inst.loader.threshold_min[6] ),
    .B(_0405_));
 sg13g2_xor2_1 _1031_ (.B(_0406_),
    .A(\system_inst.loader.threshold_min[7] ),
    .X(_0407_));
 sg13g2_nand2b_1 _1032_ (.Y(_0408_),
    .B(_0006_),
    .A_N(_0407_));
 sg13g2_xnor2_1 _1033_ (.Y(_0409_),
    .A(_0013_),
    .B(_0405_));
 sg13g2_nor2_1 _1034_ (.A(_0015_),
    .B(_0404_),
    .Y(_0410_));
 sg13g2_xnor2_1 _1035_ (.Y(_0411_),
    .A(_0014_),
    .B(_0410_));
 sg13g2_nand2_1 _1036_ (.Y(_0412_),
    .A(_0101_),
    .B(_0411_));
 sg13g2_nor2_1 _1037_ (.A(_0018_),
    .B(_0403_),
    .Y(_0413_));
 sg13g2_xor2_1 _1038_ (.B(_0413_),
    .A(_0017_),
    .X(_0414_));
 sg13g2_or2_2 _1039_ (.X(_0415_),
    .B(\system_inst.neuron.threshold[0] ),
    .A(\system_inst.neuron.threshold[1] ));
 sg13g2_nand2_1 _1040_ (.Y(_0416_),
    .A(\system_inst.neuron.threshold[1] ),
    .B(\system_inst.neuron.threshold[0] ));
 sg13g2_nor2b_1 _1041_ (.A(_0392_),
    .B_N(_0416_),
    .Y(_0417_));
 sg13g2_o21ai_1 _1042_ (.B1(_0403_),
    .Y(_0418_),
    .A1(net156),
    .A2(_0417_));
 sg13g2_nand2_1 _1043_ (.Y(_0419_),
    .A(_0415_),
    .B(_0418_));
 sg13g2_xor2_1 _1044_ (.B(_0403_),
    .A(_0018_),
    .X(_0420_));
 sg13g2_xnor2_1 _1045_ (.Y(_0421_),
    .A(_0105_),
    .B(_0420_));
 sg13g2_a22oi_1 _1046_ (.Y(_0422_),
    .B1(_0421_),
    .B2(_0419_),
    .A2(_0420_),
    .A1(_0104_));
 sg13g2_a21o_1 _1047_ (.A2(_0414_),
    .A1(net161),
    .B1(_0422_),
    .X(_0423_));
 sg13g2_xnor2_1 _1048_ (.Y(_0424_),
    .A(_0109_),
    .B(_0404_));
 sg13g2_o21ai_1 _1049_ (.B1(_0423_),
    .Y(_0425_),
    .A1(net161),
    .A2(_0414_));
 sg13g2_a21oi_1 _1050_ (.A1(_0016_),
    .A2(_0424_),
    .Y(_0426_),
    .B1(_0425_));
 sg13g2_xor2_1 _1051_ (.B(_0411_),
    .A(_0008_),
    .X(_0427_));
 sg13g2_o21ai_1 _1052_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0016_),
    .A2(_0424_));
 sg13g2_o21ai_1 _1053_ (.B1(_0412_),
    .Y(_0429_),
    .A1(_0426_),
    .A2(_0428_));
 sg13g2_xor2_1 _1054_ (.B(_0409_),
    .A(_0007_),
    .X(_0430_));
 sg13g2_a22oi_1 _1055_ (.Y(_0431_),
    .B1(_0429_),
    .B2(_0430_),
    .A2(_0409_),
    .A1(_0100_));
 sg13g2_xnor2_1 _1056_ (.Y(_0432_),
    .A(\system_inst.neuron.threshold[7] ),
    .B(_0407_));
 sg13g2_o21ai_1 _1057_ (.B1(_0408_),
    .Y(_0433_),
    .A1(_0431_),
    .A2(_0432_));
 sg13g2_nor2_1 _1058_ (.A(net162),
    .B(_0415_),
    .Y(_0434_));
 sg13g2_xnor2_1 _1059_ (.Y(_0435_),
    .A(_0104_),
    .B(_0415_));
 sg13g2_nor2_1 _1060_ (.A(net144),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_a21oi_1 _1061_ (.A1(net198),
    .A2(net144),
    .Y(_0437_),
    .B1(_0436_));
 sg13g2_a21oi_1 _1062_ (.A1(net138),
    .A2(_0437_),
    .Y(_0438_),
    .B1(net165));
 sg13g2_o21ai_1 _1063_ (.B1(_0438_),
    .Y(_0439_),
    .A1(net138),
    .A2(_0402_));
 sg13g2_a21o_1 _1064_ (.A2(_0361_),
    .A1(net139),
    .B1(net150),
    .X(_0440_));
 sg13g2_a21oi_1 _1065_ (.A1(net198),
    .A2(net165),
    .Y(_0441_),
    .B1(net135));
 sg13g2_a22oi_1 _1066_ (.Y(_0037_),
    .B1(_0441_),
    .B2(_0439_),
    .A2(net135),
    .A1(_0104_));
 sg13g2_nor2_1 _1067_ (.A(_0376_),
    .B(net146),
    .Y(_0442_));
 sg13g2_a21oi_1 _1068_ (.A1(_0093_),
    .A2(net146),
    .Y(_0443_),
    .B1(_0442_));
 sg13g2_nor3_2 _1069_ (.A(net161),
    .B(net162),
    .C(_0415_),
    .Y(_0444_));
 sg13g2_xnor2_1 _1070_ (.Y(_0445_),
    .A(net161),
    .B(_0434_));
 sg13g2_nor2_1 _1071_ (.A(net144),
    .B(_0445_),
    .Y(_0446_));
 sg13g2_a21oi_1 _1072_ (.A1(net206),
    .A2(net144),
    .Y(_0447_),
    .B1(_0446_));
 sg13g2_a21oi_1 _1073_ (.A1(net136),
    .A2(_0447_),
    .Y(_0448_),
    .B1(net164));
 sg13g2_o21ai_1 _1074_ (.B1(_0448_),
    .Y(_0449_),
    .A1(net136),
    .A2(_0443_));
 sg13g2_a21oi_1 _1075_ (.A1(net206),
    .A2(net164),
    .Y(_0450_),
    .B1(net134));
 sg13g2_a22oi_1 _1076_ (.Y(_0038_),
    .B1(_0449_),
    .B2(_0450_),
    .A2(net134),
    .A1(_0103_));
 sg13g2_nor2_1 _1077_ (.A(_0377_),
    .B(net145),
    .Y(_0451_));
 sg13g2_a21oi_1 _1078_ (.A1(\system_inst.loader.threshold_min[3] ),
    .A2(net145),
    .Y(_0452_),
    .B1(_0451_));
 sg13g2_o21ai_1 _1079_ (.B1(_0452_),
    .Y(_0453_),
    .A1(_0329_),
    .A2(_0333_));
 sg13g2_and2_1 _1080_ (.A(_0102_),
    .B(_0444_),
    .X(_0454_));
 sg13g2_xnor2_1 _1081_ (.Y(_0455_),
    .A(\system_inst.neuron.threshold[4] ),
    .B(_0444_));
 sg13g2_nor2_1 _1082_ (.A(net143),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_a21oi_1 _1083_ (.A1(\system_inst.loader.threshold_min[4] ),
    .A2(net143),
    .Y(_0457_),
    .B1(_0456_));
 sg13g2_a21oi_1 _1084_ (.A1(net136),
    .A2(_0457_),
    .Y(_0458_),
    .B1(net164));
 sg13g2_a221oi_1 _1085_ (.B2(_0458_),
    .C1(net135),
    .B1(_0453_),
    .A1(net203),
    .Y(_0459_),
    .A2(net164));
 sg13g2_a21oi_1 _1086_ (.A1(_0102_),
    .A2(net134),
    .Y(_0039_),
    .B1(_0459_));
 sg13g2_nand2_1 _1087_ (.Y(_0460_),
    .A(net203),
    .B(net145));
 sg13g2_o21ai_1 _1088_ (.B1(_0460_),
    .Y(_0461_),
    .A1(_0374_),
    .A2(net145));
 sg13g2_and2_1 _1089_ (.A(_0101_),
    .B(_0454_),
    .X(_0462_));
 sg13g2_xnor2_1 _1090_ (.Y(_0463_),
    .A(\system_inst.neuron.threshold[5] ),
    .B(_0454_));
 sg13g2_nor2_1 _1091_ (.A(net143),
    .B(_0463_),
    .Y(_0464_));
 sg13g2_a21oi_1 _1092_ (.A1(\system_inst.loader.threshold_min[5] ),
    .A2(net143),
    .Y(_0465_),
    .B1(_0464_));
 sg13g2_a21oi_1 _1093_ (.A1(net136),
    .A2(_0465_),
    .Y(_0466_),
    .B1(net164));
 sg13g2_o21ai_1 _1094_ (.B1(_0466_),
    .Y(_0467_),
    .A1(net136),
    .A2(_0461_));
 sg13g2_a21oi_1 _1095_ (.A1(net202),
    .A2(net164),
    .Y(_0468_),
    .B1(net134));
 sg13g2_a22oi_1 _1096_ (.Y(_0040_),
    .B1(_0467_),
    .B2(_0468_),
    .A2(net135),
    .A1(_0101_));
 sg13g2_nand2_1 _1097_ (.Y(_0469_),
    .A(\system_inst.loader.threshold_min[5] ),
    .B(net145));
 sg13g2_o21ai_1 _1098_ (.B1(_0469_),
    .Y(_0470_),
    .A1(_0386_),
    .A2(net145));
 sg13g2_and2_1 _1099_ (.A(_0100_),
    .B(_0462_),
    .X(_0471_));
 sg13g2_xnor2_1 _1100_ (.Y(_0472_),
    .A(\system_inst.neuron.threshold[6] ),
    .B(_0462_));
 sg13g2_nor2_1 _1101_ (.A(net143),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_a21oi_1 _1102_ (.A1(net204),
    .A2(net143),
    .Y(_0474_),
    .B1(_0473_));
 sg13g2_a21oi_1 _1103_ (.A1(net136),
    .A2(_0474_),
    .Y(_0475_),
    .B1(net166));
 sg13g2_o21ai_1 _1104_ (.B1(_0475_),
    .Y(_0476_),
    .A1(net136),
    .A2(_0470_));
 sg13g2_a21oi_1 _1105_ (.A1(net204),
    .A2(net166),
    .Y(_0477_),
    .B1(net134));
 sg13g2_a22oi_1 _1106_ (.Y(_0041_),
    .B1(_0476_),
    .B2(_0477_),
    .A2(net134),
    .A1(_0100_));
 sg13g2_xnor2_1 _1107_ (.Y(_0478_),
    .A(\system_inst.neuron.threshold[7] ),
    .B(_0471_));
 sg13g2_nor2_1 _1108_ (.A(net143),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_a21oi_1 _1109_ (.A1(\system_inst.loader.threshold_min[7] ),
    .A2(net143),
    .Y(_0480_),
    .B1(_0479_));
 sg13g2_a21oi_1 _1110_ (.A1(_0089_),
    .A2(net145),
    .Y(_0481_),
    .B1(_0399_));
 sg13g2_a21oi_1 _1111_ (.A1(net137),
    .A2(_0480_),
    .Y(_0482_),
    .B1(net166));
 sg13g2_o21ai_1 _1112_ (.B1(_0482_),
    .Y(_0483_),
    .A1(net136),
    .A2(_0481_));
 sg13g2_a21oi_1 _1113_ (.A1(\system_inst.loader.threshold_min[7] ),
    .A2(net166),
    .Y(_0484_),
    .B1(net134));
 sg13g2_a22oi_1 _1114_ (.Y(_0042_),
    .B1(_0483_),
    .B2(_0484_),
    .A2(net134),
    .A1(_0099_));
 sg13g2_nor3_1 _1115_ (.A(net166),
    .B(net138),
    .C(net146),
    .Y(_0485_));
 sg13g2_or2_1 _1116_ (.X(_0486_),
    .B(_0485_),
    .A(net135));
 sg13g2_nor2_1 _1117_ (.A(net166),
    .B(net144),
    .Y(_0487_));
 sg13g2_mux2_1 _1118_ (.A0(\system_inst.loader.threshold_min[0] ),
    .A1(_0010_),
    .S(_0487_),
    .X(_0488_));
 sg13g2_o21ai_1 _1119_ (.B1(_0488_),
    .Y(_0489_),
    .A1(net166),
    .A2(net138));
 sg13g2_o21ai_1 _1120_ (.B1(net130),
    .Y(_0490_),
    .A1(net135),
    .A2(_0485_));
 sg13g2_o21ai_1 _1121_ (.B1(_0490_),
    .Y(_0043_),
    .A1(_0486_),
    .A2(_0489_));
 sg13g2_a21oi_1 _1122_ (.A1(\system_inst.loader.threshold_min[0] ),
    .A2(net145),
    .Y(_0491_),
    .B1(net138));
 sg13g2_a21oi_1 _1123_ (.A1(_0415_),
    .A2(_0416_),
    .Y(_0492_),
    .B1(net144));
 sg13g2_a21oi_1 _1124_ (.A1(net156),
    .A2(net144),
    .Y(_0493_),
    .B1(_0492_));
 sg13g2_a21o_1 _1125_ (.A2(_0493_),
    .A1(net138),
    .B1(net165),
    .X(_0494_));
 sg13g2_nand2_1 _1126_ (.Y(_0495_),
    .A(net156),
    .B(net165));
 sg13g2_o21ai_1 _1127_ (.B1(_0495_),
    .Y(_0496_),
    .A1(_0491_),
    .A2(_0494_));
 sg13g2_mux2_1 _1128_ (.A0(_0496_),
    .A1(net215),
    .S(_0486_),
    .X(_0044_));
 sg13g2_nor3_2 _1129_ (.A(\system_inst.loader.current_state[2] ),
    .B(\system_inst.loader.current_state[5] ),
    .C(\system_inst.loader.current_state[3] ),
    .Y(_0497_));
 sg13g2_nand2_1 _1130_ (.Y(_0498_),
    .A(_0012_),
    .B(_0497_));
 sg13g2_nor2_1 _1131_ (.A(net118),
    .B(_0498_),
    .Y(_0499_));
 sg13g2_o21ai_1 _1132_ (.B1(net1),
    .Y(_0500_),
    .A1(net3),
    .A2(_0108_));
 sg13g2_nor2_1 _1133_ (.A(_0499_),
    .B(_0500_),
    .Y(_0501_));
 sg13g2_o21ai_1 _1134_ (.B1(_0497_),
    .Y(_0502_),
    .A1(_0012_),
    .A2(net155));
 sg13g2_nand2_1 _1135_ (.Y(_0503_),
    .A(net3),
    .B(_0502_));
 sg13g2_nand2_1 _1136_ (.Y(_0504_),
    .A(_0501_),
    .B(_0503_));
 sg13g2_and2_1 _1137_ (.A(_0106_),
    .B(_0497_),
    .X(_0505_));
 sg13g2_a21oi_1 _1138_ (.A1(net124),
    .A2(_0504_),
    .Y(_0506_),
    .B1(net168));
 sg13g2_o21ai_1 _1139_ (.B1(_0506_),
    .Y(_0045_),
    .A1(_0504_),
    .A2(_0505_));
 sg13g2_o21ai_1 _1140_ (.B1(net174),
    .Y(_0507_),
    .A1(net201),
    .A2(_0124_));
 sg13g2_a21oi_1 _1141_ (.A1(_0088_),
    .A2(_0124_),
    .Y(_0046_),
    .B1(_0507_));
 sg13g2_a21oi_1 _1142_ (.A1(net122),
    .A2(_0123_),
    .Y(_0508_),
    .B1(net168));
 sg13g2_o21ai_1 _1143_ (.B1(_0508_),
    .Y(_0047_),
    .A1(_0084_),
    .A2(_0123_));
 sg13g2_o21ai_1 _1144_ (.B1(net175),
    .Y(_0509_),
    .A1(net211),
    .A2(_0123_));
 sg13g2_a21oi_1 _1145_ (.A1(_0096_),
    .A2(_0123_),
    .Y(_0048_),
    .B1(_0509_));
 sg13g2_o21ai_1 _1146_ (.B1(net174),
    .Y(_0510_),
    .A1(net183),
    .A2(net152));
 sg13g2_a21oi_1 _1147_ (.A1(_0088_),
    .A2(net152),
    .Y(_0049_),
    .B1(_0510_));
 sg13g2_a21oi_1 _1148_ (.A1(net197),
    .A2(_0120_),
    .Y(_0511_),
    .B1(net169));
 sg13g2_o21ai_1 _1149_ (.B1(_0511_),
    .Y(_0050_),
    .A1(_0084_),
    .A2(_0120_));
 sg13g2_o21ai_1 _1150_ (.B1(net175),
    .Y(_0512_),
    .A1(\system_inst.loader.shift_reg[1] ),
    .A2(_0120_));
 sg13g2_a21oi_1 _1151_ (.A1(_0095_),
    .A2(_0120_),
    .Y(_0051_),
    .B1(_0512_));
 sg13g2_o21ai_1 _1152_ (.B1(net172),
    .Y(_0513_),
    .A1(\system_inst.leak_rate[3] ),
    .A2(net151));
 sg13g2_a21oi_1 _1153_ (.A1(_0083_),
    .A2(net151),
    .Y(_0052_),
    .B1(_0513_));
 sg13g2_o21ai_1 _1154_ (.B1(net174),
    .Y(_0514_),
    .A1(\system_inst.leak_rate[4] ),
    .A2(net152));
 sg13g2_a21oi_1 _1155_ (.A1(_0082_),
    .A2(net152),
    .Y(_0053_),
    .B1(_0514_));
 sg13g2_o21ai_1 _1156_ (.B1(net171),
    .Y(_0515_),
    .A1(net195),
    .A2(net151));
 sg13g2_a21oi_1 _1157_ (.A1(_0081_),
    .A2(net151),
    .Y(_0054_),
    .B1(_0515_));
 sg13g2_o21ai_1 _1158_ (.B1(net171),
    .Y(_0516_),
    .A1(net194),
    .A2(net151));
 sg13g2_a21oi_1 _1159_ (.A1(_0080_),
    .A2(net151),
    .Y(_0055_),
    .B1(_0516_));
 sg13g2_o21ai_1 _1160_ (.B1(net176),
    .Y(_0517_),
    .A1(net115),
    .A2(net151));
 sg13g2_a21oi_1 _1161_ (.A1(_0079_),
    .A2(net151),
    .Y(_0056_),
    .B1(_0517_));
 sg13g2_o21ai_1 _1162_ (.B1(net174),
    .Y(_0518_),
    .A1(net220),
    .A2(net154));
 sg13g2_a21oi_1 _1163_ (.A1(_0088_),
    .A2(net153),
    .Y(_0057_),
    .B1(_0518_));
 sg13g2_a21oi_1 _1164_ (.A1(net119),
    .A2(_0117_),
    .Y(_0519_),
    .B1(net168));
 sg13g2_o21ai_1 _1165_ (.B1(net120),
    .Y(_0058_),
    .A1(_0084_),
    .A2(_0117_));
 sg13g2_a21oi_1 _1166_ (.A1(\system_inst.loader.shift_reg[1] ),
    .A2(net154),
    .Y(_0520_),
    .B1(net168));
 sg13g2_o21ai_1 _1167_ (.B1(_0520_),
    .Y(_0059_),
    .A1(_0093_),
    .A2(net153));
 sg13g2_a21oi_1 _1168_ (.A1(net128),
    .A2(net154),
    .Y(_0521_),
    .B1(net164));
 sg13g2_o21ai_1 _1169_ (.B1(_0521_),
    .Y(_0060_),
    .A1(_0092_),
    .A2(net153));
 sg13g2_a21oi_1 _1170_ (.A1(net179),
    .A2(net154),
    .Y(_0522_),
    .B1(net164));
 sg13g2_o21ai_1 _1171_ (.B1(_0522_),
    .Y(_0061_),
    .A1(_0091_),
    .A2(net153));
 sg13g2_o21ai_1 _1172_ (.B1(net171),
    .Y(_0523_),
    .A1(net202),
    .A2(net153));
 sg13g2_a21oi_1 _1173_ (.A1(_0081_),
    .A2(net153),
    .Y(_0062_),
    .B1(_0523_));
 sg13g2_o21ai_1 _1174_ (.B1(net171),
    .Y(_0524_),
    .A1(net204),
    .A2(net153));
 sg13g2_a21oi_1 _1175_ (.A1(_0080_),
    .A2(net153),
    .Y(_0063_),
    .B1(_0524_));
 sg13g2_o21ai_1 _1176_ (.B1(net171),
    .Y(_0525_),
    .A1(\system_inst.loader.threshold_min[7] ),
    .A2(net154));
 sg13g2_a21oi_1 _1177_ (.A1(_0079_),
    .A2(net154),
    .Y(_0064_),
    .B1(_0525_));
 sg13g2_nand3_1 _1178_ (.B(net155),
    .C(_0113_),
    .A(net107),
    .Y(_0526_));
 sg13g2_o21ai_1 _1179_ (.B1(net173),
    .Y(_0527_),
    .A1(net4),
    .A2(_0526_));
 sg13g2_a21oi_1 _1180_ (.A1(_0087_),
    .A2(_0526_),
    .Y(_0065_),
    .B1(_0527_));
 sg13g2_a21oi_1 _1181_ (.A1(net181),
    .A2(_0526_),
    .Y(_0528_),
    .B1(net168));
 sg13g2_o21ai_1 _1182_ (.B1(_0528_),
    .Y(_0066_),
    .A1(_0084_),
    .A2(_0526_));
 sg13g2_o21ai_1 _1183_ (.B1(net172),
    .Y(_0529_),
    .A1(\system_inst.loader.shift_reg[1] ),
    .A2(_0526_));
 sg13g2_a21oi_1 _1184_ (.A1(_0086_),
    .A2(_0526_),
    .Y(_0067_),
    .B1(_0529_));
 sg13g2_o21ai_1 _1185_ (.B1(net172),
    .Y(_0530_),
    .A1(\system_inst.loader.shift_reg[2] ),
    .A2(_0526_));
 sg13g2_a21oi_1 _1186_ (.A1(_0085_),
    .A2(_0526_),
    .Y(_0068_),
    .B1(_0530_));
 sg13g2_nor2_1 _1187_ (.A(net3),
    .B(_0505_),
    .Y(_0531_));
 sg13g2_nor2b_2 _1188_ (.A(_0531_),
    .B_N(_0501_),
    .Y(_0532_));
 sg13g2_nand2b_1 _1189_ (.Y(_0533_),
    .B(_0501_),
    .A_N(_0531_));
 sg13g2_a21oi_2 _1190_ (.B1(_0505_),
    .Y(_0534_),
    .A2(net155),
    .A1(_0106_));
 sg13g2_a21oi_1 _1191_ (.A1(net4),
    .A2(_0534_),
    .Y(_0535_),
    .B1(_0533_));
 sg13g2_o21ai_1 _1192_ (.B1(net172),
    .Y(_0536_),
    .A1(net126),
    .A2(_0532_));
 sg13g2_nor2_1 _1193_ (.A(_0535_),
    .B(_0536_),
    .Y(_0069_));
 sg13g2_a21oi_1 _1194_ (.A1(net126),
    .A2(_0534_),
    .Y(_0537_),
    .B1(net147));
 sg13g2_o21ai_1 _1195_ (.B1(net172),
    .Y(_0538_),
    .A1(\system_inst.loader.shift_reg[1] ),
    .A2(_0532_));
 sg13g2_nor2_1 _1196_ (.A(_0537_),
    .B(_0538_),
    .Y(_0070_));
 sg13g2_a21oi_1 _1197_ (.A1(net211),
    .A2(_0534_),
    .Y(_0539_),
    .B1(net147));
 sg13g2_o21ai_1 _1198_ (.B1(net172),
    .Y(_0540_),
    .A1(net128),
    .A2(_0532_));
 sg13g2_nor2_1 _1199_ (.A(_0539_),
    .B(_0540_),
    .Y(_0071_));
 sg13g2_a21oi_1 _1200_ (.A1(net128),
    .A2(_0534_),
    .Y(_0541_),
    .B1(net147));
 sg13g2_o21ai_1 _1201_ (.B1(net172),
    .Y(_0542_),
    .A1(net179),
    .A2(_0532_));
 sg13g2_nor2_1 _1202_ (.A(_0541_),
    .B(_0542_),
    .Y(_0072_));
 sg13g2_a21oi_1 _1203_ (.A1(net179),
    .A2(_0534_),
    .Y(_0543_),
    .B1(net147));
 sg13g2_o21ai_1 _1204_ (.B1(net171),
    .Y(_0544_),
    .A1(net108),
    .A2(_0532_));
 sg13g2_nor2_1 _1205_ (.A(_0543_),
    .B(_0544_),
    .Y(_0073_));
 sg13g2_a21oi_1 _1206_ (.A1(net108),
    .A2(_0534_),
    .Y(_0545_),
    .B1(net147));
 sg13g2_o21ai_1 _1207_ (.B1(net171),
    .Y(_0546_),
    .A1(\system_inst.loader.shift_reg[5] ),
    .A2(_0532_));
 sg13g2_nor2_1 _1208_ (.A(_0545_),
    .B(_0546_),
    .Y(_0074_));
 sg13g2_a21oi_1 _1209_ (.A1(net182),
    .A2(_0534_),
    .Y(_0547_),
    .B1(net147));
 sg13g2_o21ai_1 _1210_ (.B1(net172),
    .Y(_0548_),
    .A1(net96),
    .A2(_0532_));
 sg13g2_nor2_1 _1211_ (.A(_0547_),
    .B(_0548_),
    .Y(_0075_));
 sg13g2_nor2_1 _1212_ (.A(_0505_),
    .B(_0533_),
    .Y(_0549_));
 sg13g2_o21ai_1 _1213_ (.B1(net173),
    .Y(_0550_),
    .A1(net100),
    .A2(_0549_));
 sg13g2_a21oi_1 _1214_ (.A1(net100),
    .A2(_0532_),
    .Y(_0076_),
    .B1(_0550_));
 sg13g2_o21ai_1 _1215_ (.B1(_0498_),
    .Y(_0551_),
    .A1(net113),
    .A2(net100));
 sg13g2_nor2b_1 _1216_ (.A(_0551_),
    .B_N(_0111_),
    .Y(_0552_));
 sg13g2_a22oi_1 _1217_ (.Y(_0553_),
    .B1(_0549_),
    .B2(_0552_),
    .A2(net147),
    .A1(net113));
 sg13g2_nor2_1 _1218_ (.A(net168),
    .B(net114),
    .Y(_0077_));
 sg13g2_a22oi_1 _1219_ (.Y(_0554_),
    .B1(_0497_),
    .B2(_0012_),
    .A2(_0111_),
    .A1(_0011_));
 sg13g2_nor2b_1 _1220_ (.A(net155),
    .B_N(_0554_),
    .Y(_0555_));
 sg13g2_a22oi_1 _1221_ (.Y(_0556_),
    .B1(_0549_),
    .B2(_0555_),
    .A2(net147),
    .A1(net92));
 sg13g2_nor2_1 _1222_ (.A(net168),
    .B(net93),
    .Y(_0078_));
 sg13g2_dfrbp_1 _1223_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net85),
    .D(_0019_),
    .Q_N(_0005_),
    .Q(\system_inst.neuron.v_mem[0] ));
 sg13g2_dfrbp_1 _1224_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net75),
    .D(_0020_),
    .Q_N(_0604_),
    .Q(\system_inst.neuron.v_mem[1] ));
 sg13g2_dfrbp_1 _1225_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net73),
    .D(_0021_),
    .Q_N(_0603_),
    .Q(\system_inst.neuron.v_mem[2] ));
 sg13g2_dfrbp_1 _1226_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net71),
    .D(_0022_),
    .Q_N(_0602_),
    .Q(\system_inst.neuron.v_mem[3] ));
 sg13g2_dfrbp_1 _1227_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net69),
    .D(_0023_),
    .Q_N(_0601_),
    .Q(\system_inst.neuron.v_mem[4] ));
 sg13g2_dfrbp_1 _1228_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net67),
    .D(_0024_),
    .Q_N(_0600_),
    .Q(\system_inst.neuron.v_mem[5] ));
 sg13g2_dfrbp_1 _1229_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net65),
    .D(_0025_),
    .Q_N(_0599_),
    .Q(\system_inst.neuron.v_mem[6] ));
 sg13g2_dfrbp_1 _1230_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net63),
    .D(_0026_),
    .Q_N(_0598_),
    .Q(\system_inst.neuron.v_mem[7] ));
 sg13g2_dfrbp_1 _1231_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net61),
    .D(_0027_),
    .Q_N(_0597_),
    .Q(\system_inst.neuron.v_mem[8] ));
 sg13g2_dfrbp_1 _1232_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net59),
    .D(_0028_),
    .Q_N(_0596_),
    .Q(spike_out));
 sg13g2_dfrbp_1 _1233_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net58),
    .D(net209),
    .Q_N(_0595_),
    .Q(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_dfrbp_1 _1234_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net56),
    .D(_0030_),
    .Q_N(_0594_),
    .Q(\system_inst.neuron.refr_cnt[1] ));
 sg13g2_dfrbp_1 _1235_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net54),
    .D(_0031_),
    .Q_N(_0593_),
    .Q(\system_inst.neuron.refr_cnt[2] ));
 sg13g2_dfrbp_1 _1236_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net52),
    .D(net95),
    .Q_N(_0592_),
    .Q(\system_inst.neuron.refr_cnt[3] ));
 sg13g2_dfrbp_1 _1237_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net50),
    .D(_0033_),
    .Q_N(_0591_),
    .Q(\system_inst.neuron.leak_counter[0] ));
 sg13g2_dfrbp_1 _1238_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net48),
    .D(net112),
    .Q_N(_0590_),
    .Q(\system_inst.neuron.leak_counter[1] ));
 sg13g2_dfrbp_1 _1239_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net46),
    .D(_0035_),
    .Q_N(_0589_),
    .Q(\system_inst.neuron.leak_counter[2] ));
 sg13g2_dfrbp_1 _1240_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net44),
    .D(_0036_),
    .Q_N(_0588_),
    .Q(\system_inst.neuron.leak_counter[3] ));
 sg13g2_dfrbp_1 _1241_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net42),
    .D(_0037_),
    .Q_N(_0009_),
    .Q(\system_inst.neuron.threshold[2] ));
 sg13g2_dfrbp_1 _1242_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net41),
    .D(_0038_),
    .Q_N(_0587_),
    .Q(\system_inst.neuron.threshold[3] ));
 sg13g2_dfrbp_1 _1243_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net40),
    .D(_0039_),
    .Q_N(_0016_),
    .Q(\system_inst.neuron.threshold[4] ));
 sg13g2_dfrbp_1 _1244_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net39),
    .D(net218),
    .Q_N(_0008_),
    .Q(\system_inst.neuron.threshold[5] ));
 sg13g2_dfrbp_1 _1245_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net38),
    .D(_0041_),
    .Q_N(_0007_),
    .Q(\system_inst.neuron.threshold[6] ));
 sg13g2_dfrbp_1 _1246_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net37),
    .D(net193),
    .Q_N(_0006_),
    .Q(\system_inst.neuron.threshold[7] ));
 sg13g2_dfrbp_1 _1247_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net36),
    .D(net131),
    .Q_N(_0010_),
    .Q(\system_inst.neuron.threshold[0] ));
 sg13g2_dfrbp_1 _1248_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net35),
    .D(_0044_),
    .Q_N(_0586_),
    .Q(\system_inst.neuron.threshold[1] ));
 sg13g2_dfrbp_1 _1249_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net34),
    .D(net125),
    .Q_N(_0585_),
    .Q(params_ready));
 sg13g2_dfrbp_1 _1250_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net32),
    .D(_0046_),
    .Q_N(_0584_),
    .Q(\system_inst.loader.weight_a[0] ));
 sg13g2_dfrbp_1 _1251_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net30),
    .D(net123),
    .Q_N(_0583_),
    .Q(\system_inst.loader.weight_a[1] ));
 sg13g2_dfrbp_1 _1252_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net28),
    .D(_0048_),
    .Q_N(_0582_),
    .Q(\system_inst.loader.weight_a[2] ));
 sg13g2_dfrbp_1 _1253_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net26),
    .D(_0049_),
    .Q_N(_0581_),
    .Q(\system_inst.leak_rate[0] ));
 sg13g2_dfrbp_1 _1254_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net84),
    .D(_0050_),
    .Q_N(_0580_),
    .Q(\system_inst.leak_rate[1] ));
 sg13g2_dfrbp_1 _1255_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net82),
    .D(net188),
    .Q_N(_0579_),
    .Q(\system_inst.leak_rate[2] ));
 sg13g2_dfrbp_1 _1256_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net80),
    .D(net129),
    .Q_N(_0578_),
    .Q(\system_inst.leak_rate[3] ));
 sg13g2_dfrbp_1 _1257_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net78),
    .D(net180),
    .Q_N(_0577_),
    .Q(\system_inst.leak_rate[4] ));
 sg13g2_dfrbp_1 _1258_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net76),
    .D(_0054_),
    .Q_N(_0576_),
    .Q(\system_inst.leak_rate[5] ));
 sg13g2_dfrbp_1 _1259_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net72),
    .D(_0055_),
    .Q_N(_0575_),
    .Q(\system_inst.leak_rate[6] ));
 sg13g2_dfrbp_1 _1260_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net68),
    .D(_0056_),
    .Q_N(_0574_),
    .Q(\system_inst.leak_rate[7] ));
 sg13g2_dfrbp_1 _1261_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net64),
    .D(_0057_),
    .Q_N(_0573_),
    .Q(\system_inst.loader.threshold_min[0] ));
 sg13g2_dfrbp_1 _1262_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net60),
    .D(net121),
    .Q_N(_0572_),
    .Q(\system_inst.loader.threshold_min[1] ));
 sg13g2_dfrbp_1 _1263_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net55),
    .D(net199),
    .Q_N(_0018_),
    .Q(\system_inst.loader.threshold_min[2] ));
 sg13g2_dfrbp_1 _1264_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net51),
    .D(_0060_),
    .Q_N(_0017_),
    .Q(\system_inst.loader.threshold_min[3] ));
 sg13g2_dfrbp_1 _1265_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net47),
    .D(_0061_),
    .Q_N(_0015_),
    .Q(\system_inst.loader.threshold_min[4] ));
 sg13g2_dfrbp_1 _1266_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net43),
    .D(_0062_),
    .Q_N(_0014_),
    .Q(\system_inst.loader.threshold_min[5] ));
 sg13g2_dfrbp_1 _1267_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net31),
    .D(_0063_),
    .Q_N(_0013_),
    .Q(\system_inst.loader.threshold_min[6] ));
 sg13g2_dfrbp_1 _1268_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net27),
    .D(net97),
    .Q_N(_0571_),
    .Q(\system_inst.loader.threshold_min[7] ));
 sg13g2_dfrbp_1 _1269_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net83),
    .D(net99),
    .Q_N(_0570_),
    .Q(\system_inst.leak_cycles[0] ));
 sg13g2_dfrbp_1 _1270_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net79),
    .D(_0066_),
    .Q_N(_0569_),
    .Q(\system_inst.leak_cycles[1] ));
 sg13g2_dfrbp_1 _1271_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net74),
    .D(net117),
    .Q_N(_0568_),
    .Q(\system_inst.leak_cycles[2] ));
 sg13g2_dfrbp_1 _1272_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net66),
    .D(net105),
    .Q_N(_0567_),
    .Q(\system_inst.leak_cycles[3] ));
 sg13g2_dfrbp_1 _1273_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net57),
    .D(_0069_),
    .Q_N(_0566_),
    .Q(\system_inst.loader.shift_reg[0] ));
 sg13g2_dfrbp_1 _1274_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net49),
    .D(net127),
    .Q_N(_0565_),
    .Q(\system_inst.loader.shift_reg[1] ));
 sg13g2_dfrbp_1 _1275_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net33),
    .D(_0071_),
    .Q_N(_0564_),
    .Q(\system_inst.loader.shift_reg[2] ));
 sg13g2_dfrbp_1 _1276_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net25),
    .D(_0072_),
    .Q_N(_0563_),
    .Q(\system_inst.loader.shift_reg[3] ));
 sg13g2_dfrbp_1 _1277_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net77),
    .D(_0073_),
    .Q_N(_0562_),
    .Q(\system_inst.loader.shift_reg[4] ));
 sg13g2_dfrbp_1 _1278_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net62),
    .D(net109),
    .Q_N(_0561_),
    .Q(\system_inst.loader.shift_reg[5] ));
 sg13g2_dfrbp_1 _1279_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net45),
    .D(_0075_),
    .Q_N(_0560_),
    .Q(\system_inst.loader.shift_reg[6] ));
 sg13g2_dfrbp_1 _1280_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net81),
    .D(_0076_),
    .Q_N(_0559_),
    .Q(\system_inst.loader.bit_count[0] ));
 sg13g2_dfrbp_1 _1281_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net53),
    .D(_0077_),
    .Q_N(_0558_),
    .Q(\system_inst.loader.bit_count[1] ));
 sg13g2_dfrbp_1 _1282_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net86),
    .D(_0078_),
    .Q_N(_0011_),
    .Q(\system_inst.loader.bit_count[2] ));
 sg13g2_dfrbp_1 _1283_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net87),
    .D(_0000_),
    .Q_N(_0605_),
    .Q(\system_inst.loader.current_state[0] ));
 sg13g2_dfrbp_1 _1284_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net88),
    .D(_0001_),
    .Q_N(_0012_),
    .Q(\system_inst.loader.current_state[1] ));
 sg13g2_dfrbp_1 _1285_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net89),
    .D(_0002_),
    .Q_N(_0606_),
    .Q(\system_inst.loader.current_state[2] ));
 sg13g2_dfrbp_1 _1286_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net29),
    .D(net102),
    .Q_N(_0607_),
    .Q(\system_inst.loader.current_state[3] ));
 sg13g2_dfrbp_1 _1287_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net70),
    .D(_0004_),
    .Q_N(_0557_),
    .Q(\system_inst.loader.current_state[5] ));
 sg13g2_tiehi _1253__26 (.L_HI(net26));
 sg13g2_tiehi _1268__27 (.L_HI(net27));
 sg13g2_tiehi _1252__28 (.L_HI(net28));
 sg13g2_tiehi _1286__29 (.L_HI(net29));
 sg13g2_tiehi _1251__30 (.L_HI(net30));
 sg13g2_tiehi _1267__31 (.L_HI(net31));
 sg13g2_tiehi _1250__32 (.L_HI(net32));
 sg13g2_tiehi _1275__33 (.L_HI(net33));
 sg13g2_tiehi _1249__34 (.L_HI(net34));
 sg13g2_tiehi _1248__35 (.L_HI(net35));
 sg13g2_tiehi _1247__36 (.L_HI(net36));
 sg13g2_tiehi _1246__37 (.L_HI(net37));
 sg13g2_tiehi _1245__38 (.L_HI(net38));
 sg13g2_tiehi _1244__39 (.L_HI(net39));
 sg13g2_tiehi _1243__40 (.L_HI(net40));
 sg13g2_tiehi _1242__41 (.L_HI(net41));
 sg13g2_tiehi _1241__42 (.L_HI(net42));
 sg13g2_tiehi _1266__43 (.L_HI(net43));
 sg13g2_tiehi _1240__44 (.L_HI(net44));
 sg13g2_tiehi _1279__45 (.L_HI(net45));
 sg13g2_tiehi _1239__46 (.L_HI(net46));
 sg13g2_tiehi _1265__47 (.L_HI(net47));
 sg13g2_tiehi _1238__48 (.L_HI(net48));
 sg13g2_tiehi _1274__49 (.L_HI(net49));
 sg13g2_tiehi _1237__50 (.L_HI(net50));
 sg13g2_tiehi _1264__51 (.L_HI(net51));
 sg13g2_tiehi _1236__52 (.L_HI(net52));
 sg13g2_tiehi _1281__53 (.L_HI(net53));
 sg13g2_tiehi _1235__54 (.L_HI(net54));
 sg13g2_tiehi _1263__55 (.L_HI(net55));
 sg13g2_tiehi _1234__56 (.L_HI(net56));
 sg13g2_tiehi _1273__57 (.L_HI(net57));
 sg13g2_tiehi _1233__58 (.L_HI(net58));
 sg13g2_tiehi _1232__59 (.L_HI(net59));
 sg13g2_tiehi _1262__60 (.L_HI(net60));
 sg13g2_tiehi _1231__61 (.L_HI(net61));
 sg13g2_tiehi _1278__62 (.L_HI(net62));
 sg13g2_tiehi _1230__63 (.L_HI(net63));
 sg13g2_tiehi _1261__64 (.L_HI(net64));
 sg13g2_tiehi _1229__65 (.L_HI(net65));
 sg13g2_tiehi _1272__66 (.L_HI(net66));
 sg13g2_tiehi _1228__67 (.L_HI(net67));
 sg13g2_tiehi _1260__68 (.L_HI(net68));
 sg13g2_tiehi _1227__69 (.L_HI(net69));
 sg13g2_tiehi _1287__70 (.L_HI(net70));
 sg13g2_tiehi _1226__71 (.L_HI(net71));
 sg13g2_tiehi _1259__72 (.L_HI(net72));
 sg13g2_tiehi _1225__73 (.L_HI(net73));
 sg13g2_tiehi _1271__74 (.L_HI(net74));
 sg13g2_tiehi _1224__75 (.L_HI(net75));
 sg13g2_tiehi _1258__76 (.L_HI(net76));
 sg13g2_tiehi _1277__77 (.L_HI(net77));
 sg13g2_tiehi _1257__78 (.L_HI(net78));
 sg13g2_tiehi _1270__79 (.L_HI(net79));
 sg13g2_tiehi _1256__80 (.L_HI(net80));
 sg13g2_tiehi _1280__81 (.L_HI(net81));
 sg13g2_tiehi _1255__82 (.L_HI(net82));
 sg13g2_tiehi _1269__83 (.L_HI(net83));
 sg13g2_tiehi _1254__84 (.L_HI(net84));
 sg13g2_tiehi _1223__85 (.L_HI(net85));
 sg13g2_tiehi _1282__86 (.L_HI(net86));
 sg13g2_tiehi _1283__87 (.L_HI(net87));
 sg13g2_tiehi _1284__88 (.L_HI(net88));
 sg13g2_tiehi _1285__89 (.L_HI(net89));
 sg13g2_tiehi tt_um_wokwi_434917506576906241_90 (.L_HI(net90));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_wokwi_434917506576906241_12 (.L_LO(net12));
 sg13g2_tielo tt_um_wokwi_434917506576906241_13 (.L_LO(net13));
 sg13g2_tielo tt_um_wokwi_434917506576906241_14 (.L_LO(net14));
 sg13g2_tielo tt_um_wokwi_434917506576906241_15 (.L_LO(net15));
 sg13g2_tielo tt_um_wokwi_434917506576906241_16 (.L_LO(net16));
 sg13g2_tielo tt_um_wokwi_434917506576906241_17 (.L_LO(net17));
 sg13g2_tielo tt_um_wokwi_434917506576906241_18 (.L_LO(net18));
 sg13g2_tielo tt_um_wokwi_434917506576906241_19 (.L_LO(net19));
 sg13g2_tielo tt_um_wokwi_434917506576906241_20 (.L_LO(net20));
 sg13g2_tielo tt_um_wokwi_434917506576906241_21 (.L_LO(net21));
 sg13g2_tielo tt_um_wokwi_434917506576906241_22 (.L_LO(net22));
 sg13g2_tielo tt_um_wokwi_434917506576906241_23 (.L_LO(net23));
 sg13g2_tielo tt_um_wokwi_434917506576906241_24 (.L_LO(net24));
 sg13g2_tiehi _1276__25 (.L_HI(net25));
 sg13g2_buf_2 _1368_ (.A(params_ready),
    .X(uio_out[0]));
 sg13g2_buf_1 _1369_ (.A(spike_out),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_0440_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(net140),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(net140),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(net140),
    .X(net138));
 sg13g2_buf_1 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_1 fanout140 (.A(_0334_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_0273_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_0433_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_0433_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_0400_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_0400_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_0533_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_0266_),
    .X(net148));
 sg13g2_buf_1 fanout149 (.A(_0266_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_0132_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_0119_),
    .X(net152));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(_0116_));
 sg13g2_buf_2 fanout154 (.A(_0116_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_0112_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(\system_inst.loader.threshold_min[1] ),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(net158),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(net219),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(\system_inst.loader.weight_a[1] ),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(\system_inst.loader.weight_a[0] ),
    .X(net160));
 sg13g2_buf_4 fanout161 (.X(net161),
    .A(net214));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(\system_inst.neuron.threshold[2] ));
 sg13g2_buf_2 fanout163 (.A(net216),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(net167),
    .X(net164));
 sg13g2_buf_1 fanout165 (.A(net167),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_1 fanout167 (.A(net169),
    .X(net167));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(net169));
 sg13g2_buf_2 fanout169 (.A(_0107_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(net6),
    .X(net170));
 sg13g2_buf_4 fanout171 (.X(net171),
    .A(net176));
 sg13g2_buf_2 fanout172 (.A(net174),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(rst_n),
    .X(net176));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_tielo tt_um_wokwi_434917506576906241_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_8_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\system_inst.neuron.v_mem[0] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold2 (.A(\system_inst.loader.bit_count[2] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0556_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold4 (.A(\system_inst.neuron.refr_cnt[3] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0032_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold6 (.A(\system_inst.loader.shift_reg[6] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0064_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold8 (.A(\system_inst.leak_cycles[0] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0065_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold10 (.A(\system_inst.loader.bit_count[0] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold11 (.A(\system_inst.loader.current_state[3] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0003_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold13 (.A(\system_inst.neuron.v_mem[5] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold14 (.A(\system_inst.leak_cycles[3] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0068_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold16 (.A(\system_inst.neuron.v_mem[7] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold17 (.A(\system_inst.loader.current_state[1] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold18 (.A(\system_inst.loader.shift_reg[4] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0074_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold20 (.A(\system_inst.neuron.leak_counter[1] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0364_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0034_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold23 (.A(\system_inst.loader.bit_count[1] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0553_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold25 (.A(\system_inst.leak_rate[7] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold26 (.A(\system_inst.leak_cycles[2] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0067_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold28 (.A(\system_inst.loader.current_state[0] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold29 (.A(\system_inst.loader.threshold_min[1] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0519_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0058_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold32 (.A(\system_inst.loader.weight_a[1] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0047_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold34 (.A(params_ready),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0045_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold36 (.A(\system_inst.loader.shift_reg[0] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0070_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold38 (.A(\system_inst.loader.shift_reg[2] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0052_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold40 (.A(\system_inst.neuron.threshold[0] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0043_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold42 (.A(\system_inst.loader.current_state[2] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold43 (.A(\system_inst.loader.current_state[5] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold44 (.A(\system_inst.neuron.leak_counter[3] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0368_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold46 (.A(\system_inst.loader.shift_reg[3] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0053_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold48 (.A(\system_inst.leak_cycles[1] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold49 (.A(\system_inst.loader.shift_reg[5] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold50 (.A(\system_inst.leak_rate[0] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold51 (.A(\system_inst.neuron.v_mem[6] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold52 (.A(\system_inst.neuron.leak_counter[2] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0367_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold54 (.A(\system_inst.leak_rate[2] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0051_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold56 (.A(\system_inst.neuron.leak_counter[0] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold57 (.A(\system_inst.neuron.v_mem[1] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold58 (.A(\system_inst.neuron.v_mem[4] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold59 (.A(\system_inst.neuron.threshold[7] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold60 (.A(_0042_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold61 (.A(\system_inst.leak_rate[6] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold62 (.A(\system_inst.leak_rate[5] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold63 (.A(\system_inst.neuron.v_mem[2] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold64 (.A(\system_inst.leak_rate[1] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold65 (.A(\system_inst.loader.threshold_min[2] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0059_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold67 (.A(\system_inst.neuron.v_mem[3] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold68 (.A(\system_inst.loader.weight_a[0] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold69 (.A(\system_inst.loader.threshold_min[5] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold70 (.A(\system_inst.loader.threshold_min[4] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold71 (.A(\system_inst.loader.threshold_min[6] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold72 (.A(\system_inst.neuron.threshold[4] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold73 (.A(\system_inst.loader.threshold_min[3] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0009_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold75 (.A(\system_inst.neuron.refr_cnt[0] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0029_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold77 (.A(\system_inst.neuron.threshold[6] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold78 (.A(\system_inst.loader.shift_reg[1] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold79 (.A(\system_inst.neuron.refr_cnt[2] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0359_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold81 (.A(\system_inst.neuron.threshold[3] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold82 (.A(\system_inst.neuron.threshold[1] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold83 (.A(\system_inst.neuron.v_mem[8] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold84 (.A(\system_inst.neuron.threshold[5] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0040_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold86 (.A(\system_inst.loader.weight_a[2] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold87 (.A(\system_inst.loader.threshold_min[0] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold88 (.A(\system_inst.neuron.refr_cnt[1] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0358_),
    .X(net222));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_4 FILLER_11_287 ();
 sg13g2_fill_1 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_296 ();
 sg13g2_decap_8 FILLER_11_303 ();
 sg13g2_decap_8 FILLER_11_310 ();
 sg13g2_decap_8 FILLER_11_317 ();
 sg13g2_decap_8 FILLER_11_324 ();
 sg13g2_decap_8 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_345 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_373 ();
 sg13g2_decap_8 FILLER_11_380 ();
 sg13g2_decap_8 FILLER_11_387 ();
 sg13g2_decap_8 FILLER_11_394 ();
 sg13g2_decap_8 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_fill_1 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_313 ();
 sg13g2_decap_4 FILLER_12_320 ();
 sg13g2_fill_2 FILLER_12_333 ();
 sg13g2_fill_2 FILLER_12_339 ();
 sg13g2_fill_1 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_345 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_373 ();
 sg13g2_decap_8 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_387 ();
 sg13g2_decap_8 FILLER_12_394 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_4 FILLER_13_266 ();
 sg13g2_fill_2 FILLER_13_270 ();
 sg13g2_fill_1 FILLER_13_276 ();
 sg13g2_fill_2 FILLER_13_281 ();
 sg13g2_fill_2 FILLER_13_304 ();
 sg13g2_fill_1 FILLER_13_337 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_4 FILLER_14_252 ();
 sg13g2_fill_2 FILLER_14_256 ();
 sg13g2_fill_2 FILLER_14_309 ();
 sg13g2_fill_1 FILLER_14_329 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_fill_1 FILLER_14_353 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_decap_8 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_4 FILLER_15_231 ();
 sg13g2_fill_2 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_286 ();
 sg13g2_fill_1 FILLER_15_330 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_4 FILLER_16_196 ();
 sg13g2_fill_1 FILLER_16_200 ();
 sg13g2_decap_8 FILLER_16_227 ();
 sg13g2_decap_8 FILLER_16_234 ();
 sg13g2_decap_4 FILLER_16_241 ();
 sg13g2_fill_2 FILLER_16_258 ();
 sg13g2_fill_1 FILLER_16_260 ();
 sg13g2_fill_1 FILLER_16_292 ();
 sg13g2_fill_2 FILLER_16_311 ();
 sg13g2_fill_2 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_4 FILLER_16_361 ();
 sg13g2_fill_1 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_fill_2 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_111 ();
 sg13g2_decap_8 FILLER_17_118 ();
 sg13g2_decap_8 FILLER_17_125 ();
 sg13g2_fill_2 FILLER_17_132 ();
 sg13g2_fill_1 FILLER_17_134 ();
 sg13g2_decap_8 FILLER_17_139 ();
 sg13g2_decap_8 FILLER_17_146 ();
 sg13g2_decap_8 FILLER_17_153 ();
 sg13g2_fill_2 FILLER_17_160 ();
 sg13g2_fill_1 FILLER_17_162 ();
 sg13g2_decap_8 FILLER_17_166 ();
 sg13g2_decap_8 FILLER_17_173 ();
 sg13g2_decap_8 FILLER_17_180 ();
 sg13g2_decap_8 FILLER_17_187 ();
 sg13g2_decap_8 FILLER_17_194 ();
 sg13g2_decap_8 FILLER_17_201 ();
 sg13g2_fill_1 FILLER_17_208 ();
 sg13g2_decap_4 FILLER_17_227 ();
 sg13g2_fill_2 FILLER_17_231 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_fill_2 FILLER_17_246 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_decap_4 FILLER_17_253 ();
 sg13g2_fill_1 FILLER_17_257 ();
 sg13g2_decap_8 FILLER_17_261 ();
 sg13g2_decap_8 FILLER_17_268 ();
 sg13g2_fill_2 FILLER_17_275 ();
 sg13g2_decap_4 FILLER_17_303 ();
 sg13g2_fill_2 FILLER_17_307 ();
 sg13g2_fill_1 FILLER_17_340 ();
 sg13g2_fill_2 FILLER_17_354 ();
 sg13g2_fill_1 FILLER_17_356 ();
 sg13g2_fill_2 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_4 FILLER_18_91 ();
 sg13g2_fill_2 FILLER_18_95 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_fill_1 FILLER_18_157 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_fill_2 FILLER_18_235 ();
 sg13g2_fill_1 FILLER_18_237 ();
 sg13g2_decap_4 FILLER_18_314 ();
 sg13g2_fill_2 FILLER_18_318 ();
 sg13g2_fill_2 FILLER_18_324 ();
 sg13g2_fill_1 FILLER_18_326 ();
 sg13g2_fill_1 FILLER_18_357 ();
 sg13g2_fill_2 FILLER_18_367 ();
 sg13g2_decap_4 FILLER_18_388 ();
 sg13g2_fill_2 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_85 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_fill_2 FILLER_19_112 ();
 sg13g2_fill_1 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_152 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_173 ();
 sg13g2_decap_8 FILLER_19_183 ();
 sg13g2_decap_4 FILLER_19_190 ();
 sg13g2_fill_1 FILLER_19_194 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_decap_8 FILLER_19_229 ();
 sg13g2_fill_2 FILLER_19_236 ();
 sg13g2_fill_1 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_243 ();
 sg13g2_fill_2 FILLER_19_250 ();
 sg13g2_decap_4 FILLER_19_261 ();
 sg13g2_fill_1 FILLER_19_265 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_fill_2 FILLER_19_277 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_fill_2 FILLER_19_323 ();
 sg13g2_fill_1 FILLER_19_330 ();
 sg13g2_fill_1 FILLER_19_341 ();
 sg13g2_fill_2 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_fill_2 FILLER_19_363 ();
 sg13g2_fill_1 FILLER_19_369 ();
 sg13g2_fill_2 FILLER_19_380 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_4 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_59 ();
 sg13g2_fill_1 FILLER_20_66 ();
 sg13g2_fill_2 FILLER_20_89 ();
 sg13g2_fill_1 FILLER_20_96 ();
 sg13g2_fill_1 FILLER_20_107 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_decap_4 FILLER_20_124 ();
 sg13g2_fill_2 FILLER_20_128 ();
 sg13g2_fill_2 FILLER_20_135 ();
 sg13g2_fill_2 FILLER_20_142 ();
 sg13g2_fill_1 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_157 ();
 sg13g2_fill_2 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_decap_4 FILLER_20_205 ();
 sg13g2_fill_1 FILLER_20_209 ();
 sg13g2_fill_1 FILLER_20_254 ();
 sg13g2_decap_4 FILLER_20_281 ();
 sg13g2_fill_1 FILLER_20_285 ();
 sg13g2_fill_2 FILLER_20_291 ();
 sg13g2_fill_1 FILLER_20_293 ();
 sg13g2_decap_4 FILLER_20_320 ();
 sg13g2_fill_1 FILLER_20_324 ();
 sg13g2_fill_2 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_4 FILLER_20_389 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_fill_2 FILLER_21_48 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_fill_1 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_fill_2 FILLER_21_121 ();
 sg13g2_fill_1 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_149 ();
 sg13g2_fill_2 FILLER_21_156 ();
 sg13g2_fill_1 FILLER_21_165 ();
 sg13g2_decap_4 FILLER_21_170 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_fill_2 FILLER_21_203 ();
 sg13g2_fill_1 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_213 ();
 sg13g2_decap_8 FILLER_21_220 ();
 sg13g2_fill_2 FILLER_21_227 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_fill_2 FILLER_21_283 ();
 sg13g2_fill_1 FILLER_21_285 ();
 sg13g2_fill_2 FILLER_21_300 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_decap_4 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_351 ();
 sg13g2_fill_2 FILLER_21_357 ();
 sg13g2_fill_2 FILLER_21_367 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_46 ();
 sg13g2_fill_2 FILLER_22_53 ();
 sg13g2_fill_2 FILLER_22_73 ();
 sg13g2_fill_1 FILLER_22_75 ();
 sg13g2_fill_2 FILLER_22_84 ();
 sg13g2_decap_4 FILLER_22_94 ();
 sg13g2_fill_1 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_129 ();
 sg13g2_decap_8 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_fill_2 FILLER_22_155 ();
 sg13g2_fill_1 FILLER_22_162 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_185 ();
 sg13g2_fill_2 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_229 ();
 sg13g2_fill_1 FILLER_22_231 ();
 sg13g2_fill_2 FILLER_22_258 ();
 sg13g2_fill_1 FILLER_22_317 ();
 sg13g2_decap_4 FILLER_22_356 ();
 sg13g2_fill_2 FILLER_22_360 ();
 sg13g2_fill_2 FILLER_22_372 ();
 sg13g2_fill_2 FILLER_22_388 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_23 ();
 sg13g2_fill_2 FILLER_23_62 ();
 sg13g2_decap_8 FILLER_23_69 ();
 sg13g2_fill_2 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_78 ();
 sg13g2_decap_4 FILLER_23_88 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_107 ();
 sg13g2_decap_4 FILLER_23_112 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_fill_1 FILLER_23_150 ();
 sg13g2_fill_1 FILLER_23_162 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_4 FILLER_23_214 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_244 ();
 sg13g2_fill_2 FILLER_23_255 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_decap_8 FILLER_23_281 ();
 sg13g2_decap_4 FILLER_23_288 ();
 sg13g2_fill_1 FILLER_23_292 ();
 sg13g2_fill_2 FILLER_23_316 ();
 sg13g2_fill_1 FILLER_23_318 ();
 sg13g2_decap_4 FILLER_23_325 ();
 sg13g2_decap_8 FILLER_23_352 ();
 sg13g2_fill_2 FILLER_23_359 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_4 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_46 ();
 sg13g2_fill_2 FILLER_24_71 ();
 sg13g2_decap_4 FILLER_24_89 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_fill_1 FILLER_24_109 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_125 ();
 sg13g2_fill_2 FILLER_24_144 ();
 sg13g2_fill_1 FILLER_24_146 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_fill_1 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_164 ();
 sg13g2_decap_8 FILLER_24_171 ();
 sg13g2_fill_2 FILLER_24_178 ();
 sg13g2_decap_4 FILLER_24_196 ();
 sg13g2_fill_1 FILLER_24_200 ();
 sg13g2_fill_2 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_269 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_4 FILLER_24_338 ();
 sg13g2_fill_2 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_decap_4 FILLER_24_363 ();
 sg13g2_fill_2 FILLER_24_367 ();
 sg13g2_fill_1 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_58 ();
 sg13g2_fill_1 FILLER_25_60 ();
 sg13g2_decap_8 FILLER_25_71 ();
 sg13g2_fill_2 FILLER_25_78 ();
 sg13g2_fill_1 FILLER_25_80 ();
 sg13g2_decap_8 FILLER_25_86 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_4 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_127 ();
 sg13g2_decap_4 FILLER_25_134 ();
 sg13g2_fill_2 FILLER_25_138 ();
 sg13g2_fill_2 FILLER_25_173 ();
 sg13g2_fill_1 FILLER_25_175 ();
 sg13g2_decap_4 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_185 ();
 sg13g2_decap_8 FILLER_25_190 ();
 sg13g2_decap_8 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_decap_4 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_4 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_281 ();
 sg13g2_decap_8 FILLER_25_286 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_fill_1 FILLER_25_300 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_371 ();
 sg13g2_fill_1 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_2 FILLER_26_25 ();
 sg13g2_fill_1 FILLER_26_60 ();
 sg13g2_fill_2 FILLER_26_69 ();
 sg13g2_fill_1 FILLER_26_71 ();
 sg13g2_fill_1 FILLER_26_86 ();
 sg13g2_fill_2 FILLER_26_102 ();
 sg13g2_decap_4 FILLER_26_131 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_fill_2 FILLER_26_193 ();
 sg13g2_fill_1 FILLER_26_195 ();
 sg13g2_fill_2 FILLER_26_222 ();
 sg13g2_decap_8 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_301 ();
 sg13g2_fill_2 FILLER_26_312 ();
 sg13g2_decap_4 FILLER_26_326 ();
 sg13g2_fill_2 FILLER_26_330 ();
 sg13g2_fill_2 FILLER_26_337 ();
 sg13g2_fill_1 FILLER_26_339 ();
 sg13g2_decap_4 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_fill_2 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_fill_1 FILLER_26_393 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_4 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_fill_1 FILLER_27_60 ();
 sg13g2_decap_4 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_decap_4 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_102 ();
 sg13g2_fill_1 FILLER_27_104 ();
 sg13g2_decap_4 FILLER_27_110 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_2 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_125 ();
 sg13g2_decap_4 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_134 ();
 sg13g2_fill_2 FILLER_27_148 ();
 sg13g2_fill_1 FILLER_27_150 ();
 sg13g2_decap_4 FILLER_27_156 ();
 sg13g2_fill_2 FILLER_27_160 ();
 sg13g2_decap_4 FILLER_27_167 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_decap_4 FILLER_27_203 ();
 sg13g2_fill_2 FILLER_27_207 ();
 sg13g2_decap_8 FILLER_27_229 ();
 sg13g2_decap_4 FILLER_27_236 ();
 sg13g2_decap_8 FILLER_27_253 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_fill_2 FILLER_27_324 ();
 sg13g2_decap_8 FILLER_27_362 ();
 sg13g2_fill_2 FILLER_27_377 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_44 ();
 sg13g2_fill_2 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_decap_8 FILLER_28_67 ();
 sg13g2_decap_4 FILLER_28_74 ();
 sg13g2_fill_2 FILLER_28_78 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_fill_2 FILLER_28_91 ();
 sg13g2_fill_2 FILLER_28_111 ();
 sg13g2_fill_1 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_135 ();
 sg13g2_decap_8 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_150 ();
 sg13g2_decap_8 FILLER_28_171 ();
 sg13g2_decap_4 FILLER_28_178 ();
 sg13g2_fill_2 FILLER_28_182 ();
 sg13g2_fill_1 FILLER_28_197 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_fill_1 FILLER_28_210 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_decap_8 FILLER_28_220 ();
 sg13g2_decap_8 FILLER_28_227 ();
 sg13g2_decap_8 FILLER_28_234 ();
 sg13g2_fill_2 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_decap_8 FILLER_28_267 ();
 sg13g2_decap_8 FILLER_28_274 ();
 sg13g2_fill_2 FILLER_28_281 ();
 sg13g2_decap_8 FILLER_28_293 ();
 sg13g2_decap_8 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_307 ();
 sg13g2_decap_8 FILLER_28_317 ();
 sg13g2_fill_2 FILLER_28_324 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_decap_4 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_4 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_82 ();
 sg13g2_fill_1 FILLER_29_89 ();
 sg13g2_decap_8 FILLER_29_94 ();
 sg13g2_decap_8 FILLER_29_101 ();
 sg13g2_decap_8 FILLER_29_108 ();
 sg13g2_decap_8 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_122 ();
 sg13g2_decap_8 FILLER_29_130 ();
 sg13g2_decap_4 FILLER_29_137 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_4 FILLER_29_182 ();
 sg13g2_fill_2 FILLER_29_198 ();
 sg13g2_fill_2 FILLER_29_210 ();
 sg13g2_fill_2 FILLER_29_220 ();
 sg13g2_fill_1 FILLER_29_222 ();
 sg13g2_fill_2 FILLER_29_244 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_fill_2 FILLER_29_276 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_fill_1 FILLER_29_331 ();
 sg13g2_decap_4 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_4 FILLER_30_49 ();
 sg13g2_fill_1 FILLER_30_61 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_decap_4 FILLER_30_131 ();
 sg13g2_decap_8 FILLER_30_156 ();
 sg13g2_fill_2 FILLER_30_163 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_169 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_206 ();
 sg13g2_decap_8 FILLER_30_213 ();
 sg13g2_decap_8 FILLER_30_220 ();
 sg13g2_fill_1 FILLER_30_227 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_decap_8 FILLER_30_247 ();
 sg13g2_decap_8 FILLER_30_254 ();
 sg13g2_decap_8 FILLER_30_269 ();
 sg13g2_decap_4 FILLER_30_276 ();
 sg13g2_fill_2 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_290 ();
 sg13g2_decap_8 FILLER_30_300 ();
 sg13g2_decap_8 FILLER_30_311 ();
 sg13g2_decap_4 FILLER_30_318 ();
 sg13g2_decap_8 FILLER_30_332 ();
 sg13g2_decap_4 FILLER_30_339 ();
 sg13g2_fill_1 FILLER_30_343 ();
 sg13g2_fill_1 FILLER_30_352 ();
 sg13g2_fill_2 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_fill_1 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_49 ();
 sg13g2_fill_2 FILLER_31_53 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_decap_4 FILLER_31_127 ();
 sg13g2_fill_1 FILLER_31_131 ();
 sg13g2_decap_4 FILLER_31_136 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_146 ();
 sg13g2_decap_4 FILLER_31_153 ();
 sg13g2_fill_2 FILLER_31_167 ();
 sg13g2_decap_4 FILLER_31_179 ();
 sg13g2_fill_1 FILLER_31_183 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_fill_1 FILLER_31_203 ();
 sg13g2_fill_2 FILLER_31_218 ();
 sg13g2_fill_1 FILLER_31_220 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_4 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_257 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_decap_4 FILLER_31_279 ();
 sg13g2_fill_1 FILLER_31_283 ();
 sg13g2_decap_4 FILLER_31_304 ();
 sg13g2_fill_2 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_335 ();
 sg13g2_fill_2 FILLER_31_347 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_4 FILLER_32_63 ();
 sg13g2_fill_2 FILLER_32_67 ();
 sg13g2_fill_2 FILLER_32_74 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_1 FILLER_32_107 ();
 sg13g2_fill_2 FILLER_32_113 ();
 sg13g2_decap_8 FILLER_32_120 ();
 sg13g2_decap_8 FILLER_32_127 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_fill_2 FILLER_32_155 ();
 sg13g2_decap_8 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_184 ();
 sg13g2_decap_8 FILLER_32_194 ();
 sg13g2_fill_2 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_212 ();
 sg13g2_fill_2 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_233 ();
 sg13g2_decap_4 FILLER_32_243 ();
 sg13g2_fill_1 FILLER_32_247 ();
 sg13g2_fill_2 FILLER_32_261 ();
 sg13g2_decap_8 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_278 ();
 sg13g2_decap_8 FILLER_32_285 ();
 sg13g2_fill_1 FILLER_32_292 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_decap_4 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_fill_2 FILLER_32_331 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_32_353 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_fill_1 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_4 FILLER_33_91 ();
 sg13g2_fill_1 FILLER_33_127 ();
 sg13g2_decap_8 FILLER_33_143 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_fill_1 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_decap_4 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_240 ();
 sg13g2_decap_4 FILLER_33_247 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_fill_1 FILLER_33_258 ();
 sg13g2_decap_4 FILLER_33_272 ();
 sg13g2_fill_2 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_305 ();
 sg13g2_decap_4 FILLER_33_312 ();
 sg13g2_decap_4 FILLER_33_328 ();
 sg13g2_fill_2 FILLER_33_332 ();
 sg13g2_decap_4 FILLER_33_347 ();
 sg13g2_fill_2 FILLER_33_351 ();
 sg13g2_fill_2 FILLER_33_374 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_4 FILLER_34_105 ();
 sg13g2_fill_1 FILLER_34_109 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_fill_1 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_165 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_190 ();
 sg13g2_decap_8 FILLER_34_197 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_246 ();
 sg13g2_decap_8 FILLER_34_265 ();
 sg13g2_fill_2 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_287 ();
 sg13g2_decap_4 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_330 ();
 sg13g2_fill_2 FILLER_34_337 ();
 sg13g2_fill_1 FILLER_34_339 ();
 sg13g2_fill_2 FILLER_34_345 ();
 sg13g2_decap_4 FILLER_34_357 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_fill_2 FILLER_34_367 ();
 sg13g2_fill_1 FILLER_34_369 ();
 sg13g2_fill_1 FILLER_34_397 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_127 ();
 sg13g2_fill_1 FILLER_35_129 ();
 sg13g2_decap_4 FILLER_35_136 ();
 sg13g2_decap_8 FILLER_35_148 ();
 sg13g2_fill_2 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_2 FILLER_35_167 ();
 sg13g2_decap_8 FILLER_35_199 ();
 sg13g2_decap_4 FILLER_35_218 ();
 sg13g2_fill_2 FILLER_35_222 ();
 sg13g2_fill_1 FILLER_35_228 ();
 sg13g2_decap_8 FILLER_35_242 ();
 sg13g2_decap_8 FILLER_35_249 ();
 sg13g2_fill_2 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_264 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_4 FILLER_35_280 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_decap_8 FILLER_35_298 ();
 sg13g2_decap_8 FILLER_35_305 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_fill_2 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_347 ();
 sg13g2_fill_1 FILLER_35_370 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_116 ();
 sg13g2_decap_4 FILLER_36_180 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_decap_4 FILLER_36_243 ();
 sg13g2_decap_4 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_269 ();
 sg13g2_decap_8 FILLER_36_274 ();
 sg13g2_fill_2 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_283 ();
 sg13g2_decap_8 FILLER_36_296 ();
 sg13g2_fill_2 FILLER_36_303 ();
 sg13g2_decap_4 FILLER_36_330 ();
 sg13g2_fill_1 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_fill_1 FILLER_36_346 ();
 sg13g2_fill_1 FILLER_36_350 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_357 ();
 sg13g2_fill_2 FILLER_36_371 ();
 sg13g2_fill_2 FILLER_36_392 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_127 ();
 sg13g2_fill_2 FILLER_37_147 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_fill_1 FILLER_37_163 ();
 sg13g2_fill_2 FILLER_37_195 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_fill_2 FILLER_37_206 ();
 sg13g2_decap_8 FILLER_37_221 ();
 sg13g2_decap_8 FILLER_37_228 ();
 sg13g2_fill_2 FILLER_37_240 ();
 sg13g2_fill_1 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_275 ();
 sg13g2_fill_2 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_305 ();
 sg13g2_fill_1 FILLER_37_319 ();
 sg13g2_fill_2 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_339 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_fill_2 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_183 ();
 sg13g2_fill_1 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_192 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_decap_8 FILLER_38_233 ();
 sg13g2_decap_4 FILLER_38_251 ();
 sg13g2_fill_1 FILLER_38_255 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_4 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_282 ();
 sg13g2_decap_4 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_fill_1 FILLER_38_309 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_349 ();
 assign uio_oe[0] = net90;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net12;
 assign uio_oe[3] = net13;
 assign uio_oe[4] = net14;
 assign uio_oe[5] = net15;
 assign uio_oe[6] = net16;
 assign uio_oe[7] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule
