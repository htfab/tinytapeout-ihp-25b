module tt_um_pwm_block (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \MemCell.counter[0] ;
 wire \MemCell.counter[1] ;
 wire \MemCell.counter_value[0] ;
 wire \MemCell.counter_value[10] ;
 wire \MemCell.counter_value[11] ;
 wire \MemCell.counter_value[12] ;
 wire \MemCell.counter_value[13] ;
 wire \MemCell.counter_value[14] ;
 wire \MemCell.counter_value[15] ;
 wire \MemCell.counter_value[16] ;
 wire \MemCell.counter_value[17] ;
 wire \MemCell.counter_value[18] ;
 wire \MemCell.counter_value[19] ;
 wire \MemCell.counter_value[1] ;
 wire \MemCell.counter_value[20] ;
 wire \MemCell.counter_value[21] ;
 wire \MemCell.counter_value[22] ;
 wire \MemCell.counter_value[23] ;
 wire \MemCell.counter_value[24] ;
 wire \MemCell.counter_value[25] ;
 wire \MemCell.counter_value[26] ;
 wire \MemCell.counter_value[27] ;
 wire \MemCell.counter_value[28] ;
 wire \MemCell.counter_value[29] ;
 wire \MemCell.counter_value[2] ;
 wire \MemCell.counter_value[30] ;
 wire \MemCell.counter_value[31] ;
 wire \MemCell.counter_value[3] ;
 wire \MemCell.counter_value[4] ;
 wire \MemCell.counter_value[5] ;
 wire \MemCell.counter_value[6] ;
 wire \MemCell.counter_value[7] ;
 wire \MemCell.counter_value[8] ;
 wire \MemCell.counter_value[9] ;
 wire \MemCell.curr_state[0] ;
 wire \MemCell.curr_state[1] ;
 wire \MemCell.curr_state[2] ;
 wire \MemCell.dc1_reg[0][0] ;
 wire \MemCell.dc1_reg[0][1] ;
 wire \MemCell.dc1_reg[0][2] ;
 wire \MemCell.dc1_reg[0][3] ;
 wire \MemCell.dc1_reg[0][4] ;
 wire \MemCell.dc1_reg[0][5] ;
 wire \MemCell.dc1_reg[0][6] ;
 wire \MemCell.dc1_reg[0][7] ;
 wire \MemCell.dc1_reg[1][0] ;
 wire \MemCell.dc1_reg[1][1] ;
 wire \MemCell.dc1_reg[1][2] ;
 wire \MemCell.dc1_reg[1][3] ;
 wire \MemCell.dc1_reg[1][4] ;
 wire \MemCell.dc1_reg[1][5] ;
 wire \MemCell.dc1_reg[1][6] ;
 wire \MemCell.dc1_reg[1][7] ;
 wire \MemCell.dc1_reg[2][0] ;
 wire \MemCell.dc1_reg[2][1] ;
 wire \MemCell.dc1_reg[2][2] ;
 wire \MemCell.dc1_reg[2][3] ;
 wire \MemCell.dc1_reg[2][4] ;
 wire \MemCell.dc1_reg[2][5] ;
 wire \MemCell.dc1_reg[2][6] ;
 wire \MemCell.dc1_reg[2][7] ;
 wire \MemCell.dc1_reg[3][0] ;
 wire \MemCell.dc1_reg[3][1] ;
 wire \MemCell.dc1_reg[3][2] ;
 wire \MemCell.dc1_reg[3][3] ;
 wire \MemCell.dc1_reg[3][4] ;
 wire \MemCell.dc1_reg[3][5] ;
 wire \MemCell.dc1_reg[3][6] ;
 wire \MemCell.dc1_reg[3][7] ;
 wire \MemCell.dc2_reg[0][0] ;
 wire \MemCell.dc2_reg[0][1] ;
 wire \MemCell.dc2_reg[0][2] ;
 wire \MemCell.dc2_reg[0][3] ;
 wire \MemCell.dc2_reg[0][4] ;
 wire \MemCell.dc2_reg[0][5] ;
 wire \MemCell.dc2_reg[0][6] ;
 wire \MemCell.dc2_reg[0][7] ;
 wire \MemCell.dc2_reg[1][0] ;
 wire \MemCell.dc2_reg[1][1] ;
 wire \MemCell.dc2_reg[1][2] ;
 wire \MemCell.dc2_reg[1][3] ;
 wire \MemCell.dc2_reg[1][4] ;
 wire \MemCell.dc2_reg[1][5] ;
 wire \MemCell.dc2_reg[1][6] ;
 wire \MemCell.dc2_reg[1][7] ;
 wire \MemCell.dc2_reg[2][0] ;
 wire \MemCell.dc2_reg[2][1] ;
 wire \MemCell.dc2_reg[2][2] ;
 wire \MemCell.dc2_reg[2][3] ;
 wire \MemCell.dc2_reg[2][4] ;
 wire \MemCell.dc2_reg[2][5] ;
 wire \MemCell.dc2_reg[2][6] ;
 wire \MemCell.dc2_reg[2][7] ;
 wire \MemCell.dc2_reg[3][0] ;
 wire \MemCell.dc2_reg[3][1] ;
 wire \MemCell.dc2_reg[3][2] ;
 wire \MemCell.dc2_reg[3][3] ;
 wire \MemCell.dc2_reg[3][4] ;
 wire \MemCell.dc2_reg[3][5] ;
 wire \MemCell.dc2_reg[3][6] ;
 wire \MemCell.dc2_reg[3][7] ;
 wire \MemCell.dc3_reg[0][0] ;
 wire \MemCell.dc3_reg[0][1] ;
 wire \MemCell.dc3_reg[0][2] ;
 wire \MemCell.dc3_reg[0][3] ;
 wire \MemCell.dc3_reg[0][4] ;
 wire \MemCell.dc3_reg[0][5] ;
 wire \MemCell.dc3_reg[0][6] ;
 wire \MemCell.dc3_reg[0][7] ;
 wire \MemCell.dc3_reg[1][0] ;
 wire \MemCell.dc3_reg[1][1] ;
 wire \MemCell.dc3_reg[1][2] ;
 wire \MemCell.dc3_reg[1][3] ;
 wire \MemCell.dc3_reg[1][4] ;
 wire \MemCell.dc3_reg[1][5] ;
 wire \MemCell.dc3_reg[1][6] ;
 wire \MemCell.dc3_reg[1][7] ;
 wire \MemCell.dc3_reg[2][0] ;
 wire \MemCell.dc3_reg[2][1] ;
 wire \MemCell.dc3_reg[2][2] ;
 wire \MemCell.dc3_reg[2][3] ;
 wire \MemCell.dc3_reg[2][4] ;
 wire \MemCell.dc3_reg[2][5] ;
 wire \MemCell.dc3_reg[2][6] ;
 wire \MemCell.dc3_reg[2][7] ;
 wire \MemCell.dc3_reg[3][0] ;
 wire \MemCell.dc3_reg[3][1] ;
 wire \MemCell.dc3_reg[3][2] ;
 wire \MemCell.dc3_reg[3][3] ;
 wire \MemCell.dc3_reg[3][4] ;
 wire \MemCell.dc3_reg[3][5] ;
 wire \MemCell.dc3_reg[3][6] ;
 wire \MemCell.dc3_reg[3][7] ;
 wire \MemCell.enable_pwm ;
 wire \MemCell.next_state[0] ;
 wire \MemCell.next_state[1] ;
 wire \MemCell.next_state[2] ;
 wire \MemCell.o_RX_Byte[0] ;
 wire \MemCell.o_RX_Byte[1] ;
 wire \MemCell.o_RX_Byte[2] ;
 wire \MemCell.o_RX_Byte[3] ;
 wire \MemCell.o_RX_Byte[4] ;
 wire \MemCell.o_RX_Byte[5] ;
 wire \MemCell.o_RX_Byte[6] ;
 wire \MemCell.o_RX_Byte[7] ;
 wire \MemCell.o_RX_DV ;
 wire \MemCell.prescale_reg[0][0] ;
 wire \MemCell.prescale_reg[0][1] ;
 wire \MemCell.prescale_reg[0][2] ;
 wire \MemCell.prescale_reg[0][3] ;
 wire \MemCell.prescale_reg[0][4] ;
 wire \MemCell.prescale_reg[0][5] ;
 wire \MemCell.prescale_reg[0][6] ;
 wire \MemCell.prescale_reg[0][7] ;
 wire \MemCell.prescale_reg[1][0] ;
 wire \MemCell.prescale_reg[1][1] ;
 wire \MemCell.prescale_reg[1][2] ;
 wire \MemCell.prescale_reg[1][3] ;
 wire \MemCell.prescale_reg[1][4] ;
 wire \MemCell.prescale_reg[1][5] ;
 wire \MemCell.prescale_reg[1][6] ;
 wire \MemCell.prescale_reg[1][7] ;
 wire \MemCell.prescale_reg[2][0] ;
 wire \MemCell.prescale_reg[2][1] ;
 wire \MemCell.prescale_reg[2][2] ;
 wire \MemCell.prescale_reg[2][3] ;
 wire \MemCell.prescale_reg[2][4] ;
 wire \MemCell.prescale_reg[2][5] ;
 wire \MemCell.prescale_reg[2][6] ;
 wire \MemCell.prescale_reg[2][7] ;
 wire \MemCell.prescale_reg[3][0] ;
 wire \MemCell.prescale_reg[3][1] ;
 wire \MemCell.prescale_reg[3][2] ;
 wire \MemCell.prescale_reg[3][3] ;
 wire \MemCell.prescale_reg[3][4] ;
 wire \MemCell.prescale_reg[3][5] ;
 wire \MemCell.prescale_reg[3][6] ;
 wire \MemCell.prescale_reg[3][7] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire \pwm_module.counter0[0] ;
 wire \pwm_module.counter0[10] ;
 wire \pwm_module.counter0[11] ;
 wire \pwm_module.counter0[12] ;
 wire \pwm_module.counter0[13] ;
 wire \pwm_module.counter0[14] ;
 wire \pwm_module.counter0[15] ;
 wire \pwm_module.counter0[16] ;
 wire \pwm_module.counter0[17] ;
 wire \pwm_module.counter0[18] ;
 wire \pwm_module.counter0[19] ;
 wire \pwm_module.counter0[1] ;
 wire \pwm_module.counter0[20] ;
 wire \pwm_module.counter0[21] ;
 wire \pwm_module.counter0[22] ;
 wire \pwm_module.counter0[23] ;
 wire \pwm_module.counter0[24] ;
 wire \pwm_module.counter0[25] ;
 wire \pwm_module.counter0[26] ;
 wire \pwm_module.counter0[27] ;
 wire \pwm_module.counter0[28] ;
 wire \pwm_module.counter0[29] ;
 wire \pwm_module.counter0[2] ;
 wire \pwm_module.counter0[30] ;
 wire \pwm_module.counter0[31] ;
 wire \pwm_module.counter0[3] ;
 wire \pwm_module.counter0[4] ;
 wire \pwm_module.counter0[5] ;
 wire \pwm_module.counter0[6] ;
 wire \pwm_module.counter0[7] ;
 wire \pwm_module.counter0[8] ;
 wire \pwm_module.counter0[9] ;
 wire \pwm_module.counter1[0] ;
 wire \pwm_module.counter1[10] ;
 wire \pwm_module.counter1[11] ;
 wire \pwm_module.counter1[12] ;
 wire \pwm_module.counter1[13] ;
 wire \pwm_module.counter1[14] ;
 wire \pwm_module.counter1[15] ;
 wire \pwm_module.counter1[16] ;
 wire \pwm_module.counter1[17] ;
 wire \pwm_module.counter1[18] ;
 wire \pwm_module.counter1[19] ;
 wire \pwm_module.counter1[1] ;
 wire \pwm_module.counter1[20] ;
 wire \pwm_module.counter1[21] ;
 wire \pwm_module.counter1[22] ;
 wire \pwm_module.counter1[23] ;
 wire \pwm_module.counter1[24] ;
 wire \pwm_module.counter1[25] ;
 wire \pwm_module.counter1[26] ;
 wire \pwm_module.counter1[27] ;
 wire \pwm_module.counter1[28] ;
 wire \pwm_module.counter1[29] ;
 wire \pwm_module.counter1[2] ;
 wire \pwm_module.counter1[30] ;
 wire \pwm_module.counter1[31] ;
 wire \pwm_module.counter1[3] ;
 wire \pwm_module.counter1[4] ;
 wire \pwm_module.counter1[5] ;
 wire \pwm_module.counter1[6] ;
 wire \pwm_module.counter1[7] ;
 wire \pwm_module.counter1[8] ;
 wire \pwm_module.counter1[9] ;
 wire \pwm_module.counter2[0] ;
 wire \pwm_module.counter2[10] ;
 wire \pwm_module.counter2[11] ;
 wire \pwm_module.counter2[12] ;
 wire \pwm_module.counter2[13] ;
 wire \pwm_module.counter2[14] ;
 wire \pwm_module.counter2[15] ;
 wire \pwm_module.counter2[16] ;
 wire \pwm_module.counter2[17] ;
 wire \pwm_module.counter2[18] ;
 wire \pwm_module.counter2[19] ;
 wire \pwm_module.counter2[1] ;
 wire \pwm_module.counter2[20] ;
 wire \pwm_module.counter2[21] ;
 wire \pwm_module.counter2[22] ;
 wire \pwm_module.counter2[23] ;
 wire \pwm_module.counter2[24] ;
 wire \pwm_module.counter2[25] ;
 wire \pwm_module.counter2[26] ;
 wire \pwm_module.counter2[27] ;
 wire \pwm_module.counter2[28] ;
 wire \pwm_module.counter2[29] ;
 wire \pwm_module.counter2[2] ;
 wire \pwm_module.counter2[30] ;
 wire \pwm_module.counter2[31] ;
 wire \pwm_module.counter2[3] ;
 wire \pwm_module.counter2[4] ;
 wire \pwm_module.counter2[5] ;
 wire \pwm_module.counter2[6] ;
 wire \pwm_module.counter2[7] ;
 wire \pwm_module.counter2[8] ;
 wire \pwm_module.counter2[9] ;
 wire \pwm_module.prescaler0[0] ;
 wire \pwm_module.prescaler0[10] ;
 wire \pwm_module.prescaler0[11] ;
 wire \pwm_module.prescaler0[12] ;
 wire \pwm_module.prescaler0[13] ;
 wire \pwm_module.prescaler0[14] ;
 wire \pwm_module.prescaler0[15] ;
 wire \pwm_module.prescaler0[16] ;
 wire \pwm_module.prescaler0[17] ;
 wire \pwm_module.prescaler0[18] ;
 wire \pwm_module.prescaler0[19] ;
 wire \pwm_module.prescaler0[1] ;
 wire \pwm_module.prescaler0[20] ;
 wire \pwm_module.prescaler0[21] ;
 wire \pwm_module.prescaler0[22] ;
 wire \pwm_module.prescaler0[23] ;
 wire \pwm_module.prescaler0[24] ;
 wire \pwm_module.prescaler0[25] ;
 wire \pwm_module.prescaler0[26] ;
 wire \pwm_module.prescaler0[27] ;
 wire \pwm_module.prescaler0[28] ;
 wire \pwm_module.prescaler0[29] ;
 wire \pwm_module.prescaler0[2] ;
 wire \pwm_module.prescaler0[30] ;
 wire \pwm_module.prescaler0[31] ;
 wire \pwm_module.prescaler0[3] ;
 wire \pwm_module.prescaler0[4] ;
 wire \pwm_module.prescaler0[5] ;
 wire \pwm_module.prescaler0[6] ;
 wire \pwm_module.prescaler0[7] ;
 wire \pwm_module.prescaler0[8] ;
 wire \pwm_module.prescaler0[9] ;
 wire \pwm_module.prescaler1[0] ;
 wire \pwm_module.prescaler1[10] ;
 wire \pwm_module.prescaler1[11] ;
 wire \pwm_module.prescaler1[12] ;
 wire \pwm_module.prescaler1[13] ;
 wire \pwm_module.prescaler1[14] ;
 wire \pwm_module.prescaler1[15] ;
 wire \pwm_module.prescaler1[16] ;
 wire \pwm_module.prescaler1[17] ;
 wire \pwm_module.prescaler1[18] ;
 wire \pwm_module.prescaler1[19] ;
 wire \pwm_module.prescaler1[1] ;
 wire \pwm_module.prescaler1[20] ;
 wire \pwm_module.prescaler1[21] ;
 wire \pwm_module.prescaler1[22] ;
 wire \pwm_module.prescaler1[23] ;
 wire \pwm_module.prescaler1[24] ;
 wire \pwm_module.prescaler1[25] ;
 wire \pwm_module.prescaler1[26] ;
 wire \pwm_module.prescaler1[27] ;
 wire \pwm_module.prescaler1[28] ;
 wire \pwm_module.prescaler1[29] ;
 wire \pwm_module.prescaler1[2] ;
 wire \pwm_module.prescaler1[30] ;
 wire \pwm_module.prescaler1[31] ;
 wire \pwm_module.prescaler1[3] ;
 wire \pwm_module.prescaler1[4] ;
 wire \pwm_module.prescaler1[5] ;
 wire \pwm_module.prescaler1[6] ;
 wire \pwm_module.prescaler1[7] ;
 wire \pwm_module.prescaler1[8] ;
 wire \pwm_module.prescaler1[9] ;
 wire \pwm_module.prescaler2[0] ;
 wire \pwm_module.prescaler2[10] ;
 wire \pwm_module.prescaler2[11] ;
 wire \pwm_module.prescaler2[12] ;
 wire \pwm_module.prescaler2[13] ;
 wire \pwm_module.prescaler2[14] ;
 wire \pwm_module.prescaler2[15] ;
 wire \pwm_module.prescaler2[16] ;
 wire \pwm_module.prescaler2[17] ;
 wire \pwm_module.prescaler2[18] ;
 wire \pwm_module.prescaler2[19] ;
 wire \pwm_module.prescaler2[1] ;
 wire \pwm_module.prescaler2[20] ;
 wire \pwm_module.prescaler2[21] ;
 wire \pwm_module.prescaler2[22] ;
 wire \pwm_module.prescaler2[23] ;
 wire \pwm_module.prescaler2[24] ;
 wire \pwm_module.prescaler2[25] ;
 wire \pwm_module.prescaler2[26] ;
 wire \pwm_module.prescaler2[27] ;
 wire \pwm_module.prescaler2[28] ;
 wire \pwm_module.prescaler2[29] ;
 wire \pwm_module.prescaler2[2] ;
 wire \pwm_module.prescaler2[30] ;
 wire \pwm_module.prescaler2[31] ;
 wire \pwm_module.prescaler2[3] ;
 wire \pwm_module.prescaler2[4] ;
 wire \pwm_module.prescaler2[5] ;
 wire \pwm_module.prescaler2[6] ;
 wire \pwm_module.prescaler2[7] ;
 wire \pwm_module.prescaler2[8] ;
 wire \pwm_module.prescaler2[9] ;
 wire \spi_module.r2_RX_Done ;
 wire \spi_module.r3_RX_Done ;
 wire \spi_module.r_RX_Bit_Count[0] ;
 wire \spi_module.r_RX_Bit_Count[1] ;
 wire \spi_module.r_RX_Bit_Count[2] ;
 wire \spi_module.r_RX_Byte[0] ;
 wire \spi_module.r_RX_Byte[1] ;
 wire \spi_module.r_RX_Byte[2] ;
 wire \spi_module.r_RX_Byte[3] ;
 wire \spi_module.r_RX_Byte[4] ;
 wire \spi_module.r_RX_Byte[5] ;
 wire \spi_module.r_RX_Byte[6] ;
 wire \spi_module.r_RX_Byte[7] ;
 wire \spi_module.r_RX_Done ;
 wire \spi_module.r_Temp_RX_Byte[0] ;
 wire \spi_module.r_Temp_RX_Byte[1] ;
 wire \spi_module.r_Temp_RX_Byte[2] ;
 wire \spi_module.r_Temp_RX_Byte[3] ;
 wire \spi_module.r_Temp_RX_Byte[4] ;
 wire \spi_module.r_Temp_RX_Byte[5] ;
 wire \spi_module.r_Temp_RX_Byte[6] ;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net3;
 wire clknet_leaf_0_clk;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net1;
 wire net2;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;

 sg13g2_inv_1 _2402_ (.Y(_1785_),
    .A(net490));
 sg13g2_inv_1 _2403_ (.Y(_1786_),
    .A(net473));
 sg13g2_inv_1 _2404_ (.Y(_1787_),
    .A(net185));
 sg13g2_inv_1 _2405_ (.Y(_1788_),
    .A(net391));
 sg13g2_inv_1 _2406_ (.Y(_1789_),
    .A(net197));
 sg13g2_inv_1 _2407_ (.Y(_1790_),
    .A(net183));
 sg13g2_inv_1 _2408_ (.Y(_1791_),
    .A(\pwm_module.counter1[12] ));
 sg13g2_inv_1 _2409_ (.Y(_1792_),
    .A(\pwm_module.counter1[11] ));
 sg13g2_inv_1 _2410_ (.Y(_1793_),
    .A(\pwm_module.counter1[10] ));
 sg13g2_inv_1 _2411_ (.Y(_1794_),
    .A(net143));
 sg13g2_inv_1 _2412_ (.Y(_1795_),
    .A(net559));
 sg13g2_inv_1 _2413_ (.Y(_1796_),
    .A(net141));
 sg13g2_inv_1 _2414_ (.Y(_1797_),
    .A(\pwm_module.counter1[8] ));
 sg13g2_inv_1 _2415_ (.Y(_1798_),
    .A(net485));
 sg13g2_inv_1 _2416_ (.Y(_1799_),
    .A(\pwm_module.counter1[6] ));
 sg13g2_inv_1 _2417_ (.Y(_1800_),
    .A(net138));
 sg13g2_inv_1 _2418_ (.Y(_1801_),
    .A(\pwm_module.counter1[4] ));
 sg13g2_inv_1 _2419_ (.Y(_1802_),
    .A(net67));
 sg13g2_inv_1 _2420_ (.Y(_1803_),
    .A(\pwm_module.counter1[3] ));
 sg13g2_inv_2 _2421_ (.Y(_1804_),
    .A(net188));
 sg13g2_inv_1 _2422_ (.Y(_1805_),
    .A(net146));
 sg13g2_inv_1 _2423_ (.Y(_1806_),
    .A(net163));
 sg13g2_inv_1 _2424_ (.Y(_1807_),
    .A(net450));
 sg13g2_inv_1 _2425_ (.Y(_1808_),
    .A(net98));
 sg13g2_inv_1 _2426_ (.Y(_1809_),
    .A(net531));
 sg13g2_inv_1 _2427_ (.Y(_1810_),
    .A(\pwm_module.counter2[28] ));
 sg13g2_inv_1 _2428_ (.Y(_1811_),
    .A(net217));
 sg13g2_inv_1 _2429_ (.Y(_1812_),
    .A(\pwm_module.counter2[26] ));
 sg13g2_inv_1 _2430_ (.Y(_1813_),
    .A(net196));
 sg13g2_inv_1 _2431_ (.Y(_1814_),
    .A(net463));
 sg13g2_inv_1 _2432_ (.Y(_1815_),
    .A(net214));
 sg13g2_inv_2 _2433_ (.Y(_1816_),
    .A(net524));
 sg13g2_inv_1 _2434_ (.Y(_1817_),
    .A(net427));
 sg13g2_inv_1 _2435_ (.Y(_1818_),
    .A(net195));
 sg13g2_inv_1 _2436_ (.Y(_1819_),
    .A(net194));
 sg13g2_inv_1 _2437_ (.Y(_1820_),
    .A(net542));
 sg13g2_inv_1 _2438_ (.Y(_1821_),
    .A(net526));
 sg13g2_inv_1 _2439_ (.Y(_1822_),
    .A(net535));
 sg13g2_inv_1 _2440_ (.Y(_1823_),
    .A(\pwm_module.counter2[15] ));
 sg13g2_inv_1 _2441_ (.Y(_1824_),
    .A(net184));
 sg13g2_inv_1 _2442_ (.Y(_1825_),
    .A(net377));
 sg13g2_inv_1 _2443_ (.Y(_1826_),
    .A(net182));
 sg13g2_inv_1 _2444_ (.Y(_1827_),
    .A(net482));
 sg13g2_inv_1 _2445_ (.Y(_1828_),
    .A(net140));
 sg13g2_inv_1 _2446_ (.Y(_1829_),
    .A(\pwm_module.counter2[12] ));
 sg13g2_inv_1 _2447_ (.Y(_1830_),
    .A(net340));
 sg13g2_inv_1 _2448_ (.Y(_1831_),
    .A(net129));
 sg13g2_inv_1 _2449_ (.Y(_1832_),
    .A(net295));
 sg13g2_inv_1 _2450_ (.Y(_1833_),
    .A(net161));
 sg13g2_inv_1 _2451_ (.Y(_1834_),
    .A(\pwm_module.counter2[8] ));
 sg13g2_inv_1 _2452_ (.Y(_1835_),
    .A(net464));
 sg13g2_inv_2 _2453_ (.Y(_1836_),
    .A(\pwm_module.counter2[6] ));
 sg13g2_inv_1 _2454_ (.Y(_1837_),
    .A(net121));
 sg13g2_inv_1 _2455_ (.Y(_1838_),
    .A(net360));
 sg13g2_inv_1 _2456_ (.Y(_1839_),
    .A(\pwm_module.counter2[4] ));
 sg13g2_inv_1 _2457_ (.Y(_1840_),
    .A(net187));
 sg13g2_inv_1 _2458_ (.Y(_1841_),
    .A(\pwm_module.counter2[3] ));
 sg13g2_inv_1 _2459_ (.Y(_1842_),
    .A(\pwm_module.counter2[2] ));
 sg13g2_inv_1 _2460_ (.Y(_1843_),
    .A(net649));
 sg13g2_inv_1 _2461_ (.Y(_1844_),
    .A(net362));
 sg13g2_inv_1 _2462_ (.Y(_1845_),
    .A(\MemCell.curr_state[1] ));
 sg13g2_inv_1 _2463_ (.Y(_1846_),
    .A(\MemCell.o_RX_DV ));
 sg13g2_inv_1 _2464_ (.Y(_1847_),
    .A(net429));
 sg13g2_inv_1 _2465_ (.Y(_1848_),
    .A(\pwm_module.prescaler1[2] ));
 sg13g2_inv_1 _2466_ (.Y(_1849_),
    .A(net424));
 sg13g2_inv_1 _2467_ (.Y(_1850_),
    .A(\MemCell.prescale_reg[0][4] ));
 sg13g2_inv_1 _2468_ (.Y(_1851_),
    .A(\pwm_module.prescaler1[14] ));
 sg13g2_inv_1 _2469_ (.Y(_1852_),
    .A(\pwm_module.prescaler1[13] ));
 sg13g2_inv_1 _2470_ (.Y(_1853_),
    .A(\pwm_module.prescaler1[12] ));
 sg13g2_inv_1 _2471_ (.Y(_1854_),
    .A(net345));
 sg13g2_inv_2 _2472_ (.Y(_1855_),
    .A(net364));
 sg13g2_inv_2 _2473_ (.Y(_1856_),
    .A(net298));
 sg13g2_inv_2 _2474_ (.Y(_1857_),
    .A(net442));
 sg13g2_inv_1 _2475_ (.Y(_1858_),
    .A(\MemCell.prescale_reg[3][1] ));
 sg13g2_inv_1 _2476_ (.Y(_1859_),
    .A(\MemCell.prescale_reg[3][0] ));
 sg13g2_inv_1 _2477_ (.Y(_1860_),
    .A(\MemCell.prescale_reg[2][5] ));
 sg13g2_inv_1 _2478_ (.Y(_1861_),
    .A(net280));
 sg13g2_inv_1 _2479_ (.Y(_1862_),
    .A(\MemCell.prescale_reg[2][4] ));
 sg13g2_inv_2 _2480_ (.Y(_1863_),
    .A(net385));
 sg13g2_inv_1 _2481_ (.Y(_1864_),
    .A(\pwm_module.prescaler2[4] ));
 sg13g2_inv_1 _2482_ (.Y(_1865_),
    .A(\pwm_module.prescaler2[3] ));
 sg13g2_inv_1 _2483_ (.Y(_1866_),
    .A(\pwm_module.prescaler2[2] ));
 sg13g2_inv_1 _2484_ (.Y(_1867_),
    .A(\pwm_module.prescaler0[20] ));
 sg13g2_inv_1 _2485_ (.Y(_1868_),
    .A(\pwm_module.prescaler0[16] ));
 sg13g2_inv_1 _2486_ (.Y(_1869_),
    .A(\pwm_module.prescaler0[13] ));
 sg13g2_inv_1 _2487_ (.Y(_1870_),
    .A(\pwm_module.prescaler0[6] ));
 sg13g2_inv_1 _2488_ (.Y(_1871_),
    .A(\pwm_module.prescaler0[2] ));
 sg13g2_inv_1 _2489_ (.Y(_0104_),
    .A(net683));
 sg13g2_inv_1 _2490_ (.Y(_1872_),
    .A(net290));
 sg13g2_inv_1 _2491_ (.Y(_1873_),
    .A(net440));
 sg13g2_inv_1 _2492_ (.Y(_1874_),
    .A(net471));
 sg13g2_inv_2 _2493_ (.Y(_1875_),
    .A(net335));
 sg13g2_inv_1 _2494_ (.Y(_1876_),
    .A(net546));
 sg13g2_inv_1 _2495_ (.Y(_1877_),
    .A(net342));
 sg13g2_inv_1 _2496_ (.Y(_1878_),
    .A(net434));
 sg13g2_inv_1 _2497_ (.Y(_1879_),
    .A(\pwm_module.counter0[25] ));
 sg13g2_inv_1 _2498_ (.Y(_1880_),
    .A(net443));
 sg13g2_inv_1 _2499_ (.Y(_1881_),
    .A(\pwm_module.counter0[24] ));
 sg13g2_inv_2 _2500_ (.Y(_1882_),
    .A(net409));
 sg13g2_inv_1 _2501_ (.Y(_1883_),
    .A(\pwm_module.counter0[23] ));
 sg13g2_inv_1 _2502_ (.Y(_1884_),
    .A(net502));
 sg13g2_inv_1 _2503_ (.Y(_1885_),
    .A(net373));
 sg13g2_inv_1 _2504_ (.Y(_1886_),
    .A(net513));
 sg13g2_inv_1 _2505_ (.Y(_1887_),
    .A(net367));
 sg13g2_inv_1 _2506_ (.Y(_1888_),
    .A(net483));
 sg13g2_inv_1 _2507_ (.Y(_1889_),
    .A(net503));
 sg13g2_inv_1 _2508_ (.Y(_1890_),
    .A(net398));
 sg13g2_inv_1 _2509_ (.Y(_1891_),
    .A(net497));
 sg13g2_inv_1 _2510_ (.Y(_1892_),
    .A(\pwm_module.counter0[18] ));
 sg13g2_inv_1 _2511_ (.Y(_1893_),
    .A(net478));
 sg13g2_inv_1 _2512_ (.Y(_1894_),
    .A(\pwm_module.counter0[17] ));
 sg13g2_inv_1 _2513_ (.Y(_1895_),
    .A(net461));
 sg13g2_inv_1 _2514_ (.Y(_1896_),
    .A(\pwm_module.counter0[16] ));
 sg13g2_inv_1 _2515_ (.Y(_1897_),
    .A(net457));
 sg13g2_inv_2 _2516_ (.Y(_1898_),
    .A(net462));
 sg13g2_inv_1 _2517_ (.Y(_1899_),
    .A(net488));
 sg13g2_inv_1 _2518_ (.Y(_1900_),
    .A(net408));
 sg13g2_inv_1 _2519_ (.Y(_1901_),
    .A(\pwm_module.counter0[13] ));
 sg13g2_inv_1 _2520_ (.Y(_1902_),
    .A(\pwm_module.counter0[12] ));
 sg13g2_inv_1 _2521_ (.Y(_1903_),
    .A(net510));
 sg13g2_inv_1 _2522_ (.Y(_1904_),
    .A(net380));
 sg13g2_inv_1 _2523_ (.Y(_1905_),
    .A(net288));
 sg13g2_inv_1 _2524_ (.Y(_1906_),
    .A(net351));
 sg13g2_inv_1 _2525_ (.Y(_1907_),
    .A(\pwm_module.counter0[8] ));
 sg13g2_inv_1 _2526_ (.Y(_1908_),
    .A(net469));
 sg13g2_inv_1 _2527_ (.Y(_1909_),
    .A(net394));
 sg13g2_inv_1 _2528_ (.Y(_1910_),
    .A(net511));
 sg13g2_inv_2 _2529_ (.Y(_1911_),
    .A(net305));
 sg13g2_inv_1 _2530_ (.Y(_1912_),
    .A(net498));
 sg13g2_inv_1 _2531_ (.Y(_1913_),
    .A(\pwm_module.counter0[4] ));
 sg13g2_inv_1 _2532_ (.Y(_1914_),
    .A(net530));
 sg13g2_inv_1 _2533_ (.Y(_1915_),
    .A(\pwm_module.counter0[3] ));
 sg13g2_inv_2 _2534_ (.Y(_1916_),
    .A(net215));
 sg13g2_inv_1 _2535_ (.Y(_1917_),
    .A(net240));
 sg13g2_inv_1 _2536_ (.Y(_1918_),
    .A(net500));
 sg13g2_inv_1 _2537_ (.Y(_1919_),
    .A(net515));
 sg13g2_inv_2 _2538_ (.Y(_1920_),
    .A(net383));
 sg13g2_inv_1 _2539_ (.Y(_1921_),
    .A(net369));
 sg13g2_inv_1 _2540_ (.Y(_1922_),
    .A(\pwm_module.counter1[21] ));
 sg13g2_inv_1 _2541_ (.Y(_1923_),
    .A(net514));
 sg13g2_inv_1 _2542_ (.Y(_1924_),
    .A(net402));
 sg13g2_inv_1 _2543_ (.Y(_1925_),
    .A(net459));
 sg13g2_inv_1 _2544_ (.Y(_1926_),
    .A(net160));
 sg13g2_inv_1 _2545_ (.Y(_1927_),
    .A(net153));
 sg13g2_inv_1 _2546_ (.Y(_1928_),
    .A(net294));
 sg13g2_inv_1 _2547_ (.Y(_1929_),
    .A(net297));
 sg13g2_inv_1 _2548_ (.Y(_1930_),
    .A(\MemCell.dc1_reg[3][0] ));
 sg13g2_inv_1 _2549_ (.Y(_1931_),
    .A(net144));
 sg13g2_inv_1 _2550_ (.Y(_1932_),
    .A(net177));
 sg13g2_inv_1 _2551_ (.Y(_1933_),
    .A(net125));
 sg13g2_inv_1 _2552_ (.Y(_1934_),
    .A(net169));
 sg13g2_inv_1 _2553_ (.Y(_1935_),
    .A(net108));
 sg13g2_inv_1 _2554_ (.Y(_1936_),
    .A(net227));
 sg13g2_inv_1 _2555_ (.Y(_1937_),
    .A(net130));
 sg13g2_inv_1 _2556_ (.Y(_1938_),
    .A(net151));
 sg13g2_inv_1 _2557_ (.Y(_1939_),
    .A(net156));
 sg13g2_inv_1 _2558_ (.Y(_1940_),
    .A(net210));
 sg13g2_inv_1 _2559_ (.Y(_1941_),
    .A(net242));
 sg13g2_inv_1 _2560_ (.Y(_1942_),
    .A(net109));
 sg13g2_inv_1 _2561_ (.Y(_1943_),
    .A(net272));
 sg13g2_nand2b_1 _2562_ (.Y(_1944_),
    .B(\spi_module.r_RX_Bit_Count[1] ),
    .A_N(\spi_module.r_RX_Bit_Count[0] ));
 sg13g2_nand3_1 _2563_ (.B(\spi_module.r_RX_Bit_Count[0] ),
    .C(\spi_module.r_RX_Bit_Count[2] ),
    .A(\spi_module.r_RX_Bit_Count[1] ),
    .Y(_1945_));
 sg13g2_o21ai_1 _2564_ (.B1(\spi_module.r_RX_Done ),
    .Y(_1946_),
    .A1(\spi_module.r_RX_Bit_Count[2] ),
    .A2(_1944_));
 sg13g2_nand2_1 _2565_ (.Y(_0163_),
    .A(_1945_),
    .B(_1946_));
 sg13g2_nand2b_1 _2566_ (.Y(_1947_),
    .B(\pwm_module.counter1[15] ),
    .A_N(\MemCell.dc2_reg[1][7] ));
 sg13g2_o21ai_1 _2567_ (.B1(_1947_),
    .Y(_1948_),
    .A1(\MemCell.dc2_reg[1][6] ),
    .A2(_1788_));
 sg13g2_nand2_1 _2568_ (.Y(_1949_),
    .A(\MemCell.dc2_reg[1][7] ),
    .B(_1786_));
 sg13g2_o21ai_1 _2569_ (.B1(_1949_),
    .Y(_1950_),
    .A1(_1787_),
    .A2(\pwm_module.counter1[14] ));
 sg13g2_a22oi_1 _2570_ (.Y(_1951_),
    .B1(_1790_),
    .B2(\pwm_module.counter1[12] ),
    .A2(\pwm_module.counter1[13] ),
    .A1(_1789_));
 sg13g2_nor2_1 _2571_ (.A(_1789_),
    .B(\pwm_module.counter1[13] ),
    .Y(_1952_));
 sg13g2_nand2b_1 _2572_ (.Y(_1953_),
    .B(\pwm_module.counter1[1] ),
    .A_N(\MemCell.dc2_reg[0][1] ));
 sg13g2_nor2b_1 _2573_ (.A(\pwm_module.counter1[0] ),
    .B_N(\MemCell.dc2_reg[0][0] ),
    .Y(_1954_));
 sg13g2_nor2b_1 _2574_ (.A(\pwm_module.counter1[1] ),
    .B_N(\MemCell.dc2_reg[0][1] ),
    .Y(_1955_));
 sg13g2_a221oi_1 _2575_ (.B2(_1954_),
    .C1(_1955_),
    .B1(_1953_),
    .A1(\MemCell.dc2_reg[0][2] ),
    .Y(_1956_),
    .A2(_1804_));
 sg13g2_nand2b_1 _2576_ (.Y(_1957_),
    .B(\pwm_module.counter1[3] ),
    .A_N(\MemCell.dc2_reg[0][3] ));
 sg13g2_o21ai_1 _2577_ (.B1(_1957_),
    .Y(_1958_),
    .A1(\MemCell.dc2_reg[0][2] ),
    .A2(_1804_));
 sg13g2_a22oi_1 _2578_ (.Y(_1959_),
    .B1(\MemCell.dc2_reg[0][3] ),
    .B2(_1803_),
    .A2(\MemCell.dc2_reg[0][4] ),
    .A1(_1801_));
 sg13g2_o21ai_1 _2579_ (.B1(_1959_),
    .Y(_1960_),
    .A1(_1956_),
    .A2(_1958_));
 sg13g2_a22oi_1 _2580_ (.Y(_1961_),
    .B1(\pwm_module.counter1[4] ),
    .B2(_1802_),
    .A2(net647),
    .A1(_1800_));
 sg13g2_nor2_1 _2581_ (.A(_1800_),
    .B(net647),
    .Y(_1962_));
 sg13g2_a221oi_1 _2582_ (.B2(_1961_),
    .C1(_1962_),
    .B1(_1960_),
    .A1(\MemCell.dc2_reg[0][6] ),
    .Y(_1963_),
    .A2(_1799_));
 sg13g2_nand2b_1 _2583_ (.Y(_1964_),
    .B(\pwm_module.counter1[7] ),
    .A_N(\MemCell.dc2_reg[0][7] ));
 sg13g2_o21ai_1 _2584_ (.B1(_1964_),
    .Y(_1965_),
    .A1(\MemCell.dc2_reg[0][6] ),
    .A2(_1799_));
 sg13g2_a22oi_1 _2585_ (.Y(_1966_),
    .B1(\MemCell.dc2_reg[0][7] ),
    .B2(_1798_),
    .A2(_1797_),
    .A1(\MemCell.dc2_reg[1][0] ));
 sg13g2_o21ai_1 _2586_ (.B1(_1966_),
    .Y(_1967_),
    .A1(_1963_),
    .A2(_1965_));
 sg13g2_a22oi_1 _2587_ (.Y(_1968_),
    .B1(_1796_),
    .B2(\pwm_module.counter1[8] ),
    .A2(\pwm_module.counter1[9] ),
    .A1(_1794_));
 sg13g2_nor2b_1 _2588_ (.A(\pwm_module.counter1[10] ),
    .B_N(\MemCell.dc2_reg[1][2] ),
    .Y(_1969_));
 sg13g2_a221oi_1 _2589_ (.B2(_1968_),
    .C1(_1969_),
    .B1(_1967_),
    .A1(\MemCell.dc2_reg[1][1] ),
    .Y(_1970_),
    .A2(_1795_));
 sg13g2_nand2b_1 _2590_ (.Y(_1971_),
    .B(\pwm_module.counter1[11] ),
    .A_N(\MemCell.dc2_reg[1][3] ));
 sg13g2_o21ai_1 _2591_ (.B1(_1971_),
    .Y(_1972_),
    .A1(\MemCell.dc2_reg[1][2] ),
    .A2(_1793_));
 sg13g2_a221oi_1 _2592_ (.B2(_1792_),
    .C1(_1952_),
    .B1(\MemCell.dc2_reg[1][3] ),
    .A1(\MemCell.dc2_reg[1][4] ),
    .Y(_1973_),
    .A2(_1791_));
 sg13g2_nand2_1 _2593_ (.Y(_1974_),
    .A(_1951_),
    .B(_1973_));
 sg13g2_nor3_1 _2594_ (.A(_1948_),
    .B(_1950_),
    .C(_1974_),
    .Y(_1975_));
 sg13g2_o21ai_1 _2595_ (.B1(_1975_),
    .Y(_1976_),
    .A1(_1970_),
    .A2(_1972_));
 sg13g2_nor4_1 _2596_ (.A(_1948_),
    .B(_1950_),
    .C(_1951_),
    .D(_1952_),
    .Y(_1977_));
 sg13g2_a21oi_1 _2597_ (.A1(_1948_),
    .A2(_1949_),
    .Y(_1978_),
    .B1(_1977_));
 sg13g2_nor2_1 _2598_ (.A(_1917_),
    .B(\MemCell.dc2_reg[3][7] ),
    .Y(_1979_));
 sg13g2_nor2_1 _2599_ (.A(_1918_),
    .B(\MemCell.dc2_reg[3][6] ),
    .Y(_1980_));
 sg13g2_nor2_1 _2600_ (.A(_1979_),
    .B(_1980_),
    .Y(_1981_));
 sg13g2_nand2b_1 _2601_ (.Y(_1982_),
    .B(\pwm_module.counter1[25] ),
    .A_N(\MemCell.dc2_reg[3][1] ));
 sg13g2_nand2b_1 _2602_ (.Y(_1983_),
    .B(\pwm_module.counter1[24] ),
    .A_N(\MemCell.dc2_reg[3][0] ));
 sg13g2_nor2b_1 _2603_ (.A(\pwm_module.counter1[31] ),
    .B_N(\MemCell.dc2_reg[3][7] ),
    .Y(_1984_));
 sg13g2_a21o_1 _2604_ (.A2(\MemCell.dc2_reg[3][6] ),
    .A1(_1918_),
    .B1(_1984_),
    .X(_1985_));
 sg13g2_a22oi_1 _2605_ (.Y(_1986_),
    .B1(_1940_),
    .B2(\pwm_module.counter1[28] ),
    .A2(_1939_),
    .A1(\pwm_module.counter1[29] ));
 sg13g2_nand2_1 _2606_ (.Y(_1987_),
    .A(\pwm_module.counter1[26] ),
    .B(_1941_));
 sg13g2_o21ai_1 _2607_ (.B1(_1987_),
    .Y(_1988_),
    .A1(_1919_),
    .A2(\MemCell.dc2_reg[3][3] ));
 sg13g2_nand2_1 _2608_ (.Y(_1989_),
    .A(_1919_),
    .B(\MemCell.dc2_reg[3][3] ));
 sg13g2_o21ai_1 _2609_ (.B1(_1989_),
    .Y(_1990_),
    .A1(\pwm_module.counter1[26] ),
    .A2(_1941_));
 sg13g2_nor2_1 _2610_ (.A(_1988_),
    .B(_1990_),
    .Y(_1991_));
 sg13g2_nor2_1 _2611_ (.A(\pwm_module.counter1[28] ),
    .B(_1940_),
    .Y(_1992_));
 sg13g2_nand2b_1 _2612_ (.Y(_1993_),
    .B(\MemCell.dc2_reg[3][0] ),
    .A_N(\pwm_module.counter1[24] ));
 sg13g2_nand2b_1 _2613_ (.Y(_1994_),
    .B(\MemCell.dc2_reg[3][5] ),
    .A_N(\pwm_module.counter1[29] ));
 sg13g2_nor2b_1 _2614_ (.A(\pwm_module.counter1[25] ),
    .B_N(\MemCell.dc2_reg[3][1] ),
    .Y(_1995_));
 sg13g2_nand4_1 _2615_ (.B(_1982_),
    .C(_1986_),
    .A(_1981_),
    .Y(_1996_),
    .D(_1994_));
 sg13g2_nor4_1 _2616_ (.A(_1985_),
    .B(_1992_),
    .C(_1995_),
    .D(_1996_),
    .Y(_1997_));
 sg13g2_nand4_1 _2617_ (.B(_1991_),
    .C(_1993_),
    .A(_1983_),
    .Y(_0391_),
    .D(_1997_));
 sg13g2_nand2b_1 _2618_ (.Y(_0392_),
    .B(\pwm_module.counter1[18] ),
    .A_N(\MemCell.dc2_reg[2][2] ));
 sg13g2_o21ai_1 _2619_ (.B1(_0392_),
    .Y(_0393_),
    .A1(_1924_),
    .A2(\MemCell.dc2_reg[2][3] ));
 sg13g2_nand2b_1 _2620_ (.Y(_0394_),
    .B(\MemCell.dc2_reg[2][2] ),
    .A_N(\pwm_module.counter1[18] ));
 sg13g2_nand2_1 _2621_ (.Y(_0395_),
    .A(_1924_),
    .B(\MemCell.dc2_reg[2][3] ));
 sg13g2_nand3b_1 _2622_ (.B(_0394_),
    .C(_0395_),
    .Y(_0396_),
    .A_N(_0393_));
 sg13g2_nand2b_1 _2623_ (.Y(_0397_),
    .B(\pwm_module.counter1[22] ),
    .A_N(\MemCell.dc2_reg[2][6] ));
 sg13g2_o21ai_1 _2624_ (.B1(_0397_),
    .Y(_0398_),
    .A1(_1920_),
    .A2(\MemCell.dc2_reg[2][7] ));
 sg13g2_nand2_1 _2625_ (.Y(_0399_),
    .A(_1920_),
    .B(\MemCell.dc2_reg[2][7] ));
 sg13g2_a22oi_1 _2626_ (.Y(_0400_),
    .B1(\MemCell.dc2_reg[2][6] ),
    .B2(_1921_),
    .A2(\MemCell.dc2_reg[2][7] ),
    .A1(_1920_));
 sg13g2_nand2b_1 _2627_ (.Y(_0401_),
    .B(_0400_),
    .A_N(_0398_));
 sg13g2_nand2_1 _2628_ (.Y(_0402_),
    .A(_1922_),
    .B(\MemCell.dc2_reg[2][5] ));
 sg13g2_nand2_1 _2629_ (.Y(_0403_),
    .A(_1925_),
    .B(\MemCell.dc2_reg[2][1] ));
 sg13g2_nor2_1 _2630_ (.A(\pwm_module.counter1[20] ),
    .B(_1943_),
    .Y(_0404_));
 sg13g2_a22oi_1 _2631_ (.Y(_0405_),
    .B1(_1943_),
    .B2(\pwm_module.counter1[20] ),
    .A2(_1942_),
    .A1(\pwm_module.counter1[21] ));
 sg13g2_nand2b_1 _2632_ (.Y(_0406_),
    .B(\pwm_module.counter1[17] ),
    .A_N(\MemCell.dc2_reg[2][1] ));
 sg13g2_o21ai_1 _2633_ (.B1(_0406_),
    .Y(_0407_),
    .A1(_1785_),
    .A2(\MemCell.dc2_reg[2][0] ));
 sg13g2_a221oi_1 _2634_ (.B2(\MemCell.dc2_reg[2][4] ),
    .C1(_0407_),
    .B1(_1923_),
    .A1(_1785_),
    .Y(_0408_),
    .A2(\MemCell.dc2_reg[2][0] ));
 sg13g2_nand4_1 _2635_ (.B(_0403_),
    .C(_0405_),
    .A(_0402_),
    .Y(_0409_),
    .D(_0408_));
 sg13g2_or4_1 _2636_ (.A(_0391_),
    .B(_0396_),
    .C(_0401_),
    .D(_0409_),
    .X(_0410_));
 sg13g2_a21oi_2 _2637_ (.B1(_0410_),
    .Y(_0411_),
    .A2(_1978_),
    .A1(_1976_));
 sg13g2_o21ai_1 _2638_ (.B1(_1982_),
    .Y(_0412_),
    .A1(_1983_),
    .A2(_1995_));
 sg13g2_a22oi_1 _2639_ (.Y(_0413_),
    .B1(_1991_),
    .B2(_0412_),
    .A2(_1989_),
    .A1(_1988_));
 sg13g2_o21ai_1 _2640_ (.B1(_1986_),
    .Y(_0414_),
    .A1(_1992_),
    .A2(_0413_));
 sg13g2_a21oi_1 _2641_ (.A1(_1994_),
    .A2(_0414_),
    .Y(_0415_),
    .B1(_1980_));
 sg13g2_nor2b_1 _2642_ (.A(_0396_),
    .B_N(_0403_),
    .Y(_0416_));
 sg13g2_a22oi_1 _2643_ (.Y(_0417_),
    .B1(_0407_),
    .B2(_0416_),
    .A2(_0395_),
    .A1(_0393_));
 sg13g2_o21ai_1 _2644_ (.B1(_0405_),
    .Y(_0418_),
    .A1(_0404_),
    .A2(_0417_));
 sg13g2_nor2b_1 _2645_ (.A(_0401_),
    .B_N(_0402_),
    .Y(_0419_));
 sg13g2_a22oi_1 _2646_ (.Y(_0420_),
    .B1(_0418_),
    .B2(_0419_),
    .A2(_0399_),
    .A1(_0398_));
 sg13g2_nor2_1 _2647_ (.A(_0391_),
    .B(_0420_),
    .Y(_0421_));
 sg13g2_nor2b_1 _2648_ (.A(_1979_),
    .B_N(\MemCell.enable_pwm ),
    .Y(_0422_));
 sg13g2_o21ai_1 _2649_ (.B1(_0422_),
    .Y(_0423_),
    .A1(_1985_),
    .A2(_0415_));
 sg13g2_nor3_2 _2650_ (.A(_0411_),
    .B(_0421_),
    .C(_0423_),
    .Y(_0097_));
 sg13g2_nand2b_1 _2651_ (.Y(_0424_),
    .B(\pwm_module.counter2[15] ),
    .A_N(\MemCell.dc3_reg[1][7] ));
 sg13g2_o21ai_1 _2652_ (.B1(_0424_),
    .Y(_0425_),
    .A1(\MemCell.dc3_reg[1][6] ),
    .A2(_1825_));
 sg13g2_nand2_1 _2653_ (.Y(_0426_),
    .A(\MemCell.dc3_reg[1][7] ),
    .B(_1823_));
 sg13g2_o21ai_1 _2654_ (.B1(_0426_),
    .Y(_0427_),
    .A1(_1824_),
    .A2(\pwm_module.counter2[14] ));
 sg13g2_a22oi_1 _2655_ (.Y(_0428_),
    .B1(_1828_),
    .B2(\pwm_module.counter2[12] ),
    .A2(\pwm_module.counter2[13] ),
    .A1(_1826_));
 sg13g2_nor2_1 _2656_ (.A(_1826_),
    .B(\pwm_module.counter2[13] ),
    .Y(_0429_));
 sg13g2_nand2b_1 _2657_ (.Y(_0430_),
    .B(net649),
    .A_N(\MemCell.dc3_reg[0][1] ));
 sg13g2_nor2b_1 _2658_ (.A(\pwm_module.counter2[0] ),
    .B_N(\MemCell.dc3_reg[0][0] ),
    .Y(_0431_));
 sg13g2_nor2b_1 _2659_ (.A(net649),
    .B_N(\MemCell.dc3_reg[0][1] ),
    .Y(_0432_));
 sg13g2_a221oi_1 _2660_ (.B2(_0431_),
    .C1(_0432_),
    .B1(_0430_),
    .A1(\MemCell.dc3_reg[0][2] ),
    .Y(_0433_),
    .A2(_1842_));
 sg13g2_nand2b_1 _2661_ (.Y(_0434_),
    .B(\pwm_module.counter2[2] ),
    .A_N(\MemCell.dc3_reg[0][2] ));
 sg13g2_o21ai_1 _2662_ (.B1(_0434_),
    .Y(_0435_),
    .A1(\MemCell.dc3_reg[0][3] ),
    .A2(_1841_));
 sg13g2_a22oi_1 _2663_ (.Y(_0436_),
    .B1(\MemCell.dc3_reg[0][3] ),
    .B2(_1841_),
    .A2(\MemCell.dc3_reg[0][4] ),
    .A1(_1839_));
 sg13g2_o21ai_1 _2664_ (.B1(_0436_),
    .Y(_0437_),
    .A1(_0433_),
    .A2(_0435_));
 sg13g2_a22oi_1 _2665_ (.Y(_0438_),
    .B1(\pwm_module.counter2[4] ),
    .B2(_1840_),
    .A2(\pwm_module.counter2[5] ),
    .A1(_1837_));
 sg13g2_nor2_1 _2666_ (.A(_1837_),
    .B(\pwm_module.counter2[5] ),
    .Y(_0439_));
 sg13g2_a221oi_1 _2667_ (.B2(_0438_),
    .C1(_0439_),
    .B1(_0437_),
    .A1(\MemCell.dc3_reg[0][6] ),
    .Y(_0440_),
    .A2(_1836_));
 sg13g2_nand2b_1 _2668_ (.Y(_0441_),
    .B(\pwm_module.counter2[7] ),
    .A_N(\MemCell.dc3_reg[0][7] ));
 sg13g2_o21ai_1 _2669_ (.B1(_0441_),
    .Y(_0442_),
    .A1(\MemCell.dc3_reg[0][6] ),
    .A2(_1836_));
 sg13g2_a22oi_1 _2670_ (.Y(_0443_),
    .B1(\MemCell.dc3_reg[0][7] ),
    .B2(_1835_),
    .A2(_1834_),
    .A1(\MemCell.dc3_reg[1][0] ));
 sg13g2_o21ai_1 _2671_ (.B1(_0443_),
    .Y(_0444_),
    .A1(_0440_),
    .A2(_0442_));
 sg13g2_a22oi_1 _2672_ (.Y(_0445_),
    .B1(_1833_),
    .B2(\pwm_module.counter2[8] ),
    .A2(\pwm_module.counter2[9] ),
    .A1(_1831_));
 sg13g2_nor2b_1 _2673_ (.A(\pwm_module.counter2[10] ),
    .B_N(\MemCell.dc3_reg[1][2] ),
    .Y(_0446_));
 sg13g2_a221oi_1 _2674_ (.B2(_0445_),
    .C1(_0446_),
    .B1(_0444_),
    .A1(\MemCell.dc3_reg[1][1] ),
    .Y(_0447_),
    .A2(_1832_));
 sg13g2_nand2b_1 _2675_ (.Y(_0448_),
    .B(\pwm_module.counter2[11] ),
    .A_N(\MemCell.dc3_reg[1][3] ));
 sg13g2_o21ai_1 _2676_ (.B1(_0448_),
    .Y(_0449_),
    .A1(\MemCell.dc3_reg[1][2] ),
    .A2(_1830_));
 sg13g2_nand2b_1 _2677_ (.Y(_0450_),
    .B(\MemCell.dc3_reg[1][3] ),
    .A_N(\pwm_module.counter2[11] ));
 sg13g2_a21oi_1 _2678_ (.A1(\MemCell.dc3_reg[1][4] ),
    .A2(_1829_),
    .Y(_0451_),
    .B1(_0429_));
 sg13g2_nand3_1 _2679_ (.B(_0450_),
    .C(_0451_),
    .A(_0428_),
    .Y(_0452_));
 sg13g2_nor3_1 _2680_ (.A(_0425_),
    .B(_0427_),
    .C(_0452_),
    .Y(_0453_));
 sg13g2_o21ai_1 _2681_ (.B1(_0453_),
    .Y(_0454_),
    .A1(_0447_),
    .A2(_0449_));
 sg13g2_nor4_1 _2682_ (.A(_0425_),
    .B(_0427_),
    .C(_0428_),
    .D(_0429_),
    .Y(_0455_));
 sg13g2_a21oi_1 _2683_ (.A1(_0425_),
    .A2(_0426_),
    .Y(_0456_),
    .B1(_0455_));
 sg13g2_nand2b_1 _2684_ (.Y(_0457_),
    .B(\pwm_module.counter2[27] ),
    .A_N(\MemCell.dc3_reg[3][3] ));
 sg13g2_o21ai_1 _2685_ (.B1(_0457_),
    .Y(_0458_),
    .A1(\MemCell.dc3_reg[3][2] ),
    .A2(_1812_));
 sg13g2_nand2_1 _2686_ (.Y(_0459_),
    .A(\MemCell.dc3_reg[3][2] ),
    .B(_1812_));
 sg13g2_nand2b_1 _2687_ (.Y(_0460_),
    .B(net85),
    .A_N(\pwm_module.counter2[27] ));
 sg13g2_nand3b_1 _2688_ (.B(_0459_),
    .C(_0460_),
    .Y(_0461_),
    .A_N(_0458_));
 sg13g2_nand2b_1 _2689_ (.Y(_0462_),
    .B(\pwm_module.counter2[22] ),
    .A_N(\MemCell.dc3_reg[2][6] ));
 sg13g2_o21ai_1 _2690_ (.B1(_0462_),
    .Y(_0463_),
    .A1(_1818_),
    .A2(\pwm_module.counter2[21] ));
 sg13g2_nor2b_1 _2691_ (.A(\pwm_module.counter2[23] ),
    .B_N(\MemCell.dc3_reg[2][7] ),
    .Y(_0464_));
 sg13g2_a221oi_1 _2692_ (.B2(_1817_),
    .C1(_0463_),
    .B1(\MemCell.dc3_reg[2][6] ),
    .A1(\MemCell.dc3_reg[2][7] ),
    .Y(_0465_),
    .A2(_1816_));
 sg13g2_nand2b_1 _2693_ (.Y(_0466_),
    .B(\pwm_module.counter2[18] ),
    .A_N(\MemCell.dc3_reg[2][2] ));
 sg13g2_nor2b_1 _2694_ (.A(\pwm_module.counter2[19] ),
    .B_N(\MemCell.dc3_reg[2][3] ),
    .Y(_0467_));
 sg13g2_xor2_1 _2695_ (.B(\pwm_module.counter2[18] ),
    .A(\MemCell.dc3_reg[2][2] ),
    .X(_0468_));
 sg13g2_nor2_1 _2696_ (.A(_0467_),
    .B(_0468_),
    .Y(_0469_));
 sg13g2_nor2b_1 _2697_ (.A(_0461_),
    .B_N(_0469_),
    .Y(_0470_));
 sg13g2_a22oi_1 _2698_ (.Y(_0471_),
    .B1(_1806_),
    .B2(\pwm_module.counter2[30] ),
    .A2(_1805_),
    .A1(\pwm_module.counter2[31] ));
 sg13g2_a22oi_1 _2699_ (.Y(_0472_),
    .B1(\pwm_module.counter2[28] ),
    .B2(_1811_),
    .A2(\pwm_module.counter2[29] ),
    .A1(_1808_));
 sg13g2_nand2_1 _2700_ (.Y(_0473_),
    .A(_0471_),
    .B(_0472_));
 sg13g2_nand2b_1 _2701_ (.Y(_0474_),
    .B(net146),
    .A_N(net179));
 sg13g2_o21ai_1 _2702_ (.B1(_0474_),
    .Y(_0475_),
    .A1(\pwm_module.counter2[28] ),
    .A2(_1811_));
 sg13g2_nand2_1 _2703_ (.Y(_0476_),
    .A(\MemCell.dc3_reg[3][5] ),
    .B(_1809_));
 sg13g2_o21ai_1 _2704_ (.B1(_0476_),
    .Y(_0477_),
    .A1(_1806_),
    .A2(\pwm_module.counter2[30] ));
 sg13g2_nor3_1 _2705_ (.A(_0473_),
    .B(_0475_),
    .C(_0477_),
    .Y(_0478_));
 sg13g2_nand2b_1 _2706_ (.Y(_0479_),
    .B(\pwm_module.counter2[16] ),
    .A_N(\MemCell.dc3_reg[2][0] ));
 sg13g2_nand2b_1 _2707_ (.Y(_0480_),
    .B(\pwm_module.counter2[17] ),
    .A_N(\MemCell.dc3_reg[2][1] ));
 sg13g2_a22oi_1 _2708_ (.Y(_0481_),
    .B1(_1819_),
    .B2(\pwm_module.counter2[20] ),
    .A2(\pwm_module.counter2[21] ),
    .A1(_1818_));
 sg13g2_a22oi_1 _2709_ (.Y(_0482_),
    .B1(_1815_),
    .B2(\pwm_module.counter2[24] ),
    .A2(\pwm_module.counter2[25] ),
    .A1(_1813_));
 sg13g2_nand4_1 _2710_ (.B(_0480_),
    .C(_0481_),
    .A(_0479_),
    .Y(_0483_),
    .D(_0482_));
 sg13g2_nor2b_1 _2711_ (.A(net648),
    .B_N(\MemCell.dc3_reg[2][1] ),
    .Y(_0484_));
 sg13g2_nand2b_1 _2712_ (.Y(_0485_),
    .B(\pwm_module.counter2[19] ),
    .A_N(\MemCell.dc3_reg[2][3] ));
 sg13g2_nor2b_1 _2713_ (.A(\pwm_module.counter2[16] ),
    .B_N(\MemCell.dc3_reg[2][0] ),
    .Y(_0486_));
 sg13g2_nor2_1 _2714_ (.A(_1815_),
    .B(\pwm_module.counter2[24] ),
    .Y(_0487_));
 sg13g2_nand2b_1 _2715_ (.Y(_0488_),
    .B(\pwm_module.counter2[23] ),
    .A_N(\MemCell.dc3_reg[2][7] ));
 sg13g2_nand2_1 _2716_ (.Y(_0489_),
    .A(\MemCell.dc3_reg[3][1] ),
    .B(_1814_));
 sg13g2_nor2_1 _2717_ (.A(_1819_),
    .B(\pwm_module.counter2[20] ),
    .Y(_0490_));
 sg13g2_nor4_1 _2718_ (.A(_0484_),
    .B(_0486_),
    .C(_0487_),
    .D(_0490_),
    .Y(_0491_));
 sg13g2_nand4_1 _2719_ (.B(_0488_),
    .C(_0489_),
    .A(_0485_),
    .Y(_0492_),
    .D(_0491_));
 sg13g2_nor2_1 _2720_ (.A(_0483_),
    .B(_0492_),
    .Y(_0493_));
 sg13g2_nand4_1 _2721_ (.B(_0470_),
    .C(_0478_),
    .A(_0465_),
    .Y(_0494_),
    .D(_0493_));
 sg13g2_a21oi_2 _2722_ (.B1(_0494_),
    .Y(_0495_),
    .A2(_0456_),
    .A1(_0454_));
 sg13g2_o21ai_1 _2723_ (.B1(_0485_),
    .Y(_0496_),
    .A1(_0466_),
    .A2(_0467_));
 sg13g2_a21oi_1 _2724_ (.A1(_0479_),
    .A2(_0480_),
    .Y(_0497_),
    .B1(_0484_));
 sg13g2_a21oi_1 _2725_ (.A1(_0469_),
    .A2(_0497_),
    .Y(_0498_),
    .B1(_0496_));
 sg13g2_o21ai_1 _2726_ (.B1(_0481_),
    .Y(_0499_),
    .A1(_0490_),
    .A2(_0498_));
 sg13g2_o21ai_1 _2727_ (.B1(_0488_),
    .Y(_0500_),
    .A1(_0462_),
    .A2(_0464_));
 sg13g2_a21oi_1 _2728_ (.A1(_0465_),
    .A2(_0499_),
    .Y(_0501_),
    .B1(_0500_));
 sg13g2_o21ai_1 _2729_ (.B1(_0482_),
    .Y(_0502_),
    .A1(_0487_),
    .A2(_0501_));
 sg13g2_nor2b_1 _2730_ (.A(_0461_),
    .B_N(_0489_),
    .Y(_0503_));
 sg13g2_a22oi_1 _2731_ (.Y(_0504_),
    .B1(_0502_),
    .B2(_0503_),
    .A2(_0460_),
    .A1(_0458_));
 sg13g2_nor2b_1 _2732_ (.A(_0504_),
    .B_N(_0478_),
    .Y(_0505_));
 sg13g2_o21ai_1 _2733_ (.B1(_0471_),
    .Y(_0506_),
    .A1(_0472_),
    .A2(_0477_));
 sg13g2_nand2_1 _2734_ (.Y(_0507_),
    .A(_0474_),
    .B(_0506_));
 sg13g2_nand2_1 _2735_ (.Y(_0508_),
    .A(net405),
    .B(_0507_));
 sg13g2_nor3_1 _2736_ (.A(_0495_),
    .B(_0505_),
    .C(_0508_),
    .Y(_0098_));
 sg13g2_xor2_1 _2737_ (.B(\spi_module.r_RX_Bit_Count[0] ),
    .A(\spi_module.r_RX_Bit_Count[1] ),
    .X(_0100_));
 sg13g2_a21o_1 _2738_ (.A2(\spi_module.r_RX_Bit_Count[0] ),
    .A1(\spi_module.r_RX_Bit_Count[1] ),
    .B1(\spi_module.r_RX_Bit_Count[2] ),
    .X(_0509_));
 sg13g2_and2_1 _2739_ (.A(_1945_),
    .B(_0509_),
    .X(_0101_));
 sg13g2_nor2b_1 _2740_ (.A(net436),
    .B_N(net38),
    .Y(_0099_));
 sg13g2_nand2b_1 _2741_ (.Y(_0510_),
    .B(\pwm_module.prescaler0[1] ),
    .A_N(\MemCell.prescale_reg[0][1] ));
 sg13g2_nor2b_1 _2742_ (.A(\pwm_module.prescaler0[0] ),
    .B_N(\MemCell.prescale_reg[0][0] ),
    .Y(_0511_));
 sg13g2_nor2b_1 _2743_ (.A(\pwm_module.prescaler0[1] ),
    .B_N(\MemCell.prescale_reg[0][1] ),
    .Y(_0512_));
 sg13g2_a221oi_1 _2744_ (.B2(_0511_),
    .C1(_0512_),
    .B1(_0510_),
    .A1(\MemCell.prescale_reg[0][2] ),
    .Y(_0513_),
    .A2(_1871_));
 sg13g2_nand2_1 _2745_ (.Y(_0514_),
    .A(_1847_),
    .B(\pwm_module.prescaler0[3] ));
 sg13g2_nand2_1 _2746_ (.Y(_0515_),
    .A(_1849_),
    .B(\pwm_module.prescaler0[2] ));
 sg13g2_nand3b_1 _2747_ (.B(_0514_),
    .C(_0515_),
    .Y(_0516_),
    .A_N(_0513_));
 sg13g2_nand2b_1 _2748_ (.Y(_0517_),
    .B(\pwm_module.prescaler0[7] ),
    .A_N(\MemCell.prescale_reg[0][7] ));
 sg13g2_o21ai_1 _2749_ (.B1(_0517_),
    .Y(_0518_),
    .A1(\MemCell.prescale_reg[0][6] ),
    .A2(_1870_));
 sg13g2_nor2b_1 _2750_ (.A(\MemCell.prescale_reg[0][5] ),
    .B_N(\pwm_module.prescaler0[5] ),
    .Y(_0519_));
 sg13g2_a21o_1 _2751_ (.A2(\pwm_module.prescaler0[4] ),
    .A1(_1850_),
    .B1(_0519_),
    .X(_0520_));
 sg13g2_nand2b_1 _2752_ (.Y(_0521_),
    .B(\MemCell.prescale_reg[0][7] ),
    .A_N(\pwm_module.prescaler0[7] ));
 sg13g2_nand2b_1 _2753_ (.Y(_0522_),
    .B(\MemCell.prescale_reg[0][3] ),
    .A_N(\pwm_module.prescaler0[3] ));
 sg13g2_nand2b_1 _2754_ (.Y(_0523_),
    .B(\MemCell.prescale_reg[0][4] ),
    .A_N(\pwm_module.prescaler0[4] ));
 sg13g2_nand3_1 _2755_ (.B(_0522_),
    .C(_0523_),
    .A(_0521_),
    .Y(_0524_));
 sg13g2_nor2b_1 _2756_ (.A(\pwm_module.prescaler0[5] ),
    .B_N(\MemCell.prescale_reg[0][5] ),
    .Y(_0525_));
 sg13g2_a21oi_1 _2757_ (.A1(\MemCell.prescale_reg[0][6] ),
    .A2(_1870_),
    .Y(_0526_),
    .B1(_0525_));
 sg13g2_a21o_1 _2758_ (.A2(_1870_),
    .A1(\MemCell.prescale_reg[0][6] ),
    .B1(_0525_),
    .X(_0527_));
 sg13g2_nor4_1 _2759_ (.A(_0518_),
    .B(_0520_),
    .C(_0524_),
    .D(_0527_),
    .Y(_0528_));
 sg13g2_a21o_1 _2760_ (.A2(_0526_),
    .A1(_0520_),
    .B1(_0518_),
    .X(_0529_));
 sg13g2_a22oi_1 _2761_ (.Y(_0530_),
    .B1(_0529_),
    .B2(_0521_),
    .A2(_0528_),
    .A1(_0516_));
 sg13g2_nand2b_1 _2762_ (.Y(_0531_),
    .B(\pwm_module.prescaler0[15] ),
    .A_N(\MemCell.prescale_reg[1][7] ));
 sg13g2_nand2b_1 _2763_ (.Y(_0532_),
    .B(\pwm_module.prescaler0[14] ),
    .A_N(\MemCell.prescale_reg[1][6] ));
 sg13g2_nor2b_1 _2764_ (.A(\pwm_module.prescaler0[15] ),
    .B_N(\MemCell.prescale_reg[1][7] ),
    .Y(_0533_));
 sg13g2_nand2b_1 _2765_ (.Y(_0534_),
    .B(\MemCell.prescale_reg[1][7] ),
    .A_N(\pwm_module.prescaler0[15] ));
 sg13g2_nand2b_1 _2766_ (.Y(_0535_),
    .B(\MemCell.prescale_reg[1][6] ),
    .A_N(\pwm_module.prescaler0[14] ));
 sg13g2_nor2b_1 _2767_ (.A(\pwm_module.prescaler0[13] ),
    .B_N(\MemCell.prescale_reg[1][5] ),
    .Y(_0536_));
 sg13g2_nand4_1 _2768_ (.B(_0532_),
    .C(_0534_),
    .A(_0531_),
    .Y(_0537_),
    .D(_0535_));
 sg13g2_nor2_1 _2769_ (.A(_0536_),
    .B(_0537_),
    .Y(_0538_));
 sg13g2_nand2b_1 _2770_ (.Y(_0539_),
    .B(\pwm_module.prescaler0[12] ),
    .A_N(\MemCell.prescale_reg[1][4] ));
 sg13g2_o21ai_1 _2771_ (.B1(_0539_),
    .Y(_0540_),
    .A1(\MemCell.prescale_reg[1][5] ),
    .A2(_1869_));
 sg13g2_nor2b_1 _2772_ (.A(\pwm_module.prescaler0[12] ),
    .B_N(\MemCell.prescale_reg[1][4] ),
    .Y(_0541_));
 sg13g2_nor4_1 _2773_ (.A(_0536_),
    .B(_0537_),
    .C(_0540_),
    .D(_0541_),
    .Y(_0542_));
 sg13g2_nand2b_1 _2774_ (.Y(_0543_),
    .B(\pwm_module.prescaler0[11] ),
    .A_N(net652));
 sg13g2_nand2b_1 _2775_ (.Y(_0544_),
    .B(\pwm_module.prescaler0[10] ),
    .A_N(\MemCell.prescale_reg[1][2] ));
 sg13g2_nand2b_1 _2776_ (.Y(_0545_),
    .B(\MemCell.prescale_reg[1][2] ),
    .A_N(\pwm_module.prescaler0[10] ));
 sg13g2_nor2b_1 _2777_ (.A(\pwm_module.prescaler0[11] ),
    .B_N(net652),
    .Y(_0546_));
 sg13g2_nand2b_1 _2778_ (.Y(_0547_),
    .B(net652),
    .A_N(\pwm_module.prescaler0[11] ));
 sg13g2_and4_1 _2779_ (.A(_0543_),
    .B(_0544_),
    .C(_0545_),
    .D(_0547_),
    .X(_0548_));
 sg13g2_nand2b_1 _2780_ (.Y(_0549_),
    .B(\pwm_module.prescaler0[8] ),
    .A_N(\MemCell.prescale_reg[1][0] ));
 sg13g2_nand2b_1 _2781_ (.Y(_0550_),
    .B(\pwm_module.prescaler0[9] ),
    .A_N(\MemCell.prescale_reg[1][1] ));
 sg13g2_nand2_1 _2782_ (.Y(_0551_),
    .A(_0549_),
    .B(_0550_));
 sg13g2_nor2b_1 _2783_ (.A(\pwm_module.prescaler0[9] ),
    .B_N(\MemCell.prescale_reg[1][1] ),
    .Y(_0552_));
 sg13g2_nand2b_1 _2784_ (.Y(_0553_),
    .B(\MemCell.prescale_reg[1][0] ),
    .A_N(\pwm_module.prescaler0[8] ));
 sg13g2_nor2_1 _2785_ (.A(_0551_),
    .B(_0552_),
    .Y(_0554_));
 sg13g2_nand4_1 _2786_ (.B(_0548_),
    .C(_0553_),
    .A(_0542_),
    .Y(_0555_),
    .D(_0554_));
 sg13g2_a21oi_1 _2787_ (.A1(_0543_),
    .A2(_0544_),
    .Y(_0556_),
    .B1(_0546_));
 sg13g2_a21oi_1 _2788_ (.A1(_0549_),
    .A2(_0550_),
    .Y(_0557_),
    .B1(_0552_));
 sg13g2_a21o_1 _2789_ (.A2(_0557_),
    .A1(_0548_),
    .B1(_0556_),
    .X(_0558_));
 sg13g2_a21oi_1 _2790_ (.A1(_0531_),
    .A2(_0532_),
    .Y(_0559_),
    .B1(_0533_));
 sg13g2_a221oi_1 _2791_ (.B2(_0558_),
    .C1(_0559_),
    .B1(_0542_),
    .A1(_0538_),
    .Y(_0560_),
    .A2(_0540_));
 sg13g2_o21ai_1 _2792_ (.B1(_0560_),
    .Y(_0561_),
    .A1(_0530_),
    .A2(_0555_));
 sg13g2_nor2b_1 _2793_ (.A(\MemCell.prescale_reg[3][7] ),
    .B_N(\pwm_module.prescaler0[31] ),
    .Y(_0562_));
 sg13g2_a21o_1 _2794_ (.A2(\pwm_module.prescaler0[30] ),
    .A1(_1855_),
    .B1(_0562_),
    .X(_0563_));
 sg13g2_nor2b_1 _2795_ (.A(\MemCell.prescale_reg[3][5] ),
    .B_N(\pwm_module.prescaler0[29] ),
    .Y(_0564_));
 sg13g2_a21o_1 _2796_ (.A2(\pwm_module.prescaler0[28] ),
    .A1(_1856_),
    .B1(_0564_),
    .X(_0565_));
 sg13g2_nand2b_1 _2797_ (.Y(_0566_),
    .B(\MemCell.prescale_reg[3][7] ),
    .A_N(\pwm_module.prescaler0[31] ));
 sg13g2_o21ai_1 _2798_ (.B1(_0566_),
    .Y(_0567_),
    .A1(_1856_),
    .A2(\pwm_module.prescaler0[28] ));
 sg13g2_nand2b_1 _2799_ (.Y(_0568_),
    .B(\MemCell.prescale_reg[3][5] ),
    .A_N(\pwm_module.prescaler0[29] ));
 sg13g2_o21ai_1 _2800_ (.B1(_0568_),
    .Y(_0569_),
    .A1(_1855_),
    .A2(\pwm_module.prescaler0[30] ));
 sg13g2_nor4_2 _2801_ (.A(_0563_),
    .B(_0565_),
    .C(_0567_),
    .Y(_0570_),
    .D(_0569_));
 sg13g2_nor2b_1 _2802_ (.A(\MemCell.prescale_reg[3][2] ),
    .B_N(\pwm_module.prescaler0[26] ),
    .Y(_0571_));
 sg13g2_a21oi_1 _2803_ (.A1(_1857_),
    .A2(\pwm_module.prescaler0[27] ),
    .Y(_0572_),
    .B1(_0571_));
 sg13g2_a22oi_1 _2804_ (.Y(_0573_),
    .B1(\pwm_module.prescaler0[24] ),
    .B2(_1859_),
    .A2(\pwm_module.prescaler0[25] ),
    .A1(_1858_));
 sg13g2_and2_1 _2805_ (.A(_0572_),
    .B(_0573_),
    .X(_0574_));
 sg13g2_nand2b_1 _2806_ (.Y(_0575_),
    .B(\MemCell.prescale_reg[3][2] ),
    .A_N(\pwm_module.prescaler0[26] ));
 sg13g2_nand2b_1 _2807_ (.Y(_0576_),
    .B(\MemCell.prescale_reg[3][1] ),
    .A_N(\pwm_module.prescaler0[25] ));
 sg13g2_nand2_1 _2808_ (.Y(_0577_),
    .A(_0575_),
    .B(_0576_));
 sg13g2_nor2b_1 _2809_ (.A(\pwm_module.prescaler0[24] ),
    .B_N(\MemCell.prescale_reg[3][0] ),
    .Y(_0578_));
 sg13g2_nor2_1 _2810_ (.A(_1857_),
    .B(\pwm_module.prescaler0[27] ),
    .Y(_0579_));
 sg13g2_nor3_1 _2811_ (.A(_0577_),
    .B(_0578_),
    .C(_0579_),
    .Y(_0580_));
 sg13g2_nand3_1 _2812_ (.B(_0574_),
    .C(_0580_),
    .A(_0570_),
    .Y(_0581_));
 sg13g2_nor2b_1 _2813_ (.A(net653),
    .B_N(\pwm_module.prescaler0[19] ),
    .Y(_0582_));
 sg13g2_nor2b_1 _2814_ (.A(\MemCell.prescale_reg[2][2] ),
    .B_N(\pwm_module.prescaler0[18] ),
    .Y(_0583_));
 sg13g2_nor2b_1 _2815_ (.A(\pwm_module.prescaler0[18] ),
    .B_N(\MemCell.prescale_reg[2][2] ),
    .Y(_0584_));
 sg13g2_nor2b_1 _2816_ (.A(\pwm_module.prescaler0[19] ),
    .B_N(net653),
    .Y(_0585_));
 sg13g2_nand2b_1 _2817_ (.Y(_0586_),
    .B(net653),
    .A_N(\pwm_module.prescaler0[19] ));
 sg13g2_or4_1 _2818_ (.A(_0582_),
    .B(_0583_),
    .C(_0584_),
    .D(_0585_),
    .X(_0587_));
 sg13g2_nand2b_1 _2819_ (.Y(_0588_),
    .B(\pwm_module.prescaler0[16] ),
    .A_N(\MemCell.prescale_reg[2][0] ));
 sg13g2_nand2b_1 _2820_ (.Y(_0589_),
    .B(\pwm_module.prescaler0[17] ),
    .A_N(\MemCell.prescale_reg[2][1] ));
 sg13g2_nand2_1 _2821_ (.Y(_0590_),
    .A(_0588_),
    .B(_0589_));
 sg13g2_nor2b_1 _2822_ (.A(\pwm_module.prescaler0[17] ),
    .B_N(\MemCell.prescale_reg[2][1] ),
    .Y(_0591_));
 sg13g2_nand2b_1 _2823_ (.Y(_0592_),
    .B(\pwm_module.prescaler0[23] ),
    .A_N(\MemCell.prescale_reg[2][7] ));
 sg13g2_nand2b_1 _2824_ (.Y(_0593_),
    .B(\pwm_module.prescaler0[22] ),
    .A_N(\MemCell.prescale_reg[2][6] ));
 sg13g2_nand2_1 _2825_ (.Y(_0594_),
    .A(_0592_),
    .B(_0593_));
 sg13g2_nand2b_1 _2826_ (.Y(_0595_),
    .B(\MemCell.prescale_reg[2][6] ),
    .A_N(\pwm_module.prescaler0[22] ));
 sg13g2_nand2b_1 _2827_ (.Y(_0596_),
    .B(\MemCell.prescale_reg[2][7] ),
    .A_N(\pwm_module.prescaler0[23] ));
 sg13g2_and4_1 _2828_ (.A(_0592_),
    .B(_0593_),
    .C(_0595_),
    .D(_0596_),
    .X(_0597_));
 sg13g2_a22oi_1 _2829_ (.Y(_0598_),
    .B1(\pwm_module.prescaler0[20] ),
    .B2(_1862_),
    .A2(\pwm_module.prescaler0[21] ),
    .A1(_1860_));
 sg13g2_nor2b_1 _2830_ (.A(\pwm_module.prescaler0[21] ),
    .B_N(\MemCell.prescale_reg[2][5] ),
    .Y(_0599_));
 sg13g2_a21oi_1 _2831_ (.A1(\MemCell.prescale_reg[2][4] ),
    .A2(_1867_),
    .Y(_0600_),
    .B1(_0599_));
 sg13g2_and3_1 _2832_ (.X(_0601_),
    .A(_0597_),
    .B(_0598_),
    .C(_0600_));
 sg13g2_a21oi_1 _2833_ (.A1(\MemCell.prescale_reg[2][0] ),
    .A2(_1868_),
    .Y(_0602_),
    .B1(_0587_));
 sg13g2_nand2_1 _2834_ (.Y(_0603_),
    .A(_0601_),
    .B(_0602_));
 sg13g2_nor4_1 _2835_ (.A(_0581_),
    .B(_0590_),
    .C(_0591_),
    .D(_0603_),
    .Y(_0604_));
 sg13g2_o21ai_1 _2836_ (.B1(_0586_),
    .Y(_0605_),
    .A1(_0582_),
    .A2(_0583_));
 sg13g2_a21o_1 _2837_ (.A2(_0589_),
    .A1(_0588_),
    .B1(_0591_),
    .X(_0606_));
 sg13g2_o21ai_1 _2838_ (.B1(_0605_),
    .Y(_0607_),
    .A1(_0587_),
    .A2(_0606_));
 sg13g2_and2_1 _2839_ (.A(_0594_),
    .B(_0596_),
    .X(_0608_));
 sg13g2_nor2_1 _2840_ (.A(_0598_),
    .B(_0599_),
    .Y(_0609_));
 sg13g2_a221oi_1 _2841_ (.B2(_0597_),
    .C1(_0608_),
    .B1(_0609_),
    .A1(_0601_),
    .Y(_0610_),
    .A2(_0607_));
 sg13g2_nor2b_1 _2842_ (.A(_0569_),
    .B_N(_0565_),
    .Y(_0611_));
 sg13g2_o21ai_1 _2843_ (.B1(_0566_),
    .Y(_0612_),
    .A1(_0563_),
    .A2(_0611_));
 sg13g2_a221oi_1 _2844_ (.B2(_0576_),
    .C1(_0571_),
    .B1(_0575_),
    .A1(_1857_),
    .Y(_0613_),
    .A2(\pwm_module.prescaler0[27] ));
 sg13g2_nor3_1 _2845_ (.A(_0574_),
    .B(_0579_),
    .C(_0613_),
    .Y(_0614_));
 sg13g2_o21ai_1 _2846_ (.B1(_0612_),
    .Y(_0615_),
    .A1(_0581_),
    .A2(_0610_));
 sg13g2_a221oi_1 _2847_ (.B2(_0570_),
    .C1(_0615_),
    .B1(_0614_),
    .A1(_0561_),
    .Y(_0616_),
    .A2(_0604_));
 sg13g2_nand2_2 _2848_ (.Y(_0617_),
    .A(net651),
    .B(_0616_));
 sg13g2_nor2_1 _2849_ (.A(net96),
    .B(net607),
    .Y(_0000_));
 sg13g2_xnor2_1 _2850_ (.Y(_0618_),
    .A(net382),
    .B(net96));
 sg13g2_nor2_1 _2851_ (.A(net607),
    .B(_0618_),
    .Y(_0011_));
 sg13g2_and3_1 _2852_ (.X(_0619_),
    .A(net114),
    .B(net554),
    .C(net96));
 sg13g2_a21oi_1 _2853_ (.A1(\pwm_module.prescaler0[1] ),
    .A2(net96),
    .Y(_0620_),
    .B1(net114));
 sg13g2_nor3_1 _2854_ (.A(net607),
    .B(_0619_),
    .C(net115),
    .Y(_0022_));
 sg13g2_and2_1 _2855_ (.A(net252),
    .B(_0619_),
    .X(_0621_));
 sg13g2_nand4_1 _2856_ (.B(\pwm_module.prescaler0[2] ),
    .C(\pwm_module.prescaler0[1] ),
    .A(\pwm_module.prescaler0[3] ),
    .Y(_0622_),
    .D(\pwm_module.prescaler0[0] ));
 sg13g2_nor2_1 _2857_ (.A(net252),
    .B(_0619_),
    .Y(_0623_));
 sg13g2_nor3_1 _2858_ (.A(net607),
    .B(_0621_),
    .C(net253),
    .Y(_0025_));
 sg13g2_nor2_1 _2859_ (.A(net325),
    .B(_0621_),
    .Y(_0624_));
 sg13g2_and2_1 _2860_ (.A(net325),
    .B(_0621_),
    .X(_0625_));
 sg13g2_nor3_1 _2861_ (.A(net607),
    .B(_0624_),
    .C(_0625_),
    .Y(_0026_));
 sg13g2_nor2_1 _2862_ (.A(net261),
    .B(_0625_),
    .Y(_0626_));
 sg13g2_nand2_2 _2863_ (.Y(_0627_),
    .A(net261),
    .B(net325));
 sg13g2_nor2_1 _2864_ (.A(_0622_),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_nor3_1 _2865_ (.A(net607),
    .B(net262),
    .C(_0628_),
    .Y(_0027_));
 sg13g2_xnor2_1 _2866_ (.Y(_0629_),
    .A(net258),
    .B(_0628_));
 sg13g2_nor2_1 _2867_ (.A(net607),
    .B(net259),
    .Y(_0028_));
 sg13g2_a21oi_1 _2868_ (.A1(\pwm_module.prescaler0[6] ),
    .A2(_0628_),
    .Y(_0630_),
    .B1(net116));
 sg13g2_nand2_1 _2869_ (.Y(_0631_),
    .A(net116),
    .B(net258));
 sg13g2_nor3_2 _2870_ (.A(_0622_),
    .B(_0627_),
    .C(_0631_),
    .Y(_0632_));
 sg13g2_nor3_1 _2871_ (.A(net608),
    .B(net117),
    .C(_0632_),
    .Y(_0029_));
 sg13g2_xnor2_1 _2872_ (.Y(_0633_),
    .A(net404),
    .B(_0632_));
 sg13g2_nor2_1 _2873_ (.A(net607),
    .B(_0633_),
    .Y(_0030_));
 sg13g2_a21oi_1 _2874_ (.A1(\pwm_module.prescaler0[8] ),
    .A2(_0632_),
    .Y(_0634_),
    .B1(net198));
 sg13g2_and3_1 _2875_ (.X(_0635_),
    .A(net198),
    .B(net558),
    .C(_0632_));
 sg13g2_nor3_1 _2876_ (.A(net608),
    .B(net199),
    .C(_0635_),
    .Y(_0031_));
 sg13g2_xnor2_1 _2877_ (.Y(_0636_),
    .A(net329),
    .B(_0635_));
 sg13g2_nor2_1 _2878_ (.A(net608),
    .B(net330),
    .Y(_0001_));
 sg13g2_a21oi_1 _2879_ (.A1(\pwm_module.prescaler0[10] ),
    .A2(_0635_),
    .Y(_0637_),
    .B1(net212));
 sg13g2_nand4_1 _2880_ (.B(\pwm_module.prescaler0[10] ),
    .C(\pwm_module.prescaler0[9] ),
    .A(\pwm_module.prescaler0[11] ),
    .Y(_0638_),
    .D(\pwm_module.prescaler0[8] ));
 sg13g2_nor4_2 _2881_ (.A(_0622_),
    .B(_0627_),
    .C(_0631_),
    .Y(_0639_),
    .D(_0638_));
 sg13g2_nor3_1 _2882_ (.A(net608),
    .B(net213),
    .C(_0639_),
    .Y(_0002_));
 sg13g2_xnor2_1 _2883_ (.Y(_0640_),
    .A(net333),
    .B(_0639_));
 sg13g2_nor2_1 _2884_ (.A(net608),
    .B(net334),
    .Y(_0003_));
 sg13g2_a21oi_1 _2885_ (.A1(\pwm_module.prescaler0[12] ),
    .A2(_0639_),
    .Y(_0641_),
    .B1(net132));
 sg13g2_and3_1 _2886_ (.X(_0642_),
    .A(net132),
    .B(net333),
    .C(_0639_));
 sg13g2_nor3_1 _2887_ (.A(net609),
    .B(net133),
    .C(_0642_),
    .Y(_0004_));
 sg13g2_xnor2_1 _2888_ (.Y(_0643_),
    .A(net348),
    .B(_0642_));
 sg13g2_nor2_1 _2889_ (.A(net609),
    .B(_0643_),
    .Y(_0005_));
 sg13g2_a21oi_1 _2890_ (.A1(\pwm_module.prescaler0[14] ),
    .A2(_0642_),
    .Y(_0644_),
    .B1(net154));
 sg13g2_and2_1 _2891_ (.A(\pwm_module.prescaler0[15] ),
    .B(\pwm_module.prescaler0[14] ),
    .X(_0645_));
 sg13g2_and4_2 _2892_ (.A(\pwm_module.prescaler0[13] ),
    .B(\pwm_module.prescaler0[12] ),
    .C(_0639_),
    .D(_0645_),
    .X(_0646_));
 sg13g2_nor3_1 _2893_ (.A(net609),
    .B(net155),
    .C(_0646_),
    .Y(_0006_));
 sg13g2_xnor2_1 _2894_ (.Y(_0647_),
    .A(net413),
    .B(_0646_));
 sg13g2_nor2_1 _2895_ (.A(net610),
    .B(_0647_),
    .Y(_0007_));
 sg13g2_a21oi_1 _2896_ (.A1(\pwm_module.prescaler0[16] ),
    .A2(_0646_),
    .Y(_0648_),
    .B1(net277));
 sg13g2_and3_1 _2897_ (.X(_0649_),
    .A(net277),
    .B(net553),
    .C(_0646_));
 sg13g2_nor3_1 _2898_ (.A(net610),
    .B(net278),
    .C(_0649_),
    .Y(_0008_));
 sg13g2_nand4_1 _2899_ (.B(net277),
    .C(net413),
    .A(net432),
    .Y(_0650_),
    .D(_0646_));
 sg13g2_o21ai_1 _2900_ (.B1(_0650_),
    .Y(_0651_),
    .A1(net432),
    .A2(_0649_));
 sg13g2_nor2_1 _2901_ (.A(net610),
    .B(net433),
    .Y(_0009_));
 sg13g2_a21oi_1 _2902_ (.A1(\pwm_module.prescaler0[18] ),
    .A2(_0649_),
    .Y(_0652_),
    .B1(net223));
 sg13g2_and4_1 _2903_ (.A(\pwm_module.prescaler0[19] ),
    .B(\pwm_module.prescaler0[18] ),
    .C(\pwm_module.prescaler0[17] ),
    .D(\pwm_module.prescaler0[16] ),
    .X(_0653_));
 sg13g2_and2_1 _2904_ (.A(_0646_),
    .B(_0653_),
    .X(_0654_));
 sg13g2_nor3_1 _2905_ (.A(net610),
    .B(net224),
    .C(_0654_),
    .Y(_0010_));
 sg13g2_nor2_1 _2906_ (.A(net390),
    .B(_0654_),
    .Y(_0655_));
 sg13g2_and2_1 _2907_ (.A(net390),
    .B(_0654_),
    .X(_0656_));
 sg13g2_nor3_1 _2908_ (.A(net610),
    .B(_0655_),
    .C(_0656_),
    .Y(_0012_));
 sg13g2_nor2_1 _2909_ (.A(net353),
    .B(_0656_),
    .Y(_0657_));
 sg13g2_and2_1 _2910_ (.A(net353),
    .B(_0656_),
    .X(_0658_));
 sg13g2_nor3_1 _2911_ (.A(net610),
    .B(net354),
    .C(_0658_),
    .Y(_0013_));
 sg13g2_nor2_1 _2912_ (.A(net303),
    .B(_0658_),
    .Y(_0659_));
 sg13g2_and2_1 _2913_ (.A(net303),
    .B(_0658_),
    .X(_0660_));
 sg13g2_nor3_1 _2914_ (.A(net610),
    .B(net304),
    .C(_0660_),
    .Y(_0014_));
 sg13g2_nor2_1 _2915_ (.A(net204),
    .B(_0660_),
    .Y(_0661_));
 sg13g2_and4_1 _2916_ (.A(\pwm_module.prescaler0[23] ),
    .B(\pwm_module.prescaler0[22] ),
    .C(\pwm_module.prescaler0[21] ),
    .D(\pwm_module.prescaler0[20] ),
    .X(_0662_));
 sg13g2_and2_1 _2917_ (.A(_0654_),
    .B(_0662_),
    .X(_0663_));
 sg13g2_nor3_1 _2918_ (.A(net610),
    .B(net205),
    .C(_0663_),
    .Y(_0015_));
 sg13g2_nor2_1 _2919_ (.A(net312),
    .B(_0663_),
    .Y(_0664_));
 sg13g2_and2_1 _2920_ (.A(net312),
    .B(_0663_),
    .X(_0665_));
 sg13g2_nor3_1 _2921_ (.A(net611),
    .B(_0664_),
    .C(_0665_),
    .Y(_0016_));
 sg13g2_nor2_1 _2922_ (.A(net381),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_and2_1 _2923_ (.A(net381),
    .B(_0665_),
    .X(_0667_));
 sg13g2_nor3_1 _2924_ (.A(net611),
    .B(_0666_),
    .C(_0667_),
    .Y(_0017_));
 sg13g2_nor2_1 _2925_ (.A(net265),
    .B(_0667_),
    .Y(_0668_));
 sg13g2_and3_1 _2926_ (.X(_0669_),
    .A(net265),
    .B(\pwm_module.prescaler0[25] ),
    .C(_0665_));
 sg13g2_nor3_1 _2927_ (.A(net611),
    .B(net266),
    .C(_0669_),
    .Y(_0018_));
 sg13g2_nor2_1 _2928_ (.A(net270),
    .B(_0669_),
    .Y(_0670_));
 sg13g2_and4_1 _2929_ (.A(\pwm_module.prescaler0[27] ),
    .B(\pwm_module.prescaler0[26] ),
    .C(\pwm_module.prescaler0[25] ),
    .D(\pwm_module.prescaler0[24] ),
    .X(_0671_));
 sg13g2_and2_1 _2930_ (.A(_0663_),
    .B(_0671_),
    .X(_0672_));
 sg13g2_nor3_1 _2931_ (.A(net611),
    .B(net271),
    .C(_0672_),
    .Y(_0019_));
 sg13g2_xnor2_1 _2932_ (.Y(_0673_),
    .A(net366),
    .B(_0672_));
 sg13g2_nor2_1 _2933_ (.A(net611),
    .B(_0673_),
    .Y(_0020_));
 sg13g2_a21oi_1 _2934_ (.A1(\pwm_module.prescaler0[28] ),
    .A2(_0672_),
    .Y(_0674_),
    .B1(net51));
 sg13g2_and3_1 _2935_ (.X(_0675_),
    .A(net51),
    .B(\pwm_module.prescaler0[28] ),
    .C(_0672_));
 sg13g2_nor3_1 _2936_ (.A(net611),
    .B(net52),
    .C(_0675_),
    .Y(_0021_));
 sg13g2_xnor2_1 _2937_ (.Y(_0676_),
    .A(net263),
    .B(_0675_));
 sg13g2_nor2_1 _2938_ (.A(net611),
    .B(net264),
    .Y(_0023_));
 sg13g2_a21oi_1 _2939_ (.A1(\pwm_module.prescaler0[30] ),
    .A2(_0675_),
    .Y(_0677_),
    .B1(net47));
 sg13g2_nor2_1 _2940_ (.A(_0617_),
    .B(net48),
    .Y(_0024_));
 sg13g2_nand2b_1 _2941_ (.Y(_0678_),
    .B(\pwm_module.prescaler1[1] ),
    .A_N(\MemCell.prescale_reg[0][1] ));
 sg13g2_nor2b_1 _2942_ (.A(\pwm_module.prescaler1[0] ),
    .B_N(\MemCell.prescale_reg[0][0] ),
    .Y(_0679_));
 sg13g2_nor2b_1 _2943_ (.A(\pwm_module.prescaler1[1] ),
    .B_N(\MemCell.prescale_reg[0][1] ),
    .Y(_0680_));
 sg13g2_a221oi_1 _2944_ (.B2(_0679_),
    .C1(_0680_),
    .B1(_0678_),
    .A1(_1848_),
    .Y(_0681_),
    .A2(\MemCell.prescale_reg[0][2] ));
 sg13g2_nand2_1 _2945_ (.Y(_0682_),
    .A(\pwm_module.prescaler1[3] ),
    .B(_1847_));
 sg13g2_nand2_1 _2946_ (.Y(_0683_),
    .A(\pwm_module.prescaler1[2] ),
    .B(_1849_));
 sg13g2_nand3b_1 _2947_ (.B(_0682_),
    .C(_0683_),
    .Y(_0684_),
    .A_N(_0681_));
 sg13g2_nand2b_1 _2948_ (.Y(_0685_),
    .B(\pwm_module.prescaler1[6] ),
    .A_N(\MemCell.prescale_reg[0][6] ));
 sg13g2_nand2b_1 _2949_ (.Y(_0686_),
    .B(\pwm_module.prescaler1[7] ),
    .A_N(\MemCell.prescale_reg[0][7] ));
 sg13g2_nand2_1 _2950_ (.Y(_0687_),
    .A(_0685_),
    .B(_0686_));
 sg13g2_nand2b_1 _2951_ (.Y(_0688_),
    .B(\MemCell.prescale_reg[0][7] ),
    .A_N(\pwm_module.prescaler1[7] ));
 sg13g2_nand2b_1 _2952_ (.Y(_0689_),
    .B(\MemCell.prescale_reg[0][6] ),
    .A_N(\pwm_module.prescaler1[6] ));
 sg13g2_nand4_1 _2953_ (.B(_0686_),
    .C(_0688_),
    .A(_0685_),
    .Y(_0690_),
    .D(_0689_));
 sg13g2_nor2b_1 _2954_ (.A(\MemCell.prescale_reg[0][5] ),
    .B_N(\pwm_module.prescaler1[5] ),
    .Y(_0691_));
 sg13g2_nor2b_1 _2955_ (.A(\MemCell.prescale_reg[0][4] ),
    .B_N(\pwm_module.prescaler1[4] ),
    .Y(_0692_));
 sg13g2_nand2b_1 _2956_ (.Y(_0693_),
    .B(\MemCell.prescale_reg[0][5] ),
    .A_N(\pwm_module.prescaler1[5] ));
 sg13g2_nand2b_1 _2957_ (.Y(_0694_),
    .B(\MemCell.prescale_reg[0][3] ),
    .A_N(\pwm_module.prescaler1[3] ));
 sg13g2_nand2b_1 _2958_ (.Y(_0695_),
    .B(_0694_),
    .A_N(_0691_));
 sg13g2_o21ai_1 _2959_ (.B1(_0693_),
    .Y(_0696_),
    .A1(\pwm_module.prescaler1[4] ),
    .A2(_1850_));
 sg13g2_nor4_1 _2960_ (.A(_0690_),
    .B(_0692_),
    .C(_0695_),
    .D(_0696_),
    .Y(_0697_));
 sg13g2_a21oi_1 _2961_ (.A1(_0692_),
    .A2(_0693_),
    .Y(_0698_),
    .B1(_0691_));
 sg13g2_nor2_1 _2962_ (.A(_0690_),
    .B(_0698_),
    .Y(_0699_));
 sg13g2_a221oi_1 _2963_ (.B2(_0684_),
    .C1(_0699_),
    .B1(_0697_),
    .A1(_0687_),
    .Y(_0700_),
    .A2(_0688_));
 sg13g2_nor2b_1 _2964_ (.A(\MemCell.prescale_reg[1][7] ),
    .B_N(\pwm_module.prescaler1[15] ),
    .Y(_0701_));
 sg13g2_nor2b_1 _2965_ (.A(\MemCell.prescale_reg[1][6] ),
    .B_N(\pwm_module.prescaler1[14] ),
    .Y(_0702_));
 sg13g2_nor2b_1 _2966_ (.A(\MemCell.prescale_reg[1][5] ),
    .B_N(\pwm_module.prescaler1[13] ),
    .Y(_0703_));
 sg13g2_nor2b_1 _2967_ (.A(\MemCell.prescale_reg[1][4] ),
    .B_N(\pwm_module.prescaler1[12] ),
    .Y(_0704_));
 sg13g2_nor4_1 _2968_ (.A(_0701_),
    .B(_0702_),
    .C(_0703_),
    .D(_0704_),
    .Y(_0705_));
 sg13g2_nor2b_1 _2969_ (.A(\pwm_module.prescaler1[15] ),
    .B_N(\MemCell.prescale_reg[1][7] ),
    .Y(_0706_));
 sg13g2_a21oi_1 _2970_ (.A1(_1853_),
    .A2(\MemCell.prescale_reg[1][4] ),
    .Y(_0707_),
    .B1(_0706_));
 sg13g2_a22oi_1 _2971_ (.Y(_0708_),
    .B1(_1852_),
    .B2(\MemCell.prescale_reg[1][5] ),
    .A2(\MemCell.prescale_reg[1][6] ),
    .A1(_1851_));
 sg13g2_and3_1 _2972_ (.X(_0709_),
    .A(_0705_),
    .B(_0707_),
    .C(_0708_));
 sg13g2_nor2b_1 _2973_ (.A(net652),
    .B_N(\pwm_module.prescaler1[11] ),
    .Y(_0710_));
 sg13g2_nor2b_1 _2974_ (.A(\MemCell.prescale_reg[1][2] ),
    .B_N(\pwm_module.prescaler1[10] ),
    .Y(_0711_));
 sg13g2_nor2b_1 _2975_ (.A(\pwm_module.prescaler1[10] ),
    .B_N(\MemCell.prescale_reg[1][2] ),
    .Y(_0712_));
 sg13g2_nor2b_1 _2976_ (.A(\pwm_module.prescaler1[11] ),
    .B_N(net652),
    .Y(_0713_));
 sg13g2_nand2b_1 _2977_ (.Y(_0714_),
    .B(net652),
    .A_N(\pwm_module.prescaler1[11] ));
 sg13g2_or4_1 _2978_ (.A(_0710_),
    .B(_0711_),
    .C(_0712_),
    .D(_0713_),
    .X(_0715_));
 sg13g2_nor2b_1 _2979_ (.A(\MemCell.prescale_reg[1][1] ),
    .B_N(\pwm_module.prescaler1[9] ),
    .Y(_0716_));
 sg13g2_nor2b_1 _2980_ (.A(\MemCell.prescale_reg[1][0] ),
    .B_N(\pwm_module.prescaler1[8] ),
    .Y(_0717_));
 sg13g2_nor2_1 _2981_ (.A(_0716_),
    .B(_0717_),
    .Y(_0718_));
 sg13g2_nand2b_1 _2982_ (.Y(_0719_),
    .B(\MemCell.prescale_reg[1][1] ),
    .A_N(\pwm_module.prescaler1[9] ));
 sg13g2_o21ai_1 _2983_ (.B1(_0719_),
    .Y(_0720_),
    .A1(\pwm_module.prescaler1[8] ),
    .A2(_1854_));
 sg13g2_nor2_1 _2984_ (.A(_0715_),
    .B(_0720_),
    .Y(_0721_));
 sg13g2_nand3_1 _2985_ (.B(_0718_),
    .C(_0721_),
    .A(_0709_),
    .Y(_0722_));
 sg13g2_o21ai_1 _2986_ (.B1(_0714_),
    .Y(_0723_),
    .A1(_0710_),
    .A2(_0711_));
 sg13g2_a21oi_1 _2987_ (.A1(_0717_),
    .A2(_0719_),
    .Y(_0724_),
    .B1(_0716_));
 sg13g2_o21ai_1 _2988_ (.B1(_0723_),
    .Y(_0725_),
    .A1(_0715_),
    .A2(_0724_));
 sg13g2_or3_1 _2989_ (.A(_0701_),
    .B(_0702_),
    .C(_0708_),
    .X(_0726_));
 sg13g2_nor2_1 _2990_ (.A(_0705_),
    .B(_0706_),
    .Y(_0727_));
 sg13g2_a22oi_1 _2991_ (.Y(_0728_),
    .B1(_0726_),
    .B2(_0727_),
    .A2(_0725_),
    .A1(_0709_));
 sg13g2_o21ai_1 _2992_ (.B1(_0728_),
    .Y(_0729_),
    .A1(_0700_),
    .A2(_0722_));
 sg13g2_nor2b_1 _2993_ (.A(\MemCell.prescale_reg[3][7] ),
    .B_N(\pwm_module.prescaler1[31] ),
    .Y(_0730_));
 sg13g2_a21o_1 _2994_ (.A2(_1855_),
    .A1(\pwm_module.prescaler1[30] ),
    .B1(_0730_),
    .X(_0731_));
 sg13g2_nand2b_1 _2995_ (.Y(_0732_),
    .B(\MemCell.prescale_reg[3][5] ),
    .A_N(\pwm_module.prescaler1[29] ));
 sg13g2_nand2b_1 _2996_ (.Y(_0733_),
    .B(\MemCell.prescale_reg[3][7] ),
    .A_N(\pwm_module.prescaler1[31] ));
 sg13g2_nand2b_1 _2997_ (.Y(_0734_),
    .B(\MemCell.prescale_reg[3][6] ),
    .A_N(\pwm_module.prescaler1[30] ));
 sg13g2_nand3_1 _2998_ (.B(_0733_),
    .C(_0734_),
    .A(_0732_),
    .Y(_0735_));
 sg13g2_nor2_1 _2999_ (.A(_0731_),
    .B(_0735_),
    .Y(_0736_));
 sg13g2_nor2_1 _3000_ (.A(\pwm_module.prescaler1[28] ),
    .B(_1856_),
    .Y(_0737_));
 sg13g2_nor2b_1 _3001_ (.A(\MemCell.prescale_reg[3][5] ),
    .B_N(\pwm_module.prescaler1[29] ),
    .Y(_0738_));
 sg13g2_a21o_1 _3002_ (.A2(_1856_),
    .A1(\pwm_module.prescaler1[28] ),
    .B1(_0738_),
    .X(_0739_));
 sg13g2_or4_1 _3003_ (.A(_0731_),
    .B(_0735_),
    .C(_0737_),
    .D(_0739_),
    .X(_0740_));
 sg13g2_nor2b_1 _3004_ (.A(\MemCell.prescale_reg[3][2] ),
    .B_N(\pwm_module.prescaler1[26] ),
    .Y(_0741_));
 sg13g2_nor2b_1 _3005_ (.A(\MemCell.prescale_reg[3][3] ),
    .B_N(\pwm_module.prescaler1[27] ),
    .Y(_0742_));
 sg13g2_nor2b_1 _3006_ (.A(\pwm_module.prescaler1[27] ),
    .B_N(\MemCell.prescale_reg[3][3] ),
    .Y(_0743_));
 sg13g2_nand2b_1 _3007_ (.Y(_0744_),
    .B(\MemCell.prescale_reg[3][3] ),
    .A_N(\pwm_module.prescaler1[27] ));
 sg13g2_nor2b_1 _3008_ (.A(\pwm_module.prescaler1[26] ),
    .B_N(\MemCell.prescale_reg[3][2] ),
    .Y(_0745_));
 sg13g2_nor4_1 _3009_ (.A(_0741_),
    .B(_0742_),
    .C(_0743_),
    .D(_0745_),
    .Y(_0746_));
 sg13g2_nand2b_1 _3010_ (.Y(_0747_),
    .B(\pwm_module.prescaler1[24] ),
    .A_N(\MemCell.prescale_reg[3][0] ));
 sg13g2_nand2b_1 _3011_ (.Y(_0748_),
    .B(\pwm_module.prescaler1[25] ),
    .A_N(\MemCell.prescale_reg[3][1] ));
 sg13g2_nor2b_1 _3012_ (.A(\pwm_module.prescaler1[25] ),
    .B_N(\MemCell.prescale_reg[3][1] ),
    .Y(_0749_));
 sg13g2_xor2_1 _3013_ (.B(\MemCell.prescale_reg[3][0] ),
    .A(\pwm_module.prescaler1[24] ),
    .X(_0750_));
 sg13g2_nand3b_1 _3014_ (.B(_0746_),
    .C(_0748_),
    .Y(_0751_),
    .A_N(_0749_));
 sg13g2_nor3_1 _3015_ (.A(_0740_),
    .B(_0750_),
    .C(_0751_),
    .Y(_0752_));
 sg13g2_nor2b_1 _3016_ (.A(\MemCell.prescale_reg[2][6] ),
    .B_N(\pwm_module.prescaler1[22] ),
    .Y(_0753_));
 sg13g2_nor2b_1 _3017_ (.A(\MemCell.prescale_reg[2][7] ),
    .B_N(\pwm_module.prescaler1[23] ),
    .Y(_0754_));
 sg13g2_nor2b_1 _3018_ (.A(\pwm_module.prescaler1[23] ),
    .B_N(\MemCell.prescale_reg[2][7] ),
    .Y(_0755_));
 sg13g2_nand2b_1 _3019_ (.Y(_0756_),
    .B(\MemCell.prescale_reg[2][7] ),
    .A_N(\pwm_module.prescaler1[23] ));
 sg13g2_nor2b_1 _3020_ (.A(\pwm_module.prescaler1[22] ),
    .B_N(\MemCell.prescale_reg[2][6] ),
    .Y(_0757_));
 sg13g2_nand2b_1 _3021_ (.Y(_0758_),
    .B(\MemCell.prescale_reg[2][5] ),
    .A_N(\pwm_module.prescaler1[21] ));
 sg13g2_nor4_1 _3022_ (.A(_0753_),
    .B(_0754_),
    .C(_0755_),
    .D(_0757_),
    .Y(_0759_));
 sg13g2_nand2b_1 _3023_ (.Y(_0760_),
    .B(\pwm_module.prescaler1[21] ),
    .A_N(\MemCell.prescale_reg[2][5] ));
 sg13g2_o21ai_1 _3024_ (.B1(_0760_),
    .Y(_0761_),
    .A1(_1861_),
    .A2(\MemCell.prescale_reg[2][4] ));
 sg13g2_xnor2_1 _3025_ (.Y(_0762_),
    .A(\pwm_module.prescaler1[20] ),
    .B(\MemCell.prescale_reg[2][4] ));
 sg13g2_nand4_1 _3026_ (.B(_0759_),
    .C(_0760_),
    .A(_0758_),
    .Y(_0763_),
    .D(_0762_));
 sg13g2_nand2b_1 _3027_ (.Y(_0764_),
    .B(\pwm_module.prescaler1[18] ),
    .A_N(\MemCell.prescale_reg[2][2] ));
 sg13g2_nand2b_1 _3028_ (.Y(_0765_),
    .B(\pwm_module.prescaler1[19] ),
    .A_N(net653));
 sg13g2_nand2_1 _3029_ (.Y(_0766_),
    .A(_0764_),
    .B(_0765_));
 sg13g2_nand2b_1 _3030_ (.Y(_0767_),
    .B(\MemCell.prescale_reg[2][2] ),
    .A_N(\pwm_module.prescaler1[18] ));
 sg13g2_nand2b_1 _3031_ (.Y(_0768_),
    .B(net653),
    .A_N(\pwm_module.prescaler1[19] ));
 sg13g2_and4_1 _3032_ (.A(_0764_),
    .B(_0765_),
    .C(_0767_),
    .D(_0768_),
    .X(_0769_));
 sg13g2_inv_1 _3033_ (.Y(_0770_),
    .A(_0769_));
 sg13g2_nor2b_1 _3034_ (.A(\MemCell.prescale_reg[2][0] ),
    .B_N(\pwm_module.prescaler1[16] ),
    .Y(_0771_));
 sg13g2_nand2b_1 _3035_ (.Y(_0772_),
    .B(\pwm_module.prescaler1[16] ),
    .A_N(\MemCell.prescale_reg[2][0] ));
 sg13g2_nor2b_1 _3036_ (.A(\pwm_module.prescaler1[16] ),
    .B_N(\MemCell.prescale_reg[2][0] ),
    .Y(_0773_));
 sg13g2_nand2b_1 _3037_ (.Y(_0774_),
    .B(\MemCell.prescale_reg[2][1] ),
    .A_N(\pwm_module.prescaler1[17] ));
 sg13g2_nor2b_1 _3038_ (.A(\MemCell.prescale_reg[2][1] ),
    .B_N(\pwm_module.prescaler1[17] ),
    .Y(_0775_));
 sg13g2_nor4_1 _3039_ (.A(_0763_),
    .B(_0770_),
    .C(_0773_),
    .D(_0775_),
    .Y(_0776_));
 sg13g2_and4_1 _3040_ (.A(_0752_),
    .B(_0772_),
    .C(_0774_),
    .D(_0776_),
    .X(_0777_));
 sg13g2_a21o_1 _3041_ (.A2(_0774_),
    .A1(_0771_),
    .B1(_0775_),
    .X(_0778_));
 sg13g2_a22oi_1 _3042_ (.Y(_0779_),
    .B1(_0769_),
    .B2(_0778_),
    .A2(_0768_),
    .A1(_0766_));
 sg13g2_o21ai_1 _3043_ (.B1(_0756_),
    .Y(_0780_),
    .A1(_0753_),
    .A2(_0754_));
 sg13g2_nand3_1 _3044_ (.B(_0759_),
    .C(_0761_),
    .A(_0758_),
    .Y(_0781_));
 sg13g2_o21ai_1 _3045_ (.B1(_0781_),
    .Y(_0782_),
    .A1(_0763_),
    .A2(_0779_));
 sg13g2_nand2b_1 _3046_ (.Y(_0783_),
    .B(_0780_),
    .A_N(_0782_));
 sg13g2_a22oi_1 _3047_ (.Y(_0784_),
    .B1(_0736_),
    .B2(_0739_),
    .A2(_0733_),
    .A1(_0731_));
 sg13g2_o21ai_1 _3048_ (.B1(_0744_),
    .Y(_0785_),
    .A1(_0741_),
    .A2(_0742_));
 sg13g2_o21ai_1 _3049_ (.B1(_0748_),
    .Y(_0786_),
    .A1(_0747_),
    .A2(_0749_));
 sg13g2_nand2_1 _3050_ (.Y(_0787_),
    .A(_0746_),
    .B(_0786_));
 sg13g2_and2_1 _3051_ (.A(_0785_),
    .B(_0787_),
    .X(_0788_));
 sg13g2_o21ai_1 _3052_ (.B1(_0784_),
    .Y(_0789_),
    .A1(_0740_),
    .A2(_0788_));
 sg13g2_a221oi_1 _3053_ (.B2(_0752_),
    .C1(_0789_),
    .B1(_0783_),
    .A1(_0729_),
    .Y(_0790_),
    .A2(_0777_));
 sg13g2_nand2_1 _3054_ (.Y(_0791_),
    .A(net651),
    .B(_0790_));
 sg13g2_nor2_1 _3055_ (.A(net119),
    .B(net601),
    .Y(_0032_));
 sg13g2_xnor2_1 _3056_ (.Y(_0792_),
    .A(net119),
    .B(net309));
 sg13g2_nor2_1 _3057_ (.A(net601),
    .B(_0792_),
    .Y(_0043_));
 sg13g2_and3_1 _3058_ (.X(_0793_),
    .A(net119),
    .B(\pwm_module.prescaler1[1] ),
    .C(net122));
 sg13g2_a21oi_1 _3059_ (.A1(net119),
    .A2(\pwm_module.prescaler1[1] ),
    .Y(_0794_),
    .B1(net122));
 sg13g2_nor3_1 _3060_ (.A(net601),
    .B(_0793_),
    .C(net123),
    .Y(_0054_));
 sg13g2_and4_2 _3061_ (.A(\pwm_module.prescaler1[0] ),
    .B(\pwm_module.prescaler1[1] ),
    .C(net190),
    .D(net122),
    .X(_0795_));
 sg13g2_nor2_1 _3062_ (.A(net190),
    .B(_0793_),
    .Y(_0796_));
 sg13g2_nor3_1 _3063_ (.A(net601),
    .B(_0795_),
    .C(net191),
    .Y(_0057_));
 sg13g2_nor2_1 _3064_ (.A(net320),
    .B(_0795_),
    .Y(_0797_));
 sg13g2_and2_1 _3065_ (.A(net320),
    .B(_0795_),
    .X(_0798_));
 sg13g2_nor3_1 _3066_ (.A(net601),
    .B(net321),
    .C(_0798_),
    .Y(_0058_));
 sg13g2_nor2_1 _3067_ (.A(net243),
    .B(_0798_),
    .Y(_0799_));
 sg13g2_and2_1 _3068_ (.A(\pwm_module.prescaler1[5] ),
    .B(\pwm_module.prescaler1[4] ),
    .X(_0800_));
 sg13g2_and2_1 _3069_ (.A(_0795_),
    .B(_0800_),
    .X(_0801_));
 sg13g2_nor3_1 _3070_ (.A(net601),
    .B(net244),
    .C(_0801_),
    .Y(_0059_));
 sg13g2_xnor2_1 _3071_ (.Y(_0802_),
    .A(net331),
    .B(_0801_));
 sg13g2_nor2_1 _3072_ (.A(net601),
    .B(_0802_),
    .Y(_0060_));
 sg13g2_a21oi_1 _3073_ (.A1(\pwm_module.prescaler1[6] ),
    .A2(_0801_),
    .Y(_0803_),
    .B1(net171));
 sg13g2_and4_2 _3074_ (.A(net171),
    .B(\pwm_module.prescaler1[6] ),
    .C(_0795_),
    .D(_0800_),
    .X(_0804_));
 sg13g2_nor3_1 _3075_ (.A(net601),
    .B(net172),
    .C(_0804_),
    .Y(_0061_));
 sg13g2_xnor2_1 _3076_ (.Y(_0805_),
    .A(net323),
    .B(_0804_));
 sg13g2_nor2_1 _3077_ (.A(net602),
    .B(net324),
    .Y(_0062_));
 sg13g2_a21oi_1 _3078_ (.A1(\pwm_module.prescaler1[8] ),
    .A2(_0804_),
    .Y(_0806_),
    .B1(net135));
 sg13g2_and2_1 _3079_ (.A(\pwm_module.prescaler1[9] ),
    .B(\pwm_module.prescaler1[8] ),
    .X(_0807_));
 sg13g2_and2_1 _3080_ (.A(_0804_),
    .B(_0807_),
    .X(_0808_));
 sg13g2_nor3_1 _3081_ (.A(net602),
    .B(net136),
    .C(_0808_),
    .Y(_0063_));
 sg13g2_xnor2_1 _3082_ (.Y(_0809_),
    .A(net332),
    .B(_0808_));
 sg13g2_nor2_1 _3083_ (.A(net602),
    .B(_0809_),
    .Y(_0033_));
 sg13g2_a21oi_1 _3084_ (.A1(\pwm_module.prescaler1[10] ),
    .A2(_0808_),
    .Y(_0810_),
    .B1(net147));
 sg13g2_and4_2 _3085_ (.A(net147),
    .B(net556),
    .C(_0804_),
    .D(_0807_),
    .X(_0811_));
 sg13g2_nor3_1 _3086_ (.A(net602),
    .B(net148),
    .C(_0811_),
    .Y(_0034_));
 sg13g2_nor2_1 _3087_ (.A(net186),
    .B(_0811_),
    .Y(_0812_));
 sg13g2_and2_1 _3088_ (.A(net186),
    .B(_0811_),
    .X(_0813_));
 sg13g2_nor3_1 _3089_ (.A(net602),
    .B(_0812_),
    .C(_0813_),
    .Y(_0035_));
 sg13g2_nor2_1 _3090_ (.A(net206),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_nor2_1 _3091_ (.A(_1852_),
    .B(_1853_),
    .Y(_0815_));
 sg13g2_and2_1 _3092_ (.A(_0811_),
    .B(_0815_),
    .X(_0816_));
 sg13g2_nor3_1 _3093_ (.A(net605),
    .B(_0814_),
    .C(_0816_),
    .Y(_0036_));
 sg13g2_xnor2_1 _3094_ (.Y(_0817_),
    .A(net344),
    .B(_0816_));
 sg13g2_nor2_1 _3095_ (.A(net605),
    .B(_0817_),
    .Y(_0037_));
 sg13g2_a21oi_1 _3096_ (.A1(\pwm_module.prescaler1[14] ),
    .A2(_0816_),
    .Y(_0818_),
    .B1(net88));
 sg13g2_and2_1 _3097_ (.A(\pwm_module.prescaler1[15] ),
    .B(\pwm_module.prescaler1[14] ),
    .X(_0819_));
 sg13g2_and3_1 _3098_ (.X(_0820_),
    .A(_0811_),
    .B(_0815_),
    .C(_0819_));
 sg13g2_nand3_1 _3099_ (.B(_0815_),
    .C(_0819_),
    .A(_0811_),
    .Y(_0821_));
 sg13g2_nor3_1 _3100_ (.A(net605),
    .B(net89),
    .C(_0820_),
    .Y(_0038_));
 sg13g2_nor2_1 _3101_ (.A(net419),
    .B(_0820_),
    .Y(_0822_));
 sg13g2_and2_1 _3102_ (.A(net419),
    .B(_0820_),
    .X(_0823_));
 sg13g2_nor3_1 _3103_ (.A(net605),
    .B(_0822_),
    .C(_0823_),
    .Y(_0039_));
 sg13g2_nor2_1 _3104_ (.A(net284),
    .B(_0823_),
    .Y(_0824_));
 sg13g2_and2_1 _3105_ (.A(net284),
    .B(_0823_),
    .X(_0825_));
 sg13g2_nor3_1 _3106_ (.A(net605),
    .B(net285),
    .C(_0825_),
    .Y(_0040_));
 sg13g2_nor2_1 _3107_ (.A(net420),
    .B(_0825_),
    .Y(_0826_));
 sg13g2_and2_1 _3108_ (.A(net420),
    .B(_0825_),
    .X(_0827_));
 sg13g2_nor3_1 _3109_ (.A(net605),
    .B(_0826_),
    .C(_0827_),
    .Y(_0041_));
 sg13g2_nor2_1 _3110_ (.A(net292),
    .B(_0827_),
    .Y(_0828_));
 sg13g2_nand4_1 _3111_ (.B(\pwm_module.prescaler1[18] ),
    .C(\pwm_module.prescaler1[17] ),
    .A(\pwm_module.prescaler1[19] ),
    .Y(_0829_),
    .D(\pwm_module.prescaler1[16] ));
 sg13g2_nor2_1 _3112_ (.A(_0821_),
    .B(_0829_),
    .Y(_0830_));
 sg13g2_nor3_1 _3113_ (.A(net605),
    .B(net293),
    .C(_0830_),
    .Y(_0042_));
 sg13g2_nor2_1 _3114_ (.A(net280),
    .B(_0830_),
    .Y(_0831_));
 sg13g2_nor3_2 _3115_ (.A(_1861_),
    .B(_0821_),
    .C(_0829_),
    .Y(_0832_));
 sg13g2_nor3_1 _3116_ (.A(net604),
    .B(_0831_),
    .C(_0832_),
    .Y(_0044_));
 sg13g2_nor2_1 _3117_ (.A(net363),
    .B(_0832_),
    .Y(_0833_));
 sg13g2_and2_1 _3118_ (.A(net363),
    .B(_0832_),
    .X(_0834_));
 sg13g2_nor3_1 _3119_ (.A(net604),
    .B(_0833_),
    .C(_0834_),
    .Y(_0045_));
 sg13g2_nor2_1 _3120_ (.A(net411),
    .B(_0834_),
    .Y(_0835_));
 sg13g2_and3_1 _3121_ (.X(_0836_),
    .A(net411),
    .B(net363),
    .C(_0832_));
 sg13g2_nor3_1 _3122_ (.A(net604),
    .B(_0835_),
    .C(_0836_),
    .Y(_0046_));
 sg13g2_nor2_1 _3123_ (.A(net400),
    .B(_0836_),
    .Y(_0837_));
 sg13g2_nand4_1 _3124_ (.B(\pwm_module.prescaler1[22] ),
    .C(\pwm_module.prescaler1[21] ),
    .A(net400),
    .Y(_0838_),
    .D(\pwm_module.prescaler1[20] ));
 sg13g2_nor3_2 _3125_ (.A(_0821_),
    .B(_0829_),
    .C(_0838_),
    .Y(_0839_));
 sg13g2_nor3_1 _3126_ (.A(net603),
    .B(net401),
    .C(_0839_),
    .Y(_0047_));
 sg13g2_nor2_1 _3127_ (.A(net445),
    .B(_0839_),
    .Y(_0840_));
 sg13g2_and2_1 _3128_ (.A(net445),
    .B(_0839_),
    .X(_0841_));
 sg13g2_nor3_1 _3129_ (.A(net604),
    .B(net446),
    .C(_0841_),
    .Y(_0048_));
 sg13g2_nor2_1 _3130_ (.A(net313),
    .B(_0841_),
    .Y(_0842_));
 sg13g2_and3_1 _3131_ (.X(_0843_),
    .A(net313),
    .B(net555),
    .C(_0839_));
 sg13g2_nor3_1 _3132_ (.A(net603),
    .B(net314),
    .C(_0843_),
    .Y(_0049_));
 sg13g2_nor2_1 _3133_ (.A(net379),
    .B(_0843_),
    .Y(_0844_));
 sg13g2_and2_1 _3134_ (.A(net379),
    .B(_0843_),
    .X(_0845_));
 sg13g2_nor3_1 _3135_ (.A(net603),
    .B(_0844_),
    .C(_0845_),
    .Y(_0050_));
 sg13g2_nor2_1 _3136_ (.A(net336),
    .B(_0845_),
    .Y(_0846_));
 sg13g2_nand4_1 _3137_ (.B(\pwm_module.prescaler1[26] ),
    .C(net313),
    .A(net336),
    .Y(_0847_),
    .D(\pwm_module.prescaler1[24] ));
 sg13g2_nor4_2 _3138_ (.A(_0821_),
    .B(_0829_),
    .C(_0838_),
    .Y(_0848_),
    .D(_0847_));
 sg13g2_nor3_1 _3139_ (.A(net603),
    .B(net337),
    .C(_0848_),
    .Y(_0051_));
 sg13g2_nor2_1 _3140_ (.A(net375),
    .B(_0848_),
    .Y(_0849_));
 sg13g2_and2_1 _3141_ (.A(net375),
    .B(_0848_),
    .X(_0850_));
 sg13g2_nor3_1 _3142_ (.A(net603),
    .B(net376),
    .C(_0850_),
    .Y(_0052_));
 sg13g2_nor2_1 _3143_ (.A(net174),
    .B(_0850_),
    .Y(_0851_));
 sg13g2_and3_1 _3144_ (.X(_0852_),
    .A(net174),
    .B(\pwm_module.prescaler1[28] ),
    .C(_0848_));
 sg13g2_nor3_1 _3145_ (.A(net603),
    .B(net175),
    .C(_0852_),
    .Y(_0053_));
 sg13g2_nor2_1 _3146_ (.A(net235),
    .B(_0852_),
    .Y(_0853_));
 sg13g2_a21oi_1 _3147_ (.A1(net235),
    .A2(_0852_),
    .Y(_0854_),
    .B1(net603));
 sg13g2_nor2b_1 _3148_ (.A(net236),
    .B_N(_0854_),
    .Y(_0055_));
 sg13g2_a21oi_1 _3149_ (.A1(\pwm_module.prescaler1[30] ),
    .A2(_0852_),
    .Y(_0855_),
    .B1(net41));
 sg13g2_nor2_1 _3150_ (.A(net603),
    .B(net42),
    .Y(_0056_));
 sg13g2_nand2b_1 _3151_ (.Y(_0856_),
    .B(\pwm_module.prescaler2[1] ),
    .A_N(\MemCell.prescale_reg[0][1] ));
 sg13g2_nor2b_1 _3152_ (.A(\pwm_module.prescaler2[0] ),
    .B_N(\MemCell.prescale_reg[0][0] ),
    .Y(_0857_));
 sg13g2_nor2b_1 _3153_ (.A(\pwm_module.prescaler2[1] ),
    .B_N(\MemCell.prescale_reg[0][1] ),
    .Y(_0858_));
 sg13g2_a221oi_1 _3154_ (.B2(_0857_),
    .C1(_0858_),
    .B1(_0856_),
    .A1(\MemCell.prescale_reg[0][2] ),
    .Y(_0859_),
    .A2(_1866_));
 sg13g2_a221oi_1 _3155_ (.B2(_1849_),
    .C1(_0859_),
    .B1(\pwm_module.prescaler2[2] ),
    .A1(_1847_),
    .Y(_0860_),
    .A2(\pwm_module.prescaler2[3] ));
 sg13g2_nand2b_1 _3156_ (.Y(_0861_),
    .B(\pwm_module.prescaler2[7] ),
    .A_N(\MemCell.prescale_reg[0][7] ));
 sg13g2_nand2b_1 _3157_ (.Y(_0862_),
    .B(\pwm_module.prescaler2[6] ),
    .A_N(\MemCell.prescale_reg[0][6] ));
 sg13g2_nand2_1 _3158_ (.Y(_0863_),
    .A(_0861_),
    .B(_0862_));
 sg13g2_nand2b_1 _3159_ (.Y(_0864_),
    .B(\MemCell.prescale_reg[0][6] ),
    .A_N(\pwm_module.prescaler2[6] ));
 sg13g2_nand2b_1 _3160_ (.Y(_0865_),
    .B(\MemCell.prescale_reg[0][7] ),
    .A_N(\pwm_module.prescaler2[7] ));
 sg13g2_and4_1 _3161_ (.A(_0861_),
    .B(_0862_),
    .C(_0864_),
    .D(_0865_),
    .X(_0866_));
 sg13g2_nand2b_1 _3162_ (.Y(_0867_),
    .B(\pwm_module.prescaler2[4] ),
    .A_N(\MemCell.prescale_reg[0][4] ));
 sg13g2_nand2b_1 _3163_ (.Y(_0868_),
    .B(\pwm_module.prescaler2[5] ),
    .A_N(\MemCell.prescale_reg[0][5] ));
 sg13g2_nor2b_1 _3164_ (.A(\pwm_module.prescaler2[5] ),
    .B_N(\MemCell.prescale_reg[0][5] ),
    .Y(_0869_));
 sg13g2_a221oi_1 _3165_ (.B2(\MemCell.prescale_reg[0][3] ),
    .C1(_0869_),
    .B1(_1865_),
    .A1(\MemCell.prescale_reg[0][4] ),
    .Y(_0870_),
    .A2(_1864_));
 sg13g2_nand4_1 _3166_ (.B(_0867_),
    .C(_0868_),
    .A(_0866_),
    .Y(_0871_),
    .D(_0870_));
 sg13g2_a21oi_1 _3167_ (.A1(_0867_),
    .A2(_0868_),
    .Y(_0872_),
    .B1(_0869_));
 sg13g2_a22oi_1 _3168_ (.Y(_0873_),
    .B1(_0866_),
    .B2(_0872_),
    .A2(_0865_),
    .A1(_0863_));
 sg13g2_o21ai_1 _3169_ (.B1(_0873_),
    .Y(_0874_),
    .A1(_0860_),
    .A2(_0871_));
 sg13g2_nand2b_1 _3170_ (.Y(_0875_),
    .B(\pwm_module.prescaler2[15] ),
    .A_N(\MemCell.prescale_reg[1][7] ));
 sg13g2_nand2b_1 _3171_ (.Y(_0876_),
    .B(\pwm_module.prescaler2[14] ),
    .A_N(\MemCell.prescale_reg[1][6] ));
 sg13g2_nand2_1 _3172_ (.Y(_0877_),
    .A(_0875_),
    .B(_0876_));
 sg13g2_nand2b_1 _3173_ (.Y(_0878_),
    .B(\MemCell.prescale_reg[1][7] ),
    .A_N(\pwm_module.prescaler2[15] ));
 sg13g2_nand2b_1 _3174_ (.Y(_0879_),
    .B(\MemCell.prescale_reg[1][6] ),
    .A_N(\pwm_module.prescaler2[14] ));
 sg13g2_nor2b_1 _3175_ (.A(\pwm_module.prescaler2[13] ),
    .B_N(\MemCell.prescale_reg[1][5] ),
    .Y(_0880_));
 sg13g2_nand2b_1 _3176_ (.Y(_0881_),
    .B(\MemCell.prescale_reg[1][5] ),
    .A_N(\pwm_module.prescaler2[13] ));
 sg13g2_and4_1 _3177_ (.A(_0875_),
    .B(_0876_),
    .C(_0878_),
    .D(_0879_),
    .X(_0882_));
 sg13g2_nand2b_1 _3178_ (.Y(_0883_),
    .B(\pwm_module.prescaler2[12] ),
    .A_N(\MemCell.prescale_reg[1][4] ));
 sg13g2_nand2b_1 _3179_ (.Y(_0884_),
    .B(\pwm_module.prescaler2[13] ),
    .A_N(\MemCell.prescale_reg[1][5] ));
 sg13g2_nand2b_1 _3180_ (.Y(_0885_),
    .B(\MemCell.prescale_reg[1][4] ),
    .A_N(\pwm_module.prescaler2[12] ));
 sg13g2_nand3_1 _3181_ (.B(_0884_),
    .C(_0885_),
    .A(_0883_),
    .Y(_0886_));
 sg13g2_nand3b_1 _3182_ (.B(_0881_),
    .C(_0882_),
    .Y(_0887_),
    .A_N(_0886_));
 sg13g2_nand2b_1 _3183_ (.Y(_0888_),
    .B(\pwm_module.prescaler2[11] ),
    .A_N(net652));
 sg13g2_nand2b_1 _3184_ (.Y(_0889_),
    .B(\pwm_module.prescaler2[10] ),
    .A_N(\MemCell.prescale_reg[1][2] ));
 sg13g2_nand2_1 _3185_ (.Y(_0890_),
    .A(_0888_),
    .B(_0889_));
 sg13g2_nand2b_1 _3186_ (.Y(_0891_),
    .B(\MemCell.prescale_reg[1][2] ),
    .A_N(\pwm_module.prescaler2[10] ));
 sg13g2_nand2b_1 _3187_ (.Y(_0892_),
    .B(net652),
    .A_N(\pwm_module.prescaler2[11] ));
 sg13g2_and4_1 _3188_ (.A(_0888_),
    .B(_0889_),
    .C(_0891_),
    .D(_0892_),
    .X(_0893_));
 sg13g2_nand2b_1 _3189_ (.Y(_0894_),
    .B(\pwm_module.prescaler2[8] ),
    .A_N(\MemCell.prescale_reg[1][0] ));
 sg13g2_nand2b_1 _3190_ (.Y(_0895_),
    .B(\pwm_module.prescaler2[9] ),
    .A_N(\MemCell.prescale_reg[1][1] ));
 sg13g2_nand2_1 _3191_ (.Y(_0896_),
    .A(_0894_),
    .B(_0895_));
 sg13g2_nor2b_1 _3192_ (.A(\pwm_module.prescaler2[9] ),
    .B_N(\MemCell.prescale_reg[1][1] ),
    .Y(_0897_));
 sg13g2_o21ai_1 _3193_ (.B1(_0893_),
    .Y(_0898_),
    .A1(_1854_),
    .A2(\pwm_module.prescaler2[8] ));
 sg13g2_nor4_1 _3194_ (.A(_0887_),
    .B(_0896_),
    .C(_0897_),
    .D(_0898_),
    .Y(_0899_));
 sg13g2_a21oi_1 _3195_ (.A1(_0894_),
    .A2(_0895_),
    .Y(_0900_),
    .B1(_0897_));
 sg13g2_a22oi_1 _3196_ (.Y(_0901_),
    .B1(_0893_),
    .B2(_0900_),
    .A2(_0892_),
    .A1(_0890_));
 sg13g2_a21oi_1 _3197_ (.A1(_0883_),
    .A2(_0884_),
    .Y(_0902_),
    .B1(_0880_));
 sg13g2_a22oi_1 _3198_ (.Y(_0903_),
    .B1(_0882_),
    .B2(_0902_),
    .A2(_0878_),
    .A1(_0877_));
 sg13g2_o21ai_1 _3199_ (.B1(_0903_),
    .Y(_0904_),
    .A1(_0887_),
    .A2(_0901_));
 sg13g2_a21o_2 _3200_ (.A2(_0899_),
    .A1(_0874_),
    .B1(_0904_),
    .X(_0905_));
 sg13g2_nand2b_1 _3201_ (.Y(_0906_),
    .B(\pwm_module.prescaler2[23] ),
    .A_N(\MemCell.prescale_reg[2][7] ));
 sg13g2_nand2b_1 _3202_ (.Y(_0907_),
    .B(\pwm_module.prescaler2[22] ),
    .A_N(\MemCell.prescale_reg[2][6] ));
 sg13g2_nand2_1 _3203_ (.Y(_0908_),
    .A(_0906_),
    .B(_0907_));
 sg13g2_nand2b_1 _3204_ (.Y(_0909_),
    .B(\MemCell.prescale_reg[2][7] ),
    .A_N(\pwm_module.prescaler2[23] ));
 sg13g2_nand2b_1 _3205_ (.Y(_0910_),
    .B(\MemCell.prescale_reg[2][6] ),
    .A_N(\pwm_module.prescaler2[22] ));
 sg13g2_nor2_1 _3206_ (.A(_1860_),
    .B(\pwm_module.prescaler2[21] ),
    .Y(_0911_));
 sg13g2_nand4_1 _3207_ (.B(_0907_),
    .C(_0909_),
    .A(_0906_),
    .Y(_0912_),
    .D(_0910_));
 sg13g2_nor2_1 _3208_ (.A(_0911_),
    .B(_0912_),
    .Y(_0913_));
 sg13g2_nor2b_1 _3209_ (.A(\MemCell.prescale_reg[2][4] ),
    .B_N(\pwm_module.prescaler2[20] ),
    .Y(_0914_));
 sg13g2_a21o_1 _3210_ (.A2(\pwm_module.prescaler2[21] ),
    .A1(_1860_),
    .B1(_0914_),
    .X(_0915_));
 sg13g2_nor2_1 _3211_ (.A(_1862_),
    .B(\pwm_module.prescaler2[20] ),
    .Y(_0916_));
 sg13g2_nor4_1 _3212_ (.A(_0911_),
    .B(_0912_),
    .C(_0915_),
    .D(_0916_),
    .Y(_0917_));
 sg13g2_nand2b_1 _3213_ (.Y(_0918_),
    .B(\pwm_module.prescaler2[19] ),
    .A_N(net653));
 sg13g2_nand2b_1 _3214_ (.Y(_0919_),
    .B(\pwm_module.prescaler2[18] ),
    .A_N(\MemCell.prescale_reg[2][2] ));
 sg13g2_nand2b_1 _3215_ (.Y(_0920_),
    .B(\MemCell.prescale_reg[2][2] ),
    .A_N(\pwm_module.prescaler2[18] ));
 sg13g2_nor2b_1 _3216_ (.A(\pwm_module.prescaler2[19] ),
    .B_N(net653),
    .Y(_0921_));
 sg13g2_nand2b_1 _3217_ (.Y(_0922_),
    .B(net653),
    .A_N(\pwm_module.prescaler2[19] ));
 sg13g2_and4_1 _3218_ (.A(_0918_),
    .B(_0919_),
    .C(_0920_),
    .D(_0922_),
    .X(_0923_));
 sg13g2_nand2b_1 _3219_ (.Y(_0924_),
    .B(\pwm_module.prescaler2[16] ),
    .A_N(\MemCell.prescale_reg[2][0] ));
 sg13g2_nand2b_1 _3220_ (.Y(_0925_),
    .B(\pwm_module.prescaler2[17] ),
    .A_N(\MemCell.prescale_reg[2][1] ));
 sg13g2_nand2_1 _3221_ (.Y(_0926_),
    .A(_0924_),
    .B(_0925_));
 sg13g2_nor2b_1 _3222_ (.A(\pwm_module.prescaler2[17] ),
    .B_N(\MemCell.prescale_reg[2][1] ),
    .Y(_0927_));
 sg13g2_nand2b_1 _3223_ (.Y(_0928_),
    .B(\MemCell.prescale_reg[2][0] ),
    .A_N(\pwm_module.prescaler2[16] ));
 sg13g2_nand2b_1 _3224_ (.Y(_0929_),
    .B(\pwm_module.prescaler2[31] ),
    .A_N(\MemCell.prescale_reg[3][7] ));
 sg13g2_nand2b_1 _3225_ (.Y(_0930_),
    .B(\pwm_module.prescaler2[30] ),
    .A_N(\MemCell.prescale_reg[3][6] ));
 sg13g2_nand2b_1 _3226_ (.Y(_0931_),
    .B(\pwm_module.prescaler2[29] ),
    .A_N(\MemCell.prescale_reg[3][5] ));
 sg13g2_nand2b_1 _3227_ (.Y(_0932_),
    .B(\pwm_module.prescaler2[28] ),
    .A_N(\MemCell.prescale_reg[3][4] ));
 sg13g2_nand4_1 _3228_ (.B(_0930_),
    .C(_0931_),
    .A(_0929_),
    .Y(_0933_),
    .D(_0932_));
 sg13g2_nand2b_1 _3229_ (.Y(_0934_),
    .B(\MemCell.prescale_reg[3][7] ),
    .A_N(\pwm_module.prescaler2[31] ));
 sg13g2_o21ai_1 _3230_ (.B1(_0934_),
    .Y(_0935_),
    .A1(_1856_),
    .A2(\pwm_module.prescaler2[28] ));
 sg13g2_nand2b_1 _3231_ (.Y(_0936_),
    .B(\MemCell.prescale_reg[3][5] ),
    .A_N(\pwm_module.prescaler2[29] ));
 sg13g2_o21ai_1 _3232_ (.B1(_0936_),
    .Y(_0937_),
    .A1(_1855_),
    .A2(\pwm_module.prescaler2[30] ));
 sg13g2_nor3_1 _3233_ (.A(_0933_),
    .B(_0935_),
    .C(_0937_),
    .Y(_0938_));
 sg13g2_nor2b_1 _3234_ (.A(\MemCell.prescale_reg[3][3] ),
    .B_N(\pwm_module.prescaler2[27] ),
    .Y(_0939_));
 sg13g2_nor2b_1 _3235_ (.A(\MemCell.prescale_reg[3][2] ),
    .B_N(\pwm_module.prescaler2[26] ),
    .Y(_0940_));
 sg13g2_nor2_1 _3236_ (.A(_0939_),
    .B(_0940_),
    .Y(_0941_));
 sg13g2_nor2b_1 _3237_ (.A(\MemCell.prescale_reg[3][1] ),
    .B_N(\pwm_module.prescaler2[25] ),
    .Y(_0942_));
 sg13g2_nor2b_1 _3238_ (.A(\MemCell.prescale_reg[3][0] ),
    .B_N(\pwm_module.prescaler2[24] ),
    .Y(_0943_));
 sg13g2_nor4_1 _3239_ (.A(_0939_),
    .B(_0940_),
    .C(_0942_),
    .D(_0943_),
    .Y(_0944_));
 sg13g2_nand2b_1 _3240_ (.Y(_0945_),
    .B(\MemCell.prescale_reg[3][2] ),
    .A_N(\pwm_module.prescaler2[26] ));
 sg13g2_o21ai_1 _3241_ (.B1(_0945_),
    .Y(_0946_),
    .A1(_1858_),
    .A2(\pwm_module.prescaler2[25] ));
 sg13g2_nor2b_1 _3242_ (.A(\pwm_module.prescaler2[24] ),
    .B_N(\MemCell.prescale_reg[3][0] ),
    .Y(_0947_));
 sg13g2_nor2_1 _3243_ (.A(_1857_),
    .B(\pwm_module.prescaler2[27] ),
    .Y(_0948_));
 sg13g2_nor3_1 _3244_ (.A(_0946_),
    .B(_0947_),
    .C(_0948_),
    .Y(_0949_));
 sg13g2_nand3_1 _3245_ (.B(_0944_),
    .C(_0949_),
    .A(_0938_),
    .Y(_0950_));
 sg13g2_nand3_1 _3246_ (.B(_0923_),
    .C(_0928_),
    .A(_0917_),
    .Y(_0951_));
 sg13g2_nor4_1 _3247_ (.A(_0926_),
    .B(_0927_),
    .C(_0950_),
    .D(_0951_),
    .Y(_0952_));
 sg13g2_a21oi_1 _3248_ (.A1(_0924_),
    .A2(_0925_),
    .Y(_0953_),
    .B1(_0927_));
 sg13g2_a21oi_1 _3249_ (.A1(_0918_),
    .A2(_0919_),
    .Y(_0954_),
    .B1(_0921_));
 sg13g2_a21o_1 _3250_ (.A2(_0953_),
    .A1(_0923_),
    .B1(_0954_),
    .X(_0955_));
 sg13g2_and2_1 _3251_ (.A(_0908_),
    .B(_0909_),
    .X(_0956_));
 sg13g2_a221oi_1 _3252_ (.B2(_0955_),
    .C1(_0956_),
    .B1(_0917_),
    .A1(_0913_),
    .Y(_0957_),
    .A2(_0915_));
 sg13g2_a21o_1 _3253_ (.A2(_0932_),
    .A1(_0931_),
    .B1(_0937_),
    .X(_0958_));
 sg13g2_nand3_1 _3254_ (.B(_0930_),
    .C(_0958_),
    .A(_0929_),
    .Y(_0959_));
 sg13g2_a21oi_1 _3255_ (.A1(_0941_),
    .A2(_0946_),
    .Y(_0960_),
    .B1(_0944_));
 sg13g2_nand3b_1 _3256_ (.B(_0960_),
    .C(_0938_),
    .Y(_0961_),
    .A_N(_0948_));
 sg13g2_o21ai_1 _3257_ (.B1(_0961_),
    .Y(_0962_),
    .A1(_0950_),
    .A2(_0957_));
 sg13g2_a221oi_1 _3258_ (.B2(_0934_),
    .C1(_0962_),
    .B1(_0959_),
    .A1(_0905_),
    .Y(_0963_),
    .A2(_0952_));
 sg13g2_nand2_2 _3259_ (.Y(_0964_),
    .A(net651),
    .B(net612));
 sg13g2_nor2_1 _3260_ (.A(net101),
    .B(net596),
    .Y(_0064_));
 sg13g2_xnor2_1 _3261_ (.Y(_0965_),
    .A(net384),
    .B(net101));
 sg13g2_nor2_1 _3262_ (.A(net596),
    .B(_0965_),
    .Y(_0075_));
 sg13g2_and3_1 _3263_ (.X(_0966_),
    .A(net102),
    .B(\pwm_module.prescaler2[1] ),
    .C(net101));
 sg13g2_a21oi_1 _3264_ (.A1(\pwm_module.prescaler2[1] ),
    .A2(net101),
    .Y(_0967_),
    .B1(net102));
 sg13g2_nor3_1 _3265_ (.A(net596),
    .B(_0966_),
    .C(net103),
    .Y(_0086_));
 sg13g2_and4_2 _3266_ (.A(net207),
    .B(net102),
    .C(\pwm_module.prescaler2[1] ),
    .D(\pwm_module.prescaler2[0] ),
    .X(_0968_));
 sg13g2_nor2_1 _3267_ (.A(net207),
    .B(_0966_),
    .Y(_0969_));
 sg13g2_nor3_1 _3268_ (.A(net596),
    .B(_0968_),
    .C(net208),
    .Y(_0089_));
 sg13g2_nor2_1 _3269_ (.A(net388),
    .B(_0968_),
    .Y(_0970_));
 sg13g2_and2_1 _3270_ (.A(net388),
    .B(_0968_),
    .X(_0971_));
 sg13g2_nor3_1 _3271_ (.A(net596),
    .B(net389),
    .C(_0971_),
    .Y(_0090_));
 sg13g2_nor2_1 _3272_ (.A(net310),
    .B(_0971_),
    .Y(_0972_));
 sg13g2_and2_1 _3273_ (.A(\pwm_module.prescaler2[5] ),
    .B(\pwm_module.prescaler2[4] ),
    .X(_0973_));
 sg13g2_and2_1 _3274_ (.A(_0968_),
    .B(_0973_),
    .X(_0974_));
 sg13g2_nor3_1 _3275_ (.A(net596),
    .B(net311),
    .C(_0974_),
    .Y(_0091_));
 sg13g2_xnor2_1 _3276_ (.Y(_0975_),
    .A(net355),
    .B(_0974_));
 sg13g2_nor2_1 _3277_ (.A(net596),
    .B(_0975_),
    .Y(_0092_));
 sg13g2_a21oi_1 _3278_ (.A1(\pwm_module.prescaler2[6] ),
    .A2(_0974_),
    .Y(_0976_),
    .B1(net80));
 sg13g2_and4_2 _3279_ (.A(net80),
    .B(net560),
    .C(_0968_),
    .D(_0973_),
    .X(_0977_));
 sg13g2_nor3_1 _3280_ (.A(net596),
    .B(net81),
    .C(_0977_),
    .Y(_0093_));
 sg13g2_xnor2_1 _3281_ (.Y(_0978_),
    .A(net347),
    .B(_0977_));
 sg13g2_nor2_1 _3282_ (.A(net597),
    .B(_0978_),
    .Y(_0094_));
 sg13g2_a21oi_1 _3283_ (.A1(\pwm_module.prescaler2[8] ),
    .A2(_0977_),
    .Y(_0979_),
    .B1(net110));
 sg13g2_and2_1 _3284_ (.A(\pwm_module.prescaler2[9] ),
    .B(\pwm_module.prescaler2[8] ),
    .X(_0980_));
 sg13g2_and2_1 _3285_ (.A(_0977_),
    .B(_0980_),
    .X(_0981_));
 sg13g2_nor3_1 _3286_ (.A(net597),
    .B(net111),
    .C(_0981_),
    .Y(_0095_));
 sg13g2_xnor2_1 _3287_ (.Y(_0982_),
    .A(net372),
    .B(_0981_));
 sg13g2_nor2_1 _3288_ (.A(net597),
    .B(_0982_),
    .Y(_0065_));
 sg13g2_a21oi_1 _3289_ (.A1(\pwm_module.prescaler2[10] ),
    .A2(_0981_),
    .Y(_0983_),
    .B1(net219));
 sg13g2_and3_1 _3290_ (.X(_0984_),
    .A(net219),
    .B(\pwm_module.prescaler2[10] ),
    .C(_0981_));
 sg13g2_nand4_1 _3291_ (.B(\pwm_module.prescaler2[10] ),
    .C(_0977_),
    .A(\pwm_module.prescaler2[11] ),
    .Y(_0985_),
    .D(_0980_));
 sg13g2_nor3_1 _3292_ (.A(net597),
    .B(net220),
    .C(_0984_),
    .Y(_0066_));
 sg13g2_xor2_1 _3293_ (.B(_0985_),
    .A(net393),
    .X(_0986_));
 sg13g2_nor2_1 _3294_ (.A(net600),
    .B(_0986_),
    .Y(_0067_));
 sg13g2_a21oi_1 _3295_ (.A1(\pwm_module.prescaler2[12] ),
    .A2(_0984_),
    .Y(_0987_),
    .B1(net249));
 sg13g2_nand2_2 _3296_ (.Y(_0988_),
    .A(net249),
    .B(net561));
 sg13g2_nor2_1 _3297_ (.A(_0985_),
    .B(_0988_),
    .Y(_0989_));
 sg13g2_nor3_1 _3298_ (.A(net600),
    .B(net250),
    .C(_0989_),
    .Y(_0068_));
 sg13g2_nor2_1 _3299_ (.A(net318),
    .B(_0989_),
    .Y(_0990_));
 sg13g2_and2_1 _3300_ (.A(net318),
    .B(_0989_),
    .X(_0991_));
 sg13g2_nor3_1 _3301_ (.A(net600),
    .B(net319),
    .C(_0991_),
    .Y(_0069_));
 sg13g2_nor2_1 _3302_ (.A(net231),
    .B(_0991_),
    .Y(_0992_));
 sg13g2_nand2_1 _3303_ (.Y(_0993_),
    .A(net231),
    .B(net318));
 sg13g2_nor3_2 _3304_ (.A(_0985_),
    .B(_0988_),
    .C(_0993_),
    .Y(_0994_));
 sg13g2_nor3_1 _3305_ (.A(net600),
    .B(net232),
    .C(_0994_),
    .Y(_0070_));
 sg13g2_nor2_1 _3306_ (.A(net327),
    .B(_0994_),
    .Y(_0995_));
 sg13g2_and2_1 _3307_ (.A(net327),
    .B(_0994_),
    .X(_0996_));
 sg13g2_nor3_1 _3308_ (.A(net600),
    .B(net328),
    .C(_0996_),
    .Y(_0071_));
 sg13g2_nor2_1 _3309_ (.A(net286),
    .B(_0996_),
    .Y(_0997_));
 sg13g2_and2_1 _3310_ (.A(net286),
    .B(_0996_),
    .X(_0998_));
 sg13g2_nor3_1 _3311_ (.A(net600),
    .B(net287),
    .C(_0998_),
    .Y(_0072_));
 sg13g2_nor2_1 _3312_ (.A(net273),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_a21oi_1 _3313_ (.A1(net273),
    .A2(_0998_),
    .Y(_1000_),
    .B1(net599));
 sg13g2_nor2b_1 _3314_ (.A(net274),
    .B_N(_1000_),
    .Y(_0073_));
 sg13g2_a21oi_1 _3315_ (.A1(\pwm_module.prescaler2[18] ),
    .A2(_0998_),
    .Y(_1001_),
    .B1(net225));
 sg13g2_nand4_1 _3316_ (.B(\pwm_module.prescaler2[18] ),
    .C(\pwm_module.prescaler2[17] ),
    .A(net225),
    .Y(_1002_),
    .D(\pwm_module.prescaler2[16] ));
 sg13g2_nor4_2 _3317_ (.A(_0985_),
    .B(_0988_),
    .C(_0993_),
    .Y(_1003_),
    .D(_1002_));
 sg13g2_nor3_1 _3318_ (.A(net599),
    .B(net226),
    .C(_1003_),
    .Y(_0074_));
 sg13g2_nor2_1 _3319_ (.A(net275),
    .B(_1003_),
    .Y(_1004_));
 sg13g2_and2_1 _3320_ (.A(net275),
    .B(_1003_),
    .X(_1005_));
 sg13g2_nor3_1 _3321_ (.A(net599),
    .B(net276),
    .C(_1005_),
    .Y(_0076_));
 sg13g2_nor2_1 _3322_ (.A(net256),
    .B(_1005_),
    .Y(_1006_));
 sg13g2_and2_1 _3323_ (.A(net256),
    .B(_1005_),
    .X(_1007_));
 sg13g2_nor3_1 _3324_ (.A(net598),
    .B(net257),
    .C(_1007_),
    .Y(_0077_));
 sg13g2_nor2_1 _3325_ (.A(net281),
    .B(_1007_),
    .Y(_1008_));
 sg13g2_and2_1 _3326_ (.A(net281),
    .B(_1007_),
    .X(_1009_));
 sg13g2_nor3_1 _3327_ (.A(net598),
    .B(_1008_),
    .C(_1009_),
    .Y(_0078_));
 sg13g2_nor2_1 _3328_ (.A(net237),
    .B(_1009_),
    .Y(_1010_));
 sg13g2_and4_1 _3329_ (.A(\pwm_module.prescaler2[23] ),
    .B(\pwm_module.prescaler2[22] ),
    .C(\pwm_module.prescaler2[21] ),
    .D(\pwm_module.prescaler2[20] ),
    .X(_1011_));
 sg13g2_and2_1 _3330_ (.A(_1003_),
    .B(_1011_),
    .X(_1012_));
 sg13g2_nor3_1 _3331_ (.A(net599),
    .B(net238),
    .C(_1012_),
    .Y(_0079_));
 sg13g2_nor2_1 _3332_ (.A(net359),
    .B(_1012_),
    .Y(_1013_));
 sg13g2_and2_1 _3333_ (.A(net359),
    .B(_1012_),
    .X(_1014_));
 sg13g2_nor3_1 _3334_ (.A(net599),
    .B(_1013_),
    .C(_1014_),
    .Y(_0080_));
 sg13g2_nor2_1 _3335_ (.A(net306),
    .B(_1014_),
    .Y(_1015_));
 sg13g2_and3_1 _3336_ (.X(_1016_),
    .A(net306),
    .B(\pwm_module.prescaler2[24] ),
    .C(_1012_));
 sg13g2_nor3_1 _3337_ (.A(net599),
    .B(net307),
    .C(_1016_),
    .Y(_0081_));
 sg13g2_nor2_1 _3338_ (.A(net247),
    .B(_1016_),
    .Y(_1017_));
 sg13g2_and2_1 _3339_ (.A(net247),
    .B(_1016_),
    .X(_1018_));
 sg13g2_nor3_1 _3340_ (.A(net598),
    .B(net248),
    .C(_1018_),
    .Y(_0082_));
 sg13g2_nor2_1 _3341_ (.A(net228),
    .B(_1018_),
    .Y(_1019_));
 sg13g2_and4_1 _3342_ (.A(\pwm_module.prescaler2[27] ),
    .B(\pwm_module.prescaler2[26] ),
    .C(\pwm_module.prescaler2[25] ),
    .D(\pwm_module.prescaler2[24] ),
    .X(_1020_));
 sg13g2_and2_1 _3343_ (.A(_1012_),
    .B(_1020_),
    .X(_1021_));
 sg13g2_nor3_1 _3344_ (.A(net598),
    .B(net229),
    .C(_1021_),
    .Y(_0083_));
 sg13g2_nor2_1 _3345_ (.A(net251),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_and2_1 _3346_ (.A(net251),
    .B(_1021_),
    .X(_1023_));
 sg13g2_nor3_1 _3347_ (.A(net598),
    .B(_1022_),
    .C(_1023_),
    .Y(_0084_));
 sg13g2_nor2_1 _3348_ (.A(net200),
    .B(_1023_),
    .Y(_1024_));
 sg13g2_and3_1 _3349_ (.X(_1025_),
    .A(net200),
    .B(\pwm_module.prescaler2[28] ),
    .C(_1021_));
 sg13g2_nor3_1 _3350_ (.A(net598),
    .B(net201),
    .C(_1025_),
    .Y(_0085_));
 sg13g2_nor2_1 _3351_ (.A(net245),
    .B(_1025_),
    .Y(_1026_));
 sg13g2_a21oi_1 _3352_ (.A1(net245),
    .A2(_1025_),
    .Y(_1027_),
    .B1(net598));
 sg13g2_nor2b_1 _3353_ (.A(net246),
    .B_N(_1027_),
    .Y(_0087_));
 sg13g2_a21oi_1 _3354_ (.A1(\pwm_module.prescaler2[30] ),
    .A2(_1025_),
    .Y(_1028_),
    .B1(net39));
 sg13g2_nor2_1 _3355_ (.A(net598),
    .B(net40),
    .Y(_0088_));
 sg13g2_nor2b_1 _3356_ (.A(\MemCell.curr_state[1] ),
    .B_N(\MemCell.curr_state[0] ),
    .Y(_1029_));
 sg13g2_and2_1 _3357_ (.A(\MemCell.curr_state[2] ),
    .B(_1029_),
    .X(_1030_));
 sg13g2_nand2_1 _3358_ (.Y(_1031_),
    .A(\MemCell.curr_state[0] ),
    .B(\MemCell.curr_state[1] ));
 sg13g2_nor2_1 _3359_ (.A(\MemCell.curr_state[2] ),
    .B(_1031_),
    .Y(_1032_));
 sg13g2_o21ai_1 _3360_ (.B1(_1029_),
    .Y(_1033_),
    .A1(\MemCell.curr_state[2] ),
    .A2(_0102_));
 sg13g2_nand2b_1 _3361_ (.Y(_1034_),
    .B(_1033_),
    .A_N(_1032_));
 sg13g2_and2_1 _3362_ (.A(net650),
    .B(\MemCell.counter[1] ),
    .X(_1035_));
 sg13g2_nand2_2 _3363_ (.Y(_1036_),
    .A(net650),
    .B(\MemCell.counter[1] ));
 sg13g2_nand2_1 _3364_ (.Y(_1037_),
    .A(\MemCell.o_RX_DV ),
    .B(_1035_));
 sg13g2_nand2_1 _3365_ (.Y(_1038_),
    .A(_1034_),
    .B(_1037_));
 sg13g2_nor3_1 _3366_ (.A(\MemCell.curr_state[0] ),
    .B(\MemCell.curr_state[1] ),
    .C(net550),
    .Y(_1039_));
 sg13g2_nor2_1 _3367_ (.A(_1034_),
    .B(_1039_),
    .Y(_1040_));
 sg13g2_nor2_1 _3368_ (.A(\MemCell.curr_state[0] ),
    .B(_1845_),
    .Y(_1041_));
 sg13g2_nand2_1 _3369_ (.Y(_1042_),
    .A(net550),
    .B(_1041_));
 sg13g2_or2_1 _3370_ (.X(_1043_),
    .B(_1031_),
    .A(_0102_));
 sg13g2_o21ai_1 _3371_ (.B1(_1041_),
    .Y(_1044_),
    .A1(\MemCell.curr_state[2] ),
    .A2(net550));
 sg13g2_nand4_1 _3372_ (.B(_1040_),
    .C(_1043_),
    .A(\MemCell.o_RX_DV ),
    .Y(_1045_),
    .D(_1044_));
 sg13g2_or2_1 _3373_ (.X(_1046_),
    .B(net661),
    .A(net669));
 sg13g2_nor4_2 _3374_ (.A(net666),
    .B(net655),
    .C(net660),
    .Y(_1047_),
    .D(_1046_));
 sg13g2_nand2_1 _3375_ (.Y(_1048_),
    .A(net675),
    .B(net671));
 sg13g2_xnor2_1 _3376_ (.Y(_1049_),
    .A(net680),
    .B(_1048_));
 sg13g2_nand2_1 _3377_ (.Y(_1050_),
    .A(_1047_),
    .B(_1049_));
 sg13g2_o21ai_1 _3378_ (.B1(_1038_),
    .Y(\MemCell.next_state[0] ),
    .A1(net551),
    .A2(_1050_));
 sg13g2_nand2b_1 _3379_ (.Y(_1051_),
    .B(_1042_),
    .A_N(_1032_));
 sg13g2_nand2_1 _3380_ (.Y(_1052_),
    .A(_1037_),
    .B(_1051_));
 sg13g2_nand2_1 _3381_ (.Y(_1053_),
    .A(net674),
    .B(_1047_));
 sg13g2_o21ai_1 _3382_ (.B1(_1052_),
    .Y(\MemCell.next_state[1] ),
    .A1(net551),
    .A2(_1053_));
 sg13g2_o21ai_1 _3383_ (.B1(_1037_),
    .Y(_1054_),
    .A1(_1030_),
    .A2(_1039_));
 sg13g2_nand2_1 _3384_ (.Y(_1055_),
    .A(net671),
    .B(_1047_));
 sg13g2_o21ai_1 _3385_ (.B1(_1054_),
    .Y(\MemCell.next_state[2] ),
    .A1(net551),
    .A2(_1055_));
 sg13g2_nand2b_1 _3386_ (.Y(_1056_),
    .B(\pwm_module.counter0[1] ),
    .A_N(\MemCell.dc1_reg[0][1] ));
 sg13g2_nor2b_1 _3387_ (.A(\pwm_module.counter0[0] ),
    .B_N(\MemCell.dc1_reg[0][0] ),
    .Y(_1057_));
 sg13g2_nor2b_1 _3388_ (.A(\pwm_module.counter0[1] ),
    .B_N(\MemCell.dc1_reg[0][1] ),
    .Y(_1058_));
 sg13g2_a221oi_1 _3389_ (.B2(_1057_),
    .C1(_1058_),
    .B1(_1056_),
    .A1(_1916_),
    .Y(_1059_),
    .A2(\MemCell.dc1_reg[0][2] ));
 sg13g2_nand2b_1 _3390_ (.Y(_1060_),
    .B(\pwm_module.counter0[3] ),
    .A_N(\MemCell.dc1_reg[0][3] ));
 sg13g2_o21ai_1 _3391_ (.B1(_1060_),
    .Y(_1061_),
    .A1(_1916_),
    .A2(\MemCell.dc1_reg[0][2] ));
 sg13g2_a22oi_1 _3392_ (.Y(_1062_),
    .B1(\MemCell.dc1_reg[0][3] ),
    .B2(_1915_),
    .A2(\MemCell.dc1_reg[0][4] ),
    .A1(_1913_));
 sg13g2_o21ai_1 _3393_ (.B1(_1062_),
    .Y(_1063_),
    .A1(_1059_),
    .A2(_1061_));
 sg13g2_a22oi_1 _3394_ (.Y(_1064_),
    .B1(_1938_),
    .B2(\pwm_module.counter0[4] ),
    .A2(_1937_),
    .A1(net681));
 sg13g2_nand2b_1 _3395_ (.Y(_1065_),
    .B(\MemCell.dc1_reg[0][6] ),
    .A_N(\pwm_module.counter0[6] ));
 sg13g2_o21ai_1 _3396_ (.B1(_1065_),
    .Y(_1066_),
    .A1(net681),
    .A2(_1937_));
 sg13g2_a21oi_1 _3397_ (.A1(_1063_),
    .A2(_1064_),
    .Y(_1067_),
    .B1(_1066_));
 sg13g2_nand2b_1 _3398_ (.Y(_1068_),
    .B(\pwm_module.counter0[6] ),
    .A_N(\MemCell.dc1_reg[0][6] ));
 sg13g2_o21ai_1 _3399_ (.B1(_1068_),
    .Y(_1069_),
    .A1(_1909_),
    .A2(\MemCell.dc1_reg[0][7] ));
 sg13g2_a22oi_1 _3400_ (.Y(_1070_),
    .B1(\MemCell.dc1_reg[0][7] ),
    .B2(_1909_),
    .A2(\MemCell.dc1_reg[1][0] ),
    .A1(_1907_));
 sg13g2_o21ai_1 _3401_ (.B1(_1070_),
    .Y(_1071_),
    .A1(_1067_),
    .A2(_1069_));
 sg13g2_a22oi_1 _3402_ (.Y(_1072_),
    .B1(_1936_),
    .B2(\pwm_module.counter0[8] ),
    .A2(_1935_),
    .A1(\pwm_module.counter0[9] ));
 sg13g2_nor2_1 _3403_ (.A(\pwm_module.counter0[10] ),
    .B(_1934_),
    .Y(_1073_));
 sg13g2_a221oi_1 _3404_ (.B2(_1072_),
    .C1(_1073_),
    .B1(_1071_),
    .A1(_1905_),
    .Y(_1074_),
    .A2(\MemCell.dc1_reg[1][1] ));
 sg13g2_a221oi_1 _3405_ (.B2(\pwm_module.counter0[10] ),
    .C1(_1074_),
    .B1(_1934_),
    .A1(\pwm_module.counter0[11] ),
    .Y(_1075_),
    .A2(_1933_));
 sg13g2_nand2_1 _3406_ (.Y(_1076_),
    .A(\pwm_module.counter0[14] ),
    .B(_1932_));
 sg13g2_o21ai_1 _3407_ (.B1(_1076_),
    .Y(_1077_),
    .A1(_1898_),
    .A2(\MemCell.dc1_reg[1][7] ));
 sg13g2_nand2_1 _3408_ (.Y(_1078_),
    .A(_1898_),
    .B(\MemCell.dc1_reg[1][7] ));
 sg13g2_o21ai_1 _3409_ (.B1(_1078_),
    .Y(_1079_),
    .A1(\pwm_module.counter0[14] ),
    .A2(_1932_));
 sg13g2_nor2b_1 _3410_ (.A(\pwm_module.counter0[13] ),
    .B_N(\MemCell.dc1_reg[1][5] ),
    .Y(_1080_));
 sg13g2_nor3_1 _3411_ (.A(_1077_),
    .B(_1079_),
    .C(_1080_),
    .Y(_1081_));
 sg13g2_nand2b_1 _3412_ (.Y(_1082_),
    .B(\pwm_module.counter0[12] ),
    .A_N(\MemCell.dc1_reg[1][4] ));
 sg13g2_o21ai_1 _3413_ (.B1(_1082_),
    .Y(_1083_),
    .A1(_1901_),
    .A2(\MemCell.dc1_reg[1][5] ));
 sg13g2_nand2_1 _3414_ (.Y(_1084_),
    .A(_1902_),
    .B(\MemCell.dc1_reg[1][4] ));
 sg13g2_nor2_1 _3415_ (.A(\pwm_module.counter0[11] ),
    .B(_1933_),
    .Y(_1085_));
 sg13g2_nor4_1 _3416_ (.A(_1077_),
    .B(_1079_),
    .C(_1083_),
    .D(_1085_),
    .Y(_1086_));
 sg13g2_nand3b_1 _3417_ (.B(_1084_),
    .C(_1086_),
    .Y(_1087_),
    .A_N(_1080_));
 sg13g2_a22oi_1 _3418_ (.Y(_1088_),
    .B1(_1081_),
    .B2(_1083_),
    .A2(_1078_),
    .A1(_1077_));
 sg13g2_o21ai_1 _3419_ (.B1(_1088_),
    .Y(_1089_),
    .A1(_1075_),
    .A2(_1087_));
 sg13g2_nor2_1 _3420_ (.A(_1883_),
    .B(\MemCell.dc1_reg[2][7] ),
    .Y(_1090_));
 sg13g2_nor2_1 _3421_ (.A(_1885_),
    .B(\MemCell.dc1_reg[2][6] ),
    .Y(_1091_));
 sg13g2_nand2_1 _3422_ (.Y(_1092_),
    .A(_1883_),
    .B(\MemCell.dc1_reg[2][7] ));
 sg13g2_o21ai_1 _3423_ (.B1(_1092_),
    .Y(_1093_),
    .A1(\pwm_module.counter0[22] ),
    .A2(_1931_));
 sg13g2_nor3_1 _3424_ (.A(_1090_),
    .B(_1091_),
    .C(_1093_),
    .Y(_1094_));
 sg13g2_nor2b_1 _3425_ (.A(\pwm_module.counter0[20] ),
    .B_N(\MemCell.dc1_reg[2][4] ),
    .Y(_1095_));
 sg13g2_nor2b_1 _3426_ (.A(\pwm_module.counter0[28] ),
    .B_N(\MemCell.dc1_reg[3][4] ),
    .Y(_1096_));
 sg13g2_nor2b_1 _3427_ (.A(\pwm_module.counter0[21] ),
    .B_N(\MemCell.dc1_reg[2][5] ),
    .Y(_1097_));
 sg13g2_nand2b_1 _3428_ (.Y(_1098_),
    .B(\pwm_module.counter0[29] ),
    .A_N(\MemCell.dc1_reg[3][5] ));
 sg13g2_o21ai_1 _3429_ (.B1(_1098_),
    .Y(_1099_),
    .A1(_1874_),
    .A2(\MemCell.dc1_reg[3][4] ));
 sg13g2_nand2b_1 _3430_ (.Y(_1100_),
    .B(\pwm_module.counter0[21] ),
    .A_N(\MemCell.dc1_reg[2][5] ));
 sg13g2_o21ai_1 _3431_ (.B1(_1100_),
    .Y(_1101_),
    .A1(_1888_),
    .A2(\MemCell.dc1_reg[2][4] ));
 sg13g2_a22oi_1 _3432_ (.Y(_1102_),
    .B1(_1929_),
    .B2(\pwm_module.counter0[26] ),
    .A2(_1928_),
    .A1(\pwm_module.counter0[27] ));
 sg13g2_nor2_1 _3433_ (.A(\pwm_module.counter0[27] ),
    .B(_1928_),
    .Y(_1103_));
 sg13g2_o21ai_1 _3434_ (.B1(_1102_),
    .Y(_1104_),
    .A1(\pwm_module.counter0[26] ),
    .A2(_1929_));
 sg13g2_nor2_1 _3435_ (.A(_1103_),
    .B(_1104_),
    .Y(_1105_));
 sg13g2_nand2b_1 _3436_ (.Y(_1106_),
    .B(\pwm_module.counter0[25] ),
    .A_N(\MemCell.dc1_reg[3][1] ));
 sg13g2_o21ai_1 _3437_ (.B1(_1106_),
    .Y(_1107_),
    .A1(_1881_),
    .A2(\MemCell.dc1_reg[3][0] ));
 sg13g2_nand2_1 _3438_ (.Y(_1108_),
    .A(_1879_),
    .B(\MemCell.dc1_reg[3][1] ));
 sg13g2_o21ai_1 _3439_ (.B1(_1108_),
    .Y(_1109_),
    .A1(\pwm_module.counter0[24] ),
    .A2(_1930_));
 sg13g2_nor4_1 _3440_ (.A(_1103_),
    .B(_1104_),
    .C(_1107_),
    .D(_1109_),
    .Y(_1110_));
 sg13g2_a22oi_1 _3441_ (.Y(_1111_),
    .B1(_1927_),
    .B2(\pwm_module.counter0[30] ),
    .A2(_1926_),
    .A1(\pwm_module.counter0[31] ));
 sg13g2_nor2_1 _3442_ (.A(\pwm_module.counter0[31] ),
    .B(_1926_),
    .Y(_1112_));
 sg13g2_nor2b_1 _3443_ (.A(\pwm_module.counter0[29] ),
    .B_N(\MemCell.dc1_reg[3][5] ),
    .Y(_1113_));
 sg13g2_o21ai_1 _3444_ (.B1(_1111_),
    .Y(_1114_),
    .A1(\pwm_module.counter0[30] ),
    .A2(_1927_));
 sg13g2_or2_1 _3445_ (.X(_1115_),
    .B(_1114_),
    .A(_1112_));
 sg13g2_nor2_1 _3446_ (.A(_1113_),
    .B(_1115_),
    .Y(_1116_));
 sg13g2_nor4_2 _3447_ (.A(_1096_),
    .B(_1099_),
    .C(_1113_),
    .Y(_1117_),
    .D(_1115_));
 sg13g2_and2_1 _3448_ (.A(_1110_),
    .B(_1117_),
    .X(_1118_));
 sg13g2_nor3_1 _3449_ (.A(_1095_),
    .B(_1097_),
    .C(_1101_),
    .Y(_1119_));
 sg13g2_nand3_1 _3450_ (.B(_1118_),
    .C(_1119_),
    .A(_1094_),
    .Y(_1120_));
 sg13g2_nand2b_1 _3451_ (.Y(_1121_),
    .B(\pwm_module.counter0[18] ),
    .A_N(\MemCell.dc1_reg[2][2] ));
 sg13g2_nand2b_1 _3452_ (.Y(_1122_),
    .B(\pwm_module.counter0[19] ),
    .A_N(\MemCell.dc1_reg[2][3] ));
 sg13g2_nand2_1 _3453_ (.Y(_1123_),
    .A(_1121_),
    .B(_1122_));
 sg13g2_nand2_1 _3454_ (.Y(_1124_),
    .A(_1890_),
    .B(\MemCell.dc1_reg[2][3] ));
 sg13g2_a22oi_1 _3455_ (.Y(_1125_),
    .B1(\MemCell.dc1_reg[2][1] ),
    .B2(_1894_),
    .A2(\MemCell.dc1_reg[2][2] ),
    .A1(_1892_));
 sg13g2_and4_1 _3456_ (.A(_1121_),
    .B(_1122_),
    .C(_1124_),
    .D(_1125_),
    .X(_1126_));
 sg13g2_nand4_1 _3457_ (.B(_1122_),
    .C(_1124_),
    .A(_1121_),
    .Y(_1127_),
    .D(_1125_));
 sg13g2_nor2b_1 _3458_ (.A(\pwm_module.counter0[16] ),
    .B_N(\MemCell.dc1_reg[2][0] ),
    .Y(_1128_));
 sg13g2_nand2b_1 _3459_ (.Y(_1129_),
    .B(\pwm_module.counter0[16] ),
    .A_N(\MemCell.dc1_reg[2][0] ));
 sg13g2_o21ai_1 _3460_ (.B1(_1129_),
    .Y(_1130_),
    .A1(_1894_),
    .A2(\MemCell.dc1_reg[2][1] ));
 sg13g2_nor4_2 _3461_ (.A(_1120_),
    .B(_1127_),
    .C(_1128_),
    .Y(_1131_),
    .D(_1130_));
 sg13g2_nand3_1 _3462_ (.B(_1107_),
    .C(_1108_),
    .A(_1105_),
    .Y(_1132_));
 sg13g2_o21ai_1 _3463_ (.B1(_1132_),
    .Y(_1133_),
    .A1(_1102_),
    .A2(_1103_));
 sg13g2_o21ai_1 _3464_ (.B1(_1092_),
    .Y(_1134_),
    .A1(_1090_),
    .A2(_1091_));
 sg13g2_nand3b_1 _3465_ (.B(_1101_),
    .C(_1094_),
    .Y(_1135_),
    .A_N(_1097_));
 sg13g2_nand2_1 _3466_ (.Y(_1136_),
    .A(_1134_),
    .B(_1135_));
 sg13g2_a22oi_1 _3467_ (.Y(_1137_),
    .B1(_1126_),
    .B2(_1130_),
    .A2(_1124_),
    .A1(_1123_));
 sg13g2_o21ai_1 _3468_ (.B1(net651),
    .Y(_1138_),
    .A1(_1111_),
    .A2(_1112_));
 sg13g2_a221oi_1 _3469_ (.B2(_1136_),
    .C1(_1138_),
    .B1(_1118_),
    .A1(_1099_),
    .Y(_1139_),
    .A2(_1116_));
 sg13g2_o21ai_1 _3470_ (.B1(_1139_),
    .Y(_1140_),
    .A1(_1120_),
    .A2(_1137_));
 sg13g2_a221oi_1 _3471_ (.B2(_1117_),
    .C1(_1140_),
    .B1(_1133_),
    .A1(_1089_),
    .Y(_0096_),
    .A2(_1131_));
 sg13g2_nand2_2 _3472_ (.Y(_1141_),
    .A(net644),
    .B(_0616_));
 sg13g2_nand2b_1 _3473_ (.Y(_1142_),
    .B(\MemCell.counter_value[14] ),
    .A_N(\pwm_module.counter0[14] ));
 sg13g2_nand2b_1 _3474_ (.Y(_1143_),
    .B(\MemCell.counter_value[13] ),
    .A_N(\pwm_module.counter0[13] ));
 sg13g2_nand2b_1 _3475_ (.Y(_1144_),
    .B(\MemCell.counter_value[15] ),
    .A_N(\pwm_module.counter0[15] ));
 sg13g2_nand2b_1 _3476_ (.Y(_1145_),
    .B(\MemCell.counter_value[12] ),
    .A_N(\pwm_module.counter0[12] ));
 sg13g2_nand4_1 _3477_ (.B(_1143_),
    .C(_1144_),
    .A(_1142_),
    .Y(_1146_),
    .D(_1145_));
 sg13g2_nand2b_1 _3478_ (.Y(_1147_),
    .B(\pwm_module.counter0[14] ),
    .A_N(\MemCell.counter_value[14] ));
 sg13g2_o21ai_1 _3479_ (.B1(_1147_),
    .Y(_1148_),
    .A1(_1898_),
    .A2(\MemCell.counter_value[15] ));
 sg13g2_nand2b_1 _3480_ (.Y(_1149_),
    .B(\pwm_module.counter0[13] ),
    .A_N(\MemCell.counter_value[13] ));
 sg13g2_o21ai_1 _3481_ (.B1(_1149_),
    .Y(_1150_),
    .A1(_1902_),
    .A2(\MemCell.counter_value[12] ));
 sg13g2_nor2b_1 _3482_ (.A(_1148_),
    .B_N(_1144_),
    .Y(_1151_));
 sg13g2_nor3_2 _3483_ (.A(_1146_),
    .B(_1148_),
    .C(_1150_),
    .Y(_1152_));
 sg13g2_nand2b_1 _3484_ (.Y(_1153_),
    .B(\pwm_module.counter0[10] ),
    .A_N(\MemCell.counter_value[10] ));
 sg13g2_nand2b_1 _3485_ (.Y(_1154_),
    .B(\pwm_module.counter0[11] ),
    .A_N(\MemCell.counter_value[11] ));
 sg13g2_nand2_1 _3486_ (.Y(_1155_),
    .A(_1153_),
    .B(_1154_));
 sg13g2_nand2b_1 _3487_ (.Y(_1156_),
    .B(\MemCell.counter_value[11] ),
    .A_N(\pwm_module.counter0[11] ));
 sg13g2_nand2b_1 _3488_ (.Y(_1157_),
    .B(\pwm_module.counter0[8] ),
    .A_N(\MemCell.counter_value[8] ));
 sg13g2_nand2b_1 _3489_ (.Y(_1158_),
    .B(\pwm_module.counter0[9] ),
    .A_N(\MemCell.counter_value[9] ));
 sg13g2_and2_1 _3490_ (.A(_1157_),
    .B(_1158_),
    .X(_1159_));
 sg13g2_nand2b_1 _3491_ (.Y(_1160_),
    .B(\MemCell.counter_value[10] ),
    .A_N(\pwm_module.counter0[10] ));
 sg13g2_nor2b_1 _3492_ (.A(\pwm_module.counter0[9] ),
    .B_N(\MemCell.counter_value[9] ),
    .Y(_1161_));
 sg13g2_and4_1 _3493_ (.A(_1153_),
    .B(_1154_),
    .C(_1156_),
    .D(_1160_),
    .X(_1162_));
 sg13g2_a21oi_1 _3494_ (.A1(_1157_),
    .A2(_1158_),
    .Y(_1163_),
    .B1(_1161_));
 sg13g2_a22oi_1 _3495_ (.Y(_1164_),
    .B1(_1162_),
    .B2(_1163_),
    .A2(_1156_),
    .A1(_1155_));
 sg13g2_nand2b_1 _3496_ (.Y(_1165_),
    .B(\pwm_module.counter0[1] ),
    .A_N(\MemCell.counter_value[1] ));
 sg13g2_nor2b_1 _3497_ (.A(\pwm_module.counter0[0] ),
    .B_N(\MemCell.counter_value[0] ),
    .Y(_1166_));
 sg13g2_nor2b_1 _3498_ (.A(\pwm_module.counter0[1] ),
    .B_N(\MemCell.counter_value[1] ),
    .Y(_1167_));
 sg13g2_a221oi_1 _3499_ (.B2(_1166_),
    .C1(_1167_),
    .B1(_1165_),
    .A1(_1916_),
    .Y(_1168_),
    .A2(\MemCell.counter_value[2] ));
 sg13g2_nand2b_1 _3500_ (.Y(_1169_),
    .B(\pwm_module.counter0[3] ),
    .A_N(\MemCell.counter_value[3] ));
 sg13g2_o21ai_1 _3501_ (.B1(_1169_),
    .Y(_1170_),
    .A1(_1916_),
    .A2(\MemCell.counter_value[2] ));
 sg13g2_a22oi_1 _3502_ (.Y(_1171_),
    .B1(_1915_),
    .B2(\MemCell.counter_value[3] ),
    .A2(\MemCell.counter_value[4] ),
    .A1(_1913_));
 sg13g2_o21ai_1 _3503_ (.B1(_1171_),
    .Y(_1172_),
    .A1(_1168_),
    .A2(_1170_));
 sg13g2_a22oi_1 _3504_ (.Y(_1173_),
    .B1(\pwm_module.counter0[4] ),
    .B2(_1914_),
    .A2(_1912_),
    .A1(net681));
 sg13g2_nand2b_1 _3505_ (.Y(_1174_),
    .B(\MemCell.counter_value[5] ),
    .A_N(net681));
 sg13g2_o21ai_1 _3506_ (.B1(_1174_),
    .Y(_1175_),
    .A1(\pwm_module.counter0[6] ),
    .A2(_1911_));
 sg13g2_a21o_1 _3507_ (.A2(_1173_),
    .A1(_1172_),
    .B1(_1175_),
    .X(_1176_));
 sg13g2_a22oi_1 _3508_ (.Y(_1177_),
    .B1(\pwm_module.counter0[6] ),
    .B2(_1911_),
    .A2(_1910_),
    .A1(\pwm_module.counter0[7] ));
 sg13g2_a221oi_1 _3509_ (.B2(\MemCell.counter_value[7] ),
    .C1(_1161_),
    .B1(_1909_),
    .A1(_1907_),
    .Y(_1178_),
    .A2(\MemCell.counter_value[8] ));
 sg13g2_nand2_1 _3510_ (.Y(_1179_),
    .A(_1144_),
    .B(_1148_));
 sg13g2_nand4_1 _3511_ (.B(_1143_),
    .C(_1150_),
    .A(_1142_),
    .Y(_1180_),
    .D(_1151_));
 sg13g2_nand4_1 _3512_ (.B(_1159_),
    .C(_1162_),
    .A(_1152_),
    .Y(_1181_),
    .D(_1178_));
 sg13g2_a21oi_2 _3513_ (.B1(_1181_),
    .Y(_1182_),
    .A2(_1177_),
    .A1(_1176_));
 sg13g2_nand2b_1 _3514_ (.Y(_1183_),
    .B(_1152_),
    .A_N(_1164_));
 sg13g2_nand3_1 _3515_ (.B(_1180_),
    .C(_1183_),
    .A(_1179_),
    .Y(_1184_));
 sg13g2_nand2b_1 _3516_ (.Y(_1185_),
    .B(\pwm_module.counter0[30] ),
    .A_N(\MemCell.counter_value[30] ));
 sg13g2_nand2b_1 _3517_ (.Y(_1186_),
    .B(\pwm_module.counter0[31] ),
    .A_N(\MemCell.counter_value[31] ));
 sg13g2_nand2_1 _3518_ (.Y(_1187_),
    .A(_1185_),
    .B(_1186_));
 sg13g2_nand2b_1 _3519_ (.Y(_1188_),
    .B(\MemCell.counter_value[31] ),
    .A_N(\pwm_module.counter0[31] ));
 sg13g2_nand2b_1 _3520_ (.Y(_1189_),
    .B(\MemCell.counter_value[30] ),
    .A_N(\pwm_module.counter0[30] ));
 sg13g2_and4_1 _3521_ (.A(_1185_),
    .B(_1186_),
    .C(_1188_),
    .D(_1189_),
    .X(_1190_));
 sg13g2_a22oi_1 _3522_ (.Y(_1191_),
    .B1(\pwm_module.counter0[28] ),
    .B2(_1875_),
    .A2(_1873_),
    .A1(\pwm_module.counter0[29] ));
 sg13g2_nand2b_1 _3523_ (.Y(_1192_),
    .B(\MemCell.counter_value[29] ),
    .A_N(\pwm_module.counter0[29] ));
 sg13g2_nand2_1 _3524_ (.Y(_1193_),
    .A(_1874_),
    .B(\MemCell.counter_value[28] ));
 sg13g2_and4_2 _3525_ (.A(_1190_),
    .B(_1191_),
    .C(_1192_),
    .D(_1193_),
    .X(_1194_));
 sg13g2_a22oi_1 _3526_ (.Y(_1195_),
    .B1(\pwm_module.counter0[26] ),
    .B2(_1878_),
    .A2(_1876_),
    .A1(\pwm_module.counter0[27] ));
 sg13g2_nor2b_1 _3527_ (.A(\pwm_module.counter0[27] ),
    .B_N(\MemCell.counter_value[27] ),
    .Y(_1196_));
 sg13g2_a221oi_1 _3528_ (.B2(\MemCell.counter_value[25] ),
    .C1(_1196_),
    .B1(_1879_),
    .A1(_1877_),
    .Y(_1197_),
    .A2(\MemCell.counter_value[26] ));
 sg13g2_nand2_1 _3529_ (.Y(_1198_),
    .A(_1195_),
    .B(_1197_));
 sg13g2_nor2_1 _3530_ (.A(\pwm_module.counter0[24] ),
    .B(_1882_),
    .Y(_1199_));
 sg13g2_nand2_1 _3531_ (.Y(_1200_),
    .A(\pwm_module.counter0[25] ),
    .B(_1880_));
 sg13g2_o21ai_1 _3532_ (.B1(_1200_),
    .Y(_1201_),
    .A1(_1881_),
    .A2(\MemCell.counter_value[24] ));
 sg13g2_nor3_1 _3533_ (.A(_1198_),
    .B(_1199_),
    .C(_1201_),
    .Y(_1202_));
 sg13g2_nand2b_1 _3534_ (.Y(_1203_),
    .B(\pwm_module.counter0[18] ),
    .A_N(\MemCell.counter_value[18] ));
 sg13g2_nand2b_1 _3535_ (.Y(_1204_),
    .B(\pwm_module.counter0[19] ),
    .A_N(\MemCell.counter_value[19] ));
 sg13g2_nand2_1 _3536_ (.Y(_1205_),
    .A(_1203_),
    .B(_1204_));
 sg13g2_nand2b_1 _3537_ (.Y(_1206_),
    .B(\MemCell.counter_value[19] ),
    .A_N(\pwm_module.counter0[19] ));
 sg13g2_nand2b_1 _3538_ (.Y(_1207_),
    .B(\MemCell.counter_value[18] ),
    .A_N(\pwm_module.counter0[18] ));
 sg13g2_and4_1 _3539_ (.A(_1203_),
    .B(_1204_),
    .C(_1206_),
    .D(_1207_),
    .X(_1208_));
 sg13g2_nand2b_1 _3540_ (.Y(_1209_),
    .B(\pwm_module.counter0[16] ),
    .A_N(\MemCell.counter_value[16] ));
 sg13g2_nand2b_1 _3541_ (.Y(_1210_),
    .B(\pwm_module.counter0[17] ),
    .A_N(\MemCell.counter_value[17] ));
 sg13g2_nor2b_1 _3542_ (.A(\pwm_module.counter0[17] ),
    .B_N(\MemCell.counter_value[17] ),
    .Y(_1211_));
 sg13g2_a21oi_1 _3543_ (.A1(_1896_),
    .A2(\MemCell.counter_value[16] ),
    .Y(_1212_),
    .B1(_1211_));
 sg13g2_nand4_1 _3544_ (.B(_1209_),
    .C(_1210_),
    .A(_1208_),
    .Y(_1213_),
    .D(_1212_));
 sg13g2_nor2b_1 _3545_ (.A(\pwm_module.counter0[21] ),
    .B_N(\MemCell.counter_value[21] ),
    .Y(_1214_));
 sg13g2_a21o_1 _3546_ (.A2(\MemCell.counter_value[22] ),
    .A1(_1885_),
    .B1(_1214_),
    .X(_1215_));
 sg13g2_nand2b_1 _3547_ (.Y(_1216_),
    .B(\MemCell.counter_value[23] ),
    .A_N(\pwm_module.counter0[23] ));
 sg13g2_o21ai_1 _3548_ (.B1(_1216_),
    .Y(_1217_),
    .A1(\pwm_module.counter0[20] ),
    .A2(_1889_));
 sg13g2_nand2b_1 _3549_ (.Y(_1218_),
    .B(\pwm_module.counter0[20] ),
    .A_N(\MemCell.counter_value[20] ));
 sg13g2_nand2b_1 _3550_ (.Y(_1219_),
    .B(\pwm_module.counter0[21] ),
    .A_N(\MemCell.counter_value[21] ));
 sg13g2_nand2_1 _3551_ (.Y(_1220_),
    .A(_1218_),
    .B(_1219_));
 sg13g2_nand2b_1 _3552_ (.Y(_1221_),
    .B(\pwm_module.counter0[23] ),
    .A_N(\MemCell.counter_value[23] ));
 sg13g2_o21ai_1 _3553_ (.B1(_1221_),
    .Y(_1222_),
    .A1(_1885_),
    .A2(\MemCell.counter_value[22] ));
 sg13g2_or4_1 _3554_ (.A(_1215_),
    .B(_1217_),
    .C(_1220_),
    .D(_1222_),
    .X(_1223_));
 sg13g2_nor2_1 _3555_ (.A(_1213_),
    .B(_1223_),
    .Y(_1224_));
 sg13g2_and3_1 _3556_ (.X(_1225_),
    .A(_1194_),
    .B(_1202_),
    .C(_1224_));
 sg13g2_o21ai_1 _3557_ (.B1(_1225_),
    .Y(_1226_),
    .A1(_1182_),
    .A2(_1184_));
 sg13g2_a221oi_1 _3558_ (.B2(_1219_),
    .C1(_1214_),
    .B1(_1218_),
    .A1(_1885_),
    .Y(_1227_),
    .A2(\MemCell.counter_value[22] ));
 sg13g2_o21ai_1 _3559_ (.B1(_1216_),
    .Y(_1228_),
    .A1(_1222_),
    .A2(_1227_));
 sg13g2_o21ai_1 _3560_ (.B1(_1210_),
    .Y(_1229_),
    .A1(_1209_),
    .A2(_1211_));
 sg13g2_a22oi_1 _3561_ (.Y(_1230_),
    .B1(_1208_),
    .B2(_1229_),
    .A2(_1206_),
    .A1(_1205_));
 sg13g2_o21ai_1 _3562_ (.B1(_1228_),
    .Y(_1231_),
    .A1(_1223_),
    .A2(_1230_));
 sg13g2_nand3_1 _3563_ (.B(_1202_),
    .C(_1231_),
    .A(_1194_),
    .Y(_1232_));
 sg13g2_nor2_1 _3564_ (.A(_1195_),
    .B(_1196_),
    .Y(_1233_));
 sg13g2_nor2b_1 _3565_ (.A(_1198_),
    .B_N(_1201_),
    .Y(_1234_));
 sg13g2_o21ai_1 _3566_ (.B1(_1194_),
    .Y(_1235_),
    .A1(_1233_),
    .A2(_1234_));
 sg13g2_nand3b_1 _3567_ (.B(_1192_),
    .C(_1190_),
    .Y(_1236_),
    .A_N(_1191_));
 sg13g2_nand2_1 _3568_ (.Y(_1237_),
    .A(net651),
    .B(_1236_));
 sg13g2_a21oi_1 _3569_ (.A1(_1187_),
    .A2(_1188_),
    .Y(_1238_),
    .B1(_1237_));
 sg13g2_and3_1 _3570_ (.X(_1239_),
    .A(_1232_),
    .B(_1235_),
    .C(_1238_));
 sg13g2_a22oi_1 _3571_ (.Y(_1240_),
    .B1(_1226_),
    .B2(_1239_),
    .A2(_0616_),
    .A1(net646));
 sg13g2_inv_2 _3572_ (.Y(_1241_),
    .A(net589));
 sg13g2_xnor2_1 _3573_ (.Y(_1242_),
    .A(net396),
    .B(net591));
 sg13g2_nor2_1 _3574_ (.A(net587),
    .B(_1242_),
    .Y(_0108_));
 sg13g2_a21o_1 _3575_ (.A2(net591),
    .A1(net396),
    .B1(net534),
    .X(_1243_));
 sg13g2_nand3_1 _3576_ (.B(net396),
    .C(net591),
    .A(net534),
    .Y(_1244_));
 sg13g2_and3_1 _3577_ (.X(_0109_),
    .A(net568),
    .B(_1243_),
    .C(_1244_));
 sg13g2_and3_1 _3578_ (.X(_1245_),
    .A(net215),
    .B(\pwm_module.counter0[1] ),
    .C(\pwm_module.counter0[0] ));
 sg13g2_a21o_1 _3579_ (.A2(_1245_),
    .A1(net591),
    .B1(net587),
    .X(_1246_));
 sg13g2_a21oi_1 _3580_ (.A1(_1916_),
    .A2(_1244_),
    .Y(_0110_),
    .B1(_1246_));
 sg13g2_nand3_1 _3581_ (.B(net591),
    .C(_1245_),
    .A(net465),
    .Y(_1247_));
 sg13g2_a21o_1 _3582_ (.A2(_1245_),
    .A1(net591),
    .B1(net465),
    .X(_1248_));
 sg13g2_and3_1 _3583_ (.X(_0111_),
    .A(net568),
    .B(_1247_),
    .C(_1248_));
 sg13g2_and3_1 _3584_ (.X(_1249_),
    .A(\pwm_module.counter0[4] ),
    .B(\pwm_module.counter0[3] ),
    .C(_1245_));
 sg13g2_nand3_1 _3585_ (.B(\pwm_module.counter0[3] ),
    .C(_1245_),
    .A(\pwm_module.counter0[4] ),
    .Y(_1250_));
 sg13g2_a21oi_2 _3586_ (.B1(_1250_),
    .Y(_1251_),
    .A2(_0616_),
    .A1(net644));
 sg13g2_a221oi_1 _3587_ (.B2(net591),
    .C1(net587),
    .B1(_1249_),
    .A1(_1913_),
    .Y(_0112_),
    .A2(_1247_));
 sg13g2_xnor2_1 _3588_ (.Y(_1252_),
    .A(net681),
    .B(_1251_));
 sg13g2_nor2_1 _3589_ (.A(net587),
    .B(_1252_),
    .Y(_0113_));
 sg13g2_a21o_1 _3590_ (.A2(_1251_),
    .A1(net425),
    .B1(\pwm_module.counter0[6] ),
    .X(_1253_));
 sg13g2_nand3_1 _3591_ (.B(net681),
    .C(_1251_),
    .A(\pwm_module.counter0[6] ),
    .Y(_1254_));
 sg13g2_and3_1 _3592_ (.X(_0114_),
    .A(net568),
    .B(net426),
    .C(_1254_));
 sg13g2_nand4_1 _3593_ (.B(\pwm_module.counter0[6] ),
    .C(net681),
    .A(\pwm_module.counter0[7] ),
    .Y(_1255_),
    .D(_1249_));
 sg13g2_a21oi_1 _3594_ (.A1(net644),
    .A2(_0616_),
    .Y(_1256_),
    .B1(_1255_));
 sg13g2_or2_1 _3595_ (.X(_1257_),
    .B(net586),
    .A(net587));
 sg13g2_a21oi_1 _3596_ (.A1(_1909_),
    .A2(_1254_),
    .Y(_0115_),
    .B1(_1257_));
 sg13g2_nand2_1 _3597_ (.Y(_1258_),
    .A(net529),
    .B(net586));
 sg13g2_or2_1 _3598_ (.X(_1259_),
    .B(net586),
    .A(net529));
 sg13g2_and3_1 _3599_ (.X(_0116_),
    .A(net568),
    .B(_1258_),
    .C(_1259_));
 sg13g2_and2_1 _3600_ (.A(\pwm_module.counter0[9] ),
    .B(\pwm_module.counter0[8] ),
    .X(_1260_));
 sg13g2_a21o_1 _3601_ (.A2(_1260_),
    .A1(net586),
    .B1(net590),
    .X(_1261_));
 sg13g2_a21oi_1 _3602_ (.A1(_1905_),
    .A2(_1258_),
    .Y(_0117_),
    .B1(_1261_));
 sg13g2_a21oi_1 _3603_ (.A1(net586),
    .A2(_1260_),
    .Y(_1262_),
    .B1(net166));
 sg13g2_and2_1 _3604_ (.A(net166),
    .B(_1260_),
    .X(_1263_));
 sg13g2_a21oi_1 _3605_ (.A1(_1256_),
    .A2(_1263_),
    .Y(_1264_),
    .B1(net590));
 sg13g2_nor2b_1 _3606_ (.A(net167),
    .B_N(_1264_),
    .Y(_0118_));
 sg13g2_a21oi_1 _3607_ (.A1(net586),
    .A2(_1263_),
    .Y(_1265_),
    .B1(net326));
 sg13g2_and2_1 _3608_ (.A(net326),
    .B(_1263_),
    .X(_1266_));
 sg13g2_nand2_1 _3609_ (.Y(_1267_),
    .A(\pwm_module.counter0[11] ),
    .B(_1263_));
 sg13g2_nor2_1 _3610_ (.A(_1255_),
    .B(_1267_),
    .Y(_1268_));
 sg13g2_and2_1 _3611_ (.A(net592),
    .B(_1268_),
    .X(_1269_));
 sg13g2_nor3_1 _3612_ (.A(net587),
    .B(_1265_),
    .C(_1269_),
    .Y(_0119_));
 sg13g2_a21o_1 _3613_ (.A2(_1266_),
    .A1(net586),
    .B1(net422),
    .X(_1270_));
 sg13g2_nand3_1 _3614_ (.B(net592),
    .C(_1268_),
    .A(net422),
    .Y(_1271_));
 sg13g2_and3_1 _3615_ (.X(_0120_),
    .A(net568),
    .B(_1270_),
    .C(_1271_));
 sg13g2_nor2_1 _3616_ (.A(_1901_),
    .B(_1902_),
    .Y(_1272_));
 sg13g2_nand3_1 _3617_ (.B(_1266_),
    .C(_1272_),
    .A(net586),
    .Y(_1273_));
 sg13g2_a221oi_1 _3618_ (.B2(_1269_),
    .C1(net590),
    .B1(_1272_),
    .A1(_1901_),
    .Y(_0121_),
    .A2(_1271_));
 sg13g2_nor3_2 _3619_ (.A(_1899_),
    .B(_1901_),
    .C(_1902_),
    .Y(_1274_));
 sg13g2_nand4_1 _3620_ (.B(\pwm_module.counter0[6] ),
    .C(net681),
    .A(net394),
    .Y(_1275_),
    .D(_1274_));
 sg13g2_nor3_2 _3621_ (.A(_1250_),
    .B(_1267_),
    .C(_1275_),
    .Y(_1276_));
 sg13g2_nand2_1 _3622_ (.Y(_1277_),
    .A(net592),
    .B(_1276_));
 sg13g2_a221oi_1 _3623_ (.B2(net592),
    .C1(net587),
    .B1(_1276_),
    .A1(_1899_),
    .Y(_0122_),
    .A2(_1273_));
 sg13g2_nor4_2 _3624_ (.A(_1898_),
    .B(_1250_),
    .C(_1267_),
    .Y(_1278_),
    .D(_1275_));
 sg13g2_and2_2 _3625_ (.A(net462),
    .B(_1276_),
    .X(_1279_));
 sg13g2_a221oi_1 _3626_ (.B2(net591),
    .C1(net587),
    .B1(_1279_),
    .A1(_1898_),
    .Y(_0123_),
    .A2(_1277_));
 sg13g2_nand3_1 _3627_ (.B(_1268_),
    .C(_1274_),
    .A(\pwm_module.counter0[15] ),
    .Y(_1280_));
 sg13g2_a21oi_1 _3628_ (.A1(net595),
    .A2(_1279_),
    .Y(_1281_),
    .B1(net387));
 sg13g2_nor2_1 _3629_ (.A(_1896_),
    .B(_1280_),
    .Y(_1282_));
 sg13g2_and2_1 _3630_ (.A(net595),
    .B(_1282_),
    .X(_1283_));
 sg13g2_nor3_1 _3631_ (.A(net589),
    .B(_1281_),
    .C(_1283_),
    .Y(_0124_));
 sg13g2_a21o_1 _3632_ (.A2(_1282_),
    .A1(net595),
    .B1(net453),
    .X(_1284_));
 sg13g2_nor2_1 _3633_ (.A(_1894_),
    .B(_1896_),
    .Y(_1285_));
 sg13g2_nand3_1 _3634_ (.B(net595),
    .C(_1282_),
    .A(net453),
    .Y(_1286_));
 sg13g2_and3_1 _3635_ (.X(_0125_),
    .A(_1241_),
    .B(_1284_),
    .C(_1286_));
 sg13g2_nand4_1 _3636_ (.B(net593),
    .C(_1279_),
    .A(\pwm_module.counter0[18] ),
    .Y(_1287_),
    .D(_1285_));
 sg13g2_nor2_1 _3637_ (.A(_1892_),
    .B(_1894_),
    .Y(_1288_));
 sg13g2_a221oi_1 _3638_ (.B2(_1283_),
    .C1(net589),
    .B1(_1288_),
    .A1(_1892_),
    .Y(_0126_),
    .A2(_1286_));
 sg13g2_nand3_1 _3639_ (.B(\pwm_module.counter0[18] ),
    .C(_1285_),
    .A(\pwm_module.counter0[19] ),
    .Y(_1289_));
 sg13g2_nor2_1 _3640_ (.A(_1280_),
    .B(_1289_),
    .Y(_1290_));
 sg13g2_nand2_1 _3641_ (.Y(_1291_),
    .A(net593),
    .B(_1290_));
 sg13g2_a221oi_1 _3642_ (.B2(net593),
    .C1(net588),
    .B1(_1290_),
    .A1(_1890_),
    .Y(_0127_),
    .A2(_1287_));
 sg13g2_nor3_1 _3643_ (.A(_1888_),
    .B(_1280_),
    .C(_1289_),
    .Y(_1292_));
 sg13g2_a221oi_1 _3644_ (.B2(net593),
    .C1(net588),
    .B1(_1292_),
    .A1(_1888_),
    .Y(_0128_),
    .A2(_1291_));
 sg13g2_a21o_1 _3645_ (.A2(_1292_),
    .A1(net593),
    .B1(net548),
    .X(_1293_));
 sg13g2_nand3_1 _3646_ (.B(net593),
    .C(_1292_),
    .A(\pwm_module.counter0[21] ),
    .Y(_1294_));
 sg13g2_and3_1 _3647_ (.X(_0129_),
    .A(_1241_),
    .B(_1293_),
    .C(_1294_));
 sg13g2_nand3_1 _3648_ (.B(\pwm_module.counter0[21] ),
    .C(\pwm_module.counter0[20] ),
    .A(\pwm_module.counter0[22] ),
    .Y(_1295_));
 sg13g2_nor2_1 _3649_ (.A(_1289_),
    .B(_1295_),
    .Y(_1296_));
 sg13g2_and2_1 _3650_ (.A(_1279_),
    .B(_1296_),
    .X(_1297_));
 sg13g2_a21o_1 _3651_ (.A2(_1297_),
    .A1(net593),
    .B1(net588),
    .X(_1298_));
 sg13g2_a21oi_1 _3652_ (.A1(_1885_),
    .A2(_1294_),
    .Y(_0130_),
    .B1(_1298_));
 sg13g2_a21oi_1 _3653_ (.A1(net594),
    .A2(_1297_),
    .Y(_1299_),
    .B1(net203));
 sg13g2_and4_1 _3654_ (.A(net203),
    .B(net593),
    .C(_1278_),
    .D(_1296_),
    .X(_1300_));
 sg13g2_nor3_1 _3655_ (.A(net588),
    .B(_1299_),
    .C(_1300_),
    .Y(_0131_));
 sg13g2_or3_1 _3656_ (.A(_1883_),
    .B(_1289_),
    .C(_1295_),
    .X(_1301_));
 sg13g2_or2_1 _3657_ (.X(_1302_),
    .B(_1301_),
    .A(_1280_));
 sg13g2_a21oi_2 _3658_ (.B1(_1302_),
    .Y(_1303_),
    .A2(_0616_),
    .A1(net646));
 sg13g2_xnor2_1 _3659_ (.Y(_1304_),
    .A(net371),
    .B(_1303_));
 sg13g2_nor2_1 _3660_ (.A(net589),
    .B(_1304_),
    .Y(_0132_));
 sg13g2_a21o_1 _3661_ (.A2(_1303_),
    .A1(net371),
    .B1(net518),
    .X(_1305_));
 sg13g2_nand3_1 _3662_ (.B(net371),
    .C(_1303_),
    .A(net518),
    .Y(_1306_));
 sg13g2_and3_1 _3663_ (.X(_0133_),
    .A(net568),
    .B(_1305_),
    .C(_1306_));
 sg13g2_nor3_1 _3664_ (.A(_1877_),
    .B(_1879_),
    .C(_1881_),
    .Y(_1307_));
 sg13g2_a221oi_1 _3665_ (.B2(_1300_),
    .C1(net588),
    .B1(_1307_),
    .A1(_1877_),
    .Y(_0134_),
    .A2(_1306_));
 sg13g2_a21o_1 _3666_ (.A2(_1307_),
    .A1(_1303_),
    .B1(net519),
    .X(_1308_));
 sg13g2_and2_1 _3667_ (.A(\pwm_module.counter0[27] ),
    .B(_1307_),
    .X(_1309_));
 sg13g2_inv_1 _3668_ (.Y(_1310_),
    .A(_1309_));
 sg13g2_nand2_1 _3669_ (.Y(_1311_),
    .A(_1303_),
    .B(_1309_));
 sg13g2_and3_1 _3670_ (.X(_0135_),
    .A(net568),
    .B(_1308_),
    .C(_1311_));
 sg13g2_nor4_2 _3671_ (.A(_1874_),
    .B(_1280_),
    .C(_1301_),
    .Y(_1312_),
    .D(_1310_));
 sg13g2_a221oi_1 _3672_ (.B2(net594),
    .C1(net588),
    .B1(_1312_),
    .A1(_1874_),
    .Y(_0136_),
    .A2(_1311_));
 sg13g2_a21o_1 _3673_ (.A2(_1312_),
    .A1(net594),
    .B1(net533),
    .X(_1313_));
 sg13g2_nand3_1 _3674_ (.B(net594),
    .C(_1312_),
    .A(net533),
    .Y(_1314_));
 sg13g2_and3_1 _3675_ (.X(_0137_),
    .A(net568),
    .B(_1313_),
    .C(_1314_));
 sg13g2_and3_1 _3676_ (.X(_1315_),
    .A(net290),
    .B(\pwm_module.counter0[29] ),
    .C(_1312_));
 sg13g2_a221oi_1 _3677_ (.B2(net594),
    .C1(net588),
    .B1(_1315_),
    .A1(_1872_),
    .Y(_0138_),
    .A2(_1314_));
 sg13g2_a21oi_1 _3678_ (.A1(net594),
    .A2(_1315_),
    .Y(_1316_),
    .B1(net56));
 sg13g2_nor2_1 _3679_ (.A(net588),
    .B(net57),
    .Y(_0139_));
 sg13g2_mux2_1 _3680_ (.A0(net679),
    .A1(\spi_module.r_RX_Byte[0] ),
    .S(net643),
    .X(_0140_));
 sg13g2_mux2_1 _3681_ (.A0(net676),
    .A1(\spi_module.r_RX_Byte[1] ),
    .S(net643),
    .X(_0141_));
 sg13g2_mux2_1 _3682_ (.A0(net672),
    .A1(\spi_module.r_RX_Byte[2] ),
    .S(net643),
    .X(_0142_));
 sg13g2_mux2_1 _3683_ (.A0(net669),
    .A1(\spi_module.r_RX_Byte[3] ),
    .S(net643),
    .X(_0143_));
 sg13g2_mux2_1 _3684_ (.A0(net666),
    .A1(\spi_module.r_RX_Byte[4] ),
    .S(net643),
    .X(_0144_));
 sg13g2_mux2_1 _3685_ (.A0(net663),
    .A1(\spi_module.r_RX_Byte[5] ),
    .S(_0099_),
    .X(_0145_));
 sg13g2_mux2_1 _3686_ (.A0(net659),
    .A1(\spi_module.r_RX_Byte[6] ),
    .S(net643),
    .X(_0146_));
 sg13g2_mux2_1 _3687_ (.A0(net656),
    .A1(\spi_module.r_RX_Byte[7] ),
    .S(net643),
    .X(_0147_));
 sg13g2_mux2_1 _3688_ (.A0(net1),
    .A1(\spi_module.r_Temp_RX_Byte[0] ),
    .S(net682),
    .X(_0148_));
 sg13g2_mux2_1 _3689_ (.A0(\spi_module.r_Temp_RX_Byte[0] ),
    .A1(\spi_module.r_Temp_RX_Byte[1] ),
    .S(net682),
    .X(_0149_));
 sg13g2_mux2_1 _3690_ (.A0(\spi_module.r_Temp_RX_Byte[1] ),
    .A1(\spi_module.r_Temp_RX_Byte[2] ),
    .S(net682),
    .X(_0150_));
 sg13g2_mux2_1 _3691_ (.A0(\spi_module.r_Temp_RX_Byte[2] ),
    .A1(\spi_module.r_Temp_RX_Byte[3] ),
    .S(net682),
    .X(_0151_));
 sg13g2_mux2_1 _3692_ (.A0(\spi_module.r_Temp_RX_Byte[3] ),
    .A1(\spi_module.r_Temp_RX_Byte[4] ),
    .S(net682),
    .X(_0152_));
 sg13g2_mux2_1 _3693_ (.A0(\spi_module.r_Temp_RX_Byte[4] ),
    .A1(\spi_module.r_Temp_RX_Byte[5] ),
    .S(net682),
    .X(_0153_));
 sg13g2_mux2_1 _3694_ (.A0(\spi_module.r_Temp_RX_Byte[5] ),
    .A1(\spi_module.r_Temp_RX_Byte[6] ),
    .S(net682),
    .X(_0154_));
 sg13g2_nor2_2 _3695_ (.A(net683),
    .B(_1945_),
    .Y(_1317_));
 sg13g2_mux2_1 _3696_ (.A0(\spi_module.r_RX_Byte[0] ),
    .A1(net1),
    .S(_1317_),
    .X(_0155_));
 sg13g2_mux2_1 _3697_ (.A0(\spi_module.r_RX_Byte[1] ),
    .A1(\spi_module.r_Temp_RX_Byte[0] ),
    .S(_1317_),
    .X(_0156_));
 sg13g2_mux2_1 _3698_ (.A0(\spi_module.r_RX_Byte[2] ),
    .A1(\spi_module.r_Temp_RX_Byte[1] ),
    .S(_1317_),
    .X(_0157_));
 sg13g2_mux2_1 _3699_ (.A0(\spi_module.r_RX_Byte[3] ),
    .A1(\spi_module.r_Temp_RX_Byte[2] ),
    .S(_1317_),
    .X(_0158_));
 sg13g2_mux2_1 _3700_ (.A0(\spi_module.r_RX_Byte[4] ),
    .A1(\spi_module.r_Temp_RX_Byte[3] ),
    .S(_1317_),
    .X(_0159_));
 sg13g2_mux2_1 _3701_ (.A0(\spi_module.r_RX_Byte[5] ),
    .A1(\spi_module.r_Temp_RX_Byte[4] ),
    .S(_1317_),
    .X(_0160_));
 sg13g2_mux2_1 _3702_ (.A0(\spi_module.r_RX_Byte[6] ),
    .A1(\spi_module.r_Temp_RX_Byte[5] ),
    .S(_1317_),
    .X(_0161_));
 sg13g2_mux2_1 _3703_ (.A0(\spi_module.r_RX_Byte[7] ),
    .A1(\spi_module.r_Temp_RX_Byte[6] ),
    .S(_1317_),
    .X(_0162_));
 sg13g2_nor3_1 _3704_ (.A(\MemCell.curr_state[2] ),
    .B(\MemCell.curr_state[0] ),
    .C(\MemCell.curr_state[1] ),
    .Y(_1318_));
 sg13g2_a21o_1 _3705_ (.A2(\MemCell.curr_state[1] ),
    .A1(\MemCell.curr_state[2] ),
    .B1(_1318_),
    .X(_1319_));
 sg13g2_nand3b_1 _3706_ (.B(_1039_),
    .C(\MemCell.o_RX_DV ),
    .Y(_1320_),
    .A_N(_1319_));
 sg13g2_nor2_2 _3707_ (.A(_1036_),
    .B(_1320_),
    .Y(_1321_));
 sg13g2_mux2_1 _3708_ (.A0(net149),
    .A1(net679),
    .S(net634),
    .X(_0164_));
 sg13g2_mux2_1 _3709_ (.A0(net49),
    .A1(net676),
    .S(net634),
    .X(_0165_));
 sg13g2_nand2_1 _3710_ (.Y(_1322_),
    .A(net672),
    .B(net634));
 sg13g2_o21ai_1 _3711_ (.B1(_1322_),
    .Y(_0166_),
    .A1(_1941_),
    .A2(net634));
 sg13g2_mux2_1 _3712_ (.A0(net92),
    .A1(net668),
    .S(net634),
    .X(_0167_));
 sg13g2_nand2_1 _3713_ (.Y(_1323_),
    .A(net665),
    .B(_1321_));
 sg13g2_o21ai_1 _3714_ (.B1(_1323_),
    .Y(_0168_),
    .A1(_1940_),
    .A2(net634));
 sg13g2_nand2_1 _3715_ (.Y(_1324_),
    .A(net662),
    .B(net634));
 sg13g2_o21ai_1 _3716_ (.B1(_1324_),
    .Y(_0169_),
    .A1(_1939_),
    .A2(net634));
 sg13g2_mux2_1 _3717_ (.A0(net168),
    .A1(net659),
    .S(_1321_),
    .X(_0170_));
 sg13g2_mux2_1 _3718_ (.A0(net120),
    .A1(net656),
    .S(_1321_),
    .X(_0171_));
 sg13g2_nand2b_2 _3719_ (.Y(_1325_),
    .B(\MemCell.counter[1] ),
    .A_N(net650));
 sg13g2_nand2_2 _3720_ (.Y(_1326_),
    .A(\MemCell.o_RX_DV ),
    .B(_1030_));
 sg13g2_nor2_2 _3721_ (.A(_1325_),
    .B(_1326_),
    .Y(_1327_));
 sg13g2_mux2_1 _3722_ (.A0(net58),
    .A1(net679),
    .S(net633),
    .X(_0172_));
 sg13g2_mux2_1 _3723_ (.A0(net93),
    .A1(net676),
    .S(net633),
    .X(_0173_));
 sg13g2_mux2_1 _3724_ (.A0(net173),
    .A1(net672),
    .S(net633),
    .X(_0174_));
 sg13g2_mux2_1 _3725_ (.A0(net66),
    .A1(net668),
    .S(_1327_),
    .X(_0175_));
 sg13g2_nand2_1 _3726_ (.Y(_1328_),
    .A(net665),
    .B(_1327_));
 sg13g2_o21ai_1 _3727_ (.B1(_1328_),
    .Y(_0176_),
    .A1(_1819_),
    .A2(net633));
 sg13g2_nand2_1 _3728_ (.Y(_1329_),
    .A(net662),
    .B(net633));
 sg13g2_o21ai_1 _3729_ (.B1(_1329_),
    .Y(_0177_),
    .A1(_1818_),
    .A2(net633));
 sg13g2_mux2_1 _3730_ (.A0(net71),
    .A1(net659),
    .S(net633),
    .X(_0178_));
 sg13g2_mux2_1 _3731_ (.A0(net193),
    .A1(net656),
    .S(net633),
    .X(_0179_));
 sg13g2_nor2_2 _3732_ (.A(_1320_),
    .B(_1325_),
    .Y(_1330_));
 sg13g2_mux2_1 _3733_ (.A0(net95),
    .A1(net679),
    .S(net632),
    .X(_0180_));
 sg13g2_mux2_1 _3734_ (.A0(net59),
    .A1(net676),
    .S(net632),
    .X(_0181_));
 sg13g2_mux2_1 _3735_ (.A0(net65),
    .A1(net672),
    .S(net632),
    .X(_0182_));
 sg13g2_mux2_1 _3736_ (.A0(net105),
    .A1(net668),
    .S(net632),
    .X(_0183_));
 sg13g2_nand2_1 _3737_ (.Y(_1331_),
    .A(net665),
    .B(net632));
 sg13g2_o21ai_1 _3738_ (.B1(_1331_),
    .Y(_0184_),
    .A1(_1943_),
    .A2(net632));
 sg13g2_nand2_1 _3739_ (.Y(_1332_),
    .A(net662),
    .B(net632));
 sg13g2_o21ai_1 _3740_ (.B1(_1332_),
    .Y(_0185_),
    .A1(_1942_),
    .A2(net632));
 sg13g2_mux2_1 _3741_ (.A0(net137),
    .A1(net659),
    .S(_1330_),
    .X(_0186_));
 sg13g2_mux2_1 _3742_ (.A0(net239),
    .A1(net654),
    .S(_1330_),
    .X(_0187_));
 sg13g2_nand2b_2 _3743_ (.Y(_1333_),
    .B(net650),
    .A_N(\MemCell.counter[1] ));
 sg13g2_nor2_1 _3744_ (.A(_1320_),
    .B(_1333_),
    .Y(_1334_));
 sg13g2_nand2_1 _3745_ (.Y(_1335_),
    .A(net678),
    .B(net630));
 sg13g2_o21ai_1 _3746_ (.B1(_1335_),
    .Y(_0188_),
    .A1(_1796_),
    .A2(net630));
 sg13g2_nand2_1 _3747_ (.Y(_1336_),
    .A(net674),
    .B(net630));
 sg13g2_o21ai_1 _3748_ (.B1(_1336_),
    .Y(_0189_),
    .A1(_1794_),
    .A2(net630));
 sg13g2_mux2_1 _3749_ (.A0(net73),
    .A1(net670),
    .S(net630),
    .X(_0190_));
 sg13g2_mux2_1 _3750_ (.A0(net127),
    .A1(net667),
    .S(net631),
    .X(_0191_));
 sg13g2_nand2_1 _3751_ (.Y(_1337_),
    .A(net664),
    .B(net630));
 sg13g2_o21ai_1 _3752_ (.B1(_1337_),
    .Y(_0192_),
    .A1(_1790_),
    .A2(net631));
 sg13g2_nand2_1 _3753_ (.Y(_1338_),
    .A(net661),
    .B(net630));
 sg13g2_o21ai_1 _3754_ (.B1(_1338_),
    .Y(_0193_),
    .A1(_1789_),
    .A2(net631));
 sg13g2_nand2_1 _3755_ (.Y(_1339_),
    .A(net658),
    .B(net630));
 sg13g2_o21ai_1 _3756_ (.B1(_1339_),
    .Y(_0194_),
    .A1(_1787_),
    .A2(net631));
 sg13g2_mux2_1 _3757_ (.A0(net128),
    .A1(net654),
    .S(net631),
    .X(_0195_));
 sg13g2_nor2_2 _3758_ (.A(net650),
    .B(\MemCell.counter[1] ),
    .Y(_1340_));
 sg13g2_nand2b_2 _3759_ (.Y(_1341_),
    .B(_1340_),
    .A_N(_1320_));
 sg13g2_mux2_1 _3760_ (.A0(net678),
    .A1(net76),
    .S(net629),
    .X(_0196_));
 sg13g2_mux2_1 _3761_ (.A0(net674),
    .A1(net234),
    .S(net629),
    .X(_0197_));
 sg13g2_mux2_1 _3762_ (.A0(net670),
    .A1(net218),
    .S(net629),
    .X(_0198_));
 sg13g2_mux2_1 _3763_ (.A0(net667),
    .A1(net170),
    .S(net629),
    .X(_0199_));
 sg13g2_nor2_1 _3764_ (.A(net664),
    .B(net629),
    .Y(_1342_));
 sg13g2_a21oi_1 _3765_ (.A1(_1802_),
    .A2(net629),
    .Y(_0200_),
    .B1(_1342_));
 sg13g2_nor2_1 _3766_ (.A(net661),
    .B(net629),
    .Y(_1343_));
 sg13g2_a21oi_1 _3767_ (.A1(_1800_),
    .A2(_1341_),
    .Y(_0201_),
    .B1(_1343_));
 sg13g2_mux2_1 _3768_ (.A0(net658),
    .A1(net211),
    .S(_1341_),
    .X(_0202_));
 sg13g2_mux2_1 _3769_ (.A0(net654),
    .A1(net181),
    .S(net629),
    .X(_0203_));
 sg13g2_nand2_2 _3770_ (.Y(_1344_),
    .A(\MemCell.o_RX_DV ),
    .B(_1032_));
 sg13g2_nor2_2 _3771_ (.A(_1036_),
    .B(_1344_),
    .Y(_1345_));
 sg13g2_mux2_1 _3772_ (.A0(net268),
    .A1(net680),
    .S(net628),
    .X(_0204_));
 sg13g2_mux2_1 _3773_ (.A0(net230),
    .A1(net676),
    .S(net627),
    .X(_0205_));
 sg13g2_nand2_1 _3774_ (.Y(_1346_),
    .A(net672),
    .B(net627));
 sg13g2_o21ai_1 _3775_ (.B1(_1346_),
    .Y(_0206_),
    .A1(_1929_),
    .A2(net628));
 sg13g2_nand2_1 _3776_ (.Y(_1347_),
    .A(net668),
    .B(net628));
 sg13g2_o21ai_1 _3777_ (.B1(_1347_),
    .Y(_0207_),
    .A1(_1928_),
    .A2(net628));
 sg13g2_mux2_1 _3778_ (.A0(net69),
    .A1(net665),
    .S(net627),
    .X(_0208_));
 sg13g2_mux2_1 _3779_ (.A0(net94),
    .A1(net662),
    .S(net627),
    .X(_0209_));
 sg13g2_nand2_1 _3780_ (.Y(_1348_),
    .A(net659),
    .B(net627));
 sg13g2_o21ai_1 _3781_ (.B1(_1348_),
    .Y(_0210_),
    .A1(_1927_),
    .A2(net627));
 sg13g2_nand2_1 _3782_ (.Y(_1349_),
    .A(net656),
    .B(net627));
 sg13g2_o21ai_1 _3783_ (.B1(_1349_),
    .Y(_0211_),
    .A1(_1926_),
    .A2(net627));
 sg13g2_nor2_1 _3784_ (.A(_1325_),
    .B(_1344_),
    .Y(_1350_));
 sg13g2_mux2_1 _3785_ (.A0(net54),
    .A1(net680),
    .S(net626),
    .X(_0212_));
 sg13g2_mux2_1 _3786_ (.A0(net158),
    .A1(net677),
    .S(net626),
    .X(_0213_));
 sg13g2_mux2_1 _3787_ (.A0(net90),
    .A1(net673),
    .S(net626),
    .X(_0214_));
 sg13g2_mux2_1 _3788_ (.A0(net60),
    .A1(net669),
    .S(net626),
    .X(_0215_));
 sg13g2_mux2_1 _3789_ (.A0(net84),
    .A1(net665),
    .S(net626),
    .X(_0216_));
 sg13g2_mux2_1 _3790_ (.A0(net50),
    .A1(net662),
    .S(net626),
    .X(_0217_));
 sg13g2_nand2_1 _3791_ (.Y(_1351_),
    .A(net660),
    .B(_1350_));
 sg13g2_o21ai_1 _3792_ (.B1(_1351_),
    .Y(_0218_),
    .A1(_1931_),
    .A2(net626));
 sg13g2_mux2_1 _3793_ (.A0(net64),
    .A1(net656),
    .S(net626),
    .X(_0219_));
 sg13g2_nor2_1 _3794_ (.A(_1333_),
    .B(_1344_),
    .Y(_1352_));
 sg13g2_nand2_1 _3795_ (.Y(_1353_),
    .A(net678),
    .B(net624));
 sg13g2_o21ai_1 _3796_ (.B1(_1353_),
    .Y(_0220_),
    .A1(_1936_),
    .A2(net624));
 sg13g2_nand2_1 _3797_ (.Y(_1354_),
    .A(net675),
    .B(net624));
 sg13g2_o21ai_1 _3798_ (.B1(_1354_),
    .Y(_0221_),
    .A1(_1935_),
    .A2(net624));
 sg13g2_nand2_1 _3799_ (.Y(_1355_),
    .A(net671),
    .B(net624));
 sg13g2_o21ai_1 _3800_ (.B1(_1355_),
    .Y(_0222_),
    .A1(_1934_),
    .A2(net624));
 sg13g2_nand2_1 _3801_ (.Y(_1356_),
    .A(net667),
    .B(net624));
 sg13g2_o21ai_1 _3802_ (.B1(_1356_),
    .Y(_0223_),
    .A1(_1933_),
    .A2(net624));
 sg13g2_mux2_1 _3803_ (.A0(net86),
    .A1(net666),
    .S(net625),
    .X(_0224_));
 sg13g2_mux2_1 _3804_ (.A0(net106),
    .A1(net663),
    .S(net625),
    .X(_0225_));
 sg13g2_nand2_1 _3805_ (.Y(_1357_),
    .A(net660),
    .B(net625));
 sg13g2_o21ai_1 _3806_ (.B1(_1357_),
    .Y(_0226_),
    .A1(_1932_),
    .A2(net625));
 sg13g2_mux2_1 _3807_ (.A0(net139),
    .A1(net655),
    .S(net625),
    .X(_0227_));
 sg13g2_nor3_2 _3808_ (.A(net650),
    .B(\MemCell.counter[1] ),
    .C(_1344_),
    .Y(_1358_));
 sg13g2_mux2_1 _3809_ (.A0(net43),
    .A1(net680),
    .S(net623),
    .X(_0228_));
 sg13g2_mux2_1 _3810_ (.A0(net100),
    .A1(net675),
    .S(net623),
    .X(_0229_));
 sg13g2_mux2_1 _3811_ (.A0(net83),
    .A1(net671),
    .S(net623),
    .X(_0230_));
 sg13g2_mux2_1 _3812_ (.A0(net62),
    .A1(net669),
    .S(net623),
    .X(_0231_));
 sg13g2_nand2_1 _3813_ (.Y(_1359_),
    .A(net666),
    .B(net623));
 sg13g2_o21ai_1 _3814_ (.B1(_1359_),
    .Y(_0232_),
    .A1(_1938_),
    .A2(net623));
 sg13g2_nand2_1 _3815_ (.Y(_1360_),
    .A(net663),
    .B(_1358_));
 sg13g2_o21ai_1 _3816_ (.B1(_1360_),
    .Y(_0233_),
    .A1(_1937_),
    .A2(_1358_));
 sg13g2_mux2_1 _3817_ (.A0(net77),
    .A1(net660),
    .S(net623),
    .X(_0234_));
 sg13g2_mux2_1 _3818_ (.A0(net70),
    .A1(net655),
    .S(net623),
    .X(_0235_));
 sg13g2_nor3_2 _3819_ (.A(_1846_),
    .B(_1042_),
    .C(_1319_),
    .Y(_1361_));
 sg13g2_nand2_2 _3820_ (.Y(_1362_),
    .A(_1035_),
    .B(_1361_));
 sg13g2_mux2_1 _3821_ (.A0(net679),
    .A1(net517),
    .S(net617),
    .X(_0236_));
 sg13g2_nor2_1 _3822_ (.A(net677),
    .B(net617),
    .Y(_1363_));
 sg13g2_a21oi_1 _3823_ (.A1(_1858_),
    .A2(net616),
    .Y(_0237_),
    .B1(_1363_));
 sg13g2_mux2_1 _3824_ (.A0(net673),
    .A1(net492),
    .S(net616),
    .X(_0238_));
 sg13g2_nor2_1 _3825_ (.A(net668),
    .B(net616),
    .Y(_1364_));
 sg13g2_a21oi_1 _3826_ (.A1(_1857_),
    .A2(net616),
    .Y(_0239_),
    .B1(_1364_));
 sg13g2_nor2_1 _3827_ (.A(net666),
    .B(net616),
    .Y(_1365_));
 sg13g2_a21oi_1 _3828_ (.A1(_1856_),
    .A2(net616),
    .Y(_0240_),
    .B1(_1365_));
 sg13g2_mux2_1 _3829_ (.A0(net663),
    .A1(net512),
    .S(net617),
    .X(_0241_));
 sg13g2_nor2_1 _3830_ (.A(net660),
    .B(net616),
    .Y(_1366_));
 sg13g2_a21oi_1 _3831_ (.A1(_1855_),
    .A2(net616),
    .Y(_0242_),
    .B1(_1366_));
 sg13g2_mux2_1 _3832_ (.A0(net657),
    .A1(net487),
    .S(net617),
    .X(_0243_));
 sg13g2_nand2b_2 _3833_ (.Y(_1367_),
    .B(_1361_),
    .A_N(_1325_));
 sg13g2_mux2_1 _3834_ (.A0(net680),
    .A1(\MemCell.prescale_reg[2][0] ),
    .S(_1367_),
    .X(_0244_));
 sg13g2_mux2_1 _3835_ (.A0(net677),
    .A1(net479),
    .S(_1367_),
    .X(_0245_));
 sg13g2_mux2_1 _3836_ (.A0(net673),
    .A1(\MemCell.prescale_reg[2][2] ),
    .S(net615),
    .X(_0246_));
 sg13g2_mux2_1 _3837_ (.A0(net669),
    .A1(net112),
    .S(net615),
    .X(_0247_));
 sg13g2_nor2_1 _3838_ (.A(net666),
    .B(net615),
    .Y(_1368_));
 sg13g2_a21oi_1 _3839_ (.A1(_1862_),
    .A2(net615),
    .Y(_0248_),
    .B1(_1368_));
 sg13g2_nor2_1 _3840_ (.A(net663),
    .B(net615),
    .Y(_1369_));
 sg13g2_a21oi_1 _3841_ (.A1(_1860_),
    .A2(net615),
    .Y(_0249_),
    .B1(_1369_));
 sg13g2_mux2_1 _3842_ (.A0(net660),
    .A1(net520),
    .S(net615),
    .X(_0250_));
 sg13g2_mux2_1 _3843_ (.A0(net657),
    .A1(\MemCell.prescale_reg[2][7] ),
    .S(net615),
    .X(_0251_));
 sg13g2_nor2_1 _3844_ (.A(_1326_),
    .B(_1333_),
    .Y(_1370_));
 sg13g2_nand2_1 _3845_ (.Y(_1371_),
    .A(net678),
    .B(net621));
 sg13g2_o21ai_1 _3846_ (.B1(_1371_),
    .Y(_0252_),
    .A1(_1833_),
    .A2(net621));
 sg13g2_nand2_1 _3847_ (.Y(_1372_),
    .A(net674),
    .B(net621));
 sg13g2_o21ai_1 _3848_ (.B1(_1372_),
    .Y(_0253_),
    .A1(_1831_),
    .A2(net621));
 sg13g2_mux2_1 _3849_ (.A0(net82),
    .A1(net670),
    .S(net621),
    .X(_0254_));
 sg13g2_mux2_1 _3850_ (.A0(net126),
    .A1(net667),
    .S(net621),
    .X(_0255_));
 sg13g2_nand2_1 _3851_ (.Y(_1373_),
    .A(net664),
    .B(net622));
 sg13g2_o21ai_1 _3852_ (.B1(_1373_),
    .Y(_0256_),
    .A1(_1828_),
    .A2(net622));
 sg13g2_nand2_1 _3853_ (.Y(_1374_),
    .A(net661),
    .B(net622));
 sg13g2_o21ai_1 _3854_ (.B1(_1374_),
    .Y(_0257_),
    .A1(_1826_),
    .A2(net622));
 sg13g2_nand2_1 _3855_ (.Y(_1375_),
    .A(net658),
    .B(net622));
 sg13g2_o21ai_1 _3856_ (.B1(_1375_),
    .Y(_0258_),
    .A1(_1824_),
    .A2(net621));
 sg13g2_mux2_1 _3857_ (.A0(net97),
    .A1(net654),
    .S(net621),
    .X(_0259_));
 sg13g2_nand2b_1 _3858_ (.Y(_1376_),
    .B(_1361_),
    .A_N(_1333_));
 sg13g2_nor2_1 _3859_ (.A(net680),
    .B(net614),
    .Y(_1377_));
 sg13g2_a21oi_1 _3860_ (.A1(_1854_),
    .A2(net614),
    .Y(_0260_),
    .B1(_1377_));
 sg13g2_mux2_1 _3861_ (.A0(net675),
    .A1(net406),
    .S(net614),
    .X(_0261_));
 sg13g2_mux2_1 _3862_ (.A0(net670),
    .A1(net467),
    .S(net614),
    .X(_0262_));
 sg13g2_mux2_1 _3863_ (.A0(net667),
    .A1(net74),
    .S(net614),
    .X(_0263_));
 sg13g2_mux2_1 _3864_ (.A0(net664),
    .A1(net489),
    .S(_1376_),
    .X(_0264_));
 sg13g2_mux2_1 _3865_ (.A0(net661),
    .A1(net494),
    .S(net614),
    .X(_0265_));
 sg13g2_mux2_1 _3866_ (.A0(net658),
    .A1(net468),
    .S(net614),
    .X(_0266_));
 sg13g2_mux2_1 _3867_ (.A0(net654),
    .A1(net495),
    .S(net614),
    .X(_0267_));
 sg13g2_nand2_2 _3868_ (.Y(_1378_),
    .A(_1340_),
    .B(_1361_));
 sg13g2_mux2_1 _3869_ (.A0(net678),
    .A1(net260),
    .S(net613),
    .X(_0268_));
 sg13g2_mux2_1 _3870_ (.A0(net674),
    .A1(net431),
    .S(net613),
    .X(_0269_));
 sg13g2_nor2_1 _3871_ (.A(net670),
    .B(net613),
    .Y(_1379_));
 sg13g2_a21oi_1 _3872_ (.A1(_1849_),
    .A2(net613),
    .Y(_0270_),
    .B1(_1379_));
 sg13g2_nor2_1 _3873_ (.A(net669),
    .B(net613),
    .Y(_1380_));
 sg13g2_a21oi_1 _3874_ (.A1(_1847_),
    .A2(net613),
    .Y(_0271_),
    .B1(_1380_));
 sg13g2_mux2_1 _3875_ (.A0(net664),
    .A1(net350),
    .S(net613),
    .X(_0272_));
 sg13g2_mux2_1 _3876_ (.A0(net663),
    .A1(net438),
    .S(net613),
    .X(_0273_));
 sg13g2_mux2_1 _3877_ (.A0(net658),
    .A1(net496),
    .S(_1378_),
    .X(_0274_));
 sg13g2_mux2_1 _3878_ (.A0(net655),
    .A1(net456),
    .S(_1378_),
    .X(_0275_));
 sg13g2_nand4_1 _3879_ (.B(_1845_),
    .C(_0102_),
    .A(\MemCell.curr_state[0] ),
    .Y(_1381_),
    .D(\MemCell.o_RX_DV ));
 sg13g2_nor2_2 _3880_ (.A(_1036_),
    .B(_1381_),
    .Y(_1382_));
 sg13g2_nand2_1 _3881_ (.Y(_1383_),
    .A(net679),
    .B(net641));
 sg13g2_o21ai_1 _3882_ (.B1(_1383_),
    .Y(_0276_),
    .A1(_1882_),
    .A2(net641));
 sg13g2_nand2_1 _3883_ (.Y(_1384_),
    .A(net676),
    .B(net641));
 sg13g2_o21ai_1 _3884_ (.B1(_1384_),
    .Y(_0277_),
    .A1(_1880_),
    .A2(net641));
 sg13g2_nand2_1 _3885_ (.Y(_1385_),
    .A(net672),
    .B(net641));
 sg13g2_o21ai_1 _3886_ (.B1(_1385_),
    .Y(_0278_),
    .A1(_1878_),
    .A2(net641));
 sg13g2_nand2_1 _3887_ (.Y(_1386_),
    .A(net668),
    .B(net641));
 sg13g2_o21ai_1 _3888_ (.B1(_1386_),
    .Y(_0279_),
    .A1(_1876_),
    .A2(net641));
 sg13g2_nand2_1 _3889_ (.Y(_1387_),
    .A(net665),
    .B(net642));
 sg13g2_o21ai_1 _3890_ (.B1(_1387_),
    .Y(_0280_),
    .A1(_1875_),
    .A2(net642));
 sg13g2_nand2_1 _3891_ (.Y(_1388_),
    .A(net662),
    .B(net642));
 sg13g2_o21ai_1 _3892_ (.B1(_1388_),
    .Y(_0281_),
    .A1(_1873_),
    .A2(net642));
 sg13g2_mux2_1 _3893_ (.A0(net449),
    .A1(net659),
    .S(net642),
    .X(_0282_));
 sg13g2_mux2_1 _3894_ (.A0(net368),
    .A1(net656),
    .S(net642),
    .X(_0283_));
 sg13g2_nor2_1 _3895_ (.A(_1325_),
    .B(_1381_),
    .Y(_1389_));
 sg13g2_nand2_1 _3896_ (.Y(_1390_),
    .A(net679),
    .B(net639));
 sg13g2_o21ai_1 _3897_ (.B1(_1390_),
    .Y(_0284_),
    .A1(_1897_),
    .A2(net639));
 sg13g2_nand2_1 _3898_ (.Y(_1391_),
    .A(net676),
    .B(net639));
 sg13g2_o21ai_1 _3899_ (.B1(_1391_),
    .Y(_0285_),
    .A1(_1895_),
    .A2(net639));
 sg13g2_nand2_1 _3900_ (.Y(_1392_),
    .A(net672),
    .B(net639));
 sg13g2_o21ai_1 _3901_ (.B1(_1392_),
    .Y(_0286_),
    .A1(_1893_),
    .A2(net639));
 sg13g2_nand2_1 _3902_ (.Y(_1393_),
    .A(net668),
    .B(net639));
 sg13g2_o21ai_1 _3903_ (.B1(_1393_),
    .Y(_0287_),
    .A1(_1891_),
    .A2(net639));
 sg13g2_nand2_1 _3904_ (.Y(_1394_),
    .A(net665),
    .B(net640));
 sg13g2_o21ai_1 _3905_ (.B1(_1394_),
    .Y(_0288_),
    .A1(_1889_),
    .A2(net640));
 sg13g2_nand2_1 _3906_ (.Y(_1395_),
    .A(net662),
    .B(net640));
 sg13g2_o21ai_1 _3907_ (.B1(_1395_),
    .Y(_0289_),
    .A1(_1887_),
    .A2(net640));
 sg13g2_nand2_1 _3908_ (.Y(_1396_),
    .A(net659),
    .B(net640));
 sg13g2_o21ai_1 _3909_ (.B1(_1396_),
    .Y(_0290_),
    .A1(_1886_),
    .A2(net640));
 sg13g2_nand2_1 _3910_ (.Y(_1397_),
    .A(net656),
    .B(net640));
 sg13g2_o21ai_1 _3911_ (.B1(_1397_),
    .Y(_0291_),
    .A1(_1884_),
    .A2(net640));
 sg13g2_nor2_1 _3912_ (.A(_1333_),
    .B(_1381_),
    .Y(_1398_));
 sg13g2_nand2_1 _3913_ (.Y(_1399_),
    .A(net678),
    .B(net637));
 sg13g2_o21ai_1 _3914_ (.B1(_1399_),
    .Y(_0292_),
    .A1(_1908_),
    .A2(net637));
 sg13g2_nand2_1 _3915_ (.Y(_1400_),
    .A(net674),
    .B(net637));
 sg13g2_o21ai_1 _3916_ (.B1(_1400_),
    .Y(_0293_),
    .A1(_1906_),
    .A2(net637));
 sg13g2_nand2_1 _3917_ (.Y(_1401_),
    .A(net670),
    .B(net637));
 sg13g2_o21ai_1 _3918_ (.B1(_1401_),
    .Y(_0294_),
    .A1(_1904_),
    .A2(net637));
 sg13g2_mux2_1 _3919_ (.A0(net407),
    .A1(net667),
    .S(net637),
    .X(_0295_));
 sg13g2_nand2_1 _3920_ (.Y(_1402_),
    .A(net664),
    .B(net638));
 sg13g2_o21ai_1 _3921_ (.B1(_1402_),
    .Y(_0296_),
    .A1(_1903_),
    .A2(net638));
 sg13g2_mux2_1 _3922_ (.A0(net352),
    .A1(net661),
    .S(net638),
    .X(_0297_));
 sg13g2_nand2_1 _3923_ (.Y(_1403_),
    .A(net658),
    .B(net638));
 sg13g2_o21ai_1 _3924_ (.B1(_1403_),
    .Y(_0298_),
    .A1(_1900_),
    .A2(net638));
 sg13g2_mux2_1 _3925_ (.A0(net412),
    .A1(net654),
    .S(net637),
    .X(_0299_));
 sg13g2_nor3_2 _3926_ (.A(net650),
    .B(\MemCell.counter[1] ),
    .C(_1381_),
    .Y(_1404_));
 sg13g2_mux2_1 _3927_ (.A0(net222),
    .A1(net678),
    .S(net635),
    .X(_0300_));
 sg13g2_mux2_1 _3928_ (.A0(net339),
    .A1(net674),
    .S(net635),
    .X(_0301_));
 sg13g2_mux2_1 _3929_ (.A0(net435),
    .A1(net670),
    .S(net635),
    .X(_0302_));
 sg13g2_mux2_1 _3930_ (.A0(net358),
    .A1(net667),
    .S(net635),
    .X(_0303_));
 sg13g2_nand2_1 _3931_ (.Y(_1405_),
    .A(net664),
    .B(net635));
 sg13g2_o21ai_1 _3932_ (.B1(_1405_),
    .Y(_0304_),
    .A1(_1914_),
    .A2(net635));
 sg13g2_nand2_1 _3933_ (.Y(_1406_),
    .A(net661),
    .B(net636));
 sg13g2_o21ai_1 _3934_ (.B1(_1406_),
    .Y(_0305_),
    .A1(_1912_),
    .A2(net636));
 sg13g2_nand2_1 _3935_ (.Y(_1407_),
    .A(net658),
    .B(net636));
 sg13g2_o21ai_1 _3936_ (.B1(_1407_),
    .Y(_0306_),
    .A1(_1911_),
    .A2(net636));
 sg13g2_nand2_1 _3937_ (.Y(_1408_),
    .A(net654),
    .B(net635));
 sg13g2_o21ai_1 _3938_ (.B1(_1408_),
    .Y(_0307_),
    .A1(_1910_),
    .A2(net635));
 sg13g2_a22oi_1 _3939_ (.Y(_1409_),
    .B1(_1043_),
    .B2(net651),
    .A2(_1041_),
    .A1(net474));
 sg13g2_inv_1 _3940_ (.Y(_0308_),
    .A(net475));
 sg13g2_nand2b_1 _3941_ (.Y(_1410_),
    .B(_1041_),
    .A_N(\MemCell.curr_state[2] ));
 sg13g2_a21oi_1 _3942_ (.A1(_1040_),
    .A2(_1410_),
    .Y(_1411_),
    .B1(\MemCell.o_RX_DV ));
 sg13g2_or2_1 _3943_ (.X(_1412_),
    .B(_1411_),
    .A(_1319_));
 sg13g2_nand2_1 _3944_ (.Y(_1413_),
    .A(net46),
    .B(_1411_));
 sg13g2_o21ai_1 _3945_ (.B1(_1413_),
    .Y(_0309_),
    .A1(net650),
    .A2(_1412_));
 sg13g2_nor3_1 _3946_ (.A(_1035_),
    .B(_1340_),
    .C(_1412_),
    .Y(_1414_));
 sg13g2_a21o_1 _3947_ (.A2(_1411_),
    .A1(net527),
    .B1(_1414_),
    .X(_0310_));
 sg13g2_nor2b_2 _3948_ (.A(_1326_),
    .B_N(_1340_),
    .Y(_1415_));
 sg13g2_mux2_1 _3949_ (.A0(net45),
    .A1(net678),
    .S(net620),
    .X(_0311_));
 sg13g2_mux2_1 _3950_ (.A0(net99),
    .A1(net674),
    .S(net620),
    .X(_0312_));
 sg13g2_mux2_1 _3951_ (.A0(net68),
    .A1(net670),
    .S(net620),
    .X(_0313_));
 sg13g2_mux2_1 _3952_ (.A0(net72),
    .A1(net667),
    .S(net620),
    .X(_0314_));
 sg13g2_nand2_1 _3953_ (.Y(_1416_),
    .A(net664),
    .B(net620));
 sg13g2_o21ai_1 _3954_ (.B1(_1416_),
    .Y(_0315_),
    .A1(_1840_),
    .A2(net620));
 sg13g2_nand2_1 _3955_ (.Y(_1417_),
    .A(net661),
    .B(_1415_));
 sg13g2_o21ai_1 _3956_ (.B1(_1417_),
    .Y(_0316_),
    .A1(_1837_),
    .A2(net620));
 sg13g2_mux2_1 _3957_ (.A0(net150),
    .A1(net658),
    .S(_1415_),
    .X(_0317_));
 sg13g2_mux2_1 _3958_ (.A0(net75),
    .A1(net654),
    .S(net620),
    .X(_0318_));
 sg13g2_and2_2 _3959_ (.A(_1863_),
    .B(_0963_),
    .X(_1418_));
 sg13g2_nand2_1 _3960_ (.Y(_1419_),
    .A(net644),
    .B(net612));
 sg13g2_nand2b_1 _3961_ (.Y(_1420_),
    .B(\pwm_module.counter2[13] ),
    .A_N(\MemCell.counter_value[13] ));
 sg13g2_o21ai_1 _3962_ (.B1(_1420_),
    .Y(_1421_),
    .A1(_1829_),
    .A2(\MemCell.counter_value[12] ));
 sg13g2_nand2b_1 _3963_ (.Y(_1422_),
    .B(\MemCell.counter_value[15] ),
    .A_N(\pwm_module.counter2[15] ));
 sg13g2_nor2_1 _3964_ (.A(\pwm_module.counter2[12] ),
    .B(_1903_),
    .Y(_1423_));
 sg13g2_nand2b_1 _3965_ (.Y(_1424_),
    .B(\pwm_module.counter2[14] ),
    .A_N(\MemCell.counter_value[14] ));
 sg13g2_nand2b_1 _3966_ (.Y(_1425_),
    .B(\pwm_module.counter2[15] ),
    .A_N(\MemCell.counter_value[15] ));
 sg13g2_nand2_1 _3967_ (.Y(_1426_),
    .A(_1424_),
    .B(_1425_));
 sg13g2_nand2b_1 _3968_ (.Y(_1427_),
    .B(\MemCell.counter_value[14] ),
    .A_N(\pwm_module.counter2[14] ));
 sg13g2_nor2b_1 _3969_ (.A(\pwm_module.counter2[13] ),
    .B_N(\MemCell.counter_value[13] ),
    .Y(_1428_));
 sg13g2_nand4_1 _3970_ (.B(_1424_),
    .C(_1425_),
    .A(_1422_),
    .Y(_1429_),
    .D(_1427_));
 sg13g2_nor4_2 _3971_ (.A(_1421_),
    .B(_1423_),
    .C(_1428_),
    .Y(_1430_),
    .D(_1429_));
 sg13g2_nand2b_1 _3972_ (.Y(_1431_),
    .B(\pwm_module.counter2[10] ),
    .A_N(\MemCell.counter_value[10] ));
 sg13g2_nand2b_1 _3973_ (.Y(_1432_),
    .B(\pwm_module.counter2[11] ),
    .A_N(\MemCell.counter_value[11] ));
 sg13g2_nor2b_1 _3974_ (.A(\pwm_module.counter2[11] ),
    .B_N(\MemCell.counter_value[11] ),
    .Y(_1433_));
 sg13g2_nand2b_1 _3975_ (.Y(_1434_),
    .B(\MemCell.counter_value[11] ),
    .A_N(\pwm_module.counter2[11] ));
 sg13g2_a21oi_1 _3976_ (.A1(_1431_),
    .A2(_1432_),
    .Y(_1435_),
    .B1(_1433_));
 sg13g2_nand2b_1 _3977_ (.Y(_1436_),
    .B(\pwm_module.counter2[9] ),
    .A_N(\MemCell.counter_value[9] ));
 sg13g2_nand2b_1 _3978_ (.Y(_1437_),
    .B(\pwm_module.counter2[8] ),
    .A_N(\MemCell.counter_value[8] ));
 sg13g2_and2_1 _3979_ (.A(_1436_),
    .B(_1437_),
    .X(_1438_));
 sg13g2_nand2b_1 _3980_ (.Y(_1439_),
    .B(\MemCell.counter_value[10] ),
    .A_N(\pwm_module.counter2[10] ));
 sg13g2_nor2b_1 _3981_ (.A(\pwm_module.counter2[9] ),
    .B_N(\MemCell.counter_value[9] ),
    .Y(_1440_));
 sg13g2_and4_1 _3982_ (.A(_1431_),
    .B(_1432_),
    .C(_1434_),
    .D(_1439_),
    .X(_1441_));
 sg13g2_a21oi_1 _3983_ (.A1(_1436_),
    .A2(_1437_),
    .Y(_1442_),
    .B1(_1440_));
 sg13g2_a21o_1 _3984_ (.A2(_1442_),
    .A1(_1441_),
    .B1(_1435_),
    .X(_1443_));
 sg13g2_nand2b_1 _3985_ (.Y(_1444_),
    .B(\pwm_module.counter2[7] ),
    .A_N(\MemCell.counter_value[7] ));
 sg13g2_nand2b_1 _3986_ (.Y(_1445_),
    .B(\pwm_module.counter2[6] ),
    .A_N(\MemCell.counter_value[6] ));
 sg13g2_and2_1 _3987_ (.A(_1444_),
    .B(_1445_),
    .X(_1446_));
 sg13g2_nor2b_1 _3988_ (.A(\MemCell.counter_value[4] ),
    .B_N(\pwm_module.counter2[4] ),
    .Y(_1447_));
 sg13g2_nor2b_1 _3989_ (.A(\MemCell.counter_value[5] ),
    .B_N(\pwm_module.counter2[5] ),
    .Y(_1448_));
 sg13g2_nor2_1 _3990_ (.A(_1447_),
    .B(_1448_),
    .Y(_1449_));
 sg13g2_nand2b_1 _3991_ (.Y(_1450_),
    .B(net649),
    .A_N(\MemCell.counter_value[1] ));
 sg13g2_nand3_1 _3992_ (.B(\MemCell.counter_value[0] ),
    .C(_1450_),
    .A(_1844_),
    .Y(_1451_));
 sg13g2_a22oi_1 _3993_ (.Y(_1452_),
    .B1(\MemCell.counter_value[1] ),
    .B2(_1843_),
    .A2(\MemCell.counter_value[2] ),
    .A1(_1842_));
 sg13g2_nand2b_1 _3994_ (.Y(_1453_),
    .B(\pwm_module.counter2[3] ),
    .A_N(\MemCell.counter_value[3] ));
 sg13g2_o21ai_1 _3995_ (.B1(_1453_),
    .Y(_1454_),
    .A1(_1842_),
    .A2(\MemCell.counter_value[2] ));
 sg13g2_a21o_1 _3996_ (.A2(_1452_),
    .A1(_1451_),
    .B1(_1454_),
    .X(_1455_));
 sg13g2_nand2b_1 _3997_ (.Y(_1456_),
    .B(\MemCell.counter_value[4] ),
    .A_N(\pwm_module.counter2[4] ));
 sg13g2_nand2b_1 _3998_ (.Y(_1457_),
    .B(\MemCell.counter_value[3] ),
    .A_N(\pwm_module.counter2[3] ));
 sg13g2_nand2b_1 _3999_ (.Y(_1458_),
    .B(\MemCell.counter_value[6] ),
    .A_N(\pwm_module.counter2[6] ));
 sg13g2_nand2b_1 _4000_ (.Y(_1459_),
    .B(\MemCell.counter_value[5] ),
    .A_N(\pwm_module.counter2[5] ));
 sg13g2_nand2b_1 _4001_ (.Y(_1460_),
    .B(\MemCell.counter_value[7] ),
    .A_N(\pwm_module.counter2[7] ));
 sg13g2_a21oi_1 _4002_ (.A1(_1834_),
    .A2(\MemCell.counter_value[8] ),
    .Y(_1461_),
    .B1(_1440_));
 sg13g2_and2_1 _4003_ (.A(_1422_),
    .B(_1426_),
    .X(_1462_));
 sg13g2_nor2_1 _4004_ (.A(_1428_),
    .B(_1429_),
    .Y(_1463_));
 sg13g2_a221oi_1 _4005_ (.B2(_1421_),
    .C1(_1462_),
    .B1(_1463_),
    .A1(_1430_),
    .Y(_1464_),
    .A2(_1443_));
 sg13g2_nand3_1 _4006_ (.B(_1458_),
    .C(_1459_),
    .A(_1444_),
    .Y(_1465_));
 sg13g2_o21ai_1 _4007_ (.B1(_1446_),
    .Y(_1466_),
    .A1(_1449_),
    .A2(_1465_));
 sg13g2_nand4_1 _4008_ (.B(_1456_),
    .C(_1457_),
    .A(_1445_),
    .Y(_1467_),
    .D(_1460_));
 sg13g2_nor4_1 _4009_ (.A(_1447_),
    .B(_1448_),
    .C(_1465_),
    .D(_1467_),
    .Y(_1468_));
 sg13g2_a22oi_1 _4010_ (.Y(_1469_),
    .B1(_1468_),
    .B2(_1455_),
    .A2(_1466_),
    .A1(_1460_));
 sg13g2_nand4_1 _4011_ (.B(_1438_),
    .C(_1441_),
    .A(_1430_),
    .Y(_1470_),
    .D(_1461_));
 sg13g2_o21ai_1 _4012_ (.B1(_1464_),
    .Y(_1471_),
    .A1(_1469_),
    .A2(_1470_));
 sg13g2_nand2b_1 _4013_ (.Y(_1472_),
    .B(\pwm_module.counter2[31] ),
    .A_N(\MemCell.counter_value[31] ));
 sg13g2_o21ai_1 _4014_ (.B1(_1472_),
    .Y(_1473_),
    .A1(_1807_),
    .A2(\MemCell.counter_value[30] ));
 sg13g2_nand2b_1 _4015_ (.Y(_1474_),
    .B(\MemCell.counter_value[29] ),
    .A_N(\pwm_module.counter2[29] ));
 sg13g2_nand2b_1 _4016_ (.Y(_1475_),
    .B(\MemCell.counter_value[31] ),
    .A_N(\pwm_module.counter2[31] ));
 sg13g2_nand2b_1 _4017_ (.Y(_1476_),
    .B(\MemCell.counter_value[30] ),
    .A_N(\pwm_module.counter2[30] ));
 sg13g2_nand3_1 _4018_ (.B(_1475_),
    .C(_1476_),
    .A(_1474_),
    .Y(_1477_));
 sg13g2_nor2_1 _4019_ (.A(_1473_),
    .B(_1477_),
    .Y(_1478_));
 sg13g2_nor2_1 _4020_ (.A(\pwm_module.counter2[28] ),
    .B(_1875_),
    .Y(_1479_));
 sg13g2_nand2b_1 _4021_ (.Y(_1480_),
    .B(\pwm_module.counter2[29] ),
    .A_N(\MemCell.counter_value[29] ));
 sg13g2_o21ai_1 _4022_ (.B1(_1480_),
    .Y(_1481_),
    .A1(_1810_),
    .A2(\MemCell.counter_value[28] ));
 sg13g2_nor4_2 _4023_ (.A(_1473_),
    .B(_1477_),
    .C(_1479_),
    .Y(_1482_),
    .D(_1481_));
 sg13g2_nand2b_1 _4024_ (.Y(_1483_),
    .B(\pwm_module.counter2[26] ),
    .A_N(\MemCell.counter_value[26] ));
 sg13g2_nand2b_1 _4025_ (.Y(_1484_),
    .B(\pwm_module.counter2[27] ),
    .A_N(\MemCell.counter_value[27] ));
 sg13g2_nand2_1 _4026_ (.Y(_1485_),
    .A(_1483_),
    .B(_1484_));
 sg13g2_nand2b_1 _4027_ (.Y(_1486_),
    .B(\MemCell.counter_value[27] ),
    .A_N(\pwm_module.counter2[27] ));
 sg13g2_nand2b_1 _4028_ (.Y(_1487_),
    .B(\MemCell.counter_value[26] ),
    .A_N(\pwm_module.counter2[26] ));
 sg13g2_nor2b_1 _4029_ (.A(\pwm_module.counter2[25] ),
    .B_N(\MemCell.counter_value[25] ),
    .Y(_1488_));
 sg13g2_nand2b_1 _4030_ (.Y(_1489_),
    .B(\pwm_module.counter2[24] ),
    .A_N(\MemCell.counter_value[24] ));
 sg13g2_nand2b_1 _4031_ (.Y(_1490_),
    .B(\pwm_module.counter2[25] ),
    .A_N(\MemCell.counter_value[25] ));
 sg13g2_and4_1 _4032_ (.A(_1483_),
    .B(_1484_),
    .C(_1486_),
    .D(_1487_),
    .X(_1491_));
 sg13g2_xnor2_1 _4033_ (.Y(_1492_),
    .A(\pwm_module.counter2[24] ),
    .B(\MemCell.counter_value[24] ));
 sg13g2_nor2b_1 _4034_ (.A(_1488_),
    .B_N(_1490_),
    .Y(_1493_));
 sg13g2_nand4_1 _4035_ (.B(_1491_),
    .C(_1492_),
    .A(_1482_),
    .Y(_1494_),
    .D(_1493_));
 sg13g2_inv_1 _4036_ (.Y(_1495_),
    .A(_1494_));
 sg13g2_nand2b_1 _4037_ (.Y(_1496_),
    .B(\pwm_module.counter2[18] ),
    .A_N(\MemCell.counter_value[18] ));
 sg13g2_nand2b_1 _4038_ (.Y(_1497_),
    .B(\pwm_module.counter2[19] ),
    .A_N(\MemCell.counter_value[19] ));
 sg13g2_nand2_1 _4039_ (.Y(_1498_),
    .A(_1496_),
    .B(_1497_));
 sg13g2_nand2b_1 _4040_ (.Y(_1499_),
    .B(\MemCell.counter_value[19] ),
    .A_N(\pwm_module.counter2[19] ));
 sg13g2_nand2b_1 _4041_ (.Y(_1500_),
    .B(\MemCell.counter_value[18] ),
    .A_N(\pwm_module.counter2[18] ));
 sg13g2_nor2_1 _4042_ (.A(net648),
    .B(_1895_),
    .Y(_1501_));
 sg13g2_nand4_1 _4043_ (.B(_1497_),
    .C(_1499_),
    .A(_1496_),
    .Y(_1502_),
    .D(_1500_));
 sg13g2_nand2b_1 _4044_ (.Y(_1503_),
    .B(\MemCell.counter_value[21] ),
    .A_N(\pwm_module.counter2[21] ));
 sg13g2_o21ai_1 _4045_ (.B1(_1503_),
    .Y(_1504_),
    .A1(\pwm_module.counter2[22] ),
    .A2(_1886_));
 sg13g2_a221oi_1 _4046_ (.B2(_1820_),
    .C1(_1504_),
    .B1(\MemCell.counter_value[20] ),
    .A1(_1816_),
    .Y(_1505_),
    .A2(\MemCell.counter_value[23] ));
 sg13g2_a22oi_1 _4047_ (.Y(_1506_),
    .B1(_1889_),
    .B2(\pwm_module.counter2[20] ),
    .A2(_1887_),
    .A1(\pwm_module.counter2[21] ));
 sg13g2_a22oi_1 _4048_ (.Y(_1507_),
    .B1(_1886_),
    .B2(\pwm_module.counter2[22] ),
    .A2(_1884_),
    .A1(\pwm_module.counter2[23] ));
 sg13g2_nand3_1 _4049_ (.B(_1506_),
    .C(_1507_),
    .A(_1505_),
    .Y(_1508_));
 sg13g2_nor2_1 _4050_ (.A(\pwm_module.counter2[16] ),
    .B(_1897_),
    .Y(_1509_));
 sg13g2_nor2b_1 _4051_ (.A(\MemCell.counter_value[17] ),
    .B_N(net648),
    .Y(_1510_));
 sg13g2_nor2b_1 _4052_ (.A(\MemCell.counter_value[16] ),
    .B_N(\pwm_module.counter2[16] ),
    .Y(_1511_));
 sg13g2_nor2_1 _4053_ (.A(_1510_),
    .B(_1511_),
    .Y(_1512_));
 sg13g2_or4_1 _4054_ (.A(_1501_),
    .B(_1509_),
    .C(_1510_),
    .D(_1511_),
    .X(_1513_));
 sg13g2_nor4_1 _4055_ (.A(_1494_),
    .B(_1502_),
    .C(_1508_),
    .D(_1513_),
    .Y(_1514_));
 sg13g2_nor3_1 _4056_ (.A(_1501_),
    .B(_1502_),
    .C(_1512_),
    .Y(_1515_));
 sg13g2_a21oi_1 _4057_ (.A1(_1498_),
    .A2(_1499_),
    .Y(_1516_),
    .B1(_1515_));
 sg13g2_o21ai_1 _4058_ (.B1(_1507_),
    .Y(_1517_),
    .A1(_1504_),
    .A2(_1506_));
 sg13g2_o21ai_1 _4059_ (.B1(_1517_),
    .Y(_1518_),
    .A1(\pwm_module.counter2[23] ),
    .A2(_1884_));
 sg13g2_o21ai_1 _4060_ (.B1(_1518_),
    .Y(_1519_),
    .A1(_1508_),
    .A2(_1516_));
 sg13g2_o21ai_1 _4061_ (.B1(_1490_),
    .Y(_1520_),
    .A1(_1488_),
    .A2(_1489_));
 sg13g2_a22oi_1 _4062_ (.Y(_1521_),
    .B1(_1491_),
    .B2(_1520_),
    .A2(_1486_),
    .A1(_1485_));
 sg13g2_nand2b_1 _4063_ (.Y(_1522_),
    .B(_1482_),
    .A_N(_1521_));
 sg13g2_a22oi_1 _4064_ (.Y(_1523_),
    .B1(_1478_),
    .B2(_1481_),
    .A2(_1475_),
    .A1(_1473_));
 sg13g2_nand3_1 _4065_ (.B(_1522_),
    .C(_1523_),
    .A(net651),
    .Y(_1524_));
 sg13g2_a221oi_1 _4066_ (.B2(_1495_),
    .C1(_1524_),
    .B1(_1519_),
    .A1(_1471_),
    .Y(_1525_),
    .A2(_1514_));
 sg13g2_a21oi_2 _4067_ (.B1(_1525_),
    .Y(_1526_),
    .A2(_0963_),
    .A1(net646));
 sg13g2_a21oi_2 _4068_ (.B1(_1844_),
    .Y(_1527_),
    .A2(net612),
    .A1(net644));
 sg13g2_nor2_1 _4069_ (.A(net362),
    .B(net585),
    .Y(_1528_));
 sg13g2_nor3_1 _4070_ (.A(net577),
    .B(_1527_),
    .C(_1528_),
    .Y(_0319_));
 sg13g2_xnor2_1 _4071_ (.Y(_1529_),
    .A(net649),
    .B(_1527_));
 sg13g2_nor2_1 _4072_ (.A(net577),
    .B(_1529_),
    .Y(_0320_));
 sg13g2_and3_1 _4073_ (.X(_1530_),
    .A(\pwm_module.counter2[2] ),
    .B(net649),
    .C(\pwm_module.counter2[0] ));
 sg13g2_nand3_1 _4074_ (.B(net649),
    .C(\pwm_module.counter2[0] ),
    .A(\pwm_module.counter2[2] ),
    .Y(_1531_));
 sg13g2_a21oi_2 _4075_ (.B1(_1531_),
    .Y(_1532_),
    .A2(net612),
    .A1(net645));
 sg13g2_a21oi_1 _4076_ (.A1(net164),
    .A2(_1527_),
    .Y(_1533_),
    .B1(\pwm_module.counter2[2] ));
 sg13g2_nor3_1 _4077_ (.A(net577),
    .B(_1532_),
    .C(net165),
    .Y(_0321_));
 sg13g2_xnor2_1 _4078_ (.Y(_1534_),
    .A(net441),
    .B(_1532_));
 sg13g2_nor2_1 _4079_ (.A(net577),
    .B(_1534_),
    .Y(_0322_));
 sg13g2_a21oi_1 _4080_ (.A1(\pwm_module.counter2[3] ),
    .A2(_1532_),
    .Y(_1535_),
    .B1(net300));
 sg13g2_nor4_1 _4081_ (.A(_1839_),
    .B(_1841_),
    .C(_1418_),
    .D(_1531_),
    .Y(_1536_));
 sg13g2_nand3_1 _4082_ (.B(\pwm_module.counter2[3] ),
    .C(_1532_),
    .A(net300),
    .Y(_1537_));
 sg13g2_nor3_1 _4083_ (.A(net577),
    .B(net301),
    .C(_1536_),
    .Y(_0323_));
 sg13g2_nor3_2 _4084_ (.A(_1838_),
    .B(_1839_),
    .C(_1841_),
    .Y(_1538_));
 sg13g2_a21o_1 _4085_ (.A2(_1538_),
    .A1(_1532_),
    .B1(net577),
    .X(_1539_));
 sg13g2_a21oi_1 _4086_ (.A1(_1838_),
    .A2(_1537_),
    .Y(_0324_),
    .B1(_1539_));
 sg13g2_a21oi_1 _4087_ (.A1(_1532_),
    .A2(_1538_),
    .Y(_1540_),
    .B1(net349));
 sg13g2_and3_1 _4088_ (.X(_1541_),
    .A(net349),
    .B(_1532_),
    .C(_1538_));
 sg13g2_nand3_1 _4089_ (.B(_1532_),
    .C(_1538_),
    .A(net349),
    .Y(_1542_));
 sg13g2_nor3_1 _4090_ (.A(net577),
    .B(_1540_),
    .C(_1541_),
    .Y(_0325_));
 sg13g2_nand4_1 _4091_ (.B(\pwm_module.counter2[6] ),
    .C(_1530_),
    .A(\pwm_module.counter2[7] ),
    .Y(_1543_),
    .D(_1538_));
 sg13g2_and4_1 _4092_ (.A(\pwm_module.counter2[3] ),
    .B(\pwm_module.counter2[2] ),
    .C(net649),
    .D(\pwm_module.counter2[0] ),
    .X(_1544_));
 sg13g2_nand4_1 _4093_ (.B(\pwm_module.counter2[5] ),
    .C(\pwm_module.counter2[4] ),
    .A(\pwm_module.counter2[7] ),
    .Y(_1545_),
    .D(_1544_));
 sg13g2_nor2_1 _4094_ (.A(_1836_),
    .B(_1545_),
    .Y(_1546_));
 sg13g2_inv_1 _4095_ (.Y(_1547_),
    .A(_1546_));
 sg13g2_a21oi_2 _4096_ (.B1(_1547_),
    .Y(_1548_),
    .A2(net612),
    .A1(net645));
 sg13g2_and4_1 _4097_ (.A(\pwm_module.counter2[7] ),
    .B(\pwm_module.counter2[6] ),
    .C(_1530_),
    .D(_1538_),
    .X(_1549_));
 sg13g2_inv_1 _4098_ (.Y(_1550_),
    .A(_1549_));
 sg13g2_a21oi_2 _4099_ (.B1(_1550_),
    .Y(_1551_),
    .A2(net612),
    .A1(net644));
 sg13g2_a221oi_1 _4100_ (.B2(net585),
    .C1(net577),
    .B1(_1546_),
    .A1(_1835_),
    .Y(_0326_),
    .A2(_1542_));
 sg13g2_xnor2_1 _4101_ (.Y(_1552_),
    .A(net452),
    .B(_1548_));
 sg13g2_nor2_1 _4102_ (.A(_1526_),
    .B(_1552_),
    .Y(_0327_));
 sg13g2_a21oi_1 _4103_ (.A1(\pwm_module.counter2[8] ),
    .A2(_1551_),
    .Y(_1553_),
    .B1(net295));
 sg13g2_nor4_1 _4104_ (.A(_1832_),
    .B(_1834_),
    .C(_1418_),
    .D(_1550_),
    .Y(_1554_));
 sg13g2_nand3_1 _4105_ (.B(\pwm_module.counter2[8] ),
    .C(_1548_),
    .A(net295),
    .Y(_1555_));
 sg13g2_nor3_1 _4106_ (.A(net578),
    .B(net296),
    .C(_1554_),
    .Y(_0328_));
 sg13g2_and3_1 _4107_ (.X(_1556_),
    .A(\pwm_module.counter2[10] ),
    .B(\pwm_module.counter2[9] ),
    .C(\pwm_module.counter2[8] ));
 sg13g2_a221oi_1 _4108_ (.B2(_1548_),
    .C1(net578),
    .B1(_1556_),
    .A1(_1830_),
    .Y(_0329_),
    .A2(_1555_));
 sg13g2_a21oi_1 _4109_ (.A1(_1548_),
    .A2(_1556_),
    .Y(_1557_),
    .B1(net322));
 sg13g2_and2_1 _4110_ (.A(\pwm_module.counter2[11] ),
    .B(_1556_),
    .X(_1558_));
 sg13g2_nand2_2 _4111_ (.Y(_1559_),
    .A(\pwm_module.counter2[11] ),
    .B(_1556_));
 sg13g2_nor3_2 _4112_ (.A(_1836_),
    .B(_1545_),
    .C(_1559_),
    .Y(_1560_));
 sg13g2_inv_1 _4113_ (.Y(_1561_),
    .A(_1560_));
 sg13g2_a21oi_2 _4114_ (.B1(_1561_),
    .Y(_1562_),
    .A2(net612),
    .A1(net645));
 sg13g2_nor3_1 _4115_ (.A(net578),
    .B(_1557_),
    .C(_1562_),
    .Y(_0330_));
 sg13g2_nor2_1 _4116_ (.A(net282),
    .B(_1562_),
    .Y(_1563_));
 sg13g2_nor4_2 _4117_ (.A(_1829_),
    .B(_1418_),
    .C(_1543_),
    .Y(_1564_),
    .D(_1559_));
 sg13g2_nand2_1 _4118_ (.Y(_1565_),
    .A(net282),
    .B(_1562_));
 sg13g2_nor3_1 _4119_ (.A(net578),
    .B(_1563_),
    .C(_1564_),
    .Y(_0331_));
 sg13g2_nor2_1 _4120_ (.A(_1827_),
    .B(_1829_),
    .Y(_1566_));
 sg13g2_nand2_1 _4121_ (.Y(_1567_),
    .A(_1562_),
    .B(_1566_));
 sg13g2_a221oi_1 _4122_ (.B2(_1562_),
    .C1(net578),
    .B1(_1566_),
    .A1(_1827_),
    .Y(_0332_),
    .A2(_1565_));
 sg13g2_nor2_1 _4123_ (.A(_1825_),
    .B(_1827_),
    .Y(_1568_));
 sg13g2_nand4_1 _4124_ (.B(_1551_),
    .C(_1558_),
    .A(net377),
    .Y(_1569_),
    .D(_1566_));
 sg13g2_a221oi_1 _4125_ (.B2(_1564_),
    .C1(net578),
    .B1(_1568_),
    .A1(_1825_),
    .Y(_0333_),
    .A2(_1567_));
 sg13g2_and4_2 _4126_ (.A(\pwm_module.counter2[15] ),
    .B(\pwm_module.counter2[14] ),
    .C(_1560_),
    .D(_1566_),
    .X(_1570_));
 sg13g2_a221oi_1 _4127_ (.B2(net585),
    .C1(net578),
    .B1(_1570_),
    .A1(_1823_),
    .Y(_0334_),
    .A2(_1569_));
 sg13g2_a21oi_1 _4128_ (.A1(net581),
    .A2(_1570_),
    .Y(_1571_),
    .B1(net499));
 sg13g2_and2_1 _4129_ (.A(\pwm_module.counter2[16] ),
    .B(_1570_),
    .X(_1572_));
 sg13g2_and2_1 _4130_ (.A(net581),
    .B(_1572_),
    .X(_1573_));
 sg13g2_nor3_1 _4131_ (.A(net580),
    .B(_1571_),
    .C(_1573_),
    .Y(_0335_));
 sg13g2_a21oi_1 _4132_ (.A1(net581),
    .A2(_1572_),
    .Y(_1574_),
    .B1(net648));
 sg13g2_nand2_1 _4133_ (.Y(_1575_),
    .A(net648),
    .B(\pwm_module.counter2[16] ));
 sg13g2_and3_1 _4134_ (.X(_1576_),
    .A(net648),
    .B(net581),
    .C(_1572_));
 sg13g2_nand3_1 _4135_ (.B(net581),
    .C(_1572_),
    .A(net648),
    .Y(_1577_));
 sg13g2_nor3_1 _4136_ (.A(net580),
    .B(_1574_),
    .C(_1576_),
    .Y(_0336_));
 sg13g2_and2_1 _4137_ (.A(\pwm_module.counter2[18] ),
    .B(net648),
    .X(_1578_));
 sg13g2_nand3_1 _4138_ (.B(_1572_),
    .C(_1578_),
    .A(net581),
    .Y(_1579_));
 sg13g2_a221oi_1 _4139_ (.B2(_1573_),
    .C1(net580),
    .B1(_1578_),
    .A1(_1822_),
    .Y(_0337_),
    .A2(_1577_));
 sg13g2_nor3_1 _4140_ (.A(_1821_),
    .B(_1822_),
    .C(_1575_),
    .Y(_1580_));
 sg13g2_and2_1 _4141_ (.A(_1570_),
    .B(_1580_),
    .X(_1581_));
 sg13g2_nand2_1 _4142_ (.Y(_1582_),
    .A(net581),
    .B(_1581_));
 sg13g2_a221oi_1 _4143_ (.B2(net584),
    .C1(net580),
    .B1(_1581_),
    .A1(_1821_),
    .Y(_0338_),
    .A2(_1579_));
 sg13g2_and2_1 _4144_ (.A(\pwm_module.counter2[20] ),
    .B(_1581_),
    .X(_1583_));
 sg13g2_a221oi_1 _4145_ (.B2(net581),
    .C1(net580),
    .B1(_1583_),
    .A1(_1820_),
    .Y(_0339_),
    .A2(_1582_));
 sg13g2_a21oi_1 _4146_ (.A1(net582),
    .A2(_1583_),
    .Y(_1584_),
    .B1(net455));
 sg13g2_and3_1 _4147_ (.X(_1585_),
    .A(net455),
    .B(net582),
    .C(_1583_));
 sg13g2_nand3_1 _4148_ (.B(net582),
    .C(_1583_),
    .A(\pwm_module.counter2[21] ),
    .Y(_1586_));
 sg13g2_nor3_1 _4149_ (.A(net579),
    .B(_1584_),
    .C(_1585_),
    .Y(_0340_));
 sg13g2_and3_1 _4150_ (.X(_1587_),
    .A(\pwm_module.counter2[22] ),
    .B(\pwm_module.counter2[21] ),
    .C(\pwm_module.counter2[20] ));
 sg13g2_nand2_1 _4151_ (.Y(_1588_),
    .A(_1581_),
    .B(_1587_));
 sg13g2_nand2b_1 _4152_ (.Y(_1589_),
    .B(net582),
    .A_N(_1588_));
 sg13g2_a21oi_1 _4153_ (.A1(_1525_),
    .A2(_1588_),
    .Y(_1590_),
    .B1(_1418_));
 sg13g2_a21oi_1 _4154_ (.A1(_1817_),
    .A2(_1586_),
    .Y(_0341_),
    .B1(_1590_));
 sg13g2_nand4_1 _4155_ (.B(_1570_),
    .C(_1580_),
    .A(\pwm_module.counter2[23] ),
    .Y(_1591_),
    .D(_1587_));
 sg13g2_inv_1 _4156_ (.Y(_1592_),
    .A(_1591_));
 sg13g2_a21oi_2 _4157_ (.B1(_1591_),
    .Y(_1593_),
    .A2(net612),
    .A1(net646));
 sg13g2_a221oi_1 _4158_ (.B2(net582),
    .C1(net579),
    .B1(_1592_),
    .A1(_1816_),
    .Y(_0342_),
    .A2(_1589_));
 sg13g2_nor2_1 _4159_ (.A(net523),
    .B(_1593_),
    .Y(_1594_));
 sg13g2_and2_1 _4160_ (.A(net523),
    .B(_1593_),
    .X(_1595_));
 sg13g2_nand2_1 _4161_ (.Y(_1596_),
    .A(net523),
    .B(_1593_));
 sg13g2_nor3_1 _4162_ (.A(net580),
    .B(_1594_),
    .C(_1595_),
    .Y(_0343_));
 sg13g2_and2_1 _4163_ (.A(\pwm_module.counter2[25] ),
    .B(\pwm_module.counter2[24] ),
    .X(_1597_));
 sg13g2_a221oi_1 _4164_ (.B2(_1593_),
    .C1(net579),
    .B1(_1597_),
    .A1(_1814_),
    .Y(_0344_),
    .A2(_1596_));
 sg13g2_a21oi_1 _4165_ (.A1(_1593_),
    .A2(_1597_),
    .Y(_1598_),
    .B1(net315));
 sg13g2_and3_1 _4166_ (.X(_1599_),
    .A(net315),
    .B(_1592_),
    .C(_1597_));
 sg13g2_a21oi_1 _4167_ (.A1(net583),
    .A2(_1599_),
    .Y(_1600_),
    .B1(net579));
 sg13g2_nor2b_1 _4168_ (.A(_1598_),
    .B_N(_1600_),
    .Y(_0345_));
 sg13g2_a21oi_1 _4169_ (.A1(net583),
    .A2(_1599_),
    .Y(_1601_),
    .B1(net316));
 sg13g2_and3_1 _4170_ (.X(_1602_),
    .A(net316),
    .B(net583),
    .C(_1599_));
 sg13g2_nand3_1 _4171_ (.B(net582),
    .C(_1599_),
    .A(net316),
    .Y(_1603_));
 sg13g2_nor3_1 _4172_ (.A(net579),
    .B(_1601_),
    .C(_1602_),
    .Y(_0346_));
 sg13g2_nand4_1 _4173_ (.B(net316),
    .C(net315),
    .A(\pwm_module.counter2[28] ),
    .Y(_1604_),
    .D(_1597_));
 sg13g2_nor2_1 _4174_ (.A(_1591_),
    .B(_1604_),
    .Y(_1605_));
 sg13g2_or2_1 _4175_ (.X(_1606_),
    .B(_1604_),
    .A(_1591_));
 sg13g2_a21oi_1 _4176_ (.A1(net646),
    .A2(_0963_),
    .Y(_1607_),
    .B1(_1606_));
 sg13g2_or2_1 _4177_ (.X(_1608_),
    .B(_1607_),
    .A(net579));
 sg13g2_a21oi_1 _4178_ (.A1(_1810_),
    .A2(_1603_),
    .Y(_0347_),
    .B1(_1608_));
 sg13g2_nand4_1 _4179_ (.B(net583),
    .C(_1525_),
    .A(_1809_),
    .Y(_1609_),
    .D(_1605_));
 sg13g2_o21ai_1 _4180_ (.B1(_1609_),
    .Y(_0348_),
    .A1(_1809_),
    .A2(_1608_));
 sg13g2_nand2_1 _4181_ (.Y(_1610_),
    .A(\pwm_module.counter2[29] ),
    .B(_1607_));
 sg13g2_nor3_1 _4182_ (.A(_1807_),
    .B(_1809_),
    .C(_1606_),
    .Y(_1611_));
 sg13g2_a221oi_1 _4183_ (.B2(net582),
    .C1(net579),
    .B1(_1611_),
    .A1(_1807_),
    .Y(_0349_),
    .A2(_1610_));
 sg13g2_a21oi_1 _4184_ (.A1(net582),
    .A2(_1611_),
    .Y(_1612_),
    .B1(net179));
 sg13g2_nor2_1 _4185_ (.A(net579),
    .B(net180),
    .Y(_0350_));
 sg13g2_nor2_2 _4186_ (.A(_1036_),
    .B(_1326_),
    .Y(_1613_));
 sg13g2_nand2_1 _4187_ (.Y(_1614_),
    .A(net679),
    .B(net618));
 sg13g2_o21ai_1 _4188_ (.B1(_1614_),
    .Y(_0351_),
    .A1(_1815_),
    .A2(net618));
 sg13g2_nand2_1 _4189_ (.Y(_1615_),
    .A(net676),
    .B(net618));
 sg13g2_o21ai_1 _4190_ (.B1(_1615_),
    .Y(_0352_),
    .A1(_1813_),
    .A2(net618));
 sg13g2_mux2_1 _4191_ (.A0(net157),
    .A1(net672),
    .S(net618),
    .X(_0353_));
 sg13g2_mux2_1 _4192_ (.A0(net85),
    .A1(net668),
    .S(net618),
    .X(_0354_));
 sg13g2_nand2_1 _4193_ (.Y(_1616_),
    .A(net665),
    .B(net619));
 sg13g2_o21ai_1 _4194_ (.B1(_1616_),
    .Y(_0355_),
    .A1(_1811_),
    .A2(net619));
 sg13g2_nand2_1 _4195_ (.Y(_1617_),
    .A(net662),
    .B(net619));
 sg13g2_o21ai_1 _4196_ (.B1(_1617_),
    .Y(_0356_),
    .A1(_1808_),
    .A2(net619));
 sg13g2_nand2_1 _4197_ (.Y(_1618_),
    .A(net659),
    .B(net619));
 sg13g2_o21ai_1 _4198_ (.B1(_1618_),
    .Y(_0357_),
    .A1(_1806_),
    .A2(net619));
 sg13g2_nand2_1 _4199_ (.Y(_1619_),
    .A(net656),
    .B(net618));
 sg13g2_o21ai_1 _4200_ (.B1(_1619_),
    .Y(_0358_),
    .A1(_1805_),
    .A2(net618));
 sg13g2_nand2_1 _4201_ (.Y(_1620_),
    .A(net646),
    .B(_0790_));
 sg13g2_nand2b_1 _4202_ (.Y(_1621_),
    .B(\pwm_module.counter1[31] ),
    .A_N(\MemCell.counter_value[31] ));
 sg13g2_o21ai_1 _4203_ (.B1(_1621_),
    .Y(_1622_),
    .A1(\MemCell.counter_value[30] ),
    .A2(_1918_));
 sg13g2_nand2b_1 _4204_ (.Y(_1623_),
    .B(\MemCell.counter_value[30] ),
    .A_N(\pwm_module.counter1[30] ));
 sg13g2_nand2b_1 _4205_ (.Y(_1624_),
    .B(\MemCell.counter_value[31] ),
    .A_N(\pwm_module.counter1[31] ));
 sg13g2_nand2b_1 _4206_ (.Y(_1625_),
    .B(\MemCell.counter_value[29] ),
    .A_N(\pwm_module.counter1[29] ));
 sg13g2_nand3_1 _4207_ (.B(_1624_),
    .C(_1625_),
    .A(_1623_),
    .Y(_1626_));
 sg13g2_nor2_1 _4208_ (.A(_1622_),
    .B(_1626_),
    .Y(_1627_));
 sg13g2_nor2b_1 _4209_ (.A(\MemCell.counter_value[29] ),
    .B_N(\pwm_module.counter1[29] ),
    .Y(_1628_));
 sg13g2_a21o_1 _4210_ (.A2(\pwm_module.counter1[28] ),
    .A1(_1875_),
    .B1(_1628_),
    .X(_1629_));
 sg13g2_nor2_1 _4211_ (.A(_1875_),
    .B(\pwm_module.counter1[28] ),
    .Y(_1630_));
 sg13g2_nor4_2 _4212_ (.A(_1622_),
    .B(_1626_),
    .C(_1629_),
    .Y(_1631_),
    .D(_1630_));
 sg13g2_nand2b_1 _4213_ (.Y(_1632_),
    .B(\pwm_module.counter1[26] ),
    .A_N(\MemCell.counter_value[26] ));
 sg13g2_nor2_1 _4214_ (.A(_1876_),
    .B(\pwm_module.counter1[27] ),
    .Y(_1633_));
 sg13g2_o21ai_1 _4215_ (.B1(_1632_),
    .Y(_1634_),
    .A1(_1876_),
    .A2(\pwm_module.counter1[27] ));
 sg13g2_nand2b_1 _4216_ (.Y(_1635_),
    .B(\MemCell.counter_value[26] ),
    .A_N(\pwm_module.counter1[26] ));
 sg13g2_nand2b_1 _4217_ (.Y(_1636_),
    .B(\MemCell.counter_value[25] ),
    .A_N(\pwm_module.counter1[25] ));
 sg13g2_nand2b_1 _4218_ (.Y(_1637_),
    .B(\pwm_module.counter1[27] ),
    .A_N(\MemCell.counter_value[27] ));
 sg13g2_nand3_1 _4219_ (.B(_1636_),
    .C(_1637_),
    .A(_1635_),
    .Y(_1638_));
 sg13g2_nor2b_1 _4220_ (.A(\MemCell.counter_value[25] ),
    .B_N(\pwm_module.counter1[25] ),
    .Y(_1639_));
 sg13g2_a21oi_1 _4221_ (.A1(_1882_),
    .A2(\pwm_module.counter1[24] ),
    .Y(_1640_),
    .B1(_1639_));
 sg13g2_a21o_1 _4222_ (.A2(\pwm_module.counter1[24] ),
    .A1(_1882_),
    .B1(_1639_),
    .X(_1641_));
 sg13g2_nor2_1 _4223_ (.A(_1882_),
    .B(\pwm_module.counter1[24] ),
    .Y(_1642_));
 sg13g2_nor4_2 _4224_ (.A(_1634_),
    .B(_1638_),
    .C(_1641_),
    .Y(_1643_),
    .D(_1642_));
 sg13g2_nand2_2 _4225_ (.Y(_1644_),
    .A(_1631_),
    .B(_1643_));
 sg13g2_nor2b_1 _4226_ (.A(\MemCell.counter_value[23] ),
    .B_N(\pwm_module.counter1[23] ),
    .Y(_1645_));
 sg13g2_nor2b_1 _4227_ (.A(\MemCell.counter_value[22] ),
    .B_N(\pwm_module.counter1[22] ),
    .Y(_1646_));
 sg13g2_nor2_1 _4228_ (.A(_1645_),
    .B(_1646_),
    .Y(_1647_));
 sg13g2_nand2b_1 _4229_ (.Y(_1648_),
    .B(\MemCell.counter_value[22] ),
    .A_N(\pwm_module.counter1[22] ));
 sg13g2_o21ai_1 _4230_ (.B1(_1648_),
    .Y(_1649_),
    .A1(_1887_),
    .A2(\pwm_module.counter1[21] ));
 sg13g2_nor2b_1 _4231_ (.A(\MemCell.counter_value[20] ),
    .B_N(\pwm_module.counter1[20] ),
    .Y(_1650_));
 sg13g2_nor2b_1 _4232_ (.A(\MemCell.counter_value[21] ),
    .B_N(\pwm_module.counter1[21] ),
    .Y(_1651_));
 sg13g2_nor4_1 _4233_ (.A(_1645_),
    .B(_1646_),
    .C(_1650_),
    .D(_1651_),
    .Y(_1652_));
 sg13g2_a221oi_1 _4234_ (.B2(_1649_),
    .C1(_1652_),
    .B1(_1647_),
    .A1(\MemCell.counter_value[23] ),
    .Y(_1653_),
    .A2(_1920_));
 sg13g2_nand3_1 _4235_ (.B(_1643_),
    .C(_1653_),
    .A(_1631_),
    .Y(_1654_));
 sg13g2_nor3_1 _4236_ (.A(_1634_),
    .B(_1638_),
    .C(_1640_),
    .Y(_1655_));
 sg13g2_o21ai_1 _4237_ (.B1(_1637_),
    .Y(_1656_),
    .A1(_1632_),
    .A2(_1633_));
 sg13g2_o21ai_1 _4238_ (.B1(_1631_),
    .Y(_1657_),
    .A1(_1655_),
    .A2(_1656_));
 sg13g2_a22oi_1 _4239_ (.Y(_1658_),
    .B1(_1627_),
    .B2(_1629_),
    .A2(_1624_),
    .A1(_1622_));
 sg13g2_nand4_1 _4240_ (.B(_1654_),
    .C(_1657_),
    .A(net651),
    .Y(_1659_),
    .D(_1658_));
 sg13g2_a22oi_1 _4241_ (.Y(_1660_),
    .B1(_1923_),
    .B2(\MemCell.counter_value[20] ),
    .A2(_1920_),
    .A1(\MemCell.counter_value[23] ));
 sg13g2_nand2_1 _4242_ (.Y(_1661_),
    .A(_1652_),
    .B(_1660_));
 sg13g2_nor3_1 _4243_ (.A(_1644_),
    .B(_1649_),
    .C(_1661_),
    .Y(_1662_));
 sg13g2_nor2_1 _4244_ (.A(_1891_),
    .B(\pwm_module.counter1[19] ),
    .Y(_1663_));
 sg13g2_a22oi_1 _4245_ (.Y(_1664_),
    .B1(\pwm_module.counter1[18] ),
    .B2(_1893_),
    .A2(\pwm_module.counter1[19] ),
    .A1(_1891_));
 sg13g2_a22oi_1 _4246_ (.Y(_1665_),
    .B1(\pwm_module.counter1[17] ),
    .B2(_1895_),
    .A2(_1897_),
    .A1(\pwm_module.counter1[16] ));
 sg13g2_nor2_1 _4247_ (.A(_1893_),
    .B(\pwm_module.counter1[18] ),
    .Y(_1666_));
 sg13g2_nor2_1 _4248_ (.A(_1895_),
    .B(\pwm_module.counter1[17] ),
    .Y(_1667_));
 sg13g2_or3_1 _4249_ (.A(_1665_),
    .B(_1666_),
    .C(_1667_),
    .X(_1668_));
 sg13g2_a21oi_1 _4250_ (.A1(_1664_),
    .A2(_1668_),
    .Y(_1669_),
    .B1(_1663_));
 sg13g2_nand2b_1 _4251_ (.Y(_1670_),
    .B(\pwm_module.counter1[1] ),
    .A_N(\MemCell.counter_value[1] ));
 sg13g2_nor2b_1 _4252_ (.A(\pwm_module.counter1[0] ),
    .B_N(\MemCell.counter_value[0] ),
    .Y(_1671_));
 sg13g2_nor2b_1 _4253_ (.A(\pwm_module.counter1[1] ),
    .B_N(\MemCell.counter_value[1] ),
    .Y(_1672_));
 sg13g2_a221oi_1 _4254_ (.B2(_1671_),
    .C1(_1672_),
    .B1(_1670_),
    .A1(_1804_),
    .Y(_1673_),
    .A2(\MemCell.counter_value[2] ));
 sg13g2_nand2b_1 _4255_ (.Y(_1674_),
    .B(\pwm_module.counter1[3] ),
    .A_N(\MemCell.counter_value[3] ));
 sg13g2_o21ai_1 _4256_ (.B1(_1674_),
    .Y(_1675_),
    .A1(_1804_),
    .A2(\MemCell.counter_value[2] ));
 sg13g2_a22oi_1 _4257_ (.Y(_1676_),
    .B1(\MemCell.counter_value[3] ),
    .B2(_1803_),
    .A2(\MemCell.counter_value[4] ),
    .A1(_1801_));
 sg13g2_o21ai_1 _4258_ (.B1(_1676_),
    .Y(_1677_),
    .A1(_1673_),
    .A2(_1675_));
 sg13g2_a22oi_1 _4259_ (.Y(_1678_),
    .B1(_1914_),
    .B2(\pwm_module.counter1[4] ),
    .A2(_1912_),
    .A1(net647));
 sg13g2_nand2b_1 _4260_ (.Y(_1679_),
    .B(\MemCell.counter_value[5] ),
    .A_N(net647));
 sg13g2_o21ai_1 _4261_ (.B1(_1679_),
    .Y(_1680_),
    .A1(\pwm_module.counter1[6] ),
    .A2(_1911_));
 sg13g2_a21o_1 _4262_ (.A2(_1678_),
    .A1(_1677_),
    .B1(_1680_),
    .X(_1681_));
 sg13g2_a22oi_1 _4263_ (.Y(_1682_),
    .B1(_1911_),
    .B2(\pwm_module.counter1[6] ),
    .A2(_1910_),
    .A1(\pwm_module.counter1[7] ));
 sg13g2_nand2b_1 _4264_ (.Y(_1683_),
    .B(\pwm_module.counter1[14] ),
    .A_N(\MemCell.counter_value[14] ));
 sg13g2_o21ai_1 _4265_ (.B1(_1683_),
    .Y(_1684_),
    .A1(_1786_),
    .A2(\MemCell.counter_value[15] ));
 sg13g2_nand2b_1 _4266_ (.Y(_1685_),
    .B(\MemCell.counter_value[15] ),
    .A_N(\pwm_module.counter1[15] ));
 sg13g2_o21ai_1 _4267_ (.B1(_1685_),
    .Y(_1686_),
    .A1(\pwm_module.counter1[14] ),
    .A2(_1900_));
 sg13g2_nor2_1 _4268_ (.A(_1684_),
    .B(_1686_),
    .Y(_1687_));
 sg13g2_nand2b_1 _4269_ (.Y(_1688_),
    .B(\pwm_module.counter1[13] ),
    .A_N(\MemCell.counter_value[13] ));
 sg13g2_o21ai_1 _4270_ (.B1(_1688_),
    .Y(_1689_),
    .A1(_1791_),
    .A2(\MemCell.counter_value[12] ));
 sg13g2_nand2b_1 _4271_ (.Y(_1690_),
    .B(\MemCell.counter_value[13] ),
    .A_N(\pwm_module.counter1[13] ));
 sg13g2_o21ai_1 _4272_ (.B1(_1690_),
    .Y(_1691_),
    .A1(\pwm_module.counter1[12] ),
    .A2(_1903_));
 sg13g2_nor4_2 _4273_ (.A(_1684_),
    .B(_1686_),
    .C(_1689_),
    .Y(_1692_),
    .D(_1691_));
 sg13g2_nand2b_1 _4274_ (.Y(_1693_),
    .B(\pwm_module.counter1[10] ),
    .A_N(\MemCell.counter_value[10] ));
 sg13g2_o21ai_1 _4275_ (.B1(_1693_),
    .Y(_1694_),
    .A1(_1792_),
    .A2(\MemCell.counter_value[11] ));
 sg13g2_nor2_1 _4276_ (.A(\pwm_module.counter1[9] ),
    .B(_1906_),
    .Y(_1695_));
 sg13g2_nand2b_1 _4277_ (.Y(_1696_),
    .B(\MemCell.counter_value[11] ),
    .A_N(\pwm_module.counter1[11] ));
 sg13g2_o21ai_1 _4278_ (.B1(_1696_),
    .Y(_1697_),
    .A1(\pwm_module.counter1[10] ),
    .A2(_1904_));
 sg13g2_nor3_1 _4279_ (.A(_1694_),
    .B(_1695_),
    .C(_1697_),
    .Y(_1698_));
 sg13g2_a22oi_1 _4280_ (.Y(_1699_),
    .B1(_1908_),
    .B2(\pwm_module.counter1[8] ),
    .A2(_1906_),
    .A1(\pwm_module.counter1[9] ));
 sg13g2_a22oi_1 _4281_ (.Y(_1700_),
    .B1(\MemCell.counter_value[7] ),
    .B2(_1798_),
    .A2(\MemCell.counter_value[8] ),
    .A1(_1797_));
 sg13g2_nand4_1 _4282_ (.B(_1698_),
    .C(_1699_),
    .A(_1692_),
    .Y(_1701_),
    .D(_1700_));
 sg13g2_a21oi_2 _4283_ (.B1(_1701_),
    .Y(_1702_),
    .A2(_1682_),
    .A1(_1681_));
 sg13g2_and2_1 _4284_ (.A(_1694_),
    .B(_1696_),
    .X(_1703_));
 sg13g2_nor4_1 _4285_ (.A(_1694_),
    .B(_1695_),
    .C(_1697_),
    .D(_1699_),
    .Y(_1704_));
 sg13g2_o21ai_1 _4286_ (.B1(_1692_),
    .Y(_1705_),
    .A1(_1703_),
    .A2(_1704_));
 sg13g2_nand2_1 _4287_ (.Y(_1706_),
    .A(_1684_),
    .B(_1685_));
 sg13g2_nand3_1 _4288_ (.B(_1689_),
    .C(_1690_),
    .A(_1687_),
    .Y(_1707_));
 sg13g2_nand3_1 _4289_ (.B(_1706_),
    .C(_1707_),
    .A(_1705_),
    .Y(_1708_));
 sg13g2_nor2_1 _4290_ (.A(\pwm_module.counter1[16] ),
    .B(_1897_),
    .Y(_1709_));
 sg13g2_nor4_1 _4291_ (.A(_1663_),
    .B(_1666_),
    .C(_1667_),
    .D(_1709_),
    .Y(_1710_));
 sg13g2_nand3_1 _4292_ (.B(_1665_),
    .C(_1710_),
    .A(_1664_),
    .Y(_1711_));
 sg13g2_nor4_2 _4293_ (.A(_1644_),
    .B(_1649_),
    .C(_1661_),
    .Y(_1712_),
    .D(_1711_));
 sg13g2_o21ai_1 _4294_ (.B1(_1712_),
    .Y(_1713_),
    .A1(_1702_),
    .A2(_1708_));
 sg13g2_a21oi_2 _4295_ (.B1(_1659_),
    .Y(_1714_),
    .A2(_1669_),
    .A1(_1662_));
 sg13g2_nand2_1 _4296_ (.Y(_1715_),
    .A(_1713_),
    .B(_1714_));
 sg13g2_a22oi_1 _4297_ (.Y(_1716_),
    .B1(_1713_),
    .B2(_1714_),
    .A2(_0790_),
    .A1(net646));
 sg13g2_nand2_2 _4298_ (.Y(_1717_),
    .A(net574),
    .B(_1715_));
 sg13g2_xnor2_1 _4299_ (.Y(_1718_),
    .A(net421),
    .B(net572));
 sg13g2_nor2_1 _4300_ (.A(net569),
    .B(_1718_),
    .Y(_0359_));
 sg13g2_a21o_1 _4301_ (.A2(net572),
    .A1(net421),
    .B1(net541),
    .X(_1719_));
 sg13g2_nand3_1 _4302_ (.B(net528),
    .C(net572),
    .A(net541),
    .Y(_1720_));
 sg13g2_and3_1 _4303_ (.X(_0360_),
    .A(net567),
    .B(_1719_),
    .C(_1720_));
 sg13g2_and3_1 _4304_ (.X(_1721_),
    .A(net188),
    .B(\pwm_module.counter1[1] ),
    .C(\pwm_module.counter1[0] ));
 sg13g2_a21o_1 _4305_ (.A2(_1721_),
    .A1(net572),
    .B1(net569),
    .X(_1722_));
 sg13g2_a21oi_1 _4306_ (.A1(_1804_),
    .A2(_1720_),
    .Y(_0361_),
    .B1(_1722_));
 sg13g2_a21o_1 _4307_ (.A2(_1721_),
    .A1(net572),
    .B1(net417),
    .X(_1723_));
 sg13g2_nand3_1 _4308_ (.B(net572),
    .C(_1721_),
    .A(net417),
    .Y(_1724_));
 sg13g2_and3_1 _4309_ (.X(_0362_),
    .A(net567),
    .B(_1723_),
    .C(_1724_));
 sg13g2_and3_2 _4310_ (.X(_1725_),
    .A(\pwm_module.counter1[4] ),
    .B(\pwm_module.counter1[3] ),
    .C(_1721_));
 sg13g2_inv_1 _4311_ (.Y(_1726_),
    .A(_1725_));
 sg13g2_a21oi_2 _4312_ (.B1(_1726_),
    .Y(_1727_),
    .A2(_0790_),
    .A1(net644));
 sg13g2_a221oi_1 _4313_ (.B2(net572),
    .C1(net569),
    .B1(_1725_),
    .A1(_1801_),
    .Y(_0363_),
    .A2(_1724_));
 sg13g2_xnor2_1 _4314_ (.Y(_1728_),
    .A(net79),
    .B(_1727_));
 sg13g2_nor2_1 _4315_ (.A(net569),
    .B(_1728_),
    .Y(_0364_));
 sg13g2_a21o_1 _4316_ (.A2(_1727_),
    .A1(net647),
    .B1(net543),
    .X(_1729_));
 sg13g2_nand3_1 _4317_ (.B(net647),
    .C(_1727_),
    .A(net543),
    .Y(_1730_));
 sg13g2_and3_1 _4318_ (.X(_0365_),
    .A(net567),
    .B(_1729_),
    .C(_1730_));
 sg13g2_and3_1 _4319_ (.X(_1731_),
    .A(net485),
    .B(\pwm_module.counter1[6] ),
    .C(net647));
 sg13g2_and4_1 _4320_ (.A(\pwm_module.counter1[7] ),
    .B(\pwm_module.counter1[6] ),
    .C(net647),
    .D(_1725_),
    .X(_1732_));
 sg13g2_inv_1 _4321_ (.Y(_1733_),
    .A(_1732_));
 sg13g2_a21oi_2 _4322_ (.B1(_1733_),
    .Y(_1734_),
    .A2(_0790_),
    .A1(net644));
 sg13g2_a221oi_1 _4323_ (.B2(_1727_),
    .C1(net569),
    .B1(_1731_),
    .A1(_1798_),
    .Y(_0366_),
    .A2(_1730_));
 sg13g2_or2_1 _4324_ (.X(_1735_),
    .B(_1734_),
    .A(net522));
 sg13g2_nand2_1 _4325_ (.Y(_1736_),
    .A(net522),
    .B(_1734_));
 sg13g2_and3_1 _4326_ (.X(_0367_),
    .A(net567),
    .B(_1735_),
    .C(_1736_));
 sg13g2_a21o_1 _4327_ (.A2(_1734_),
    .A1(net522),
    .B1(net414),
    .X(_1737_));
 sg13g2_nand3_1 _4328_ (.B(\pwm_module.counter1[8] ),
    .C(_1734_),
    .A(net414),
    .Y(_1738_));
 sg13g2_and3_1 _4329_ (.X(_0368_),
    .A(net567),
    .B(_1737_),
    .C(net415));
 sg13g2_nor3_2 _4330_ (.A(_1793_),
    .B(_1795_),
    .C(_1797_),
    .Y(_1739_));
 sg13g2_a221oi_1 _4331_ (.B2(_1734_),
    .C1(net571),
    .B1(_1739_),
    .A1(_1793_),
    .Y(_0369_),
    .A2(net415));
 sg13g2_a21oi_1 _4332_ (.A1(_1734_),
    .A2(_1739_),
    .Y(_1740_),
    .B1(net279));
 sg13g2_nand4_1 _4333_ (.B(_1725_),
    .C(_1731_),
    .A(net279),
    .Y(_1741_),
    .D(_1739_));
 sg13g2_a21oi_2 _4334_ (.B1(_1741_),
    .Y(_1742_),
    .A2(_0790_),
    .A1(net645));
 sg13g2_nor3_1 _4335_ (.A(net569),
    .B(_1740_),
    .C(_1742_),
    .Y(_0370_));
 sg13g2_nor2_1 _4336_ (.A(net397),
    .B(_1742_),
    .Y(_1743_));
 sg13g2_a221oi_1 _4337_ (.B2(net397),
    .C1(_1743_),
    .B1(_1742_),
    .A1(net572),
    .Y(_0371_),
    .A2(_1715_));
 sg13g2_a21o_1 _4338_ (.A2(_1742_),
    .A1(net397),
    .B1(net539),
    .X(_1744_));
 sg13g2_nand3_1 _4339_ (.B(\pwm_module.counter1[12] ),
    .C(_1742_),
    .A(net539),
    .Y(_1745_));
 sg13g2_and3_1 _4340_ (.X(_0372_),
    .A(net567),
    .B(_1744_),
    .C(_1745_));
 sg13g2_and3_1 _4341_ (.X(_1746_),
    .A(net391),
    .B(net557),
    .C(\pwm_module.counter1[12] ));
 sg13g2_nand4_1 _4342_ (.B(_1732_),
    .C(_1739_),
    .A(\pwm_module.counter1[11] ),
    .Y(_1747_),
    .D(_1746_));
 sg13g2_nand2_1 _4343_ (.Y(_1748_),
    .A(_1742_),
    .B(_1746_));
 sg13g2_a221oi_1 _4344_ (.B2(_1742_),
    .C1(net569),
    .B1(_1746_),
    .A1(_1788_),
    .Y(_0373_),
    .A2(_1745_));
 sg13g2_nor2_2 _4345_ (.A(_1786_),
    .B(_1747_),
    .Y(_1749_));
 sg13g2_nand2_1 _4346_ (.Y(_1750_),
    .A(net574),
    .B(_1749_));
 sg13g2_a221oi_1 _4347_ (.B2(net576),
    .C1(net569),
    .B1(_1749_),
    .A1(_1786_),
    .Y(_0374_),
    .A2(_1748_));
 sg13g2_and2_1 _4348_ (.A(net490),
    .B(_1749_),
    .X(_1751_));
 sg13g2_nand2_1 _4349_ (.Y(_1752_),
    .A(net574),
    .B(_1751_));
 sg13g2_a221oi_1 _4350_ (.B2(net574),
    .C1(net570),
    .B1(_1751_),
    .A1(_1785_),
    .Y(_0375_),
    .A2(_1750_));
 sg13g2_and2_1 _4351_ (.A(net459),
    .B(_1751_),
    .X(_1753_));
 sg13g2_a221oi_1 _4352_ (.B2(net574),
    .C1(net570),
    .B1(_1753_),
    .A1(_1925_),
    .Y(_0376_),
    .A2(_1752_));
 sg13g2_a21o_1 _4353_ (.A2(_1753_),
    .A1(net574),
    .B1(net545),
    .X(_1754_));
 sg13g2_nand3_1 _4354_ (.B(net574),
    .C(_1753_),
    .A(\pwm_module.counter1[18] ),
    .Y(_1755_));
 sg13g2_and3_1 _4355_ (.X(_0377_),
    .A(_1717_),
    .B(_1754_),
    .C(_1755_));
 sg13g2_nand4_1 _4356_ (.B(\pwm_module.counter1[19] ),
    .C(\pwm_module.counter1[18] ),
    .A(\pwm_module.counter1[16] ),
    .Y(_1756_),
    .D(\pwm_module.counter1[17] ));
 sg13g2_inv_1 _4357_ (.Y(_1757_),
    .A(_1756_));
 sg13g2_and2_1 _4358_ (.A(_1749_),
    .B(_1757_),
    .X(_1758_));
 sg13g2_nand2_1 _4359_ (.Y(_1759_),
    .A(net573),
    .B(_1758_));
 sg13g2_a221oi_1 _4360_ (.B2(net574),
    .C1(net570),
    .B1(_1758_),
    .A1(_1924_),
    .Y(_0378_),
    .A2(_1755_));
 sg13g2_and2_1 _4361_ (.A(net514),
    .B(_1758_),
    .X(_1760_));
 sg13g2_a221oi_1 _4362_ (.B2(net573),
    .C1(net571),
    .B1(_1760_),
    .A1(_1923_),
    .Y(_0379_),
    .A2(_1759_));
 sg13g2_a21o_1 _4363_ (.A2(_1760_),
    .A1(net573),
    .B1(net537),
    .X(_1761_));
 sg13g2_nand3_1 _4364_ (.B(net573),
    .C(_1760_),
    .A(net537),
    .Y(_1762_));
 sg13g2_and3_1 _4365_ (.X(_0380_),
    .A(_1717_),
    .B(_1761_),
    .C(_1762_));
 sg13g2_nor3_1 _4366_ (.A(_1921_),
    .B(_1922_),
    .C(_1923_),
    .Y(_1763_));
 sg13g2_and2_1 _4367_ (.A(_1758_),
    .B(_1763_),
    .X(_1764_));
 sg13g2_nand2_1 _4368_ (.Y(_1765_),
    .A(net573),
    .B(_1764_));
 sg13g2_a21o_1 _4369_ (.A2(_1764_),
    .A1(net573),
    .B1(net571),
    .X(_1766_));
 sg13g2_a21oi_1 _4370_ (.A1(_1921_),
    .A2(_1762_),
    .Y(_0381_),
    .B1(_1766_));
 sg13g2_nand3_1 _4371_ (.B(_1713_),
    .C(_1714_),
    .A(_1920_),
    .Y(_1767_));
 sg13g2_a22oi_1 _4372_ (.Y(_0382_),
    .B1(_1766_),
    .B2(_1767_),
    .A2(_1765_),
    .A1(_1920_));
 sg13g2_nand4_1 _4373_ (.B(_1749_),
    .C(_1757_),
    .A(\pwm_module.counter1[23] ),
    .Y(_1768_),
    .D(_1763_));
 sg13g2_a21oi_2 _4374_ (.B1(_1768_),
    .Y(_1769_),
    .A2(_0790_),
    .A1(net646));
 sg13g2_xnor2_1 _4375_ (.Y(_1770_),
    .A(net525),
    .B(_1769_));
 sg13g2_nor2_1 _4376_ (.A(net570),
    .B(_1770_),
    .Y(_0383_));
 sg13g2_a21oi_1 _4377_ (.A1(\pwm_module.counter1[24] ),
    .A2(_1769_),
    .Y(_1771_),
    .B1(net254));
 sg13g2_and2_1 _4378_ (.A(\pwm_module.counter1[25] ),
    .B(\pwm_module.counter1[24] ),
    .X(_1772_));
 sg13g2_a21oi_1 _4379_ (.A1(_1769_),
    .A2(_1772_),
    .Y(_1773_),
    .B1(net570));
 sg13g2_nor2b_1 _4380_ (.A(net255),
    .B_N(_1773_),
    .Y(_0384_));
 sg13g2_a21o_1 _4381_ (.A2(_1772_),
    .A1(_1769_),
    .B1(net549),
    .X(_1774_));
 sg13g2_nand3_1 _4382_ (.B(_1769_),
    .C(_1772_),
    .A(\pwm_module.counter1[26] ),
    .Y(_1775_));
 sg13g2_and3_1 _4383_ (.X(_0385_),
    .A(net567),
    .B(_1774_),
    .C(_1775_));
 sg13g2_and3_1 _4384_ (.X(_1776_),
    .A(net515),
    .B(\pwm_module.counter1[26] ),
    .C(_1772_));
 sg13g2_a221oi_1 _4385_ (.B2(_1769_),
    .C1(net571),
    .B1(_1776_),
    .A1(_1919_),
    .Y(_0386_),
    .A2(_1775_));
 sg13g2_a21oi_1 _4386_ (.A1(_1769_),
    .A2(_1776_),
    .Y(_1777_),
    .B1(net356));
 sg13g2_nand2_1 _4387_ (.Y(_1778_),
    .A(\pwm_module.counter1[28] ),
    .B(_1776_));
 sg13g2_nor2_2 _4388_ (.A(_1768_),
    .B(_1778_),
    .Y(_1779_));
 sg13g2_a21oi_1 _4389_ (.A1(net575),
    .A2(_1779_),
    .Y(_1780_),
    .B1(net570));
 sg13g2_nor2b_1 _4390_ (.A(net357),
    .B_N(_1780_),
    .Y(_0387_));
 sg13g2_a21o_1 _4391_ (.A2(_1779_),
    .A1(net575),
    .B1(net547),
    .X(_1781_));
 sg13g2_nand3_1 _4392_ (.B(net575),
    .C(_1779_),
    .A(\pwm_module.counter1[29] ),
    .Y(_1782_));
 sg13g2_and3_1 _4393_ (.X(_0388_),
    .A(net567),
    .B(_1781_),
    .C(_1782_));
 sg13g2_and3_1 _4394_ (.X(_1783_),
    .A(net500),
    .B(\pwm_module.counter1[29] ),
    .C(_1779_));
 sg13g2_nand4_1 _4395_ (.B(\pwm_module.counter1[29] ),
    .C(net573),
    .A(\pwm_module.counter1[30] ),
    .Y(_1784_),
    .D(_1779_));
 sg13g2_a221oi_1 _4396_ (.B2(net573),
    .C1(net570),
    .B1(_1783_),
    .A1(_1918_),
    .Y(_0389_),
    .A2(_1782_));
 sg13g2_a21oi_1 _4397_ (.A1(_1917_),
    .A2(_1784_),
    .Y(_0390_),
    .B1(net570));
 sg13g2_inv_1 _4398_ (.Y(_0105_),
    .A(net683));
 sg13g2_inv_1 _4399_ (.Y(_0106_),
    .A(net683));
 sg13g2_inv_1 _4400_ (.Y(_0107_),
    .A(net682));
 sg13g2_dfrbp_1 _4401_ (.CLK(net685),
    .RESET_B(_0104_),
    .D(_1998_),
    .Q_N(_1998_),
    .Q(\spi_module.r_RX_Bit_Count[0] ));
 sg13g2_dfrbp_1 _4402_ (.CLK(net685),
    .RESET_B(_0105_),
    .D(_0100_),
    .Q_N(_2281_),
    .Q(\spi_module.r_RX_Bit_Count[1] ));
 sg13g2_dfrbp_1 _4403_ (.CLK(net685),
    .RESET_B(_0106_),
    .D(_0101_),
    .Q_N(_2280_),
    .Q(\spi_module.r_RX_Bit_Count[2] ));
 sg13g2_dfrbp_1 _4404_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net692),
    .D(_0108_),
    .Q_N(_2279_),
    .Q(\pwm_module.counter0[0] ));
 sg13g2_dfrbp_1 _4405_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net692),
    .D(_0109_),
    .Q_N(_2278_),
    .Q(\pwm_module.counter0[1] ));
 sg13g2_dfrbp_1 _4406_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net692),
    .D(net216),
    .Q_N(_2277_),
    .Q(\pwm_module.counter0[2] ));
 sg13g2_dfrbp_1 _4407_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net694),
    .D(_0111_),
    .Q_N(_2276_),
    .Q(\pwm_module.counter0[3] ));
 sg13g2_dfrbp_1 _4408_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net694),
    .D(net466),
    .Q_N(_2275_),
    .Q(\pwm_module.counter0[4] ));
 sg13g2_dfrbp_1 _4409_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net693),
    .D(_0113_),
    .Q_N(_2274_),
    .Q(\pwm_module.counter0[5] ));
 sg13g2_dfrbp_1 _4410_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net694),
    .D(_0114_),
    .Q_N(_2273_),
    .Q(\pwm_module.counter0[6] ));
 sg13g2_dfrbp_1 _4411_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net693),
    .D(net395),
    .Q_N(_2272_),
    .Q(\pwm_module.counter0[7] ));
 sg13g2_dfrbp_1 _4412_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net705),
    .D(_0116_),
    .Q_N(_2271_),
    .Q(\pwm_module.counter0[8] ));
 sg13g2_dfrbp_1 _4413_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net693),
    .D(net289),
    .Q_N(_2270_),
    .Q(\pwm_module.counter0[9] ));
 sg13g2_dfrbp_1 _4414_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net712),
    .D(_0118_),
    .Q_N(_2269_),
    .Q(\pwm_module.counter0[10] ));
 sg13g2_dfrbp_1 _4415_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net699),
    .D(_0119_),
    .Q_N(_2268_),
    .Q(\pwm_module.counter0[11] ));
 sg13g2_dfrbp_1 _4416_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net701),
    .D(_0120_),
    .Q_N(_2267_),
    .Q(\pwm_module.counter0[12] ));
 sg13g2_dfrbp_1 _4417_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net699),
    .D(net423),
    .Q_N(_2266_),
    .Q(\pwm_module.counter0[13] ));
 sg13g2_dfrbp_1 _4418_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net699),
    .D(_0122_),
    .Q_N(_2265_),
    .Q(\pwm_module.counter0[14] ));
 sg13g2_dfrbp_1 _4419_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net701),
    .D(_0123_),
    .Q_N(_2264_),
    .Q(\pwm_module.counter0[15] ));
 sg13g2_dfrbp_1 _4420_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net725),
    .D(_0124_),
    .Q_N(_2263_),
    .Q(\pwm_module.counter0[16] ));
 sg13g2_dfrbp_1 _4421_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net725),
    .D(_0125_),
    .Q_N(_2262_),
    .Q(\pwm_module.counter0[17] ));
 sg13g2_dfrbp_1 _4422_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net725),
    .D(net454),
    .Q_N(_2261_),
    .Q(\pwm_module.counter0[18] ));
 sg13g2_dfrbp_1 _4423_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net725),
    .D(net399),
    .Q_N(_2260_),
    .Q(\pwm_module.counter0[19] ));
 sg13g2_dfrbp_1 _4424_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net727),
    .D(net484),
    .Q_N(_2259_),
    .Q(\pwm_module.counter0[20] ));
 sg13g2_dfrbp_1 _4425_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net726),
    .D(_0129_),
    .Q_N(_2258_),
    .Q(\pwm_module.counter0[21] ));
 sg13g2_dfrbp_1 _4426_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net726),
    .D(net374),
    .Q_N(_2257_),
    .Q(\pwm_module.counter0[22] ));
 sg13g2_dfrbp_1 _4427_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net724),
    .D(_0131_),
    .Q_N(_2256_),
    .Q(\pwm_module.counter0[23] ));
 sg13g2_dfrbp_1 _4428_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net731),
    .D(_0132_),
    .Q_N(_2255_),
    .Q(\pwm_module.counter0[24] ));
 sg13g2_dfrbp_1 _4429_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net731),
    .D(_0133_),
    .Q_N(_2254_),
    .Q(\pwm_module.counter0[25] ));
 sg13g2_dfrbp_1 _4430_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net731),
    .D(net343),
    .Q_N(_2253_),
    .Q(\pwm_module.counter0[26] ));
 sg13g2_dfrbp_1 _4431_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net726),
    .D(_0135_),
    .Q_N(_2252_),
    .Q(\pwm_module.counter0[27] ));
 sg13g2_dfrbp_1 _4432_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net738),
    .D(net472),
    .Q_N(_2251_),
    .Q(\pwm_module.counter0[28] ));
 sg13g2_dfrbp_1 _4433_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net738),
    .D(_0137_),
    .Q_N(_2250_),
    .Q(\pwm_module.counter0[29] ));
 sg13g2_dfrbp_1 _4434_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net738),
    .D(net291),
    .Q_N(_2249_),
    .Q(\pwm_module.counter0[30] ));
 sg13g2_dfrbp_1 _4435_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net745),
    .D(_0139_),
    .Q_N(_2282_),
    .Q(\pwm_module.counter0[31] ));
 sg13g2_dfrbp_1 _4436_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net751),
    .D(net38),
    .Q_N(_2283_),
    .Q(\spi_module.r3_RX_Done ));
 sg13g2_dfrbp_1 _4437_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net745),
    .D(net643),
    .Q_N(_2248_),
    .Q(\MemCell.o_RX_DV ));
 sg13g2_dfrbp_1 _4438_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net747),
    .D(_0140_),
    .Q_N(_2247_),
    .Q(\MemCell.o_RX_Byte[0] ));
 sg13g2_dfrbp_1 _4439_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net747),
    .D(_0141_),
    .Q_N(_2246_),
    .Q(\MemCell.o_RX_Byte[1] ));
 sg13g2_dfrbp_1 _4440_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net747),
    .D(_0142_),
    .Q_N(_2245_),
    .Q(\MemCell.o_RX_Byte[2] ));
 sg13g2_dfrbp_1 _4441_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net747),
    .D(_0143_),
    .Q_N(_2244_),
    .Q(\MemCell.o_RX_Byte[3] ));
 sg13g2_dfrbp_1 _4442_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net750),
    .D(_0144_),
    .Q_N(_2243_),
    .Q(\MemCell.o_RX_Byte[4] ));
 sg13g2_dfrbp_1 _4443_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net750),
    .D(net437),
    .Q_N(_2242_),
    .Q(\MemCell.o_RX_Byte[5] ));
 sg13g2_dfrbp_1 _4444_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net750),
    .D(_0146_),
    .Q_N(_2241_),
    .Q(\MemCell.o_RX_Byte[6] ));
 sg13g2_dfrbp_1 _4445_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net750),
    .D(_0147_),
    .Q_N(_2240_),
    .Q(\MemCell.o_RX_Byte[7] ));
 sg13g2_dfrbp_1 _4446_ (.CLK(net684),
    .RESET_B(net31),
    .D(_0148_),
    .Q_N(_2239_),
    .Q(\spi_module.r_Temp_RX_Byte[0] ));
 sg13g2_dfrbp_1 _4447_ (.CLK(net684),
    .RESET_B(net30),
    .D(_0149_),
    .Q_N(_2238_),
    .Q(\spi_module.r_Temp_RX_Byte[1] ));
 sg13g2_dfrbp_1 _4448_ (.CLK(net684),
    .RESET_B(net29),
    .D(_0150_),
    .Q_N(_2237_),
    .Q(\spi_module.r_Temp_RX_Byte[2] ));
 sg13g2_dfrbp_1 _4449_ (.CLK(net684),
    .RESET_B(net28),
    .D(_0151_),
    .Q_N(_2236_),
    .Q(\spi_module.r_Temp_RX_Byte[3] ));
 sg13g2_dfrbp_1 _4450_ (.CLK(net684),
    .RESET_B(net27),
    .D(_0152_),
    .Q_N(_2235_),
    .Q(\spi_module.r_Temp_RX_Byte[4] ));
 sg13g2_dfrbp_1 _4451_ (.CLK(net685),
    .RESET_B(net26),
    .D(_0153_),
    .Q_N(_2234_),
    .Q(\spi_module.r_Temp_RX_Byte[5] ));
 sg13g2_dfrbp_1 _4452_ (.CLK(net686),
    .RESET_B(net32),
    .D(_0154_),
    .Q_N(_2284_),
    .Q(\spi_module.r_Temp_RX_Byte[6] ));
 sg13g2_dfrbp_1 _4453_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net750),
    .D(\spi_module.r_RX_Done ),
    .Q_N(_2233_),
    .Q(\spi_module.r2_RX_Done ));
 sg13g2_dfrbp_1 _4454_ (.CLK(net684),
    .RESET_B(net25),
    .D(_0155_),
    .Q_N(_2232_),
    .Q(\spi_module.r_RX_Byte[0] ));
 sg13g2_dfrbp_1 _4455_ (.CLK(net684),
    .RESET_B(net24),
    .D(_0156_),
    .Q_N(_2231_),
    .Q(\spi_module.r_RX_Byte[1] ));
 sg13g2_dfrbp_1 _4456_ (.CLK(net684),
    .RESET_B(net23),
    .D(_0157_),
    .Q_N(_2230_),
    .Q(\spi_module.r_RX_Byte[2] ));
 sg13g2_dfrbp_1 _4457_ (.CLK(net686),
    .RESET_B(net22),
    .D(_0158_),
    .Q_N(_2229_),
    .Q(\spi_module.r_RX_Byte[3] ));
 sg13g2_dfrbp_1 _4458_ (.CLK(net686),
    .RESET_B(net21),
    .D(_0159_),
    .Q_N(_2228_),
    .Q(\spi_module.r_RX_Byte[4] ));
 sg13g2_dfrbp_1 _4459_ (.CLK(net685),
    .RESET_B(net20),
    .D(_0160_),
    .Q_N(_2227_),
    .Q(\spi_module.r_RX_Byte[5] ));
 sg13g2_dfrbp_1 _4460_ (.CLK(net685),
    .RESET_B(net19),
    .D(_0161_),
    .Q_N(_2226_),
    .Q(\spi_module.r_RX_Byte[6] ));
 sg13g2_dfrbp_1 _4461_ (.CLK(net685),
    .RESET_B(net18),
    .D(_0162_),
    .Q_N(_2225_),
    .Q(\spi_module.r_RX_Byte[7] ));
 sg13g2_dfrbp_1 _4462_ (.CLK(net685),
    .RESET_B(_0107_),
    .D(_0163_),
    .Q_N(_2224_),
    .Q(\spi_module.r_RX_Done ));
 sg13g2_dfrbp_1 _4463_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net728),
    .D(_0164_),
    .Q_N(_2223_),
    .Q(\MemCell.dc2_reg[3][0] ));
 sg13g2_dfrbp_1 _4464_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net728),
    .D(_0165_),
    .Q_N(_2222_),
    .Q(\MemCell.dc2_reg[3][1] ));
 sg13g2_dfrbp_1 _4465_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net728),
    .D(_0166_),
    .Q_N(_2221_),
    .Q(\MemCell.dc2_reg[3][2] ));
 sg13g2_dfrbp_1 _4466_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net728),
    .D(_0167_),
    .Q_N(_2220_),
    .Q(\MemCell.dc2_reg[3][3] ));
 sg13g2_dfrbp_1 _4467_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net728),
    .D(_0168_),
    .Q_N(_2219_),
    .Q(\MemCell.dc2_reg[3][4] ));
 sg13g2_dfrbp_1 _4468_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net729),
    .D(_0169_),
    .Q_N(_2218_),
    .Q(\MemCell.dc2_reg[3][5] ));
 sg13g2_dfrbp_1 _4469_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net728),
    .D(_0170_),
    .Q_N(_2217_),
    .Q(\MemCell.dc2_reg[3][6] ));
 sg13g2_dfrbp_1 _4470_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net728),
    .D(_0171_),
    .Q_N(_2216_),
    .Q(\MemCell.dc2_reg[3][7] ));
 sg13g2_dfrbp_1 _4471_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net730),
    .D(_0172_),
    .Q_N(_2215_),
    .Q(\MemCell.dc3_reg[2][0] ));
 sg13g2_dfrbp_1 _4472_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net730),
    .D(_0173_),
    .Q_N(_2214_),
    .Q(\MemCell.dc3_reg[2][1] ));
 sg13g2_dfrbp_1 _4473_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net730),
    .D(_0174_),
    .Q_N(_2213_),
    .Q(\MemCell.dc3_reg[2][2] ));
 sg13g2_dfrbp_1 _4474_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net730),
    .D(_0175_),
    .Q_N(_2212_),
    .Q(\MemCell.dc3_reg[2][3] ));
 sg13g2_dfrbp_1 _4475_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net730),
    .D(_0176_),
    .Q_N(_2211_),
    .Q(\MemCell.dc3_reg[2][4] ));
 sg13g2_dfrbp_1 _4476_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net730),
    .D(_0177_),
    .Q_N(_2210_),
    .Q(\MemCell.dc3_reg[2][5] ));
 sg13g2_dfrbp_1 _4477_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net729),
    .D(_0178_),
    .Q_N(_2209_),
    .Q(\MemCell.dc3_reg[2][6] ));
 sg13g2_dfrbp_1 _4478_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net730),
    .D(_0179_),
    .Q_N(_2208_),
    .Q(\MemCell.dc3_reg[2][7] ));
 sg13g2_dfrbp_1 _4479_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net720),
    .D(_0180_),
    .Q_N(_2207_),
    .Q(\MemCell.dc2_reg[2][0] ));
 sg13g2_dfrbp_1 _4480_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net720),
    .D(_0181_),
    .Q_N(_2206_),
    .Q(\MemCell.dc2_reg[2][1] ));
 sg13g2_dfrbp_1 _4481_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net720),
    .D(_0182_),
    .Q_N(_2205_),
    .Q(\MemCell.dc2_reg[2][2] ));
 sg13g2_dfrbp_1 _4482_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net720),
    .D(_0183_),
    .Q_N(_2204_),
    .Q(\MemCell.dc2_reg[2][3] ));
 sg13g2_dfrbp_1 _4483_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net721),
    .D(_0184_),
    .Q_N(_2203_),
    .Q(\MemCell.dc2_reg[2][4] ));
 sg13g2_dfrbp_1 _4484_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net721),
    .D(_0185_),
    .Q_N(_2202_),
    .Q(\MemCell.dc2_reg[2][5] ));
 sg13g2_dfrbp_1 _4485_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net721),
    .D(_0186_),
    .Q_N(_2201_),
    .Q(\MemCell.dc2_reg[2][6] ));
 sg13g2_dfrbp_1 _4486_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net721),
    .D(_0187_),
    .Q_N(_2200_),
    .Q(\MemCell.dc2_reg[2][7] ));
 sg13g2_dfrbp_1 _4487_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net689),
    .D(net142),
    .Q_N(_2199_),
    .Q(\MemCell.dc2_reg[1][0] ));
 sg13g2_dfrbp_1 _4488_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net695),
    .D(_0189_),
    .Q_N(_2198_),
    .Q(\MemCell.dc2_reg[1][1] ));
 sg13g2_dfrbp_1 _4489_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net695),
    .D(_0190_),
    .Q_N(_2197_),
    .Q(\MemCell.dc2_reg[1][2] ));
 sg13g2_dfrbp_1 _4490_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net695),
    .D(_0191_),
    .Q_N(_2196_),
    .Q(\MemCell.dc2_reg[1][3] ));
 sg13g2_dfrbp_1 _4491_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net697),
    .D(_0192_),
    .Q_N(_2195_),
    .Q(\MemCell.dc2_reg[1][4] ));
 sg13g2_dfrbp_1 _4492_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net697),
    .D(_0193_),
    .Q_N(_2194_),
    .Q(\MemCell.dc2_reg[1][5] ));
 sg13g2_dfrbp_1 _4493_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net697),
    .D(_0194_),
    .Q_N(_2193_),
    .Q(\MemCell.dc2_reg[1][6] ));
 sg13g2_dfrbp_1 _4494_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net698),
    .D(_0195_),
    .Q_N(_2192_),
    .Q(\MemCell.dc2_reg[1][7] ));
 sg13g2_dfrbp_1 _4495_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net687),
    .D(_0196_),
    .Q_N(_2191_),
    .Q(\MemCell.dc2_reg[0][0] ));
 sg13g2_dfrbp_1 _4496_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net687),
    .D(_0197_),
    .Q_N(_2190_),
    .Q(\MemCell.dc2_reg[0][1] ));
 sg13g2_dfrbp_1 _4497_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net687),
    .D(_0198_),
    .Q_N(_2189_),
    .Q(\MemCell.dc2_reg[0][2] ));
 sg13g2_dfrbp_1 _4498_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net687),
    .D(_0199_),
    .Q_N(_2188_),
    .Q(\MemCell.dc2_reg[0][3] ));
 sg13g2_dfrbp_1 _4499_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net687),
    .D(_0200_),
    .Q_N(_2187_),
    .Q(\MemCell.dc2_reg[0][4] ));
 sg13g2_dfrbp_1 _4500_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net689),
    .D(_0201_),
    .Q_N(_2186_),
    .Q(\MemCell.dc2_reg[0][5] ));
 sg13g2_dfrbp_1 _4501_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net689),
    .D(_0202_),
    .Q_N(_2185_),
    .Q(\MemCell.dc2_reg[0][6] ));
 sg13g2_dfrbp_1 _4502_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net689),
    .D(_0203_),
    .Q_N(_2184_),
    .Q(\MemCell.dc2_reg[0][7] ));
 sg13g2_dfrbp_1 _4503_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net745),
    .D(net269),
    .Q_N(_2183_),
    .Q(\MemCell.dc1_reg[3][0] ));
 sg13g2_dfrbp_1 _4504_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net745),
    .D(_0205_),
    .Q_N(_2182_),
    .Q(\MemCell.dc1_reg[3][1] ));
 sg13g2_dfrbp_1 _4505_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net745),
    .D(_0206_),
    .Q_N(_2181_),
    .Q(\MemCell.dc1_reg[3][2] ));
 sg13g2_dfrbp_1 _4506_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net745),
    .D(_0207_),
    .Q_N(_2180_),
    .Q(\MemCell.dc1_reg[3][3] ));
 sg13g2_dfrbp_1 _4507_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net738),
    .D(_0208_),
    .Q_N(_2179_),
    .Q(\MemCell.dc1_reg[3][4] ));
 sg13g2_dfrbp_1 _4508_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net738),
    .D(_0209_),
    .Q_N(_2178_),
    .Q(\MemCell.dc1_reg[3][5] ));
 sg13g2_dfrbp_1 _4509_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net745),
    .D(_0210_),
    .Q_N(_2177_),
    .Q(\MemCell.dc1_reg[3][6] ));
 sg13g2_dfrbp_1 _4510_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net745),
    .D(_0211_),
    .Q_N(_2176_),
    .Q(\MemCell.dc1_reg[3][7] ));
 sg13g2_dfrbp_1 _4511_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net736),
    .D(net55),
    .Q_N(_2175_),
    .Q(\MemCell.dc1_reg[2][0] ));
 sg13g2_dfrbp_1 _4512_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net736),
    .D(net159),
    .Q_N(_2174_),
    .Q(\MemCell.dc1_reg[2][1] ));
 sg13g2_dfrbp_1 _4513_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net736),
    .D(net91),
    .Q_N(_2173_),
    .Q(\MemCell.dc1_reg[2][2] ));
 sg13g2_dfrbp_1 _4514_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net724),
    .D(net61),
    .Q_N(_2172_),
    .Q(\MemCell.dc1_reg[2][3] ));
 sg13g2_dfrbp_1 _4515_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net736),
    .D(_0216_),
    .Q_N(_2171_),
    .Q(\MemCell.dc1_reg[2][4] ));
 sg13g2_dfrbp_1 _4516_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net736),
    .D(_0217_),
    .Q_N(_2170_),
    .Q(\MemCell.dc1_reg[2][5] ));
 sg13g2_dfrbp_1 _4517_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net736),
    .D(net145),
    .Q_N(_2169_),
    .Q(\MemCell.dc1_reg[2][6] ));
 sg13g2_dfrbp_1 _4518_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net736),
    .D(_0219_),
    .Q_N(_2168_),
    .Q(\MemCell.dc1_reg[2][7] ));
 sg13g2_dfrbp_1 _4519_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net705),
    .D(_0220_),
    .Q_N(_2167_),
    .Q(\MemCell.dc1_reg[1][0] ));
 sg13g2_dfrbp_1 _4520_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net705),
    .D(_0221_),
    .Q_N(_2166_),
    .Q(\MemCell.dc1_reg[1][1] ));
 sg13g2_dfrbp_1 _4521_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net712),
    .D(_0222_),
    .Q_N(_2165_),
    .Q(\MemCell.dc1_reg[1][2] ));
 sg13g2_dfrbp_1 _4522_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net712),
    .D(_0223_),
    .Q_N(_2164_),
    .Q(\MemCell.dc1_reg[1][3] ));
 sg13g2_dfrbp_1 _4523_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net712),
    .D(net87),
    .Q_N(_2163_),
    .Q(\MemCell.dc1_reg[1][4] ));
 sg13g2_dfrbp_1 _4524_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net712),
    .D(net107),
    .Q_N(_2162_),
    .Q(\MemCell.dc1_reg[1][5] ));
 sg13g2_dfrbp_1 _4525_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net712),
    .D(net178),
    .Q_N(_2161_),
    .Q(\MemCell.dc1_reg[1][6] ));
 sg13g2_dfrbp_1 _4526_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net712),
    .D(_0227_),
    .Q_N(_2160_),
    .Q(\MemCell.dc1_reg[1][7] ));
 sg13g2_dfrbp_1 _4527_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net703),
    .D(net44),
    .Q_N(_2159_),
    .Q(\MemCell.dc1_reg[0][0] ));
 sg13g2_dfrbp_1 _4528_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net703),
    .D(_0229_),
    .Q_N(_2158_),
    .Q(\MemCell.dc1_reg[0][1] ));
 sg13g2_dfrbp_1 _4529_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net703),
    .D(_0230_),
    .Q_N(_2157_),
    .Q(\MemCell.dc1_reg[0][2] ));
 sg13g2_dfrbp_1 _4530_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net703),
    .D(net63),
    .Q_N(_2156_),
    .Q(\MemCell.dc1_reg[0][3] ));
 sg13g2_dfrbp_1 _4531_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net703),
    .D(net152),
    .Q_N(_2155_),
    .Q(\MemCell.dc1_reg[0][4] ));
 sg13g2_dfrbp_1 _4532_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net703),
    .D(net131),
    .Q_N(_2154_),
    .Q(\MemCell.dc1_reg[0][5] ));
 sg13g2_dfrbp_1 _4533_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net705),
    .D(net78),
    .Q_N(_2153_),
    .Q(\MemCell.dc1_reg[0][6] ));
 sg13g2_dfrbp_1 _4534_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net705),
    .D(_0235_),
    .Q_N(_2152_),
    .Q(\MemCell.dc1_reg[0][7] ));
 sg13g2_dfrbp_1 _4535_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net748),
    .D(_0236_),
    .Q_N(_2151_),
    .Q(\MemCell.prescale_reg[3][0] ));
 sg13g2_dfrbp_1 _4536_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net742),
    .D(net448),
    .Q_N(_2150_),
    .Q(\MemCell.prescale_reg[3][1] ));
 sg13g2_dfrbp_1 _4537_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net748),
    .D(net493),
    .Q_N(_2149_),
    .Q(\MemCell.prescale_reg[3][2] ));
 sg13g2_dfrbp_1 _4538_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net742),
    .D(_0239_),
    .Q_N(_2148_),
    .Q(\MemCell.prescale_reg[3][3] ));
 sg13g2_dfrbp_1 _4539_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net739),
    .D(net299),
    .Q_N(_2147_),
    .Q(\MemCell.prescale_reg[3][4] ));
 sg13g2_dfrbp_1 _4540_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net746),
    .D(_0241_),
    .Q_N(_2146_),
    .Q(\MemCell.prescale_reg[3][5] ));
 sg13g2_dfrbp_1 _4541_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net738),
    .D(net365),
    .Q_N(_2145_),
    .Q(\MemCell.prescale_reg[3][6] ));
 sg13g2_dfrbp_1 _4542_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net738),
    .D(_0243_),
    .Q_N(_2144_),
    .Q(\MemCell.prescale_reg[3][7] ));
 sg13g2_dfrbp_1 _4543_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net742),
    .D(net477),
    .Q_N(_2143_),
    .Q(\MemCell.prescale_reg[2][0] ));
 sg13g2_dfrbp_1 _4544_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net740),
    .D(_0245_),
    .Q_N(_2142_),
    .Q(\MemCell.prescale_reg[2][1] ));
 sg13g2_dfrbp_1 _4545_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net743),
    .D(net505),
    .Q_N(_2141_),
    .Q(\MemCell.prescale_reg[2][2] ));
 sg13g2_dfrbp_1 _4546_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net749),
    .D(net113),
    .Q_N(_2140_),
    .Q(\MemCell.prescale_reg[2][3] ));
 sg13g2_dfrbp_1 _4547_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net743),
    .D(net507),
    .Q_N(_2139_),
    .Q(\MemCell.prescale_reg[2][4] ));
 sg13g2_dfrbp_1 _4548_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net743),
    .D(net509),
    .Q_N(_2138_),
    .Q(\MemCell.prescale_reg[2][5] ));
 sg13g2_dfrbp_1 _4549_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net749),
    .D(net521),
    .Q_N(_2137_),
    .Q(\MemCell.prescale_reg[2][6] ));
 sg13g2_dfrbp_1 _4550_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net749),
    .D(net481),
    .Q_N(_2136_),
    .Q(\MemCell.prescale_reg[2][7] ));
 sg13g2_dfrbp_1 _4551_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net693),
    .D(net162),
    .Q_N(_2135_),
    .Q(\MemCell.dc3_reg[1][0] ));
 sg13g2_dfrbp_1 _4552_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net699),
    .D(_0253_),
    .Q_N(_2134_),
    .Q(\MemCell.dc3_reg[1][1] ));
 sg13g2_dfrbp_1 _4553_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net701),
    .D(_0254_),
    .Q_N(_2133_),
    .Q(\MemCell.dc3_reg[1][2] ));
 sg13g2_dfrbp_1 _4554_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net701),
    .D(_0255_),
    .Q_N(_2132_),
    .Q(\MemCell.dc3_reg[1][3] ));
 sg13g2_dfrbp_1 _4555_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net700),
    .D(_0256_),
    .Q_N(_2131_),
    .Q(\MemCell.dc3_reg[1][4] ));
 sg13g2_dfrbp_1 _4556_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net700),
    .D(_0257_),
    .Q_N(_2130_),
    .Q(\MemCell.dc3_reg[1][5] ));
 sg13g2_dfrbp_1 _4557_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net700),
    .D(_0258_),
    .Q_N(_2129_),
    .Q(\MemCell.dc3_reg[1][6] ));
 sg13g2_dfrbp_1 _4558_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net700),
    .D(_0259_),
    .Q_N(_2128_),
    .Q(\MemCell.dc3_reg[1][7] ));
 sg13g2_dfrbp_1 _4559_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net715),
    .D(net346),
    .Q_N(_2127_),
    .Q(\MemCell.prescale_reg[1][0] ));
 sg13g2_dfrbp_1 _4560_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net715),
    .D(_0261_),
    .Q_N(_2126_),
    .Q(\MemCell.prescale_reg[1][1] ));
 sg13g2_dfrbp_1 _4561_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net715),
    .D(_0262_),
    .Q_N(_2125_),
    .Q(\MemCell.prescale_reg[1][2] ));
 sg13g2_dfrbp_1 _4562_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net715),
    .D(_0263_),
    .Q_N(_2124_),
    .Q(\MemCell.prescale_reg[1][3] ));
 sg13g2_dfrbp_1 _4563_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net715),
    .D(_0264_),
    .Q_N(_2123_),
    .Q(\MemCell.prescale_reg[1][4] ));
 sg13g2_dfrbp_1 _4564_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net716),
    .D(_0265_),
    .Q_N(_2122_),
    .Q(\MemCell.prescale_reg[1][5] ));
 sg13g2_dfrbp_1 _4565_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net718),
    .D(_0266_),
    .Q_N(_2121_),
    .Q(\MemCell.prescale_reg[1][6] ));
 sg13g2_dfrbp_1 _4566_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net718),
    .D(_0267_),
    .Q_N(_2120_),
    .Q(\MemCell.prescale_reg[1][7] ));
 sg13g2_dfrbp_1 _4567_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net704),
    .D(_0268_),
    .Q_N(_2119_),
    .Q(\MemCell.prescale_reg[0][0] ));
 sg13g2_dfrbp_1 _4568_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net704),
    .D(_0269_),
    .Q_N(_2118_),
    .Q(\MemCell.prescale_reg[0][1] ));
 sg13g2_dfrbp_1 _4569_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net704),
    .D(_0270_),
    .Q_N(_2117_),
    .Q(\MemCell.prescale_reg[0][2] ));
 sg13g2_dfrbp_1 _4570_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net703),
    .D(net430),
    .Q_N(_2116_),
    .Q(\MemCell.prescale_reg[0][3] ));
 sg13g2_dfrbp_1 _4571_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net709),
    .D(_0272_),
    .Q_N(_2115_),
    .Q(\MemCell.prescale_reg[0][4] ));
 sg13g2_dfrbp_1 _4572_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net710),
    .D(net439),
    .Q_N(_2114_),
    .Q(\MemCell.prescale_reg[0][5] ));
 sg13g2_dfrbp_1 _4573_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net710),
    .D(_0274_),
    .Q_N(_2113_),
    .Q(\MemCell.prescale_reg[0][6] ));
 sg13g2_dfrbp_1 _4574_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net710),
    .D(_0275_),
    .Q_N(_2112_),
    .Q(\MemCell.prescale_reg[0][7] ));
 sg13g2_dfrbp_1 _4575_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net726),
    .D(net410),
    .Q_N(_2111_),
    .Q(\MemCell.counter_value[24] ));
 sg13g2_dfrbp_1 _4576_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net731),
    .D(net444),
    .Q_N(_2110_),
    .Q(\MemCell.counter_value[25] ));
 sg13g2_dfrbp_1 _4577_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net726),
    .D(_0278_),
    .Q_N(_2109_),
    .Q(\MemCell.counter_value[26] ));
 sg13g2_dfrbp_1 _4578_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net726),
    .D(_0279_),
    .Q_N(_2108_),
    .Q(\MemCell.counter_value[27] ));
 sg13g2_dfrbp_1 _4579_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net731),
    .D(_0280_),
    .Q_N(_2107_),
    .Q(\MemCell.counter_value[28] ));
 sg13g2_dfrbp_1 _4580_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net732),
    .D(_0281_),
    .Q_N(_2106_),
    .Q(\MemCell.counter_value[29] ));
 sg13g2_dfrbp_1 _4581_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net731),
    .D(_0282_),
    .Q_N(_2105_),
    .Q(\MemCell.counter_value[30] ));
 sg13g2_dfrbp_1 _4582_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net731),
    .D(_0283_),
    .Q_N(_2104_),
    .Q(\MemCell.counter_value[31] ));
 sg13g2_dfrbp_1 _4583_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net724),
    .D(net458),
    .Q_N(_2103_),
    .Q(\MemCell.counter_value[16] ));
 sg13g2_dfrbp_1 _4584_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net724),
    .D(_0285_),
    .Q_N(_2102_),
    .Q(\MemCell.counter_value[17] ));
 sg13g2_dfrbp_1 _4585_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net724),
    .D(_0286_),
    .Q_N(_2101_),
    .Q(\MemCell.counter_value[18] ));
 sg13g2_dfrbp_1 _4586_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net724),
    .D(_0287_),
    .Q_N(_2100_),
    .Q(\MemCell.counter_value[19] ));
 sg13g2_dfrbp_1 _4587_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net724),
    .D(_0288_),
    .Q_N(_2099_),
    .Q(\MemCell.counter_value[20] ));
 sg13g2_dfrbp_1 _4588_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net721),
    .D(_0289_),
    .Q_N(_2098_),
    .Q(\MemCell.counter_value[21] ));
 sg13g2_dfrbp_1 _4589_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net724),
    .D(_0290_),
    .Q_N(_2097_),
    .Q(\MemCell.counter_value[22] ));
 sg13g2_dfrbp_1 _4590_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net727),
    .D(_0291_),
    .Q_N(_2096_),
    .Q(\MemCell.counter_value[23] ));
 sg13g2_dfrbp_1 _4591_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net696),
    .D(net470),
    .Q_N(_2095_),
    .Q(\MemCell.counter_value[8] ));
 sg13g2_dfrbp_1 _4592_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net696),
    .D(_0293_),
    .Q_N(_2094_),
    .Q(\MemCell.counter_value[9] ));
 sg13g2_dfrbp_1 _4593_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net695),
    .D(_0294_),
    .Q_N(_2093_),
    .Q(\MemCell.counter_value[10] ));
 sg13g2_dfrbp_1 _4594_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net696),
    .D(_0295_),
    .Q_N(_2092_),
    .Q(\MemCell.counter_value[11] ));
 sg13g2_dfrbp_1 _4595_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net696),
    .D(_0296_),
    .Q_N(_2091_),
    .Q(\MemCell.counter_value[12] ));
 sg13g2_dfrbp_1 _4596_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net698),
    .D(_0297_),
    .Q_N(_2090_),
    .Q(\MemCell.counter_value[13] ));
 sg13g2_dfrbp_1 _4597_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net698),
    .D(_0298_),
    .Q_N(_2089_),
    .Q(\MemCell.counter_value[14] ));
 sg13g2_dfrbp_1 _4598_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net697),
    .D(_0299_),
    .Q_N(_2088_),
    .Q(\MemCell.counter_value[15] ));
 sg13g2_dfrbp_1 _4599_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net688),
    .D(_0300_),
    .Q_N(_2087_),
    .Q(\MemCell.counter_value[0] ));
 sg13g2_dfrbp_1 _4600_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net688),
    .D(_0301_),
    .Q_N(_2086_),
    .Q(\MemCell.counter_value[1] ));
 sg13g2_dfrbp_1 _4601_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net688),
    .D(_0302_),
    .Q_N(_2085_),
    .Q(\MemCell.counter_value[2] ));
 sg13g2_dfrbp_1 _4602_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net688),
    .D(_0303_),
    .Q_N(_2084_),
    .Q(\MemCell.counter_value[3] ));
 sg13g2_dfrbp_1 _4603_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net688),
    .D(_0304_),
    .Q_N(_2083_),
    .Q(\MemCell.counter_value[4] ));
 sg13g2_dfrbp_1 _4604_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net689),
    .D(_0305_),
    .Q_N(_2082_),
    .Q(\MemCell.counter_value[5] ));
 sg13g2_dfrbp_1 _4605_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net689),
    .D(_0306_),
    .Q_N(_2081_),
    .Q(\MemCell.counter_value[6] ));
 sg13g2_dfrbp_1 _4606_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net689),
    .D(_0307_),
    .Q_N(_2080_),
    .Q(\MemCell.counter_value[7] ));
 sg13g2_dfrbp_1 _4607_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net736),
    .D(_0308_),
    .Q_N(_0103_),
    .Q(\MemCell.enable_pwm ));
 sg13g2_dfrbp_1 _4608_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net714),
    .D(_0309_),
    .Q_N(_2079_),
    .Q(\MemCell.counter[0] ));
 sg13g2_dfrbp_1 _4609_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net714),
    .D(_0310_),
    .Q_N(_2078_),
    .Q(\MemCell.counter[1] ));
 sg13g2_dfrbp_1 _4610_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net691),
    .D(_0311_),
    .Q_N(_2077_),
    .Q(\MemCell.dc3_reg[0][0] ));
 sg13g2_dfrbp_1 _4611_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net691),
    .D(_0312_),
    .Q_N(_2076_),
    .Q(\MemCell.dc3_reg[0][1] ));
 sg13g2_dfrbp_1 _4612_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net691),
    .D(_0313_),
    .Q_N(_2075_),
    .Q(\MemCell.dc3_reg[0][2] ));
 sg13g2_dfrbp_1 _4613_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net691),
    .D(_0314_),
    .Q_N(_2074_),
    .Q(\MemCell.dc3_reg[0][3] ));
 sg13g2_dfrbp_1 _4614_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net691),
    .D(_0315_),
    .Q_N(_2073_),
    .Q(\MemCell.dc3_reg[0][4] ));
 sg13g2_dfrbp_1 _4615_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net692),
    .D(_0316_),
    .Q_N(_2072_),
    .Q(\MemCell.dc3_reg[0][5] ));
 sg13g2_dfrbp_1 _4616_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net693),
    .D(_0317_),
    .Q_N(_2071_),
    .Q(\MemCell.dc3_reg[0][6] ));
 sg13g2_dfrbp_1 _4617_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net693),
    .D(_0318_),
    .Q_N(_2285_),
    .Q(\MemCell.dc3_reg[0][7] ));
 sg13g2_dfrbp_1 _4618_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net714),
    .D(net552),
    .Q_N(_2286_),
    .Q(\MemCell.curr_state[0] ));
 sg13g2_dfrbp_1 _4619_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net714),
    .D(\MemCell.next_state[1] ),
    .Q_N(_2287_),
    .Q(\MemCell.curr_state[1] ));
 sg13g2_dfrbp_1 _4620_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net714),
    .D(\MemCell.next_state[2] ),
    .Q_N(_0102_),
    .Q(\MemCell.curr_state[2] ));
 sg13g2_dfrbp_1 _4621_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net692),
    .D(_0319_),
    .Q_N(_2070_),
    .Q(\pwm_module.counter2[0] ));
 sg13g2_dfrbp_1 _4622_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net691),
    .D(_0320_),
    .Q_N(_2069_),
    .Q(\pwm_module.counter2[1] ));
 sg13g2_dfrbp_1 _4623_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net691),
    .D(_0321_),
    .Q_N(_2068_),
    .Q(\pwm_module.counter2[2] ));
 sg13g2_dfrbp_1 _4624_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net691),
    .D(_0322_),
    .Q_N(_2067_),
    .Q(\pwm_module.counter2[3] ));
 sg13g2_dfrbp_1 _4625_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net692),
    .D(net302),
    .Q_N(_2066_),
    .Q(\pwm_module.counter2[4] ));
 sg13g2_dfrbp_1 _4626_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net692),
    .D(net361),
    .Q_N(_2065_),
    .Q(\pwm_module.counter2[5] ));
 sg13g2_dfrbp_1 _4627_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net693),
    .D(_0325_),
    .Q_N(_2064_),
    .Q(\pwm_module.counter2[6] ));
 sg13g2_dfrbp_1 _4628_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net693),
    .D(_0326_),
    .Q_N(_2063_),
    .Q(\pwm_module.counter2[7] ));
 sg13g2_dfrbp_1 _4629_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net699),
    .D(_0327_),
    .Q_N(_2062_),
    .Q(\pwm_module.counter2[8] ));
 sg13g2_dfrbp_1 _4630_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net699),
    .D(_0328_),
    .Q_N(_2061_),
    .Q(\pwm_module.counter2[9] ));
 sg13g2_dfrbp_1 _4631_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net699),
    .D(net341),
    .Q_N(_2060_),
    .Q(\pwm_module.counter2[10] ));
 sg13g2_dfrbp_1 _4632_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net699),
    .D(net386),
    .Q_N(_2059_),
    .Q(\pwm_module.counter2[11] ));
 sg13g2_dfrbp_1 _4633_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net700),
    .D(_0331_),
    .Q_N(_2058_),
    .Q(\pwm_module.counter2[12] ));
 sg13g2_dfrbp_1 _4634_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net700),
    .D(net283),
    .Q_N(_2057_),
    .Q(\pwm_module.counter2[13] ));
 sg13g2_dfrbp_1 _4635_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net700),
    .D(_0333_),
    .Q_N(_2056_),
    .Q(\pwm_module.counter2[14] ));
 sg13g2_dfrbp_1 _4636_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net700),
    .D(net378),
    .Q_N(_2055_),
    .Q(\pwm_module.counter2[15] ));
 sg13g2_dfrbp_1 _4637_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net723),
    .D(_0335_),
    .Q_N(_2054_),
    .Q(\pwm_module.counter2[16] ));
 sg13g2_dfrbp_1 _4638_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net723),
    .D(_0336_),
    .Q_N(_2053_),
    .Q(\pwm_module.counter2[17] ));
 sg13g2_dfrbp_1 _4639_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net723),
    .D(net536),
    .Q_N(_2052_),
    .Q(\pwm_module.counter2[18] ));
 sg13g2_dfrbp_1 _4640_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net729),
    .D(_0338_),
    .Q_N(_2051_),
    .Q(\pwm_module.counter2[19] ));
 sg13g2_dfrbp_1 _4641_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net729),
    .D(_0339_),
    .Q_N(_2050_),
    .Q(\pwm_module.counter2[20] ));
 sg13g2_dfrbp_1 _4642_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net729),
    .D(_0340_),
    .Q_N(_2049_),
    .Q(\pwm_module.counter2[21] ));
 sg13g2_dfrbp_1 _4643_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net729),
    .D(net428),
    .Q_N(_2048_),
    .Q(\pwm_module.counter2[22] ));
 sg13g2_dfrbp_1 _4644_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net732),
    .D(_0342_),
    .Q_N(_2047_),
    .Q(\pwm_module.counter2[23] ));
 sg13g2_dfrbp_1 _4645_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net733),
    .D(_0343_),
    .Q_N(_2046_),
    .Q(\pwm_module.counter2[24] ));
 sg13g2_dfrbp_1 _4646_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net732),
    .D(_0344_),
    .Q_N(_2045_),
    .Q(\pwm_module.counter2[25] ));
 sg13g2_dfrbp_1 _4647_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net732),
    .D(_0345_),
    .Q_N(_2044_),
    .Q(\pwm_module.counter2[26] ));
 sg13g2_dfrbp_1 _4648_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net733),
    .D(_0346_),
    .Q_N(_2043_),
    .Q(\pwm_module.counter2[27] ));
 sg13g2_dfrbp_1 _4649_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net731),
    .D(net317),
    .Q_N(_2042_),
    .Q(\pwm_module.counter2[28] ));
 sg13g2_dfrbp_1 _4650_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net732),
    .D(net532),
    .Q_N(_2041_),
    .Q(\pwm_module.counter2[29] ));
 sg13g2_dfrbp_1 _4651_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net734),
    .D(net451),
    .Q_N(_2040_),
    .Q(\pwm_module.counter2[30] ));
 sg13g2_dfrbp_1 _4652_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net734),
    .D(_0350_),
    .Q_N(_2288_),
    .Q(\pwm_module.counter2[31] ));
 sg13g2_dfrbp_1 _4653_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net706),
    .D(_0032_),
    .Q_N(_2289_),
    .Q(\pwm_module.prescaler1[0] ));
 sg13g2_dfrbp_1 _4654_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net706),
    .D(_0043_),
    .Q_N(_2290_),
    .Q(\pwm_module.prescaler1[1] ));
 sg13g2_dfrbp_1 _4655_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net706),
    .D(net124),
    .Q_N(_2291_),
    .Q(\pwm_module.prescaler1[2] ));
 sg13g2_dfrbp_1 _4656_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net706),
    .D(net192),
    .Q_N(_2292_),
    .Q(\pwm_module.prescaler1[3] ));
 sg13g2_dfrbp_1 _4657_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net706),
    .D(_0058_),
    .Q_N(_2293_),
    .Q(\pwm_module.prescaler1[4] ));
 sg13g2_dfrbp_1 _4658_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net705),
    .D(_0059_),
    .Q_N(_2294_),
    .Q(\pwm_module.prescaler1[5] ));
 sg13g2_dfrbp_1 _4659_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net705),
    .D(_0060_),
    .Q_N(_2295_),
    .Q(\pwm_module.prescaler1[6] ));
 sg13g2_dfrbp_1 _4660_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net705),
    .D(_0061_),
    .Q_N(_2296_),
    .Q(\pwm_module.prescaler1[7] ));
 sg13g2_dfrbp_1 _4661_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net713),
    .D(_0062_),
    .Q_N(_2297_),
    .Q(\pwm_module.prescaler1[8] ));
 sg13g2_dfrbp_1 _4662_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net713),
    .D(_0063_),
    .Q_N(_2298_),
    .Q(\pwm_module.prescaler1[9] ));
 sg13g2_dfrbp_1 _4663_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net713),
    .D(_0033_),
    .Q_N(_2299_),
    .Q(\pwm_module.prescaler1[10] ));
 sg13g2_dfrbp_1 _4664_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net712),
    .D(_0034_),
    .Q_N(_2300_),
    .Q(\pwm_module.prescaler1[11] ));
 sg13g2_dfrbp_1 _4665_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net713),
    .D(_0035_),
    .Q_N(_2301_),
    .Q(\pwm_module.prescaler1[12] ));
 sg13g2_dfrbp_1 _4666_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net715),
    .D(_0036_),
    .Q_N(_2302_),
    .Q(\pwm_module.prescaler1[13] ));
 sg13g2_dfrbp_1 _4667_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net714),
    .D(_0037_),
    .Q_N(_2303_),
    .Q(\pwm_module.prescaler1[14] ));
 sg13g2_dfrbp_1 _4668_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net717),
    .D(_0038_),
    .Q_N(_2304_),
    .Q(\pwm_module.prescaler1[15] ));
 sg13g2_dfrbp_1 _4669_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net717),
    .D(_0039_),
    .Q_N(_2305_),
    .Q(\pwm_module.prescaler1[16] ));
 sg13g2_dfrbp_1 _4670_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net717),
    .D(_0040_),
    .Q_N(_2306_),
    .Q(\pwm_module.prescaler1[17] ));
 sg13g2_dfrbp_1 _4671_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net717),
    .D(_0041_),
    .Q_N(_2307_),
    .Q(\pwm_module.prescaler1[18] ));
 sg13g2_dfrbp_1 _4672_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net717),
    .D(_0042_),
    .Q_N(_2308_),
    .Q(\pwm_module.prescaler1[19] ));
 sg13g2_dfrbp_1 _4673_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net741),
    .D(_0044_),
    .Q_N(_2309_),
    .Q(\pwm_module.prescaler1[20] ));
 sg13g2_dfrbp_1 _4674_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net740),
    .D(_0045_),
    .Q_N(_2310_),
    .Q(\pwm_module.prescaler1[21] ));
 sg13g2_dfrbp_1 _4675_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net741),
    .D(_0046_),
    .Q_N(_2311_),
    .Q(\pwm_module.prescaler1[22] ));
 sg13g2_dfrbp_1 _4676_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net741),
    .D(_0047_),
    .Q_N(_2312_),
    .Q(\pwm_module.prescaler1[23] ));
 sg13g2_dfrbp_1 _4677_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net740),
    .D(_0048_),
    .Q_N(_2313_),
    .Q(\pwm_module.prescaler1[24] ));
 sg13g2_dfrbp_1 _4678_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net740),
    .D(_0049_),
    .Q_N(_2314_),
    .Q(\pwm_module.prescaler1[25] ));
 sg13g2_dfrbp_1 _4679_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net740),
    .D(_0050_),
    .Q_N(_2315_),
    .Q(\pwm_module.prescaler1[26] ));
 sg13g2_dfrbp_1 _4680_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net740),
    .D(net338),
    .Q_N(_2316_),
    .Q(\pwm_module.prescaler1[27] ));
 sg13g2_dfrbp_1 _4681_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net737),
    .D(_0052_),
    .Q_N(_2317_),
    .Q(\pwm_module.prescaler1[28] ));
 sg13g2_dfrbp_1 _4682_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net737),
    .D(net176),
    .Q_N(_2318_),
    .Q(\pwm_module.prescaler1[29] ));
 sg13g2_dfrbp_1 _4683_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net737),
    .D(_0055_),
    .Q_N(_2319_),
    .Q(\pwm_module.prescaler1[30] ));
 sg13g2_dfrbp_1 _4684_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net737),
    .D(_0056_),
    .Q_N(_2320_),
    .Q(\pwm_module.prescaler1[31] ));
 sg13g2_dfrbp_1 _4685_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net747),
    .D(_0097_),
    .Q_N(_2321_),
    .Q(uo_out[1]));
 sg13g2_dfrbp_1 _4686_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net747),
    .D(_0096_),
    .Q_N(_2322_),
    .Q(uo_out[0]));
 sg13g2_dfrbp_1 _4687_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net704),
    .D(_0064_),
    .Q_N(_2323_),
    .Q(\pwm_module.prescaler2[0] ));
 sg13g2_dfrbp_1 _4688_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net704),
    .D(_0075_),
    .Q_N(_2324_),
    .Q(\pwm_module.prescaler2[1] ));
 sg13g2_dfrbp_1 _4689_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net703),
    .D(net104),
    .Q_N(_2325_),
    .Q(\pwm_module.prescaler2[2] ));
 sg13g2_dfrbp_1 _4690_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net704),
    .D(net209),
    .Q_N(_2326_),
    .Q(\pwm_module.prescaler2[3] ));
 sg13g2_dfrbp_1 _4691_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net708),
    .D(_0090_),
    .Q_N(_2327_),
    .Q(\pwm_module.prescaler2[4] ));
 sg13g2_dfrbp_1 _4692_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net708),
    .D(_0091_),
    .Q_N(_2328_),
    .Q(\pwm_module.prescaler2[5] ));
 sg13g2_dfrbp_1 _4693_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net708),
    .D(_0092_),
    .Q_N(_2329_),
    .Q(\pwm_module.prescaler2[6] ));
 sg13g2_dfrbp_1 _4694_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net709),
    .D(_0093_),
    .Q_N(_2330_),
    .Q(\pwm_module.prescaler2[7] ));
 sg13g2_dfrbp_1 _4695_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net710),
    .D(_0094_),
    .Q_N(_2331_),
    .Q(\pwm_module.prescaler2[8] ));
 sg13g2_dfrbp_1 _4696_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net711),
    .D(_0095_),
    .Q_N(_2332_),
    .Q(\pwm_module.prescaler2[9] ));
 sg13g2_dfrbp_1 _4697_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net716),
    .D(_0065_),
    .Q_N(_2333_),
    .Q(\pwm_module.prescaler2[10] ));
 sg13g2_dfrbp_1 _4698_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net716),
    .D(net221),
    .Q_N(_2334_),
    .Q(\pwm_module.prescaler2[11] ));
 sg13g2_dfrbp_1 _4699_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net715),
    .D(_0067_),
    .Q_N(_2335_),
    .Q(\pwm_module.prescaler2[12] ));
 sg13g2_dfrbp_1 _4700_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net716),
    .D(_0068_),
    .Q_N(_2336_),
    .Q(\pwm_module.prescaler2[13] ));
 sg13g2_dfrbp_1 _4701_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net717),
    .D(_0069_),
    .Q_N(_2337_),
    .Q(\pwm_module.prescaler2[14] ));
 sg13g2_dfrbp_1 _4702_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net717),
    .D(net233),
    .Q_N(_2338_),
    .Q(\pwm_module.prescaler2[15] ));
 sg13g2_dfrbp_1 _4703_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net717),
    .D(_0071_),
    .Q_N(_2339_),
    .Q(\pwm_module.prescaler2[16] ));
 sg13g2_dfrbp_1 _4704_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net741),
    .D(_0072_),
    .Q_N(_2340_),
    .Q(\pwm_module.prescaler2[17] ));
 sg13g2_dfrbp_1 _4705_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net740),
    .D(_0073_),
    .Q_N(_2341_),
    .Q(\pwm_module.prescaler2[18] ));
 sg13g2_dfrbp_1 _4706_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net740),
    .D(_0074_),
    .Q_N(_2342_),
    .Q(\pwm_module.prescaler2[19] ));
 sg13g2_dfrbp_1 _4707_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net743),
    .D(_0076_),
    .Q_N(_2343_),
    .Q(\pwm_module.prescaler2[20] ));
 sg13g2_dfrbp_1 _4708_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net742),
    .D(_0077_),
    .Q_N(_2344_),
    .Q(\pwm_module.prescaler2[21] ));
 sg13g2_dfrbp_1 _4709_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net743),
    .D(_0078_),
    .Q_N(_2345_),
    .Q(\pwm_module.prescaler2[22] ));
 sg13g2_dfrbp_1 _4710_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net743),
    .D(_0079_),
    .Q_N(_2346_),
    .Q(\pwm_module.prescaler2[23] ));
 sg13g2_dfrbp_1 _4711_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net742),
    .D(_0080_),
    .Q_N(_2347_),
    .Q(\pwm_module.prescaler2[24] ));
 sg13g2_dfrbp_1 _4712_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net742),
    .D(net308),
    .Q_N(_2348_),
    .Q(\pwm_module.prescaler2[25] ));
 sg13g2_dfrbp_1 _4713_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net742),
    .D(_0082_),
    .Q_N(_2349_),
    .Q(\pwm_module.prescaler2[26] ));
 sg13g2_dfrbp_1 _4714_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net742),
    .D(_0083_),
    .Q_N(_2350_),
    .Q(\pwm_module.prescaler2[27] ));
 sg13g2_dfrbp_1 _4715_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net738),
    .D(_0084_),
    .Q_N(_2351_),
    .Q(\pwm_module.prescaler2[28] ));
 sg13g2_dfrbp_1 _4716_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net737),
    .D(net202),
    .Q_N(_2352_),
    .Q(\pwm_module.prescaler2[29] ));
 sg13g2_dfrbp_1 _4717_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net737),
    .D(_0087_),
    .Q_N(_2353_),
    .Q(\pwm_module.prescaler2[30] ));
 sg13g2_dfrbp_1 _4718_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net737),
    .D(_0088_),
    .Q_N(_2039_),
    .Q(\pwm_module.prescaler2[31] ));
 sg13g2_dfrbp_1 _4719_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net733),
    .D(_0351_),
    .Q_N(_2038_),
    .Q(\MemCell.dc3_reg[3][0] ));
 sg13g2_dfrbp_1 _4720_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net733),
    .D(_0352_),
    .Q_N(_2037_),
    .Q(\MemCell.dc3_reg[3][1] ));
 sg13g2_dfrbp_1 _4721_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net733),
    .D(_0353_),
    .Q_N(_2036_),
    .Q(\MemCell.dc3_reg[3][2] ));
 sg13g2_dfrbp_1 _4722_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net733),
    .D(_0354_),
    .Q_N(_2035_),
    .Q(\MemCell.dc3_reg[3][3] ));
 sg13g2_dfrbp_1 _4723_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net734),
    .D(_0355_),
    .Q_N(_2034_),
    .Q(\MemCell.dc3_reg[3][4] ));
 sg13g2_dfrbp_1 _4724_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net734),
    .D(_0356_),
    .Q_N(_2033_),
    .Q(\MemCell.dc3_reg[3][5] ));
 sg13g2_dfrbp_1 _4725_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net734),
    .D(_0357_),
    .Q_N(_2032_),
    .Q(\MemCell.dc3_reg[3][6] ));
 sg13g2_dfrbp_1 _4726_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net733),
    .D(_0358_),
    .Q_N(_2354_),
    .Q(\MemCell.dc3_reg[3][7] ));
 sg13g2_dfrbp_1 _4727_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net733),
    .D(_0098_),
    .Q_N(_2031_),
    .Q(uo_out[2]));
 sg13g2_dfrbp_1 _4728_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net687),
    .D(_0359_),
    .Q_N(_2030_),
    .Q(\pwm_module.counter1[0] ));
 sg13g2_dfrbp_1 _4729_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net687),
    .D(_0360_),
    .Q_N(_2029_),
    .Q(\pwm_module.counter1[1] ));
 sg13g2_dfrbp_1 _4730_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net687),
    .D(net189),
    .Q_N(_2028_),
    .Q(\pwm_module.counter1[2] ));
 sg13g2_dfrbp_1 _4731_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net688),
    .D(_0362_),
    .Q_N(_2027_),
    .Q(\pwm_module.counter1[3] ));
 sg13g2_dfrbp_1 _4732_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net690),
    .D(net418),
    .Q_N(_2026_),
    .Q(\pwm_module.counter1[4] ));
 sg13g2_dfrbp_1 _4733_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net689),
    .D(_0364_),
    .Q_N(_2025_),
    .Q(\pwm_module.counter1[5] ));
 sg13g2_dfrbp_1 _4734_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net690),
    .D(_0365_),
    .Q_N(_2024_),
    .Q(\pwm_module.counter1[6] ));
 sg13g2_dfrbp_1 _4735_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net690),
    .D(net486),
    .Q_N(_2023_),
    .Q(\pwm_module.counter1[7] ));
 sg13g2_dfrbp_1 _4736_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net695),
    .D(_0367_),
    .Q_N(_2022_),
    .Q(\pwm_module.counter1[8] ));
 sg13g2_dfrbp_1 _4737_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net695),
    .D(_0368_),
    .Q_N(_2021_),
    .Q(\pwm_module.counter1[9] ));
 sg13g2_dfrbp_1 _4738_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net695),
    .D(net416),
    .Q_N(_2020_),
    .Q(\pwm_module.counter1[10] ));
 sg13g2_dfrbp_1 _4739_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net695),
    .D(_0370_),
    .Q_N(_2019_),
    .Q(\pwm_module.counter1[11] ));
 sg13g2_dfrbp_1 _4740_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net697),
    .D(_0371_),
    .Q_N(_2018_),
    .Q(\pwm_module.counter1[12] ));
 sg13g2_dfrbp_1 _4741_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net697),
    .D(net540),
    .Q_N(_2017_),
    .Q(\pwm_module.counter1[13] ));
 sg13g2_dfrbp_1 _4742_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net697),
    .D(net392),
    .Q_N(_2016_),
    .Q(\pwm_module.counter1[14] ));
 sg13g2_dfrbp_1 _4743_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net697),
    .D(_0374_),
    .Q_N(_2015_),
    .Q(\pwm_module.counter1[15] ));
 sg13g2_dfrbp_1 _4744_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net720),
    .D(net491),
    .Q_N(_2014_),
    .Q(\pwm_module.counter1[16] ));
 sg13g2_dfrbp_1 _4745_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net720),
    .D(net460),
    .Q_N(_2013_),
    .Q(\pwm_module.counter1[17] ));
 sg13g2_dfrbp_1 _4746_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net720),
    .D(_0377_),
    .Q_N(_2012_),
    .Q(\pwm_module.counter1[18] ));
 sg13g2_dfrbp_1 _4747_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net720),
    .D(net403),
    .Q_N(_2011_),
    .Q(\pwm_module.counter1[19] ));
 sg13g2_dfrbp_1 _4748_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net721),
    .D(_0379_),
    .Q_N(_2010_),
    .Q(\pwm_module.counter1[20] ));
 sg13g2_dfrbp_1 _4749_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net722),
    .D(_0380_),
    .Q_N(_2009_),
    .Q(\pwm_module.counter1[21] ));
 sg13g2_dfrbp_1 _4750_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net723),
    .D(net370),
    .Q_N(_2008_),
    .Q(\pwm_module.counter1[22] ));
 sg13g2_dfrbp_1 _4751_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net721),
    .D(_0382_),
    .Q_N(_2007_),
    .Q(\pwm_module.counter1[23] ));
 sg13g2_dfrbp_1 _4752_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net722),
    .D(_0383_),
    .Q_N(_2006_),
    .Q(\pwm_module.counter1[24] ));
 sg13g2_dfrbp_1 _4753_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net722),
    .D(_0384_),
    .Q_N(_2005_),
    .Q(\pwm_module.counter1[25] ));
 sg13g2_dfrbp_1 _4754_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net722),
    .D(_0385_),
    .Q_N(_2004_),
    .Q(\pwm_module.counter1[26] ));
 sg13g2_dfrbp_1 _4755_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net722),
    .D(net516),
    .Q_N(_2003_),
    .Q(\pwm_module.counter1[27] ));
 sg13g2_dfrbp_1 _4756_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net722),
    .D(_0387_),
    .Q_N(_2002_),
    .Q(\pwm_module.counter1[28] ));
 sg13g2_dfrbp_1 _4757_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net722),
    .D(_0388_),
    .Q_N(_2001_),
    .Q(\pwm_module.counter1[29] ));
 sg13g2_dfrbp_1 _4758_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net722),
    .D(net501),
    .Q_N(_2000_),
    .Q(\pwm_module.counter1[30] ));
 sg13g2_dfrbp_1 _4759_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net728),
    .D(net241),
    .Q_N(_2355_),
    .Q(\pwm_module.counter1[31] ));
 sg13g2_dfrbp_1 _4760_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net708),
    .D(_0000_),
    .Q_N(_2356_),
    .Q(\pwm_module.prescaler0[0] ));
 sg13g2_dfrbp_1 _4761_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net708),
    .D(_0011_),
    .Q_N(_2357_),
    .Q(\pwm_module.prescaler0[1] ));
 sg13g2_dfrbp_1 _4762_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net708),
    .D(_0022_),
    .Q_N(_2358_),
    .Q(\pwm_module.prescaler0[2] ));
 sg13g2_dfrbp_1 _4763_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net708),
    .D(_0025_),
    .Q_N(_2359_),
    .Q(\pwm_module.prescaler0[3] ));
 sg13g2_dfrbp_1 _4764_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net708),
    .D(_0026_),
    .Q_N(_2360_),
    .Q(\pwm_module.prescaler0[4] ));
 sg13g2_dfrbp_1 _4765_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net709),
    .D(_0027_),
    .Q_N(_2361_),
    .Q(\pwm_module.prescaler0[5] ));
 sg13g2_dfrbp_1 _4766_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net709),
    .D(_0028_),
    .Q_N(_2362_),
    .Q(\pwm_module.prescaler0[6] ));
 sg13g2_dfrbp_1 _4767_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net709),
    .D(net118),
    .Q_N(_2363_),
    .Q(\pwm_module.prescaler0[7] ));
 sg13g2_dfrbp_1 _4768_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net709),
    .D(_0030_),
    .Q_N(_2364_),
    .Q(\pwm_module.prescaler0[8] ));
 sg13g2_dfrbp_1 _4769_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net710),
    .D(_0031_),
    .Q_N(_2365_),
    .Q(\pwm_module.prescaler0[9] ));
 sg13g2_dfrbp_1 _4770_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net710),
    .D(_0001_),
    .Q_N(_2366_),
    .Q(\pwm_module.prescaler0[10] ));
 sg13g2_dfrbp_1 _4771_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net711),
    .D(_0002_),
    .Q_N(_2367_),
    .Q(\pwm_module.prescaler0[11] ));
 sg13g2_dfrbp_1 _4772_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net710),
    .D(_0003_),
    .Q_N(_2368_),
    .Q(\pwm_module.prescaler0[12] ));
 sg13g2_dfrbp_1 _4773_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net710),
    .D(net134),
    .Q_N(_2369_),
    .Q(\pwm_module.prescaler0[13] ));
 sg13g2_dfrbp_1 _4774_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net716),
    .D(_0005_),
    .Q_N(_2370_),
    .Q(\pwm_module.prescaler0[14] ));
 sg13g2_dfrbp_1 _4775_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net715),
    .D(_0006_),
    .Q_N(_2371_),
    .Q(\pwm_module.prescaler0[15] ));
 sg13g2_dfrbp_1 _4776_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net749),
    .D(_0007_),
    .Q_N(_2372_),
    .Q(\pwm_module.prescaler0[16] ));
 sg13g2_dfrbp_1 _4777_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net749),
    .D(_0008_),
    .Q_N(_2373_),
    .Q(\pwm_module.prescaler0[17] ));
 sg13g2_dfrbp_1 _4778_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net748),
    .D(_0009_),
    .Q_N(_2374_),
    .Q(\pwm_module.prescaler0[18] ));
 sg13g2_dfrbp_1 _4779_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net748),
    .D(_0010_),
    .Q_N(_2375_),
    .Q(\pwm_module.prescaler0[19] ));
 sg13g2_dfrbp_1 _4780_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net750),
    .D(_0012_),
    .Q_N(_2376_),
    .Q(\pwm_module.prescaler0[20] ));
 sg13g2_dfrbp_1 _4781_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net750),
    .D(_0013_),
    .Q_N(_2377_),
    .Q(\pwm_module.prescaler0[21] ));
 sg13g2_dfrbp_1 _4782_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net750),
    .D(_0014_),
    .Q_N(_2378_),
    .Q(\pwm_module.prescaler0[22] ));
 sg13g2_dfrbp_1 _4783_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net751),
    .D(_0015_),
    .Q_N(_2379_),
    .Q(\pwm_module.prescaler0[23] ));
 sg13g2_dfrbp_1 _4784_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net748),
    .D(_0016_),
    .Q_N(_2380_),
    .Q(\pwm_module.prescaler0[24] ));
 sg13g2_dfrbp_1 _4785_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net748),
    .D(_0017_),
    .Q_N(_2381_),
    .Q(\pwm_module.prescaler0[25] ));
 sg13g2_dfrbp_1 _4786_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net748),
    .D(net267),
    .Q_N(_2382_),
    .Q(\pwm_module.prescaler0[26] ));
 sg13g2_dfrbp_1 _4787_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net748),
    .D(_0019_),
    .Q_N(_2383_),
    .Q(\pwm_module.prescaler0[27] ));
 sg13g2_dfrbp_1 _4788_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net746),
    .D(_0020_),
    .Q_N(_2384_),
    .Q(\pwm_module.prescaler0[28] ));
 sg13g2_dfrbp_1 _4789_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net746),
    .D(net53),
    .Q_N(_2385_),
    .Q(\pwm_module.prescaler0[29] ));
 sg13g2_dfrbp_1 _4790_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net746),
    .D(_0023_),
    .Q_N(_2386_),
    .Q(\pwm_module.prescaler0[30] ));
 sg13g2_dfrbp_1 _4791_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net746),
    .D(_0024_),
    .Q_N(_1999_),
    .Q(\pwm_module.prescaler0[31] ));
 sg13g2_tiehi _4460__19 (.L_HI(net19));
 sg13g2_tiehi _4459__20 (.L_HI(net20));
 sg13g2_tiehi _4458__21 (.L_HI(net21));
 sg13g2_tiehi _4457__22 (.L_HI(net22));
 sg13g2_tiehi _4456__23 (.L_HI(net23));
 sg13g2_tiehi _4455__24 (.L_HI(net24));
 sg13g2_tiehi _4454__25 (.L_HI(net25));
 sg13g2_tiehi _4451__26 (.L_HI(net26));
 sg13g2_tiehi _4450__27 (.L_HI(net27));
 sg13g2_tiehi _4449__28 (.L_HI(net28));
 sg13g2_tiehi _4448__29 (.L_HI(net29));
 sg13g2_tiehi _4447__30 (.L_HI(net30));
 sg13g2_tiehi _4446__31 (.L_HI(net31));
 sg13g2_tiehi _4452__32 (.L_HI(net32));
 sg13g2_tiehi tt_um_pwm_block_33 (.L_HI(net33));
 sg13g2_tiehi tt_um_pwm_block_34 (.L_HI(net34));
 sg13g2_tiehi tt_um_pwm_block_35 (.L_HI(net35));
 sg13g2_tiehi tt_um_pwm_block_36 (.L_HI(net36));
 sg13g2_tiehi tt_um_pwm_block_37 (.L_HI(net37));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_pwm_block_3 (.L_LO(net3));
 sg13g2_tielo tt_um_pwm_block_4 (.L_LO(net4));
 sg13g2_tielo tt_um_pwm_block_5 (.L_LO(net5));
 sg13g2_tielo tt_um_pwm_block_6 (.L_LO(net6));
 sg13g2_tielo tt_um_pwm_block_7 (.L_LO(net7));
 sg13g2_tielo tt_um_pwm_block_8 (.L_LO(net8));
 sg13g2_tielo tt_um_pwm_block_9 (.L_LO(net9));
 sg13g2_tielo tt_um_pwm_block_10 (.L_LO(net10));
 sg13g2_tielo tt_um_pwm_block_11 (.L_LO(net11));
 sg13g2_tielo tt_um_pwm_block_12 (.L_LO(net12));
 sg13g2_tielo tt_um_pwm_block_13 (.L_LO(net13));
 sg13g2_tielo tt_um_pwm_block_14 (.L_LO(net14));
 sg13g2_tielo tt_um_pwm_block_15 (.L_LO(net15));
 sg13g2_tielo tt_um_pwm_block_16 (.L_LO(net16));
 sg13g2_tielo tt_um_pwm_block_17 (.L_LO(net17));
 sg13g2_tiehi _4461__18 (.L_HI(net18));
 sg13g2_buf_4 fanout567 (.X(net567),
    .A(_1717_));
 sg13g2_buf_4 fanout568 (.X(net568),
    .A(_1241_));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(net571));
 sg13g2_buf_2 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_1716_),
    .X(net571));
 sg13g2_buf_4 fanout572 (.X(net572),
    .A(net576));
 sg13g2_buf_2 fanout573 (.A(net575),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(net576),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_1620_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_1526_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_1526_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(net584),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net584),
    .X(net582));
 sg13g2_buf_1 fanout583 (.A(net584),
    .X(net583));
 sg13g2_buf_1 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_4 fanout585 (.X(net585),
    .A(_1419_));
 sg13g2_buf_2 fanout586 (.A(_1256_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(net590),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_1240_),
    .X(net590));
 sg13g2_buf_4 fanout591 (.X(net591),
    .A(_1141_));
 sg13g2_buf_1 fanout592 (.A(_1141_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(net595),
    .X(net594));
 sg13g2_buf_1 fanout595 (.A(_1141_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_0964_),
    .X(net596));
 sg13g2_buf_1 fanout597 (.A(_0964_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(net600),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(net600),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_0964_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(net606),
    .X(net601));
 sg13g2_buf_1 fanout602 (.A(net606),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(net606),
    .X(net603));
 sg13g2_buf_1 fanout604 (.A(net605),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(net606),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_0791_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(net609),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_0617_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(net611),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_0617_),
    .X(net611));
 sg13g2_buf_8 fanout612 (.A(_0963_),
    .X(net612));
 sg13g2_buf_4 fanout613 (.X(net613),
    .A(_1378_));
 sg13g2_buf_4 fanout614 (.X(net614),
    .A(_1376_));
 sg13g2_buf_2 fanout615 (.A(_1367_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_1362_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_1362_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_1613_),
    .X(net618));
 sg13g2_buf_1 fanout619 (.A(_1613_),
    .X(net619));
 sg13g2_buf_4 fanout620 (.X(net620),
    .A(_1415_));
 sg13g2_buf_4 fanout621 (.X(net621),
    .A(_1370_));
 sg13g2_buf_1 fanout622 (.A(_1370_),
    .X(net622));
 sg13g2_buf_4 fanout623 (.X(net623),
    .A(_1358_));
 sg13g2_buf_2 fanout624 (.A(_1352_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_1352_),
    .X(net625));
 sg13g2_buf_4 fanout626 (.X(net626),
    .A(_1350_));
 sg13g2_buf_2 fanout627 (.A(_1345_),
    .X(net627));
 sg13g2_buf_1 fanout628 (.A(_1345_),
    .X(net628));
 sg13g2_buf_4 fanout629 (.X(net629),
    .A(_1341_));
 sg13g2_buf_2 fanout630 (.A(_1334_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_1334_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_1330_),
    .X(net632));
 sg13g2_buf_4 fanout633 (.X(net633),
    .A(_1327_));
 sg13g2_buf_2 fanout634 (.A(_1321_),
    .X(net634));
 sg13g2_buf_4 fanout635 (.X(net635),
    .A(_1404_));
 sg13g2_buf_1 fanout636 (.A(_1404_),
    .X(net636));
 sg13g2_buf_4 fanout637 (.X(net637),
    .A(_1398_));
 sg13g2_buf_2 fanout638 (.A(_1398_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_1389_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_1389_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_1382_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_1382_),
    .X(net642));
 sg13g2_buf_4 fanout643 (.X(net643),
    .A(_0099_));
 sg13g2_buf_4 fanout644 (.X(net644),
    .A(net645));
 sg13g2_buf_4 fanout645 (.X(net645),
    .A(_1863_));
 sg13g2_buf_4 fanout646 (.X(net646),
    .A(_1863_));
 sg13g2_buf_2 fanout647 (.A(net79),
    .X(net647));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(net538));
 sg13g2_buf_2 fanout649 (.A(net164),
    .X(net649));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(net46));
 sg13g2_buf_4 fanout651 (.X(net651),
    .A(\MemCell.enable_pwm ));
 sg13g2_buf_2 fanout652 (.A(\MemCell.prescale_reg[1][3] ),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(\MemCell.prescale_reg[2][3] ),
    .X(net653));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(net657));
 sg13g2_buf_2 fanout655 (.A(net657),
    .X(net655));
 sg13g2_buf_4 fanout656 (.X(net656),
    .A(net657));
 sg13g2_buf_4 fanout657 (.X(net657),
    .A(net480));
 sg13g2_buf_4 fanout658 (.X(net658),
    .A(net660));
 sg13g2_buf_4 fanout659 (.X(net659),
    .A(net660));
 sg13g2_buf_4 fanout660 (.X(net660),
    .A(\MemCell.o_RX_Byte[6] ));
 sg13g2_buf_4 fanout661 (.X(net661),
    .A(net663));
 sg13g2_buf_4 fanout662 (.X(net662),
    .A(net663));
 sg13g2_buf_8 fanout663 (.A(net508),
    .X(net663));
 sg13g2_buf_4 fanout664 (.X(net664),
    .A(net666));
 sg13g2_buf_4 fanout665 (.X(net665),
    .A(net666));
 sg13g2_buf_8 fanout666 (.A(net506),
    .X(net666));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(net669));
 sg13g2_buf_8 fanout668 (.A(net669),
    .X(net668));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(net544));
 sg13g2_buf_4 fanout670 (.X(net670),
    .A(net673));
 sg13g2_buf_2 fanout671 (.A(net673),
    .X(net671));
 sg13g2_buf_4 fanout672 (.X(net672),
    .A(net673));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(net504));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(net677));
 sg13g2_buf_2 fanout675 (.A(net677),
    .X(net675));
 sg13g2_buf_8 fanout676 (.A(net677),
    .X(net676));
 sg13g2_buf_4 fanout677 (.X(net677),
    .A(net447));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(net680));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(net680));
 sg13g2_buf_8 fanout680 (.A(net476),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(net425),
    .X(net681));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(uio_in[7]));
 sg13g2_buf_1 fanout683 (.A(uio_in[7]),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(net686),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(net686),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(uio_in[4]),
    .X(net686));
 sg13g2_buf_4 fanout687 (.X(net687),
    .A(net690));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(net690));
 sg13g2_buf_4 fanout689 (.X(net689),
    .A(net690));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(net702));
 sg13g2_buf_4 fanout691 (.X(net691),
    .A(net692));
 sg13g2_buf_4 fanout692 (.X(net692),
    .A(net694));
 sg13g2_buf_4 fanout693 (.X(net693),
    .A(net694));
 sg13g2_buf_2 fanout694 (.A(net702),
    .X(net694));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(net698));
 sg13g2_buf_2 fanout696 (.A(net698),
    .X(net696));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(net698));
 sg13g2_buf_2 fanout698 (.A(net702),
    .X(net698));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(net701));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(net701));
 sg13g2_buf_2 fanout701 (.A(net702),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(net753),
    .X(net702));
 sg13g2_buf_4 fanout703 (.X(net703),
    .A(net707));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(net707));
 sg13g2_buf_4 fanout705 (.X(net705),
    .A(net707));
 sg13g2_buf_2 fanout706 (.A(net707),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(net719),
    .X(net707));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(net709));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(net711));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(net711));
 sg13g2_buf_2 fanout711 (.A(net719),
    .X(net711));
 sg13g2_buf_4 fanout712 (.X(net712),
    .A(net714));
 sg13g2_buf_2 fanout713 (.A(net714),
    .X(net713));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(net719));
 sg13g2_buf_4 fanout715 (.X(net715),
    .A(net718));
 sg13g2_buf_2 fanout716 (.A(net718),
    .X(net716));
 sg13g2_buf_4 fanout717 (.X(net717),
    .A(net718));
 sg13g2_buf_2 fanout718 (.A(net719),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(net753),
    .X(net719));
 sg13g2_buf_4 fanout720 (.X(net720),
    .A(net721));
 sg13g2_buf_4 fanout721 (.X(net721),
    .A(net723));
 sg13g2_buf_4 fanout722 (.X(net722),
    .A(net723));
 sg13g2_buf_4 fanout723 (.X(net723),
    .A(net727));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(net726));
 sg13g2_buf_2 fanout725 (.A(net726),
    .X(net725));
 sg13g2_buf_4 fanout726 (.X(net726),
    .A(net727));
 sg13g2_buf_2 fanout727 (.A(net753),
    .X(net727));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(net729));
 sg13g2_buf_4 fanout729 (.X(net729),
    .A(net730));
 sg13g2_buf_4 fanout730 (.X(net730),
    .A(net735));
 sg13g2_buf_4 fanout731 (.X(net731),
    .A(net732));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(net735));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(net735));
 sg13g2_buf_2 fanout734 (.A(net735),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(net753),
    .X(net735));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(net739));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(net739));
 sg13g2_buf_4 fanout738 (.X(net738),
    .A(net739));
 sg13g2_buf_2 fanout739 (.A(net752),
    .X(net739));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(net744));
 sg13g2_buf_2 fanout741 (.A(net744),
    .X(net741));
 sg13g2_buf_4 fanout742 (.X(net742),
    .A(net744));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(net744));
 sg13g2_buf_2 fanout744 (.A(net752),
    .X(net744));
 sg13g2_buf_4 fanout745 (.X(net745),
    .A(net747));
 sg13g2_buf_2 fanout746 (.A(net747),
    .X(net746));
 sg13g2_buf_4 fanout747 (.X(net747),
    .A(net752));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(net751));
 sg13g2_buf_2 fanout749 (.A(net751),
    .X(net749));
 sg13g2_buf_4 fanout750 (.X(net750),
    .A(net751));
 sg13g2_buf_2 fanout751 (.A(net752),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(net753),
    .X(net752));
 sg13g2_buf_4 fanout753 (.X(net753),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(uio_in[6]),
    .X(net1));
 sg13g2_tielo tt_um_pwm_block_2 (.L_LO(net2));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_47_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_50_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_3_clk));
 sg13g2_inv_4 clkload8 (.A(clknet_leaf_43_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_35_clk));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_39_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_leaf_42_clk));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_6_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_20_clk));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_17_clk));
 sg13g2_inv_4 clkload15 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_28_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_25_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\spi_module.r2_RX_Done ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold2 (.A(\pwm_module.prescaler2[31] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold3 (.A(_1028_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold4 (.A(\pwm_module.prescaler1[31] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0855_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold6 (.A(\MemCell.dc1_reg[0][0] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0228_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold8 (.A(\MemCell.dc3_reg[0][0] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold9 (.A(\MemCell.counter[0] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold10 (.A(\pwm_module.prescaler0[31] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0677_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold12 (.A(\MemCell.dc2_reg[3][1] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold13 (.A(\MemCell.dc1_reg[2][5] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold14 (.A(\pwm_module.prescaler0[29] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0674_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0021_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold17 (.A(\MemCell.dc1_reg[2][0] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0212_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold19 (.A(\pwm_module.counter0[31] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold20 (.A(_1316_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold21 (.A(\MemCell.dc3_reg[2][0] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold22 (.A(\MemCell.dc2_reg[2][1] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold23 (.A(\MemCell.dc1_reg[2][3] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0215_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold25 (.A(\MemCell.dc1_reg[0][3] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0231_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold27 (.A(\MemCell.dc1_reg[2][7] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold28 (.A(\MemCell.dc2_reg[2][2] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold29 (.A(\MemCell.dc3_reg[2][3] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold30 (.A(\MemCell.dc2_reg[0][4] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold31 (.A(\MemCell.dc3_reg[0][2] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold32 (.A(\MemCell.dc1_reg[3][4] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold33 (.A(\MemCell.dc1_reg[0][7] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold34 (.A(\MemCell.dc3_reg[2][6] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold35 (.A(\MemCell.dc3_reg[0][3] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold36 (.A(\MemCell.dc2_reg[1][2] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold37 (.A(\MemCell.prescale_reg[1][3] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold38 (.A(\MemCell.dc3_reg[0][7] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold39 (.A(\MemCell.dc2_reg[0][0] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold40 (.A(\MemCell.dc1_reg[0][6] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0234_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold42 (.A(\pwm_module.counter1[5] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold43 (.A(\pwm_module.prescaler2[7] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0976_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold45 (.A(\MemCell.dc3_reg[1][2] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold46 (.A(\MemCell.dc1_reg[0][2] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold47 (.A(\MemCell.dc1_reg[2][4] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold48 (.A(\MemCell.dc3_reg[3][3] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold49 (.A(\MemCell.dc1_reg[1][4] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0224_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold51 (.A(\pwm_module.prescaler1[15] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0818_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold53 (.A(\MemCell.dc1_reg[2][2] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0214_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold55 (.A(\MemCell.dc2_reg[3][3] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold56 (.A(\MemCell.dc3_reg[2][1] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold57 (.A(\MemCell.dc1_reg[3][5] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold58 (.A(\MemCell.dc2_reg[2][0] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold59 (.A(\pwm_module.prescaler0[0] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold60 (.A(\MemCell.dc3_reg[1][7] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold61 (.A(\MemCell.dc3_reg[3][5] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold62 (.A(\MemCell.dc3_reg[0][1] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold63 (.A(\MemCell.dc1_reg[0][1] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold64 (.A(\pwm_module.prescaler2[0] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold65 (.A(\pwm_module.prescaler2[2] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0967_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0086_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold68 (.A(\MemCell.dc2_reg[2][3] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold69 (.A(\MemCell.dc1_reg[1][5] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0225_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold71 (.A(\MemCell.dc1_reg[1][1] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold72 (.A(\MemCell.dc2_reg[2][5] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold73 (.A(\pwm_module.prescaler2[9] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0979_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold75 (.A(\MemCell.prescale_reg[2][3] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0247_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold77 (.A(\pwm_module.prescaler0[2] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0620_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold79 (.A(\pwm_module.prescaler0[7] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0630_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0029_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold82 (.A(\pwm_module.prescaler1[0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold83 (.A(\MemCell.dc2_reg[3][7] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold84 (.A(\MemCell.dc3_reg[0][5] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold85 (.A(\pwm_module.prescaler1[2] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0794_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0054_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold88 (.A(\MemCell.dc1_reg[1][3] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold89 (.A(\MemCell.dc3_reg[1][3] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold90 (.A(\MemCell.dc2_reg[1][3] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold91 (.A(\MemCell.dc2_reg[1][7] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold92 (.A(\MemCell.dc3_reg[1][1] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold93 (.A(\MemCell.dc1_reg[0][5] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0233_),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold95 (.A(\pwm_module.prescaler0[13] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0641_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0004_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold98 (.A(\pwm_module.prescaler1[9] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0806_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold100 (.A(\MemCell.dc2_reg[2][6] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold101 (.A(\MemCell.dc2_reg[0][5] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold102 (.A(\MemCell.dc1_reg[1][7] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold103 (.A(\MemCell.dc3_reg[1][4] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold104 (.A(\MemCell.dc2_reg[1][0] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0188_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold106 (.A(\MemCell.dc2_reg[1][1] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold107 (.A(\MemCell.dc1_reg[2][6] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0218_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold109 (.A(\MemCell.dc3_reg[3][7] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold110 (.A(\pwm_module.prescaler1[11] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0810_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold112 (.A(\MemCell.dc2_reg[3][0] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold113 (.A(\MemCell.dc3_reg[0][6] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold114 (.A(\MemCell.dc1_reg[0][4] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0232_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold116 (.A(\MemCell.dc1_reg[3][6] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold117 (.A(\pwm_module.prescaler0[15] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0644_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold119 (.A(\MemCell.dc2_reg[3][5] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold120 (.A(\MemCell.dc3_reg[3][2] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold121 (.A(\MemCell.dc1_reg[2][1] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0213_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold123 (.A(\MemCell.dc1_reg[3][7] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold124 (.A(\MemCell.dc3_reg[1][0] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0252_),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold126 (.A(\MemCell.dc3_reg[3][6] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold127 (.A(\pwm_module.counter2[1] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold128 (.A(_1533_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold129 (.A(\pwm_module.counter0[10] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold130 (.A(_1262_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold131 (.A(\MemCell.dc2_reg[3][6] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold132 (.A(\MemCell.dc1_reg[1][2] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold133 (.A(\MemCell.dc2_reg[0][3] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold134 (.A(\pwm_module.prescaler1[7] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0803_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold136 (.A(\MemCell.dc3_reg[2][2] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold137 (.A(\pwm_module.prescaler1[29] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0851_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0053_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold140 (.A(\MemCell.dc1_reg[1][6] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0226_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold142 (.A(\pwm_module.counter2[31] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold143 (.A(_1612_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold144 (.A(\MemCell.dc2_reg[0][7] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold145 (.A(\MemCell.dc3_reg[1][5] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold146 (.A(\MemCell.dc2_reg[1][4] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold147 (.A(\MemCell.dc3_reg[1][6] ),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold148 (.A(\MemCell.dc2_reg[1][6] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold149 (.A(\pwm_module.prescaler1[12] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold150 (.A(\MemCell.dc3_reg[0][4] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold151 (.A(\pwm_module.counter1[2] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0361_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold153 (.A(\pwm_module.prescaler1[3] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0796_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0057_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold156 (.A(\MemCell.dc3_reg[2][7] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold157 (.A(\MemCell.dc3_reg[2][4] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold158 (.A(\MemCell.dc3_reg[2][5] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold159 (.A(\MemCell.dc3_reg[3][1] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold160 (.A(\MemCell.dc2_reg[1][5] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold161 (.A(\pwm_module.prescaler0[9] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0634_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold163 (.A(\pwm_module.prescaler2[29] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold164 (.A(_1024_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0085_),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold166 (.A(\pwm_module.counter0[23] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold167 (.A(\pwm_module.prescaler0[23] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0661_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold169 (.A(\pwm_module.prescaler1[13] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold170 (.A(\pwm_module.prescaler2[3] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0969_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0089_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold173 (.A(\MemCell.dc2_reg[3][4] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold174 (.A(\MemCell.dc2_reg[0][6] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold175 (.A(\pwm_module.prescaler0[11] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0637_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold177 (.A(\MemCell.dc3_reg[3][0] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold178 (.A(\pwm_module.counter0[2] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0110_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold180 (.A(\MemCell.dc3_reg[3][4] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold181 (.A(\MemCell.dc2_reg[0][2] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold182 (.A(\pwm_module.prescaler2[11] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0983_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0066_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold185 (.A(\MemCell.counter_value[0] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold186 (.A(\pwm_module.prescaler0[19] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0652_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold188 (.A(\pwm_module.prescaler2[19] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold189 (.A(_1001_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold190 (.A(\MemCell.dc1_reg[1][0] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold191 (.A(\pwm_module.prescaler2[27] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold192 (.A(_1019_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold193 (.A(\MemCell.dc1_reg[3][1] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold194 (.A(\pwm_module.prescaler2[15] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0992_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0070_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold197 (.A(\MemCell.dc2_reg[0][1] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold198 (.A(\pwm_module.prescaler1[30] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0853_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold200 (.A(\pwm_module.prescaler2[23] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold201 (.A(_1010_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold202 (.A(\MemCell.dc2_reg[2][7] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold203 (.A(\pwm_module.counter1[31] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0390_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold205 (.A(\MemCell.dc2_reg[3][2] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold206 (.A(\pwm_module.prescaler1[5] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0799_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold208 (.A(\pwm_module.prescaler2[30] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold209 (.A(_1026_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold210 (.A(\pwm_module.prescaler2[26] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold211 (.A(_1017_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold212 (.A(\pwm_module.prescaler2[13] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0987_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold214 (.A(\pwm_module.prescaler2[28] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold215 (.A(\pwm_module.prescaler0[3] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0623_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold217 (.A(\pwm_module.counter1[25] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold218 (.A(_1771_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold219 (.A(\pwm_module.prescaler2[21] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold220 (.A(_1006_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold221 (.A(\pwm_module.prescaler0[6] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0629_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold223 (.A(\MemCell.prescale_reg[0][0] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold224 (.A(\pwm_module.prescaler0[5] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0626_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold226 (.A(\pwm_module.prescaler0[30] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0676_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold228 (.A(\pwm_module.prescaler0[26] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0668_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0018_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold231 (.A(\MemCell.dc1_reg[3][0] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0204_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold233 (.A(\pwm_module.prescaler0[27] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0670_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold235 (.A(\MemCell.dc2_reg[2][4] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold236 (.A(\pwm_module.prescaler2[18] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0999_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold238 (.A(\pwm_module.prescaler2[20] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold239 (.A(_1004_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold240 (.A(\pwm_module.prescaler0[17] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0648_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold242 (.A(\pwm_module.counter1[11] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold243 (.A(\pwm_module.prescaler1[20] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold244 (.A(\pwm_module.prescaler2[22] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold245 (.A(\pwm_module.counter2[12] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0332_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold247 (.A(\pwm_module.prescaler1[17] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0824_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold249 (.A(\pwm_module.prescaler2[17] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0997_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold251 (.A(\pwm_module.counter0[9] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0117_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold253 (.A(\pwm_module.counter0[30] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0138_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold255 (.A(\pwm_module.prescaler1[19] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0828_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold257 (.A(\MemCell.dc1_reg[3][3] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold258 (.A(\pwm_module.counter2[9] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold259 (.A(_1553_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold260 (.A(\MemCell.dc1_reg[3][2] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold261 (.A(\MemCell.prescale_reg[3][4] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0240_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold263 (.A(\pwm_module.counter2[4] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold264 (.A(_1535_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold265 (.A(_0323_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold266 (.A(\pwm_module.prescaler0[22] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0659_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold268 (.A(\MemCell.counter_value[6] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold269 (.A(\pwm_module.prescaler2[25] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold270 (.A(_1015_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0081_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold272 (.A(\pwm_module.prescaler1[1] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold273 (.A(\pwm_module.prescaler2[5] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0972_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold275 (.A(\pwm_module.prescaler0[24] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold276 (.A(\pwm_module.prescaler1[25] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0842_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold278 (.A(\pwm_module.counter2[26] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold279 (.A(\pwm_module.counter2[27] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0347_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold281 (.A(\pwm_module.prescaler2[14] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0990_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold283 (.A(\pwm_module.prescaler1[4] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0797_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold285 (.A(\pwm_module.counter2[11] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold286 (.A(\pwm_module.prescaler1[8] ),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0805_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold288 (.A(\pwm_module.prescaler0[4] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold289 (.A(\pwm_module.counter0[11] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold290 (.A(\pwm_module.prescaler2[16] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0995_),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold292 (.A(\pwm_module.prescaler0[10] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0636_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold294 (.A(\pwm_module.prescaler1[6] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold295 (.A(\pwm_module.prescaler1[10] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold296 (.A(\pwm_module.prescaler0[12] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0640_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold298 (.A(\MemCell.counter_value[28] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold299 (.A(\pwm_module.prescaler1[27] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0846_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0051_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold302 (.A(\MemCell.counter_value[1] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold303 (.A(\pwm_module.counter2[10] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0329_),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold305 (.A(\pwm_module.counter0[26] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0134_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold307 (.A(\pwm_module.prescaler1[14] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold308 (.A(\MemCell.prescale_reg[1][0] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0260_),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold310 (.A(\pwm_module.prescaler2[8] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold311 (.A(\pwm_module.prescaler0[14] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold312 (.A(\pwm_module.counter2[6] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold313 (.A(\MemCell.prescale_reg[0][4] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold314 (.A(\MemCell.counter_value[9] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold315 (.A(\MemCell.counter_value[13] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold316 (.A(\pwm_module.prescaler0[21] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0657_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold318 (.A(\pwm_module.prescaler2[6] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold319 (.A(\pwm_module.counter1[28] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold320 (.A(_1777_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold321 (.A(\MemCell.counter_value[3] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold322 (.A(\pwm_module.prescaler2[24] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold323 (.A(\pwm_module.counter2[5] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0324_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold325 (.A(\pwm_module.counter2[0] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold326 (.A(\pwm_module.prescaler1[21] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold327 (.A(\MemCell.prescale_reg[3][6] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0242_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold329 (.A(\pwm_module.prescaler0[28] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold330 (.A(\MemCell.counter_value[21] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold331 (.A(\MemCell.counter_value[31] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold332 (.A(\pwm_module.counter1[22] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0381_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold334 (.A(\pwm_module.counter0[24] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold335 (.A(\pwm_module.prescaler2[10] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold336 (.A(\pwm_module.counter0[22] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0130_),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold338 (.A(\pwm_module.prescaler1[28] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0849_),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold340 (.A(\pwm_module.counter2[14] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0334_),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold342 (.A(\pwm_module.prescaler1[26] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold343 (.A(\MemCell.counter_value[10] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold344 (.A(\pwm_module.prescaler0[25] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold345 (.A(\pwm_module.prescaler0[1] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold346 (.A(\pwm_module.counter1[23] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold347 (.A(\pwm_module.prescaler2[1] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0103_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0330_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold350 (.A(\pwm_module.counter0[16] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold351 (.A(\pwm_module.prescaler2[4] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0970_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold353 (.A(\pwm_module.prescaler0[20] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold354 (.A(\pwm_module.counter1[14] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0373_),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold356 (.A(\pwm_module.prescaler2[12] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold357 (.A(\pwm_module.counter0[7] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0115_),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold359 (.A(\pwm_module.counter0[0] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold360 (.A(\pwm_module.counter1[12] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold361 (.A(\pwm_module.counter0[19] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0127_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold363 (.A(\pwm_module.prescaler1[23] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0837_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold365 (.A(\pwm_module.counter1[19] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0378_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold367 (.A(\pwm_module.prescaler0[8] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold368 (.A(\MemCell.enable_pwm ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold369 (.A(\MemCell.prescale_reg[1][1] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold370 (.A(\MemCell.counter_value[11] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold371 (.A(\MemCell.counter_value[14] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold372 (.A(\MemCell.counter_value[24] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0276_),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold374 (.A(\pwm_module.prescaler1[22] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold375 (.A(\MemCell.counter_value[15] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold376 (.A(\pwm_module.prescaler0[16] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold377 (.A(\pwm_module.counter1[9] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold378 (.A(_1738_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0369_),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold380 (.A(\pwm_module.counter1[3] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0363_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold382 (.A(\pwm_module.prescaler1[16] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold383 (.A(\pwm_module.prescaler1[18] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold384 (.A(\pwm_module.counter1[0] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold385 (.A(\pwm_module.counter0[12] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0121_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold387 (.A(\MemCell.prescale_reg[0][2] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold388 (.A(\pwm_module.counter0[5] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold389 (.A(_1253_),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold390 (.A(\pwm_module.counter2[22] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0341_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold392 (.A(\MemCell.prescale_reg[0][3] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0271_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold394 (.A(\MemCell.prescale_reg[0][1] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold395 (.A(\pwm_module.prescaler0[18] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0651_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold397 (.A(\MemCell.counter_value[26] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold398 (.A(\MemCell.counter_value[2] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold399 (.A(\spi_module.r3_RX_Done ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0145_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold401 (.A(\MemCell.prescale_reg[0][5] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0273_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold403 (.A(\MemCell.counter_value[29] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold404 (.A(\pwm_module.counter2[3] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold405 (.A(\MemCell.prescale_reg[3][3] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold406 (.A(\MemCell.counter_value[25] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0277_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold408 (.A(\pwm_module.prescaler1[24] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0840_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold410 (.A(\MemCell.o_RX_Byte[1] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0237_),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold412 (.A(\MemCell.counter_value[30] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold413 (.A(\pwm_module.counter2[30] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold414 (.A(_0349_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold415 (.A(\pwm_module.counter2[8] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold416 (.A(\pwm_module.counter0[17] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0126_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold418 (.A(\pwm_module.counter2[21] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold419 (.A(\MemCell.prescale_reg[0][7] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold420 (.A(\MemCell.counter_value[16] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0284_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold422 (.A(\pwm_module.counter1[17] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0376_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold424 (.A(\MemCell.counter_value[17] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold425 (.A(\pwm_module.counter0[15] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold426 (.A(\pwm_module.counter2[25] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold427 (.A(\pwm_module.counter2[7] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold428 (.A(\pwm_module.counter0[3] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold429 (.A(_0112_),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold430 (.A(\MemCell.prescale_reg[1][2] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold431 (.A(\MemCell.prescale_reg[1][6] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold432 (.A(\MemCell.counter_value[8] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold433 (.A(_0292_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold434 (.A(\pwm_module.counter0[28] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0136_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold436 (.A(\pwm_module.counter1[15] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold437 (.A(\MemCell.curr_state[2] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold438 (.A(_1409_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold439 (.A(\MemCell.o_RX_Byte[0] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold440 (.A(_0244_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold441 (.A(\MemCell.counter_value[18] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold442 (.A(\MemCell.prescale_reg[2][1] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold443 (.A(\MemCell.o_RX_Byte[7] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0251_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold445 (.A(\pwm_module.counter2[13] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold446 (.A(\pwm_module.counter0[20] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0128_),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold448 (.A(\pwm_module.counter1[7] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold449 (.A(_0366_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold450 (.A(\MemCell.prescale_reg[3][7] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold451 (.A(\pwm_module.counter0[14] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold452 (.A(\MemCell.prescale_reg[1][4] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold453 (.A(\pwm_module.counter1[16] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0375_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold455 (.A(\MemCell.prescale_reg[3][2] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0238_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold457 (.A(\MemCell.prescale_reg[1][5] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold458 (.A(\MemCell.prescale_reg[1][7] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold459 (.A(\MemCell.prescale_reg[0][6] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold460 (.A(\MemCell.counter_value[19] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold461 (.A(\MemCell.counter_value[5] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold462 (.A(\pwm_module.counter2[16] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold463 (.A(\pwm_module.counter1[30] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0389_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold465 (.A(\MemCell.counter_value[23] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold466 (.A(\MemCell.counter_value[20] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold467 (.A(\MemCell.o_RX_Byte[2] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0246_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold469 (.A(\MemCell.o_RX_Byte[4] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold470 (.A(_0248_),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold471 (.A(\MemCell.o_RX_Byte[5] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0249_),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold473 (.A(\MemCell.counter_value[12] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold474 (.A(\MemCell.counter_value[7] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold475 (.A(\MemCell.prescale_reg[3][5] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold476 (.A(\MemCell.counter_value[22] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold477 (.A(\pwm_module.counter1[20] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold478 (.A(\pwm_module.counter1[27] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0386_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold480 (.A(\MemCell.prescale_reg[3][0] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold481 (.A(\pwm_module.counter0[25] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold482 (.A(\pwm_module.counter0[27] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold483 (.A(\MemCell.prescale_reg[2][6] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0250_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold485 (.A(\pwm_module.counter1[8] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold486 (.A(\pwm_module.counter2[24] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold487 (.A(\pwm_module.counter2[23] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold488 (.A(\pwm_module.counter1[24] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold489 (.A(\pwm_module.counter2[19] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold490 (.A(\MemCell.counter[1] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold491 (.A(\pwm_module.counter1[0] ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold492 (.A(\pwm_module.counter0[8] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold493 (.A(\MemCell.counter_value[4] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold494 (.A(\pwm_module.counter2[29] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0348_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold496 (.A(\pwm_module.counter0[29] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold497 (.A(\pwm_module.counter0[1] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold498 (.A(\pwm_module.counter2[18] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0337_),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold500 (.A(\pwm_module.counter1[21] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold501 (.A(\pwm_module.counter2[17] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold502 (.A(\pwm_module.counter1[13] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0372_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold504 (.A(\pwm_module.counter1[1] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold505 (.A(\pwm_module.counter2[20] ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold506 (.A(\pwm_module.counter1[6] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold507 (.A(\MemCell.o_RX_Byte[3] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold508 (.A(\pwm_module.counter1[18] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold509 (.A(\MemCell.counter_value[27] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold510 (.A(\pwm_module.counter1[29] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold511 (.A(\pwm_module.counter0[21] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold512 (.A(\pwm_module.counter1[26] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold513 (.A(_0102_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold514 (.A(_1045_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold515 (.A(\MemCell.next_state[0] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold516 (.A(\pwm_module.prescaler0[16] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold517 (.A(\pwm_module.prescaler0[1] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold518 (.A(\pwm_module.prescaler1[24] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold519 (.A(\pwm_module.prescaler1[10] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold520 (.A(\pwm_module.counter1[13] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold521 (.A(\pwm_module.prescaler0[8] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold522 (.A(\pwm_module.counter1[9] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold523 (.A(\pwm_module.prescaler2[6] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold524 (.A(\pwm_module.prescaler2[12] ),
    .X(net561));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_4 FILLER_0_56 ();
 sg13g2_fill_2 FILLER_0_60 ();
 sg13g2_decap_8 FILLER_0_67 ();
 sg13g2_decap_8 FILLER_0_74 ();
 sg13g2_decap_8 FILLER_0_81 ();
 sg13g2_decap_8 FILLER_0_88 ();
 sg13g2_decap_8 FILLER_0_95 ();
 sg13g2_decap_8 FILLER_0_102 ();
 sg13g2_decap_8 FILLER_0_109 ();
 sg13g2_decap_8 FILLER_0_116 ();
 sg13g2_decap_8 FILLER_0_123 ();
 sg13g2_fill_1 FILLER_0_135 ();
 sg13g2_decap_8 FILLER_0_160 ();
 sg13g2_decap_8 FILLER_0_167 ();
 sg13g2_decap_8 FILLER_0_174 ();
 sg13g2_decap_8 FILLER_0_181 ();
 sg13g2_decap_8 FILLER_0_188 ();
 sg13g2_decap_8 FILLER_0_195 ();
 sg13g2_decap_8 FILLER_0_202 ();
 sg13g2_decap_8 FILLER_0_209 ();
 sg13g2_decap_8 FILLER_0_216 ();
 sg13g2_decap_8 FILLER_0_223 ();
 sg13g2_decap_8 FILLER_0_230 ();
 sg13g2_decap_8 FILLER_0_237 ();
 sg13g2_decap_8 FILLER_0_244 ();
 sg13g2_decap_8 FILLER_0_251 ();
 sg13g2_decap_8 FILLER_0_258 ();
 sg13g2_decap_8 FILLER_0_265 ();
 sg13g2_decap_8 FILLER_0_272 ();
 sg13g2_decap_8 FILLER_0_279 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_fill_2 FILLER_0_293 ();
 sg13g2_fill_2 FILLER_0_303 ();
 sg13g2_fill_1 FILLER_0_305 ();
 sg13g2_fill_1 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_fill_1 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_83 ();
 sg13g2_decap_8 FILLER_1_90 ();
 sg13g2_decap_8 FILLER_1_97 ();
 sg13g2_decap_8 FILLER_1_104 ();
 sg13g2_decap_4 FILLER_1_111 ();
 sg13g2_fill_1 FILLER_1_115 ();
 sg13g2_fill_2 FILLER_1_151 ();
 sg13g2_decap_8 FILLER_1_179 ();
 sg13g2_decap_8 FILLER_1_186 ();
 sg13g2_decap_8 FILLER_1_193 ();
 sg13g2_decap_8 FILLER_1_200 ();
 sg13g2_decap_8 FILLER_1_207 ();
 sg13g2_decap_8 FILLER_1_214 ();
 sg13g2_decap_8 FILLER_1_221 ();
 sg13g2_decap_8 FILLER_1_228 ();
 sg13g2_decap_8 FILLER_1_235 ();
 sg13g2_decap_8 FILLER_1_242 ();
 sg13g2_decap_8 FILLER_1_249 ();
 sg13g2_decap_8 FILLER_1_256 ();
 sg13g2_decap_8 FILLER_1_263 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_277 ();
 sg13g2_decap_4 FILLER_1_284 ();
 sg13g2_fill_1 FILLER_1_288 ();
 sg13g2_fill_1 FILLER_1_349 ();
 sg13g2_decap_8 FILLER_1_376 ();
 sg13g2_decap_8 FILLER_1_383 ();
 sg13g2_decap_8 FILLER_1_390 ();
 sg13g2_decap_8 FILLER_1_397 ();
 sg13g2_decap_4 FILLER_1_404 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_fill_1 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_fill_2 FILLER_2_98 ();
 sg13g2_fill_1 FILLER_2_100 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_fill_2 FILLER_2_277 ();
 sg13g2_fill_1 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_4 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_25 ();
 sg13g2_fill_2 FILLER_3_98 ();
 sg13g2_decap_4 FILLER_3_114 ();
 sg13g2_decap_8 FILLER_3_185 ();
 sg13g2_decap_8 FILLER_3_192 ();
 sg13g2_decap_8 FILLER_3_199 ();
 sg13g2_decap_8 FILLER_3_206 ();
 sg13g2_decap_8 FILLER_3_213 ();
 sg13g2_decap_8 FILLER_3_220 ();
 sg13g2_decap_8 FILLER_3_227 ();
 sg13g2_decap_8 FILLER_3_234 ();
 sg13g2_decap_8 FILLER_3_241 ();
 sg13g2_decap_8 FILLER_3_248 ();
 sg13g2_decap_8 FILLER_3_255 ();
 sg13g2_decap_4 FILLER_3_262 ();
 sg13g2_fill_1 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_4 FILLER_4_28 ();
 sg13g2_fill_2 FILLER_4_32 ();
 sg13g2_fill_2 FILLER_4_42 ();
 sg13g2_fill_1 FILLER_4_44 ();
 sg13g2_decap_4 FILLER_4_54 ();
 sg13g2_fill_2 FILLER_4_82 ();
 sg13g2_fill_1 FILLER_4_84 ();
 sg13g2_fill_2 FILLER_4_121 ();
 sg13g2_fill_1 FILLER_4_129 ();
 sg13g2_decap_8 FILLER_4_183 ();
 sg13g2_decap_8 FILLER_4_190 ();
 sg13g2_decap_8 FILLER_4_197 ();
 sg13g2_decap_8 FILLER_4_204 ();
 sg13g2_decap_8 FILLER_4_211 ();
 sg13g2_decap_8 FILLER_4_218 ();
 sg13g2_decap_8 FILLER_4_225 ();
 sg13g2_decap_8 FILLER_4_232 ();
 sg13g2_decap_8 FILLER_4_239 ();
 sg13g2_decap_8 FILLER_4_246 ();
 sg13g2_fill_2 FILLER_4_253 ();
 sg13g2_fill_1 FILLER_4_338 ();
 sg13g2_fill_2 FILLER_4_353 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_fill_2 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_23 ();
 sg13g2_fill_2 FILLER_5_63 ();
 sg13g2_fill_1 FILLER_5_65 ();
 sg13g2_fill_1 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_212 ();
 sg13g2_decap_8 FILLER_5_219 ();
 sg13g2_decap_8 FILLER_5_226 ();
 sg13g2_decap_8 FILLER_5_233 ();
 sg13g2_decap_8 FILLER_5_240 ();
 sg13g2_decap_4 FILLER_5_247 ();
 sg13g2_fill_1 FILLER_5_251 ();
 sg13g2_fill_2 FILLER_5_273 ();
 sg13g2_fill_1 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_4 FILLER_6_21 ();
 sg13g2_fill_1 FILLER_6_25 ();
 sg13g2_fill_1 FILLER_6_75 ();
 sg13g2_fill_1 FILLER_6_84 ();
 sg13g2_fill_1 FILLER_6_164 ();
 sg13g2_fill_2 FILLER_6_178 ();
 sg13g2_fill_1 FILLER_6_180 ();
 sg13g2_fill_1 FILLER_6_196 ();
 sg13g2_fill_2 FILLER_6_270 ();
 sg13g2_fill_1 FILLER_6_272 ();
 sg13g2_fill_2 FILLER_6_281 ();
 sg13g2_fill_1 FILLER_6_283 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_4 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_4 FILLER_7_21 ();
 sg13g2_fill_1 FILLER_7_39 ();
 sg13g2_fill_1 FILLER_7_52 ();
 sg13g2_decap_4 FILLER_7_81 ();
 sg13g2_fill_2 FILLER_7_103 ();
 sg13g2_decap_4 FILLER_7_114 ();
 sg13g2_fill_1 FILLER_7_130 ();
 sg13g2_fill_2 FILLER_7_144 ();
 sg13g2_decap_8 FILLER_7_169 ();
 sg13g2_fill_1 FILLER_7_176 ();
 sg13g2_fill_2 FILLER_7_185 ();
 sg13g2_fill_1 FILLER_7_227 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_274 ();
 sg13g2_fill_1 FILLER_7_356 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_4 FILLER_8_47 ();
 sg13g2_fill_1 FILLER_8_51 ();
 sg13g2_decap_4 FILLER_8_92 ();
 sg13g2_decap_8 FILLER_8_106 ();
 sg13g2_fill_1 FILLER_8_113 ();
 sg13g2_fill_2 FILLER_8_124 ();
 sg13g2_decap_4 FILLER_8_183 ();
 sg13g2_fill_1 FILLER_8_233 ();
 sg13g2_fill_1 FILLER_8_262 ();
 sg13g2_fill_2 FILLER_8_315 ();
 sg13g2_fill_1 FILLER_8_330 ();
 sg13g2_fill_1 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_28 ();
 sg13g2_fill_1 FILLER_9_72 ();
 sg13g2_fill_2 FILLER_9_84 ();
 sg13g2_fill_1 FILLER_9_132 ();
 sg13g2_decap_4 FILLER_9_154 ();
 sg13g2_fill_1 FILLER_9_194 ();
 sg13g2_fill_1 FILLER_9_222 ();
 sg13g2_fill_1 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_4 FILLER_10_21 ();
 sg13g2_fill_2 FILLER_10_57 ();
 sg13g2_fill_2 FILLER_10_128 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_fill_1 FILLER_10_177 ();
 sg13g2_fill_1 FILLER_10_206 ();
 sg13g2_fill_1 FILLER_10_226 ();
 sg13g2_fill_1 FILLER_10_242 ();
 sg13g2_fill_2 FILLER_10_252 ();
 sg13g2_fill_1 FILLER_10_289 ();
 sg13g2_fill_2 FILLER_10_299 ();
 sg13g2_fill_1 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_35 ();
 sg13g2_fill_2 FILLER_11_62 ();
 sg13g2_fill_1 FILLER_11_96 ();
 sg13g2_decap_4 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_fill_1 FILLER_11_294 ();
 sg13g2_fill_1 FILLER_11_348 ();
 sg13g2_fill_1 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_fill_2 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_45 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_fill_2 FILLER_12_59 ();
 sg13g2_fill_1 FILLER_12_88 ();
 sg13g2_fill_2 FILLER_12_124 ();
 sg13g2_decap_4 FILLER_12_185 ();
 sg13g2_decap_4 FILLER_12_223 ();
 sg13g2_fill_2 FILLER_12_241 ();
 sg13g2_fill_1 FILLER_12_243 ();
 sg13g2_fill_1 FILLER_12_258 ();
 sg13g2_fill_2 FILLER_12_298 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_35 ();
 sg13g2_fill_1 FILLER_13_37 ();
 sg13g2_fill_1 FILLER_13_85 ();
 sg13g2_fill_2 FILLER_13_93 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_fill_2 FILLER_13_126 ();
 sg13g2_fill_1 FILLER_13_128 ();
 sg13g2_decap_4 FILLER_13_175 ();
 sg13g2_fill_1 FILLER_13_188 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_fill_1 FILLER_13_217 ();
 sg13g2_fill_2 FILLER_13_258 ();
 sg13g2_fill_1 FILLER_13_260 ();
 sg13g2_fill_2 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_fill_1 FILLER_13_323 ();
 sg13g2_fill_2 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_21 ();
 sg13g2_fill_1 FILLER_14_23 ();
 sg13g2_fill_2 FILLER_14_55 ();
 sg13g2_fill_1 FILLER_14_57 ();
 sg13g2_fill_2 FILLER_14_89 ();
 sg13g2_fill_1 FILLER_14_91 ();
 sg13g2_fill_1 FILLER_14_118 ();
 sg13g2_decap_8 FILLER_14_138 ();
 sg13g2_decap_8 FILLER_14_145 ();
 sg13g2_decap_4 FILLER_14_152 ();
 sg13g2_fill_2 FILLER_14_160 ();
 sg13g2_fill_1 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_195 ();
 sg13g2_fill_2 FILLER_14_223 ();
 sg13g2_fill_1 FILLER_14_225 ();
 sg13g2_fill_1 FILLER_14_261 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_28 ();
 sg13g2_fill_2 FILLER_15_59 ();
 sg13g2_fill_2 FILLER_15_84 ();
 sg13g2_fill_1 FILLER_15_132 ();
 sg13g2_fill_1 FILLER_15_141 ();
 sg13g2_fill_1 FILLER_15_256 ();
 sg13g2_fill_1 FILLER_15_314 ();
 sg13g2_fill_2 FILLER_15_348 ();
 sg13g2_fill_1 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_88 ();
 sg13g2_fill_1 FILLER_16_95 ();
 sg13g2_fill_2 FILLER_16_108 ();
 sg13g2_fill_1 FILLER_16_110 ();
 sg13g2_fill_1 FILLER_16_159 ();
 sg13g2_fill_2 FILLER_16_220 ();
 sg13g2_fill_1 FILLER_16_222 ();
 sg13g2_fill_1 FILLER_16_267 ();
 sg13g2_fill_1 FILLER_16_314 ();
 sg13g2_fill_1 FILLER_16_348 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_23 ();
 sg13g2_fill_1 FILLER_17_86 ();
 sg13g2_fill_2 FILLER_17_122 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_decap_4 FILLER_17_184 ();
 sg13g2_fill_2 FILLER_17_188 ();
 sg13g2_decap_4 FILLER_17_193 ();
 sg13g2_fill_1 FILLER_17_197 ();
 sg13g2_decap_8 FILLER_17_213 ();
 sg13g2_fill_2 FILLER_17_229 ();
 sg13g2_fill_2 FILLER_17_310 ();
 sg13g2_fill_1 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_339 ();
 sg13g2_decap_4 FILLER_17_346 ();
 sg13g2_fill_1 FILLER_17_366 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_47 ();
 sg13g2_fill_1 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_72 ();
 sg13g2_decap_4 FILLER_18_79 ();
 sg13g2_fill_2 FILLER_18_83 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_184 ();
 sg13g2_fill_2 FILLER_18_215 ();
 sg13g2_decap_4 FILLER_18_220 ();
 sg13g2_fill_1 FILLER_18_229 ();
 sg13g2_fill_2 FILLER_18_274 ();
 sg13g2_decap_4 FILLER_18_307 ();
 sg13g2_fill_2 FILLER_18_337 ();
 sg13g2_fill_1 FILLER_18_339 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_57 ();
 sg13g2_fill_1 FILLER_19_85 ();
 sg13g2_fill_2 FILLER_19_127 ();
 sg13g2_fill_1 FILLER_19_140 ();
 sg13g2_fill_2 FILLER_19_170 ();
 sg13g2_decap_8 FILLER_19_257 ();
 sg13g2_fill_2 FILLER_19_264 ();
 sg13g2_decap_4 FILLER_19_315 ();
 sg13g2_fill_2 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_1 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_34 ();
 sg13g2_fill_2 FILLER_20_41 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_4 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_96 ();
 sg13g2_decap_8 FILLER_20_103 ();
 sg13g2_decap_8 FILLER_20_110 ();
 sg13g2_fill_2 FILLER_20_117 ();
 sg13g2_fill_1 FILLER_20_119 ();
 sg13g2_decap_4 FILLER_20_146 ();
 sg13g2_fill_1 FILLER_20_179 ();
 sg13g2_fill_2 FILLER_20_196 ();
 sg13g2_fill_1 FILLER_20_213 ();
 sg13g2_fill_1 FILLER_20_240 ();
 sg13g2_decap_4 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_79 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_fill_2 FILLER_21_160 ();
 sg13g2_fill_1 FILLER_21_162 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_fill_1 FILLER_21_179 ();
 sg13g2_decap_4 FILLER_21_186 ();
 sg13g2_fill_1 FILLER_21_239 ();
 sg13g2_fill_2 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_fill_2 FILLER_21_334 ();
 sg13g2_fill_1 FILLER_21_336 ();
 sg13g2_fill_1 FILLER_21_358 ();
 sg13g2_fill_2 FILLER_21_373 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_169 ();
 sg13g2_fill_2 FILLER_22_186 ();
 sg13g2_fill_1 FILLER_22_203 ();
 sg13g2_fill_2 FILLER_22_211 ();
 sg13g2_fill_1 FILLER_22_213 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_decap_4 FILLER_22_267 ();
 sg13g2_fill_2 FILLER_22_338 ();
 sg13g2_fill_2 FILLER_22_350 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_fill_2 FILLER_22_375 ();
 sg13g2_fill_1 FILLER_22_377 ();
 sg13g2_fill_1 FILLER_22_398 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_18 ();
 sg13g2_fill_1 FILLER_23_60 ();
 sg13g2_fill_2 FILLER_23_107 ();
 sg13g2_fill_1 FILLER_23_123 ();
 sg13g2_fill_2 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_decap_4 FILLER_23_190 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_280 ();
 sg13g2_fill_2 FILLER_23_341 ();
 sg13g2_fill_2 FILLER_23_373 ();
 sg13g2_fill_1 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_23 ();
 sg13g2_fill_2 FILLER_24_41 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_97 ();
 sg13g2_fill_2 FILLER_24_103 ();
 sg13g2_decap_4 FILLER_24_135 ();
 sg13g2_fill_1 FILLER_24_162 ();
 sg13g2_fill_2 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_fill_1 FILLER_24_291 ();
 sg13g2_fill_1 FILLER_24_316 ();
 sg13g2_fill_2 FILLER_24_358 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_fill_2 FILLER_24_366 ();
 sg13g2_fill_2 FILLER_24_380 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_4 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_77 ();
 sg13g2_fill_2 FILLER_25_107 ();
 sg13g2_fill_1 FILLER_25_109 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_169 ();
 sg13g2_fill_2 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_188 ();
 sg13g2_fill_1 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_257 ();
 sg13g2_fill_2 FILLER_25_293 ();
 sg13g2_fill_2 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_fill_2 FILLER_26_21 ();
 sg13g2_fill_1 FILLER_26_23 ();
 sg13g2_fill_1 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_111 ();
 sg13g2_fill_1 FILLER_26_133 ();
 sg13g2_fill_1 FILLER_26_143 ();
 sg13g2_fill_1 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_decap_8 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_decap_4 FILLER_26_217 ();
 sg13g2_fill_2 FILLER_26_230 ();
 sg13g2_fill_2 FILLER_26_236 ();
 sg13g2_fill_2 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_fill_2 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_128 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_decap_4 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_fill_2 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_34 ();
 sg13g2_fill_2 FILLER_28_41 ();
 sg13g2_fill_1 FILLER_28_43 ();
 sg13g2_decap_8 FILLER_28_50 ();
 sg13g2_decap_4 FILLER_28_57 ();
 sg13g2_fill_2 FILLER_28_66 ();
 sg13g2_fill_2 FILLER_28_94 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_decap_4 FILLER_28_210 ();
 sg13g2_fill_2 FILLER_28_318 ();
 sg13g2_decap_4 FILLER_28_330 ();
 sg13g2_fill_2 FILLER_28_334 ();
 sg13g2_fill_1 FILLER_28_374 ();
 sg13g2_fill_2 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_382 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_4 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_32 ();
 sg13g2_decap_8 FILLER_29_38 ();
 sg13g2_decap_8 FILLER_29_45 ();
 sg13g2_fill_1 FILLER_29_55 ();
 sg13g2_fill_2 FILLER_29_68 ();
 sg13g2_decap_4 FILLER_29_97 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_decap_4 FILLER_29_168 ();
 sg13g2_fill_2 FILLER_29_172 ();
 sg13g2_fill_2 FILLER_29_220 ();
 sg13g2_fill_1 FILLER_29_297 ();
 sg13g2_fill_2 FILLER_29_332 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_18 ();
 sg13g2_decap_8 FILLER_30_94 ();
 sg13g2_fill_1 FILLER_30_101 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_190 ();
 sg13g2_fill_2 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_284 ();
 sg13g2_fill_2 FILLER_30_330 ();
 sg13g2_fill_2 FILLER_30_374 ();
 sg13g2_fill_2 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_75 ();
 sg13g2_fill_1 FILLER_31_86 ();
 sg13g2_fill_2 FILLER_31_92 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_130 ();
 sg13g2_fill_2 FILLER_31_153 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_decap_8 FILLER_31_169 ();
 sg13g2_decap_8 FILLER_31_176 ();
 sg13g2_decap_8 FILLER_31_183 ();
 sg13g2_fill_2 FILLER_31_195 ();
 sg13g2_fill_1 FILLER_31_207 ();
 sg13g2_fill_1 FILLER_31_230 ();
 sg13g2_fill_2 FILLER_31_244 ();
 sg13g2_fill_1 FILLER_31_246 ();
 sg13g2_decap_4 FILLER_31_256 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_277 ();
 sg13g2_fill_1 FILLER_31_312 ();
 sg13g2_fill_2 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_18 ();
 sg13g2_fill_1 FILLER_32_46 ();
 sg13g2_fill_1 FILLER_32_74 ();
 sg13g2_fill_1 FILLER_32_83 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_167 ();
 sg13g2_fill_2 FILLER_32_177 ();
 sg13g2_fill_2 FILLER_32_199 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_fill_2 FILLER_32_237 ();
 sg13g2_decap_4 FILLER_32_259 ();
 sg13g2_fill_2 FILLER_32_263 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_fill_2 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_282 ();
 sg13g2_fill_2 FILLER_32_297 ();
 sg13g2_fill_1 FILLER_32_308 ();
 sg13g2_fill_1 FILLER_32_318 ();
 sg13g2_fill_1 FILLER_32_338 ();
 sg13g2_fill_2 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_360 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_11 ();
 sg13g2_fill_2 FILLER_33_36 ();
 sg13g2_fill_2 FILLER_33_60 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_fill_2 FILLER_33_139 ();
 sg13g2_fill_2 FILLER_33_155 ();
 sg13g2_decap_4 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_236 ();
 sg13g2_fill_2 FILLER_33_246 ();
 sg13g2_fill_1 FILLER_33_253 ();
 sg13g2_decap_4 FILLER_33_292 ();
 sg13g2_fill_2 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_330 ();
 sg13g2_fill_2 FILLER_33_358 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_fill_2 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_18 ();
 sg13g2_fill_1 FILLER_34_78 ();
 sg13g2_fill_2 FILLER_34_94 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_fill_2 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_4 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_25 ();
 sg13g2_fill_1 FILLER_35_32 ();
 sg13g2_fill_2 FILLER_35_99 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_1 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_215 ();
 sg13g2_decap_8 FILLER_35_222 ();
 sg13g2_decap_8 FILLER_35_229 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_fill_1 FILLER_35_282 ();
 sg13g2_fill_2 FILLER_35_288 ();
 sg13g2_fill_1 FILLER_35_290 ();
 sg13g2_decap_8 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_35_333 ();
 sg13g2_fill_1 FILLER_35_340 ();
 sg13g2_fill_1 FILLER_35_363 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_28 ();
 sg13g2_fill_1 FILLER_36_32 ();
 sg13g2_fill_2 FILLER_36_41 ();
 sg13g2_fill_1 FILLER_36_87 ();
 sg13g2_fill_1 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_decap_4 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_2 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_fill_1 FILLER_36_314 ();
 sg13g2_decap_8 FILLER_36_327 ();
 sg13g2_decap_8 FILLER_36_334 ();
 sg13g2_fill_1 FILLER_36_341 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_4 FILLER_37_21 ();
 sg13g2_decap_4 FILLER_37_58 ();
 sg13g2_fill_1 FILLER_37_62 ();
 sg13g2_fill_2 FILLER_37_68 ();
 sg13g2_fill_1 FILLER_37_120 ();
 sg13g2_fill_2 FILLER_37_189 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_fill_2 FILLER_37_247 ();
 sg13g2_fill_1 FILLER_37_249 ();
 sg13g2_fill_1 FILLER_37_297 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_fill_1 FILLER_37_313 ();
 sg13g2_decap_4 FILLER_37_340 ();
 sg13g2_decap_8 FILLER_37_348 ();
 sg13g2_decap_4 FILLER_37_355 ();
 sg13g2_fill_1 FILLER_37_359 ();
 sg13g2_decap_4 FILLER_38_26 ();
 sg13g2_fill_1 FILLER_38_30 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_fill_2 FILLER_38_64 ();
 sg13g2_fill_1 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_124 ();
 sg13g2_fill_2 FILLER_38_181 ();
 sg13g2_fill_1 FILLER_38_197 ();
 sg13g2_fill_2 FILLER_38_256 ();
 sg13g2_fill_2 FILLER_38_322 ();
 sg13g2_fill_2 FILLER_38_362 ();
 sg13g2_fill_1 FILLER_38_364 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_1 FILLER_39_59 ();
 sg13g2_fill_1 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_106 ();
 sg13g2_decap_4 FILLER_39_113 ();
 sg13g2_fill_1 FILLER_39_121 ();
 sg13g2_fill_2 FILLER_39_151 ();
 sg13g2_fill_1 FILLER_39_179 ();
 sg13g2_decap_4 FILLER_39_218 ();
 sg13g2_fill_2 FILLER_39_222 ();
 sg13g2_fill_2 FILLER_39_233 ();
 sg13g2_fill_1 FILLER_39_241 ();
 sg13g2_fill_2 FILLER_39_258 ();
 sg13g2_fill_1 FILLER_39_377 ();
 sg13g2_fill_2 FILLER_39_383 ();
 sg13g2_fill_1 FILLER_39_385 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_4 ();
 sg13g2_fill_2 FILLER_40_24 ();
 sg13g2_fill_1 FILLER_40_44 ();
 sg13g2_fill_1 FILLER_40_59 ();
 sg13g2_fill_1 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_80 ();
 sg13g2_decap_8 FILLER_40_87 ();
 sg13g2_decap_8 FILLER_40_94 ();
 sg13g2_decap_8 FILLER_40_101 ();
 sg13g2_decap_8 FILLER_40_108 ();
 sg13g2_decap_8 FILLER_40_115 ();
 sg13g2_decap_8 FILLER_40_122 ();
 sg13g2_decap_8 FILLER_40_129 ();
 sg13g2_decap_4 FILLER_40_136 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_fill_2 FILLER_40_175 ();
 sg13g2_fill_1 FILLER_40_177 ();
 sg13g2_decap_8 FILLER_40_190 ();
 sg13g2_decap_8 FILLER_40_197 ();
 sg13g2_fill_2 FILLER_40_204 ();
 sg13g2_fill_1 FILLER_40_206 ();
 sg13g2_fill_2 FILLER_40_216 ();
 sg13g2_fill_2 FILLER_40_221 ();
 sg13g2_decap_8 FILLER_40_229 ();
 sg13g2_decap_4 FILLER_40_236 ();
 sg13g2_fill_2 FILLER_40_240 ();
 sg13g2_fill_2 FILLER_40_297 ();
 sg13g2_fill_1 FILLER_40_299 ();
 sg13g2_fill_2 FILLER_40_318 ();
 sg13g2_fill_1 FILLER_40_320 ();
 sg13g2_fill_1 FILLER_40_398 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_21 ();
 sg13g2_fill_2 FILLER_41_98 ();
 sg13g2_fill_1 FILLER_41_106 ();
 sg13g2_fill_1 FILLER_41_110 ();
 sg13g2_decap_8 FILLER_41_115 ();
 sg13g2_decap_8 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_129 ();
 sg13g2_decap_8 FILLER_41_136 ();
 sg13g2_fill_2 FILLER_41_143 ();
 sg13g2_decap_8 FILLER_41_149 ();
 sg13g2_fill_2 FILLER_41_156 ();
 sg13g2_decap_8 FILLER_41_163 ();
 sg13g2_decap_8 FILLER_41_170 ();
 sg13g2_fill_1 FILLER_41_177 ();
 sg13g2_decap_8 FILLER_41_215 ();
 sg13g2_fill_1 FILLER_41_222 ();
 sg13g2_decap_4 FILLER_41_238 ();
 sg13g2_fill_2 FILLER_41_242 ();
 sg13g2_fill_1 FILLER_41_256 ();
 sg13g2_decap_4 FILLER_41_264 ();
 sg13g2_fill_1 FILLER_41_268 ();
 sg13g2_decap_4 FILLER_41_288 ();
 sg13g2_decap_8 FILLER_41_302 ();
 sg13g2_fill_2 FILLER_41_327 ();
 sg13g2_fill_2 FILLER_41_357 ();
 sg13g2_fill_1 FILLER_41_368 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_4 ();
 sg13g2_fill_1 FILLER_42_31 ();
 sg13g2_fill_1 FILLER_42_41 ();
 sg13g2_fill_2 FILLER_42_51 ();
 sg13g2_fill_1 FILLER_42_53 ();
 sg13g2_fill_2 FILLER_42_94 ();
 sg13g2_fill_1 FILLER_42_100 ();
 sg13g2_fill_1 FILLER_42_117 ();
 sg13g2_decap_4 FILLER_42_152 ();
 sg13g2_decap_8 FILLER_42_173 ();
 sg13g2_decap_8 FILLER_42_180 ();
 sg13g2_fill_2 FILLER_42_187 ();
 sg13g2_fill_1 FILLER_42_189 ();
 sg13g2_decap_4 FILLER_42_204 ();
 sg13g2_fill_1 FILLER_42_208 ();
 sg13g2_fill_1 FILLER_42_225 ();
 sg13g2_fill_2 FILLER_42_235 ();
 sg13g2_fill_2 FILLER_42_274 ();
 sg13g2_fill_1 FILLER_42_276 ();
 sg13g2_fill_2 FILLER_42_330 ();
 sg13g2_fill_1 FILLER_42_332 ();
 sg13g2_fill_1 FILLER_42_361 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_4 FILLER_43_68 ();
 sg13g2_fill_2 FILLER_43_72 ();
 sg13g2_fill_1 FILLER_43_83 ();
 sg13g2_fill_1 FILLER_43_162 ();
 sg13g2_fill_2 FILLER_43_169 ();
 sg13g2_fill_1 FILLER_43_171 ();
 sg13g2_fill_2 FILLER_43_180 ();
 sg13g2_fill_2 FILLER_43_242 ();
 sg13g2_fill_1 FILLER_43_283 ();
 sg13g2_fill_1 FILLER_43_312 ();
 sg13g2_fill_2 FILLER_43_362 ();
 sg13g2_fill_1 FILLER_43_399 ();
 sg13g2_fill_1 FILLER_44_26 ();
 sg13g2_decap_8 FILLER_44_64 ();
 sg13g2_decap_8 FILLER_44_71 ();
 sg13g2_fill_2 FILLER_44_116 ();
 sg13g2_fill_1 FILLER_44_144 ();
 sg13g2_fill_2 FILLER_44_158 ();
 sg13g2_fill_1 FILLER_44_160 ();
 sg13g2_decap_4 FILLER_44_175 ();
 sg13g2_fill_2 FILLER_44_270 ();
 sg13g2_fill_1 FILLER_44_272 ();
 sg13g2_fill_2 FILLER_44_299 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_56 ();
 sg13g2_fill_1 FILLER_45_62 ();
 sg13g2_decap_4 FILLER_45_72 ();
 sg13g2_fill_2 FILLER_45_76 ();
 sg13g2_fill_1 FILLER_45_111 ();
 sg13g2_fill_2 FILLER_45_153 ();
 sg13g2_fill_2 FILLER_45_241 ();
 sg13g2_fill_1 FILLER_45_243 ();
 sg13g2_fill_2 FILLER_45_296 ();
 sg13g2_fill_1 FILLER_45_298 ();
 sg13g2_fill_1 FILLER_45_382 ();
 sg13g2_fill_2 FILLER_46_59 ();
 sg13g2_fill_2 FILLER_46_80 ();
 sg13g2_decap_4 FILLER_46_87 ();
 sg13g2_fill_2 FILLER_46_116 ();
 sg13g2_decap_8 FILLER_46_145 ();
 sg13g2_fill_1 FILLER_46_152 ();
 sg13g2_decap_4 FILLER_46_157 ();
 sg13g2_fill_1 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_167 ();
 sg13g2_fill_2 FILLER_46_174 ();
 sg13g2_fill_1 FILLER_46_176 ();
 sg13g2_fill_1 FILLER_46_194 ();
 sg13g2_fill_2 FILLER_46_204 ();
 sg13g2_fill_2 FILLER_46_211 ();
 sg13g2_fill_1 FILLER_46_230 ();
 sg13g2_fill_2 FILLER_46_267 ();
 sg13g2_fill_1 FILLER_46_269 ();
 sg13g2_fill_2 FILLER_46_286 ();
 sg13g2_fill_1 FILLER_46_288 ();
 sg13g2_fill_1 FILLER_46_303 ();
 sg13g2_fill_1 FILLER_47_26 ();
 sg13g2_fill_1 FILLER_47_108 ();
 sg13g2_fill_1 FILLER_47_181 ();
 sg13g2_fill_1 FILLER_47_252 ();
 sg13g2_fill_2 FILLER_47_262 ();
 sg13g2_fill_1 FILLER_47_264 ();
 sg13g2_fill_2 FILLER_47_312 ();
 sg13g2_fill_1 FILLER_47_323 ();
 sg13g2_fill_1 FILLER_47_342 ();
 sg13g2_fill_1 FILLER_47_363 ();
 sg13g2_fill_1 FILLER_47_382 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_7 ();
 sg13g2_fill_1 FILLER_48_9 ();
 sg13g2_fill_2 FILLER_48_46 ();
 sg13g2_fill_1 FILLER_48_68 ();
 sg13g2_fill_1 FILLER_48_78 ();
 sg13g2_fill_2 FILLER_48_102 ();
 sg13g2_fill_1 FILLER_48_143 ();
 sg13g2_fill_1 FILLER_48_164 ();
 sg13g2_fill_1 FILLER_48_234 ();
 sg13g2_fill_1 FILLER_48_261 ();
 sg13g2_fill_2 FILLER_48_317 ();
 sg13g2_fill_1 FILLER_48_362 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_48 ();
 sg13g2_fill_1 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_112 ();
 sg13g2_fill_1 FILLER_49_119 ();
 sg13g2_fill_1 FILLER_49_150 ();
 sg13g2_fill_2 FILLER_49_172 ();
 sg13g2_fill_2 FILLER_49_183 ();
 sg13g2_fill_1 FILLER_49_185 ();
 sg13g2_fill_1 FILLER_49_264 ();
 sg13g2_fill_2 FILLER_49_319 ();
 sg13g2_fill_1 FILLER_49_321 ();
 sg13g2_fill_2 FILLER_49_339 ();
 sg13g2_fill_1 FILLER_49_341 ();
 sg13g2_fill_2 FILLER_49_359 ();
 sg13g2_fill_1 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_38 ();
 sg13g2_fill_1 FILLER_50_105 ();
 sg13g2_fill_2 FILLER_50_134 ();
 sg13g2_fill_2 FILLER_50_151 ();
 sg13g2_fill_2 FILLER_50_161 ();
 sg13g2_decap_4 FILLER_50_168 ();
 sg13g2_fill_1 FILLER_50_179 ();
 sg13g2_fill_1 FILLER_50_190 ();
 sg13g2_fill_1 FILLER_50_212 ();
 sg13g2_fill_1 FILLER_50_218 ();
 sg13g2_decap_8 FILLER_50_264 ();
 sg13g2_decap_4 FILLER_50_271 ();
 sg13g2_fill_2 FILLER_50_275 ();
 sg13g2_fill_1 FILLER_50_315 ();
 sg13g2_fill_2 FILLER_50_383 ();
 sg13g2_fill_1 FILLER_50_385 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_4 FILLER_51_21 ();
 sg13g2_fill_2 FILLER_51_25 ();
 sg13g2_fill_2 FILLER_51_77 ();
 sg13g2_fill_2 FILLER_51_93 ();
 sg13g2_fill_2 FILLER_51_120 ();
 sg13g2_fill_1 FILLER_51_156 ();
 sg13g2_decap_8 FILLER_51_165 ();
 sg13g2_decap_8 FILLER_51_172 ();
 sg13g2_decap_8 FILLER_51_179 ();
 sg13g2_fill_2 FILLER_51_186 ();
 sg13g2_fill_1 FILLER_51_188 ();
 sg13g2_fill_1 FILLER_51_202 ();
 sg13g2_fill_2 FILLER_51_227 ();
 sg13g2_fill_2 FILLER_51_282 ();
 sg13g2_fill_1 FILLER_51_284 ();
 sg13g2_fill_1 FILLER_51_314 ();
 sg13g2_fill_2 FILLER_51_351 ();
 sg13g2_fill_2 FILLER_51_397 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_4 FILLER_52_21 ();
 sg13g2_fill_2 FILLER_52_25 ();
 sg13g2_fill_1 FILLER_52_40 ();
 sg13g2_fill_2 FILLER_52_52 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_fill_1 FILLER_52_116 ();
 sg13g2_fill_2 FILLER_52_136 ();
 sg13g2_fill_2 FILLER_52_164 ();
 sg13g2_fill_1 FILLER_52_175 ();
 sg13g2_fill_1 FILLER_52_183 ();
 sg13g2_fill_2 FILLER_52_229 ();
 sg13g2_decap_4 FILLER_52_267 ();
 sg13g2_fill_1 FILLER_52_271 ();
 sg13g2_fill_2 FILLER_52_312 ();
 sg13g2_decap_8 FILLER_52_338 ();
 sg13g2_decap_4 FILLER_52_345 ();
 sg13g2_fill_2 FILLER_52_349 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_4 FILLER_53_14 ();
 sg13g2_fill_2 FILLER_53_66 ();
 sg13g2_fill_1 FILLER_53_78 ();
 sg13g2_fill_1 FILLER_53_165 ();
 sg13g2_fill_2 FILLER_53_176 ();
 sg13g2_fill_1 FILLER_53_178 ();
 sg13g2_fill_1 FILLER_53_222 ();
 sg13g2_fill_1 FILLER_53_263 ();
 sg13g2_fill_1 FILLER_53_290 ();
 sg13g2_fill_2 FILLER_53_296 ();
 sg13g2_fill_1 FILLER_53_298 ();
 sg13g2_fill_2 FILLER_53_329 ();
 sg13g2_fill_2 FILLER_53_354 ();
 sg13g2_fill_1 FILLER_53_356 ();
 sg13g2_fill_2 FILLER_53_384 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_7 ();
 sg13g2_fill_1 FILLER_54_9 ();
 sg13g2_fill_1 FILLER_54_36 ();
 sg13g2_fill_2 FILLER_54_71 ();
 sg13g2_decap_4 FILLER_54_96 ();
 sg13g2_fill_1 FILLER_54_100 ();
 sg13g2_fill_1 FILLER_54_106 ();
 sg13g2_decap_4 FILLER_54_114 ();
 sg13g2_fill_2 FILLER_54_118 ();
 sg13g2_fill_2 FILLER_54_128 ();
 sg13g2_fill_2 FILLER_54_138 ();
 sg13g2_fill_2 FILLER_54_149 ();
 sg13g2_fill_1 FILLER_54_170 ();
 sg13g2_fill_2 FILLER_54_195 ();
 sg13g2_fill_2 FILLER_54_213 ();
 sg13g2_fill_2 FILLER_54_220 ();
 sg13g2_fill_1 FILLER_54_227 ();
 sg13g2_fill_2 FILLER_54_334 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_4 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_37 ();
 sg13g2_fill_2 FILLER_55_73 ();
 sg13g2_decap_8 FILLER_55_118 ();
 sg13g2_fill_2 FILLER_55_149 ();
 sg13g2_fill_2 FILLER_55_183 ();
 sg13g2_fill_1 FILLER_55_235 ();
 sg13g2_fill_1 FILLER_55_275 ();
 sg13g2_fill_2 FILLER_55_346 ();
 sg13g2_fill_1 FILLER_55_348 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_37 ();
 sg13g2_decap_4 FILLER_56_59 ();
 sg13g2_fill_2 FILLER_56_63 ();
 sg13g2_decap_4 FILLER_56_95 ();
 sg13g2_fill_2 FILLER_56_99 ();
 sg13g2_fill_1 FILLER_56_106 ();
 sg13g2_fill_1 FILLER_56_188 ();
 sg13g2_fill_2 FILLER_56_228 ();
 sg13g2_fill_2 FILLER_56_235 ();
 sg13g2_decap_4 FILLER_56_253 ();
 sg13g2_fill_1 FILLER_56_257 ();
 sg13g2_decap_8 FILLER_56_271 ();
 sg13g2_fill_2 FILLER_56_278 ();
 sg13g2_fill_1 FILLER_56_307 ();
 sg13g2_fill_2 FILLER_56_355 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_fill_2 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_16 ();
 sg13g2_decap_4 FILLER_57_30 ();
 sg13g2_fill_2 FILLER_57_42 ();
 sg13g2_fill_1 FILLER_57_44 ();
 sg13g2_decap_8 FILLER_57_55 ();
 sg13g2_decap_8 FILLER_57_62 ();
 sg13g2_fill_1 FILLER_57_88 ();
 sg13g2_fill_1 FILLER_57_127 ();
 sg13g2_fill_2 FILLER_57_174 ();
 sg13g2_fill_1 FILLER_57_224 ();
 sg13g2_decap_8 FILLER_57_246 ();
 sg13g2_decap_8 FILLER_57_253 ();
 sg13g2_fill_2 FILLER_57_260 ();
 sg13g2_fill_1 FILLER_57_262 ();
 sg13g2_fill_2 FILLER_57_327 ();
 sg13g2_fill_1 FILLER_57_329 ();
 sg13g2_fill_1 FILLER_57_372 ();
 sg13g2_fill_1 FILLER_57_399 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_61 ();
 sg13g2_decap_4 FILLER_58_68 ();
 sg13g2_fill_1 FILLER_58_72 ();
 sg13g2_decap_4 FILLER_58_99 ();
 sg13g2_decap_8 FILLER_58_167 ();
 sg13g2_fill_2 FILLER_58_174 ();
 sg13g2_fill_1 FILLER_58_216 ();
 sg13g2_fill_2 FILLER_58_260 ();
 sg13g2_fill_2 FILLER_58_292 ();
 sg13g2_fill_1 FILLER_58_330 ();
 sg13g2_fill_1 FILLER_58_340 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_72 ();
 sg13g2_decap_4 FILLER_59_79 ();
 sg13g2_fill_1 FILLER_59_83 ();
 sg13g2_fill_2 FILLER_59_118 ();
 sg13g2_fill_1 FILLER_59_134 ();
 sg13g2_decap_4 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_162 ();
 sg13g2_decap_8 FILLER_59_169 ();
 sg13g2_decap_4 FILLER_59_176 ();
 sg13g2_decap_4 FILLER_59_184 ();
 sg13g2_fill_1 FILLER_59_188 ();
 sg13g2_fill_1 FILLER_59_223 ();
 sg13g2_fill_2 FILLER_59_300 ();
 sg13g2_fill_1 FILLER_59_346 ();
 sg13g2_fill_1 FILLER_59_373 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_92 ();
 sg13g2_fill_2 FILLER_60_99 ();
 sg13g2_fill_1 FILLER_60_101 ();
 sg13g2_fill_1 FILLER_60_107 ();
 sg13g2_decap_8 FILLER_60_129 ();
 sg13g2_fill_2 FILLER_60_136 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_fill_2 FILLER_60_162 ();
 sg13g2_decap_4 FILLER_60_191 ();
 sg13g2_fill_1 FILLER_60_195 ();
 sg13g2_fill_1 FILLER_60_217 ();
 sg13g2_decap_8 FILLER_60_246 ();
 sg13g2_decap_8 FILLER_60_253 ();
 sg13g2_decap_8 FILLER_60_260 ();
 sg13g2_fill_1 FILLER_60_267 ();
 sg13g2_fill_1 FILLER_60_373 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_4 FILLER_61_14 ();
 sg13g2_fill_2 FILLER_61_18 ();
 sg13g2_fill_1 FILLER_61_24 ();
 sg13g2_fill_1 FILLER_61_44 ();
 sg13g2_fill_2 FILLER_61_133 ();
 sg13g2_fill_1 FILLER_61_135 ();
 sg13g2_fill_1 FILLER_61_154 ();
 sg13g2_fill_2 FILLER_61_190 ();
 sg13g2_decap_4 FILLER_61_204 ();
 sg13g2_fill_2 FILLER_61_208 ();
 sg13g2_fill_2 FILLER_61_239 ();
 sg13g2_fill_2 FILLER_61_302 ();
 sg13g2_fill_1 FILLER_61_304 ();
 sg13g2_fill_2 FILLER_61_318 ();
 sg13g2_fill_1 FILLER_61_333 ();
 sg13g2_fill_2 FILLER_61_361 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_4 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_46 ();
 sg13g2_decap_4 FILLER_62_85 ();
 sg13g2_fill_1 FILLER_62_89 ();
 sg13g2_fill_2 FILLER_62_125 ();
 sg13g2_fill_1 FILLER_62_127 ();
 sg13g2_fill_2 FILLER_62_132 ();
 sg13g2_fill_1 FILLER_62_169 ();
 sg13g2_fill_2 FILLER_62_190 ();
 sg13g2_decap_4 FILLER_62_256 ();
 sg13g2_fill_2 FILLER_62_260 ();
 sg13g2_fill_2 FILLER_62_276 ();
 sg13g2_fill_1 FILLER_62_303 ();
 sg13g2_fill_1 FILLER_62_342 ();
 sg13g2_fill_1 FILLER_62_353 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_4 FILLER_63_21 ();
 sg13g2_fill_1 FILLER_63_25 ();
 sg13g2_fill_1 FILLER_63_66 ();
 sg13g2_fill_2 FILLER_63_117 ();
 sg13g2_fill_1 FILLER_63_119 ();
 sg13g2_fill_2 FILLER_63_136 ();
 sg13g2_fill_1 FILLER_63_272 ();
 sg13g2_fill_2 FILLER_63_299 ();
 sg13g2_fill_1 FILLER_63_301 ();
 sg13g2_fill_2 FILLER_63_342 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_14 ();
 sg13g2_fill_2 FILLER_64_28 ();
 sg13g2_fill_1 FILLER_64_51 ();
 sg13g2_fill_1 FILLER_64_78 ();
 sg13g2_fill_1 FILLER_64_110 ();
 sg13g2_fill_1 FILLER_64_162 ();
 sg13g2_fill_2 FILLER_64_366 ();
 sg13g2_fill_2 FILLER_64_384 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_7 ();
 sg13g2_decap_4 FILLER_65_43 ();
 sg13g2_fill_2 FILLER_65_65 ();
 sg13g2_decap_8 FILLER_65_85 ();
 sg13g2_fill_2 FILLER_65_92 ();
 sg13g2_fill_1 FILLER_65_94 ();
 sg13g2_fill_2 FILLER_65_113 ();
 sg13g2_fill_1 FILLER_65_131 ();
 sg13g2_fill_1 FILLER_65_145 ();
 sg13g2_fill_2 FILLER_65_165 ();
 sg13g2_fill_1 FILLER_65_177 ();
 sg13g2_fill_2 FILLER_65_210 ();
 sg13g2_decap_4 FILLER_65_233 ();
 sg13g2_fill_1 FILLER_65_237 ();
 sg13g2_fill_1 FILLER_65_242 ();
 sg13g2_fill_2 FILLER_65_287 ();
 sg13g2_fill_2 FILLER_65_298 ();
 sg13g2_fill_1 FILLER_65_347 ();
 sg13g2_fill_1 FILLER_65_371 ();
 sg13g2_fill_1 FILLER_65_387 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_75 ();
 sg13g2_decap_4 FILLER_66_82 ();
 sg13g2_fill_1 FILLER_66_86 ();
 sg13g2_fill_2 FILLER_66_113 ();
 sg13g2_fill_1 FILLER_66_145 ();
 sg13g2_fill_2 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_240 ();
 sg13g2_decap_4 FILLER_66_247 ();
 sg13g2_fill_2 FILLER_66_251 ();
 sg13g2_fill_2 FILLER_66_258 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_4 FILLER_67_14 ();
 sg13g2_fill_1 FILLER_67_28 ();
 sg13g2_fill_2 FILLER_67_38 ();
 sg13g2_fill_2 FILLER_67_139 ();
 sg13g2_fill_2 FILLER_67_167 ();
 sg13g2_fill_2 FILLER_67_345 ();
 sg13g2_fill_1 FILLER_67_347 ();
 sg13g2_fill_1 FILLER_67_358 ();
 sg13g2_fill_1 FILLER_67_392 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_21 ();
 sg13g2_fill_2 FILLER_68_101 ();
 sg13g2_fill_1 FILLER_68_103 ();
 sg13g2_fill_1 FILLER_68_125 ();
 sg13g2_fill_1 FILLER_68_182 ();
 sg13g2_fill_2 FILLER_68_228 ();
 sg13g2_fill_2 FILLER_68_339 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_14 ();
 sg13g2_fill_1 FILLER_69_102 ();
 sg13g2_decap_8 FILLER_69_185 ();
 sg13g2_decap_4 FILLER_69_192 ();
 sg13g2_fill_1 FILLER_69_268 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_7 ();
 sg13g2_fill_1 FILLER_70_11 ();
 sg13g2_fill_2 FILLER_70_43 ();
 sg13g2_fill_2 FILLER_70_68 ();
 sg13g2_fill_1 FILLER_70_80 ();
 sg13g2_fill_1 FILLER_70_95 ();
 sg13g2_fill_2 FILLER_70_111 ();
 sg13g2_fill_2 FILLER_70_180 ();
 sg13g2_decap_8 FILLER_70_191 ();
 sg13g2_decap_4 FILLER_70_198 ();
 sg13g2_fill_2 FILLER_70_202 ();
 sg13g2_fill_1 FILLER_70_221 ();
 sg13g2_decap_8 FILLER_70_249 ();
 sg13g2_decap_8 FILLER_70_256 ();
 sg13g2_decap_4 FILLER_70_263 ();
 sg13g2_fill_2 FILLER_70_267 ();
 sg13g2_fill_2 FILLER_70_278 ();
 sg13g2_fill_1 FILLER_70_280 ();
 sg13g2_fill_1 FILLER_70_344 ();
 sg13g2_fill_2 FILLER_70_381 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_4 FILLER_71_14 ();
 sg13g2_fill_1 FILLER_71_18 ();
 sg13g2_fill_1 FILLER_71_70 ();
 sg13g2_fill_2 FILLER_71_197 ();
 sg13g2_decap_4 FILLER_71_209 ();
 sg13g2_decap_8 FILLER_71_254 ();
 sg13g2_decap_4 FILLER_71_271 ();
 sg13g2_fill_2 FILLER_71_275 ();
 sg13g2_fill_1 FILLER_71_295 ();
 sg13g2_fill_2 FILLER_71_311 ();
 sg13g2_fill_2 FILLER_71_373 ();
 sg13g2_fill_1 FILLER_71_375 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_4 FILLER_72_28 ();
 sg13g2_fill_2 FILLER_72_32 ();
 sg13g2_fill_2 FILLER_72_109 ();
 sg13g2_fill_1 FILLER_72_160 ();
 sg13g2_decap_4 FILLER_72_196 ();
 sg13g2_fill_2 FILLER_72_200 ();
 sg13g2_decap_8 FILLER_72_238 ();
 sg13g2_fill_2 FILLER_72_291 ();
 sg13g2_fill_1 FILLER_72_293 ();
 sg13g2_fill_2 FILLER_72_333 ();
 sg13g2_fill_1 FILLER_72_335 ();
 sg13g2_fill_1 FILLER_72_367 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_4 FILLER_73_28 ();
 sg13g2_fill_1 FILLER_73_32 ();
 sg13g2_fill_1 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_48 ();
 sg13g2_fill_1 FILLER_73_55 ();
 sg13g2_fill_2 FILLER_73_103 ();
 sg13g2_fill_1 FILLER_73_105 ();
 sg13g2_fill_2 FILLER_73_141 ();
 sg13g2_fill_2 FILLER_73_163 ();
 sg13g2_fill_1 FILLER_73_196 ();
 sg13g2_fill_2 FILLER_73_233 ();
 sg13g2_fill_1 FILLER_73_235 ();
 sg13g2_fill_2 FILLER_73_241 ();
 sg13g2_fill_2 FILLER_73_330 ();
 sg13g2_fill_1 FILLER_73_389 ();
 sg13g2_fill_1 FILLER_73_399 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_4 FILLER_74_56 ();
 sg13g2_fill_1 FILLER_74_60 ();
 sg13g2_fill_2 FILLER_74_69 ();
 sg13g2_fill_1 FILLER_74_71 ();
 sg13g2_decap_4 FILLER_74_99 ();
 sg13g2_fill_2 FILLER_74_115 ();
 sg13g2_fill_1 FILLER_74_117 ();
 sg13g2_fill_1 FILLER_74_124 ();
 sg13g2_fill_1 FILLER_74_134 ();
 sg13g2_fill_2 FILLER_74_138 ();
 sg13g2_fill_1 FILLER_74_176 ();
 sg13g2_fill_1 FILLER_74_212 ();
 sg13g2_fill_2 FILLER_74_217 ();
 sg13g2_fill_1 FILLER_74_219 ();
 sg13g2_fill_2 FILLER_74_251 ();
 sg13g2_fill_2 FILLER_74_267 ();
 sg13g2_fill_1 FILLER_74_269 ();
 sg13g2_fill_1 FILLER_74_322 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_4 FILLER_75_66 ();
 sg13g2_fill_2 FILLER_75_70 ();
 sg13g2_fill_2 FILLER_75_89 ();
 sg13g2_fill_1 FILLER_75_91 ();
 sg13g2_fill_2 FILLER_75_103 ();
 sg13g2_decap_4 FILLER_75_110 ();
 sg13g2_fill_1 FILLER_75_179 ();
 sg13g2_decap_4 FILLER_75_209 ();
 sg13g2_fill_2 FILLER_75_213 ();
 sg13g2_decap_4 FILLER_75_229 ();
 sg13g2_fill_1 FILLER_75_233 ();
 sg13g2_fill_2 FILLER_75_253 ();
 sg13g2_fill_1 FILLER_75_255 ();
 sg13g2_decap_8 FILLER_75_260 ();
 sg13g2_decap_4 FILLER_75_267 ();
 sg13g2_fill_2 FILLER_75_275 ();
 sg13g2_decap_8 FILLER_75_291 ();
 sg13g2_fill_1 FILLER_75_368 ();
 sg13g2_fill_2 FILLER_75_379 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_4 FILLER_76_42 ();
 sg13g2_fill_1 FILLER_76_46 ();
 sg13g2_fill_2 FILLER_76_93 ();
 sg13g2_fill_1 FILLER_76_105 ();
 sg13g2_fill_2 FILLER_76_116 ();
 sg13g2_fill_1 FILLER_76_123 ();
 sg13g2_fill_1 FILLER_76_132 ();
 sg13g2_fill_1 FILLER_76_143 ();
 sg13g2_decap_8 FILLER_76_177 ();
 sg13g2_decap_8 FILLER_76_184 ();
 sg13g2_fill_2 FILLER_76_191 ();
 sg13g2_fill_1 FILLER_76_193 ();
 sg13g2_decap_8 FILLER_76_204 ();
 sg13g2_decap_8 FILLER_76_211 ();
 sg13g2_decap_8 FILLER_76_218 ();
 sg13g2_decap_4 FILLER_76_225 ();
 sg13g2_decap_8 FILLER_76_239 ();
 sg13g2_decap_8 FILLER_76_246 ();
 sg13g2_decap_8 FILLER_76_253 ();
 sg13g2_decap_8 FILLER_76_260 ();
 sg13g2_decap_8 FILLER_76_267 ();
 sg13g2_fill_2 FILLER_76_274 ();
 sg13g2_fill_1 FILLER_76_276 ();
 sg13g2_fill_2 FILLER_76_283 ();
 sg13g2_fill_2 FILLER_76_300 ();
 sg13g2_fill_2 FILLER_76_307 ();
 sg13g2_fill_2 FILLER_76_319 ();
 sg13g2_fill_2 FILLER_76_353 ();
 sg13g2_fill_2 FILLER_76_387 ();
 sg13g2_fill_2 FILLER_76_398 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_fill_2 FILLER_77_49 ();
 sg13g2_fill_1 FILLER_77_112 ();
 sg13g2_fill_1 FILLER_77_189 ();
 sg13g2_fill_2 FILLER_77_216 ();
 sg13g2_fill_1 FILLER_77_218 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_fill_2 FILLER_77_294 ();
 sg13g2_fill_2 FILLER_77_331 ();
 sg13g2_fill_1 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_fill_2 FILLER_78_49 ();
 sg13g2_fill_2 FILLER_78_78 ();
 sg13g2_fill_1 FILLER_78_80 ();
 sg13g2_fill_1 FILLER_78_115 ();
 sg13g2_fill_1 FILLER_78_316 ();
 sg13g2_fill_2 FILLER_78_400 ();
 sg13g2_fill_1 FILLER_78_402 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_fill_2 FILLER_79_56 ();
 sg13g2_fill_1 FILLER_79_58 ();
 sg13g2_fill_2 FILLER_79_95 ();
 sg13g2_fill_1 FILLER_79_97 ();
 sg13g2_fill_1 FILLER_79_137 ();
 sg13g2_decap_8 FILLER_79_164 ();
 sg13g2_decap_8 FILLER_79_171 ();
 sg13g2_decap_8 FILLER_79_178 ();
 sg13g2_fill_2 FILLER_79_185 ();
 sg13g2_fill_1 FILLER_79_187 ();
 sg13g2_fill_2 FILLER_79_244 ();
 sg13g2_fill_1 FILLER_79_266 ();
 sg13g2_fill_2 FILLER_79_357 ();
 sg13g2_fill_2 FILLER_79_395 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_fill_2 FILLER_80_60 ();
 sg13g2_fill_2 FILLER_80_83 ();
 sg13g2_fill_2 FILLER_80_107 ();
 sg13g2_fill_2 FILLER_80_150 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_4 FILLER_80_180 ();
 sg13g2_decap_4 FILLER_80_188 ();
 sg13g2_fill_1 FILLER_80_196 ();
 sg13g2_fill_2 FILLER_80_205 ();
 sg13g2_fill_1 FILLER_80_207 ();
 sg13g2_decap_4 FILLER_80_212 ();
 sg13g2_decap_8 FILLER_80_220 ();
 sg13g2_decap_8 FILLER_80_227 ();
 sg13g2_decap_8 FILLER_80_234 ();
 sg13g2_decap_8 FILLER_80_241 ();
 sg13g2_decap_4 FILLER_80_248 ();
 sg13g2_fill_2 FILLER_80_252 ();
 sg13g2_fill_1 FILLER_80_262 ();
 sg13g2_decap_8 FILLER_80_267 ();
 sg13g2_fill_1 FILLER_80_274 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_fill_1 FILLER_80_292 ();
 sg13g2_fill_2 FILLER_80_302 ();
 sg13g2_decap_8 FILLER_80_309 ();
 sg13g2_decap_8 FILLER_80_316 ();
 sg13g2_decap_8 FILLER_80_323 ();
 sg13g2_fill_2 FILLER_80_330 ();
 sg13g2_decap_8 FILLER_80_336 ();
 sg13g2_fill_2 FILLER_80_343 ();
 sg13g2_fill_2 FILLER_80_362 ();
 sg13g2_decap_4 FILLER_80_405 ();
 assign uio_oe[0] = net33;
 assign uio_oe[1] = net34;
 assign uio_oe[2] = net35;
 assign uio_oe[3] = net36;
 assign uio_oe[4] = net2;
 assign uio_oe[5] = net37;
 assign uio_oe[6] = net3;
 assign uio_oe[7] = net4;
 assign uio_out[0] = net5;
 assign uio_out[1] = net6;
 assign uio_out[2] = net7;
 assign uio_out[3] = net8;
 assign uio_out[4] = net9;
 assign uio_out[5] = net10;
 assign uio_out[6] = net11;
 assign uio_out[7] = net12;
 assign uo_out[3] = net13;
 assign uo_out[4] = net14;
 assign uo_out[5] = net15;
 assign uo_out[6] = net16;
 assign uo_out[7] = net17;
endmodule
