module tt_um_bleeptrack_prism (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \dist_x[0] ;
 wire \dist_y[0] ;
 wire hsync;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;

 sg13g2_inv_1 _455_ (.Y(_056_),
    .A(net67));
 sg13g2_inv_1 _456_ (.Y(_057_),
    .A(\hvsync_gen.vpos[3] ));
 sg13g2_inv_1 _457_ (.Y(_058_),
    .A(net37));
 sg13g2_inv_1 _458_ (.Y(_059_),
    .A(net38));
 sg13g2_inv_1 _459_ (.Y(_060_),
    .A(\hvsync_gen.hpos[7] ));
 sg13g2_inv_1 _460_ (.Y(_061_),
    .A(\hvsync_gen.hpos[6] ));
 sg13g2_inv_1 _461_ (.Y(_062_),
    .A(net101));
 sg13g2_inv_1 _462_ (.Y(_063_),
    .A(_004_));
 sg13g2_inv_1 _463_ (.Y(_064_),
    .A(_003_));
 sg13g2_inv_1 _464_ (.Y(_065_),
    .A(_012_));
 sg13g2_inv_1 _465_ (.Y(_066_),
    .A(_015_));
 sg13g2_inv_1 _466_ (.Y(_067_),
    .A(\counter[4] ));
 sg13g2_inv_1 _467_ (.Y(_068_),
    .A(_019_));
 sg13g2_inv_2 _468_ (.Y(_069_),
    .A(\counter[6] ));
 sg13g2_inv_1 _469_ (.Y(_070_),
    .A(_022_));
 sg13g2_inv_1 _470_ (.Y(_071_),
    .A(\counter[9] ));
 sg13g2_and4_1 _471_ (.A(\hvsync_gen.vpos[7] ),
    .B(\hvsync_gen.vpos[6] ),
    .C(net37),
    .D(net92),
    .X(_072_));
 sg13g2_nor3_1 _472_ (.A(\hvsync_gen.vpos[2] ),
    .B(net38),
    .C(\hvsync_gen.vpos[9] ),
    .Y(_073_));
 sg13g2_and4_1 _473_ (.A(net89),
    .B(net93),
    .C(_072_),
    .D(_073_),
    .X(_001_));
 sg13g2_nand2_1 _474_ (.Y(_074_),
    .A(net40),
    .B(\hvsync_gen.hpos[8] ));
 sg13g2_nor2_1 _475_ (.A(\hvsync_gen.hpos[5] ),
    .B(\hvsync_gen.hpos[4] ),
    .Y(_075_));
 sg13g2_nand2_1 _476_ (.Y(_076_),
    .A(\hvsync_gen.hpos[7] ),
    .B(net40));
 sg13g2_a21o_1 _477_ (.A2(_075_),
    .A1(_061_),
    .B1(_076_),
    .X(_077_));
 sg13g2_nor2_1 _478_ (.A(_060_),
    .B(_061_),
    .Y(_078_));
 sg13g2_nand3_1 _479_ (.B(\hvsync_gen.hpos[4] ),
    .C(_078_),
    .A(\hvsync_gen.hpos[5] ),
    .Y(_079_));
 sg13g2_nor2b_1 _480_ (.A(\hvsync_gen.hpos[8] ),
    .B_N(net40),
    .Y(_080_));
 sg13g2_a21oi_1 _481_ (.A1(_079_),
    .A2(_080_),
    .Y(_081_),
    .B1(net70));
 sg13g2_a21oi_1 _482_ (.A1(_074_),
    .A2(_077_),
    .Y(_000_),
    .B1(net71));
 sg13g2_a21oi_2 _483_ (.B1(_002_),
    .Y(_082_),
    .A2(_062_),
    .A1(_060_));
 sg13g2_nor3_2 _484_ (.A(\hvsync_gen.vpos[9] ),
    .B(_072_),
    .C(_082_),
    .Y(_083_));
 sg13g2_and2_1 _485_ (.A(net37),
    .B(net38),
    .X(_084_));
 sg13g2_nand2_1 _486_ (.Y(_085_),
    .A(net37),
    .B(net38));
 sg13g2_nand4_1 _487_ (.B(\hvsync_gen.vpos[6] ),
    .C(net37),
    .A(\hvsync_gen.vpos[7] ),
    .Y(_086_),
    .D(net38));
 sg13g2_nor2_2 _488_ (.A(\hvsync_gen.vpos[8] ),
    .B(\hvsync_gen.vpos[9] ),
    .Y(_087_));
 sg13g2_or2_1 _489_ (.X(_088_),
    .B(\hvsync_gen.vpos[9] ),
    .A(\hvsync_gen.vpos[8] ));
 sg13g2_and2_1 _490_ (.A(_086_),
    .B(_087_),
    .X(_089_));
 sg13g2_or2_1 _491_ (.X(_090_),
    .B(\hvsync_gen.vpos[1] ),
    .A(net39));
 sg13g2_nor3_1 _492_ (.A(net39),
    .B(\hvsync_gen.vpos[1] ),
    .C(\hvsync_gen.vpos[2] ),
    .Y(_091_));
 sg13g2_nor4_2 _493_ (.A(net39),
    .B(\hvsync_gen.vpos[1] ),
    .C(\hvsync_gen.vpos[3] ),
    .Y(_092_),
    .D(\hvsync_gen.vpos[2] ));
 sg13g2_o21ai_1 _494_ (.B1(_010_),
    .Y(_093_),
    .A1(_086_),
    .A2(_092_));
 sg13g2_nor3_1 _495_ (.A(_010_),
    .B(_086_),
    .C(_092_),
    .Y(_094_));
 sg13g2_o21ai_1 _496_ (.B1(_087_),
    .Y(_095_),
    .A1(_086_),
    .A2(_092_));
 sg13g2_nor2b_1 _497_ (.A(_094_),
    .B_N(_095_),
    .Y(_096_));
 sg13g2_a21o_2 _498_ (.A2(_096_),
    .A1(_093_),
    .B1(_089_),
    .X(_097_));
 sg13g2_nor2_1 _499_ (.A(\hvsync_gen.hpos[7] ),
    .B(\hvsync_gen.hpos[6] ),
    .Y(_098_));
 sg13g2_nand2_1 _500_ (.Y(_099_),
    .A(_060_),
    .B(_061_));
 sg13g2_or2_1 _501_ (.X(_100_),
    .B(\hvsync_gen.hpos[1] ),
    .A(net41));
 sg13g2_nor4_2 _502_ (.A(net41),
    .B(\hvsync_gen.hpos[3] ),
    .C(\hvsync_gen.hpos[2] ),
    .Y(_101_),
    .D(\hvsync_gen.hpos[1] ));
 sg13g2_nor3_1 _503_ (.A(\hvsync_gen.hpos[5] ),
    .B(\hvsync_gen.hpos[4] ),
    .C(\hvsync_gen.hpos[7] ),
    .Y(_102_));
 sg13g2_a21oi_1 _504_ (.A1(_101_),
    .A2(_102_),
    .Y(_103_),
    .B1(_098_));
 sg13g2_inv_1 _505_ (.Y(_104_),
    .A(_103_));
 sg13g2_a221oi_1 _506_ (.B2(_102_),
    .C1(_062_),
    .B1(_101_),
    .A1(_060_),
    .Y(_105_),
    .A2(_061_));
 sg13g2_nor2_2 _507_ (.A(net40),
    .B(_105_),
    .Y(_106_));
 sg13g2_a22oi_1 _508_ (.Y(_107_),
    .B1(_106_),
    .B2(_099_),
    .A2(_104_),
    .A1(net40));
 sg13g2_xnor2_1 _509_ (.Y(_108_),
    .A(\hvsync_gen.hpos[8] ),
    .B(_107_));
 sg13g2_nand2_1 _510_ (.Y(_109_),
    .A(_097_),
    .B(_108_));
 sg13g2_a21oi_2 _511_ (.B1(_092_),
    .Y(_110_),
    .A2(_087_),
    .A1(_086_));
 sg13g2_a22oi_1 _512_ (.Y(_111_),
    .B1(_110_),
    .B2(_066_),
    .A2(_087_),
    .A1(_059_));
 sg13g2_xnor2_1 _513_ (.Y(_112_),
    .A(\hvsync_gen.vpos[5] ),
    .B(_111_));
 sg13g2_inv_1 _514_ (.Y(_113_),
    .A(_112_));
 sg13g2_nand2b_1 _515_ (.Y(_114_),
    .B(_101_),
    .A_N(\hvsync_gen.hpos[4] ));
 sg13g2_nand2_1 _516_ (.Y(_115_),
    .A(_075_),
    .B(_101_));
 sg13g2_xnor2_1 _517_ (.Y(_116_),
    .A(\hvsync_gen.hpos[5] ),
    .B(_114_));
 sg13g2_mux2_2 _518_ (.A0(_116_),
    .A1(_014_),
    .S(_106_),
    .X(_117_));
 sg13g2_and2_1 _519_ (.A(_112_),
    .B(_117_),
    .X(_118_));
 sg13g2_xnor2_1 _520_ (.Y(_119_),
    .A(\hvsync_gen.vpos[4] ),
    .B(_110_));
 sg13g2_xor2_1 _521_ (.B(_101_),
    .A(\hvsync_gen.hpos[4] ),
    .X(_120_));
 sg13g2_mux2_2 _522_ (.A0(_120_),
    .A1(_016_),
    .S(_106_),
    .X(_121_));
 sg13g2_inv_1 _523_ (.Y(_122_),
    .A(_121_));
 sg13g2_nand2_1 _524_ (.Y(_123_),
    .A(_119_),
    .B(_122_));
 sg13g2_xnor2_1 _525_ (.Y(_124_),
    .A(_119_),
    .B(_121_));
 sg13g2_and2_1 _526_ (.A(net41),
    .B(\hvsync_gen.hpos[1] ),
    .X(_125_));
 sg13g2_xnor2_1 _527_ (.Y(_126_),
    .A(net84),
    .B(\hvsync_gen.hpos[1] ));
 sg13g2_inv_1 _528_ (.Y(_127_),
    .A(_126_));
 sg13g2_or3_1 _529_ (.A(\hvsync_gen.hpos[9] ),
    .B(_007_),
    .C(_105_),
    .X(_128_));
 sg13g2_o21ai_1 _530_ (.B1(_127_),
    .Y(_129_),
    .A1(\hvsync_gen.hpos[9] ),
    .A2(_105_));
 sg13g2_and2_1 _531_ (.A(_128_),
    .B(_129_),
    .X(_130_));
 sg13g2_nand2_1 _532_ (.Y(_131_),
    .A(net39),
    .B(\hvsync_gen.vpos[1] ));
 sg13g2_nand2_1 _533_ (.Y(_132_),
    .A(_090_),
    .B(_131_));
 sg13g2_mux2_1 _534_ (.A0(_008_),
    .A1(_132_),
    .S(_095_),
    .X(_133_));
 sg13g2_inv_1 _535_ (.Y(_134_),
    .A(_133_));
 sg13g2_a21oi_1 _536_ (.A1(_128_),
    .A2(_129_),
    .Y(_135_),
    .B1(_133_));
 sg13g2_nand3_1 _537_ (.B(_129_),
    .C(_133_),
    .A(_128_),
    .Y(_136_));
 sg13g2_nand2b_1 _538_ (.Y(_137_),
    .B(_136_),
    .A_N(_135_));
 sg13g2_and2_1 _539_ (.A(\dist_y[0] ),
    .B(net41),
    .X(_138_));
 sg13g2_a21oi_1 _540_ (.A1(_136_),
    .A2(_138_),
    .Y(_139_),
    .B1(_135_));
 sg13g2_o21ai_1 _541_ (.B1(_100_),
    .Y(_140_),
    .A1(\hvsync_gen.hpos[9] ),
    .A2(_105_));
 sg13g2_xnor2_1 _542_ (.Y(_141_),
    .A(_004_),
    .B(_140_));
 sg13g2_xnor2_1 _543_ (.Y(_142_),
    .A(\hvsync_gen.vpos[2] ),
    .B(_090_));
 sg13g2_mux2_2 _544_ (.A0(_005_),
    .A1(_142_),
    .S(_095_),
    .X(_143_));
 sg13g2_inv_1 _545_ (.Y(_144_),
    .A(_143_));
 sg13g2_nand2b_1 _546_ (.Y(_145_),
    .B(\hvsync_gen.vpos[3] ),
    .A_N(_091_));
 sg13g2_nor2_1 _547_ (.A(_018_),
    .B(_095_),
    .Y(_146_));
 sg13g2_a21oi_2 _548_ (.B1(_146_),
    .Y(_147_),
    .A2(_145_),
    .A1(_110_));
 sg13g2_inv_1 _549_ (.Y(_148_),
    .A(_147_));
 sg13g2_nor2_1 _550_ (.A(_063_),
    .B(_100_),
    .Y(_149_));
 sg13g2_xor2_1 _551_ (.B(_149_),
    .A(\hvsync_gen.hpos[3] ),
    .X(_150_));
 sg13g2_mux2_2 _552_ (.A0(_150_),
    .A1(_017_),
    .S(_106_),
    .X(_151_));
 sg13g2_or2_1 _553_ (.X(_152_),
    .B(_151_),
    .A(_147_));
 sg13g2_xnor2_1 _554_ (.Y(_153_),
    .A(_147_),
    .B(_151_));
 sg13g2_nand2b_1 _555_ (.Y(_154_),
    .B(_144_),
    .A_N(_141_));
 sg13g2_xnor2_1 _556_ (.Y(_155_),
    .A(_141_),
    .B(_143_));
 sg13g2_nor3_2 _557_ (.A(_139_),
    .B(_153_),
    .C(_155_),
    .Y(_156_));
 sg13g2_o21ai_1 _558_ (.B1(_152_),
    .Y(_157_),
    .A1(_153_),
    .A2(_154_));
 sg13g2_o21ai_1 _559_ (.B1(_124_),
    .Y(_158_),
    .A1(_156_),
    .A2(_157_));
 sg13g2_nor2_1 _560_ (.A(_112_),
    .B(_117_),
    .Y(_159_));
 sg13g2_a21oi_1 _561_ (.A1(_119_),
    .A2(_122_),
    .Y(_160_),
    .B1(_159_));
 sg13g2_a21oi_1 _562_ (.A1(_158_),
    .A2(_160_),
    .Y(_161_),
    .B1(_118_));
 sg13g2_a21o_1 _563_ (.A2(_160_),
    .A1(_158_),
    .B1(_118_),
    .X(_162_));
 sg13g2_a221oi_1 _564_ (.B2(_057_),
    .C1(_085_),
    .B1(_091_),
    .A1(_086_),
    .Y(_163_),
    .A2(_087_));
 sg13g2_a21o_1 _565_ (.A2(_087_),
    .A1(_085_),
    .B1(_163_),
    .X(_164_));
 sg13g2_xor2_1 _566_ (.B(_164_),
    .A(\hvsync_gen.vpos[6] ),
    .X(_165_));
 sg13g2_xnor2_1 _567_ (.Y(_166_),
    .A(_013_),
    .B(_115_));
 sg13g2_mux2_2 _568_ (.A0(_166_),
    .A1(\hvsync_gen.hpos[6] ),
    .S(_106_),
    .X(_167_));
 sg13g2_nand2_1 _569_ (.Y(_168_),
    .A(_165_),
    .B(_167_));
 sg13g2_or4_1 _570_ (.A(net40),
    .B(_078_),
    .C(_098_),
    .D(_105_),
    .X(_169_));
 sg13g2_a21oi_1 _571_ (.A1(_075_),
    .A2(_101_),
    .Y(_170_),
    .B1(_061_));
 sg13g2_xnor2_1 _572_ (.Y(_171_),
    .A(_011_),
    .B(_170_));
 sg13g2_o21ai_1 _573_ (.B1(_169_),
    .Y(_172_),
    .A1(_106_),
    .A2(_171_));
 sg13g2_inv_1 _574_ (.Y(_173_),
    .A(_172_));
 sg13g2_a21oi_1 _575_ (.A1(\hvsync_gen.vpos[6] ),
    .A2(_084_),
    .Y(_174_),
    .B1(_088_));
 sg13g2_a21oi_1 _576_ (.A1(_065_),
    .A2(_163_),
    .Y(_175_),
    .B1(_174_));
 sg13g2_xnor2_1 _577_ (.Y(_176_),
    .A(\hvsync_gen.vpos[7] ),
    .B(_175_));
 sg13g2_nand2_1 _578_ (.Y(_177_),
    .A(_172_),
    .B(_176_));
 sg13g2_inv_1 _579_ (.Y(_178_),
    .A(_177_));
 sg13g2_nor2_1 _580_ (.A(_165_),
    .B(_167_),
    .Y(_179_));
 sg13g2_nor2_1 _581_ (.A(_172_),
    .B(_176_),
    .Y(_180_));
 sg13g2_or2_1 _582_ (.X(_181_),
    .B(_180_),
    .A(_179_));
 sg13g2_nor2_1 _583_ (.A(_178_),
    .B(_180_),
    .Y(_182_));
 sg13g2_nor2_1 _584_ (.A(_178_),
    .B(_181_),
    .Y(_183_));
 sg13g2_nand3b_1 _585_ (.B(_177_),
    .C(_168_),
    .Y(_184_),
    .A_N(_181_));
 sg13g2_a221oi_1 _586_ (.B2(_160_),
    .C1(_184_),
    .B1(_158_),
    .A1(_112_),
    .Y(_185_),
    .A2(_117_));
 sg13g2_and2_1 _587_ (.A(_177_),
    .B(_181_),
    .X(_186_));
 sg13g2_or2_1 _588_ (.X(_187_),
    .B(_186_),
    .A(_185_));
 sg13g2_nand3_1 _589_ (.B(_099_),
    .C(_106_),
    .A(\hvsync_gen.hpos[8] ),
    .Y(_188_));
 sg13g2_nor2_1 _590_ (.A(_009_),
    .B(_104_),
    .Y(_189_));
 sg13g2_xnor2_1 _591_ (.Y(_190_),
    .A(_002_),
    .B(_189_));
 sg13g2_o21ai_1 _592_ (.B1(_188_),
    .Y(_191_),
    .A1(_106_),
    .A2(_190_));
 sg13g2_xor2_1 _593_ (.B(_093_),
    .A(\hvsync_gen.vpos[9] ),
    .X(_192_));
 sg13g2_a22oi_1 _594_ (.Y(_193_),
    .B1(_095_),
    .B2(_192_),
    .A2(_089_),
    .A1(_010_));
 sg13g2_xor2_1 _595_ (.B(_193_),
    .A(_191_),
    .X(_194_));
 sg13g2_o21ai_1 _596_ (.B1(_194_),
    .Y(_195_),
    .A1(_185_),
    .A2(_186_));
 sg13g2_and2_1 _597_ (.A(_109_),
    .B(_195_),
    .X(_196_));
 sg13g2_o21ai_1 _598_ (.B1(_194_),
    .Y(_197_),
    .A1(_097_),
    .A2(_108_));
 sg13g2_a22oi_1 _599_ (.Y(_198_),
    .B1(_197_),
    .B2(_187_),
    .A2(_195_),
    .A1(_109_));
 sg13g2_a22oi_1 _600_ (.Y(_199_),
    .B1(_182_),
    .B2(_162_),
    .A2(_167_),
    .A1(_165_));
 sg13g2_nor2_1 _601_ (.A(_161_),
    .B(_183_),
    .Y(_200_));
 sg13g2_or3_1 _602_ (.A(_124_),
    .B(_156_),
    .C(_157_),
    .X(_201_));
 sg13g2_and2_1 _603_ (.A(_158_),
    .B(_201_),
    .X(_202_));
 sg13g2_nand3_1 _604_ (.B(_143_),
    .C(_153_),
    .A(_141_),
    .Y(_203_));
 sg13g2_o21ai_1 _605_ (.B1(_203_),
    .Y(_204_),
    .A1(_153_),
    .A2(_154_));
 sg13g2_a21oi_1 _606_ (.A1(_139_),
    .A2(_204_),
    .Y(_205_),
    .B1(_156_));
 sg13g2_nor2_1 _607_ (.A(\dist_y[0] ),
    .B(net41),
    .Y(_206_));
 sg13g2_mux2_1 _608_ (.A0(_138_),
    .A1(_206_),
    .S(_137_),
    .X(_207_));
 sg13g2_nand2b_1 _609_ (.Y(_208_),
    .B(_207_),
    .A_N(_205_));
 sg13g2_or2_1 _610_ (.X(_209_),
    .B(_159_),
    .A(_118_));
 sg13g2_nand2_1 _611_ (.Y(_210_),
    .A(_123_),
    .B(_158_));
 sg13g2_xnor2_1 _612_ (.Y(_211_),
    .A(_209_),
    .B(_210_));
 sg13g2_o21ai_1 _613_ (.B1(_211_),
    .Y(_212_),
    .A1(_202_),
    .A2(_208_));
 sg13g2_mux2_1 _614_ (.A0(_200_),
    .A1(_183_),
    .S(_199_),
    .X(_213_));
 sg13g2_a221oi_1 _615_ (.B2(_213_),
    .C1(_198_),
    .B1(_212_),
    .A1(_196_),
    .Y(_214_),
    .A2(_197_));
 sg13g2_nor2_1 _616_ (.A(_057_),
    .B(net4),
    .Y(_215_));
 sg13g2_xnor2_1 _617_ (.Y(_216_),
    .A(_017_),
    .B(_215_));
 sg13g2_nand2b_1 _618_ (.Y(_217_),
    .B(net39),
    .A_N(net1));
 sg13g2_o21ai_1 _619_ (.B1(\counter[0] ),
    .Y(_218_),
    .A1(_025_),
    .A2(_217_));
 sg13g2_a21o_1 _620_ (.A2(_217_),
    .A1(_025_),
    .B1(_218_),
    .X(_219_));
 sg13g2_nor2b_1 _621_ (.A(net2),
    .B_N(\hvsync_gen.vpos[1] ),
    .Y(_220_));
 sg13g2_xnor2_1 _622_ (.Y(_221_),
    .A(_007_),
    .B(_220_));
 sg13g2_xor2_1 _623_ (.B(_221_),
    .A(_006_),
    .X(_222_));
 sg13g2_nand2_1 _624_ (.Y(_223_),
    .A(\counter[1] ),
    .B(_221_));
 sg13g2_o21ai_1 _625_ (.B1(_223_),
    .Y(_224_),
    .A1(_219_),
    .A2(_222_));
 sg13g2_nor2b_1 _626_ (.A(net3),
    .B_N(\hvsync_gen.vpos[2] ),
    .Y(_225_));
 sg13g2_xnor2_1 _627_ (.Y(_226_),
    .A(_004_),
    .B(_225_));
 sg13g2_xor2_1 _628_ (.B(_226_),
    .A(\counter[2] ),
    .X(_227_));
 sg13g2_a22oi_1 _629_ (.Y(_228_),
    .B1(_227_),
    .B2(_224_),
    .A2(_226_),
    .A1(_064_));
 sg13g2_xnor2_1 _630_ (.Y(_229_),
    .A(\counter[3] ),
    .B(_216_));
 sg13g2_nor2_1 _631_ (.A(_228_),
    .B(_229_),
    .Y(_230_));
 sg13g2_a21oi_2 _632_ (.B1(_230_),
    .Y(_231_),
    .A2(_216_),
    .A1(_068_));
 sg13g2_nand2_1 _633_ (.Y(_232_),
    .A(net38),
    .B(net5));
 sg13g2_xor2_1 _634_ (.B(_016_),
    .A(net41),
    .X(_233_));
 sg13g2_xnor2_1 _635_ (.Y(_234_),
    .A(_232_),
    .B(_233_));
 sg13g2_or2_1 _636_ (.X(_235_),
    .B(_234_),
    .A(_020_));
 sg13g2_xnor2_1 _637_ (.Y(_236_),
    .A(\hvsync_gen.hpos[2] ),
    .B(_013_));
 sg13g2_nand2_1 _638_ (.Y(_237_),
    .A(\hvsync_gen.vpos[6] ),
    .B(net7));
 sg13g2_xnor2_1 _639_ (.Y(_238_),
    .A(_236_),
    .B(_237_));
 sg13g2_xnor2_1 _640_ (.Y(_239_),
    .A(_069_),
    .B(_238_));
 sg13g2_nand2_1 _641_ (.Y(_240_),
    .A(net37),
    .B(net6));
 sg13g2_xnor2_1 _642_ (.Y(_241_),
    .A(\hvsync_gen.hpos[1] ),
    .B(_014_));
 sg13g2_xnor2_1 _643_ (.Y(_242_),
    .A(_240_),
    .B(_241_));
 sg13g2_xor2_1 _644_ (.B(_242_),
    .A(\counter[5] ),
    .X(_243_));
 sg13g2_a22oi_1 _645_ (.Y(_244_),
    .B1(_239_),
    .B2(_243_),
    .A2(_235_),
    .A1(_231_));
 sg13g2_xnor2_1 _646_ (.Y(_245_),
    .A(\counter[4] ),
    .B(_234_));
 sg13g2_nand2b_1 _647_ (.Y(_246_),
    .B(_242_),
    .A_N(_021_));
 sg13g2_a21o_1 _648_ (.A2(_246_),
    .A1(_239_),
    .B1(_243_),
    .X(_247_));
 sg13g2_a21oi_1 _649_ (.A1(_235_),
    .A2(_247_),
    .Y(_248_),
    .B1(_245_));
 sg13g2_nand2b_1 _650_ (.Y(_249_),
    .B(_231_),
    .A_N(_248_));
 sg13g2_nor2_1 _651_ (.A(_231_),
    .B(_245_),
    .Y(_250_));
 sg13g2_xor2_1 _652_ (.B(_229_),
    .A(_228_),
    .X(_251_));
 sg13g2_a21oi_1 _653_ (.A1(\counter[6] ),
    .A2(_070_),
    .Y(_252_),
    .B1(_239_));
 sg13g2_nand2_1 _654_ (.Y(_253_),
    .A(\hvsync_gen.vpos[7] ),
    .B(net8));
 sg13g2_xnor2_1 _655_ (.Y(_254_),
    .A(\counter[7] ),
    .B(_253_));
 sg13g2_xnor2_1 _656_ (.Y(_255_),
    .A(\hvsync_gen.hpos[3] ),
    .B(_011_));
 sg13g2_xnor2_1 _657_ (.Y(_256_),
    .A(_254_),
    .B(_255_));
 sg13g2_xnor2_1 _658_ (.Y(_257_),
    .A(_252_),
    .B(_256_));
 sg13g2_o21ai_1 _659_ (.B1(_257_),
    .Y(_258_),
    .A1(_239_),
    .A2(_246_));
 sg13g2_nor3_1 _660_ (.A(_250_),
    .B(_251_),
    .C(_258_),
    .Y(_259_));
 sg13g2_nand3b_1 _661_ (.B(_249_),
    .C(_259_),
    .Y(_260_),
    .A_N(_244_));
 sg13g2_xnor2_1 _662_ (.Y(_261_),
    .A(_219_),
    .B(_222_));
 sg13g2_nor2_1 _663_ (.A(_260_),
    .B(_261_),
    .Y(_262_));
 sg13g2_o21ai_1 _664_ (.B1(_083_),
    .Y(_263_),
    .A1(_214_),
    .A2(_262_));
 sg13g2_xnor2_1 _665_ (.Y(_264_),
    .A(\counter[1] ),
    .B(_130_));
 sg13g2_o21ai_1 _666_ (.B1(\counter[0] ),
    .Y(_265_),
    .A1(net39),
    .A2(net41));
 sg13g2_nand2b_1 _667_ (.Y(_266_),
    .B(_265_),
    .A_N(_138_));
 sg13g2_o21ai_1 _668_ (.B1(_266_),
    .Y(_267_),
    .A1(_134_),
    .A2(_264_));
 sg13g2_a21oi_1 _669_ (.A1(_134_),
    .A2(_264_),
    .Y(_268_),
    .B1(_267_));
 sg13g2_nor2_1 _670_ (.A(_006_),
    .B(_130_),
    .Y(_269_));
 sg13g2_a21oi_1 _671_ (.A1(_134_),
    .A2(_264_),
    .Y(_270_),
    .B1(_269_));
 sg13g2_nor2_1 _672_ (.A(_003_),
    .B(_141_),
    .Y(_271_));
 sg13g2_xnor2_1 _673_ (.Y(_272_),
    .A(_064_),
    .B(_141_));
 sg13g2_xnor2_1 _674_ (.Y(_273_),
    .A(_143_),
    .B(_272_));
 sg13g2_nor2b_1 _675_ (.A(_270_),
    .B_N(_273_),
    .Y(_274_));
 sg13g2_xnor2_1 _676_ (.Y(_275_),
    .A(_270_),
    .B(_273_));
 sg13g2_nand2_1 _677_ (.Y(_276_),
    .A(_268_),
    .B(_275_));
 sg13g2_o21ai_1 _678_ (.B1(net1),
    .Y(_277_),
    .A1(_268_),
    .A2(_275_));
 sg13g2_nand2b_1 _679_ (.Y(_278_),
    .B(_276_),
    .A_N(_277_));
 sg13g2_a21oi_2 _680_ (.B1(_263_),
    .Y(uo_out[4]),
    .A2(_278_),
    .A1(_214_));
 sg13g2_xnor2_1 _681_ (.Y(_279_),
    .A(_224_),
    .B(_227_));
 sg13g2_nor2_1 _682_ (.A(_260_),
    .B(_279_),
    .Y(_280_));
 sg13g2_o21ai_1 _683_ (.B1(_083_),
    .Y(_281_),
    .A1(_214_),
    .A2(_280_));
 sg13g2_xnor2_1 _684_ (.Y(_282_),
    .A(_023_),
    .B(net41));
 sg13g2_o21ai_1 _685_ (.B1(net2),
    .Y(_283_),
    .A1(\counter[0] ),
    .A2(_282_));
 sg13g2_a21o_1 _686_ (.A2(_282_),
    .A1(\counter[0] ),
    .B1(_283_),
    .X(_284_));
 sg13g2_a21oi_2 _687_ (.B1(_281_),
    .Y(uo_out[0]),
    .A2(_284_),
    .A1(_214_));
 sg13g2_xnor2_1 _688_ (.Y(_285_),
    .A(_069_),
    .B(_167_));
 sg13g2_nor2_1 _689_ (.A(_165_),
    .B(_285_),
    .Y(_286_));
 sg13g2_nor2_1 _690_ (.A(_022_),
    .B(_167_),
    .Y(_287_));
 sg13g2_nand2_1 _691_ (.Y(_288_),
    .A(\counter[7] ),
    .B(_173_));
 sg13g2_xor2_1 _692_ (.B(_172_),
    .A(\counter[7] ),
    .X(_289_));
 sg13g2_xor2_1 _693_ (.B(_289_),
    .A(_176_),
    .X(_290_));
 sg13g2_or3_1 _694_ (.A(_286_),
    .B(_287_),
    .C(_290_),
    .X(_291_));
 sg13g2_o21ai_1 _695_ (.B1(_290_),
    .Y(_292_),
    .A1(_286_),
    .A2(_287_));
 sg13g2_nand2_1 _696_ (.Y(_293_),
    .A(_291_),
    .B(_292_));
 sg13g2_xnor2_1 _697_ (.Y(_294_),
    .A(_165_),
    .B(_285_));
 sg13g2_xnor2_1 _698_ (.Y(_295_),
    .A(\counter[5] ),
    .B(_117_));
 sg13g2_nor2_1 _699_ (.A(_021_),
    .B(_117_),
    .Y(_296_));
 sg13g2_a21oi_1 _700_ (.A1(_113_),
    .A2(_295_),
    .Y(_297_),
    .B1(_296_));
 sg13g2_or2_1 _701_ (.X(_298_),
    .B(_297_),
    .A(_294_));
 sg13g2_xnor2_1 _702_ (.Y(_299_),
    .A(_294_),
    .B(_297_));
 sg13g2_inv_1 _703_ (.Y(_300_),
    .A(_299_));
 sg13g2_xnor2_1 _704_ (.Y(_301_),
    .A(\counter[3] ),
    .B(_151_));
 sg13g2_xnor2_1 _705_ (.Y(_302_),
    .A(_148_),
    .B(_301_));
 sg13g2_a21oi_1 _706_ (.A1(_144_),
    .A2(_272_),
    .Y(_303_),
    .B1(_271_));
 sg13g2_nor2_1 _707_ (.A(_302_),
    .B(_303_),
    .Y(_304_));
 sg13g2_nor2_1 _708_ (.A(_274_),
    .B(_304_),
    .Y(_305_));
 sg13g2_a22oi_1 _709_ (.Y(_306_),
    .B1(_305_),
    .B2(_276_),
    .A2(_303_),
    .A1(_302_));
 sg13g2_xnor2_1 _710_ (.Y(_307_),
    .A(\counter[4] ),
    .B(_121_));
 sg13g2_nand2_1 _711_ (.Y(_308_),
    .A(_119_),
    .B(_307_));
 sg13g2_xor2_1 _712_ (.B(_307_),
    .A(_119_),
    .X(_309_));
 sg13g2_nor2_1 _713_ (.A(_019_),
    .B(_151_),
    .Y(_310_));
 sg13g2_a21oi_1 _714_ (.A1(_148_),
    .A2(_301_),
    .Y(_311_),
    .B1(_310_));
 sg13g2_nand2b_1 _715_ (.Y(_312_),
    .B(_309_),
    .A_N(_311_));
 sg13g2_xnor2_1 _716_ (.Y(_313_),
    .A(_309_),
    .B(_311_));
 sg13g2_or2_1 _717_ (.X(_314_),
    .B(_121_),
    .A(_020_));
 sg13g2_xnor2_1 _718_ (.Y(_315_),
    .A(_113_),
    .B(_295_));
 sg13g2_a21o_1 _719_ (.A2(_314_),
    .A1(_308_),
    .B1(_315_),
    .X(_316_));
 sg13g2_and3_1 _720_ (.X(_317_),
    .A(_308_),
    .B(_314_),
    .C(_315_));
 sg13g2_nand3b_1 _721_ (.B(_313_),
    .C(_316_),
    .Y(_318_),
    .A_N(_317_));
 sg13g2_a221oi_1 _722_ (.B2(_276_),
    .C1(_318_),
    .B1(_305_),
    .A1(_302_),
    .Y(_319_),
    .A2(_303_));
 sg13g2_a21oi_2 _723_ (.B1(_317_),
    .Y(_320_),
    .A2(_316_),
    .A1(_312_));
 sg13g2_o21ai_1 _724_ (.B1(_300_),
    .Y(_321_),
    .A1(_319_),
    .A2(_320_));
 sg13g2_a21o_1 _725_ (.A2(_321_),
    .A1(_298_),
    .B1(_293_),
    .X(_322_));
 sg13g2_nand3_1 _726_ (.B(_298_),
    .C(_321_),
    .A(_293_),
    .Y(_323_));
 sg13g2_nand3_1 _727_ (.B(_322_),
    .C(_323_),
    .A(net3),
    .Y(_324_));
 sg13g2_a21oi_2 _728_ (.B1(_263_),
    .Y(uo_out[5]),
    .A2(_324_),
    .A1(_214_));
 sg13g2_o21ai_1 _729_ (.B1(net4),
    .Y(_325_),
    .A1(_306_),
    .A2(_313_));
 sg13g2_a21o_1 _730_ (.A2(_313_),
    .A1(_306_),
    .B1(_325_),
    .X(_326_));
 sg13g2_a21oi_2 _731_ (.B1(_281_),
    .Y(uo_out[1]),
    .A2(_326_),
    .A1(_214_));
 sg13g2_o21ai_1 _732_ (.B1(_288_),
    .Y(_327_),
    .A1(_176_),
    .A2(_289_));
 sg13g2_xnor2_1 _733_ (.Y(_328_),
    .A(\counter[8] ),
    .B(_108_));
 sg13g2_nor2b_1 _734_ (.A(_328_),
    .B_N(_097_),
    .Y(_329_));
 sg13g2_xnor2_1 _735_ (.Y(_330_),
    .A(_097_),
    .B(_328_));
 sg13g2_nor2_1 _736_ (.A(_327_),
    .B(_330_),
    .Y(_331_));
 sg13g2_nor3_1 _737_ (.A(_293_),
    .B(_299_),
    .C(_331_),
    .Y(_332_));
 sg13g2_o21ai_1 _738_ (.B1(_332_),
    .Y(_333_),
    .A1(_319_),
    .A2(_320_));
 sg13g2_nand2b_1 _739_ (.Y(_334_),
    .B(_291_),
    .A_N(_298_));
 sg13g2_nand2_1 _740_ (.Y(_335_),
    .A(_327_),
    .B(_330_));
 sg13g2_nand3_1 _741_ (.B(_334_),
    .C(_335_),
    .A(_292_),
    .Y(_336_));
 sg13g2_nand2b_1 _742_ (.Y(_337_),
    .B(_336_),
    .A_N(_331_));
 sg13g2_a21oi_1 _743_ (.A1(\counter[8] ),
    .A2(_108_),
    .Y(_338_),
    .B1(_329_));
 sg13g2_xnor2_1 _744_ (.Y(_339_),
    .A(\counter[9] ),
    .B(_194_));
 sg13g2_xnor2_1 _745_ (.Y(_340_),
    .A(_338_),
    .B(_339_));
 sg13g2_a21o_1 _746_ (.A2(_337_),
    .A1(_333_),
    .B1(_340_),
    .X(_341_));
 sg13g2_nand3_1 _747_ (.B(_337_),
    .C(_340_),
    .A(_333_),
    .Y(_342_));
 sg13g2_nand3_1 _748_ (.B(_341_),
    .C(_342_),
    .A(net5),
    .Y(_343_));
 sg13g2_a21oi_2 _749_ (.B1(_263_),
    .Y(uo_out[6]),
    .A2(_343_),
    .A1(_214_));
 sg13g2_nor3_1 _750_ (.A(_300_),
    .B(_319_),
    .C(_320_),
    .Y(_344_));
 sg13g2_nand3b_1 _751_ (.B(net6),
    .C(_321_),
    .Y(_345_),
    .A_N(_344_));
 sg13g2_a21oi_2 _752_ (.B1(_281_),
    .Y(uo_out[2]),
    .A2(_345_),
    .A1(_214_));
 sg13g2_and3_1 _753_ (.X(_346_),
    .A(\hvsync_gen.hpos[3] ),
    .B(\hvsync_gen.hpos[2] ),
    .C(_125_));
 sg13g2_nand2_1 _754_ (.Y(_347_),
    .A(\hvsync_gen.hpos[4] ),
    .B(_346_));
 sg13g2_nor4_2 _755_ (.A(\hvsync_gen.hpos[5] ),
    .B(_074_),
    .C(_099_),
    .Y(_348_),
    .D(_347_));
 sg13g2_nor2b_1 _756_ (.A(_348_),
    .B_N(net43),
    .Y(_349_));
 sg13g2_nand2b_1 _757_ (.Y(_350_),
    .B(net43),
    .A_N(_348_));
 sg13g2_and2_1 _758_ (.A(net69),
    .B(net34),
    .X(_026_));
 sg13g2_nor2_1 _759_ (.A(net85),
    .B(_350_),
    .Y(_027_));
 sg13g2_o21ai_1 _760_ (.B1(net42),
    .Y(_351_),
    .A1(net78),
    .A2(_125_));
 sg13g2_a21oi_1 _761_ (.A1(net78),
    .A2(_125_),
    .Y(_028_),
    .B1(_351_));
 sg13g2_nand2_1 _762_ (.Y(_352_),
    .A(_063_),
    .B(_125_));
 sg13g2_xor2_1 _763_ (.B(_352_),
    .A(net98),
    .X(_353_));
 sg13g2_nor2_1 _764_ (.A(_350_),
    .B(net99),
    .Y(_029_));
 sg13g2_o21ai_1 _765_ (.B1(net42),
    .Y(_354_),
    .A1(net102),
    .A2(_346_));
 sg13g2_nor2b_1 _766_ (.A(_354_),
    .B_N(_347_),
    .Y(_030_));
 sg13g2_nor2b_1 _767_ (.A(net90),
    .B_N(_346_),
    .Y(_355_));
 sg13g2_o21ai_1 _768_ (.B1(net35),
    .Y(_356_),
    .A1(\hvsync_gen.hpos[5] ),
    .A2(_355_));
 sg13g2_a21oi_1 _769_ (.A1(\hvsync_gen.hpos[5] ),
    .A2(_355_),
    .Y(_031_),
    .B1(_356_));
 sg13g2_and3_1 _770_ (.X(_357_),
    .A(\hvsync_gen.hpos[5] ),
    .B(\hvsync_gen.hpos[4] ),
    .C(_346_));
 sg13g2_o21ai_1 _771_ (.B1(net35),
    .Y(_358_),
    .A1(net73),
    .A2(_357_));
 sg13g2_a21oi_1 _772_ (.A1(net73),
    .A2(_357_),
    .Y(_032_),
    .B1(_358_));
 sg13g2_nor2b_1 _773_ (.A(_013_),
    .B_N(_357_),
    .Y(_359_));
 sg13g2_o21ai_1 _774_ (.B1(net35),
    .Y(_360_),
    .A1(net76),
    .A2(_359_));
 sg13g2_a21oi_1 _775_ (.A1(net76),
    .A2(_359_),
    .Y(_033_),
    .B1(_360_));
 sg13g2_nand2_1 _776_ (.Y(_361_),
    .A(_078_),
    .B(_357_));
 sg13g2_o21ai_1 _777_ (.B1(net35),
    .Y(_362_),
    .A1(_062_),
    .A2(_361_));
 sg13g2_a21oi_1 _778_ (.A1(_062_),
    .A2(_361_),
    .Y(_034_),
    .B1(_362_));
 sg13g2_nor2_1 _779_ (.A(net79),
    .B(_361_),
    .Y(_363_));
 sg13g2_o21ai_1 _780_ (.B1(net35),
    .Y(_364_),
    .A1(net40),
    .A2(_363_));
 sg13g2_a21oi_1 _781_ (.A1(net40),
    .A2(_363_),
    .Y(_035_),
    .B1(_364_));
 sg13g2_and2_1 _782_ (.A(net43),
    .B(_024_),
    .X(_036_));
 sg13g2_nand2_1 _783_ (.Y(_365_),
    .A(\counter[1] ),
    .B(\counter[0] ));
 sg13g2_o21ai_1 _784_ (.B1(net43),
    .Y(_366_),
    .A1(\counter[1] ),
    .A2(\counter[0] ));
 sg13g2_nor2b_1 _785_ (.A(_366_),
    .B_N(_365_),
    .Y(_037_));
 sg13g2_xnor2_1 _786_ (.Y(_367_),
    .A(\counter[2] ),
    .B(_365_));
 sg13g2_and2_1 _787_ (.A(net43),
    .B(_367_),
    .X(_038_));
 sg13g2_nor2_1 _788_ (.A(_003_),
    .B(_365_),
    .Y(_368_));
 sg13g2_o21ai_1 _789_ (.B1(net43),
    .Y(_369_),
    .A1(\counter[3] ),
    .A2(_368_));
 sg13g2_a21oi_1 _790_ (.A1(\counter[3] ),
    .A2(_368_),
    .Y(_039_),
    .B1(_369_));
 sg13g2_nand4_1 _791_ (.B(\counter[1] ),
    .C(\counter[0] ),
    .A(\counter[2] ),
    .Y(_370_),
    .D(\counter[3] ));
 sg13g2_nor2_1 _792_ (.A(_067_),
    .B(_370_),
    .Y(_371_));
 sg13g2_o21ai_1 _793_ (.B1(net42),
    .Y(_372_),
    .A1(_067_),
    .A2(_370_));
 sg13g2_a21oi_1 _794_ (.A1(_067_),
    .A2(_370_),
    .Y(_040_),
    .B1(_372_));
 sg13g2_nor2_1 _795_ (.A(_020_),
    .B(_370_),
    .Y(_373_));
 sg13g2_o21ai_1 _796_ (.B1(net42),
    .Y(_374_),
    .A1(\counter[5] ),
    .A2(_373_));
 sg13g2_a21oi_1 _797_ (.A1(\counter[5] ),
    .A2(_373_),
    .Y(_041_),
    .B1(_374_));
 sg13g2_nand2_1 _798_ (.Y(_375_),
    .A(\counter[5] ),
    .B(_371_));
 sg13g2_o21ai_1 _799_ (.B1(net42),
    .Y(_376_),
    .A1(_069_),
    .A2(_375_));
 sg13g2_a21oi_1 _800_ (.A1(_069_),
    .A2(_375_),
    .Y(_042_),
    .B1(_376_));
 sg13g2_nor2_1 _801_ (.A(_022_),
    .B(_375_),
    .Y(_377_));
 sg13g2_o21ai_1 _802_ (.B1(net42),
    .Y(_378_),
    .A1(\counter[7] ),
    .A2(_377_));
 sg13g2_a21oi_1 _803_ (.A1(\counter[7] ),
    .A2(_377_),
    .Y(_043_),
    .B1(_378_));
 sg13g2_and4_1 _804_ (.A(\counter[5] ),
    .B(\counter[6] ),
    .C(\counter[7] ),
    .D(_371_),
    .X(_379_));
 sg13g2_or2_1 _805_ (.X(_380_),
    .B(_379_),
    .A(\counter[8] ));
 sg13g2_nand2_1 _806_ (.Y(_381_),
    .A(\counter[8] ),
    .B(_379_));
 sg13g2_and3_1 _807_ (.X(_044_),
    .A(net42),
    .B(_380_),
    .C(_381_));
 sg13g2_o21ai_1 _808_ (.B1(net42),
    .Y(_382_),
    .A1(_071_),
    .A2(_381_));
 sg13g2_a21oi_1 _809_ (.A1(_071_),
    .A2(_381_),
    .Y(_045_),
    .B1(_382_));
 sg13g2_nand2_1 _810_ (.Y(_383_),
    .A(net39),
    .B(net34));
 sg13g2_nor3_1 _811_ (.A(net37),
    .B(net38),
    .C(\hvsync_gen.vpos[8] ),
    .Y(_384_));
 sg13g2_nand2_1 _812_ (.Y(_385_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_384_));
 sg13g2_nor3_1 _813_ (.A(\hvsync_gen.vpos[7] ),
    .B(\hvsync_gen.vpos[6] ),
    .C(_090_),
    .Y(_386_));
 sg13g2_nand3_1 _814_ (.B(\hvsync_gen.vpos[2] ),
    .C(_386_),
    .A(\hvsync_gen.vpos[3] ),
    .Y(_387_));
 sg13g2_o21ai_1 _815_ (.B1(net43),
    .Y(_388_),
    .A1(_385_),
    .A2(_387_));
 sg13g2_inv_1 _816_ (.Y(_389_),
    .A(_388_));
 sg13g2_nand2_2 _817_ (.Y(_390_),
    .A(_348_),
    .B(_389_));
 sg13g2_o21ai_1 _818_ (.B1(_383_),
    .Y(_046_),
    .A1(_056_),
    .A2(_390_));
 sg13g2_nand2_1 _819_ (.Y(_391_),
    .A(net89),
    .B(net35));
 sg13g2_o21ai_1 _820_ (.B1(_391_),
    .Y(_047_),
    .A1(_132_),
    .A2(_390_));
 sg13g2_nor2_1 _821_ (.A(_131_),
    .B(net34),
    .Y(_392_));
 sg13g2_nor2_2 _822_ (.A(net34),
    .B(_389_),
    .Y(_393_));
 sg13g2_xnor2_1 _823_ (.Y(_394_),
    .A(net103),
    .B(_392_));
 sg13g2_nor2_1 _824_ (.A(_393_),
    .B(_394_),
    .Y(_048_));
 sg13g2_nand2_1 _825_ (.Y(_395_),
    .A(\hvsync_gen.vpos[3] ),
    .B(_349_));
 sg13g2_nor2_1 _826_ (.A(net86),
    .B(_131_),
    .Y(_396_));
 sg13g2_xnor2_1 _827_ (.Y(_397_),
    .A(\hvsync_gen.vpos[3] ),
    .B(_396_));
 sg13g2_o21ai_1 _828_ (.B1(_395_),
    .Y(_049_),
    .A1(_390_),
    .A2(net87));
 sg13g2_nand2_1 _829_ (.Y(_398_),
    .A(net38),
    .B(net34));
 sg13g2_nand4_1 _830_ (.B(\hvsync_gen.vpos[1] ),
    .C(\hvsync_gen.vpos[3] ),
    .A(net39),
    .Y(_399_),
    .D(\hvsync_gen.vpos[2] ));
 sg13g2_xnor2_1 _831_ (.Y(_400_),
    .A(net74),
    .B(_399_));
 sg13g2_o21ai_1 _832_ (.B1(_398_),
    .Y(_050_),
    .A1(_390_),
    .A2(_400_));
 sg13g2_nand2_1 _833_ (.Y(_401_),
    .A(net37),
    .B(net34));
 sg13g2_o21ai_1 _834_ (.B1(_058_),
    .Y(_402_),
    .A1(_059_),
    .A2(_399_));
 sg13g2_or2_1 _835_ (.X(_403_),
    .B(_399_),
    .A(_085_));
 sg13g2_nand2_1 _836_ (.Y(_404_),
    .A(_402_),
    .B(_403_));
 sg13g2_o21ai_1 _837_ (.B1(_401_),
    .Y(_051_),
    .A1(_390_),
    .A2(_404_));
 sg13g2_nor2_1 _838_ (.A(net34),
    .B(_403_),
    .Y(_405_));
 sg13g2_xnor2_1 _839_ (.Y(_406_),
    .A(net97),
    .B(_405_));
 sg13g2_nor2_1 _840_ (.A(_393_),
    .B(_406_),
    .Y(_052_));
 sg13g2_nand2_1 _841_ (.Y(_407_),
    .A(\hvsync_gen.vpos[7] ),
    .B(net34));
 sg13g2_nor2_1 _842_ (.A(net81),
    .B(_403_),
    .Y(_408_));
 sg13g2_xnor2_1 _843_ (.Y(_409_),
    .A(\hvsync_gen.vpos[7] ),
    .B(_408_));
 sg13g2_o21ai_1 _844_ (.B1(_407_),
    .Y(_053_),
    .A1(_390_),
    .A2(net82));
 sg13g2_nand3_1 _845_ (.B(net104),
    .C(_405_),
    .A(\hvsync_gen.vpos[7] ),
    .Y(_410_));
 sg13g2_xor2_1 _846_ (.B(_410_),
    .A(net92),
    .X(_411_));
 sg13g2_nor2_1 _847_ (.A(_393_),
    .B(_411_),
    .Y(_054_));
 sg13g2_nand2_1 _848_ (.Y(_412_),
    .A(net95),
    .B(net35));
 sg13g2_nor3_1 _849_ (.A(_010_),
    .B(_086_),
    .C(_399_),
    .Y(_413_));
 sg13g2_xnor2_1 _850_ (.Y(_414_),
    .A(net95),
    .B(_413_));
 sg13g2_o21ai_1 _851_ (.B1(_412_),
    .Y(_055_),
    .A1(_390_),
    .A2(_414_));
 sg13g2_dfrbp_1 _852_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net55),
    .D(_026_),
    .Q_N(_025_),
    .Q(\dist_x[0] ));
 sg13g2_dfrbp_1 _853_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net30),
    .D(_027_),
    .Q_N(_007_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 _854_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net29),
    .D(_028_),
    .Q_N(_004_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 _855_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net28),
    .D(_029_),
    .Q_N(_017_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 _856_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net27),
    .D(_030_),
    .Q_N(_016_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 _857_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net26),
    .D(net91),
    .Q_N(_014_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 _858_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net25),
    .D(_032_),
    .Q_N(_013_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 _859_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net65),
    .D(net77),
    .Q_N(_011_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 _860_ (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net64),
    .D(_034_),
    .Q_N(_009_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 _861_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net63),
    .D(net80),
    .Q_N(_002_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 _862_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net62),
    .D(_036_),
    .Q_N(_024_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 _863_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net61),
    .D(_037_),
    .Q_N(_006_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 _864_ (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net60),
    .D(_038_),
    .Q_N(_003_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 _865_ (.CLK(net36),
    .RESET_B(net59),
    .D(_039_),
    .Q_N(_019_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 _866_ (.CLK(net36),
    .RESET_B(net58),
    .D(_040_),
    .Q_N(_020_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 _867_ (.CLK(net36),
    .RESET_B(net57),
    .D(_041_),
    .Q_N(_021_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 _868_ (.CLK(net36),
    .RESET_B(net56),
    .D(_042_),
    .Q_N(_022_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 _869_ (.CLK(net36),
    .RESET_B(net54),
    .D(_043_),
    .Q_N(_420_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 _870_ (.CLK(net36),
    .RESET_B(net53),
    .D(_044_),
    .Q_N(_419_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 _871_ (.CLK(net36),
    .RESET_B(net66),
    .D(_045_),
    .Q_N(_421_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 _872_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net52),
    .D(net72),
    .Q_N(_418_),
    .Q(hsync));
 sg13g2_dfrbp_1 _873_ (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net51),
    .D(net68),
    .Q_N(_023_),
    .Q(\dist_y[0] ));
 sg13g2_dfrbp_1 _874_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net49),
    .D(_047_),
    .Q_N(_008_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 _875_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net47),
    .D(_048_),
    .Q_N(_005_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 _876_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net45),
    .D(net88),
    .Q_N(_018_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 _877_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net33),
    .D(net75),
    .Q_N(_015_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 _878_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net31),
    .D(_051_),
    .Q_N(_417_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 _879_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net48),
    .D(_052_),
    .Q_N(_012_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 _880_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net44),
    .D(net83),
    .Q_N(_416_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 _881_ (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net50),
    .D(_054_),
    .Q_N(_010_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 _882_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net46),
    .D(net96),
    .Q_N(_422_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 _883_ (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net32),
    .D(net94),
    .Q_N(_415_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_tiehi _857__26 (.L_HI(net26));
 sg13g2_tiehi _856__27 (.L_HI(net27));
 sg13g2_tiehi _855__28 (.L_HI(net28));
 sg13g2_tiehi _854__29 (.L_HI(net29));
 sg13g2_tiehi _853__30 (.L_HI(net30));
 sg13g2_tiehi _878__31 (.L_HI(net31));
 sg13g2_tiehi _883__32 (.L_HI(net32));
 sg13g2_tiehi _877__33 (.L_HI(net33));
 sg13g2_tiehi _880__34 (.L_HI(net44));
 sg13g2_tiehi _876__35 (.L_HI(net45));
 sg13g2_tiehi _882__36 (.L_HI(net46));
 sg13g2_tiehi _875__37 (.L_HI(net47));
 sg13g2_tiehi _879__38 (.L_HI(net48));
 sg13g2_tiehi _874__39 (.L_HI(net49));
 sg13g2_tiehi _881__40 (.L_HI(net50));
 sg13g2_tiehi _873__41 (.L_HI(net51));
 sg13g2_tiehi _872__42 (.L_HI(net52));
 sg13g2_tiehi _870__43 (.L_HI(net53));
 sg13g2_tiehi _869__44 (.L_HI(net54));
 sg13g2_tiehi _852__45 (.L_HI(net55));
 sg13g2_tiehi _868__46 (.L_HI(net56));
 sg13g2_tiehi _867__47 (.L_HI(net57));
 sg13g2_tiehi _866__48 (.L_HI(net58));
 sg13g2_tiehi _865__49 (.L_HI(net59));
 sg13g2_tiehi _864__50 (.L_HI(net60));
 sg13g2_tiehi _863__51 (.L_HI(net61));
 sg13g2_tiehi _862__52 (.L_HI(net62));
 sg13g2_tiehi _861__53 (.L_HI(net63));
 sg13g2_tiehi _860__54 (.L_HI(net64));
 sg13g2_tiehi _859__55 (.L_HI(net65));
 sg13g2_tiehi _871__56 (.L_HI(net66));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_bleeptrack_prism_10 (.L_LO(net10));
 sg13g2_tielo tt_um_bleeptrack_prism_11 (.L_LO(net11));
 sg13g2_tielo tt_um_bleeptrack_prism_12 (.L_LO(net12));
 sg13g2_tielo tt_um_bleeptrack_prism_13 (.L_LO(net13));
 sg13g2_tielo tt_um_bleeptrack_prism_14 (.L_LO(net14));
 sg13g2_tielo tt_um_bleeptrack_prism_15 (.L_LO(net15));
 sg13g2_tielo tt_um_bleeptrack_prism_16 (.L_LO(net16));
 sg13g2_tielo tt_um_bleeptrack_prism_17 (.L_LO(net17));
 sg13g2_tielo tt_um_bleeptrack_prism_18 (.L_LO(net18));
 sg13g2_tielo tt_um_bleeptrack_prism_19 (.L_LO(net19));
 sg13g2_tielo tt_um_bleeptrack_prism_20 (.L_LO(net20));
 sg13g2_tielo tt_um_bleeptrack_prism_21 (.L_LO(net21));
 sg13g2_tielo tt_um_bleeptrack_prism_22 (.L_LO(net22));
 sg13g2_tielo tt_um_bleeptrack_prism_23 (.L_LO(net23));
 sg13g2_tielo tt_um_bleeptrack_prism_24 (.L_LO(net24));
 sg13g2_tiehi _858__25 (.L_HI(net25));
 sg13g2_buf_1 _932_ (.A(net36),
    .X(uo_out[3]));
 sg13g2_buf_1 _933_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout34 (.A(net35),
    .X(net34));
 sg13g2_buf_4 fanout35 (.X(net35),
    .A(_349_));
 sg13g2_buf_2 fanout36 (.A(\hvsync_gen.vsync ),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(net100),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(\hvsync_gen.vpos[4] ),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(\dist_y[0] ),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(\hvsync_gen.hpos[9] ),
    .X(net40));
 sg13g2_buf_4 fanout41 (.X(net41),
    .A(\dist_x[0] ));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(net43));
 sg13g2_buf_4 fanout43 (.X(net43),
    .A(rst_n));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_bleeptrack_prism_9 (.L_LO(net9));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(_023_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold2 (.A(_046_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold3 (.A(_025_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold4 (.A(_002_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold5 (.A(_081_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold6 (.A(_000_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold7 (.A(\hvsync_gen.hpos[6] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold8 (.A(_015_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold9 (.A(_050_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold10 (.A(\hvsync_gen.hpos[7] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold11 (.A(_033_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold12 (.A(\hvsync_gen.hpos[2] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold13 (.A(_009_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold14 (.A(_035_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold15 (.A(_012_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold16 (.A(_409_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold17 (.A(_053_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold18 (.A(\dist_x[0] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold19 (.A(_126_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold20 (.A(_005_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold21 (.A(_397_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold22 (.A(_049_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold23 (.A(\hvsync_gen.vpos[1] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold24 (.A(_016_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold25 (.A(_031_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold26 (.A(\hvsync_gen.vpos[8] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold27 (.A(\hvsync_gen.vpos[3] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold28 (.A(_001_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold29 (.A(\hvsync_gen.vpos[9] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold30 (.A(_055_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold31 (.A(\hvsync_gen.vpos[6] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold32 (.A(\hvsync_gen.hpos[3] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold33 (.A(_353_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold34 (.A(\hvsync_gen.vpos[5] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold35 (.A(\hvsync_gen.hpos[8] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold36 (.A(\hvsync_gen.hpos[4] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold37 (.A(\hvsync_gen.vpos[2] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold38 (.A(\hvsync_gen.vpos[6] ),
    .X(net104));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_215 ();
 sg13g2_decap_8 FILLER_17_222 ();
 sg13g2_decap_8 FILLER_17_229 ();
 sg13g2_decap_4 FILLER_17_236 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_4 FILLER_18_196 ();
 sg13g2_decap_4 FILLER_18_226 ();
 sg13g2_fill_2 FILLER_18_256 ();
 sg13g2_fill_1 FILLER_18_258 ();
 sg13g2_decap_4 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_296 ();
 sg13g2_decap_8 FILLER_18_303 ();
 sg13g2_fill_2 FILLER_18_310 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_8 FILLER_18_332 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_360 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_388 ();
 sg13g2_decap_8 FILLER_18_395 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_fill_2 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_174 ();
 sg13g2_decap_8 FILLER_19_181 ();
 sg13g2_decap_4 FILLER_19_188 ();
 sg13g2_fill_2 FILLER_19_192 ();
 sg13g2_fill_2 FILLER_19_225 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_decap_4 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_248 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_decap_4 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_331 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_4 FILLER_20_140 ();
 sg13g2_fill_2 FILLER_20_144 ();
 sg13g2_fill_2 FILLER_20_172 ();
 sg13g2_fill_1 FILLER_20_174 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_2 FILLER_20_224 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_fill_1 FILLER_20_232 ();
 sg13g2_fill_2 FILLER_20_249 ();
 sg13g2_decap_4 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_292 ();
 sg13g2_fill_2 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_303 ();
 sg13g2_fill_2 FILLER_20_312 ();
 sg13g2_fill_2 FILLER_20_337 ();
 sg13g2_fill_1 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_fill_1 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_384 ();
 sg13g2_decap_8 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_fill_1 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_fill_2 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_193 ();
 sg13g2_fill_2 FILLER_21_225 ();
 sg13g2_decap_8 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_decap_4 FILLER_21_284 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_fill_2 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_395 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_4 FILLER_22_133 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_164 ();
 sg13g2_fill_2 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_216 ();
 sg13g2_decap_4 FILLER_22_239 ();
 sg13g2_fill_1 FILLER_22_243 ();
 sg13g2_fill_1 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_254 ();
 sg13g2_fill_2 FILLER_22_261 ();
 sg13g2_fill_1 FILLER_22_263 ();
 sg13g2_fill_2 FILLER_22_310 ();
 sg13g2_decap_8 FILLER_22_381 ();
 sg13g2_decap_4 FILLER_22_388 ();
 sg13g2_fill_1 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_4 FILLER_23_112 ();
 sg13g2_fill_1 FILLER_23_116 ();
 sg13g2_decap_4 FILLER_23_121 ();
 sg13g2_fill_1 FILLER_23_125 ();
 sg13g2_fill_2 FILLER_23_157 ();
 sg13g2_fill_1 FILLER_23_159 ();
 sg13g2_decap_8 FILLER_23_173 ();
 sg13g2_decap_8 FILLER_23_195 ();
 sg13g2_fill_2 FILLER_23_226 ();
 sg13g2_decap_8 FILLER_23_236 ();
 sg13g2_fill_2 FILLER_23_243 ();
 sg13g2_decap_4 FILLER_23_250 ();
 sg13g2_fill_1 FILLER_23_254 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_fill_1 FILLER_23_274 ();
 sg13g2_fill_2 FILLER_23_279 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_decap_8 FILLER_23_290 ();
 sg13g2_decap_4 FILLER_23_297 ();
 sg13g2_decap_4 FILLER_23_306 ();
 sg13g2_fill_1 FILLER_23_314 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_fill_2 FILLER_23_336 ();
 sg13g2_decap_4 FILLER_23_351 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_fill_2 FILLER_23_371 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_105 ();
 sg13g2_fill_1 FILLER_24_132 ();
 sg13g2_fill_2 FILLER_24_142 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_201 ();
 sg13g2_decap_8 FILLER_24_218 ();
 sg13g2_decap_4 FILLER_24_225 ();
 sg13g2_fill_1 FILLER_24_229 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_fill_2 FILLER_24_271 ();
 sg13g2_fill_1 FILLER_24_273 ();
 sg13g2_fill_1 FILLER_24_279 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_fill_1 FILLER_24_369 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_4 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_123 ();
 sg13g2_fill_1 FILLER_25_156 ();
 sg13g2_fill_1 FILLER_25_174 ();
 sg13g2_decap_8 FILLER_25_179 ();
 sg13g2_decap_8 FILLER_25_186 ();
 sg13g2_decap_8 FILLER_25_193 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_decap_8 FILLER_25_207 ();
 sg13g2_decap_4 FILLER_25_214 ();
 sg13g2_fill_2 FILLER_25_218 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_4 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_decap_4 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_254 ();
 sg13g2_decap_8 FILLER_25_274 ();
 sg13g2_fill_2 FILLER_25_281 ();
 sg13g2_fill_1 FILLER_25_283 ();
 sg13g2_decap_4 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_4 FILLER_25_333 ();
 sg13g2_fill_1 FILLER_25_337 ();
 sg13g2_fill_2 FILLER_25_376 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_fill_2 FILLER_26_98 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_fill_2 FILLER_26_127 ();
 sg13g2_fill_1 FILLER_26_129 ();
 sg13g2_fill_2 FILLER_26_139 ();
 sg13g2_fill_2 FILLER_26_158 ();
 sg13g2_decap_4 FILLER_26_180 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_decap_8 FILLER_26_208 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_fill_1 FILLER_26_304 ();
 sg13g2_fill_1 FILLER_26_331 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_decap_4 FILLER_26_364 ();
 sg13g2_fill_1 FILLER_26_368 ();
 sg13g2_decap_4 FILLER_26_372 ();
 sg13g2_fill_2 FILLER_26_376 ();
 sg13g2_fill_2 FILLER_26_386 ();
 sg13g2_fill_1 FILLER_26_388 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_105 ();
 sg13g2_fill_2 FILLER_27_124 ();
 sg13g2_fill_1 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_149 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_fill_2 FILLER_27_174 ();
 sg13g2_fill_1 FILLER_27_181 ();
 sg13g2_decap_8 FILLER_27_187 ();
 sg13g2_fill_2 FILLER_27_194 ();
 sg13g2_fill_1 FILLER_27_196 ();
 sg13g2_fill_1 FILLER_27_208 ();
 sg13g2_decap_8 FILLER_27_213 ();
 sg13g2_fill_2 FILLER_27_227 ();
 sg13g2_fill_1 FILLER_27_256 ();
 sg13g2_decap_4 FILLER_27_261 ();
 sg13g2_fill_2 FILLER_27_265 ();
 sg13g2_decap_8 FILLER_27_275 ();
 sg13g2_fill_2 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_292 ();
 sg13g2_fill_2 FILLER_27_299 ();
 sg13g2_fill_1 FILLER_27_301 ();
 sg13g2_decap_4 FILLER_27_305 ();
 sg13g2_decap_8 FILLER_27_320 ();
 sg13g2_decap_8 FILLER_27_331 ();
 sg13g2_fill_2 FILLER_27_338 ();
 sg13g2_decap_4 FILLER_27_348 ();
 sg13g2_fill_1 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_4 FILLER_27_365 ();
 sg13g2_fill_1 FILLER_27_369 ();
 sg13g2_fill_2 FILLER_27_382 ();
 sg13g2_fill_2 FILLER_27_394 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_4 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_183 ();
 sg13g2_fill_2 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_199 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_decap_8 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_229 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_decap_4 FILLER_28_249 ();
 sg13g2_fill_2 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_fill_2 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_decap_4 FILLER_28_342 ();
 sg13g2_fill_2 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_375 ();
 sg13g2_fill_1 FILLER_28_381 ();
 sg13g2_fill_1 FILLER_28_392 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_4 FILLER_29_112 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_fill_2 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_decap_4 FILLER_29_181 ();
 sg13g2_decap_8 FILLER_29_199 ();
 sg13g2_fill_1 FILLER_29_206 ();
 sg13g2_fill_1 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_fill_1 FILLER_29_222 ();
 sg13g2_fill_2 FILLER_29_237 ();
 sg13g2_fill_1 FILLER_29_239 ();
 sg13g2_decap_8 FILLER_29_260 ();
 sg13g2_fill_2 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_269 ();
 sg13g2_fill_2 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_276 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_decap_8 FILLER_29_292 ();
 sg13g2_fill_2 FILLER_29_299 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_decap_8 FILLER_29_324 ();
 sg13g2_decap_4 FILLER_29_331 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_decap_8 FILLER_29_359 ();
 sg13g2_decap_4 FILLER_29_366 ();
 sg13g2_fill_2 FILLER_29_370 ();
 sg13g2_fill_2 FILLER_29_385 ();
 sg13g2_fill_1 FILLER_29_387 ();
 sg13g2_fill_1 FILLER_29_396 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_decap_8 FILLER_30_179 ();
 sg13g2_fill_2 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_188 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_220 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_decap_4 FILLER_30_251 ();
 sg13g2_decap_4 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_fill_2 FILLER_30_275 ();
 sg13g2_fill_1 FILLER_30_277 ();
 sg13g2_decap_8 FILLER_30_286 ();
 sg13g2_decap_8 FILLER_30_293 ();
 sg13g2_decap_4 FILLER_30_300 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_decap_4 FILLER_30_319 ();
 sg13g2_fill_2 FILLER_30_323 ();
 sg13g2_fill_2 FILLER_30_337 ();
 sg13g2_fill_1 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_fill_2 FILLER_30_350 ();
 sg13g2_fill_1 FILLER_30_352 ();
 sg13g2_decap_4 FILLER_30_361 ();
 sg13g2_fill_2 FILLER_30_365 ();
 sg13g2_fill_2 FILLER_30_372 ();
 sg13g2_fill_1 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_fill_1 FILLER_30_396 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_197 ();
 sg13g2_fill_2 FILLER_31_204 ();
 sg13g2_decap_8 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_220 ();
 sg13g2_fill_2 FILLER_31_227 ();
 sg13g2_decap_8 FILLER_31_239 ();
 sg13g2_decap_8 FILLER_31_246 ();
 sg13g2_decap_8 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_267 ();
 sg13g2_fill_1 FILLER_31_269 ();
 sg13g2_decap_8 FILLER_31_277 ();
 sg13g2_decap_8 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_291 ();
 sg13g2_fill_1 FILLER_31_293 ();
 sg13g2_decap_4 FILLER_31_315 ();
 sg13g2_fill_1 FILLER_31_319 ();
 sg13g2_decap_8 FILLER_31_332 ();
 sg13g2_fill_2 FILLER_31_339 ();
 sg13g2_fill_1 FILLER_31_341 ();
 sg13g2_fill_2 FILLER_31_356 ();
 sg13g2_decap_4 FILLER_31_366 ();
 sg13g2_fill_1 FILLER_31_378 ();
 sg13g2_fill_2 FILLER_31_388 ();
 sg13g2_fill_1 FILLER_31_390 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_4 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_decap_4 FILLER_32_195 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_4 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_240 ();
 sg13g2_decap_4 FILLER_32_246 ();
 sg13g2_decap_4 FILLER_32_282 ();
 sg13g2_decap_8 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_decap_4 FILLER_32_372 ();
 sg13g2_fill_1 FILLER_32_376 ();
 sg13g2_fill_2 FILLER_32_394 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_4 FILLER_33_182 ();
 sg13g2_fill_1 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_fill_2 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_242 ();
 sg13g2_fill_2 FILLER_33_249 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_fill_1 FILLER_33_258 ();
 sg13g2_decap_8 FILLER_33_262 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_fill_1 FILLER_33_282 ();
 sg13g2_decap_4 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_292 ();
 sg13g2_fill_1 FILLER_33_306 ();
 sg13g2_fill_2 FILLER_33_328 ();
 sg13g2_fill_1 FILLER_33_330 ();
 sg13g2_decap_8 FILLER_33_349 ();
 sg13g2_fill_1 FILLER_33_356 ();
 sg13g2_decap_8 FILLER_33_365 ();
 sg13g2_decap_4 FILLER_33_372 ();
 sg13g2_fill_1 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_187 ();
 sg13g2_decap_8 FILLER_34_202 ();
 sg13g2_fill_2 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_211 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_fill_1 FILLER_34_231 ();
 sg13g2_decap_4 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_253 ();
 sg13g2_decap_4 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_272 ();
 sg13g2_decap_8 FILLER_34_278 ();
 sg13g2_decap_4 FILLER_34_285 ();
 sg13g2_fill_2 FILLER_34_289 ();
 sg13g2_decap_8 FILLER_34_298 ();
 sg13g2_decap_4 FILLER_34_323 ();
 sg13g2_fill_2 FILLER_34_327 ();
 sg13g2_fill_1 FILLER_34_337 ();
 sg13g2_decap_4 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_354 ();
 sg13g2_decap_4 FILLER_34_373 ();
 sg13g2_fill_1 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_387 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_4 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_176 ();
 sg13g2_decap_8 FILLER_35_183 ();
 sg13g2_decap_8 FILLER_35_194 ();
 sg13g2_decap_8 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_fill_2 FILLER_35_231 ();
 sg13g2_fill_1 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_247 ();
 sg13g2_fill_1 FILLER_35_280 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_decap_4 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_decap_8 FILLER_35_313 ();
 sg13g2_decap_8 FILLER_35_320 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_fill_2 FILLER_35_355 ();
 sg13g2_fill_1 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_4 FILLER_36_154 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_fill_2 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_decap_4 FILLER_36_207 ();
 sg13g2_fill_2 FILLER_36_211 ();
 sg13g2_decap_8 FILLER_36_225 ();
 sg13g2_fill_2 FILLER_36_232 ();
 sg13g2_decap_8 FILLER_36_237 ();
 sg13g2_decap_4 FILLER_36_244 ();
 sg13g2_decap_8 FILLER_36_253 ();
 sg13g2_decap_8 FILLER_36_260 ();
 sg13g2_decap_8 FILLER_36_267 ();
 sg13g2_fill_2 FILLER_36_274 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_decap_4 FILLER_36_281 ();
 sg13g2_decap_8 FILLER_36_295 ();
 sg13g2_decap_4 FILLER_36_302 ();
 sg13g2_decap_8 FILLER_36_314 ();
 sg13g2_decap_8 FILLER_36_321 ();
 sg13g2_fill_2 FILLER_36_328 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_fill_2 FILLER_36_366 ();
 sg13g2_fill_1 FILLER_36_374 ();
 sg13g2_decap_4 FILLER_36_379 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_fill_2 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_178 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_decap_8 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_fill_2 FILLER_37_241 ();
 sg13g2_fill_1 FILLER_37_243 ();
 sg13g2_fill_2 FILLER_37_270 ();
 sg13g2_fill_1 FILLER_37_272 ();
 sg13g2_fill_1 FILLER_37_290 ();
 sg13g2_fill_2 FILLER_37_348 ();
 sg13g2_fill_1 FILLER_37_350 ();
 sg13g2_fill_1 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_fill_1 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_fill_2 FILLER_38_223 ();
 sg13g2_fill_1 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_230 ();
 sg13g2_decap_8 FILLER_38_237 ();
 sg13g2_fill_2 FILLER_38_244 ();
 sg13g2_fill_1 FILLER_38_246 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_254 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_fill_2 FILLER_38_280 ();
 sg13g2_fill_1 FILLER_38_282 ();
 sg13g2_decap_8 FILLER_38_291 ();
 sg13g2_decap_4 FILLER_38_298 ();
 sg13g2_decap_4 FILLER_38_306 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_decap_4 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_376 ();
 sg13g2_decap_8 FILLER_38_383 ();
 sg13g2_decap_4 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule
