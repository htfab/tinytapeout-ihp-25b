module tt_um_urish_sic1 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \A[0] ;
 wire \A[1] ;
 wire \A[2] ;
 wire \A[3] ;
 wire \A[4] ;
 wire \A[5] ;
 wire \A[6] ;
 wire \A[7] ;
 wire \B[0] ;
 wire \B[1] ;
 wire \B[2] ;
 wire \B[3] ;
 wire \B[4] ;
 wire \B[5] ;
 wire \B[6] ;
 wire \B[7] ;
 wire \C[0] ;
 wire \C[1] ;
 wire \C[2] ;
 wire \C[3] ;
 wire \C[4] ;
 wire \C[5] ;
 wire \C[6] ;
 wire \C[7] ;
 wire \PC[0] ;
 wire \PC[1] ;
 wire \PC[2] ;
 wire \PC[3] ;
 wire \PC[4] ;
 wire \PC[5] ;
 wire \PC[6] ;
 wire \PC[7] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire halted;
 wire \mem.addr[0] ;
 wire \mem.addr[1] ;
 wire \mem.addr[2] ;
 wire \mem.addr[3] ;
 wire \mem.addr[4] ;
 wire \mem.addr[5] ;
 wire \mem.addr[6] ;
 wire \mem.addr[7] ;
 wire \mem.data_in[0] ;
 wire \mem.data_in[1] ;
 wire \mem.data_in[2] ;
 wire \mem.data_in[3] ;
 wire \mem.data_in[4] ;
 wire \mem.data_in[5] ;
 wire \mem.data_in[6] ;
 wire \mem.data_in[7] ;
 wire \mem.mem[0][0] ;
 wire \mem.mem[0][1] ;
 wire \mem.mem[0][2] ;
 wire \mem.mem[0][3] ;
 wire \mem.mem[0][4] ;
 wire \mem.mem[0][5] ;
 wire \mem.mem[0][6] ;
 wire \mem.mem[0][7] ;
 wire \mem.mem[100][0] ;
 wire \mem.mem[100][1] ;
 wire \mem.mem[100][2] ;
 wire \mem.mem[100][3] ;
 wire \mem.mem[100][4] ;
 wire \mem.mem[100][5] ;
 wire \mem.mem[100][6] ;
 wire \mem.mem[100][7] ;
 wire \mem.mem[101][0] ;
 wire \mem.mem[101][1] ;
 wire \mem.mem[101][2] ;
 wire \mem.mem[101][3] ;
 wire \mem.mem[101][4] ;
 wire \mem.mem[101][5] ;
 wire \mem.mem[101][6] ;
 wire \mem.mem[101][7] ;
 wire \mem.mem[102][0] ;
 wire \mem.mem[102][1] ;
 wire \mem.mem[102][2] ;
 wire \mem.mem[102][3] ;
 wire \mem.mem[102][4] ;
 wire \mem.mem[102][5] ;
 wire \mem.mem[102][6] ;
 wire \mem.mem[102][7] ;
 wire \mem.mem[103][0] ;
 wire \mem.mem[103][1] ;
 wire \mem.mem[103][2] ;
 wire \mem.mem[103][3] ;
 wire \mem.mem[103][4] ;
 wire \mem.mem[103][5] ;
 wire \mem.mem[103][6] ;
 wire \mem.mem[103][7] ;
 wire \mem.mem[104][0] ;
 wire \mem.mem[104][1] ;
 wire \mem.mem[104][2] ;
 wire \mem.mem[104][3] ;
 wire \mem.mem[104][4] ;
 wire \mem.mem[104][5] ;
 wire \mem.mem[104][6] ;
 wire \mem.mem[104][7] ;
 wire \mem.mem[105][0] ;
 wire \mem.mem[105][1] ;
 wire \mem.mem[105][2] ;
 wire \mem.mem[105][3] ;
 wire \mem.mem[105][4] ;
 wire \mem.mem[105][5] ;
 wire \mem.mem[105][6] ;
 wire \mem.mem[105][7] ;
 wire \mem.mem[106][0] ;
 wire \mem.mem[106][1] ;
 wire \mem.mem[106][2] ;
 wire \mem.mem[106][3] ;
 wire \mem.mem[106][4] ;
 wire \mem.mem[106][5] ;
 wire \mem.mem[106][6] ;
 wire \mem.mem[106][7] ;
 wire \mem.mem[107][0] ;
 wire \mem.mem[107][1] ;
 wire \mem.mem[107][2] ;
 wire \mem.mem[107][3] ;
 wire \mem.mem[107][4] ;
 wire \mem.mem[107][5] ;
 wire \mem.mem[107][6] ;
 wire \mem.mem[107][7] ;
 wire \mem.mem[108][0] ;
 wire \mem.mem[108][1] ;
 wire \mem.mem[108][2] ;
 wire \mem.mem[108][3] ;
 wire \mem.mem[108][4] ;
 wire \mem.mem[108][5] ;
 wire \mem.mem[108][6] ;
 wire \mem.mem[108][7] ;
 wire \mem.mem[109][0] ;
 wire \mem.mem[109][1] ;
 wire \mem.mem[109][2] ;
 wire \mem.mem[109][3] ;
 wire \mem.mem[109][4] ;
 wire \mem.mem[109][5] ;
 wire \mem.mem[109][6] ;
 wire \mem.mem[109][7] ;
 wire \mem.mem[10][0] ;
 wire \mem.mem[10][1] ;
 wire \mem.mem[10][2] ;
 wire \mem.mem[10][3] ;
 wire \mem.mem[10][4] ;
 wire \mem.mem[10][5] ;
 wire \mem.mem[10][6] ;
 wire \mem.mem[10][7] ;
 wire \mem.mem[110][0] ;
 wire \mem.mem[110][1] ;
 wire \mem.mem[110][2] ;
 wire \mem.mem[110][3] ;
 wire \mem.mem[110][4] ;
 wire \mem.mem[110][5] ;
 wire \mem.mem[110][6] ;
 wire \mem.mem[110][7] ;
 wire \mem.mem[111][0] ;
 wire \mem.mem[111][1] ;
 wire \mem.mem[111][2] ;
 wire \mem.mem[111][3] ;
 wire \mem.mem[111][4] ;
 wire \mem.mem[111][5] ;
 wire \mem.mem[111][6] ;
 wire \mem.mem[111][7] ;
 wire \mem.mem[112][0] ;
 wire \mem.mem[112][1] ;
 wire \mem.mem[112][2] ;
 wire \mem.mem[112][3] ;
 wire \mem.mem[112][4] ;
 wire \mem.mem[112][5] ;
 wire \mem.mem[112][6] ;
 wire \mem.mem[112][7] ;
 wire \mem.mem[113][0] ;
 wire \mem.mem[113][1] ;
 wire \mem.mem[113][2] ;
 wire \mem.mem[113][3] ;
 wire \mem.mem[113][4] ;
 wire \mem.mem[113][5] ;
 wire \mem.mem[113][6] ;
 wire \mem.mem[113][7] ;
 wire \mem.mem[114][0] ;
 wire \mem.mem[114][1] ;
 wire \mem.mem[114][2] ;
 wire \mem.mem[114][3] ;
 wire \mem.mem[114][4] ;
 wire \mem.mem[114][5] ;
 wire \mem.mem[114][6] ;
 wire \mem.mem[114][7] ;
 wire \mem.mem[115][0] ;
 wire \mem.mem[115][1] ;
 wire \mem.mem[115][2] ;
 wire \mem.mem[115][3] ;
 wire \mem.mem[115][4] ;
 wire \mem.mem[115][5] ;
 wire \mem.mem[115][6] ;
 wire \mem.mem[115][7] ;
 wire \mem.mem[116][0] ;
 wire \mem.mem[116][1] ;
 wire \mem.mem[116][2] ;
 wire \mem.mem[116][3] ;
 wire \mem.mem[116][4] ;
 wire \mem.mem[116][5] ;
 wire \mem.mem[116][6] ;
 wire \mem.mem[116][7] ;
 wire \mem.mem[117][0] ;
 wire \mem.mem[117][1] ;
 wire \mem.mem[117][2] ;
 wire \mem.mem[117][3] ;
 wire \mem.mem[117][4] ;
 wire \mem.mem[117][5] ;
 wire \mem.mem[117][6] ;
 wire \mem.mem[117][7] ;
 wire \mem.mem[118][0] ;
 wire \mem.mem[118][1] ;
 wire \mem.mem[118][2] ;
 wire \mem.mem[118][3] ;
 wire \mem.mem[118][4] ;
 wire \mem.mem[118][5] ;
 wire \mem.mem[118][6] ;
 wire \mem.mem[118][7] ;
 wire \mem.mem[119][0] ;
 wire \mem.mem[119][1] ;
 wire \mem.mem[119][2] ;
 wire \mem.mem[119][3] ;
 wire \mem.mem[119][4] ;
 wire \mem.mem[119][5] ;
 wire \mem.mem[119][6] ;
 wire \mem.mem[119][7] ;
 wire \mem.mem[11][0] ;
 wire \mem.mem[11][1] ;
 wire \mem.mem[11][2] ;
 wire \mem.mem[11][3] ;
 wire \mem.mem[11][4] ;
 wire \mem.mem[11][5] ;
 wire \mem.mem[11][6] ;
 wire \mem.mem[11][7] ;
 wire \mem.mem[120][0] ;
 wire \mem.mem[120][1] ;
 wire \mem.mem[120][2] ;
 wire \mem.mem[120][3] ;
 wire \mem.mem[120][4] ;
 wire \mem.mem[120][5] ;
 wire \mem.mem[120][6] ;
 wire \mem.mem[120][7] ;
 wire \mem.mem[121][0] ;
 wire \mem.mem[121][1] ;
 wire \mem.mem[121][2] ;
 wire \mem.mem[121][3] ;
 wire \mem.mem[121][4] ;
 wire \mem.mem[121][5] ;
 wire \mem.mem[121][6] ;
 wire \mem.mem[121][7] ;
 wire \mem.mem[122][0] ;
 wire \mem.mem[122][1] ;
 wire \mem.mem[122][2] ;
 wire \mem.mem[122][3] ;
 wire \mem.mem[122][4] ;
 wire \mem.mem[122][5] ;
 wire \mem.mem[122][6] ;
 wire \mem.mem[122][7] ;
 wire \mem.mem[123][0] ;
 wire \mem.mem[123][1] ;
 wire \mem.mem[123][2] ;
 wire \mem.mem[123][3] ;
 wire \mem.mem[123][4] ;
 wire \mem.mem[123][5] ;
 wire \mem.mem[123][6] ;
 wire \mem.mem[123][7] ;
 wire \mem.mem[124][0] ;
 wire \mem.mem[124][1] ;
 wire \mem.mem[124][2] ;
 wire \mem.mem[124][3] ;
 wire \mem.mem[124][4] ;
 wire \mem.mem[124][5] ;
 wire \mem.mem[124][6] ;
 wire \mem.mem[124][7] ;
 wire \mem.mem[125][0] ;
 wire \mem.mem[125][1] ;
 wire \mem.mem[125][2] ;
 wire \mem.mem[125][3] ;
 wire \mem.mem[125][4] ;
 wire \mem.mem[125][5] ;
 wire \mem.mem[125][6] ;
 wire \mem.mem[125][7] ;
 wire \mem.mem[126][0] ;
 wire \mem.mem[126][1] ;
 wire \mem.mem[126][2] ;
 wire \mem.mem[126][3] ;
 wire \mem.mem[126][4] ;
 wire \mem.mem[126][5] ;
 wire \mem.mem[126][6] ;
 wire \mem.mem[126][7] ;
 wire \mem.mem[127][0] ;
 wire \mem.mem[127][1] ;
 wire \mem.mem[127][2] ;
 wire \mem.mem[127][3] ;
 wire \mem.mem[127][4] ;
 wire \mem.mem[127][5] ;
 wire \mem.mem[127][6] ;
 wire \mem.mem[127][7] ;
 wire \mem.mem[128][0] ;
 wire \mem.mem[128][1] ;
 wire \mem.mem[128][2] ;
 wire \mem.mem[128][3] ;
 wire \mem.mem[128][4] ;
 wire \mem.mem[128][5] ;
 wire \mem.mem[128][6] ;
 wire \mem.mem[128][7] ;
 wire \mem.mem[129][0] ;
 wire \mem.mem[129][1] ;
 wire \mem.mem[129][2] ;
 wire \mem.mem[129][3] ;
 wire \mem.mem[129][4] ;
 wire \mem.mem[129][5] ;
 wire \mem.mem[129][6] ;
 wire \mem.mem[129][7] ;
 wire \mem.mem[12][0] ;
 wire \mem.mem[12][1] ;
 wire \mem.mem[12][2] ;
 wire \mem.mem[12][3] ;
 wire \mem.mem[12][4] ;
 wire \mem.mem[12][5] ;
 wire \mem.mem[12][6] ;
 wire \mem.mem[12][7] ;
 wire \mem.mem[130][0] ;
 wire \mem.mem[130][1] ;
 wire \mem.mem[130][2] ;
 wire \mem.mem[130][3] ;
 wire \mem.mem[130][4] ;
 wire \mem.mem[130][5] ;
 wire \mem.mem[130][6] ;
 wire \mem.mem[130][7] ;
 wire \mem.mem[131][0] ;
 wire \mem.mem[131][1] ;
 wire \mem.mem[131][2] ;
 wire \mem.mem[131][3] ;
 wire \mem.mem[131][4] ;
 wire \mem.mem[131][5] ;
 wire \mem.mem[131][6] ;
 wire \mem.mem[131][7] ;
 wire \mem.mem[132][0] ;
 wire \mem.mem[132][1] ;
 wire \mem.mem[132][2] ;
 wire \mem.mem[132][3] ;
 wire \mem.mem[132][4] ;
 wire \mem.mem[132][5] ;
 wire \mem.mem[132][6] ;
 wire \mem.mem[132][7] ;
 wire \mem.mem[133][0] ;
 wire \mem.mem[133][1] ;
 wire \mem.mem[133][2] ;
 wire \mem.mem[133][3] ;
 wire \mem.mem[133][4] ;
 wire \mem.mem[133][5] ;
 wire \mem.mem[133][6] ;
 wire \mem.mem[133][7] ;
 wire \mem.mem[134][0] ;
 wire \mem.mem[134][1] ;
 wire \mem.mem[134][2] ;
 wire \mem.mem[134][3] ;
 wire \mem.mem[134][4] ;
 wire \mem.mem[134][5] ;
 wire \mem.mem[134][6] ;
 wire \mem.mem[134][7] ;
 wire \mem.mem[135][0] ;
 wire \mem.mem[135][1] ;
 wire \mem.mem[135][2] ;
 wire \mem.mem[135][3] ;
 wire \mem.mem[135][4] ;
 wire \mem.mem[135][5] ;
 wire \mem.mem[135][6] ;
 wire \mem.mem[135][7] ;
 wire \mem.mem[136][0] ;
 wire \mem.mem[136][1] ;
 wire \mem.mem[136][2] ;
 wire \mem.mem[136][3] ;
 wire \mem.mem[136][4] ;
 wire \mem.mem[136][5] ;
 wire \mem.mem[136][6] ;
 wire \mem.mem[136][7] ;
 wire \mem.mem[137][0] ;
 wire \mem.mem[137][1] ;
 wire \mem.mem[137][2] ;
 wire \mem.mem[137][3] ;
 wire \mem.mem[137][4] ;
 wire \mem.mem[137][5] ;
 wire \mem.mem[137][6] ;
 wire \mem.mem[137][7] ;
 wire \mem.mem[138][0] ;
 wire \mem.mem[138][1] ;
 wire \mem.mem[138][2] ;
 wire \mem.mem[138][3] ;
 wire \mem.mem[138][4] ;
 wire \mem.mem[138][5] ;
 wire \mem.mem[138][6] ;
 wire \mem.mem[138][7] ;
 wire \mem.mem[139][0] ;
 wire \mem.mem[139][1] ;
 wire \mem.mem[139][2] ;
 wire \mem.mem[139][3] ;
 wire \mem.mem[139][4] ;
 wire \mem.mem[139][5] ;
 wire \mem.mem[139][6] ;
 wire \mem.mem[139][7] ;
 wire \mem.mem[13][0] ;
 wire \mem.mem[13][1] ;
 wire \mem.mem[13][2] ;
 wire \mem.mem[13][3] ;
 wire \mem.mem[13][4] ;
 wire \mem.mem[13][5] ;
 wire \mem.mem[13][6] ;
 wire \mem.mem[13][7] ;
 wire \mem.mem[140][0] ;
 wire \mem.mem[140][1] ;
 wire \mem.mem[140][2] ;
 wire \mem.mem[140][3] ;
 wire \mem.mem[140][4] ;
 wire \mem.mem[140][5] ;
 wire \mem.mem[140][6] ;
 wire \mem.mem[140][7] ;
 wire \mem.mem[141][0] ;
 wire \mem.mem[141][1] ;
 wire \mem.mem[141][2] ;
 wire \mem.mem[141][3] ;
 wire \mem.mem[141][4] ;
 wire \mem.mem[141][5] ;
 wire \mem.mem[141][6] ;
 wire \mem.mem[141][7] ;
 wire \mem.mem[142][0] ;
 wire \mem.mem[142][1] ;
 wire \mem.mem[142][2] ;
 wire \mem.mem[142][3] ;
 wire \mem.mem[142][4] ;
 wire \mem.mem[142][5] ;
 wire \mem.mem[142][6] ;
 wire \mem.mem[142][7] ;
 wire \mem.mem[143][0] ;
 wire \mem.mem[143][1] ;
 wire \mem.mem[143][2] ;
 wire \mem.mem[143][3] ;
 wire \mem.mem[143][4] ;
 wire \mem.mem[143][5] ;
 wire \mem.mem[143][6] ;
 wire \mem.mem[143][7] ;
 wire \mem.mem[144][0] ;
 wire \mem.mem[144][1] ;
 wire \mem.mem[144][2] ;
 wire \mem.mem[144][3] ;
 wire \mem.mem[144][4] ;
 wire \mem.mem[144][5] ;
 wire \mem.mem[144][6] ;
 wire \mem.mem[144][7] ;
 wire \mem.mem[145][0] ;
 wire \mem.mem[145][1] ;
 wire \mem.mem[145][2] ;
 wire \mem.mem[145][3] ;
 wire \mem.mem[145][4] ;
 wire \mem.mem[145][5] ;
 wire \mem.mem[145][6] ;
 wire \mem.mem[145][7] ;
 wire \mem.mem[146][0] ;
 wire \mem.mem[146][1] ;
 wire \mem.mem[146][2] ;
 wire \mem.mem[146][3] ;
 wire \mem.mem[146][4] ;
 wire \mem.mem[146][5] ;
 wire \mem.mem[146][6] ;
 wire \mem.mem[146][7] ;
 wire \mem.mem[147][0] ;
 wire \mem.mem[147][1] ;
 wire \mem.mem[147][2] ;
 wire \mem.mem[147][3] ;
 wire \mem.mem[147][4] ;
 wire \mem.mem[147][5] ;
 wire \mem.mem[147][6] ;
 wire \mem.mem[147][7] ;
 wire \mem.mem[148][0] ;
 wire \mem.mem[148][1] ;
 wire \mem.mem[148][2] ;
 wire \mem.mem[148][3] ;
 wire \mem.mem[148][4] ;
 wire \mem.mem[148][5] ;
 wire \mem.mem[148][6] ;
 wire \mem.mem[148][7] ;
 wire \mem.mem[149][0] ;
 wire \mem.mem[149][1] ;
 wire \mem.mem[149][2] ;
 wire \mem.mem[149][3] ;
 wire \mem.mem[149][4] ;
 wire \mem.mem[149][5] ;
 wire \mem.mem[149][6] ;
 wire \mem.mem[149][7] ;
 wire \mem.mem[14][0] ;
 wire \mem.mem[14][1] ;
 wire \mem.mem[14][2] ;
 wire \mem.mem[14][3] ;
 wire \mem.mem[14][4] ;
 wire \mem.mem[14][5] ;
 wire \mem.mem[14][6] ;
 wire \mem.mem[14][7] ;
 wire \mem.mem[150][0] ;
 wire \mem.mem[150][1] ;
 wire \mem.mem[150][2] ;
 wire \mem.mem[150][3] ;
 wire \mem.mem[150][4] ;
 wire \mem.mem[150][5] ;
 wire \mem.mem[150][6] ;
 wire \mem.mem[150][7] ;
 wire \mem.mem[151][0] ;
 wire \mem.mem[151][1] ;
 wire \mem.mem[151][2] ;
 wire \mem.mem[151][3] ;
 wire \mem.mem[151][4] ;
 wire \mem.mem[151][5] ;
 wire \mem.mem[151][6] ;
 wire \mem.mem[151][7] ;
 wire \mem.mem[152][0] ;
 wire \mem.mem[152][1] ;
 wire \mem.mem[152][2] ;
 wire \mem.mem[152][3] ;
 wire \mem.mem[152][4] ;
 wire \mem.mem[152][5] ;
 wire \mem.mem[152][6] ;
 wire \mem.mem[152][7] ;
 wire \mem.mem[153][0] ;
 wire \mem.mem[153][1] ;
 wire \mem.mem[153][2] ;
 wire \mem.mem[153][3] ;
 wire \mem.mem[153][4] ;
 wire \mem.mem[153][5] ;
 wire \mem.mem[153][6] ;
 wire \mem.mem[153][7] ;
 wire \mem.mem[154][0] ;
 wire \mem.mem[154][1] ;
 wire \mem.mem[154][2] ;
 wire \mem.mem[154][3] ;
 wire \mem.mem[154][4] ;
 wire \mem.mem[154][5] ;
 wire \mem.mem[154][6] ;
 wire \mem.mem[154][7] ;
 wire \mem.mem[155][0] ;
 wire \mem.mem[155][1] ;
 wire \mem.mem[155][2] ;
 wire \mem.mem[155][3] ;
 wire \mem.mem[155][4] ;
 wire \mem.mem[155][5] ;
 wire \mem.mem[155][6] ;
 wire \mem.mem[155][7] ;
 wire \mem.mem[156][0] ;
 wire \mem.mem[156][1] ;
 wire \mem.mem[156][2] ;
 wire \mem.mem[156][3] ;
 wire \mem.mem[156][4] ;
 wire \mem.mem[156][5] ;
 wire \mem.mem[156][6] ;
 wire \mem.mem[156][7] ;
 wire \mem.mem[157][0] ;
 wire \mem.mem[157][1] ;
 wire \mem.mem[157][2] ;
 wire \mem.mem[157][3] ;
 wire \mem.mem[157][4] ;
 wire \mem.mem[157][5] ;
 wire \mem.mem[157][6] ;
 wire \mem.mem[157][7] ;
 wire \mem.mem[158][0] ;
 wire \mem.mem[158][1] ;
 wire \mem.mem[158][2] ;
 wire \mem.mem[158][3] ;
 wire \mem.mem[158][4] ;
 wire \mem.mem[158][5] ;
 wire \mem.mem[158][6] ;
 wire \mem.mem[158][7] ;
 wire \mem.mem[159][0] ;
 wire \mem.mem[159][1] ;
 wire \mem.mem[159][2] ;
 wire \mem.mem[159][3] ;
 wire \mem.mem[159][4] ;
 wire \mem.mem[159][5] ;
 wire \mem.mem[159][6] ;
 wire \mem.mem[159][7] ;
 wire \mem.mem[15][0] ;
 wire \mem.mem[15][1] ;
 wire \mem.mem[15][2] ;
 wire \mem.mem[15][3] ;
 wire \mem.mem[15][4] ;
 wire \mem.mem[15][5] ;
 wire \mem.mem[15][6] ;
 wire \mem.mem[15][7] ;
 wire \mem.mem[160][0] ;
 wire \mem.mem[160][1] ;
 wire \mem.mem[160][2] ;
 wire \mem.mem[160][3] ;
 wire \mem.mem[160][4] ;
 wire \mem.mem[160][5] ;
 wire \mem.mem[160][6] ;
 wire \mem.mem[160][7] ;
 wire \mem.mem[161][0] ;
 wire \mem.mem[161][1] ;
 wire \mem.mem[161][2] ;
 wire \mem.mem[161][3] ;
 wire \mem.mem[161][4] ;
 wire \mem.mem[161][5] ;
 wire \mem.mem[161][6] ;
 wire \mem.mem[161][7] ;
 wire \mem.mem[162][0] ;
 wire \mem.mem[162][1] ;
 wire \mem.mem[162][2] ;
 wire \mem.mem[162][3] ;
 wire \mem.mem[162][4] ;
 wire \mem.mem[162][5] ;
 wire \mem.mem[162][6] ;
 wire \mem.mem[162][7] ;
 wire \mem.mem[163][0] ;
 wire \mem.mem[163][1] ;
 wire \mem.mem[163][2] ;
 wire \mem.mem[163][3] ;
 wire \mem.mem[163][4] ;
 wire \mem.mem[163][5] ;
 wire \mem.mem[163][6] ;
 wire \mem.mem[163][7] ;
 wire \mem.mem[164][0] ;
 wire \mem.mem[164][1] ;
 wire \mem.mem[164][2] ;
 wire \mem.mem[164][3] ;
 wire \mem.mem[164][4] ;
 wire \mem.mem[164][5] ;
 wire \mem.mem[164][6] ;
 wire \mem.mem[164][7] ;
 wire \mem.mem[165][0] ;
 wire \mem.mem[165][1] ;
 wire \mem.mem[165][2] ;
 wire \mem.mem[165][3] ;
 wire \mem.mem[165][4] ;
 wire \mem.mem[165][5] ;
 wire \mem.mem[165][6] ;
 wire \mem.mem[165][7] ;
 wire \mem.mem[166][0] ;
 wire \mem.mem[166][1] ;
 wire \mem.mem[166][2] ;
 wire \mem.mem[166][3] ;
 wire \mem.mem[166][4] ;
 wire \mem.mem[166][5] ;
 wire \mem.mem[166][6] ;
 wire \mem.mem[166][7] ;
 wire \mem.mem[167][0] ;
 wire \mem.mem[167][1] ;
 wire \mem.mem[167][2] ;
 wire \mem.mem[167][3] ;
 wire \mem.mem[167][4] ;
 wire \mem.mem[167][5] ;
 wire \mem.mem[167][6] ;
 wire \mem.mem[167][7] ;
 wire \mem.mem[168][0] ;
 wire \mem.mem[168][1] ;
 wire \mem.mem[168][2] ;
 wire \mem.mem[168][3] ;
 wire \mem.mem[168][4] ;
 wire \mem.mem[168][5] ;
 wire \mem.mem[168][6] ;
 wire \mem.mem[168][7] ;
 wire \mem.mem[169][0] ;
 wire \mem.mem[169][1] ;
 wire \mem.mem[169][2] ;
 wire \mem.mem[169][3] ;
 wire \mem.mem[169][4] ;
 wire \mem.mem[169][5] ;
 wire \mem.mem[169][6] ;
 wire \mem.mem[169][7] ;
 wire \mem.mem[16][0] ;
 wire \mem.mem[16][1] ;
 wire \mem.mem[16][2] ;
 wire \mem.mem[16][3] ;
 wire \mem.mem[16][4] ;
 wire \mem.mem[16][5] ;
 wire \mem.mem[16][6] ;
 wire \mem.mem[16][7] ;
 wire \mem.mem[170][0] ;
 wire \mem.mem[170][1] ;
 wire \mem.mem[170][2] ;
 wire \mem.mem[170][3] ;
 wire \mem.mem[170][4] ;
 wire \mem.mem[170][5] ;
 wire \mem.mem[170][6] ;
 wire \mem.mem[170][7] ;
 wire \mem.mem[171][0] ;
 wire \mem.mem[171][1] ;
 wire \mem.mem[171][2] ;
 wire \mem.mem[171][3] ;
 wire \mem.mem[171][4] ;
 wire \mem.mem[171][5] ;
 wire \mem.mem[171][6] ;
 wire \mem.mem[171][7] ;
 wire \mem.mem[172][0] ;
 wire \mem.mem[172][1] ;
 wire \mem.mem[172][2] ;
 wire \mem.mem[172][3] ;
 wire \mem.mem[172][4] ;
 wire \mem.mem[172][5] ;
 wire \mem.mem[172][6] ;
 wire \mem.mem[172][7] ;
 wire \mem.mem[173][0] ;
 wire \mem.mem[173][1] ;
 wire \mem.mem[173][2] ;
 wire \mem.mem[173][3] ;
 wire \mem.mem[173][4] ;
 wire \mem.mem[173][5] ;
 wire \mem.mem[173][6] ;
 wire \mem.mem[173][7] ;
 wire \mem.mem[174][0] ;
 wire \mem.mem[174][1] ;
 wire \mem.mem[174][2] ;
 wire \mem.mem[174][3] ;
 wire \mem.mem[174][4] ;
 wire \mem.mem[174][5] ;
 wire \mem.mem[174][6] ;
 wire \mem.mem[174][7] ;
 wire \mem.mem[175][0] ;
 wire \mem.mem[175][1] ;
 wire \mem.mem[175][2] ;
 wire \mem.mem[175][3] ;
 wire \mem.mem[175][4] ;
 wire \mem.mem[175][5] ;
 wire \mem.mem[175][6] ;
 wire \mem.mem[175][7] ;
 wire \mem.mem[176][0] ;
 wire \mem.mem[176][1] ;
 wire \mem.mem[176][2] ;
 wire \mem.mem[176][3] ;
 wire \mem.mem[176][4] ;
 wire \mem.mem[176][5] ;
 wire \mem.mem[176][6] ;
 wire \mem.mem[176][7] ;
 wire \mem.mem[177][0] ;
 wire \mem.mem[177][1] ;
 wire \mem.mem[177][2] ;
 wire \mem.mem[177][3] ;
 wire \mem.mem[177][4] ;
 wire \mem.mem[177][5] ;
 wire \mem.mem[177][6] ;
 wire \mem.mem[177][7] ;
 wire \mem.mem[178][0] ;
 wire \mem.mem[178][1] ;
 wire \mem.mem[178][2] ;
 wire \mem.mem[178][3] ;
 wire \mem.mem[178][4] ;
 wire \mem.mem[178][5] ;
 wire \mem.mem[178][6] ;
 wire \mem.mem[178][7] ;
 wire \mem.mem[179][0] ;
 wire \mem.mem[179][1] ;
 wire \mem.mem[179][2] ;
 wire \mem.mem[179][3] ;
 wire \mem.mem[179][4] ;
 wire \mem.mem[179][5] ;
 wire \mem.mem[179][6] ;
 wire \mem.mem[179][7] ;
 wire \mem.mem[17][0] ;
 wire \mem.mem[17][1] ;
 wire \mem.mem[17][2] ;
 wire \mem.mem[17][3] ;
 wire \mem.mem[17][4] ;
 wire \mem.mem[17][5] ;
 wire \mem.mem[17][6] ;
 wire \mem.mem[17][7] ;
 wire \mem.mem[180][0] ;
 wire \mem.mem[180][1] ;
 wire \mem.mem[180][2] ;
 wire \mem.mem[180][3] ;
 wire \mem.mem[180][4] ;
 wire \mem.mem[180][5] ;
 wire \mem.mem[180][6] ;
 wire \mem.mem[180][7] ;
 wire \mem.mem[181][0] ;
 wire \mem.mem[181][1] ;
 wire \mem.mem[181][2] ;
 wire \mem.mem[181][3] ;
 wire \mem.mem[181][4] ;
 wire \mem.mem[181][5] ;
 wire \mem.mem[181][6] ;
 wire \mem.mem[181][7] ;
 wire \mem.mem[182][0] ;
 wire \mem.mem[182][1] ;
 wire \mem.mem[182][2] ;
 wire \mem.mem[182][3] ;
 wire \mem.mem[182][4] ;
 wire \mem.mem[182][5] ;
 wire \mem.mem[182][6] ;
 wire \mem.mem[182][7] ;
 wire \mem.mem[183][0] ;
 wire \mem.mem[183][1] ;
 wire \mem.mem[183][2] ;
 wire \mem.mem[183][3] ;
 wire \mem.mem[183][4] ;
 wire \mem.mem[183][5] ;
 wire \mem.mem[183][6] ;
 wire \mem.mem[183][7] ;
 wire \mem.mem[184][0] ;
 wire \mem.mem[184][1] ;
 wire \mem.mem[184][2] ;
 wire \mem.mem[184][3] ;
 wire \mem.mem[184][4] ;
 wire \mem.mem[184][5] ;
 wire \mem.mem[184][6] ;
 wire \mem.mem[184][7] ;
 wire \mem.mem[185][0] ;
 wire \mem.mem[185][1] ;
 wire \mem.mem[185][2] ;
 wire \mem.mem[185][3] ;
 wire \mem.mem[185][4] ;
 wire \mem.mem[185][5] ;
 wire \mem.mem[185][6] ;
 wire \mem.mem[185][7] ;
 wire \mem.mem[186][0] ;
 wire \mem.mem[186][1] ;
 wire \mem.mem[186][2] ;
 wire \mem.mem[186][3] ;
 wire \mem.mem[186][4] ;
 wire \mem.mem[186][5] ;
 wire \mem.mem[186][6] ;
 wire \mem.mem[186][7] ;
 wire \mem.mem[187][0] ;
 wire \mem.mem[187][1] ;
 wire \mem.mem[187][2] ;
 wire \mem.mem[187][3] ;
 wire \mem.mem[187][4] ;
 wire \mem.mem[187][5] ;
 wire \mem.mem[187][6] ;
 wire \mem.mem[187][7] ;
 wire \mem.mem[188][0] ;
 wire \mem.mem[188][1] ;
 wire \mem.mem[188][2] ;
 wire \mem.mem[188][3] ;
 wire \mem.mem[188][4] ;
 wire \mem.mem[188][5] ;
 wire \mem.mem[188][6] ;
 wire \mem.mem[188][7] ;
 wire \mem.mem[189][0] ;
 wire \mem.mem[189][1] ;
 wire \mem.mem[189][2] ;
 wire \mem.mem[189][3] ;
 wire \mem.mem[189][4] ;
 wire \mem.mem[189][5] ;
 wire \mem.mem[189][6] ;
 wire \mem.mem[189][7] ;
 wire \mem.mem[18][0] ;
 wire \mem.mem[18][1] ;
 wire \mem.mem[18][2] ;
 wire \mem.mem[18][3] ;
 wire \mem.mem[18][4] ;
 wire \mem.mem[18][5] ;
 wire \mem.mem[18][6] ;
 wire \mem.mem[18][7] ;
 wire \mem.mem[190][0] ;
 wire \mem.mem[190][1] ;
 wire \mem.mem[190][2] ;
 wire \mem.mem[190][3] ;
 wire \mem.mem[190][4] ;
 wire \mem.mem[190][5] ;
 wire \mem.mem[190][6] ;
 wire \mem.mem[190][7] ;
 wire \mem.mem[191][0] ;
 wire \mem.mem[191][1] ;
 wire \mem.mem[191][2] ;
 wire \mem.mem[191][3] ;
 wire \mem.mem[191][4] ;
 wire \mem.mem[191][5] ;
 wire \mem.mem[191][6] ;
 wire \mem.mem[191][7] ;
 wire \mem.mem[192][0] ;
 wire \mem.mem[192][1] ;
 wire \mem.mem[192][2] ;
 wire \mem.mem[192][3] ;
 wire \mem.mem[192][4] ;
 wire \mem.mem[192][5] ;
 wire \mem.mem[192][6] ;
 wire \mem.mem[192][7] ;
 wire \mem.mem[193][0] ;
 wire \mem.mem[193][1] ;
 wire \mem.mem[193][2] ;
 wire \mem.mem[193][3] ;
 wire \mem.mem[193][4] ;
 wire \mem.mem[193][5] ;
 wire \mem.mem[193][6] ;
 wire \mem.mem[193][7] ;
 wire \mem.mem[194][0] ;
 wire \mem.mem[194][1] ;
 wire \mem.mem[194][2] ;
 wire \mem.mem[194][3] ;
 wire \mem.mem[194][4] ;
 wire \mem.mem[194][5] ;
 wire \mem.mem[194][6] ;
 wire \mem.mem[194][7] ;
 wire \mem.mem[195][0] ;
 wire \mem.mem[195][1] ;
 wire \mem.mem[195][2] ;
 wire \mem.mem[195][3] ;
 wire \mem.mem[195][4] ;
 wire \mem.mem[195][5] ;
 wire \mem.mem[195][6] ;
 wire \mem.mem[195][7] ;
 wire \mem.mem[196][0] ;
 wire \mem.mem[196][1] ;
 wire \mem.mem[196][2] ;
 wire \mem.mem[196][3] ;
 wire \mem.mem[196][4] ;
 wire \mem.mem[196][5] ;
 wire \mem.mem[196][6] ;
 wire \mem.mem[196][7] ;
 wire \mem.mem[197][0] ;
 wire \mem.mem[197][1] ;
 wire \mem.mem[197][2] ;
 wire \mem.mem[197][3] ;
 wire \mem.mem[197][4] ;
 wire \mem.mem[197][5] ;
 wire \mem.mem[197][6] ;
 wire \mem.mem[197][7] ;
 wire \mem.mem[198][0] ;
 wire \mem.mem[198][1] ;
 wire \mem.mem[198][2] ;
 wire \mem.mem[198][3] ;
 wire \mem.mem[198][4] ;
 wire \mem.mem[198][5] ;
 wire \mem.mem[198][6] ;
 wire \mem.mem[198][7] ;
 wire \mem.mem[199][0] ;
 wire \mem.mem[199][1] ;
 wire \mem.mem[199][2] ;
 wire \mem.mem[199][3] ;
 wire \mem.mem[199][4] ;
 wire \mem.mem[199][5] ;
 wire \mem.mem[199][6] ;
 wire \mem.mem[199][7] ;
 wire \mem.mem[19][0] ;
 wire \mem.mem[19][1] ;
 wire \mem.mem[19][2] ;
 wire \mem.mem[19][3] ;
 wire \mem.mem[19][4] ;
 wire \mem.mem[19][5] ;
 wire \mem.mem[19][6] ;
 wire \mem.mem[19][7] ;
 wire \mem.mem[1][0] ;
 wire \mem.mem[1][1] ;
 wire \mem.mem[1][2] ;
 wire \mem.mem[1][3] ;
 wire \mem.mem[1][4] ;
 wire \mem.mem[1][5] ;
 wire \mem.mem[1][6] ;
 wire \mem.mem[1][7] ;
 wire \mem.mem[200][0] ;
 wire \mem.mem[200][1] ;
 wire \mem.mem[200][2] ;
 wire \mem.mem[200][3] ;
 wire \mem.mem[200][4] ;
 wire \mem.mem[200][5] ;
 wire \mem.mem[200][6] ;
 wire \mem.mem[200][7] ;
 wire \mem.mem[201][0] ;
 wire \mem.mem[201][1] ;
 wire \mem.mem[201][2] ;
 wire \mem.mem[201][3] ;
 wire \mem.mem[201][4] ;
 wire \mem.mem[201][5] ;
 wire \mem.mem[201][6] ;
 wire \mem.mem[201][7] ;
 wire \mem.mem[202][0] ;
 wire \mem.mem[202][1] ;
 wire \mem.mem[202][2] ;
 wire \mem.mem[202][3] ;
 wire \mem.mem[202][4] ;
 wire \mem.mem[202][5] ;
 wire \mem.mem[202][6] ;
 wire \mem.mem[202][7] ;
 wire \mem.mem[203][0] ;
 wire \mem.mem[203][1] ;
 wire \mem.mem[203][2] ;
 wire \mem.mem[203][3] ;
 wire \mem.mem[203][4] ;
 wire \mem.mem[203][5] ;
 wire \mem.mem[203][6] ;
 wire \mem.mem[203][7] ;
 wire \mem.mem[204][0] ;
 wire \mem.mem[204][1] ;
 wire \mem.mem[204][2] ;
 wire \mem.mem[204][3] ;
 wire \mem.mem[204][4] ;
 wire \mem.mem[204][5] ;
 wire \mem.mem[204][6] ;
 wire \mem.mem[204][7] ;
 wire \mem.mem[205][0] ;
 wire \mem.mem[205][1] ;
 wire \mem.mem[205][2] ;
 wire \mem.mem[205][3] ;
 wire \mem.mem[205][4] ;
 wire \mem.mem[205][5] ;
 wire \mem.mem[205][6] ;
 wire \mem.mem[205][7] ;
 wire \mem.mem[206][0] ;
 wire \mem.mem[206][1] ;
 wire \mem.mem[206][2] ;
 wire \mem.mem[206][3] ;
 wire \mem.mem[206][4] ;
 wire \mem.mem[206][5] ;
 wire \mem.mem[206][6] ;
 wire \mem.mem[206][7] ;
 wire \mem.mem[207][0] ;
 wire \mem.mem[207][1] ;
 wire \mem.mem[207][2] ;
 wire \mem.mem[207][3] ;
 wire \mem.mem[207][4] ;
 wire \mem.mem[207][5] ;
 wire \mem.mem[207][6] ;
 wire \mem.mem[207][7] ;
 wire \mem.mem[208][0] ;
 wire \mem.mem[208][1] ;
 wire \mem.mem[208][2] ;
 wire \mem.mem[208][3] ;
 wire \mem.mem[208][4] ;
 wire \mem.mem[208][5] ;
 wire \mem.mem[208][6] ;
 wire \mem.mem[208][7] ;
 wire \mem.mem[209][0] ;
 wire \mem.mem[209][1] ;
 wire \mem.mem[209][2] ;
 wire \mem.mem[209][3] ;
 wire \mem.mem[209][4] ;
 wire \mem.mem[209][5] ;
 wire \mem.mem[209][6] ;
 wire \mem.mem[209][7] ;
 wire \mem.mem[20][0] ;
 wire \mem.mem[20][1] ;
 wire \mem.mem[20][2] ;
 wire \mem.mem[20][3] ;
 wire \mem.mem[20][4] ;
 wire \mem.mem[20][5] ;
 wire \mem.mem[20][6] ;
 wire \mem.mem[20][7] ;
 wire \mem.mem[210][0] ;
 wire \mem.mem[210][1] ;
 wire \mem.mem[210][2] ;
 wire \mem.mem[210][3] ;
 wire \mem.mem[210][4] ;
 wire \mem.mem[210][5] ;
 wire \mem.mem[210][6] ;
 wire \mem.mem[210][7] ;
 wire \mem.mem[211][0] ;
 wire \mem.mem[211][1] ;
 wire \mem.mem[211][2] ;
 wire \mem.mem[211][3] ;
 wire \mem.mem[211][4] ;
 wire \mem.mem[211][5] ;
 wire \mem.mem[211][6] ;
 wire \mem.mem[211][7] ;
 wire \mem.mem[212][0] ;
 wire \mem.mem[212][1] ;
 wire \mem.mem[212][2] ;
 wire \mem.mem[212][3] ;
 wire \mem.mem[212][4] ;
 wire \mem.mem[212][5] ;
 wire \mem.mem[212][6] ;
 wire \mem.mem[212][7] ;
 wire \mem.mem[213][0] ;
 wire \mem.mem[213][1] ;
 wire \mem.mem[213][2] ;
 wire \mem.mem[213][3] ;
 wire \mem.mem[213][4] ;
 wire \mem.mem[213][5] ;
 wire \mem.mem[213][6] ;
 wire \mem.mem[213][7] ;
 wire \mem.mem[214][0] ;
 wire \mem.mem[214][1] ;
 wire \mem.mem[214][2] ;
 wire \mem.mem[214][3] ;
 wire \mem.mem[214][4] ;
 wire \mem.mem[214][5] ;
 wire \mem.mem[214][6] ;
 wire \mem.mem[214][7] ;
 wire \mem.mem[215][0] ;
 wire \mem.mem[215][1] ;
 wire \mem.mem[215][2] ;
 wire \mem.mem[215][3] ;
 wire \mem.mem[215][4] ;
 wire \mem.mem[215][5] ;
 wire \mem.mem[215][6] ;
 wire \mem.mem[215][7] ;
 wire \mem.mem[216][0] ;
 wire \mem.mem[216][1] ;
 wire \mem.mem[216][2] ;
 wire \mem.mem[216][3] ;
 wire \mem.mem[216][4] ;
 wire \mem.mem[216][5] ;
 wire \mem.mem[216][6] ;
 wire \mem.mem[216][7] ;
 wire \mem.mem[217][0] ;
 wire \mem.mem[217][1] ;
 wire \mem.mem[217][2] ;
 wire \mem.mem[217][3] ;
 wire \mem.mem[217][4] ;
 wire \mem.mem[217][5] ;
 wire \mem.mem[217][6] ;
 wire \mem.mem[217][7] ;
 wire \mem.mem[218][0] ;
 wire \mem.mem[218][1] ;
 wire \mem.mem[218][2] ;
 wire \mem.mem[218][3] ;
 wire \mem.mem[218][4] ;
 wire \mem.mem[218][5] ;
 wire \mem.mem[218][6] ;
 wire \mem.mem[218][7] ;
 wire \mem.mem[219][0] ;
 wire \mem.mem[219][1] ;
 wire \mem.mem[219][2] ;
 wire \mem.mem[219][3] ;
 wire \mem.mem[219][4] ;
 wire \mem.mem[219][5] ;
 wire \mem.mem[219][6] ;
 wire \mem.mem[219][7] ;
 wire \mem.mem[21][0] ;
 wire \mem.mem[21][1] ;
 wire \mem.mem[21][2] ;
 wire \mem.mem[21][3] ;
 wire \mem.mem[21][4] ;
 wire \mem.mem[21][5] ;
 wire \mem.mem[21][6] ;
 wire \mem.mem[21][7] ;
 wire \mem.mem[220][0] ;
 wire \mem.mem[220][1] ;
 wire \mem.mem[220][2] ;
 wire \mem.mem[220][3] ;
 wire \mem.mem[220][4] ;
 wire \mem.mem[220][5] ;
 wire \mem.mem[220][6] ;
 wire \mem.mem[220][7] ;
 wire \mem.mem[221][0] ;
 wire \mem.mem[221][1] ;
 wire \mem.mem[221][2] ;
 wire \mem.mem[221][3] ;
 wire \mem.mem[221][4] ;
 wire \mem.mem[221][5] ;
 wire \mem.mem[221][6] ;
 wire \mem.mem[221][7] ;
 wire \mem.mem[222][0] ;
 wire \mem.mem[222][1] ;
 wire \mem.mem[222][2] ;
 wire \mem.mem[222][3] ;
 wire \mem.mem[222][4] ;
 wire \mem.mem[222][5] ;
 wire \mem.mem[222][6] ;
 wire \mem.mem[222][7] ;
 wire \mem.mem[223][0] ;
 wire \mem.mem[223][1] ;
 wire \mem.mem[223][2] ;
 wire \mem.mem[223][3] ;
 wire \mem.mem[223][4] ;
 wire \mem.mem[223][5] ;
 wire \mem.mem[223][6] ;
 wire \mem.mem[223][7] ;
 wire \mem.mem[224][0] ;
 wire \mem.mem[224][1] ;
 wire \mem.mem[224][2] ;
 wire \mem.mem[224][3] ;
 wire \mem.mem[224][4] ;
 wire \mem.mem[224][5] ;
 wire \mem.mem[224][6] ;
 wire \mem.mem[224][7] ;
 wire \mem.mem[225][0] ;
 wire \mem.mem[225][1] ;
 wire \mem.mem[225][2] ;
 wire \mem.mem[225][3] ;
 wire \mem.mem[225][4] ;
 wire \mem.mem[225][5] ;
 wire \mem.mem[225][6] ;
 wire \mem.mem[225][7] ;
 wire \mem.mem[226][0] ;
 wire \mem.mem[226][1] ;
 wire \mem.mem[226][2] ;
 wire \mem.mem[226][3] ;
 wire \mem.mem[226][4] ;
 wire \mem.mem[226][5] ;
 wire \mem.mem[226][6] ;
 wire \mem.mem[226][7] ;
 wire \mem.mem[227][0] ;
 wire \mem.mem[227][1] ;
 wire \mem.mem[227][2] ;
 wire \mem.mem[227][3] ;
 wire \mem.mem[227][4] ;
 wire \mem.mem[227][5] ;
 wire \mem.mem[227][6] ;
 wire \mem.mem[227][7] ;
 wire \mem.mem[228][0] ;
 wire \mem.mem[228][1] ;
 wire \mem.mem[228][2] ;
 wire \mem.mem[228][3] ;
 wire \mem.mem[228][4] ;
 wire \mem.mem[228][5] ;
 wire \mem.mem[228][6] ;
 wire \mem.mem[228][7] ;
 wire \mem.mem[229][0] ;
 wire \mem.mem[229][1] ;
 wire \mem.mem[229][2] ;
 wire \mem.mem[229][3] ;
 wire \mem.mem[229][4] ;
 wire \mem.mem[229][5] ;
 wire \mem.mem[229][6] ;
 wire \mem.mem[229][7] ;
 wire \mem.mem[22][0] ;
 wire \mem.mem[22][1] ;
 wire \mem.mem[22][2] ;
 wire \mem.mem[22][3] ;
 wire \mem.mem[22][4] ;
 wire \mem.mem[22][5] ;
 wire \mem.mem[22][6] ;
 wire \mem.mem[22][7] ;
 wire \mem.mem[230][0] ;
 wire \mem.mem[230][1] ;
 wire \mem.mem[230][2] ;
 wire \mem.mem[230][3] ;
 wire \mem.mem[230][4] ;
 wire \mem.mem[230][5] ;
 wire \mem.mem[230][6] ;
 wire \mem.mem[230][7] ;
 wire \mem.mem[231][0] ;
 wire \mem.mem[231][1] ;
 wire \mem.mem[231][2] ;
 wire \mem.mem[231][3] ;
 wire \mem.mem[231][4] ;
 wire \mem.mem[231][5] ;
 wire \mem.mem[231][6] ;
 wire \mem.mem[231][7] ;
 wire \mem.mem[232][0] ;
 wire \mem.mem[232][1] ;
 wire \mem.mem[232][2] ;
 wire \mem.mem[232][3] ;
 wire \mem.mem[232][4] ;
 wire \mem.mem[232][5] ;
 wire \mem.mem[232][6] ;
 wire \mem.mem[232][7] ;
 wire \mem.mem[233][0] ;
 wire \mem.mem[233][1] ;
 wire \mem.mem[233][2] ;
 wire \mem.mem[233][3] ;
 wire \mem.mem[233][4] ;
 wire \mem.mem[233][5] ;
 wire \mem.mem[233][6] ;
 wire \mem.mem[233][7] ;
 wire \mem.mem[234][0] ;
 wire \mem.mem[234][1] ;
 wire \mem.mem[234][2] ;
 wire \mem.mem[234][3] ;
 wire \mem.mem[234][4] ;
 wire \mem.mem[234][5] ;
 wire \mem.mem[234][6] ;
 wire \mem.mem[234][7] ;
 wire \mem.mem[235][0] ;
 wire \mem.mem[235][1] ;
 wire \mem.mem[235][2] ;
 wire \mem.mem[235][3] ;
 wire \mem.mem[235][4] ;
 wire \mem.mem[235][5] ;
 wire \mem.mem[235][6] ;
 wire \mem.mem[235][7] ;
 wire \mem.mem[236][0] ;
 wire \mem.mem[236][1] ;
 wire \mem.mem[236][2] ;
 wire \mem.mem[236][3] ;
 wire \mem.mem[236][4] ;
 wire \mem.mem[236][5] ;
 wire \mem.mem[236][6] ;
 wire \mem.mem[236][7] ;
 wire \mem.mem[237][0] ;
 wire \mem.mem[237][1] ;
 wire \mem.mem[237][2] ;
 wire \mem.mem[237][3] ;
 wire \mem.mem[237][4] ;
 wire \mem.mem[237][5] ;
 wire \mem.mem[237][6] ;
 wire \mem.mem[237][7] ;
 wire \mem.mem[238][0] ;
 wire \mem.mem[238][1] ;
 wire \mem.mem[238][2] ;
 wire \mem.mem[238][3] ;
 wire \mem.mem[238][4] ;
 wire \mem.mem[238][5] ;
 wire \mem.mem[238][6] ;
 wire \mem.mem[238][7] ;
 wire \mem.mem[239][0] ;
 wire \mem.mem[239][1] ;
 wire \mem.mem[239][2] ;
 wire \mem.mem[239][3] ;
 wire \mem.mem[239][4] ;
 wire \mem.mem[239][5] ;
 wire \mem.mem[239][6] ;
 wire \mem.mem[239][7] ;
 wire \mem.mem[23][0] ;
 wire \mem.mem[23][1] ;
 wire \mem.mem[23][2] ;
 wire \mem.mem[23][3] ;
 wire \mem.mem[23][4] ;
 wire \mem.mem[23][5] ;
 wire \mem.mem[23][6] ;
 wire \mem.mem[23][7] ;
 wire \mem.mem[240][0] ;
 wire \mem.mem[240][1] ;
 wire \mem.mem[240][2] ;
 wire \mem.mem[240][3] ;
 wire \mem.mem[240][4] ;
 wire \mem.mem[240][5] ;
 wire \mem.mem[240][6] ;
 wire \mem.mem[240][7] ;
 wire \mem.mem[241][0] ;
 wire \mem.mem[241][1] ;
 wire \mem.mem[241][2] ;
 wire \mem.mem[241][3] ;
 wire \mem.mem[241][4] ;
 wire \mem.mem[241][5] ;
 wire \mem.mem[241][6] ;
 wire \mem.mem[241][7] ;
 wire \mem.mem[242][0] ;
 wire \mem.mem[242][1] ;
 wire \mem.mem[242][2] ;
 wire \mem.mem[242][3] ;
 wire \mem.mem[242][4] ;
 wire \mem.mem[242][5] ;
 wire \mem.mem[242][6] ;
 wire \mem.mem[242][7] ;
 wire \mem.mem[243][0] ;
 wire \mem.mem[243][1] ;
 wire \mem.mem[243][2] ;
 wire \mem.mem[243][3] ;
 wire \mem.mem[243][4] ;
 wire \mem.mem[243][5] ;
 wire \mem.mem[243][6] ;
 wire \mem.mem[243][7] ;
 wire \mem.mem[244][0] ;
 wire \mem.mem[244][1] ;
 wire \mem.mem[244][2] ;
 wire \mem.mem[244][3] ;
 wire \mem.mem[244][4] ;
 wire \mem.mem[244][5] ;
 wire \mem.mem[244][6] ;
 wire \mem.mem[244][7] ;
 wire \mem.mem[245][0] ;
 wire \mem.mem[245][1] ;
 wire \mem.mem[245][2] ;
 wire \mem.mem[245][3] ;
 wire \mem.mem[245][4] ;
 wire \mem.mem[245][5] ;
 wire \mem.mem[245][6] ;
 wire \mem.mem[245][7] ;
 wire \mem.mem[246][0] ;
 wire \mem.mem[246][1] ;
 wire \mem.mem[246][2] ;
 wire \mem.mem[246][3] ;
 wire \mem.mem[246][4] ;
 wire \mem.mem[246][5] ;
 wire \mem.mem[246][6] ;
 wire \mem.mem[246][7] ;
 wire \mem.mem[247][0] ;
 wire \mem.mem[247][1] ;
 wire \mem.mem[247][2] ;
 wire \mem.mem[247][3] ;
 wire \mem.mem[247][4] ;
 wire \mem.mem[247][5] ;
 wire \mem.mem[247][6] ;
 wire \mem.mem[247][7] ;
 wire \mem.mem[248][0] ;
 wire \mem.mem[248][1] ;
 wire \mem.mem[248][2] ;
 wire \mem.mem[248][3] ;
 wire \mem.mem[248][4] ;
 wire \mem.mem[248][5] ;
 wire \mem.mem[248][6] ;
 wire \mem.mem[248][7] ;
 wire \mem.mem[249][0] ;
 wire \mem.mem[249][1] ;
 wire \mem.mem[249][2] ;
 wire \mem.mem[249][3] ;
 wire \mem.mem[249][4] ;
 wire \mem.mem[249][5] ;
 wire \mem.mem[249][6] ;
 wire \mem.mem[249][7] ;
 wire \mem.mem[24][0] ;
 wire \mem.mem[24][1] ;
 wire \mem.mem[24][2] ;
 wire \mem.mem[24][3] ;
 wire \mem.mem[24][4] ;
 wire \mem.mem[24][5] ;
 wire \mem.mem[24][6] ;
 wire \mem.mem[24][7] ;
 wire \mem.mem[250][0] ;
 wire \mem.mem[250][1] ;
 wire \mem.mem[250][2] ;
 wire \mem.mem[250][3] ;
 wire \mem.mem[250][4] ;
 wire \mem.mem[250][5] ;
 wire \mem.mem[250][6] ;
 wire \mem.mem[250][7] ;
 wire \mem.mem[251][0] ;
 wire \mem.mem[251][1] ;
 wire \mem.mem[251][2] ;
 wire \mem.mem[251][3] ;
 wire \mem.mem[251][4] ;
 wire \mem.mem[251][5] ;
 wire \mem.mem[251][6] ;
 wire \mem.mem[251][7] ;
 wire \mem.mem[252][0] ;
 wire \mem.mem[252][1] ;
 wire \mem.mem[252][2] ;
 wire \mem.mem[252][3] ;
 wire \mem.mem[252][4] ;
 wire \mem.mem[252][5] ;
 wire \mem.mem[252][6] ;
 wire \mem.mem[252][7] ;
 wire \mem.mem[25][0] ;
 wire \mem.mem[25][1] ;
 wire \mem.mem[25][2] ;
 wire \mem.mem[25][3] ;
 wire \mem.mem[25][4] ;
 wire \mem.mem[25][5] ;
 wire \mem.mem[25][6] ;
 wire \mem.mem[25][7] ;
 wire \mem.mem[26][0] ;
 wire \mem.mem[26][1] ;
 wire \mem.mem[26][2] ;
 wire \mem.mem[26][3] ;
 wire \mem.mem[26][4] ;
 wire \mem.mem[26][5] ;
 wire \mem.mem[26][6] ;
 wire \mem.mem[26][7] ;
 wire \mem.mem[27][0] ;
 wire \mem.mem[27][1] ;
 wire \mem.mem[27][2] ;
 wire \mem.mem[27][3] ;
 wire \mem.mem[27][4] ;
 wire \mem.mem[27][5] ;
 wire \mem.mem[27][6] ;
 wire \mem.mem[27][7] ;
 wire \mem.mem[28][0] ;
 wire \mem.mem[28][1] ;
 wire \mem.mem[28][2] ;
 wire \mem.mem[28][3] ;
 wire \mem.mem[28][4] ;
 wire \mem.mem[28][5] ;
 wire \mem.mem[28][6] ;
 wire \mem.mem[28][7] ;
 wire \mem.mem[29][0] ;
 wire \mem.mem[29][1] ;
 wire \mem.mem[29][2] ;
 wire \mem.mem[29][3] ;
 wire \mem.mem[29][4] ;
 wire \mem.mem[29][5] ;
 wire \mem.mem[29][6] ;
 wire \mem.mem[29][7] ;
 wire \mem.mem[2][0] ;
 wire \mem.mem[2][1] ;
 wire \mem.mem[2][2] ;
 wire \mem.mem[2][3] ;
 wire \mem.mem[2][4] ;
 wire \mem.mem[2][5] ;
 wire \mem.mem[2][6] ;
 wire \mem.mem[2][7] ;
 wire \mem.mem[30][0] ;
 wire \mem.mem[30][1] ;
 wire \mem.mem[30][2] ;
 wire \mem.mem[30][3] ;
 wire \mem.mem[30][4] ;
 wire \mem.mem[30][5] ;
 wire \mem.mem[30][6] ;
 wire \mem.mem[30][7] ;
 wire \mem.mem[31][0] ;
 wire \mem.mem[31][1] ;
 wire \mem.mem[31][2] ;
 wire \mem.mem[31][3] ;
 wire \mem.mem[31][4] ;
 wire \mem.mem[31][5] ;
 wire \mem.mem[31][6] ;
 wire \mem.mem[31][7] ;
 wire \mem.mem[32][0] ;
 wire \mem.mem[32][1] ;
 wire \mem.mem[32][2] ;
 wire \mem.mem[32][3] ;
 wire \mem.mem[32][4] ;
 wire \mem.mem[32][5] ;
 wire \mem.mem[32][6] ;
 wire \mem.mem[32][7] ;
 wire \mem.mem[33][0] ;
 wire \mem.mem[33][1] ;
 wire \mem.mem[33][2] ;
 wire \mem.mem[33][3] ;
 wire \mem.mem[33][4] ;
 wire \mem.mem[33][5] ;
 wire \mem.mem[33][6] ;
 wire \mem.mem[33][7] ;
 wire \mem.mem[34][0] ;
 wire \mem.mem[34][1] ;
 wire \mem.mem[34][2] ;
 wire \mem.mem[34][3] ;
 wire \mem.mem[34][4] ;
 wire \mem.mem[34][5] ;
 wire \mem.mem[34][6] ;
 wire \mem.mem[34][7] ;
 wire \mem.mem[35][0] ;
 wire \mem.mem[35][1] ;
 wire \mem.mem[35][2] ;
 wire \mem.mem[35][3] ;
 wire \mem.mem[35][4] ;
 wire \mem.mem[35][5] ;
 wire \mem.mem[35][6] ;
 wire \mem.mem[35][7] ;
 wire \mem.mem[36][0] ;
 wire \mem.mem[36][1] ;
 wire \mem.mem[36][2] ;
 wire \mem.mem[36][3] ;
 wire \mem.mem[36][4] ;
 wire \mem.mem[36][5] ;
 wire \mem.mem[36][6] ;
 wire \mem.mem[36][7] ;
 wire \mem.mem[37][0] ;
 wire \mem.mem[37][1] ;
 wire \mem.mem[37][2] ;
 wire \mem.mem[37][3] ;
 wire \mem.mem[37][4] ;
 wire \mem.mem[37][5] ;
 wire \mem.mem[37][6] ;
 wire \mem.mem[37][7] ;
 wire \mem.mem[38][0] ;
 wire \mem.mem[38][1] ;
 wire \mem.mem[38][2] ;
 wire \mem.mem[38][3] ;
 wire \mem.mem[38][4] ;
 wire \mem.mem[38][5] ;
 wire \mem.mem[38][6] ;
 wire \mem.mem[38][7] ;
 wire \mem.mem[39][0] ;
 wire \mem.mem[39][1] ;
 wire \mem.mem[39][2] ;
 wire \mem.mem[39][3] ;
 wire \mem.mem[39][4] ;
 wire \mem.mem[39][5] ;
 wire \mem.mem[39][6] ;
 wire \mem.mem[39][7] ;
 wire \mem.mem[3][0] ;
 wire \mem.mem[3][1] ;
 wire \mem.mem[3][2] ;
 wire \mem.mem[3][3] ;
 wire \mem.mem[3][4] ;
 wire \mem.mem[3][5] ;
 wire \mem.mem[3][6] ;
 wire \mem.mem[3][7] ;
 wire \mem.mem[40][0] ;
 wire \mem.mem[40][1] ;
 wire \mem.mem[40][2] ;
 wire \mem.mem[40][3] ;
 wire \mem.mem[40][4] ;
 wire \mem.mem[40][5] ;
 wire \mem.mem[40][6] ;
 wire \mem.mem[40][7] ;
 wire \mem.mem[41][0] ;
 wire \mem.mem[41][1] ;
 wire \mem.mem[41][2] ;
 wire \mem.mem[41][3] ;
 wire \mem.mem[41][4] ;
 wire \mem.mem[41][5] ;
 wire \mem.mem[41][6] ;
 wire \mem.mem[41][7] ;
 wire \mem.mem[42][0] ;
 wire \mem.mem[42][1] ;
 wire \mem.mem[42][2] ;
 wire \mem.mem[42][3] ;
 wire \mem.mem[42][4] ;
 wire \mem.mem[42][5] ;
 wire \mem.mem[42][6] ;
 wire \mem.mem[42][7] ;
 wire \mem.mem[43][0] ;
 wire \mem.mem[43][1] ;
 wire \mem.mem[43][2] ;
 wire \mem.mem[43][3] ;
 wire \mem.mem[43][4] ;
 wire \mem.mem[43][5] ;
 wire \mem.mem[43][6] ;
 wire \mem.mem[43][7] ;
 wire \mem.mem[44][0] ;
 wire \mem.mem[44][1] ;
 wire \mem.mem[44][2] ;
 wire \mem.mem[44][3] ;
 wire \mem.mem[44][4] ;
 wire \mem.mem[44][5] ;
 wire \mem.mem[44][6] ;
 wire \mem.mem[44][7] ;
 wire \mem.mem[45][0] ;
 wire \mem.mem[45][1] ;
 wire \mem.mem[45][2] ;
 wire \mem.mem[45][3] ;
 wire \mem.mem[45][4] ;
 wire \mem.mem[45][5] ;
 wire \mem.mem[45][6] ;
 wire \mem.mem[45][7] ;
 wire \mem.mem[46][0] ;
 wire \mem.mem[46][1] ;
 wire \mem.mem[46][2] ;
 wire \mem.mem[46][3] ;
 wire \mem.mem[46][4] ;
 wire \mem.mem[46][5] ;
 wire \mem.mem[46][6] ;
 wire \mem.mem[46][7] ;
 wire \mem.mem[47][0] ;
 wire \mem.mem[47][1] ;
 wire \mem.mem[47][2] ;
 wire \mem.mem[47][3] ;
 wire \mem.mem[47][4] ;
 wire \mem.mem[47][5] ;
 wire \mem.mem[47][6] ;
 wire \mem.mem[47][7] ;
 wire \mem.mem[48][0] ;
 wire \mem.mem[48][1] ;
 wire \mem.mem[48][2] ;
 wire \mem.mem[48][3] ;
 wire \mem.mem[48][4] ;
 wire \mem.mem[48][5] ;
 wire \mem.mem[48][6] ;
 wire \mem.mem[48][7] ;
 wire \mem.mem[49][0] ;
 wire \mem.mem[49][1] ;
 wire \mem.mem[49][2] ;
 wire \mem.mem[49][3] ;
 wire \mem.mem[49][4] ;
 wire \mem.mem[49][5] ;
 wire \mem.mem[49][6] ;
 wire \mem.mem[49][7] ;
 wire \mem.mem[4][0] ;
 wire \mem.mem[4][1] ;
 wire \mem.mem[4][2] ;
 wire \mem.mem[4][3] ;
 wire \mem.mem[4][4] ;
 wire \mem.mem[4][5] ;
 wire \mem.mem[4][6] ;
 wire \mem.mem[4][7] ;
 wire \mem.mem[50][0] ;
 wire \mem.mem[50][1] ;
 wire \mem.mem[50][2] ;
 wire \mem.mem[50][3] ;
 wire \mem.mem[50][4] ;
 wire \mem.mem[50][5] ;
 wire \mem.mem[50][6] ;
 wire \mem.mem[50][7] ;
 wire \mem.mem[51][0] ;
 wire \mem.mem[51][1] ;
 wire \mem.mem[51][2] ;
 wire \mem.mem[51][3] ;
 wire \mem.mem[51][4] ;
 wire \mem.mem[51][5] ;
 wire \mem.mem[51][6] ;
 wire \mem.mem[51][7] ;
 wire \mem.mem[52][0] ;
 wire \mem.mem[52][1] ;
 wire \mem.mem[52][2] ;
 wire \mem.mem[52][3] ;
 wire \mem.mem[52][4] ;
 wire \mem.mem[52][5] ;
 wire \mem.mem[52][6] ;
 wire \mem.mem[52][7] ;
 wire \mem.mem[53][0] ;
 wire \mem.mem[53][1] ;
 wire \mem.mem[53][2] ;
 wire \mem.mem[53][3] ;
 wire \mem.mem[53][4] ;
 wire \mem.mem[53][5] ;
 wire \mem.mem[53][6] ;
 wire \mem.mem[53][7] ;
 wire \mem.mem[54][0] ;
 wire \mem.mem[54][1] ;
 wire \mem.mem[54][2] ;
 wire \mem.mem[54][3] ;
 wire \mem.mem[54][4] ;
 wire \mem.mem[54][5] ;
 wire \mem.mem[54][6] ;
 wire \mem.mem[54][7] ;
 wire \mem.mem[55][0] ;
 wire \mem.mem[55][1] ;
 wire \mem.mem[55][2] ;
 wire \mem.mem[55][3] ;
 wire \mem.mem[55][4] ;
 wire \mem.mem[55][5] ;
 wire \mem.mem[55][6] ;
 wire \mem.mem[55][7] ;
 wire \mem.mem[56][0] ;
 wire \mem.mem[56][1] ;
 wire \mem.mem[56][2] ;
 wire \mem.mem[56][3] ;
 wire \mem.mem[56][4] ;
 wire \mem.mem[56][5] ;
 wire \mem.mem[56][6] ;
 wire \mem.mem[56][7] ;
 wire \mem.mem[57][0] ;
 wire \mem.mem[57][1] ;
 wire \mem.mem[57][2] ;
 wire \mem.mem[57][3] ;
 wire \mem.mem[57][4] ;
 wire \mem.mem[57][5] ;
 wire \mem.mem[57][6] ;
 wire \mem.mem[57][7] ;
 wire \mem.mem[58][0] ;
 wire \mem.mem[58][1] ;
 wire \mem.mem[58][2] ;
 wire \mem.mem[58][3] ;
 wire \mem.mem[58][4] ;
 wire \mem.mem[58][5] ;
 wire \mem.mem[58][6] ;
 wire \mem.mem[58][7] ;
 wire \mem.mem[59][0] ;
 wire \mem.mem[59][1] ;
 wire \mem.mem[59][2] ;
 wire \mem.mem[59][3] ;
 wire \mem.mem[59][4] ;
 wire \mem.mem[59][5] ;
 wire \mem.mem[59][6] ;
 wire \mem.mem[59][7] ;
 wire \mem.mem[5][0] ;
 wire \mem.mem[5][1] ;
 wire \mem.mem[5][2] ;
 wire \mem.mem[5][3] ;
 wire \mem.mem[5][4] ;
 wire \mem.mem[5][5] ;
 wire \mem.mem[5][6] ;
 wire \mem.mem[5][7] ;
 wire \mem.mem[60][0] ;
 wire \mem.mem[60][1] ;
 wire \mem.mem[60][2] ;
 wire \mem.mem[60][3] ;
 wire \mem.mem[60][4] ;
 wire \mem.mem[60][5] ;
 wire \mem.mem[60][6] ;
 wire \mem.mem[60][7] ;
 wire \mem.mem[61][0] ;
 wire \mem.mem[61][1] ;
 wire \mem.mem[61][2] ;
 wire \mem.mem[61][3] ;
 wire \mem.mem[61][4] ;
 wire \mem.mem[61][5] ;
 wire \mem.mem[61][6] ;
 wire \mem.mem[61][7] ;
 wire \mem.mem[62][0] ;
 wire \mem.mem[62][1] ;
 wire \mem.mem[62][2] ;
 wire \mem.mem[62][3] ;
 wire \mem.mem[62][4] ;
 wire \mem.mem[62][5] ;
 wire \mem.mem[62][6] ;
 wire \mem.mem[62][7] ;
 wire \mem.mem[63][0] ;
 wire \mem.mem[63][1] ;
 wire \mem.mem[63][2] ;
 wire \mem.mem[63][3] ;
 wire \mem.mem[63][4] ;
 wire \mem.mem[63][5] ;
 wire \mem.mem[63][6] ;
 wire \mem.mem[63][7] ;
 wire \mem.mem[64][0] ;
 wire \mem.mem[64][1] ;
 wire \mem.mem[64][2] ;
 wire \mem.mem[64][3] ;
 wire \mem.mem[64][4] ;
 wire \mem.mem[64][5] ;
 wire \mem.mem[64][6] ;
 wire \mem.mem[64][7] ;
 wire \mem.mem[65][0] ;
 wire \mem.mem[65][1] ;
 wire \mem.mem[65][2] ;
 wire \mem.mem[65][3] ;
 wire \mem.mem[65][4] ;
 wire \mem.mem[65][5] ;
 wire \mem.mem[65][6] ;
 wire \mem.mem[65][7] ;
 wire \mem.mem[66][0] ;
 wire \mem.mem[66][1] ;
 wire \mem.mem[66][2] ;
 wire \mem.mem[66][3] ;
 wire \mem.mem[66][4] ;
 wire \mem.mem[66][5] ;
 wire \mem.mem[66][6] ;
 wire \mem.mem[66][7] ;
 wire \mem.mem[67][0] ;
 wire \mem.mem[67][1] ;
 wire \mem.mem[67][2] ;
 wire \mem.mem[67][3] ;
 wire \mem.mem[67][4] ;
 wire \mem.mem[67][5] ;
 wire \mem.mem[67][6] ;
 wire \mem.mem[67][7] ;
 wire \mem.mem[68][0] ;
 wire \mem.mem[68][1] ;
 wire \mem.mem[68][2] ;
 wire \mem.mem[68][3] ;
 wire \mem.mem[68][4] ;
 wire \mem.mem[68][5] ;
 wire \mem.mem[68][6] ;
 wire \mem.mem[68][7] ;
 wire \mem.mem[69][0] ;
 wire \mem.mem[69][1] ;
 wire \mem.mem[69][2] ;
 wire \mem.mem[69][3] ;
 wire \mem.mem[69][4] ;
 wire \mem.mem[69][5] ;
 wire \mem.mem[69][6] ;
 wire \mem.mem[69][7] ;
 wire \mem.mem[6][0] ;
 wire \mem.mem[6][1] ;
 wire \mem.mem[6][2] ;
 wire \mem.mem[6][3] ;
 wire \mem.mem[6][4] ;
 wire \mem.mem[6][5] ;
 wire \mem.mem[6][6] ;
 wire \mem.mem[6][7] ;
 wire \mem.mem[70][0] ;
 wire \mem.mem[70][1] ;
 wire \mem.mem[70][2] ;
 wire \mem.mem[70][3] ;
 wire \mem.mem[70][4] ;
 wire \mem.mem[70][5] ;
 wire \mem.mem[70][6] ;
 wire \mem.mem[70][7] ;
 wire \mem.mem[71][0] ;
 wire \mem.mem[71][1] ;
 wire \mem.mem[71][2] ;
 wire \mem.mem[71][3] ;
 wire \mem.mem[71][4] ;
 wire \mem.mem[71][5] ;
 wire \mem.mem[71][6] ;
 wire \mem.mem[71][7] ;
 wire \mem.mem[72][0] ;
 wire \mem.mem[72][1] ;
 wire \mem.mem[72][2] ;
 wire \mem.mem[72][3] ;
 wire \mem.mem[72][4] ;
 wire \mem.mem[72][5] ;
 wire \mem.mem[72][6] ;
 wire \mem.mem[72][7] ;
 wire \mem.mem[73][0] ;
 wire \mem.mem[73][1] ;
 wire \mem.mem[73][2] ;
 wire \mem.mem[73][3] ;
 wire \mem.mem[73][4] ;
 wire \mem.mem[73][5] ;
 wire \mem.mem[73][6] ;
 wire \mem.mem[73][7] ;
 wire \mem.mem[74][0] ;
 wire \mem.mem[74][1] ;
 wire \mem.mem[74][2] ;
 wire \mem.mem[74][3] ;
 wire \mem.mem[74][4] ;
 wire \mem.mem[74][5] ;
 wire \mem.mem[74][6] ;
 wire \mem.mem[74][7] ;
 wire \mem.mem[75][0] ;
 wire \mem.mem[75][1] ;
 wire \mem.mem[75][2] ;
 wire \mem.mem[75][3] ;
 wire \mem.mem[75][4] ;
 wire \mem.mem[75][5] ;
 wire \mem.mem[75][6] ;
 wire \mem.mem[75][7] ;
 wire \mem.mem[76][0] ;
 wire \mem.mem[76][1] ;
 wire \mem.mem[76][2] ;
 wire \mem.mem[76][3] ;
 wire \mem.mem[76][4] ;
 wire \mem.mem[76][5] ;
 wire \mem.mem[76][6] ;
 wire \mem.mem[76][7] ;
 wire \mem.mem[77][0] ;
 wire \mem.mem[77][1] ;
 wire \mem.mem[77][2] ;
 wire \mem.mem[77][3] ;
 wire \mem.mem[77][4] ;
 wire \mem.mem[77][5] ;
 wire \mem.mem[77][6] ;
 wire \mem.mem[77][7] ;
 wire \mem.mem[78][0] ;
 wire \mem.mem[78][1] ;
 wire \mem.mem[78][2] ;
 wire \mem.mem[78][3] ;
 wire \mem.mem[78][4] ;
 wire \mem.mem[78][5] ;
 wire \mem.mem[78][6] ;
 wire \mem.mem[78][7] ;
 wire \mem.mem[79][0] ;
 wire \mem.mem[79][1] ;
 wire \mem.mem[79][2] ;
 wire \mem.mem[79][3] ;
 wire \mem.mem[79][4] ;
 wire \mem.mem[79][5] ;
 wire \mem.mem[79][6] ;
 wire \mem.mem[79][7] ;
 wire \mem.mem[7][0] ;
 wire \mem.mem[7][1] ;
 wire \mem.mem[7][2] ;
 wire \mem.mem[7][3] ;
 wire \mem.mem[7][4] ;
 wire \mem.mem[7][5] ;
 wire \mem.mem[7][6] ;
 wire \mem.mem[7][7] ;
 wire \mem.mem[80][0] ;
 wire \mem.mem[80][1] ;
 wire \mem.mem[80][2] ;
 wire \mem.mem[80][3] ;
 wire \mem.mem[80][4] ;
 wire \mem.mem[80][5] ;
 wire \mem.mem[80][6] ;
 wire \mem.mem[80][7] ;
 wire \mem.mem[81][0] ;
 wire \mem.mem[81][1] ;
 wire \mem.mem[81][2] ;
 wire \mem.mem[81][3] ;
 wire \mem.mem[81][4] ;
 wire \mem.mem[81][5] ;
 wire \mem.mem[81][6] ;
 wire \mem.mem[81][7] ;
 wire \mem.mem[82][0] ;
 wire \mem.mem[82][1] ;
 wire \mem.mem[82][2] ;
 wire \mem.mem[82][3] ;
 wire \mem.mem[82][4] ;
 wire \mem.mem[82][5] ;
 wire \mem.mem[82][6] ;
 wire \mem.mem[82][7] ;
 wire \mem.mem[83][0] ;
 wire \mem.mem[83][1] ;
 wire \mem.mem[83][2] ;
 wire \mem.mem[83][3] ;
 wire \mem.mem[83][4] ;
 wire \mem.mem[83][5] ;
 wire \mem.mem[83][6] ;
 wire \mem.mem[83][7] ;
 wire \mem.mem[84][0] ;
 wire \mem.mem[84][1] ;
 wire \mem.mem[84][2] ;
 wire \mem.mem[84][3] ;
 wire \mem.mem[84][4] ;
 wire \mem.mem[84][5] ;
 wire \mem.mem[84][6] ;
 wire \mem.mem[84][7] ;
 wire \mem.mem[85][0] ;
 wire \mem.mem[85][1] ;
 wire \mem.mem[85][2] ;
 wire \mem.mem[85][3] ;
 wire \mem.mem[85][4] ;
 wire \mem.mem[85][5] ;
 wire \mem.mem[85][6] ;
 wire \mem.mem[85][7] ;
 wire \mem.mem[86][0] ;
 wire \mem.mem[86][1] ;
 wire \mem.mem[86][2] ;
 wire \mem.mem[86][3] ;
 wire \mem.mem[86][4] ;
 wire \mem.mem[86][5] ;
 wire \mem.mem[86][6] ;
 wire \mem.mem[86][7] ;
 wire \mem.mem[87][0] ;
 wire \mem.mem[87][1] ;
 wire \mem.mem[87][2] ;
 wire \mem.mem[87][3] ;
 wire \mem.mem[87][4] ;
 wire \mem.mem[87][5] ;
 wire \mem.mem[87][6] ;
 wire \mem.mem[87][7] ;
 wire \mem.mem[88][0] ;
 wire \mem.mem[88][1] ;
 wire \mem.mem[88][2] ;
 wire \mem.mem[88][3] ;
 wire \mem.mem[88][4] ;
 wire \mem.mem[88][5] ;
 wire \mem.mem[88][6] ;
 wire \mem.mem[88][7] ;
 wire \mem.mem[89][0] ;
 wire \mem.mem[89][1] ;
 wire \mem.mem[89][2] ;
 wire \mem.mem[89][3] ;
 wire \mem.mem[89][4] ;
 wire \mem.mem[89][5] ;
 wire \mem.mem[89][6] ;
 wire \mem.mem[89][7] ;
 wire \mem.mem[8][0] ;
 wire \mem.mem[8][1] ;
 wire \mem.mem[8][2] ;
 wire \mem.mem[8][3] ;
 wire \mem.mem[8][4] ;
 wire \mem.mem[8][5] ;
 wire \mem.mem[8][6] ;
 wire \mem.mem[8][7] ;
 wire \mem.mem[90][0] ;
 wire \mem.mem[90][1] ;
 wire \mem.mem[90][2] ;
 wire \mem.mem[90][3] ;
 wire \mem.mem[90][4] ;
 wire \mem.mem[90][5] ;
 wire \mem.mem[90][6] ;
 wire \mem.mem[90][7] ;
 wire \mem.mem[91][0] ;
 wire \mem.mem[91][1] ;
 wire \mem.mem[91][2] ;
 wire \mem.mem[91][3] ;
 wire \mem.mem[91][4] ;
 wire \mem.mem[91][5] ;
 wire \mem.mem[91][6] ;
 wire \mem.mem[91][7] ;
 wire \mem.mem[92][0] ;
 wire \mem.mem[92][1] ;
 wire \mem.mem[92][2] ;
 wire \mem.mem[92][3] ;
 wire \mem.mem[92][4] ;
 wire \mem.mem[92][5] ;
 wire \mem.mem[92][6] ;
 wire \mem.mem[92][7] ;
 wire \mem.mem[93][0] ;
 wire \mem.mem[93][1] ;
 wire \mem.mem[93][2] ;
 wire \mem.mem[93][3] ;
 wire \mem.mem[93][4] ;
 wire \mem.mem[93][5] ;
 wire \mem.mem[93][6] ;
 wire \mem.mem[93][7] ;
 wire \mem.mem[94][0] ;
 wire \mem.mem[94][1] ;
 wire \mem.mem[94][2] ;
 wire \mem.mem[94][3] ;
 wire \mem.mem[94][4] ;
 wire \mem.mem[94][5] ;
 wire \mem.mem[94][6] ;
 wire \mem.mem[94][7] ;
 wire \mem.mem[95][0] ;
 wire \mem.mem[95][1] ;
 wire \mem.mem[95][2] ;
 wire \mem.mem[95][3] ;
 wire \mem.mem[95][4] ;
 wire \mem.mem[95][5] ;
 wire \mem.mem[95][6] ;
 wire \mem.mem[95][7] ;
 wire \mem.mem[96][0] ;
 wire \mem.mem[96][1] ;
 wire \mem.mem[96][2] ;
 wire \mem.mem[96][3] ;
 wire \mem.mem[96][4] ;
 wire \mem.mem[96][5] ;
 wire \mem.mem[96][6] ;
 wire \mem.mem[96][7] ;
 wire \mem.mem[97][0] ;
 wire \mem.mem[97][1] ;
 wire \mem.mem[97][2] ;
 wire \mem.mem[97][3] ;
 wire \mem.mem[97][4] ;
 wire \mem.mem[97][5] ;
 wire \mem.mem[97][6] ;
 wire \mem.mem[97][7] ;
 wire \mem.mem[98][0] ;
 wire \mem.mem[98][1] ;
 wire \mem.mem[98][2] ;
 wire \mem.mem[98][3] ;
 wire \mem.mem[98][4] ;
 wire \mem.mem[98][5] ;
 wire \mem.mem[98][6] ;
 wire \mem.mem[98][7] ;
 wire \mem.mem[99][0] ;
 wire \mem.mem[99][1] ;
 wire \mem.mem[99][2] ;
 wire \mem.mem[99][3] ;
 wire \mem.mem[99][4] ;
 wire \mem.mem[99][5] ;
 wire \mem.mem[99][6] ;
 wire \mem.mem[99][7] ;
 wire \mem.mem[9][0] ;
 wire \mem.mem[9][1] ;
 wire \mem.mem[9][2] ;
 wire \mem.mem[9][3] ;
 wire \mem.mem[9][4] ;
 wire \mem.mem[9][5] ;
 wire \mem.mem[9][6] ;
 wire \mem.mem[9][7] ;
 wire \mem.out_strobe ;
 wire \mem.uo_out[0] ;
 wire \mem.uo_out[1] ;
 wire \mem.uo_out[2] ;
 wire \mem.uo_out[3] ;
 wire \mem.uo_out[4] ;
 wire \mem.uo_out[5] ;
 wire \mem.uo_out[6] ;
 wire \mem.uo_out[7] ;
 wire \mem.wr_en ;
 wire \mem_A[0] ;
 wire \mem_A[1] ;
 wire \mem_A[2] ;
 wire \mem_A[3] ;
 wire \mem_A[4] ;
 wire \mem_A[5] ;
 wire \mem_A[6] ;
 wire \mem_A[7] ;
 wire prev_run;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net15;
 wire net2129;
 wire net16;
 wire net17;
 wire clknet_leaf_0_clk;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;

 sg13g2_inv_1 _09387_ (.Y(_02120_),
    .A(net2631));
 sg13g2_inv_1 _09388_ (.Y(_02121_),
    .A(net2177));
 sg13g2_inv_1 _09389_ (.Y(_02122_),
    .A(net2167));
 sg13g2_inv_1 _09390_ (.Y(_02123_),
    .A(net2361));
 sg13g2_inv_1 _09391_ (.Y(_02124_),
    .A(net4581));
 sg13g2_inv_1 _09392_ (.Y(_02125_),
    .A(net2148));
 sg13g2_inv_1 _09393_ (.Y(_02126_),
    .A(net5040));
 sg13g2_inv_1 _09394_ (.Y(_02127_),
    .A(net2203));
 sg13g2_inv_1 _09395_ (.Y(_02128_),
    .A(net5098));
 sg13g2_inv_1 _09396_ (.Y(_02129_),
    .A(net5201));
 sg13g2_inv_2 _09397_ (.Y(_02130_),
    .A(net4850));
 sg13g2_inv_1 _09398_ (.Y(_02131_),
    .A(\PC[7] ));
 sg13g2_inv_1 _09399_ (.Y(_02132_),
    .A(\PC[3] ));
 sg13g2_inv_1 _09400_ (.Y(_02133_),
    .A(\PC[2] ));
 sg13g2_inv_1 _09401_ (.Y(_02134_),
    .A(\PC[1] ));
 sg13g2_inv_1 _09402_ (.Y(_02135_),
    .A(\PC[0] ));
 sg13g2_inv_1 _09403_ (.Y(_02136_),
    .A(\state[2] ));
 sg13g2_inv_1 _09404_ (.Y(_02137_),
    .A(net2133));
 sg13g2_inv_1 _09405_ (.Y(_02138_),
    .A(net2616));
 sg13g2_inv_1 _09406_ (.Y(_02139_),
    .A(net2141));
 sg13g2_inv_1 _09407_ (.Y(_02140_),
    .A(net2655));
 sg13g2_inv_1 _09408_ (.Y(_02141_),
    .A(net2782));
 sg13g2_inv_1 _09409_ (.Y(_02142_),
    .A(net2673));
 sg13g2_inv_2 _09410_ (.Y(_02143_),
    .A(net3742));
 sg13g2_inv_2 _09411_ (.Y(_02144_),
    .A(net3686));
 sg13g2_inv_1 _09412_ (.Y(_02145_),
    .A(net3648));
 sg13g2_inv_4 _09413_ (.A(net3626),
    .Y(_02146_));
 sg13g2_inv_8 _09414_ (.Y(_02147_),
    .A(net3619));
 sg13g2_inv_4 _09415_ (.A(net3614),
    .Y(_02148_));
 sg13g2_inv_2 _09416_ (.Y(_02149_),
    .A(_00007_));
 sg13g2_inv_1 _09417_ (.Y(_02150_),
    .A(net2));
 sg13g2_inv_1 _09418_ (.Y(_02151_),
    .A(net2222));
 sg13g2_inv_1 _09419_ (.Y(_02152_),
    .A(\mem.mem[14][2] ));
 sg13g2_inv_1 _09420_ (.Y(_02153_),
    .A(net2164));
 sg13g2_inv_1 _09421_ (.Y(_02154_),
    .A(\mem.mem[102][2] ));
 sg13g2_inv_1 _09422_ (.Y(_02155_),
    .A(\mem.mem[132][2] ));
 sg13g2_inv_1 _09423_ (.Y(_02156_),
    .A(net4));
 sg13g2_inv_1 _09424_ (.Y(_02157_),
    .A(\mem.mem[190][3] ));
 sg13g2_inv_2 _09425_ (.Y(_02158_),
    .A(net5));
 sg13g2_inv_1 _09426_ (.Y(_02159_),
    .A(\mem.mem[126][4] ));
 sg13g2_inv_2 _09427_ (.Y(_02160_),
    .A(net6));
 sg13g2_inv_1 _09428_ (.Y(_02161_),
    .A(net2171));
 sg13g2_inv_1 _09429_ (.Y(_02162_),
    .A(net2221));
 sg13g2_inv_1 _09430_ (.Y(_02163_),
    .A(\mem.mem[190][5] ));
 sg13g2_inv_1 _09431_ (.Y(_02164_),
    .A(net2183));
 sg13g2_inv_1 _09432_ (.Y(_02165_),
    .A(net2166));
 sg13g2_inv_1 _09433_ (.Y(_02166_),
    .A(net2226));
 sg13g2_inv_1 _09434_ (.Y(_02167_),
    .A(\mem.mem[126][6] ));
 sg13g2_inv_1 _09435_ (.Y(_02168_),
    .A(\mem.mem[14][7] ));
 sg13g2_inv_1 _09436_ (.Y(_02169_),
    .A(net2732));
 sg13g2_inv_1 _09437_ (.Y(_02170_),
    .A(net2173));
 sg13g2_inv_1 _09438_ (.Y(_02171_),
    .A(net2180));
 sg13g2_inv_1 _09439_ (.Y(_02172_),
    .A(net2776));
 sg13g2_inv_1 _09440_ (.Y(_02173_),
    .A(net4035));
 sg13g2_inv_1 _09441_ (.Y(_02174_),
    .A(\mem.mem[110][7] ));
 sg13g2_inv_1 _09442_ (.Y(_02175_),
    .A(\mem.mem[126][7] ));
 sg13g2_inv_1 _09443_ (.Y(_02176_),
    .A(\mem.mem[142][7] ));
 sg13g2_inv_1 _09444_ (.Y(_02177_),
    .A(\mem.mem[174][7] ));
 sg13g2_inv_1 _09445_ (.Y(_02178_),
    .A(net2458));
 sg13g2_inv_1 _09446_ (.Y(_02179_),
    .A(\mem.mem[206][7] ));
 sg13g2_inv_1 _09447_ (.Y(_02180_),
    .A(net2191));
 sg13g2_inv_1 _09448_ (.Y(_02181_),
    .A(net9));
 sg13g2_inv_1 _09449_ (.Y(_02182_),
    .A(net12));
 sg13g2_inv_1 _09450_ (.Y(_02183_),
    .A(net11));
 sg13g2_inv_1 _09451_ (.Y(_02184_),
    .A(net4008));
 sg13g2_inv_1 _09452_ (.Y(_02185_),
    .A(_00013_));
 sg13g2_inv_1 _09453_ (.Y(_02186_),
    .A(\mem.mem[30][0] ));
 sg13g2_inv_1 _09454_ (.Y(_02187_),
    .A(net2617));
 sg13g2_inv_1 _09455_ (.Y(_02188_),
    .A(net2714));
 sg13g2_nor2_2 _09456_ (.A(net3609),
    .B(net3610),
    .Y(_02189_));
 sg13g2_or2_2 _09457_ (.X(_02190_),
    .B(\state[0] ),
    .A(net3609));
 sg13g2_nand2_2 _09458_ (.Y(_02191_),
    .A(_02136_),
    .B(_02189_));
 sg13g2_inv_1 _09459_ (.Y(halted),
    .A(_02191_));
 sg13g2_and3_1 _09460_ (.X(_02192_),
    .A(net13),
    .B(net12),
    .C(net11));
 sg13g2_nor3_2 _09461_ (.A(net3999),
    .B(_02182_),
    .C(_02183_),
    .Y(_02193_));
 sg13g2_nor2_2 _09462_ (.A(net12),
    .B(net11),
    .Y(_02194_));
 sg13g2_and2_2 _09463_ (.A(net3999),
    .B(_02194_),
    .X(_02195_));
 sg13g2_nor3_2 _09464_ (.A(net3999),
    .B(net12),
    .C(_02183_),
    .Y(_02196_));
 sg13g2_and3_2 _09465_ (.X(_02197_),
    .A(net3999),
    .B(_02182_),
    .C(net11));
 sg13g2_nor3_2 _09466_ (.A(net3999),
    .B(net12),
    .C(net11),
    .Y(_02198_));
 sg13g2_nand2b_2 _09467_ (.Y(_02199_),
    .B(_02194_),
    .A_N(net3999));
 sg13g2_nor3_2 _09468_ (.A(net3999),
    .B(_02182_),
    .C(net11),
    .Y(_02200_));
 sg13g2_and3_2 _09469_ (.X(_02201_),
    .A(net3999),
    .B(net12),
    .C(_02183_));
 sg13g2_a22oi_1 _09470_ (.Y(_02202_),
    .B1(_02197_),
    .B2(\mem_A[0] ),
    .A2(_02192_),
    .A1(net3610));
 sg13g2_a22oi_1 _09471_ (.Y(_02203_),
    .B1(_02200_),
    .B2(\A[0] ),
    .A2(_02196_),
    .A1(\PC[0] ));
 sg13g2_a22oi_1 _09472_ (.Y(_02204_),
    .B1(_02195_),
    .B2(\C[0] ),
    .A2(_02193_),
    .A1(\B[0] ));
 sg13g2_a21oi_1 _09473_ (.A1(net3570),
    .A2(_02201_),
    .Y(_02205_),
    .B1(_02198_));
 sg13g2_nand4_1 _09474_ (.B(_02203_),
    .C(_02204_),
    .A(_02202_),
    .Y(_02206_),
    .D(_02205_));
 sg13g2_o21ai_1 _09475_ (.B1(_02206_),
    .Y(_02207_),
    .A1(\mem.uo_out[0] ),
    .A2(_02199_));
 sg13g2_inv_2 _09476_ (.Y(uo_out[0]),
    .A(_02207_));
 sg13g2_a22oi_1 _09477_ (.Y(_02208_),
    .B1(_02193_),
    .B2(\B[1] ),
    .A2(_02192_),
    .A1(net3609));
 sg13g2_a22oi_1 _09478_ (.Y(_02209_),
    .B1(_02200_),
    .B2(\A[1] ),
    .A2(_02197_),
    .A1(\mem_A[1] ));
 sg13g2_a221oi_1 _09479_ (.B2(net3523),
    .C1(_02198_),
    .B1(_02201_),
    .A1(\C[1] ),
    .Y(_02210_),
    .A2(_02194_));
 sg13g2_nand3_1 _09480_ (.B(_02209_),
    .C(_02210_),
    .A(_02208_),
    .Y(_02211_));
 sg13g2_a21oi_1 _09481_ (.A1(\PC[1] ),
    .A2(_02196_),
    .Y(_02212_),
    .B1(_02211_));
 sg13g2_a21oi_2 _09482_ (.B1(_02212_),
    .Y(uo_out[1]),
    .A2(net3993),
    .A1(_02126_));
 sg13g2_a22oi_1 _09483_ (.Y(_02213_),
    .B1(_02200_),
    .B2(\A[2] ),
    .A2(_02197_),
    .A1(\mem_A[2] ));
 sg13g2_a22oi_1 _09484_ (.Y(_02214_),
    .B1(_02201_),
    .B2(net3476),
    .A2(_02196_),
    .A1(\PC[2] ));
 sg13g2_a22oi_1 _09485_ (.Y(_02215_),
    .B1(_02195_),
    .B2(\C[2] ),
    .A2(_02192_),
    .A1(\state[2] ));
 sg13g2_a21oi_1 _09486_ (.A1(\B[2] ),
    .A2(_02193_),
    .Y(_02216_),
    .B1(net3993));
 sg13g2_nand4_1 _09487_ (.B(_02214_),
    .C(_02215_),
    .A(_02213_),
    .Y(_02217_),
    .D(_02216_));
 sg13g2_o21ai_1 _09488_ (.B1(_02217_),
    .Y(_02218_),
    .A1(\mem.uo_out[2] ),
    .A2(_02199_));
 sg13g2_inv_2 _09489_ (.Y(uo_out[2]),
    .A(_02218_));
 sg13g2_a22oi_1 _09490_ (.Y(_02219_),
    .B1(_02200_),
    .B2(\A[3] ),
    .A2(_02193_),
    .A1(\B[3] ));
 sg13g2_a22oi_1 _09491_ (.Y(_02220_),
    .B1(_02201_),
    .B2(net3431),
    .A2(_02195_),
    .A1(\C[3] ));
 sg13g2_a21oi_1 _09492_ (.A1(\PC[3] ),
    .A2(_02196_),
    .Y(_02221_),
    .B1(net3993));
 sg13g2_nand3_1 _09493_ (.B(_02220_),
    .C(_02221_),
    .A(_02219_),
    .Y(_02222_));
 sg13g2_a21oi_1 _09494_ (.A1(\mem_A[3] ),
    .A2(_02197_),
    .Y(_02223_),
    .B1(_02222_));
 sg13g2_a21oi_2 _09495_ (.B1(_02223_),
    .Y(uo_out[3]),
    .A2(net3993),
    .A1(_02124_));
 sg13g2_a221oi_1 _09496_ (.B2(\PC[4] ),
    .C1(_02198_),
    .B1(_02196_),
    .A1(\C[4] ),
    .Y(_02224_),
    .A2(_02194_));
 sg13g2_a22oi_1 _09497_ (.Y(_02225_),
    .B1(_02200_),
    .B2(\A[4] ),
    .A2(_02197_),
    .A1(\mem_A[4] ));
 sg13g2_a22oi_1 _09498_ (.Y(_02226_),
    .B1(_02201_),
    .B2(net3385),
    .A2(_02193_),
    .A1(\B[4] ));
 sg13g2_nand3_1 _09499_ (.B(_02225_),
    .C(_02226_),
    .A(_02224_),
    .Y(_02227_));
 sg13g2_o21ai_1 _09500_ (.B1(_02227_),
    .Y(_02228_),
    .A1(\mem.uo_out[4] ),
    .A2(_02199_));
 sg13g2_inv_2 _09501_ (.Y(uo_out[4]),
    .A(_02228_));
 sg13g2_a221oi_1 _09502_ (.B2(\A[5] ),
    .C1(net3993),
    .B1(_02200_),
    .A1(\C[5] ),
    .Y(_02229_),
    .A2(_02195_));
 sg13g2_a22oi_1 _09503_ (.Y(_02230_),
    .B1(_02201_),
    .B2(net3339),
    .A2(_02196_),
    .A1(\PC[5] ));
 sg13g2_a22oi_1 _09504_ (.Y(_02231_),
    .B1(_02197_),
    .B2(\mem_A[5] ),
    .A2(_02193_),
    .A1(\B[5] ));
 sg13g2_nand3_1 _09505_ (.B(_02230_),
    .C(_02231_),
    .A(_02229_),
    .Y(_02232_));
 sg13g2_o21ai_1 _09506_ (.B1(_02232_),
    .Y(_02233_),
    .A1(\mem.uo_out[5] ),
    .A2(_02199_));
 sg13g2_inv_2 _09507_ (.Y(uo_out[5]),
    .A(_02233_));
 sg13g2_a221oi_1 _09508_ (.B2(\C[6] ),
    .C1(net3993),
    .B1(_02194_),
    .A1(\B[6] ),
    .Y(_02234_),
    .A2(_02193_));
 sg13g2_a22oi_1 _09509_ (.Y(_02235_),
    .B1(_02200_),
    .B2(\A[6] ),
    .A2(_02196_),
    .A1(\PC[6] ));
 sg13g2_a22oi_1 _09510_ (.Y(_02236_),
    .B1(_02201_),
    .B2(net3293),
    .A2(_02197_),
    .A1(\mem_A[6] ));
 sg13g2_nand3_1 _09511_ (.B(_02235_),
    .C(_02236_),
    .A(_02234_),
    .Y(_02237_));
 sg13g2_o21ai_1 _09512_ (.B1(_02237_),
    .Y(_02238_),
    .A1(\mem.uo_out[6] ),
    .A2(_02199_));
 sg13g2_inv_1 _09513_ (.Y(uo_out[6]),
    .A(_02238_));
 sg13g2_a22oi_1 _09514_ (.Y(_02239_),
    .B1(_02201_),
    .B2(net3247),
    .A2(_02195_),
    .A1(\C[7] ));
 sg13g2_a22oi_1 _09515_ (.Y(_02240_),
    .B1(_02197_),
    .B2(\mem_A[7] ),
    .A2(_02193_),
    .A1(\B[7] ));
 sg13g2_a21oi_1 _09516_ (.A1(\PC[7] ),
    .A2(_02196_),
    .Y(_02241_),
    .B1(net3993));
 sg13g2_nand3_1 _09517_ (.B(_02240_),
    .C(_02241_),
    .A(_02239_),
    .Y(_02242_));
 sg13g2_a21oi_1 _09518_ (.A1(\A[7] ),
    .A2(_02200_),
    .Y(_02243_),
    .B1(_02242_));
 sg13g2_a21oi_2 _09519_ (.B1(_02243_),
    .Y(uo_out[7]),
    .A2(net3993),
    .A1(_02120_));
 sg13g2_and2_2 _09520_ (.A(\mem.addr[3] ),
    .B(net3606),
    .X(_02244_));
 sg13g2_nand2_2 _09521_ (.Y(_02245_),
    .A(\mem.addr[3] ),
    .B(\mem.addr[2] ));
 sg13g2_nor2b_2 _09522_ (.A(net3608),
    .B_N(net3607),
    .Y(_02246_));
 sg13g2_nand2b_2 _09523_ (.Y(_02247_),
    .B(net3607),
    .A_N(net3608));
 sg13g2_nor2_2 _09524_ (.A(_02245_),
    .B(_02247_),
    .Y(_02248_));
 sg13g2_nand2_2 _09525_ (.Y(_02249_),
    .A(_02244_),
    .B(_02246_));
 sg13g2_nor2b_2 _09526_ (.A(\mem.addr[5] ),
    .B_N(net3604),
    .Y(_02250_));
 sg13g2_nand2b_2 _09527_ (.Y(_02251_),
    .B(net3604),
    .A_N(\mem.addr[5] ));
 sg13g2_nand2_1 _09528_ (.Y(_02252_),
    .A(\mem.addr[5] ),
    .B(net3604));
 sg13g2_nand2_2 _09529_ (.Y(_02253_),
    .A(\mem.addr[7] ),
    .B(\mem.addr[6] ));
 sg13g2_nor2_2 _09530_ (.A(net3088),
    .B(_02253_),
    .Y(_02254_));
 sg13g2_or2_1 _09531_ (.X(_02255_),
    .B(_02253_),
    .A(_02252_));
 sg13g2_nor2_1 _09532_ (.A(net3607),
    .B(net3608),
    .Y(_02256_));
 sg13g2_nand2_2 _09533_ (.Y(_02257_),
    .A(_02244_),
    .B(_02254_));
 sg13g2_nor2_2 _09534_ (.A(net3087),
    .B(_02257_),
    .Y(_02258_));
 sg13g2_or2_2 _09535_ (.X(_02259_),
    .B(_02257_),
    .A(net3087));
 sg13g2_nor2_2 _09536_ (.A(_00008_),
    .B(net3996),
    .Y(_02260_));
 sg13g2_nand2b_2 _09537_ (.Y(_02261_),
    .B(net4008),
    .A_N(_00008_));
 sg13g2_nor2_1 _09538_ (.A(_02258_),
    .B(_02261_),
    .Y(_02262_));
 sg13g2_nand2_2 _09539_ (.Y(_02263_),
    .A(_02259_),
    .B(_02260_));
 sg13g2_nor2b_1 _09540_ (.A(\mem.addr[7] ),
    .B_N(net3603),
    .Y(_02264_));
 sg13g2_nand2b_2 _09541_ (.Y(_02265_),
    .B(net3603),
    .A_N(\mem.addr[7] ));
 sg13g2_nor2_2 _09542_ (.A(_02251_),
    .B(_02265_),
    .Y(_02266_));
 sg13g2_nand2_2 _09543_ (.Y(_02267_),
    .A(_02250_),
    .B(_02264_));
 sg13g2_nand2_2 _09544_ (.Y(_02268_),
    .A(net3041),
    .B(net3083));
 sg13g2_nor2_2 _09545_ (.A(_02249_),
    .B(_02268_),
    .Y(_02269_));
 sg13g2_nand2_1 _09546_ (.Y(_02270_),
    .A(net3568),
    .B(_02269_));
 sg13g2_o21ai_1 _09547_ (.B1(_02270_),
    .Y(_00018_),
    .A1(_02188_),
    .A2(_02269_));
 sg13g2_mux2_1 _09548_ (.A0(net2271),
    .A1(net3520),
    .S(net3023),
    .X(_00019_));
 sg13g2_mux2_1 _09549_ (.A0(net2905),
    .A1(net3474),
    .S(net3023),
    .X(_00020_));
 sg13g2_mux2_1 _09550_ (.A0(net2439),
    .A1(net3428),
    .S(net3023),
    .X(_00021_));
 sg13g2_mux2_1 _09551_ (.A0(net2290),
    .A1(net3382),
    .S(net3023),
    .X(_00022_));
 sg13g2_mux2_1 _09552_ (.A0(net2155),
    .A1(net3337),
    .S(net3023),
    .X(_00023_));
 sg13g2_mux2_1 _09553_ (.A0(net2185),
    .A1(net3292),
    .S(net3023),
    .X(_00024_));
 sg13g2_nand2_1 _09554_ (.Y(_02271_),
    .A(net3244),
    .B(net3023));
 sg13g2_o21ai_1 _09555_ (.B1(_02271_),
    .Y(_00025_),
    .A1(_02173_),
    .A2(net3023));
 sg13g2_nor2_2 _09556_ (.A(\mem.addr[5] ),
    .B(net3604),
    .Y(_02272_));
 sg13g2_nor2_2 _09557_ (.A(\mem.addr[7] ),
    .B(net3603),
    .Y(_02273_));
 sg13g2_and2_2 _09558_ (.A(_02272_),
    .B(_02273_),
    .X(_02274_));
 sg13g2_nor2b_2 _09559_ (.A(net3605),
    .B_N(\mem.addr[2] ),
    .Y(_02275_));
 sg13g2_nand2b_2 _09560_ (.Y(_02276_),
    .B(net3606),
    .A_N(net3605));
 sg13g2_and2_2 _09561_ (.A(_02256_),
    .B(_02275_),
    .X(_02277_));
 sg13g2_nand2_2 _09562_ (.Y(_02278_),
    .A(net3087),
    .B(_02275_));
 sg13g2_nand3_1 _09563_ (.B(net3082),
    .C(_02277_),
    .A(_02260_),
    .Y(_02279_));
 sg13g2_mux2_1 _09564_ (.A0(net3582),
    .A1(net2874),
    .S(net3050),
    .X(_00026_));
 sg13g2_mux2_1 _09565_ (.A0(net3538),
    .A1(net4054),
    .S(net3050),
    .X(_00027_));
 sg13g2_nor2_1 _09566_ (.A(net3493),
    .B(net3050),
    .Y(_02280_));
 sg13g2_a21oi_1 _09567_ (.A1(_02151_),
    .A2(net3050),
    .Y(_00028_),
    .B1(_02280_));
 sg13g2_mux2_1 _09568_ (.A0(net3445),
    .A1(net4131),
    .S(net3050),
    .X(_00029_));
 sg13g2_mux2_1 _09569_ (.A0(net3400),
    .A1(net4938),
    .S(_02279_),
    .X(_00030_));
 sg13g2_mux2_1 _09570_ (.A0(net3355),
    .A1(net2828),
    .S(net3050),
    .X(_00031_));
 sg13g2_mux2_1 _09571_ (.A0(net3310),
    .A1(net2735),
    .S(net3050),
    .X(_00032_));
 sg13g2_mux2_1 _09572_ (.A0(net3262),
    .A1(net4162),
    .S(net3050),
    .X(_00033_));
 sg13g2_nor2_2 _09573_ (.A(net3605),
    .B(net3606),
    .Y(_02281_));
 sg13g2_and2_2 _09574_ (.A(net3087),
    .B(_02281_),
    .X(_02282_));
 sg13g2_and2_2 _09575_ (.A(_02260_),
    .B(net3079),
    .X(_02283_));
 sg13g2_nor2b_2 _09576_ (.A(net3088),
    .B_N(_02273_),
    .Y(_02284_));
 sg13g2_nand2b_2 _09577_ (.Y(_02285_),
    .B(_02273_),
    .A_N(net3088));
 sg13g2_nand2_2 _09578_ (.Y(_02286_),
    .A(_02283_),
    .B(_02284_));
 sg13g2_mux2_1 _09579_ (.A0(net3597),
    .A1(net4665),
    .S(_02286_),
    .X(_00034_));
 sg13g2_mux2_1 _09580_ (.A0(net3552),
    .A1(net4509),
    .S(_02286_),
    .X(_00035_));
 sg13g2_mux2_1 _09581_ (.A0(net3505),
    .A1(net2731),
    .S(_02286_),
    .X(_00036_));
 sg13g2_mux2_1 _09582_ (.A0(net3461),
    .A1(net2641),
    .S(_02286_),
    .X(_00037_));
 sg13g2_mux2_1 _09583_ (.A0(net3413),
    .A1(net2911),
    .S(_02286_),
    .X(_00038_));
 sg13g2_mux2_1 _09584_ (.A0(net3369),
    .A1(net4029),
    .S(_02286_),
    .X(_00039_));
 sg13g2_mux2_1 _09585_ (.A0(net3323),
    .A1(net2926),
    .S(_02286_),
    .X(_00040_));
 sg13g2_mux2_1 _09586_ (.A0(net3277),
    .A1(net5057),
    .S(_02286_),
    .X(_00041_));
 sg13g2_nand2_2 _09587_ (.Y(_02287_),
    .A(net3083),
    .B(_02283_));
 sg13g2_mux2_1 _09588_ (.A0(net3569),
    .A1(net4127),
    .S(_02287_),
    .X(_00042_));
 sg13g2_mux2_1 _09589_ (.A0(net3520),
    .A1(net4960),
    .S(_02287_),
    .X(_00043_));
 sg13g2_mux2_1 _09590_ (.A0(net3473),
    .A1(net4303),
    .S(_02287_),
    .X(_00044_));
 sg13g2_mux2_1 _09591_ (.A0(net3429),
    .A1(net2851),
    .S(_02287_),
    .X(_00045_));
 sg13g2_mux2_1 _09592_ (.A0(net3381),
    .A1(net5085),
    .S(_02287_),
    .X(_00046_));
 sg13g2_mux2_1 _09593_ (.A0(net3336),
    .A1(net4571),
    .S(_02287_),
    .X(_00047_));
 sg13g2_mux2_1 _09594_ (.A0(net3291),
    .A1(net5150),
    .S(_02287_),
    .X(_00048_));
 sg13g2_mux2_1 _09595_ (.A0(net3245),
    .A1(net4392),
    .S(_02287_),
    .X(_00049_));
 sg13g2_and2_2 _09596_ (.A(_02246_),
    .B(_02281_),
    .X(_02288_));
 sg13g2_nand2_2 _09597_ (.Y(_02289_),
    .A(_02246_),
    .B(_02281_));
 sg13g2_nand2b_2 _09598_ (.Y(_02290_),
    .B(\mem.addr[5] ),
    .A_N(net3604));
 sg13g2_or3_2 _09599_ (.A(\mem.addr[7] ),
    .B(\mem.addr[6] ),
    .C(_02290_),
    .X(_02291_));
 sg13g2_nor2_2 _09600_ (.A(net3040),
    .B(_02291_),
    .Y(_02292_));
 sg13g2_nor2_2 _09601_ (.A(net3040),
    .B(_02289_),
    .Y(_02293_));
 sg13g2_nand2_2 _09602_ (.Y(_02294_),
    .A(_02288_),
    .B(net3037));
 sg13g2_mux2_1 _09603_ (.A0(net3591),
    .A1(net5114),
    .S(_02294_),
    .X(_00050_));
 sg13g2_mux2_1 _09604_ (.A0(net3547),
    .A1(net4754),
    .S(_02294_),
    .X(_00051_));
 sg13g2_mux2_1 _09605_ (.A0(net3500),
    .A1(net4588),
    .S(_02294_),
    .X(_00052_));
 sg13g2_mux2_1 _09606_ (.A0(net3465),
    .A1(net5013),
    .S(_02294_),
    .X(_00053_));
 sg13g2_mux2_1 _09607_ (.A0(net3409),
    .A1(net4566),
    .S(_02294_),
    .X(_00054_));
 sg13g2_mux2_1 _09608_ (.A0(net3365),
    .A1(net4269),
    .S(_02294_),
    .X(_00055_));
 sg13g2_mux2_1 _09609_ (.A0(net3319),
    .A1(net4870),
    .S(_02294_),
    .X(_00056_));
 sg13g2_mux2_1 _09610_ (.A0(net3270),
    .A1(net4792),
    .S(_02294_),
    .X(_00057_));
 sg13g2_nor2b_2 _09611_ (.A(net3607),
    .B_N(net3608),
    .Y(_02295_));
 sg13g2_nand2b_2 _09612_ (.Y(_02296_),
    .B(net3608),
    .A_N(net3607));
 sg13g2_and2_2 _09613_ (.A(_02281_),
    .B(_02295_),
    .X(_02297_));
 sg13g2_nand2_2 _09614_ (.Y(_02298_),
    .A(_02281_),
    .B(_02295_));
 sg13g2_nor2_2 _09615_ (.A(_02251_),
    .B(_02253_),
    .Y(_02299_));
 sg13g2_and2_2 _09616_ (.A(net3041),
    .B(_02299_),
    .X(_02300_));
 sg13g2_nand2_2 _09617_ (.Y(_02301_),
    .A(net3041),
    .B(net3078));
 sg13g2_nor2_2 _09618_ (.A(_02298_),
    .B(_02301_),
    .Y(_02302_));
 sg13g2_mux2_1 _09619_ (.A0(net2588),
    .A1(net3560),
    .S(_02302_),
    .X(_00058_));
 sg13g2_mux2_1 _09620_ (.A0(net2528),
    .A1(net3516),
    .S(_02302_),
    .X(_00059_));
 sg13g2_mux2_1 _09621_ (.A0(net2524),
    .A1(net3470),
    .S(_02302_),
    .X(_00060_));
 sg13g2_mux2_1 _09622_ (.A0(net2248),
    .A1(net3425),
    .S(_02302_),
    .X(_00061_));
 sg13g2_mux2_1 _09623_ (.A0(net2835),
    .A1(net3377),
    .S(_02302_),
    .X(_00062_));
 sg13g2_mux2_1 _09624_ (.A0(net2696),
    .A1(net3332),
    .S(_02302_),
    .X(_00063_));
 sg13g2_mux2_1 _09625_ (.A0(net2315),
    .A1(net3284),
    .S(_02302_),
    .X(_00064_));
 sg13g2_mux2_1 _09626_ (.A0(net2324),
    .A1(net3241),
    .S(_02302_),
    .X(_00065_));
 sg13g2_nor2_1 _09627_ (.A(_02181_),
    .B(net3994),
    .Y(_00066_));
 sg13g2_and2_2 _09628_ (.A(net3607),
    .B(net3608),
    .X(_02303_));
 sg13g2_nand2_2 _09629_ (.Y(_02304_),
    .A(net3607),
    .B(net3608));
 sg13g2_nand2_2 _09630_ (.Y(_02305_),
    .A(net3606),
    .B(_02303_));
 sg13g2_nor2_2 _09631_ (.A(_02245_),
    .B(_02304_),
    .Y(_02306_));
 sg13g2_nand2_2 _09632_ (.Y(_02307_),
    .A(_02244_),
    .B(_02303_));
 sg13g2_nand2_2 _09633_ (.Y(_02308_),
    .A(net3037),
    .B(_02306_));
 sg13g2_mux2_1 _09634_ (.A0(net3592),
    .A1(net5025),
    .S(_02308_),
    .X(_00067_));
 sg13g2_mux2_1 _09635_ (.A0(net3547),
    .A1(net4094),
    .S(_02308_),
    .X(_00068_));
 sg13g2_mux2_1 _09636_ (.A0(net3506),
    .A1(net4919),
    .S(_02308_),
    .X(_00069_));
 sg13g2_mux2_1 _09637_ (.A0(net3458),
    .A1(net4123),
    .S(_02308_),
    .X(_00070_));
 sg13g2_mux2_1 _09638_ (.A0(net3416),
    .A1(net4831),
    .S(_02308_),
    .X(_00071_));
 sg13g2_mux2_1 _09639_ (.A0(net3371),
    .A1(net4939),
    .S(_02308_),
    .X(_00072_));
 sg13g2_mux2_1 _09640_ (.A0(net3325),
    .A1(net5164),
    .S(_02308_),
    .X(_00073_));
 sg13g2_mux2_1 _09641_ (.A0(net3273),
    .A1(net4832),
    .S(_02308_),
    .X(_00074_));
 sg13g2_nor2_2 _09642_ (.A(_02276_),
    .B(_02304_),
    .Y(_02309_));
 sg13g2_nor3_2 _09643_ (.A(net3605),
    .B(_02261_),
    .C(_02305_),
    .Y(_02310_));
 sg13g2_and2_2 _09644_ (.A(net3043),
    .B(_02274_),
    .X(_02311_));
 sg13g2_nand2_2 _09645_ (.Y(_02312_),
    .A(_02309_),
    .B(_02311_));
 sg13g2_mux2_1 _09646_ (.A0(net3582),
    .A1(net4081),
    .S(_02312_),
    .X(_00075_));
 sg13g2_mux2_1 _09647_ (.A0(net3536),
    .A1(net5157),
    .S(_02312_),
    .X(_00076_));
 sg13g2_mux2_1 _09648_ (.A0(net3493),
    .A1(net4350),
    .S(_02312_),
    .X(_00077_));
 sg13g2_mux2_1 _09649_ (.A0(net3445),
    .A1(net5022),
    .S(_02312_),
    .X(_00078_));
 sg13g2_mux2_1 _09650_ (.A0(net3400),
    .A1(net5134),
    .S(_02312_),
    .X(_00079_));
 sg13g2_mux2_1 _09651_ (.A0(net3358),
    .A1(net4258),
    .S(_02312_),
    .X(_00080_));
 sg13g2_mux2_1 _09652_ (.A0(net3312),
    .A1(net5165),
    .S(_02312_),
    .X(_00081_));
 sg13g2_mux2_1 _09653_ (.A0(net3262),
    .A1(net4142),
    .S(_02312_),
    .X(_00082_));
 sg13g2_and2_2 _09654_ (.A(_02264_),
    .B(_02272_),
    .X(_02313_));
 sg13g2_nand2_2 _09655_ (.Y(_02314_),
    .A(net3041),
    .B(_02313_));
 sg13g2_nor2_2 _09656_ (.A(_02249_),
    .B(_02314_),
    .Y(_02315_));
 sg13g2_nand2_1 _09657_ (.Y(_02316_),
    .A(net3565),
    .B(_02315_));
 sg13g2_o21ai_1 _09658_ (.B1(_02316_),
    .Y(_00083_),
    .A1(_02187_),
    .A2(_02315_));
 sg13g2_mux2_1 _09659_ (.A0(net2594),
    .A1(net3522),
    .S(net3022),
    .X(_00084_));
 sg13g2_mux2_1 _09660_ (.A0(net2375),
    .A1(net3475),
    .S(net3022),
    .X(_00085_));
 sg13g2_mux2_1 _09661_ (.A0(net2475),
    .A1(net3429),
    .S(net3022),
    .X(_00086_));
 sg13g2_mux2_1 _09662_ (.A0(net2495),
    .A1(net3380),
    .S(net3022),
    .X(_00087_));
 sg13g2_mux2_1 _09663_ (.A0(net2344),
    .A1(net3338),
    .S(net3022),
    .X(_00088_));
 sg13g2_mux2_1 _09664_ (.A0(net2136),
    .A1(net3290),
    .S(net3022),
    .X(_00089_));
 sg13g2_nand2_1 _09665_ (.Y(_02317_),
    .A(net3245),
    .B(net3022));
 sg13g2_o21ai_1 _09666_ (.B1(_02317_),
    .Y(_00090_),
    .A1(_02172_),
    .A2(net3022));
 sg13g2_nor2_2 _09667_ (.A(_02245_),
    .B(_02296_),
    .Y(_02318_));
 sg13g2_nor4_2 _09668_ (.A(_02245_),
    .B(net3039),
    .C(_02267_),
    .Y(_02319_),
    .D(_02296_));
 sg13g2_mux2_1 _09669_ (.A0(net2337),
    .A1(net3569),
    .S(_02319_),
    .X(_00091_));
 sg13g2_mux2_1 _09670_ (.A0(net2262),
    .A1(net3522),
    .S(_02319_),
    .X(_00092_));
 sg13g2_mux2_1 _09671_ (.A0(net2314),
    .A1(net3474),
    .S(_02319_),
    .X(_00093_));
 sg13g2_mux2_1 _09672_ (.A0(net2658),
    .A1(net3428),
    .S(_02319_),
    .X(_00094_));
 sg13g2_mux2_1 _09673_ (.A0(net2481),
    .A1(net3382),
    .S(_02319_),
    .X(_00095_));
 sg13g2_mux2_1 _09674_ (.A0(net2682),
    .A1(net3340),
    .S(_02319_),
    .X(_00096_));
 sg13g2_mux2_1 _09675_ (.A0(net2741),
    .A1(net3293),
    .S(_02319_),
    .X(_00097_));
 sg13g2_mux2_1 _09676_ (.A0(net2521),
    .A1(net3244),
    .S(_02319_),
    .X(_00098_));
 sg13g2_nand3_1 _09677_ (.B(net3075),
    .C(net3073),
    .A(net3041),
    .Y(_02320_));
 sg13g2_mux2_1 _09678_ (.A0(net3567),
    .A1(net4349),
    .S(_02320_),
    .X(_00099_));
 sg13g2_mux2_1 _09679_ (.A0(net3522),
    .A1(net4169),
    .S(_02320_),
    .X(_00100_));
 sg13g2_mux2_1 _09680_ (.A0(net3475),
    .A1(net4563),
    .S(_02320_),
    .X(_00101_));
 sg13g2_mux2_1 _09681_ (.A0(net3429),
    .A1(net4466),
    .S(_02320_),
    .X(_00102_));
 sg13g2_mux2_1 _09682_ (.A0(net3380),
    .A1(net4357),
    .S(_02320_),
    .X(_00103_));
 sg13g2_mux2_1 _09683_ (.A0(net3338),
    .A1(net4618),
    .S(_02320_),
    .X(_00104_));
 sg13g2_mux2_1 _09684_ (.A0(net3290),
    .A1(net5140),
    .S(_02320_),
    .X(_00105_));
 sg13g2_mux2_1 _09685_ (.A0(net3245),
    .A1(net4769),
    .S(_02320_),
    .X(_00106_));
 sg13g2_nor4_2 _09686_ (.A(\mem.addr[1] ),
    .B(net3608),
    .C(_02245_),
    .Y(_02321_),
    .D(_02261_));
 sg13g2_nand3_1 _09687_ (.B(net3087),
    .C(_02260_),
    .A(_02244_),
    .Y(_02322_));
 sg13g2_nand2_2 _09688_ (.Y(_02323_),
    .A(net3083),
    .B(net3072));
 sg13g2_mux2_1 _09689_ (.A0(net3568),
    .A1(net4329),
    .S(_02323_),
    .X(_00107_));
 sg13g2_mux2_1 _09690_ (.A0(net3520),
    .A1(net4439),
    .S(_02323_),
    .X(_00108_));
 sg13g2_mux2_1 _09691_ (.A0(net3474),
    .A1(net4656),
    .S(_02323_),
    .X(_00109_));
 sg13g2_mux2_1 _09692_ (.A0(net3428),
    .A1(net2915),
    .S(_02323_),
    .X(_00110_));
 sg13g2_mux2_1 _09693_ (.A0(net3382),
    .A1(net2739),
    .S(_02323_),
    .X(_00111_));
 sg13g2_mux2_1 _09694_ (.A0(net3336),
    .A1(net2704),
    .S(_02323_),
    .X(_00112_));
 sg13g2_mux2_1 _09695_ (.A0(net3292),
    .A1(net2781),
    .S(_02323_),
    .X(_00113_));
 sg13g2_mux2_1 _09696_ (.A0(net3244),
    .A1(net2868),
    .S(_02323_),
    .X(_00114_));
 sg13g2_and2_2 _09697_ (.A(net3075),
    .B(net3072),
    .X(_02324_));
 sg13g2_mux2_1 _09698_ (.A0(net2293),
    .A1(net3567),
    .S(_02324_),
    .X(_00115_));
 sg13g2_mux2_1 _09699_ (.A0(net2373),
    .A1(net3522),
    .S(_02324_),
    .X(_00116_));
 sg13g2_mux2_1 _09700_ (.A0(net2156),
    .A1(net3475),
    .S(_02324_),
    .X(_00117_));
 sg13g2_mux2_1 _09701_ (.A0(net2435),
    .A1(net3429),
    .S(_02324_),
    .X(_00118_));
 sg13g2_mux2_1 _09702_ (.A0(net2366),
    .A1(net3380),
    .S(_02324_),
    .X(_00119_));
 sg13g2_mux2_1 _09703_ (.A0(net2636),
    .A1(net3338),
    .S(_02324_),
    .X(_00120_));
 sg13g2_mux2_1 _09704_ (.A0(net2144),
    .A1(net3290),
    .S(_02324_),
    .X(_00121_));
 sg13g2_mux2_1 _09705_ (.A0(net2660),
    .A1(net3245),
    .S(_02324_),
    .X(_00122_));
 sg13g2_nor2b_2 _09706_ (.A(net3606),
    .B_N(net3605),
    .Y(_02325_));
 sg13g2_nand2b_2 _09707_ (.Y(_02326_),
    .B(net3605),
    .A_N(net3606));
 sg13g2_nor2_2 _09708_ (.A(_02304_),
    .B(_02326_),
    .Y(_02327_));
 sg13g2_and2_2 _09709_ (.A(net3044),
    .B(net3071),
    .X(_02328_));
 sg13g2_nand2_2 _09710_ (.Y(_02329_),
    .A(net3075),
    .B(_02328_));
 sg13g2_mux2_1 _09711_ (.A0(net3565),
    .A1(net4836),
    .S(_02329_),
    .X(_00123_));
 sg13g2_mux2_1 _09712_ (.A0(net3514),
    .A1(net4790),
    .S(_02329_),
    .X(_00124_));
 sg13g2_mux2_1 _09713_ (.A0(net3469),
    .A1(net4354),
    .S(_02329_),
    .X(_00125_));
 sg13g2_mux2_1 _09714_ (.A0(net3424),
    .A1(net4646),
    .S(_02329_),
    .X(_00126_));
 sg13g2_mux2_1 _09715_ (.A0(net3380),
    .A1(net4860),
    .S(_02329_),
    .X(_00127_));
 sg13g2_mux2_1 _09716_ (.A0(net3330),
    .A1(net4456),
    .S(_02329_),
    .X(_00128_));
 sg13g2_mux2_1 _09717_ (.A0(net3290),
    .A1(net4529),
    .S(_02329_),
    .X(_00129_));
 sg13g2_mux2_1 _09718_ (.A0(net3240),
    .A1(net4511),
    .S(_02329_),
    .X(_00130_));
 sg13g2_nor2_2 _09719_ (.A(_02247_),
    .B(_02326_),
    .Y(_02330_));
 sg13g2_nand2_2 _09720_ (.Y(_02331_),
    .A(_02246_),
    .B(_02325_));
 sg13g2_nor2_2 _09721_ (.A(net3039),
    .B(_02331_),
    .Y(_02332_));
 sg13g2_nand2_2 _09722_ (.Y(_02333_),
    .A(net3075),
    .B(_02332_));
 sg13g2_mux2_1 _09723_ (.A0(net3565),
    .A1(net4568),
    .S(_02333_),
    .X(_00131_));
 sg13g2_mux2_1 _09724_ (.A0(net3514),
    .A1(net2787),
    .S(_02333_),
    .X(_00132_));
 sg13g2_mux2_1 _09725_ (.A0(net3469),
    .A1(net4908),
    .S(_02333_),
    .X(_00133_));
 sg13g2_mux2_1 _09726_ (.A0(net3424),
    .A1(net2939),
    .S(_02333_),
    .X(_00134_));
 sg13g2_mux2_1 _09727_ (.A0(net3380),
    .A1(net4944),
    .S(_02333_),
    .X(_00135_));
 sg13g2_mux2_1 _09728_ (.A0(net3330),
    .A1(net2956),
    .S(_02333_),
    .X(_00136_));
 sg13g2_mux2_1 _09729_ (.A0(net3290),
    .A1(net4988),
    .S(_02333_),
    .X(_00137_));
 sg13g2_mux2_1 _09730_ (.A0(net3240),
    .A1(net4308),
    .S(_02333_),
    .X(_00138_));
 sg13g2_nor2_2 _09731_ (.A(_02296_),
    .B(_02326_),
    .Y(_02334_));
 sg13g2_nand2_2 _09732_ (.Y(_02335_),
    .A(_02295_),
    .B(_02325_));
 sg13g2_nor2_2 _09733_ (.A(_02314_),
    .B(_02335_),
    .Y(_02336_));
 sg13g2_mux2_1 _09734_ (.A0(net2477),
    .A1(net3565),
    .S(_02336_),
    .X(_00139_));
 sg13g2_mux2_1 _09735_ (.A0(net2501),
    .A1(net3515),
    .S(_02336_),
    .X(_00140_));
 sg13g2_mux2_1 _09736_ (.A0(net2496),
    .A1(net3469),
    .S(_02336_),
    .X(_00141_));
 sg13g2_mux2_1 _09737_ (.A0(net2511),
    .A1(net3424),
    .S(_02336_),
    .X(_00142_));
 sg13g2_mux2_1 _09738_ (.A0(net2385),
    .A1(net3380),
    .S(_02336_),
    .X(_00143_));
 sg13g2_mux2_1 _09739_ (.A0(net2339),
    .A1(net3330),
    .S(_02336_),
    .X(_00144_));
 sg13g2_mux2_1 _09740_ (.A0(net2291),
    .A1(net3290),
    .S(_02336_),
    .X(_00145_));
 sg13g2_mux2_1 _09741_ (.A0(net2469),
    .A1(net3240),
    .S(_02336_),
    .X(_00146_));
 sg13g2_and2_2 _09742_ (.A(net3087),
    .B(_02325_),
    .X(_02337_));
 sg13g2_nand2_2 _09743_ (.Y(_02338_),
    .A(net3087),
    .B(_02325_));
 sg13g2_nor2_2 _09744_ (.A(_02261_),
    .B(_02338_),
    .Y(_02339_));
 sg13g2_nand2_2 _09745_ (.Y(_02340_),
    .A(_02260_),
    .B(_02337_));
 sg13g2_and2_2 _09746_ (.A(net3075),
    .B(_02339_),
    .X(_02341_));
 sg13g2_mux2_1 _09747_ (.A0(net2351),
    .A1(net3565),
    .S(_02341_),
    .X(_00147_));
 sg13g2_mux2_1 _09748_ (.A0(net2153),
    .A1(net3514),
    .S(_02341_),
    .X(_00148_));
 sg13g2_mux2_1 _09749_ (.A0(net2620),
    .A1(net3469),
    .S(_02341_),
    .X(_00149_));
 sg13g2_mux2_1 _09750_ (.A0(net2551),
    .A1(net3424),
    .S(_02341_),
    .X(_00150_));
 sg13g2_mux2_1 _09751_ (.A0(net2536),
    .A1(net3380),
    .S(_02341_),
    .X(_00151_));
 sg13g2_mux2_1 _09752_ (.A0(net2578),
    .A1(net3330),
    .S(_02341_),
    .X(_00152_));
 sg13g2_mux2_1 _09753_ (.A0(net2436),
    .A1(net3290),
    .S(_02341_),
    .X(_00153_));
 sg13g2_mux2_1 _09754_ (.A0(net2323),
    .A1(net3240),
    .S(_02341_),
    .X(_00154_));
 sg13g2_nand2_1 _09755_ (.Y(_02342_),
    .A(net3085),
    .B(net3037));
 sg13g2_mux2_1 _09756_ (.A0(net3594),
    .A1(net2826),
    .S(net3021),
    .X(_00155_));
 sg13g2_mux2_1 _09757_ (.A0(net3548),
    .A1(net4949),
    .S(net3021),
    .X(_00156_));
 sg13g2_mux2_1 _09758_ (.A0(net3506),
    .A1(net4384),
    .S(net3021),
    .X(_00157_));
 sg13g2_mux2_1 _09759_ (.A0(net3458),
    .A1(net4838),
    .S(net3021),
    .X(_00158_));
 sg13g2_mux2_1 _09760_ (.A0(net3416),
    .A1(net4207),
    .S(net3021),
    .X(_00159_));
 sg13g2_mux2_1 _09761_ (.A0(net3371),
    .A1(net2717),
    .S(net3021),
    .X(_00160_));
 sg13g2_nor2_1 _09762_ (.A(net3324),
    .B(net3021),
    .Y(_02343_));
 sg13g2_a21oi_1 _09763_ (.A1(_02164_),
    .A2(net3021),
    .Y(_00161_),
    .B1(_02343_));
 sg13g2_nor2_1 _09764_ (.A(net3273),
    .B(_02342_),
    .Y(_02344_));
 sg13g2_a21oi_1 _09765_ (.A1(_02170_),
    .A2(_02342_),
    .Y(_00162_),
    .B1(_02344_));
 sg13g2_nor2_2 _09766_ (.A(_02276_),
    .B(_02296_),
    .Y(_02345_));
 sg13g2_and2_2 _09767_ (.A(net3043),
    .B(_02345_),
    .X(_02346_));
 sg13g2_nor2b_2 _09768_ (.A(_02314_),
    .B_N(net3069),
    .Y(_02347_));
 sg13g2_mux2_1 _09769_ (.A0(net2359),
    .A1(net3570),
    .S(_02347_),
    .X(_00163_));
 sg13g2_mux2_1 _09770_ (.A0(net2556),
    .A1(net3523),
    .S(_02347_),
    .X(_00164_));
 sg13g2_mux2_1 _09771_ (.A0(net2520),
    .A1(net3476),
    .S(_02347_),
    .X(_00165_));
 sg13g2_mux2_1 _09772_ (.A0(net2581),
    .A1(net3430),
    .S(_02347_),
    .X(_00166_));
 sg13g2_mux2_1 _09773_ (.A0(net2194),
    .A1(net3384),
    .S(_02347_),
    .X(_00167_));
 sg13g2_mux2_1 _09774_ (.A0(net2675),
    .A1(net3339),
    .S(_02347_),
    .X(_00168_));
 sg13g2_mux2_1 _09775_ (.A0(net2754),
    .A1(net3295),
    .S(_02347_),
    .X(_00169_));
 sg13g2_mux2_1 _09776_ (.A0(net2585),
    .A1(net3246),
    .S(_02347_),
    .X(_00170_));
 sg13g2_nand2_2 _09777_ (.Y(_02348_),
    .A(net3037),
    .B(net3074));
 sg13g2_mux2_1 _09778_ (.A0(net3592),
    .A1(net4266),
    .S(_02348_),
    .X(_00171_));
 sg13g2_mux2_1 _09779_ (.A0(net3552),
    .A1(net4858),
    .S(_02348_),
    .X(_00172_));
 sg13g2_mux2_1 _09780_ (.A0(net3506),
    .A1(net4355),
    .S(_02348_),
    .X(_00173_));
 sg13g2_mux2_1 _09781_ (.A0(net3462),
    .A1(net4877),
    .S(_02348_),
    .X(_00174_));
 sg13g2_mux2_1 _09782_ (.A0(net3416),
    .A1(net4572),
    .S(_02348_),
    .X(_00175_));
 sg13g2_mux2_1 _09783_ (.A0(net3371),
    .A1(net4996),
    .S(_02348_),
    .X(_00176_));
 sg13g2_mux2_1 _09784_ (.A0(net3324),
    .A1(net5068),
    .S(_02348_),
    .X(_00177_));
 sg13g2_mux2_1 _09785_ (.A0(net3273),
    .A1(net4323),
    .S(_02348_),
    .X(_00178_));
 sg13g2_and2_2 _09786_ (.A(_02281_),
    .B(_02303_),
    .X(_02349_));
 sg13g2_nand2_2 _09787_ (.Y(_02350_),
    .A(_02250_),
    .B(_02273_));
 sg13g2_nor2_2 _09788_ (.A(net3040),
    .B(_02350_),
    .Y(_02351_));
 sg13g2_nand2_2 _09789_ (.Y(_02352_),
    .A(_02349_),
    .B(net3034));
 sg13g2_and2_2 _09790_ (.A(net3043),
    .B(_02349_),
    .X(_02353_));
 sg13g2_mux2_1 _09791_ (.A0(net3591),
    .A1(net4450),
    .S(_02352_),
    .X(_00179_));
 sg13g2_mux2_1 _09792_ (.A0(net3545),
    .A1(net4770),
    .S(_02352_),
    .X(_00180_));
 sg13g2_mux2_1 _09793_ (.A0(net3499),
    .A1(net4684),
    .S(_02352_),
    .X(_00181_));
 sg13g2_mux2_1 _09794_ (.A0(net3454),
    .A1(net4578),
    .S(_02352_),
    .X(_00182_));
 sg13g2_mux2_1 _09795_ (.A0(net3408),
    .A1(net4958),
    .S(_02352_),
    .X(_00183_));
 sg13g2_mux2_1 _09796_ (.A0(net3366),
    .A1(net4512),
    .S(_02352_),
    .X(_00184_));
 sg13g2_mux2_1 _09797_ (.A0(net3320),
    .A1(net5044),
    .S(_02352_),
    .X(_00185_));
 sg13g2_mux2_1 _09798_ (.A0(net3270),
    .A1(net4159),
    .S(_02352_),
    .X(_00186_));
 sg13g2_nand2b_2 _09799_ (.Y(_02354_),
    .B(\mem.addr[7] ),
    .A_N(net3603));
 sg13g2_nor3_1 _09800_ (.A(net3088),
    .B(net3039),
    .C(_02354_),
    .Y(_02355_));
 sg13g2_nand2_2 _09801_ (.Y(_02356_),
    .A(_02349_),
    .B(net3031));
 sg13g2_mux2_1 _09802_ (.A0(net3579),
    .A1(net4208),
    .S(_02356_),
    .X(_00187_));
 sg13g2_mux2_1 _09803_ (.A0(net3532),
    .A1(net4716),
    .S(_02356_),
    .X(_00188_));
 sg13g2_mux2_1 _09804_ (.A0(net3486),
    .A1(net4363),
    .S(_02356_),
    .X(_00189_));
 sg13g2_mux2_1 _09805_ (.A0(net3448),
    .A1(net4676),
    .S(_02356_),
    .X(_00190_));
 sg13g2_mux2_1 _09806_ (.A0(net3404),
    .A1(net5067),
    .S(_02356_),
    .X(_00191_));
 sg13g2_mux2_1 _09807_ (.A0(net3350),
    .A1(net4088),
    .S(_02356_),
    .X(_00192_));
 sg13g2_mux2_1 _09808_ (.A0(net3305),
    .A1(net5065),
    .S(_02356_),
    .X(_00193_));
 sg13g2_mux2_1 _09809_ (.A0(net3264),
    .A1(net5180),
    .S(_02356_),
    .X(_00194_));
 sg13g2_nor2_2 _09810_ (.A(_02291_),
    .B(_02322_),
    .Y(_02357_));
 sg13g2_mux2_1 _09811_ (.A0(net2408),
    .A1(net3594),
    .S(_02357_),
    .X(_00195_));
 sg13g2_mux2_1 _09812_ (.A0(net2810),
    .A1(net3552),
    .S(_02357_),
    .X(_00196_));
 sg13g2_mux2_1 _09813_ (.A0(net2539),
    .A1(net3506),
    .S(_02357_),
    .X(_00197_));
 sg13g2_mux2_1 _09814_ (.A0(net2645),
    .A1(net3458),
    .S(_02357_),
    .X(_00198_));
 sg13g2_mux2_1 _09815_ (.A0(net2340),
    .A1(net3416),
    .S(_02357_),
    .X(_00199_));
 sg13g2_mux2_1 _09816_ (.A0(net2158),
    .A1(net3371),
    .S(_02357_),
    .X(_00200_));
 sg13g2_mux2_1 _09817_ (.A0(net2140),
    .A1(net3324),
    .S(_02357_),
    .X(_00201_));
 sg13g2_mux2_1 _09818_ (.A0(net2440),
    .A1(net3273),
    .S(_02357_),
    .X(_00202_));
 sg13g2_nor2_1 _09819_ (.A(net3088),
    .B(_02265_),
    .Y(_02358_));
 sg13g2_nand2_2 _09820_ (.Y(_02359_),
    .A(net3042),
    .B(net3068));
 sg13g2_nand2_2 _09821_ (.Y(_02360_),
    .A(net3049),
    .B(net3067));
 sg13g2_mux2_1 _09822_ (.A0(net3563),
    .A1(net4536),
    .S(_02360_),
    .X(_00203_));
 sg13g2_mux2_1 _09823_ (.A0(net3525),
    .A1(net4444),
    .S(_02360_),
    .X(_00204_));
 sg13g2_mux2_1 _09824_ (.A0(net3481),
    .A1(net4200),
    .S(_02360_),
    .X(_00205_));
 sg13g2_mux2_1 _09825_ (.A0(net3435),
    .A1(net4946),
    .S(_02360_),
    .X(_00206_));
 sg13g2_mux2_1 _09826_ (.A0(net3389),
    .A1(net4634),
    .S(_02360_),
    .X(_00207_));
 sg13g2_mux2_1 _09827_ (.A0(net3342),
    .A1(net4455),
    .S(_02360_),
    .X(_00208_));
 sg13g2_mux2_1 _09828_ (.A0(net3302),
    .A1(net4708),
    .S(_02360_),
    .X(_00209_));
 sg13g2_mux2_1 _09829_ (.A0(net3248),
    .A1(net4503),
    .S(_02360_),
    .X(_00210_));
 sg13g2_nand2_2 _09830_ (.Y(_02361_),
    .A(net3038),
    .B(net3071));
 sg13g2_mux2_1 _09831_ (.A0(net3594),
    .A1(net4078),
    .S(_02361_),
    .X(_00211_));
 sg13g2_mux2_1 _09832_ (.A0(net3548),
    .A1(net4687),
    .S(_02361_),
    .X(_00212_));
 sg13g2_mux2_1 _09833_ (.A0(net3507),
    .A1(net4623),
    .S(_02361_),
    .X(_00213_));
 sg13g2_mux2_1 _09834_ (.A0(net3459),
    .A1(net4977),
    .S(_02361_),
    .X(_00214_));
 sg13g2_mux2_1 _09835_ (.A0(net3416),
    .A1(net2995),
    .S(_02361_),
    .X(_00215_));
 sg13g2_mux2_1 _09836_ (.A0(net3373),
    .A1(net5092),
    .S(_02361_),
    .X(_00216_));
 sg13g2_mux2_1 _09837_ (.A0(net3325),
    .A1(net4018),
    .S(_02361_),
    .X(_00217_));
 sg13g2_mux2_1 _09838_ (.A0(net3274),
    .A1(net4233),
    .S(_02361_),
    .X(_00218_));
 sg13g2_nor2_2 _09839_ (.A(_02290_),
    .B(_02354_),
    .Y(_02362_));
 sg13g2_and2_1 _09840_ (.A(net3043),
    .B(_02362_),
    .X(_02363_));
 sg13g2_nand2_2 _09841_ (.Y(_02364_),
    .A(net3070),
    .B(net3030));
 sg13g2_mux2_1 _09842_ (.A0(net3579),
    .A1(net4399),
    .S(_02364_),
    .X(_00219_));
 sg13g2_mux2_1 _09843_ (.A0(net3540),
    .A1(net4577),
    .S(_02364_),
    .X(_00220_));
 sg13g2_mux2_1 _09844_ (.A0(net3485),
    .A1(net4979),
    .S(_02364_),
    .X(_00221_));
 sg13g2_mux2_1 _09845_ (.A0(net3447),
    .A1(net4758),
    .S(_02364_),
    .X(_00222_));
 sg13g2_mux2_1 _09846_ (.A0(net3395),
    .A1(net4852),
    .S(_02364_),
    .X(_00223_));
 sg13g2_mux2_1 _09847_ (.A0(net3349),
    .A1(net4817),
    .S(_02364_),
    .X(_00224_));
 sg13g2_mux2_1 _09848_ (.A0(net3305),
    .A1(net4446),
    .S(_02364_),
    .X(_00225_));
 sg13g2_mux2_1 _09849_ (.A0(net3254),
    .A1(net4324),
    .S(_02364_),
    .X(_00226_));
 sg13g2_nor2_2 _09850_ (.A(_02251_),
    .B(_02354_),
    .Y(_02365_));
 sg13g2_and2_1 _09851_ (.A(net3043),
    .B(_02365_),
    .X(_02366_));
 sg13g2_and2_2 _09852_ (.A(_02306_),
    .B(net3027),
    .X(_02367_));
 sg13g2_mux2_1 _09853_ (.A0(net2219),
    .A1(net3597),
    .S(_02367_),
    .X(_00227_));
 sg13g2_mux2_1 _09854_ (.A0(net2621),
    .A1(net3551),
    .S(_02367_),
    .X(_00228_));
 sg13g2_mux2_1 _09855_ (.A0(net2600),
    .A1(net3505),
    .S(_02367_),
    .X(_00229_));
 sg13g2_mux2_1 _09856_ (.A0(net2667),
    .A1(net3460),
    .S(_02367_),
    .X(_00230_));
 sg13g2_mux2_1 _09857_ (.A0(net2780),
    .A1(net3415),
    .S(_02367_),
    .X(_00231_));
 sg13g2_mux2_1 _09858_ (.A0(net2389),
    .A1(net3362),
    .S(_02367_),
    .X(_00232_));
 sg13g2_mux2_1 _09859_ (.A0(net2519),
    .A1(net3317),
    .S(_02367_),
    .X(_00233_));
 sg13g2_mux2_1 _09860_ (.A0(net2560),
    .A1(net3276),
    .S(_02367_),
    .X(_00234_));
 sg13g2_nor2_2 _09861_ (.A(net3076),
    .B(_02314_),
    .Y(_02368_));
 sg13g2_mux2_1 _09862_ (.A0(net2303),
    .A1(net3565),
    .S(_02368_),
    .X(_00235_));
 sg13g2_mux2_1 _09863_ (.A0(net2498),
    .A1(net3522),
    .S(_02368_),
    .X(_00236_));
 sg13g2_mux2_1 _09864_ (.A0(net2611),
    .A1(net3475),
    .S(_02368_),
    .X(_00237_));
 sg13g2_mux2_1 _09865_ (.A0(net2414),
    .A1(net3429),
    .S(_02368_),
    .X(_00238_));
 sg13g2_mux2_1 _09866_ (.A0(net2543),
    .A1(net3380),
    .S(_02368_),
    .X(_00239_));
 sg13g2_mux2_1 _09867_ (.A0(net2295),
    .A1(net3338),
    .S(_02368_),
    .X(_00240_));
 sg13g2_mux2_1 _09868_ (.A0(net2434),
    .A1(net3290),
    .S(_02368_),
    .X(_00241_));
 sg13g2_mux2_1 _09869_ (.A0(net2494),
    .A1(net3245),
    .S(_02368_),
    .X(_00242_));
 sg13g2_nand3b_1 _09870_ (.B(_02272_),
    .C(\mem.addr[7] ),
    .Y(_02369_),
    .A_N(net3603));
 sg13g2_nor2_2 _09871_ (.A(net3040),
    .B(_02369_),
    .Y(_02370_));
 sg13g2_or2_2 _09872_ (.X(_02371_),
    .B(_02369_),
    .A(net3040));
 sg13g2_nor2_2 _09873_ (.A(_02298_),
    .B(_02371_),
    .Y(_02372_));
 sg13g2_mux2_1 _09874_ (.A0(net2744),
    .A1(net3584),
    .S(_02372_),
    .X(_00243_));
 sg13g2_mux2_1 _09875_ (.A0(net2227),
    .A1(net3537),
    .S(_02372_),
    .X(_00244_));
 sg13g2_mux2_1 _09876_ (.A0(net2489),
    .A1(net3492),
    .S(_02372_),
    .X(_00245_));
 sg13g2_mux2_1 _09877_ (.A0(net2367),
    .A1(net3448),
    .S(_02372_),
    .X(_00246_));
 sg13g2_mux2_1 _09878_ (.A0(net2765),
    .A1(net3405),
    .S(_02372_),
    .X(_00247_));
 sg13g2_mux2_1 _09879_ (.A0(net2792),
    .A1(net3356),
    .S(_02372_),
    .X(_00248_));
 sg13g2_mux2_1 _09880_ (.A0(net2534),
    .A1(net3311),
    .S(_02372_),
    .X(_00249_));
 sg13g2_mux2_1 _09881_ (.A0(net2297),
    .A1(net3261),
    .S(_02372_),
    .X(_00250_));
 sg13g2_nand2_2 _09882_ (.Y(_02373_),
    .A(_02345_),
    .B(net3028));
 sg13g2_mux2_1 _09883_ (.A0(net3598),
    .A1(net4471),
    .S(_02373_),
    .X(_00251_));
 sg13g2_mux2_1 _09884_ (.A0(net3553),
    .A1(net4136),
    .S(_02373_),
    .X(_00252_));
 sg13g2_mux2_1 _09885_ (.A0(net3508),
    .A1(net5124),
    .S(_02373_),
    .X(_00253_));
 sg13g2_mux2_1 _09886_ (.A0(net3463),
    .A1(net4514),
    .S(_02373_),
    .X(_00254_));
 sg13g2_mux2_1 _09887_ (.A0(net3418),
    .A1(net4589),
    .S(_02373_),
    .X(_00255_));
 sg13g2_mux2_1 _09888_ (.A0(net3372),
    .A1(net2892),
    .S(_02373_),
    .X(_00256_));
 sg13g2_mux2_1 _09889_ (.A0(net3326),
    .A1(net4291),
    .S(_02373_),
    .X(_00257_));
 sg13g2_mux2_1 _09890_ (.A0(net3278),
    .A1(net2984),
    .S(_02373_),
    .X(_00258_));
 sg13g2_nand2_2 _09891_ (.Y(_02374_),
    .A(net3038),
    .B(_02330_));
 sg13g2_mux2_1 _09892_ (.A0(net3594),
    .A1(net4398),
    .S(_02374_),
    .X(_00259_));
 sg13g2_mux2_1 _09893_ (.A0(net3548),
    .A1(net4847),
    .S(_02374_),
    .X(_00260_));
 sg13g2_mux2_1 _09894_ (.A0(net3507),
    .A1(net4261),
    .S(_02374_),
    .X(_00261_));
 sg13g2_mux2_1 _09895_ (.A0(net3459),
    .A1(net4408),
    .S(_02374_),
    .X(_00262_));
 sg13g2_mux2_1 _09896_ (.A0(net3416),
    .A1(net4336),
    .S(_02374_),
    .X(_00263_));
 sg13g2_mux2_1 _09897_ (.A0(net3373),
    .A1(net4394),
    .S(_02374_),
    .X(_00264_));
 sg13g2_mux2_1 _09898_ (.A0(net3325),
    .A1(net2987),
    .S(_02374_),
    .X(_00265_));
 sg13g2_mux2_1 _09899_ (.A0(net3274),
    .A1(net4249),
    .S(_02374_),
    .X(_00266_));
 sg13g2_nor2_2 _09900_ (.A(net3039),
    .B(_02285_),
    .Y(_02375_));
 sg13g2_nand2_2 _09901_ (.Y(_02376_),
    .A(net3071),
    .B(_02375_));
 sg13g2_mux2_1 _09902_ (.A0(net3599),
    .A1(net2957),
    .S(_02376_),
    .X(_00267_));
 sg13g2_mux2_1 _09903_ (.A0(net3554),
    .A1(net4376),
    .S(_02376_),
    .X(_00268_));
 sg13g2_mux2_1 _09904_ (.A0(net3507),
    .A1(net4055),
    .S(_02376_),
    .X(_00269_));
 sg13g2_mux2_1 _09905_ (.A0(net3464),
    .A1(net5090),
    .S(_02376_),
    .X(_00270_));
 sg13g2_mux2_1 _09906_ (.A0(net3417),
    .A1(net4779),
    .S(_02376_),
    .X(_00271_));
 sg13g2_mux2_1 _09907_ (.A0(net3373),
    .A1(net5036),
    .S(_02376_),
    .X(_00272_));
 sg13g2_mux2_1 _09908_ (.A0(net3327),
    .A1(net2930),
    .S(_02376_),
    .X(_00273_));
 sg13g2_mux2_1 _09909_ (.A0(net3280),
    .A1(net5039),
    .S(_02376_),
    .X(_00274_));
 sg13g2_nand2_2 _09910_ (.Y(_02377_),
    .A(net3038),
    .B(_02334_));
 sg13g2_mux2_1 _09911_ (.A0(net3593),
    .A1(net4679),
    .S(_02377_),
    .X(_00275_));
 sg13g2_mux2_1 _09912_ (.A0(net3548),
    .A1(net5108),
    .S(_02377_),
    .X(_00276_));
 sg13g2_mux2_1 _09913_ (.A0(net3506),
    .A1(net4741),
    .S(_02377_),
    .X(_00277_));
 sg13g2_mux2_1 _09914_ (.A0(net3458),
    .A1(net4898),
    .S(_02377_),
    .X(_00278_));
 sg13g2_mux2_1 _09915_ (.A0(net3416),
    .A1(net4429),
    .S(_02377_),
    .X(_00279_));
 sg13g2_mux2_1 _09916_ (.A0(net3371),
    .A1(net5176),
    .S(_02377_),
    .X(_00280_));
 sg13g2_mux2_1 _09917_ (.A0(net3325),
    .A1(net4906),
    .S(_02377_),
    .X(_00281_));
 sg13g2_mux2_1 _09918_ (.A0(net3274),
    .A1(net4968),
    .S(_02377_),
    .X(_00282_));
 sg13g2_nor2_2 _09919_ (.A(_02291_),
    .B(_02340_),
    .Y(_02378_));
 sg13g2_mux2_1 _09920_ (.A0(net2546),
    .A1(net3593),
    .S(_02378_),
    .X(_00283_));
 sg13g2_mux2_1 _09921_ (.A0(net2508),
    .A1(net3548),
    .S(_02378_),
    .X(_00284_));
 sg13g2_mux2_1 _09922_ (.A0(net2187),
    .A1(net3506),
    .S(_02378_),
    .X(_00285_));
 sg13g2_mux2_1 _09923_ (.A0(net2453),
    .A1(net3459),
    .S(_02378_),
    .X(_00286_));
 sg13g2_mux2_1 _09924_ (.A0(net2393),
    .A1(net3416),
    .S(_02378_),
    .X(_00287_));
 sg13g2_mux2_1 _09925_ (.A0(net2470),
    .A1(net3371),
    .S(_02378_),
    .X(_00288_));
 sg13g2_mux2_1 _09926_ (.A0(net2418),
    .A1(net3325),
    .S(_02378_),
    .X(_00289_));
 sg13g2_mux2_1 _09927_ (.A0(net2584),
    .A1(net3274),
    .S(_02378_),
    .X(_00290_));
 sg13g2_nor2b_2 _09928_ (.A(_02253_),
    .B_N(_02272_),
    .Y(_02379_));
 sg13g2_nand2_2 _09929_ (.Y(_02380_),
    .A(net3049),
    .B(net3066));
 sg13g2_nand2_2 _09930_ (.Y(_02381_),
    .A(net3041),
    .B(_02379_));
 sg13g2_mux2_1 _09931_ (.A0(net3558),
    .A1(net4913),
    .S(_02380_),
    .X(_00291_));
 sg13g2_mux2_1 _09932_ (.A0(net3513),
    .A1(net2983),
    .S(_02380_),
    .X(_00292_));
 sg13g2_mux2_1 _09933_ (.A0(net3468),
    .A1(net4062),
    .S(_02380_),
    .X(_00293_));
 sg13g2_mux2_1 _09934_ (.A0(net3423),
    .A1(net4063),
    .S(_02380_),
    .X(_00294_));
 sg13g2_mux2_1 _09935_ (.A0(net3375),
    .A1(net4751),
    .S(_02380_),
    .X(_00295_));
 sg13g2_mux2_1 _09936_ (.A0(net3331),
    .A1(net4404),
    .S(_02380_),
    .X(_00296_));
 sg13g2_mux2_1 _09937_ (.A0(net3283),
    .A1(net4659),
    .S(_02380_),
    .X(_00297_));
 sg13g2_mux2_1 _09938_ (.A0(net3239),
    .A1(net4468),
    .S(_02380_),
    .X(_00298_));
 sg13g2_nand2_2 _09939_ (.Y(_02382_),
    .A(_02274_),
    .B(_02353_));
 sg13g2_mux2_1 _09940_ (.A0(net3590),
    .A1(net5075),
    .S(_02382_),
    .X(_00299_));
 sg13g2_mux2_1 _09941_ (.A0(net3545),
    .A1(net4599),
    .S(_02382_),
    .X(_00300_));
 sg13g2_mux2_1 _09942_ (.A0(net3501),
    .A1(net5080),
    .S(_02382_),
    .X(_00301_));
 sg13g2_mux2_1 _09943_ (.A0(net3454),
    .A1(net4373),
    .S(_02382_),
    .X(_00302_));
 sg13g2_mux2_1 _09944_ (.A0(net3408),
    .A1(net4881),
    .S(_02382_),
    .X(_00303_));
 sg13g2_mux2_1 _09945_ (.A0(net3355),
    .A1(net5131),
    .S(_02382_),
    .X(_00304_));
 sg13g2_mux2_1 _09946_ (.A0(net3320),
    .A1(net5005),
    .S(_02382_),
    .X(_00305_));
 sg13g2_mux2_1 _09947_ (.A0(net3269),
    .A1(net5016),
    .S(_02382_),
    .X(_00306_));
 sg13g2_nor2_2 _09948_ (.A(_02247_),
    .B(_02276_),
    .Y(_02383_));
 sg13g2_nand2_2 _09949_ (.Y(_02384_),
    .A(net3037),
    .B(net3065));
 sg13g2_and2_2 _09950_ (.A(net3044),
    .B(net3065),
    .X(_02385_));
 sg13g2_mux2_1 _09951_ (.A0(net3592),
    .A1(net4150),
    .S(net3020),
    .X(_00307_));
 sg13g2_mux2_1 _09952_ (.A0(net3550),
    .A1(net2777),
    .S(net3020),
    .X(_00308_));
 sg13g2_nor2_1 _09953_ (.A(net3503),
    .B(net3020),
    .Y(_02386_));
 sg13g2_a21oi_1 _09954_ (.A1(_02153_),
    .A2(net3020),
    .Y(_00309_),
    .B1(_02386_));
 sg13g2_mux2_1 _09955_ (.A0(net3458),
    .A1(net4307),
    .S(net3020),
    .X(_00310_));
 sg13g2_mux2_1 _09956_ (.A0(net3412),
    .A1(net4202),
    .S(net3020),
    .X(_00311_));
 sg13g2_mux2_1 _09957_ (.A0(net3368),
    .A1(net4041),
    .S(_02384_),
    .X(_00312_));
 sg13g2_mux2_1 _09958_ (.A0(net3322),
    .A1(net4819),
    .S(net3020),
    .X(_00313_));
 sg13g2_mux2_1 _09959_ (.A0(net3273),
    .A1(net2972),
    .S(net3020),
    .X(_00314_));
 sg13g2_nand2_2 _09960_ (.Y(_02387_),
    .A(net3073),
    .B(net3031));
 sg13g2_mux2_1 _09961_ (.A0(net3578),
    .A1(net4742),
    .S(_02387_),
    .X(_00315_));
 sg13g2_mux2_1 _09962_ (.A0(net3530),
    .A1(net4795),
    .S(_02387_),
    .X(_00316_));
 sg13g2_mux2_1 _09963_ (.A0(net3484),
    .A1(net5073),
    .S(_02387_),
    .X(_00317_));
 sg13g2_mux2_1 _09964_ (.A0(net3439),
    .A1(net5097),
    .S(_02387_),
    .X(_00318_));
 sg13g2_mux2_1 _09965_ (.A0(net3394),
    .A1(net4228),
    .S(_02387_),
    .X(_00319_));
 sg13g2_mux2_1 _09966_ (.A0(net3347),
    .A1(net4984),
    .S(_02387_),
    .X(_00320_));
 sg13g2_mux2_1 _09967_ (.A0(net3304),
    .A1(net4579),
    .S(_02387_),
    .X(_00321_));
 sg13g2_mux2_1 _09968_ (.A0(net3256),
    .A1(net4991),
    .S(_02387_),
    .X(_00322_));
 sg13g2_nand2_2 _09969_ (.Y(_02388_),
    .A(net3609),
    .B(net5187));
 sg13g2_a22oi_1 _09970_ (.Y(_02389_),
    .B1(_02388_),
    .B2(\state[2] ),
    .A2(_02190_),
    .A1(_00011_));
 sg13g2_nor2_2 _09971_ (.A(net10),
    .B(_02191_),
    .Y(_02390_));
 sg13g2_o21ai_1 _09972_ (.B1(\PC[2] ),
    .Y(_02391_),
    .A1(\PC[1] ),
    .A2(\PC[0] ));
 sg13g2_nor2_1 _09973_ (.A(_02132_),
    .B(_02391_),
    .Y(_02392_));
 sg13g2_and2_1 _09974_ (.A(\PC[4] ),
    .B(_02392_),
    .X(_02393_));
 sg13g2_and3_1 _09975_ (.X(_02394_),
    .A(\PC[6] ),
    .B(\PC[5] ),
    .C(_02393_));
 sg13g2_a21oi_1 _09976_ (.A1(\PC[7] ),
    .A2(_02394_),
    .Y(_02395_),
    .B1(_02181_));
 sg13g2_nand2b_2 _09977_ (.Y(_02396_),
    .B(_02395_),
    .A_N(net5210));
 sg13g2_a22oi_1 _09978_ (.Y(_02397_),
    .B1(_02390_),
    .B2(_02396_),
    .A2(net3063),
    .A1(_02190_));
 sg13g2_nand2_1 _09979_ (.Y(_02398_),
    .A(\state[2] ),
    .B(\state[1] ));
 sg13g2_nor2_2 _09980_ (.A(net3610),
    .B(_02398_),
    .Y(_02399_));
 sg13g2_or2_2 _09981_ (.X(_02400_),
    .B(_02398_),
    .A(net3610));
 sg13g2_nor3_1 _09982_ (.A(net3476),
    .B(net3523),
    .C(net3570),
    .Y(_02401_));
 sg13g2_nor4_1 _09983_ (.A(net3296),
    .B(net3339),
    .C(net3385),
    .D(net3431),
    .Y(_02402_));
 sg13g2_a21oi_2 _09984_ (.B1(net3247),
    .Y(_02403_),
    .A2(_02402_),
    .A1(_02401_));
 sg13g2_mux2_1 _09985_ (.A0(net5200),
    .A1(_00010_),
    .S(net3062),
    .X(_02404_));
 sg13g2_nand2_1 _09986_ (.Y(_02405_),
    .A(_02399_),
    .B(_02404_));
 sg13g2_nor2b_2 _09987_ (.A(net3609),
    .B_N(net3610),
    .Y(_02406_));
 sg13g2_and2_1 _09988_ (.A(\state[2] ),
    .B(_02406_),
    .X(_02407_));
 sg13g2_nand2_2 _09989_ (.Y(_02408_),
    .A(\state[2] ),
    .B(_02406_));
 sg13g2_nand2_1 _09990_ (.Y(_02409_),
    .A(net3609),
    .B(_00011_));
 sg13g2_and3_1 _09991_ (.X(_02410_),
    .A(net3609),
    .B(net3610),
    .C(_00011_));
 sg13g2_nand3_1 _09992_ (.B(net3610),
    .C(_00011_),
    .A(net3609),
    .Y(_02411_));
 sg13g2_nand2_2 _09993_ (.Y(_02412_),
    .A(net3059),
    .B(_02411_));
 sg13g2_nor2_1 _09994_ (.A(_02136_),
    .B(_02190_),
    .Y(_02413_));
 sg13g2_nand2_2 _09995_ (.Y(_02414_),
    .A(\state[2] ),
    .B(_02189_));
 sg13g2_a21oi_1 _09996_ (.A1(\B[0] ),
    .A2(net3057),
    .Y(_02415_),
    .B1(net3063));
 sg13g2_and3_2 _09997_ (.X(_02416_),
    .A(_00011_),
    .B(_02190_),
    .C(_02388_));
 sg13g2_nand3_1 _09998_ (.B(_02190_),
    .C(_02388_),
    .A(_00011_),
    .Y(_02417_));
 sg13g2_o21ai_1 _09999_ (.B1(_02415_),
    .Y(_02418_),
    .A1(\mem.addr[0] ),
    .A2(_02417_));
 sg13g2_a21oi_1 _10000_ (.A1(\A[0] ),
    .A2(_02412_),
    .Y(_02419_),
    .B1(_02418_));
 sg13g2_a22oi_1 _10001_ (.Y(_02420_),
    .B1(_02405_),
    .B2(_02419_),
    .A2(net3063),
    .A1(_02135_));
 sg13g2_nor2b_1 _10002_ (.A(_02420_),
    .B_N(net3019),
    .Y(_02421_));
 sg13g2_nor2_1 _10003_ (.A(net5215),
    .B(net3019),
    .Y(_02422_));
 sg13g2_nor3_1 _10004_ (.A(net3996),
    .B(_02421_),
    .C(_02422_),
    .Y(_00323_));
 sg13g2_nand2_1 _10005_ (.Y(_02423_),
    .A(_02134_),
    .B(net3063));
 sg13g2_nor2_1 _10006_ (.A(_02134_),
    .B(_02135_),
    .Y(_02424_));
 sg13g2_xnor2_1 _10007_ (.Y(_02425_),
    .A(\PC[1] ),
    .B(\PC[0] ));
 sg13g2_mux2_1 _10008_ (.A0(net5198),
    .A1(_02425_),
    .S(net3061),
    .X(_02426_));
 sg13g2_nand2_2 _10009_ (.Y(_02427_),
    .A(_02399_),
    .B(_02426_));
 sg13g2_nand2_1 _10010_ (.Y(_02428_),
    .A(_02247_),
    .B(_02296_));
 sg13g2_a21oi_1 _10011_ (.A1(\B[1] ),
    .A2(net3057),
    .Y(_02429_),
    .B1(net3063));
 sg13g2_a22oi_1 _10012_ (.Y(_02430_),
    .B1(_02416_),
    .B2(_02428_),
    .A2(_02412_),
    .A1(\A[1] ));
 sg13g2_nand3_1 _10013_ (.B(_02429_),
    .C(_02430_),
    .A(_02427_),
    .Y(_02431_));
 sg13g2_nand2b_1 _10014_ (.Y(_02432_),
    .B(net3607),
    .A_N(net3019));
 sg13g2_nand3_1 _10015_ (.B(_02423_),
    .C(_02431_),
    .A(net3018),
    .Y(_02433_));
 sg13g2_a21oi_1 _10016_ (.A1(_02432_),
    .A2(_02433_),
    .Y(_00324_),
    .B1(net3996));
 sg13g2_nand3_1 _10017_ (.B(_02134_),
    .C(_02135_),
    .A(_02133_),
    .Y(_02434_));
 sg13g2_and2_1 _10018_ (.A(_02391_),
    .B(_02434_),
    .X(_02435_));
 sg13g2_nor2_1 _10019_ (.A(net5220),
    .B(net3061),
    .Y(_02436_));
 sg13g2_a21oi_1 _10020_ (.A1(net3062),
    .A2(_02435_),
    .Y(_02437_),
    .B1(_02436_));
 sg13g2_or2_1 _10021_ (.X(_02438_),
    .B(_02437_),
    .A(_02400_));
 sg13g2_o21ai_1 _10022_ (.B1(_02416_),
    .Y(_02439_),
    .A1(net3606),
    .A2(_02303_));
 sg13g2_nor2b_1 _10023_ (.A(_02439_),
    .B_N(_02305_),
    .Y(_02440_));
 sg13g2_a221oi_1 _10024_ (.B2(\B[2] ),
    .C1(net3064),
    .B1(net3058),
    .A1(\A[2] ),
    .Y(_02441_),
    .A2(_02412_));
 sg13g2_nor2b_1 _10025_ (.A(_02440_),
    .B_N(_02441_),
    .Y(_02442_));
 sg13g2_a22oi_1 _10026_ (.Y(_02443_),
    .B1(_02438_),
    .B2(_02442_),
    .A2(net3063),
    .A1(_02133_));
 sg13g2_nand2b_1 _10027_ (.Y(_02444_),
    .B(net3606),
    .A_N(net3017));
 sg13g2_nand2_1 _10028_ (.Y(_02445_),
    .A(net3017),
    .B(_02443_));
 sg13g2_a21oi_1 _10029_ (.A1(_02444_),
    .A2(_02445_),
    .Y(_00325_),
    .B1(net3995));
 sg13g2_nand2_1 _10030_ (.Y(_02446_),
    .A(_02132_),
    .B(net3063));
 sg13g2_xnor2_1 _10031_ (.Y(_02447_),
    .A(\PC[3] ),
    .B(_02391_));
 sg13g2_nor2_1 _10032_ (.A(net5225),
    .B(net3062),
    .Y(_02448_));
 sg13g2_a21oi_1 _10033_ (.A1(net3062),
    .A2(_02447_),
    .Y(_02449_),
    .B1(_02448_));
 sg13g2_nor2_2 _10034_ (.A(_02400_),
    .B(_02449_),
    .Y(_02450_));
 sg13g2_xor2_1 _10035_ (.B(_02305_),
    .A(net3605),
    .X(_02451_));
 sg13g2_a221oi_1 _10036_ (.B2(\B[3] ),
    .C1(net3064),
    .B1(net3058),
    .A1(\A[3] ),
    .Y(_02452_),
    .A2(_02412_));
 sg13g2_o21ai_1 _10037_ (.B1(_02452_),
    .Y(_02453_),
    .A1(_02417_),
    .A2(_02451_));
 sg13g2_o21ai_1 _10038_ (.B1(_02446_),
    .Y(_02454_),
    .A1(_02450_),
    .A2(_02453_));
 sg13g2_o21ai_1 _10039_ (.B1(net4008),
    .Y(_02455_),
    .A1(net3605),
    .A2(net3017));
 sg13g2_a21oi_1 _10040_ (.A1(net3018),
    .A2(_02454_),
    .Y(_00326_),
    .B1(_02455_));
 sg13g2_xor2_1 _10041_ (.B(_02392_),
    .A(\PC[4] ),
    .X(_02456_));
 sg13g2_nor2_1 _10042_ (.A(_00015_),
    .B(net3062),
    .Y(_02457_));
 sg13g2_a21oi_1 _10043_ (.A1(net3061),
    .A2(_02456_),
    .Y(_02458_),
    .B1(_02457_));
 sg13g2_nor2_2 _10044_ (.A(_02400_),
    .B(_02458_),
    .Y(_02459_));
 sg13g2_xnor2_1 _10045_ (.Y(_02460_),
    .A(net3604),
    .B(net3076));
 sg13g2_a22oi_1 _10046_ (.Y(_02461_),
    .B1(_02412_),
    .B2(net5193),
    .A2(net3063),
    .A1(\PC[4] ));
 sg13g2_a22oi_1 _10047_ (.Y(_02462_),
    .B1(_02416_),
    .B2(_02460_),
    .A2(net3057),
    .A1(\B[4] ));
 sg13g2_nand2_1 _10048_ (.Y(_02463_),
    .A(_02461_),
    .B(_02462_));
 sg13g2_nor2_2 _10049_ (.A(_02459_),
    .B(_02463_),
    .Y(_02464_));
 sg13g2_o21ai_1 _10050_ (.B1(net4008),
    .Y(_02465_),
    .A1(net5206),
    .A2(net3019));
 sg13g2_a21oi_1 _10051_ (.A1(net3019),
    .A2(_02464_),
    .Y(_00327_),
    .B1(_02465_));
 sg13g2_xor2_1 _10052_ (.B(_02393_),
    .A(\PC[5] ),
    .X(_02466_));
 sg13g2_nor2_1 _10053_ (.A(_00014_),
    .B(net3061),
    .Y(_02467_));
 sg13g2_a21oi_1 _10054_ (.A1(net3061),
    .A2(_02466_),
    .Y(_02468_),
    .B1(_02467_));
 sg13g2_nor2_2 _10055_ (.A(_02400_),
    .B(_02468_),
    .Y(_02469_));
 sg13g2_a21oi_1 _10056_ (.A1(net3604),
    .A2(net3077),
    .Y(_02470_),
    .B1(\mem.addr[5] ));
 sg13g2_o21ai_1 _10057_ (.B1(_02416_),
    .Y(_02471_),
    .A1(net3088),
    .A2(net3076));
 sg13g2_a221oi_1 _10058_ (.B2(\B[5] ),
    .C1(net3064),
    .B1(net3058),
    .A1(\A[5] ),
    .Y(_02472_),
    .A2(_02412_));
 sg13g2_o21ai_1 _10059_ (.B1(_02472_),
    .Y(_02473_),
    .A1(_02470_),
    .A2(_02471_));
 sg13g2_nand2b_1 _10060_ (.Y(_02474_),
    .B(net3064),
    .A_N(\PC[5] ));
 sg13g2_o21ai_1 _10061_ (.B1(_02474_),
    .Y(_02475_),
    .A1(_02469_),
    .A2(_02473_));
 sg13g2_o21ai_1 _10062_ (.B1(net4008),
    .Y(_02476_),
    .A1(net5224),
    .A2(net3018));
 sg13g2_a21oi_1 _10063_ (.A1(net3017),
    .A2(_02475_),
    .Y(_00328_),
    .B1(_02476_));
 sg13g2_nand4_1 _10064_ (.B(\mem.addr[5] ),
    .C(net3604),
    .A(net3603),
    .Y(_02477_),
    .D(net3077));
 sg13g2_inv_1 _10065_ (.Y(_02478_),
    .A(_02477_));
 sg13g2_o21ai_1 _10066_ (.B1(net3017),
    .Y(_02479_),
    .A1(_02417_),
    .A2(_02478_));
 sg13g2_a21oi_1 _10067_ (.A1(\PC[5] ),
    .A2(_02393_),
    .Y(_02480_),
    .B1(\PC[6] ));
 sg13g2_o21ai_1 _10068_ (.B1(net3061),
    .Y(_02481_),
    .A1(_02394_),
    .A2(_02480_));
 sg13g2_o21ai_1 _10069_ (.B1(_02481_),
    .Y(_02482_),
    .A1(_02185_),
    .A2(net3061));
 sg13g2_nor2_1 _10070_ (.A(_02400_),
    .B(_02482_),
    .Y(_02483_));
 sg13g2_nor4_2 _10071_ (.A(net3603),
    .B(net3088),
    .C(net3076),
    .Y(_02484_),
    .D(_02417_));
 sg13g2_nand2_1 _10072_ (.Y(_02485_),
    .A(\B[6] ),
    .B(net3058));
 sg13g2_a221oi_1 _10073_ (.B2(\A[6] ),
    .C1(_02484_),
    .B1(_02412_),
    .A1(\PC[6] ),
    .Y(_02486_),
    .A2(net3064));
 sg13g2_nand3b_1 _10074_ (.B(_02485_),
    .C(_02486_),
    .Y(_02487_),
    .A_N(_02483_));
 sg13g2_a22oi_1 _10075_ (.Y(_02488_),
    .B1(_02487_),
    .B2(net3018),
    .A2(_02479_),
    .A1(net3603));
 sg13g2_nor2_1 _10076_ (.A(net3996),
    .B(_02488_),
    .Y(_00329_));
 sg13g2_xnor2_1 _10077_ (.Y(_02489_),
    .A(\PC[7] ),
    .B(_02394_));
 sg13g2_mux2_1 _10078_ (.A0(net5219),
    .A1(_02489_),
    .S(net3061),
    .X(_02490_));
 sg13g2_nand2b_1 _10079_ (.Y(_02491_),
    .B(_02399_),
    .A_N(_02490_));
 sg13g2_a21oi_1 _10080_ (.A1(\B[7] ),
    .A2(net3058),
    .Y(_02492_),
    .B1(net3064));
 sg13g2_nand3_1 _10081_ (.B(net3068),
    .C(_02416_),
    .A(net3077),
    .Y(_02493_));
 sg13g2_nand2_1 _10082_ (.Y(_02494_),
    .A(_02492_),
    .B(_02493_));
 sg13g2_a21oi_1 _10083_ (.A1(\A[7] ),
    .A2(_02412_),
    .Y(_02495_),
    .B1(_02494_));
 sg13g2_a22oi_1 _10084_ (.Y(_02496_),
    .B1(_02491_),
    .B2(_02495_),
    .A2(net3064),
    .A1(_02131_));
 sg13g2_a22oi_1 _10085_ (.Y(_02497_),
    .B1(_02496_),
    .B2(net3017),
    .A2(_02479_),
    .A1(net5226));
 sg13g2_nor2_1 _10086_ (.A(net3996),
    .B(_02497_),
    .Y(_00330_));
 sg13g2_nand2_2 _10087_ (.Y(_02498_),
    .A(net3038),
    .B(net3069));
 sg13g2_mux2_1 _10088_ (.A0(net3592),
    .A1(net5017),
    .S(_02498_),
    .X(_00331_));
 sg13g2_mux2_1 _10089_ (.A0(net3548),
    .A1(net2953),
    .S(_02498_),
    .X(_00332_));
 sg13g2_mux2_1 _10090_ (.A0(net3503),
    .A1(net4531),
    .S(_02498_),
    .X(_00333_));
 sg13g2_mux2_1 _10091_ (.A0(net3458),
    .A1(net4783),
    .S(_02498_),
    .X(_00334_));
 sg13g2_mux2_1 _10092_ (.A0(net3412),
    .A1(net4331),
    .S(_02498_),
    .X(_00335_));
 sg13g2_mux2_1 _10093_ (.A0(net3368),
    .A1(net4251),
    .S(_02498_),
    .X(_00336_));
 sg13g2_mux2_1 _10094_ (.A0(net3322),
    .A1(net5113),
    .S(_02498_),
    .X(_00337_));
 sg13g2_mux2_1 _10095_ (.A0(net3273),
    .A1(net5042),
    .S(_02498_),
    .X(_00338_));
 sg13g2_nand2_2 _10096_ (.Y(_02499_),
    .A(net3069),
    .B(_02375_));
 sg13g2_mux2_1 _10097_ (.A0(net3599),
    .A1(net4160),
    .S(_02499_),
    .X(_00339_));
 sg13g2_mux2_1 _10098_ (.A0(net3554),
    .A1(net4433),
    .S(_02499_),
    .X(_00340_));
 sg13g2_mux2_1 _10099_ (.A0(net3508),
    .A1(net5173),
    .S(_02499_),
    .X(_00341_));
 sg13g2_mux2_1 _10100_ (.A0(net3462),
    .A1(net2895),
    .S(_02499_),
    .X(_00342_));
 sg13g2_mux2_1 _10101_ (.A0(net3413),
    .A1(net4652),
    .S(_02499_),
    .X(_00343_));
 sg13g2_mux2_1 _10102_ (.A0(net3369),
    .A1(net4752),
    .S(_02499_),
    .X(_00344_));
 sg13g2_mux2_1 _10103_ (.A0(net3323),
    .A1(net4365),
    .S(_02499_),
    .X(_00345_));
 sg13g2_mux2_1 _10104_ (.A0(net3277),
    .A1(net4627),
    .S(_02499_),
    .X(_00346_));
 sg13g2_nand2_2 _10105_ (.Y(_02500_),
    .A(_02277_),
    .B(net3038));
 sg13g2_mux2_1 _10106_ (.A0(net3592),
    .A1(net4598),
    .S(_02500_),
    .X(_00347_));
 sg13g2_mux2_1 _10107_ (.A0(net3548),
    .A1(net4158),
    .S(_02500_),
    .X(_00348_));
 sg13g2_mux2_1 _10108_ (.A0(net3503),
    .A1(net4969),
    .S(_02500_),
    .X(_00349_));
 sg13g2_mux2_1 _10109_ (.A0(net3458),
    .A1(net4546),
    .S(_02500_),
    .X(_00350_));
 sg13g2_mux2_1 _10110_ (.A0(net3412),
    .A1(net2923),
    .S(_02500_),
    .X(_00351_));
 sg13g2_mux2_1 _10111_ (.A0(net3368),
    .A1(net2884),
    .S(_02500_),
    .X(_00352_));
 sg13g2_mux2_1 _10112_ (.A0(net3322),
    .A1(net2867),
    .S(_02500_),
    .X(_00353_));
 sg13g2_mux2_1 _10113_ (.A0(net3273),
    .A1(net2891),
    .S(_02500_),
    .X(_00354_));
 sg13g2_nor3_2 _10114_ (.A(_02261_),
    .B(_02278_),
    .C(_02285_),
    .Y(_02501_));
 sg13g2_mux2_1 _10115_ (.A0(net2179),
    .A1(net3599),
    .S(_02501_),
    .X(_00355_));
 sg13g2_mux2_1 _10116_ (.A0(net2809),
    .A1(net3553),
    .S(_02501_),
    .X(_00356_));
 sg13g2_mux2_1 _10117_ (.A0(net2242),
    .A1(net3504),
    .S(_02501_),
    .X(_00357_));
 sg13g2_mux2_1 _10118_ (.A0(net2437),
    .A1(net3462),
    .S(_02501_),
    .X(_00358_));
 sg13g2_mux2_1 _10119_ (.A0(net2333),
    .A1(net3415),
    .S(_02501_),
    .X(_00359_));
 sg13g2_mux2_1 _10120_ (.A0(net2184),
    .A1(net3369),
    .S(_02501_),
    .X(_00360_));
 sg13g2_mux2_1 _10121_ (.A0(net2182),
    .A1(net3323),
    .S(_02501_),
    .X(_00361_));
 sg13g2_mux2_1 _10122_ (.A0(net2410),
    .A1(net3277),
    .S(_02501_),
    .X(_00362_));
 sg13g2_nand2_2 _10123_ (.Y(_02502_),
    .A(net3037),
    .B(_02349_));
 sg13g2_mux2_1 _10124_ (.A0(net3591),
    .A1(net4680),
    .S(_02502_),
    .X(_00363_));
 sg13g2_mux2_1 _10125_ (.A0(net3547),
    .A1(net4585),
    .S(_02502_),
    .X(_00364_));
 sg13g2_mux2_1 _10126_ (.A0(net3500),
    .A1(net5122),
    .S(_02502_),
    .X(_00365_));
 sg13g2_mux2_1 _10127_ (.A0(net3455),
    .A1(net4556),
    .S(_02502_),
    .X(_00366_));
 sg13g2_mux2_1 _10128_ (.A0(net3409),
    .A1(net4467),
    .S(_02502_),
    .X(_00367_));
 sg13g2_mux2_1 _10129_ (.A0(net3365),
    .A1(net4839),
    .S(_02502_),
    .X(_00368_));
 sg13g2_mux2_1 _10130_ (.A0(net3319),
    .A1(net4138),
    .S(_02502_),
    .X(_00369_));
 sg13g2_mux2_1 _10131_ (.A0(net3270),
    .A1(net4595),
    .S(_02502_),
    .X(_00370_));
 sg13g2_nand2_2 _10132_ (.Y(_02503_),
    .A(_02284_),
    .B(net3033));
 sg13g2_mux2_1 _10133_ (.A0(net3597),
    .A1(net4872),
    .S(_02503_),
    .X(_00371_));
 sg13g2_mux2_1 _10134_ (.A0(net3552),
    .A1(net4516),
    .S(_02503_),
    .X(_00372_));
 sg13g2_mux2_1 _10135_ (.A0(net3505),
    .A1(net5009),
    .S(_02503_),
    .X(_00373_));
 sg13g2_mux2_1 _10136_ (.A0(net3461),
    .A1(net4874),
    .S(_02503_),
    .X(_00374_));
 sg13g2_mux2_1 _10137_ (.A0(net3413),
    .A1(net4313),
    .S(_02503_),
    .X(_00375_));
 sg13g2_mux2_1 _10138_ (.A0(net3369),
    .A1(net5087),
    .S(_02503_),
    .X(_00376_));
 sg13g2_mux2_1 _10139_ (.A0(net3323),
    .A1(net4260),
    .S(_02503_),
    .X(_00377_));
 sg13g2_mux2_1 _10140_ (.A0(net3277),
    .A1(net4826),
    .S(_02503_),
    .X(_00378_));
 sg13g2_nand2_2 _10141_ (.Y(_02504_),
    .A(net3049),
    .B(net3075));
 sg13g2_mux2_1 _10142_ (.A0(net3566),
    .A1(net4236),
    .S(_02504_),
    .X(_00379_));
 sg13g2_mux2_1 _10143_ (.A0(net3523),
    .A1(net4697),
    .S(_02504_),
    .X(_00380_));
 sg13g2_mux2_1 _10144_ (.A0(net3476),
    .A1(net4650),
    .S(_02504_),
    .X(_00381_));
 sg13g2_mux2_1 _10145_ (.A0(net3430),
    .A1(net5037),
    .S(_02504_),
    .X(_00382_));
 sg13g2_mux2_1 _10146_ (.A0(net3384),
    .A1(net5003),
    .S(_02504_),
    .X(_00383_));
 sg13g2_mux2_1 _10147_ (.A0(net3339),
    .A1(net4948),
    .S(_02504_),
    .X(_00384_));
 sg13g2_mux2_1 _10148_ (.A0(net3294),
    .A1(net4842),
    .S(_02504_),
    .X(_00385_));
 sg13g2_mux2_1 _10149_ (.A0(net3246),
    .A1(net5120),
    .S(_02504_),
    .X(_00386_));
 sg13g2_nand2_2 _10150_ (.Y(_02505_),
    .A(net3083),
    .B(_02328_));
 sg13g2_mux2_1 _10151_ (.A0(net3568),
    .A1(net4980),
    .S(_02505_),
    .X(_00387_));
 sg13g2_mux2_1 _10152_ (.A0(net3520),
    .A1(net4432),
    .S(_02505_),
    .X(_00388_));
 sg13g2_mux2_1 _10153_ (.A0(net3473),
    .A1(net4347),
    .S(_02505_),
    .X(_00389_));
 sg13g2_mux2_1 _10154_ (.A0(net3428),
    .A1(net4420),
    .S(_02505_),
    .X(_00390_));
 sg13g2_mux2_1 _10155_ (.A0(net3382),
    .A1(net5052),
    .S(_02505_),
    .X(_00391_));
 sg13g2_mux2_1 _10156_ (.A0(net3337),
    .A1(net5030),
    .S(_02505_),
    .X(_00392_));
 sg13g2_mux2_1 _10157_ (.A0(net3292),
    .A1(net4840),
    .S(_02505_),
    .X(_00393_));
 sg13g2_mux2_1 _10158_ (.A0(net3244),
    .A1(net4934),
    .S(_02505_),
    .X(_00394_));
 sg13g2_and2_2 _10159_ (.A(net3075),
    .B(_02385_),
    .X(_02506_));
 sg13g2_mux2_1 _10160_ (.A0(net2399),
    .A1(net3567),
    .S(_02506_),
    .X(_00395_));
 sg13g2_mux2_1 _10161_ (.A0(net2478),
    .A1(net3523),
    .S(_02506_),
    .X(_00396_));
 sg13g2_mux2_1 _10162_ (.A0(net2720),
    .A1(net3476),
    .S(_02506_),
    .X(_00397_));
 sg13g2_mux2_1 _10163_ (.A0(net2624),
    .A1(net3430),
    .S(_02506_),
    .X(_00398_));
 sg13g2_mux2_1 _10164_ (.A0(net2160),
    .A1(net3384),
    .S(_02506_),
    .X(_00399_));
 sg13g2_mux2_1 _10165_ (.A0(net2161),
    .A1(net3339),
    .S(_02506_),
    .X(_00400_));
 sg13g2_mux2_1 _10166_ (.A0(net2137),
    .A1(net3294),
    .S(_02506_),
    .X(_00401_));
 sg13g2_mux2_1 _10167_ (.A0(net2252),
    .A1(net3246),
    .S(_02506_),
    .X(_00402_));
 sg13g2_nand2_2 _10168_ (.Y(_02507_),
    .A(net3082),
    .B(_02385_));
 sg13g2_mux2_1 _10169_ (.A0(net3582),
    .A1(net4911),
    .S(_02507_),
    .X(_00403_));
 sg13g2_mux2_1 _10170_ (.A0(net3536),
    .A1(net4900),
    .S(_02507_),
    .X(_00404_));
 sg13g2_mux2_1 _10171_ (.A0(net3493),
    .A1(net4353),
    .S(_02507_),
    .X(_00405_));
 sg13g2_mux2_1 _10172_ (.A0(net3445),
    .A1(net4335),
    .S(_02507_),
    .X(_00406_));
 sg13g2_mux2_1 _10173_ (.A0(net3400),
    .A1(net2710),
    .S(_02507_),
    .X(_00407_));
 sg13g2_mux2_1 _10174_ (.A0(net3358),
    .A1(net2625),
    .S(_02507_),
    .X(_00408_));
 sg13g2_mux2_1 _10175_ (.A0(net3312),
    .A1(net2779),
    .S(_02507_),
    .X(_00409_));
 sg13g2_mux2_1 _10176_ (.A0(net3262),
    .A1(net4902),
    .S(_02507_),
    .X(_00410_));
 sg13g2_nand2_2 _10177_ (.Y(_02508_),
    .A(net3083),
    .B(_02332_));
 sg13g2_mux2_1 _10178_ (.A0(net3568),
    .A1(net4074),
    .S(_02508_),
    .X(_00411_));
 sg13g2_mux2_1 _10179_ (.A0(net3520),
    .A1(net5014),
    .S(_02508_),
    .X(_00412_));
 sg13g2_mux2_1 _10180_ (.A0(net3473),
    .A1(net4857),
    .S(_02508_),
    .X(_00413_));
 sg13g2_mux2_1 _10181_ (.A0(net3428),
    .A1(net5093),
    .S(_02508_),
    .X(_00414_));
 sg13g2_mux2_1 _10182_ (.A0(net3382),
    .A1(net4403),
    .S(_02508_),
    .X(_00415_));
 sg13g2_mux2_1 _10183_ (.A0(net3336),
    .A1(net4145),
    .S(_02508_),
    .X(_00416_));
 sg13g2_mux2_1 _10184_ (.A0(net3292),
    .A1(net2862),
    .S(_02508_),
    .X(_00417_));
 sg13g2_mux2_1 _10185_ (.A0(net3244),
    .A1(net5125),
    .S(_02508_),
    .X(_00418_));
 sg13g2_nor2_2 _10186_ (.A(net3081),
    .B(_02314_),
    .Y(_02509_));
 sg13g2_mux2_1 _10187_ (.A0(net2500),
    .A1(net3566),
    .S(_02509_),
    .X(_00419_));
 sg13g2_mux2_1 _10188_ (.A0(net2386),
    .A1(net3523),
    .S(_02509_),
    .X(_00420_));
 sg13g2_mux2_1 _10189_ (.A0(net2455),
    .A1(net3476),
    .S(_02509_),
    .X(_00421_));
 sg13g2_mux2_1 _10190_ (.A0(net2547),
    .A1(net3430),
    .S(_02509_),
    .X(_00422_));
 sg13g2_mux2_1 _10191_ (.A0(net2579),
    .A1(net3384),
    .S(_02509_),
    .X(_00423_));
 sg13g2_mux2_1 _10192_ (.A0(net2135),
    .A1(net3339),
    .S(_02509_),
    .X(_00424_));
 sg13g2_mux2_1 _10193_ (.A0(net2147),
    .A1(net3295),
    .S(_02509_),
    .X(_00425_));
 sg13g2_mux2_1 _10194_ (.A0(net2289),
    .A1(net3246),
    .S(_02509_),
    .X(_00426_));
 sg13g2_nand2_2 _10195_ (.Y(_02510_),
    .A(_02313_),
    .B(net3033));
 sg13g2_mux2_1 _10196_ (.A0(net3566),
    .A1(net5169),
    .S(_02510_),
    .X(_00427_));
 sg13g2_mux2_1 _10197_ (.A0(net3518),
    .A1(net4105),
    .S(_02510_),
    .X(_00428_));
 sg13g2_mux2_1 _10198_ (.A0(net3470),
    .A1(net4894),
    .S(_02510_),
    .X(_00429_));
 sg13g2_mux2_1 _10199_ (.A0(net3426),
    .A1(net4224),
    .S(_02510_),
    .X(_00430_));
 sg13g2_mux2_1 _10200_ (.A0(net3379),
    .A1(net4452),
    .S(_02510_),
    .X(_00431_));
 sg13g2_mux2_1 _10201_ (.A0(net3339),
    .A1(net4893),
    .S(_02510_),
    .X(_00432_));
 sg13g2_mux2_1 _10202_ (.A0(net3294),
    .A1(net4813),
    .S(_02510_),
    .X(_00433_));
 sg13g2_mux2_1 _10203_ (.A0(net3242),
    .A1(net4280),
    .S(_02510_),
    .X(_00434_));
 sg13g2_nand2_2 _10204_ (.Y(_02511_),
    .A(net3082),
    .B(_02339_));
 sg13g2_mux2_1 _10205_ (.A0(net3589),
    .A1(net4296),
    .S(_02511_),
    .X(_00435_));
 sg13g2_mux2_1 _10206_ (.A0(net3537),
    .A1(net4478),
    .S(_02511_),
    .X(_00436_));
 sg13g2_mux2_1 _10207_ (.A0(net3492),
    .A1(net4211),
    .S(_02511_),
    .X(_00437_));
 sg13g2_mux2_1 _10208_ (.A0(net3445),
    .A1(net4865),
    .S(_02511_),
    .X(_00438_));
 sg13g2_mux2_1 _10209_ (.A0(net3401),
    .A1(net5153),
    .S(_02511_),
    .X(_00439_));
 sg13g2_mux2_1 _10210_ (.A0(net3356),
    .A1(net4289),
    .S(_02511_),
    .X(_00440_));
 sg13g2_mux2_1 _10211_ (.A0(net3309),
    .A1(net4172),
    .S(_02511_),
    .X(_00441_));
 sg13g2_mux2_1 _10212_ (.A0(net3261),
    .A1(net4714),
    .S(_02511_),
    .X(_00442_));
 sg13g2_nand2_2 _10213_ (.Y(_02512_),
    .A(net3036),
    .B(_02313_));
 sg13g2_mux2_1 _10214_ (.A0(net3566),
    .A1(net4867),
    .S(_02512_),
    .X(_00443_));
 sg13g2_mux2_1 _10215_ (.A0(net3518),
    .A1(net5053),
    .S(_02512_),
    .X(_00444_));
 sg13g2_mux2_1 _10216_ (.A0(net3470),
    .A1(net5004),
    .S(_02512_),
    .X(_00445_));
 sg13g2_mux2_1 _10217_ (.A0(net3426),
    .A1(net4535),
    .S(_02512_),
    .X(_00446_));
 sg13g2_mux2_1 _10218_ (.A0(net3379),
    .A1(net4505),
    .S(_02512_),
    .X(_00447_));
 sg13g2_mux2_1 _10219_ (.A0(net3339),
    .A1(net4019),
    .S(_02512_),
    .X(_00448_));
 sg13g2_mux2_1 _10220_ (.A0(net3294),
    .A1(net2813),
    .S(_02512_),
    .X(_00449_));
 sg13g2_mux2_1 _10221_ (.A0(net3243),
    .A1(net4668),
    .S(_02512_),
    .X(_00450_));
 sg13g2_nor2_2 _10222_ (.A(_02298_),
    .B(_02314_),
    .Y(_02513_));
 sg13g2_mux2_1 _10223_ (.A0(net2296),
    .A1(net3566),
    .S(_02513_),
    .X(_00451_));
 sg13g2_mux2_1 _10224_ (.A0(net2635),
    .A1(net3517),
    .S(_02513_),
    .X(_00452_));
 sg13g2_mux2_1 _10225_ (.A0(net2454),
    .A1(net3470),
    .S(_02513_),
    .X(_00453_));
 sg13g2_mux2_1 _10226_ (.A0(net2395),
    .A1(net3425),
    .S(_02513_),
    .X(_00454_));
 sg13g2_mux2_1 _10227_ (.A0(net2678),
    .A1(net3378),
    .S(_02513_),
    .X(_00455_));
 sg13g2_mux2_1 _10228_ (.A0(net2349),
    .A1(net3334),
    .S(_02513_),
    .X(_00456_));
 sg13g2_mux2_1 _10229_ (.A0(net2758),
    .A1(net3294),
    .S(_02513_),
    .X(_00457_));
 sg13g2_mux2_1 _10230_ (.A0(net2446),
    .A1(net3243),
    .S(_02513_),
    .X(_00458_));
 sg13g2_nor2_2 _10231_ (.A(_02267_),
    .B(_02340_),
    .Y(_02514_));
 sg13g2_mux2_1 _10232_ (.A0(net2596),
    .A1(net3568),
    .S(_02514_),
    .X(_00459_));
 sg13g2_mux2_1 _10233_ (.A0(net2267),
    .A1(net3520),
    .S(_02514_),
    .X(_00460_));
 sg13g2_mux2_1 _10234_ (.A0(net2292),
    .A1(net3473),
    .S(_02514_),
    .X(_00461_));
 sg13g2_mux2_1 _10235_ (.A0(net2213),
    .A1(net3428),
    .S(_02514_),
    .X(_00462_));
 sg13g2_mux2_1 _10236_ (.A0(net2736),
    .A1(net3382),
    .S(_02514_),
    .X(_00463_));
 sg13g2_mux2_1 _10237_ (.A0(net2843),
    .A1(net3336),
    .S(_02514_),
    .X(_00464_));
 sg13g2_mux2_1 _10238_ (.A0(net2162),
    .A1(net3292),
    .S(_02514_),
    .X(_00465_));
 sg13g2_mux2_1 _10239_ (.A0(net2628),
    .A1(net3244),
    .S(_02514_),
    .X(_00466_));
 sg13g2_nand3_1 _10240_ (.B(net3079),
    .C(net3075),
    .A(net3041),
    .Y(_02515_));
 sg13g2_mux2_1 _10241_ (.A0(net3566),
    .A1(net4184),
    .S(_02515_),
    .X(_00467_));
 sg13g2_mux2_1 _10242_ (.A0(net3517),
    .A1(net4217),
    .S(_02515_),
    .X(_00468_));
 sg13g2_mux2_1 _10243_ (.A0(net3470),
    .A1(net4843),
    .S(_02515_),
    .X(_00469_));
 sg13g2_mux2_1 _10244_ (.A0(net3425),
    .A1(net4271),
    .S(_02515_),
    .X(_00470_));
 sg13g2_mux2_1 _10245_ (.A0(net3378),
    .A1(net4352),
    .S(_02515_),
    .X(_00471_));
 sg13g2_mux2_1 _10246_ (.A0(net3334),
    .A1(net2683),
    .S(_02515_),
    .X(_00472_));
 sg13g2_mux2_1 _10247_ (.A0(net3295),
    .A1(net2921),
    .S(_02515_),
    .X(_00473_));
 sg13g2_mux2_1 _10248_ (.A0(net3243),
    .A1(net4472),
    .S(_02515_),
    .X(_00474_));
 sg13g2_nor3_2 _10249_ (.A(net3039),
    .B(_02285_),
    .C(net3076),
    .Y(_02516_));
 sg13g2_mux2_1 _10250_ (.A0(net2601),
    .A1(net3598),
    .S(_02516_),
    .X(_00475_));
 sg13g2_mux2_1 _10251_ (.A0(net2251),
    .A1(net3553),
    .S(_02516_),
    .X(_00476_));
 sg13g2_mux2_1 _10252_ (.A0(net2650),
    .A1(net3509),
    .S(_02516_),
    .X(_00477_));
 sg13g2_mux2_1 _10253_ (.A0(net2426),
    .A1(net3464),
    .S(_02516_),
    .X(_00478_));
 sg13g2_mux2_1 _10254_ (.A0(net2211),
    .A1(net3419),
    .S(_02516_),
    .X(_00479_));
 sg13g2_mux2_1 _10255_ (.A0(net2299),
    .A1(net3373),
    .S(_02516_),
    .X(_00480_));
 sg13g2_mux2_1 _10256_ (.A0(net2283),
    .A1(net3327),
    .S(_02516_),
    .X(_00481_));
 sg13g2_mux2_1 _10257_ (.A0(net2257),
    .A1(net3280),
    .S(_02516_),
    .X(_00482_));
 sg13g2_nand2_2 _10258_ (.Y(_02517_),
    .A(_02266_),
    .B(net3049));
 sg13g2_mux2_1 _10259_ (.A0(net3566),
    .A1(net4221),
    .S(_02517_),
    .X(_00483_));
 sg13g2_mux2_1 _10260_ (.A0(net3524),
    .A1(net4814),
    .S(_02517_),
    .X(_00484_));
 sg13g2_mux2_1 _10261_ (.A0(net3477),
    .A1(net4745),
    .S(_02517_),
    .X(_00485_));
 sg13g2_mux2_1 _10262_ (.A0(net3430),
    .A1(net4636),
    .S(_02517_),
    .X(_00486_));
 sg13g2_mux2_1 _10263_ (.A0(net3384),
    .A1(net4569),
    .S(_02517_),
    .X(_00487_));
 sg13g2_mux2_1 _10264_ (.A0(net3340),
    .A1(net4892),
    .S(_02517_),
    .X(_00488_));
 sg13g2_mux2_1 _10265_ (.A0(net3294),
    .A1(net4587),
    .S(_02517_),
    .X(_00489_));
 sg13g2_mux2_1 _10266_ (.A0(net3246),
    .A1(net4737),
    .S(_02517_),
    .X(_00490_));
 sg13g2_nand2_1 _10267_ (.Y(_02518_),
    .A(net3085),
    .B(_02375_));
 sg13g2_mux2_1 _10268_ (.A0(net3598),
    .A1(net2791),
    .S(net3016),
    .X(_00491_));
 sg13g2_mux2_1 _10269_ (.A0(net3553),
    .A1(net5071),
    .S(net3016),
    .X(_00492_));
 sg13g2_mux2_1 _10270_ (.A0(net3508),
    .A1(net2707),
    .S(net3015),
    .X(_00493_));
 sg13g2_mux2_1 _10271_ (.A0(net3463),
    .A1(net4648),
    .S(net3015),
    .X(_00494_));
 sg13g2_mux2_1 _10272_ (.A0(net3418),
    .A1(net4185),
    .S(net3016),
    .X(_00495_));
 sg13g2_nor2_1 _10273_ (.A(net3373),
    .B(net3015),
    .Y(_02519_));
 sg13g2_a21oi_1 _10274_ (.A1(_02161_),
    .A2(net3015),
    .Y(_00496_),
    .B1(_02519_));
 sg13g2_nor2_1 _10275_ (.A(net3327),
    .B(net3015),
    .Y(_02520_));
 sg13g2_a21oi_1 _10276_ (.A1(_02165_),
    .A2(net3015),
    .Y(_00497_),
    .B1(_02520_));
 sg13g2_nor2_1 _10277_ (.A(net3279),
    .B(net3015),
    .Y(_02521_));
 sg13g2_a21oi_1 _10278_ (.A1(_02171_),
    .A2(net3015),
    .Y(_00498_),
    .B1(_02521_));
 sg13g2_nand2_2 _10279_ (.Y(_02522_),
    .A(net3074),
    .B(_02375_));
 sg13g2_mux2_1 _10280_ (.A0(net3598),
    .A1(net4299),
    .S(_02522_),
    .X(_00499_));
 sg13g2_mux2_1 _10281_ (.A0(net3553),
    .A1(net4558),
    .S(_02522_),
    .X(_00500_));
 sg13g2_mux2_1 _10282_ (.A0(net3508),
    .A1(net4482),
    .S(_02522_),
    .X(_00501_));
 sg13g2_mux2_1 _10283_ (.A0(net3463),
    .A1(net4912),
    .S(_02522_),
    .X(_00502_));
 sg13g2_mux2_1 _10284_ (.A0(net3418),
    .A1(net4091),
    .S(_02522_),
    .X(_00503_));
 sg13g2_mux2_1 _10285_ (.A0(net3372),
    .A1(net4999),
    .S(_02522_),
    .X(_00504_));
 sg13g2_mux2_1 _10286_ (.A0(net3326),
    .A1(net4360),
    .S(_02522_),
    .X(_00505_));
 sg13g2_mux2_1 _10287_ (.A0(net3279),
    .A1(net5159),
    .S(_02522_),
    .X(_00506_));
 sg13g2_nand2_2 _10288_ (.Y(_02523_),
    .A(_02266_),
    .B(_02385_));
 sg13g2_mux2_1 _10289_ (.A0(net3566),
    .A1(net4415),
    .S(_02523_),
    .X(_00507_));
 sg13g2_mux2_1 _10290_ (.A0(net3524),
    .A1(net2729),
    .S(_02523_),
    .X(_00508_));
 sg13g2_mux2_1 _10291_ (.A0(net3476),
    .A1(net4950),
    .S(_02523_),
    .X(_00509_));
 sg13g2_mux2_1 _10292_ (.A0(net3430),
    .A1(net4767),
    .S(_02523_),
    .X(_00510_));
 sg13g2_mux2_1 _10293_ (.A0(net3384),
    .A1(net2818),
    .S(_02523_),
    .X(_00511_));
 sg13g2_mux2_1 _10294_ (.A0(net3340),
    .A1(net5100),
    .S(_02523_),
    .X(_00512_));
 sg13g2_mux2_1 _10295_ (.A0(net3294),
    .A1(net4092),
    .S(_02523_),
    .X(_00513_));
 sg13g2_mux2_1 _10296_ (.A0(net3246),
    .A1(net4173),
    .S(_02523_),
    .X(_00514_));
 sg13g2_nand2_2 _10297_ (.Y(_02524_),
    .A(_02284_),
    .B(_02321_));
 sg13g2_mux2_1 _10298_ (.A0(net3600),
    .A1(net2985),
    .S(_02524_),
    .X(_00515_));
 sg13g2_mux2_1 _10299_ (.A0(net3553),
    .A1(net4231),
    .S(_02524_),
    .X(_00516_));
 sg13g2_mux2_1 _10300_ (.A0(net3508),
    .A1(net2876),
    .S(_02524_),
    .X(_00517_));
 sg13g2_mux2_1 _10301_ (.A0(net3464),
    .A1(net4240),
    .S(_02524_),
    .X(_00518_));
 sg13g2_mux2_1 _10302_ (.A0(net3418),
    .A1(net4389),
    .S(_02524_),
    .X(_00519_));
 sg13g2_mux2_1 _10303_ (.A0(net3372),
    .A1(net4500),
    .S(_02524_),
    .X(_00520_));
 sg13g2_mux2_1 _10304_ (.A0(net3326),
    .A1(net4023),
    .S(_02524_),
    .X(_00521_));
 sg13g2_mux2_1 _10305_ (.A0(net3279),
    .A1(net2733),
    .S(_02524_),
    .X(_00522_));
 sg13g2_nand2_2 _10306_ (.Y(_02525_),
    .A(net3082),
    .B(_02346_));
 sg13g2_mux2_1 _10307_ (.A0(net3582),
    .A1(net2927),
    .S(_02525_),
    .X(_00523_));
 sg13g2_mux2_1 _10308_ (.A0(net3536),
    .A1(net4755),
    .S(_02525_),
    .X(_00524_));
 sg13g2_mux2_1 _10309_ (.A0(net3493),
    .A1(net4785),
    .S(_02525_),
    .X(_00525_));
 sg13g2_mux2_1 _10310_ (.A0(net3445),
    .A1(net4937),
    .S(_02525_),
    .X(_00526_));
 sg13g2_mux2_1 _10311_ (.A0(net3400),
    .A1(net5095),
    .S(_02525_),
    .X(_00527_));
 sg13g2_mux2_1 _10312_ (.A0(net3355),
    .A1(net4951),
    .S(_02525_),
    .X(_00528_));
 sg13g2_mux2_1 _10313_ (.A0(net3310),
    .A1(net4823),
    .S(_02525_),
    .X(_00529_));
 sg13g2_mux2_1 _10314_ (.A0(net3262),
    .A1(net5007),
    .S(_02525_),
    .X(_00530_));
 sg13g2_nand2_2 _10315_ (.Y(_02526_),
    .A(net3083),
    .B(_02346_));
 sg13g2_mux2_1 _10316_ (.A0(net3567),
    .A1(net4784),
    .S(_02526_),
    .X(_00531_));
 sg13g2_mux2_1 _10317_ (.A0(net3523),
    .A1(net4242),
    .S(_02526_),
    .X(_00532_));
 sg13g2_mux2_1 _10318_ (.A0(net3476),
    .A1(net4706),
    .S(_02526_),
    .X(_00533_));
 sg13g2_mux2_1 _10319_ (.A0(net3430),
    .A1(net4909),
    .S(_02526_),
    .X(_00534_));
 sg13g2_mux2_1 _10320_ (.A0(net3384),
    .A1(net4524),
    .S(_02526_),
    .X(_00535_));
 sg13g2_mux2_1 _10321_ (.A0(net3340),
    .A1(net5138),
    .S(_02526_),
    .X(_00536_));
 sg13g2_mux2_1 _10322_ (.A0(net3296),
    .A1(net4397),
    .S(_02526_),
    .X(_00537_));
 sg13g2_mux2_1 _10323_ (.A0(net3246),
    .A1(net4547),
    .S(_02526_),
    .X(_00538_));
 sg13g2_nand2_2 _10324_ (.Y(_02527_),
    .A(_02330_),
    .B(_02375_));
 sg13g2_mux2_1 _10325_ (.A0(net3599),
    .A1(net4440),
    .S(_02527_),
    .X(_00539_));
 sg13g2_mux2_1 _10326_ (.A0(net3554),
    .A1(net4527),
    .S(_02527_),
    .X(_00540_));
 sg13g2_mux2_1 _10327_ (.A0(net3507),
    .A1(net4681),
    .S(_02527_),
    .X(_00541_));
 sg13g2_mux2_1 _10328_ (.A0(net3462),
    .A1(net2814),
    .S(_02527_),
    .X(_00542_));
 sg13g2_mux2_1 _10329_ (.A0(net3417),
    .A1(net4917),
    .S(_02527_),
    .X(_00543_));
 sg13g2_mux2_1 _10330_ (.A0(net3373),
    .A1(net4244),
    .S(_02527_),
    .X(_00544_));
 sg13g2_mux2_1 _10331_ (.A0(net3325),
    .A1(net4930),
    .S(_02527_),
    .X(_00545_));
 sg13g2_mux2_1 _10332_ (.A0(net3280),
    .A1(net4526),
    .S(_02527_),
    .X(_00546_));
 sg13g2_nand2_2 _10333_ (.Y(_02528_),
    .A(net3070),
    .B(_02375_));
 sg13g2_mux2_1 _10334_ (.A0(net3599),
    .A1(net2959),
    .S(_02528_),
    .X(_00547_));
 sg13g2_mux2_1 _10335_ (.A0(net3554),
    .A1(net4140),
    .S(_02528_),
    .X(_00548_));
 sg13g2_mux2_1 _10336_ (.A0(net3506),
    .A1(net4476),
    .S(_02528_),
    .X(_00549_));
 sg13g2_mux2_1 _10337_ (.A0(net3462),
    .A1(net4345),
    .S(_02528_),
    .X(_00550_));
 sg13g2_mux2_1 _10338_ (.A0(net3417),
    .A1(net4090),
    .S(_02528_),
    .X(_00551_));
 sg13g2_mux2_1 _10339_ (.A0(net3371),
    .A1(net4761),
    .S(_02528_),
    .X(_00552_));
 sg13g2_mux2_1 _10340_ (.A0(net3325),
    .A1(net4393),
    .S(_02528_),
    .X(_00553_));
 sg13g2_mux2_1 _10341_ (.A0(net3280),
    .A1(net4396),
    .S(_02528_),
    .X(_00554_));
 sg13g2_nor3_2 _10342_ (.A(_02261_),
    .B(_02267_),
    .C(net3081),
    .Y(_02529_));
 sg13g2_mux2_1 _10343_ (.A0(net2413),
    .A1(net3567),
    .S(_02529_),
    .X(_00555_));
 sg13g2_mux2_1 _10344_ (.A0(net2535),
    .A1(net3523),
    .S(_02529_),
    .X(_00556_));
 sg13g2_mux2_1 _10345_ (.A0(net2718),
    .A1(net3477),
    .S(_02529_),
    .X(_00557_));
 sg13g2_mux2_1 _10346_ (.A0(net2433),
    .A1(net3430),
    .S(_02529_),
    .X(_00558_));
 sg13g2_mux2_1 _10347_ (.A0(net2152),
    .A1(net3384),
    .S(_02529_),
    .X(_00559_));
 sg13g2_mux2_1 _10348_ (.A0(net2727),
    .A1(net3340),
    .S(_02529_),
    .X(_00560_));
 sg13g2_mux2_1 _10349_ (.A0(net2175),
    .A1(net3294),
    .S(_02529_),
    .X(_00561_));
 sg13g2_mux2_1 _10350_ (.A0(net2288),
    .A1(net3246),
    .S(_02529_),
    .X(_00562_));
 sg13g2_nor2_2 _10351_ (.A(_02285_),
    .B(_02340_),
    .Y(_02530_));
 sg13g2_mux2_1 _10352_ (.A0(net2201),
    .A1(net3599),
    .S(_02530_),
    .X(_00563_));
 sg13g2_mux2_1 _10353_ (.A0(net2327),
    .A1(net3554),
    .S(_02530_),
    .X(_00564_));
 sg13g2_mux2_1 _10354_ (.A0(net2595),
    .A1(net3507),
    .S(_02530_),
    .X(_00565_));
 sg13g2_mux2_1 _10355_ (.A0(net2174),
    .A1(net3462),
    .S(_02530_),
    .X(_00566_));
 sg13g2_mux2_1 _10356_ (.A0(net2442),
    .A1(net3417),
    .S(_02530_),
    .X(_00567_));
 sg13g2_mux2_1 _10357_ (.A0(net2590),
    .A1(net3371),
    .S(_02530_),
    .X(_00568_));
 sg13g2_mux2_1 _10358_ (.A0(net2282),
    .A1(net3325),
    .S(_02530_),
    .X(_00569_));
 sg13g2_mux2_1 _10359_ (.A0(net2680),
    .A1(net3280),
    .S(_02530_),
    .X(_00570_));
 sg13g2_nand2_2 _10360_ (.Y(_02531_),
    .A(_02284_),
    .B(_02310_));
 sg13g2_mux2_1 _10361_ (.A0(net3599),
    .A1(net4555),
    .S(_02531_),
    .X(_00571_));
 sg13g2_mux2_1 _10362_ (.A0(net3554),
    .A1(net4733),
    .S(_02531_),
    .X(_00572_));
 sg13g2_mux2_1 _10363_ (.A0(net3504),
    .A1(net4590),
    .S(_02531_),
    .X(_00573_));
 sg13g2_mux2_1 _10364_ (.A0(net3462),
    .A1(net4375),
    .S(_02531_),
    .X(_00574_));
 sg13g2_mux2_1 _10365_ (.A0(net3415),
    .A1(net4561),
    .S(_02531_),
    .X(_00575_));
 sg13g2_mux2_1 _10366_ (.A0(net3369),
    .A1(net4201),
    .S(_02531_),
    .X(_00576_));
 sg13g2_mux2_1 _10367_ (.A0(net3323),
    .A1(net4171),
    .S(_02531_),
    .X(_00577_));
 sg13g2_mux2_1 _10368_ (.A0(net3277),
    .A1(net4044),
    .S(_02531_),
    .X(_00578_));
 sg13g2_nand2_2 _10369_ (.Y(_02532_),
    .A(net3083),
    .B(net3033));
 sg13g2_mux2_1 _10370_ (.A0(net3565),
    .A1(net5066),
    .S(_02532_),
    .X(_00579_));
 sg13g2_mux2_1 _10371_ (.A0(net3521),
    .A1(net4330),
    .S(_02532_),
    .X(_00580_));
 sg13g2_mux2_1 _10372_ (.A0(net3473),
    .A1(net4584),
    .S(_02532_),
    .X(_00581_));
 sg13g2_mux2_1 _10373_ (.A0(net3429),
    .A1(net4861),
    .S(_02532_),
    .X(_00582_));
 sg13g2_mux2_1 _10374_ (.A0(net3381),
    .A1(net4175),
    .S(_02532_),
    .X(_00583_));
 sg13g2_mux2_1 _10375_ (.A0(net3336),
    .A1(net4093),
    .S(_02532_),
    .X(_00584_));
 sg13g2_mux2_1 _10376_ (.A0(net3291),
    .A1(net4419),
    .S(_02532_),
    .X(_00585_));
 sg13g2_mux2_1 _10377_ (.A0(net3245),
    .A1(net4887),
    .S(_02532_),
    .X(_00586_));
 sg13g2_nand2_2 _10378_ (.Y(_02533_),
    .A(_02375_),
    .B(_02383_));
 sg13g2_mux2_1 _10379_ (.A0(net3599),
    .A1(net4495),
    .S(_02533_),
    .X(_00587_));
 sg13g2_mux2_1 _10380_ (.A0(net3554),
    .A1(net2852),
    .S(_02533_),
    .X(_00588_));
 sg13g2_mux2_1 _10381_ (.A0(net3506),
    .A1(net5175),
    .S(_02533_),
    .X(_00589_));
 sg13g2_mux2_1 _10382_ (.A0(net3462),
    .A1(net4321),
    .S(_02533_),
    .X(_00590_));
 sg13g2_mux2_1 _10383_ (.A0(net3415),
    .A1(net4226),
    .S(_02533_),
    .X(_00591_));
 sg13g2_mux2_1 _10384_ (.A0(net3369),
    .A1(net4366),
    .S(_02533_),
    .X(_00592_));
 sg13g2_mux2_1 _10385_ (.A0(net3323),
    .A1(net4449),
    .S(_02533_),
    .X(_00593_));
 sg13g2_mux2_1 _10386_ (.A0(net3277),
    .A1(net2886),
    .S(_02533_),
    .X(_00594_));
 sg13g2_and2_1 _10387_ (.A(_00011_),
    .B(_02406_),
    .X(_02534_));
 sg13g2_nand2_2 _10388_ (.Y(_02535_),
    .A(_00011_),
    .B(_02406_));
 sg13g2_nor2_2 _10389_ (.A(_02257_),
    .B(_02296_),
    .Y(_02536_));
 sg13g2_nor2b_1 _10390_ (.A(net3810),
    .B_N(\mem.mem[68][0] ),
    .Y(_02537_));
 sg13g2_a21oi_1 _10391_ (.A1(net3809),
    .A2(\mem.mem[69][0] ),
    .Y(_02538_),
    .B1(_02537_));
 sg13g2_nand2b_1 _10392_ (.Y(_02539_),
    .B(\mem.mem[70][0] ),
    .A_N(net3809));
 sg13g2_a21oi_1 _10393_ (.A1(net3809),
    .A2(\mem.mem[71][0] ),
    .Y(_02540_),
    .B1(net3184));
 sg13g2_a221oi_1 _10394_ (.B2(_02540_),
    .C1(net3132),
    .B1(_02539_),
    .A1(net3184),
    .Y(_02541_),
    .A2(_02538_));
 sg13g2_nor2b_1 _10395_ (.A(net3808),
    .B_N(\mem.mem[64][0] ),
    .Y(_02542_));
 sg13g2_a21oi_1 _10396_ (.A1(net3808),
    .A2(\mem.mem[65][0] ),
    .Y(_02543_),
    .B1(_02542_));
 sg13g2_nand2b_1 _10397_ (.Y(_02544_),
    .B(\mem.mem[66][0] ),
    .A_N(net3811));
 sg13g2_a21oi_1 _10398_ (.A1(net3811),
    .A2(\mem.mem[67][0] ),
    .Y(_02545_),
    .B1(net3184));
 sg13g2_a221oi_1 _10399_ (.B2(_02545_),
    .C1(net3664),
    .B1(_02544_),
    .A1(net3184),
    .Y(_02546_),
    .A2(_02543_));
 sg13g2_nor3_1 _10400_ (.A(net3636),
    .B(_02541_),
    .C(_02546_),
    .Y(_02547_));
 sg13g2_mux4_1 _10401_ (.S0(net3800),
    .A0(\mem.mem[72][0] ),
    .A1(\mem.mem[73][0] ),
    .A2(\mem.mem[74][0] ),
    .A3(\mem.mem[75][0] ),
    .S1(net3704),
    .X(_02548_));
 sg13g2_a21oi_1 _10402_ (.A1(net3800),
    .A2(\mem.mem[79][0] ),
    .Y(_02549_),
    .B1(net3182));
 sg13g2_o21ai_1 _10403_ (.B1(_02549_),
    .Y(_02550_),
    .A1(net3800),
    .A2(_02187_));
 sg13g2_nand2b_1 _10404_ (.Y(_02551_),
    .B(\mem.mem[76][0] ),
    .A_N(net3801));
 sg13g2_a21oi_1 _10405_ (.A1(net3801),
    .A2(\mem.mem[77][0] ),
    .Y(_02552_),
    .B1(net3704));
 sg13g2_a21oi_1 _10406_ (.A1(_02551_),
    .A2(_02552_),
    .Y(_02553_),
    .B1(net3131));
 sg13g2_a221oi_1 _10407_ (.B2(_02553_),
    .C1(net3103),
    .B1(_02550_),
    .A1(net3131),
    .Y(_02554_),
    .A2(_02548_));
 sg13g2_o21ai_1 _10408_ (.B1(net3096),
    .Y(_02555_),
    .A1(_02547_),
    .A2(_02554_));
 sg13g2_nand2b_1 _10409_ (.Y(_02556_),
    .B(\mem.mem[86][0] ),
    .A_N(net3810));
 sg13g2_a21oi_1 _10410_ (.A1(net3810),
    .A2(\mem.mem[87][0] ),
    .Y(_02557_),
    .B1(net3184));
 sg13g2_nor2b_1 _10411_ (.A(net3810),
    .B_N(\mem.mem[84][0] ),
    .Y(_02558_));
 sg13g2_a21oi_1 _10412_ (.A1(net3810),
    .A2(\mem.mem[85][0] ),
    .Y(_02559_),
    .B1(_02558_));
 sg13g2_a221oi_1 _10413_ (.B2(net3184),
    .C1(net3132),
    .B1(_02559_),
    .A1(_02556_),
    .Y(_02560_),
    .A2(_02557_));
 sg13g2_nor2b_1 _10414_ (.A(net3801),
    .B_N(\mem.mem[80][0] ),
    .Y(_02561_));
 sg13g2_a21oi_1 _10415_ (.A1(net3801),
    .A2(\mem.mem[81][0] ),
    .Y(_02562_),
    .B1(_02561_));
 sg13g2_nand2b_1 _10416_ (.Y(_02563_),
    .B(\mem.mem[82][0] ),
    .A_N(net3800));
 sg13g2_a21oi_1 _10417_ (.A1(net3801),
    .A2(\mem.mem[83][0] ),
    .Y(_02564_),
    .B1(net3182));
 sg13g2_a221oi_1 _10418_ (.B2(_02564_),
    .C1(net3662),
    .B1(_02563_),
    .A1(net3182),
    .Y(_02565_),
    .A2(_02562_));
 sg13g2_nor3_1 _10419_ (.A(net3634),
    .B(_02560_),
    .C(_02565_),
    .Y(_02566_));
 sg13g2_mux4_1 _10420_ (.S0(net3804),
    .A0(\mem.mem[88][0] ),
    .A1(\mem.mem[89][0] ),
    .A2(\mem.mem[90][0] ),
    .A3(\mem.mem[91][0] ),
    .S1(net3707),
    .X(_02567_));
 sg13g2_nand2b_1 _10421_ (.Y(_02568_),
    .B(\mem.mem[92][0] ),
    .A_N(net3805));
 sg13g2_a21oi_1 _10422_ (.A1(net3805),
    .A2(\mem.mem[93][0] ),
    .Y(_02569_),
    .B1(net3707));
 sg13g2_a21oi_1 _10423_ (.A1(net3805),
    .A2(\mem.mem[95][0] ),
    .Y(_02570_),
    .B1(net3183));
 sg13g2_o21ai_1 _10424_ (.B1(_02570_),
    .Y(_02571_),
    .A1(net3805),
    .A2(_02188_));
 sg13g2_a21oi_1 _10425_ (.A1(_02568_),
    .A2(_02569_),
    .Y(_02572_),
    .B1(net3130));
 sg13g2_a221oi_1 _10426_ (.B2(_02572_),
    .C1(net3104),
    .B1(_02571_),
    .A1(net3130),
    .Y(_02573_),
    .A2(_02567_));
 sg13g2_o21ai_1 _10427_ (.B1(net3624),
    .Y(_02574_),
    .A1(_02566_),
    .A2(_02573_));
 sg13g2_nand3_1 _10428_ (.B(_02555_),
    .C(_02574_),
    .A(net3090),
    .Y(_02575_));
 sg13g2_nand2b_1 _10429_ (.Y(_02576_),
    .B(\mem.mem[102][0] ),
    .A_N(net3915));
 sg13g2_a21oi_1 _10430_ (.A1(net3915),
    .A2(\mem.mem[103][0] ),
    .Y(_02577_),
    .B1(net3216));
 sg13g2_nor2b_1 _10431_ (.A(net3919),
    .B_N(\mem.mem[100][0] ),
    .Y(_02578_));
 sg13g2_a21oi_1 _10432_ (.A1(net3919),
    .A2(\mem.mem[101][0] ),
    .Y(_02579_),
    .B1(_02578_));
 sg13g2_a221oi_1 _10433_ (.B2(net3216),
    .C1(net3158),
    .B1(_02579_),
    .A1(_02576_),
    .Y(_02580_),
    .A2(_02577_));
 sg13g2_mux4_1 _10434_ (.S0(net3903),
    .A0(\mem.mem[96][0] ),
    .A1(\mem.mem[97][0] ),
    .A2(\mem.mem[98][0] ),
    .A3(\mem.mem[99][0] ),
    .S1(net3745),
    .X(_02581_));
 sg13g2_a21oi_1 _10435_ (.A1(net3154),
    .A2(_02581_),
    .Y(_02582_),
    .B1(_02580_));
 sg13g2_nor2b_1 _10436_ (.A(net3918),
    .B_N(\mem.mem[104][0] ),
    .Y(_02583_));
 sg13g2_a21oi_1 _10437_ (.A1(net3917),
    .A2(\mem.mem[105][0] ),
    .Y(_02584_),
    .B1(_02583_));
 sg13g2_nand2b_1 _10438_ (.Y(_02585_),
    .B(\mem.mem[106][0] ),
    .A_N(net3917));
 sg13g2_a21oi_1 _10439_ (.A1(net3917),
    .A2(\mem.mem[107][0] ),
    .Y(_02586_),
    .B1(net3215));
 sg13g2_a221oi_1 _10440_ (.B2(_02586_),
    .C1(net3679),
    .B1(_02585_),
    .A1(net3215),
    .Y(_02587_),
    .A2(_02584_));
 sg13g2_nand2b_1 _10441_ (.Y(_02588_),
    .B(\mem.mem[108][0] ),
    .A_N(net3904));
 sg13g2_a21oi_1 _10442_ (.A1(net3904),
    .A2(\mem.mem[109][0] ),
    .Y(_02589_),
    .B1(net3744));
 sg13g2_mux2_1 _10443_ (.A0(\mem.mem[110][0] ),
    .A1(\mem.mem[111][0] ),
    .S(net3904),
    .X(_02590_));
 sg13g2_a21oi_1 _10444_ (.A1(_02588_),
    .A2(_02589_),
    .Y(_02591_),
    .B1(net3159));
 sg13g2_o21ai_1 _10445_ (.B1(_02591_),
    .Y(_02592_),
    .A1(net3211),
    .A2(_02590_));
 sg13g2_nor2_1 _10446_ (.A(net3113),
    .B(_02587_),
    .Y(_02593_));
 sg13g2_a22oi_1 _10447_ (.Y(_02594_),
    .B1(_02592_),
    .B2(_02593_),
    .A2(_02582_),
    .A1(net3112));
 sg13g2_nor2b_1 _10448_ (.A(net3822),
    .B_N(\mem.mem[116][0] ),
    .Y(_02595_));
 sg13g2_a21oi_1 _10449_ (.A1(net3822),
    .A2(\mem.mem[117][0] ),
    .Y(_02596_),
    .B1(_02595_));
 sg13g2_nand2b_1 _10450_ (.Y(_02597_),
    .B(\mem.mem[118][0] ),
    .A_N(net3823));
 sg13g2_a21oi_1 _10451_ (.A1(net3823),
    .A2(\mem.mem[119][0] ),
    .Y(_02598_),
    .B1(net3188));
 sg13g2_a221oi_1 _10452_ (.B2(_02598_),
    .C1(net3134),
    .B1(_02597_),
    .A1(net3188),
    .Y(_02599_),
    .A2(_02596_));
 sg13g2_mux2_1 _10453_ (.A0(\mem.mem[112][0] ),
    .A1(\mem.mem[113][0] ),
    .S(net3825),
    .X(_02600_));
 sg13g2_nor2_1 _10454_ (.A(net3714),
    .B(_02600_),
    .Y(_02601_));
 sg13g2_mux2_1 _10455_ (.A0(\mem.mem[114][0] ),
    .A1(\mem.mem[115][0] ),
    .S(net3825),
    .X(_02602_));
 sg13g2_o21ai_1 _10456_ (.B1(net3134),
    .Y(_02603_),
    .A1(net3188),
    .A2(_02602_));
 sg13g2_o21ai_1 _10457_ (.B1(net3106),
    .Y(_02604_),
    .A1(_02601_),
    .A2(_02603_));
 sg13g2_mux4_1 _10458_ (.S0(net3845),
    .A0(\mem.mem[120][0] ),
    .A1(\mem.mem[121][0] ),
    .A2(\mem.mem[122][0] ),
    .A3(\mem.mem[123][0] ),
    .S1(net3721),
    .X(_02605_));
 sg13g2_mux2_1 _10459_ (.A0(\mem.mem[126][0] ),
    .A1(\mem.mem[127][0] ),
    .S(net3844),
    .X(_02606_));
 sg13g2_nor2_1 _10460_ (.A(net3192),
    .B(_02606_),
    .Y(_02607_));
 sg13g2_mux2_1 _10461_ (.A0(\mem.mem[124][0] ),
    .A1(\mem.mem[125][0] ),
    .S(net3842),
    .X(_02608_));
 sg13g2_o21ai_1 _10462_ (.B1(net3671),
    .Y(_02609_),
    .A1(net3721),
    .A2(_02608_));
 sg13g2_a21oi_1 _10463_ (.A1(net3139),
    .A2(_02605_),
    .Y(_02610_),
    .B1(net3109));
 sg13g2_o21ai_1 _10464_ (.B1(_02610_),
    .Y(_02611_),
    .A1(_02607_),
    .A2(_02609_));
 sg13g2_o21ai_1 _10465_ (.B1(_02611_),
    .Y(_02612_),
    .A1(_02599_),
    .A2(_02604_));
 sg13g2_a21oi_1 _10466_ (.A1(net3622),
    .A2(_02612_),
    .Y(_02613_),
    .B1(_02147_));
 sg13g2_o21ai_1 _10467_ (.B1(_02613_),
    .Y(_02614_),
    .A1(net3622),
    .A2(_02594_));
 sg13g2_nand2_1 _10468_ (.Y(_02615_),
    .A(_02575_),
    .B(_02614_));
 sg13g2_nand2b_1 _10469_ (.Y(_02616_),
    .B(\mem.mem[38][0] ),
    .A_N(net3933));
 sg13g2_a21oi_1 _10470_ (.A1(net3933),
    .A2(\mem.mem[39][0] ),
    .Y(_02617_),
    .B1(net3226));
 sg13g2_nor2b_1 _10471_ (.A(net3947),
    .B_N(\mem.mem[36][0] ),
    .Y(_02618_));
 sg13g2_a21oi_1 _10472_ (.A1(net3947),
    .A2(\mem.mem[37][0] ),
    .Y(_02619_),
    .B1(_02618_));
 sg13g2_a221oi_1 _10473_ (.B2(net3226),
    .C1(net3162),
    .B1(_02619_),
    .A1(_02616_),
    .Y(_02620_),
    .A2(_02617_));
 sg13g2_mux4_1 _10474_ (.S0(net3932),
    .A0(\mem.mem[32][0] ),
    .A1(\mem.mem[33][0] ),
    .A2(\mem.mem[34][0] ),
    .A3(\mem.mem[35][0] ),
    .S1(net3753),
    .X(_02621_));
 sg13g2_a21oi_1 _10475_ (.A1(net3162),
    .A2(_02621_),
    .Y(_02622_),
    .B1(_02620_));
 sg13g2_nor2b_1 _10476_ (.A(net3951),
    .B_N(\mem.mem[40][0] ),
    .Y(_02623_));
 sg13g2_a21oi_1 _10477_ (.A1(net3951),
    .A2(\mem.mem[41][0] ),
    .Y(_02624_),
    .B1(_02623_));
 sg13g2_nand2b_1 _10478_ (.Y(_02625_),
    .B(\mem.mem[42][0] ),
    .A_N(net3950));
 sg13g2_a21oi_1 _10479_ (.A1(net3950),
    .A2(\mem.mem[43][0] ),
    .Y(_02626_),
    .B1(net3225));
 sg13g2_a221oi_1 _10480_ (.B2(_02626_),
    .C1(net3684),
    .B1(_02625_),
    .A1(net3225),
    .Y(_02627_),
    .A2(_02624_));
 sg13g2_nand2b_1 _10481_ (.Y(_02628_),
    .B(\mem.mem[44][0] ),
    .A_N(net3945));
 sg13g2_a21oi_1 _10482_ (.A1(net3945),
    .A2(\mem.mem[45][0] ),
    .Y(_02629_),
    .B1(net3757));
 sg13g2_mux2_1 _10483_ (.A0(\mem.mem[46][0] ),
    .A1(\mem.mem[47][0] ),
    .S(net3936),
    .X(_02630_));
 sg13g2_a21oi_1 _10484_ (.A1(_02628_),
    .A2(_02629_),
    .Y(_02631_),
    .B1(net3162));
 sg13g2_o21ai_1 _10485_ (.B1(_02631_),
    .Y(_02632_),
    .A1(net3226),
    .A2(_02630_));
 sg13g2_nor2_1 _10486_ (.A(net3116),
    .B(_02627_),
    .Y(_02633_));
 sg13g2_a22oi_1 _10487_ (.Y(_02634_),
    .B1(_02632_),
    .B2(_02633_),
    .A2(_02622_),
    .A1(net3116));
 sg13g2_nor2b_1 _10488_ (.A(net3976),
    .B_N(\mem.mem[52][0] ),
    .Y(_02635_));
 sg13g2_a21oi_1 _10489_ (.A1(net3976),
    .A2(\mem.mem[53][0] ),
    .Y(_02636_),
    .B1(_02635_));
 sg13g2_nand2b_1 _10490_ (.Y(_02637_),
    .B(\mem.mem[54][0] ),
    .A_N(net3976));
 sg13g2_a21oi_1 _10491_ (.A1(net3976),
    .A2(\mem.mem[55][0] ),
    .Y(_02638_),
    .B1(net3232));
 sg13g2_a221oi_1 _10492_ (.B2(_02638_),
    .C1(net3170),
    .B1(_02637_),
    .A1(net3232),
    .Y(_02639_),
    .A2(_02636_));
 sg13g2_mux4_1 _10493_ (.S0(net3957),
    .A0(\mem.mem[48][0] ),
    .A1(\mem.mem[49][0] ),
    .A2(\mem.mem[50][0] ),
    .A3(\mem.mem[51][0] ),
    .S1(net3760),
    .X(_02640_));
 sg13g2_nand2_1 _10494_ (.Y(_02641_),
    .A(net3166),
    .B(_02640_));
 sg13g2_nor2_1 _10495_ (.A(net3653),
    .B(_02639_),
    .Y(_02642_));
 sg13g2_nor2b_1 _10496_ (.A(net3978),
    .B_N(\mem.mem[56][0] ),
    .Y(_02643_));
 sg13g2_a21oi_1 _10497_ (.A1(net3978),
    .A2(\mem.mem[57][0] ),
    .Y(_02644_),
    .B1(_02643_));
 sg13g2_nand2b_1 _10498_ (.Y(_02645_),
    .B(\mem.mem[58][0] ),
    .A_N(net3975));
 sg13g2_a21oi_1 _10499_ (.A1(net3977),
    .A2(\mem.mem[59][0] ),
    .Y(_02646_),
    .B1(net3233));
 sg13g2_a221oi_1 _10500_ (.B2(_02646_),
    .C1(net3689),
    .B1(_02645_),
    .A1(net3233),
    .Y(_02647_),
    .A2(_02644_));
 sg13g2_mux2_1 _10501_ (.A0(\mem.mem[62][0] ),
    .A1(\mem.mem[63][0] ),
    .S(net3983),
    .X(_02648_));
 sg13g2_nand2b_1 _10502_ (.Y(_02649_),
    .B(\mem.mem[60][0] ),
    .A_N(net3983));
 sg13g2_a21oi_1 _10503_ (.A1(net3983),
    .A2(\mem.mem[61][0] ),
    .Y(_02650_),
    .B1(net3768));
 sg13g2_a21oi_1 _10504_ (.A1(_02649_),
    .A2(_02650_),
    .Y(_02651_),
    .B1(net3173));
 sg13g2_o21ai_1 _10505_ (.B1(_02651_),
    .Y(_02652_),
    .A1(net3234),
    .A2(_02648_));
 sg13g2_nor2_1 _10506_ (.A(net3118),
    .B(_02647_),
    .Y(_02653_));
 sg13g2_a22oi_1 _10507_ (.Y(_02654_),
    .B1(_02652_),
    .B2(_02653_),
    .A2(_02642_),
    .A1(_02641_));
 sg13g2_nor2b_1 _10508_ (.A(net3884),
    .B_N(\mem.mem[4][0] ),
    .Y(_02655_));
 sg13g2_a21oi_1 _10509_ (.A1(net3883),
    .A2(\mem.mem[5][0] ),
    .Y(_02656_),
    .B1(_02655_));
 sg13g2_nand2b_1 _10510_ (.Y(_02657_),
    .B(\mem.mem[6][0] ),
    .A_N(net3883));
 sg13g2_a21oi_1 _10511_ (.A1(net3883),
    .A2(\mem.mem[7][0] ),
    .Y(_02658_),
    .B1(net3205));
 sg13g2_a221oi_1 _10512_ (.B2(_02658_),
    .C1(net3150),
    .B1(_02657_),
    .A1(net3205),
    .Y(_02659_),
    .A2(_02656_));
 sg13g2_mux4_1 _10513_ (.S0(net3926),
    .A0(\mem.mem[0][0] ),
    .A1(\mem.mem[1][0] ),
    .A2(\mem.mem[2][0] ),
    .A3(\mem.mem[3][0] ),
    .S1(net3752),
    .X(_02660_));
 sg13g2_nand2_1 _10514_ (.Y(_02661_),
    .A(net3160),
    .B(_02660_));
 sg13g2_nor2_1 _10515_ (.A(net3650),
    .B(_02659_),
    .Y(_02662_));
 sg13g2_nor2b_1 _10516_ (.A(net3887),
    .B_N(\mem.mem[8][0] ),
    .Y(_02663_));
 sg13g2_a21oi_1 _10517_ (.A1(net3888),
    .A2(\mem.mem[9][0] ),
    .Y(_02664_),
    .B1(_02663_));
 sg13g2_nand2b_1 _10518_ (.Y(_02665_),
    .B(\mem.mem[10][0] ),
    .A_N(net3888));
 sg13g2_a21oi_1 _10519_ (.A1(net3888),
    .A2(\mem.mem[11][0] ),
    .Y(_02666_),
    .B1(net3207));
 sg13g2_a221oi_1 _10520_ (.B2(_02666_),
    .C1(net3676),
    .B1(_02665_),
    .A1(net3208),
    .Y(_02667_),
    .A2(_02664_));
 sg13g2_mux2_1 _10521_ (.A0(\mem.mem[14][0] ),
    .A1(\mem.mem[15][0] ),
    .S(net3932),
    .X(_02668_));
 sg13g2_nand2b_1 _10522_ (.Y(_02669_),
    .B(\mem.mem[12][0] ),
    .A_N(net3925));
 sg13g2_a21oi_1 _10523_ (.A1(net3925),
    .A2(\mem.mem[13][0] ),
    .Y(_02670_),
    .B1(net3752));
 sg13g2_a21oi_1 _10524_ (.A1(_02669_),
    .A2(_02670_),
    .Y(_02671_),
    .B1(net3160));
 sg13g2_o21ai_1 _10525_ (.B1(_02671_),
    .Y(_02672_),
    .A1(net3221),
    .A2(_02668_));
 sg13g2_nor2_2 _10526_ (.A(net3114),
    .B(_02667_),
    .Y(_02673_));
 sg13g2_a22oi_1 _10527_ (.Y(_02674_),
    .B1(_02672_),
    .B2(_02673_),
    .A2(_02662_),
    .A1(_02661_));
 sg13g2_nand2b_1 _10528_ (.Y(_02675_),
    .B(\mem.mem[22][0] ),
    .A_N(net3939));
 sg13g2_a21oi_1 _10529_ (.A1(net3943),
    .A2(\mem.mem[23][0] ),
    .Y(_02676_),
    .B1(net3223));
 sg13g2_nor2b_1 _10530_ (.A(net3943),
    .B_N(\mem.mem[20][0] ),
    .Y(_02677_));
 sg13g2_a21oi_1 _10531_ (.A1(net3943),
    .A2(\mem.mem[21][0] ),
    .Y(_02678_),
    .B1(_02677_));
 sg13g2_a221oi_1 _10532_ (.B2(net3223),
    .C1(net3164),
    .B1(_02678_),
    .A1(_02675_),
    .Y(_02679_),
    .A2(_02676_));
 sg13g2_nor2b_1 _10533_ (.A(net3927),
    .B_N(\mem.mem[16][0] ),
    .Y(_02680_));
 sg13g2_a21oi_1 _10534_ (.A1(net3928),
    .A2(\mem.mem[17][0] ),
    .Y(_02681_),
    .B1(_02680_));
 sg13g2_nand2b_1 _10535_ (.Y(_02682_),
    .B(\mem.mem[18][0] ),
    .A_N(net3928));
 sg13g2_a21oi_1 _10536_ (.A1(net3928),
    .A2(\mem.mem[19][0] ),
    .Y(_02683_),
    .B1(net3222));
 sg13g2_a221oi_1 _10537_ (.B2(_02683_),
    .C1(net3683),
    .B1(_02682_),
    .A1(net3222),
    .Y(_02684_),
    .A2(_02681_));
 sg13g2_nor3_2 _10538_ (.A(net3648),
    .B(_02679_),
    .C(_02684_),
    .Y(_02685_));
 sg13g2_mux4_1 _10539_ (.S0(net3948),
    .A0(\mem.mem[24][0] ),
    .A1(\mem.mem[25][0] ),
    .A2(\mem.mem[26][0] ),
    .A3(\mem.mem[27][0] ),
    .S1(net3758),
    .X(_02686_));
 sg13g2_nand2b_1 _10540_ (.Y(_02687_),
    .B(\mem.mem[28][0] ),
    .A_N(net3947));
 sg13g2_a21oi_1 _10541_ (.A1(net3947),
    .A2(\mem.mem[29][0] ),
    .Y(_02688_),
    .B1(net3757));
 sg13g2_a21oi_1 _10542_ (.A1(net3947),
    .A2(\mem.mem[31][0] ),
    .Y(_02689_),
    .B1(net3224));
 sg13g2_o21ai_1 _10543_ (.B1(_02689_),
    .Y(_02690_),
    .A1(net3947),
    .A2(_02186_));
 sg13g2_a21oi_1 _10544_ (.A1(_02687_),
    .A2(_02688_),
    .Y(_02691_),
    .B1(net3162));
 sg13g2_a221oi_1 _10545_ (.B2(_02691_),
    .C1(net3115),
    .B1(_02690_),
    .A1(net3162),
    .Y(_02692_),
    .A2(_02686_));
 sg13g2_nor2_1 _10546_ (.A(_02685_),
    .B(_02692_),
    .Y(_02693_));
 sg13g2_mux4_1 _10547_ (.S0(net3627),
    .A0(_02634_),
    .A1(_02654_),
    .A2(_02674_),
    .A3(_02693_),
    .S1(net3092),
    .X(_02694_));
 sg13g2_mux4_1 _10548_ (.S0(net3838),
    .A0(\mem.mem[160][0] ),
    .A1(\mem.mem[161][0] ),
    .A2(\mem.mem[162][0] ),
    .A3(\mem.mem[163][0] ),
    .S1(net3718),
    .X(_02695_));
 sg13g2_nand2_1 _10549_ (.Y(_02696_),
    .A(net3137),
    .B(_02695_));
 sg13g2_nand2_1 _10550_ (.Y(_02697_),
    .A(net3895),
    .B(\mem.mem[165][0] ));
 sg13g2_nand2b_1 _10551_ (.Y(_02698_),
    .B(\mem.mem[164][0] ),
    .A_N(net3895));
 sg13g2_nand3_1 _10552_ (.B(_02697_),
    .C(_02698_),
    .A(net3203),
    .Y(_02699_));
 sg13g2_nor2b_1 _10553_ (.A(net3874),
    .B_N(\mem.mem[166][0] ),
    .Y(_02700_));
 sg13g2_a21oi_1 _10554_ (.A1(net3878),
    .A2(\mem.mem[167][0] ),
    .Y(_02701_),
    .B1(_02700_));
 sg13g2_a21oi_1 _10555_ (.A1(net3734),
    .A2(_02701_),
    .Y(_02702_),
    .B1(net3149));
 sg13g2_a21oi_1 _10556_ (.A1(_02699_),
    .A2(_02702_),
    .Y(_02703_),
    .B1(net3643));
 sg13g2_mux2_1 _10557_ (.A0(\mem.mem[172][0] ),
    .A1(\mem.mem[173][0] ),
    .S(net3836),
    .X(_02704_));
 sg13g2_nor2b_1 _10558_ (.A(net3835),
    .B_N(\mem.mem[174][0] ),
    .Y(_02705_));
 sg13g2_a21oi_1 _10559_ (.A1(net3835),
    .A2(\mem.mem[175][0] ),
    .Y(_02706_),
    .B1(_02705_));
 sg13g2_a21oi_1 _10560_ (.A1(net3718),
    .A2(_02706_),
    .Y(_02707_),
    .B1(net3137));
 sg13g2_o21ai_1 _10561_ (.B1(_02707_),
    .Y(_02708_),
    .A1(net3718),
    .A2(_02704_));
 sg13g2_nand2_1 _10562_ (.Y(_02709_),
    .A(net3851),
    .B(\mem.mem[169][0] ));
 sg13g2_nand2b_1 _10563_ (.Y(_02710_),
    .B(\mem.mem[168][0] ),
    .A_N(net3851));
 sg13g2_nand3_1 _10564_ (.B(_02709_),
    .C(_02710_),
    .A(net3196),
    .Y(_02711_));
 sg13g2_nor2b_1 _10565_ (.A(net3852),
    .B_N(\mem.mem[170][0] ),
    .Y(_02712_));
 sg13g2_a21oi_1 _10566_ (.A1(net3852),
    .A2(\mem.mem[171][0] ),
    .Y(_02713_),
    .B1(_02712_));
 sg13g2_a21oi_1 _10567_ (.A1(net3726),
    .A2(_02713_),
    .Y(_02714_),
    .B1(net3672));
 sg13g2_a21oi_2 _10568_ (.B1(net3110),
    .Y(_02715_),
    .A2(_02714_),
    .A1(_02711_));
 sg13g2_a221oi_1 _10569_ (.B2(_02715_),
    .C1(net3625),
    .B1(_02708_),
    .A1(_02696_),
    .Y(_02716_),
    .A2(_02703_));
 sg13g2_nor2b_1 _10570_ (.A(net3854),
    .B_N(\mem.mem[182][0] ),
    .Y(_02717_));
 sg13g2_a21oi_1 _10571_ (.A1(net3854),
    .A2(\mem.mem[183][0] ),
    .Y(_02718_),
    .B1(_02717_));
 sg13g2_mux2_1 _10572_ (.A0(\mem.mem[180][0] ),
    .A1(\mem.mem[181][0] ),
    .S(net3860),
    .X(_02719_));
 sg13g2_a21oi_1 _10573_ (.A1(net3727),
    .A2(_02718_),
    .Y(_02720_),
    .B1(net3141));
 sg13g2_o21ai_1 _10574_ (.B1(_02720_),
    .Y(_02721_),
    .A1(net3727),
    .A2(_02719_));
 sg13g2_nand2_1 _10575_ (.Y(_02722_),
    .A(net3849),
    .B(\mem.mem[177][0] ));
 sg13g2_nand2b_1 _10576_ (.Y(_02723_),
    .B(\mem.mem[176][0] ),
    .A_N(net3850));
 sg13g2_nand3_1 _10577_ (.B(_02722_),
    .C(_02723_),
    .A(net3196),
    .Y(_02724_));
 sg13g2_nor2b_1 _10578_ (.A(net3850),
    .B_N(\mem.mem[178][0] ),
    .Y(_02725_));
 sg13g2_a21oi_1 _10579_ (.A1(net3850),
    .A2(\mem.mem[179][0] ),
    .Y(_02726_),
    .B1(_02725_));
 sg13g2_a21oi_1 _10580_ (.A1(net3725),
    .A2(_02726_),
    .Y(_02727_),
    .B1(net3672));
 sg13g2_a21oi_1 _10581_ (.A1(_02724_),
    .A2(_02727_),
    .Y(_02728_),
    .B1(net3640));
 sg13g2_mux2_1 _10582_ (.A0(\mem.mem[184][0] ),
    .A1(\mem.mem[185][0] ),
    .S(net3857),
    .X(_02729_));
 sg13g2_nor2_1 _10583_ (.A(net3727),
    .B(_02729_),
    .Y(_02730_));
 sg13g2_mux2_1 _10584_ (.A0(\mem.mem[186][0] ),
    .A1(\mem.mem[187][0] ),
    .S(net3857),
    .X(_02731_));
 sg13g2_o21ai_1 _10585_ (.B1(net3141),
    .Y(_02732_),
    .A1(net3194),
    .A2(_02731_));
 sg13g2_nor2b_1 _10586_ (.A(net3856),
    .B_N(\mem.mem[188][0] ),
    .Y(_02733_));
 sg13g2_a21oi_1 _10587_ (.A1(net3856),
    .A2(\mem.mem[189][0] ),
    .Y(_02734_),
    .B1(_02733_));
 sg13g2_nand2b_1 _10588_ (.Y(_02735_),
    .B(\mem.mem[190][0] ),
    .A_N(net3856));
 sg13g2_a21oi_1 _10589_ (.A1(net3856),
    .A2(\mem.mem[191][0] ),
    .Y(_02736_),
    .B1(net3193));
 sg13g2_a221oi_1 _10590_ (.B2(_02736_),
    .C1(net3140),
    .B1(_02735_),
    .A1(net3193),
    .Y(_02737_),
    .A2(_02734_));
 sg13g2_o21ai_1 _10591_ (.B1(net3641),
    .Y(_02738_),
    .A1(_02730_),
    .A2(_02732_));
 sg13g2_o21ai_1 _10592_ (.B1(net3622),
    .Y(_02739_),
    .A1(_02737_),
    .A2(_02738_));
 sg13g2_a21oi_2 _10593_ (.B1(_02739_),
    .Y(_02740_),
    .A2(_02728_),
    .A1(_02721_));
 sg13g2_o21ai_1 _10594_ (.B1(net3616),
    .Y(_02741_),
    .A1(_02716_),
    .A2(_02740_));
 sg13g2_mux4_1 _10595_ (.S0(net3910),
    .A0(\mem.mem[128][0] ),
    .A1(\mem.mem[129][0] ),
    .A2(\mem.mem[130][0] ),
    .A3(\mem.mem[131][0] ),
    .S1(net3746),
    .X(_02742_));
 sg13g2_nand2_1 _10596_ (.Y(_02743_),
    .A(net3155),
    .B(_02742_));
 sg13g2_nand2_1 _10597_ (.Y(_02744_),
    .A(net3912),
    .B(\mem.mem[133][0] ));
 sg13g2_nand2b_1 _10598_ (.Y(_02745_),
    .B(\mem.mem[132][0] ),
    .A_N(net3912));
 sg13g2_nand3_1 _10599_ (.B(_02744_),
    .C(_02745_),
    .A(net3228),
    .Y(_02746_));
 sg13g2_nor2b_1 _10600_ (.A(net3912),
    .B_N(\mem.mem[134][0] ),
    .Y(_02747_));
 sg13g2_a21oi_1 _10601_ (.A1(net3912),
    .A2(\mem.mem[135][0] ),
    .Y(_02748_),
    .B1(_02747_));
 sg13g2_a21oi_1 _10602_ (.A1(net3747),
    .A2(_02748_),
    .Y(_02749_),
    .B1(net3157));
 sg13g2_a21oi_1 _10603_ (.A1(_02746_),
    .A2(_02749_),
    .Y(_02750_),
    .B1(net3652));
 sg13g2_mux2_1 _10604_ (.A0(\mem.mem[140][0] ),
    .A1(\mem.mem[141][0] ),
    .S(net3909),
    .X(_02751_));
 sg13g2_nor2b_1 _10605_ (.A(net3910),
    .B_N(\mem.mem[142][0] ),
    .Y(_02752_));
 sg13g2_a21oi_1 _10606_ (.A1(net3910),
    .A2(\mem.mem[143][0] ),
    .Y(_02753_),
    .B1(_02752_));
 sg13g2_a21oi_1 _10607_ (.A1(net3746),
    .A2(_02753_),
    .Y(_02754_),
    .B1(net3155));
 sg13g2_o21ai_1 _10608_ (.B1(_02754_),
    .Y(_02755_),
    .A1(net3746),
    .A2(_02751_));
 sg13g2_nand2_1 _10609_ (.Y(_02756_),
    .A(net3897),
    .B(\mem.mem[137][0] ));
 sg13g2_nand2b_1 _10610_ (.Y(_02757_),
    .B(\mem.mem[136][0] ),
    .A_N(net3897));
 sg13g2_nand3_1 _10611_ (.B(_02756_),
    .C(_02757_),
    .A(net3209),
    .Y(_02758_));
 sg13g2_nor2b_1 _10612_ (.A(net3897),
    .B_N(\mem.mem[138][0] ),
    .Y(_02759_));
 sg13g2_a21oi_1 _10613_ (.A1(net3897),
    .A2(\mem.mem[139][0] ),
    .Y(_02760_),
    .B1(_02759_));
 sg13g2_a21oi_1 _10614_ (.A1(net3742),
    .A2(_02760_),
    .Y(_02761_),
    .B1(net3677));
 sg13g2_a21oi_1 _10615_ (.A1(_02758_),
    .A2(_02761_),
    .Y(_02762_),
    .B1(net3112));
 sg13g2_a221oi_1 _10616_ (.B2(_02762_),
    .C1(net3631),
    .B1(_02755_),
    .A1(_02743_),
    .Y(_02763_),
    .A2(_02750_));
 sg13g2_mux4_1 _10617_ (.S0(net3967),
    .A0(\mem.mem[144][0] ),
    .A1(\mem.mem[145][0] ),
    .A2(\mem.mem[146][0] ),
    .A3(\mem.mem[147][0] ),
    .S1(net3762),
    .X(_02764_));
 sg13g2_nand2_1 _10618_ (.Y(_02765_),
    .A(net3968),
    .B(\mem.mem[149][0] ));
 sg13g2_nand2b_1 _10619_ (.Y(_02766_),
    .B(\mem.mem[148][0] ),
    .A_N(net3968));
 sg13g2_nand3_1 _10620_ (.B(_02765_),
    .C(_02766_),
    .A(net3234),
    .Y(_02767_));
 sg13g2_nor2b_1 _10621_ (.A(net3968),
    .B_N(\mem.mem[150][0] ),
    .Y(_02768_));
 sg13g2_a21oi_1 _10622_ (.A1(net3968),
    .A2(\mem.mem[151][0] ),
    .Y(_02769_),
    .B1(_02768_));
 sg13g2_a21oi_1 _10623_ (.A1(net3764),
    .A2(_02769_),
    .Y(_02770_),
    .B1(net3167));
 sg13g2_a221oi_1 _10624_ (.B2(_02770_),
    .C1(net3651),
    .B1(_02767_),
    .A1(net3167),
    .Y(_02771_),
    .A2(_02764_));
 sg13g2_nand2b_1 _10625_ (.Y(_02772_),
    .B(\mem.mem[158][0] ),
    .A_N(net3969));
 sg13g2_a21oi_1 _10626_ (.A1(net3969),
    .A2(\mem.mem[159][0] ),
    .Y(_02773_),
    .B1(net3231));
 sg13g2_nor2b_1 _10627_ (.A(net3969),
    .B_N(\mem.mem[156][0] ),
    .Y(_02774_));
 sg13g2_a21oi_1 _10628_ (.A1(net3969),
    .A2(\mem.mem[157][0] ),
    .Y(_02775_),
    .B1(_02774_));
 sg13g2_a221oi_1 _10629_ (.B2(net3231),
    .C1(net3167),
    .B1(_02775_),
    .A1(_02772_),
    .Y(_02776_),
    .A2(_02773_));
 sg13g2_mux4_1 _10630_ (.S0(net3986),
    .A0(\mem.mem[152][0] ),
    .A1(\mem.mem[153][0] ),
    .A2(\mem.mem[154][0] ),
    .A3(\mem.mem[155][0] ),
    .S1(net3769),
    .X(_02777_));
 sg13g2_a21o_1 _10631_ (.A2(_02777_),
    .A1(net3172),
    .B1(net3119),
    .X(_02778_));
 sg13g2_o21ai_1 _10632_ (.B1(net3629),
    .Y(_02779_),
    .A1(_02776_),
    .A2(_02778_));
 sg13g2_nor2_2 _10633_ (.A(_02771_),
    .B(_02779_),
    .Y(_02780_));
 sg13g2_o21ai_1 _10634_ (.B1(net3093),
    .Y(_02781_),
    .A1(_02763_),
    .A2(_02780_));
 sg13g2_nand2b_1 _10635_ (.Y(_02782_),
    .B(net3783),
    .A_N(\mem.mem[197][0] ));
 sg13g2_o21ai_1 _10636_ (.B1(_02782_),
    .Y(_02783_),
    .A1(net3774),
    .A2(\mem.mem[196][0] ));
 sg13g2_nand2b_1 _10637_ (.Y(_02784_),
    .B(\mem.mem[198][0] ),
    .A_N(net3775));
 sg13g2_a21oi_1 _10638_ (.A1(net3775),
    .A2(\mem.mem[199][0] ),
    .Y(_02785_),
    .B1(net3176));
 sg13g2_a221oi_1 _10639_ (.B2(_02785_),
    .C1(net3122),
    .B1(_02784_),
    .A1(net3176),
    .Y(_02786_),
    .A2(_02783_));
 sg13g2_mux4_1 _10640_ (.S0(net3775),
    .A0(\mem.mem[192][0] ),
    .A1(\mem.mem[193][0] ),
    .A2(\mem.mem[194][0] ),
    .A3(\mem.mem[195][0] ),
    .S1(net3692),
    .X(_02787_));
 sg13g2_a21oi_2 _10641_ (.B1(_02786_),
    .Y(_02788_),
    .A2(_02787_),
    .A1(net3122));
 sg13g2_mux4_1 _10642_ (.S0(net3782),
    .A0(\mem.mem[200][0] ),
    .A1(\mem.mem[201][0] ),
    .A2(\mem.mem[202][0] ),
    .A3(\mem.mem[203][0] ),
    .S1(net3701),
    .X(_02789_));
 sg13g2_nand2_1 _10643_ (.Y(_02790_),
    .A(net3122),
    .B(_02789_));
 sg13g2_nand2b_1 _10644_ (.Y(_02791_),
    .B(\mem.mem[206][0] ),
    .A_N(net3779));
 sg13g2_a21oi_1 _10645_ (.A1(net3779),
    .A2(\mem.mem[207][0] ),
    .Y(_02792_),
    .B1(net3177));
 sg13g2_nor2b_1 _10646_ (.A(net3779),
    .B_N(\mem.mem[204][0] ),
    .Y(_02793_));
 sg13g2_a21oi_1 _10647_ (.A1(net3779),
    .A2(\mem.mem[205][0] ),
    .Y(_02794_),
    .B1(_02793_));
 sg13g2_a221oi_1 _10648_ (.B2(net3177),
    .C1(net3123),
    .B1(_02794_),
    .A1(_02791_),
    .Y(_02795_),
    .A2(_02792_));
 sg13g2_mux4_1 _10649_ (.S0(net3790),
    .A0(\mem.mem[212][0] ),
    .A1(\mem.mem[213][0] ),
    .A2(\mem.mem[214][0] ),
    .A3(\mem.mem[215][0] ),
    .S1(net3698),
    .X(_02796_));
 sg13g2_nor2b_1 _10650_ (.A(net3783),
    .B_N(\mem.mem[210][0] ),
    .Y(_02797_));
 sg13g2_a21oi_1 _10651_ (.A1(net3784),
    .A2(\mem.mem[211][0] ),
    .Y(_02798_),
    .B1(_02797_));
 sg13g2_nand2_1 _10652_ (.Y(_02799_),
    .A(net3785),
    .B(\mem.mem[209][0] ));
 sg13g2_nand2b_1 _10653_ (.Y(_02800_),
    .B(\mem.mem[208][0] ),
    .A_N(net3784));
 sg13g2_nand3_1 _10654_ (.B(_02799_),
    .C(_02800_),
    .A(net3178),
    .Y(_02801_));
 sg13g2_a21oi_1 _10655_ (.A1(net3697),
    .A2(_02798_),
    .Y(_02802_),
    .B1(net3659));
 sg13g2_mux4_1 _10656_ (.S0(net3788),
    .A0(\mem.mem[216][0] ),
    .A1(\mem.mem[217][0] ),
    .A2(\mem.mem[218][0] ),
    .A3(\mem.mem[219][0] ),
    .S1(net3696),
    .X(_02803_));
 sg13g2_nor2_1 _10657_ (.A(net3101),
    .B(_02795_),
    .Y(_02804_));
 sg13g2_a221oi_1 _10658_ (.B2(_02804_),
    .C1(net3620),
    .B1(_02790_),
    .A1(net3101),
    .Y(_02805_),
    .A2(_02788_));
 sg13g2_a221oi_1 _10659_ (.B2(_02802_),
    .C1(net3637),
    .B1(_02801_),
    .A1(net3659),
    .Y(_02806_),
    .A2(_02796_));
 sg13g2_nand2b_1 _10660_ (.Y(_02807_),
    .B(\mem.mem[222][0] ),
    .A_N(net3788));
 sg13g2_a21oi_1 _10661_ (.A1(net3789),
    .A2(\mem.mem[223][0] ),
    .Y(_02808_),
    .B1(net3180));
 sg13g2_nor2b_1 _10662_ (.A(net3787),
    .B_N(\mem.mem[220][0] ),
    .Y(_02809_));
 sg13g2_a21oi_1 _10663_ (.A1(net3789),
    .A2(\mem.mem[221][0] ),
    .Y(_02810_),
    .B1(_02809_));
 sg13g2_a221oi_1 _10664_ (.B2(net3180),
    .C1(net3126),
    .B1(_02810_),
    .A1(_02807_),
    .Y(_02811_),
    .A2(_02808_));
 sg13g2_a21o_1 _10665_ (.A2(_02803_),
    .A1(net3126),
    .B1(net3102),
    .X(_02812_));
 sg13g2_o21ai_1 _10666_ (.B1(net3620),
    .Y(_02813_),
    .A1(_02811_),
    .A2(_02812_));
 sg13g2_nor2_1 _10667_ (.A(_02806_),
    .B(_02813_),
    .Y(_02814_));
 sg13g2_o21ai_1 _10668_ (.B1(net3090),
    .Y(_02815_),
    .A1(_02805_),
    .A2(_02814_));
 sg13g2_mux2_1 _10669_ (.A0(\mem.mem[236][0] ),
    .A1(\mem.mem[237][0] ),
    .S(net3831),
    .X(_02816_));
 sg13g2_nor2b_1 _10670_ (.A(\mem.mem[239][0] ),
    .B_N(net3831),
    .Y(_02817_));
 sg13g2_o21ai_1 _10671_ (.B1(net3716),
    .Y(_02818_),
    .A1(net3830),
    .A2(\mem.mem[238][0] ));
 sg13g2_o21ai_1 _10672_ (.B1(net3668),
    .Y(_02819_),
    .A1(_02817_),
    .A2(_02818_));
 sg13g2_a21oi_1 _10673_ (.A1(net3190),
    .A2(_02816_),
    .Y(_02820_),
    .B1(_02819_));
 sg13g2_mux4_1 _10674_ (.S0(net3832),
    .A0(\mem.mem[232][0] ),
    .A1(\mem.mem[233][0] ),
    .A2(\mem.mem[234][0] ),
    .A3(\mem.mem[235][0] ),
    .S1(net3716),
    .X(_02821_));
 sg13g2_o21ai_1 _10675_ (.B1(net3639),
    .Y(_02822_),
    .A1(net3669),
    .A2(_02821_));
 sg13g2_nand2b_1 _10676_ (.Y(_02823_),
    .B(net3869),
    .A_N(\mem.mem[231][0] ));
 sg13g2_o21ai_1 _10677_ (.B1(_02823_),
    .Y(_02824_),
    .A1(net3869),
    .A2(\mem.mem[230][0] ));
 sg13g2_mux2_1 _10678_ (.A0(\mem.mem[228][0] ),
    .A1(\mem.mem[229][0] ),
    .S(net3880),
    .X(_02825_));
 sg13g2_a21oi_1 _10679_ (.A1(net3205),
    .A2(_02825_),
    .Y(_02826_),
    .B1(net3147));
 sg13g2_o21ai_1 _10680_ (.B1(_02826_),
    .Y(_02827_),
    .A1(net3205),
    .A2(_02824_));
 sg13g2_mux2_1 _10681_ (.A0(\mem.mem[226][0] ),
    .A1(\mem.mem[227][0] ),
    .S(net3879),
    .X(_02828_));
 sg13g2_nand2_1 _10682_ (.Y(_02829_),
    .A(net3732),
    .B(_02828_));
 sg13g2_mux2_1 _10683_ (.A0(\mem.mem[224][0] ),
    .A1(\mem.mem[225][0] ),
    .S(net3870),
    .X(_02830_));
 sg13g2_a21oi_1 _10684_ (.A1(net3205),
    .A2(_02830_),
    .Y(_02831_),
    .B1(net3681));
 sg13g2_a21oi_1 _10685_ (.A1(_02829_),
    .A2(_02831_),
    .Y(_02832_),
    .B1(net3644));
 sg13g2_a21oi_2 _10686_ (.B1(net3625),
    .Y(_02833_),
    .A2(_02832_),
    .A1(_02827_));
 sg13g2_o21ai_1 _10687_ (.B1(_02833_),
    .Y(_02834_),
    .A1(_02820_),
    .A2(_02822_));
 sg13g2_mux4_1 _10688_ (.S0(net3819),
    .A0(\mem.mem[240][0] ),
    .A1(\mem.mem[241][0] ),
    .A2(\mem.mem[242][0] ),
    .A3(\mem.mem[243][0] ),
    .S1(net3713),
    .X(_02835_));
 sg13g2_mux4_1 _10689_ (.S0(net3819),
    .A0(\mem.mem[244][0] ),
    .A1(\mem.mem[245][0] ),
    .A2(\mem.mem[246][0] ),
    .A3(\mem.mem[247][0] ),
    .S1(net3713),
    .X(_02836_));
 sg13g2_mux2_1 _10690_ (.A0(_02835_),
    .A1(_02836_),
    .S(net3667),
    .X(_02837_));
 sg13g2_mux4_1 _10691_ (.S0(net3818),
    .A0(\mem.mem[248][0] ),
    .A1(\mem.mem[249][0] ),
    .A2(\mem.mem[250][0] ),
    .A3(\mem.mem[251][0] ),
    .S1(net3712),
    .X(_02838_));
 sg13g2_nor2_1 _10692_ (.A(net3667),
    .B(_02838_),
    .Y(_02839_));
 sg13g2_o21ai_1 _10693_ (.B1(net3638),
    .Y(_02840_),
    .A1(net3133),
    .A2(\mem.mem[252][0] ));
 sg13g2_a21oi_1 _10694_ (.A1(net3106),
    .A2(_02837_),
    .Y(_02841_),
    .B1(net3095));
 sg13g2_o21ai_1 _10695_ (.B1(_02841_),
    .Y(_02842_),
    .A1(_02839_),
    .A2(_02840_));
 sg13g2_nand3_1 _10696_ (.B(_02834_),
    .C(_02842_),
    .A(net3615),
    .Y(_02843_));
 sg13g2_nand2_1 _10697_ (.Y(_02844_),
    .A(_02741_),
    .B(_02781_));
 sg13g2_nand2_2 _10698_ (.Y(_02845_),
    .A(_02815_),
    .B(_02843_));
 sg13g2_mux4_1 _10699_ (.S0(net3089),
    .A0(_02615_),
    .A1(_02694_),
    .A2(_02845_),
    .A3(_02844_),
    .S1(net3611),
    .X(_02846_));
 sg13g2_a22oi_1 _10700_ (.Y(_02847_),
    .B1(_02846_),
    .B2(_02259_),
    .A2(_02536_),
    .A1(net1));
 sg13g2_o21ai_1 _10701_ (.B1(net4006),
    .Y(_02848_),
    .A1(net5182),
    .A2(net3055));
 sg13g2_a21oi_1 _10702_ (.A1(net3055),
    .A2(_02847_),
    .Y(_00595_),
    .B1(_02848_));
 sg13g2_mux4_1 _10703_ (.S0(net3887),
    .A0(\mem.mem[8][1] ),
    .A1(\mem.mem[9][1] ),
    .A2(\mem.mem[10][1] ),
    .A3(\mem.mem[11][1] ),
    .S1(net3740),
    .X(_02849_));
 sg13g2_nand2b_1 _10704_ (.Y(_02850_),
    .B(\mem.mem[12][1] ),
    .A_N(net3883));
 sg13g2_nand2_1 _10705_ (.Y(_02851_),
    .A(net3883),
    .B(\mem.mem[13][1] ));
 sg13g2_nand3_1 _10706_ (.B(_02850_),
    .C(_02851_),
    .A(net3206),
    .Y(_02852_));
 sg13g2_nor2b_1 _10707_ (.A(net3889),
    .B_N(\mem.mem[14][1] ),
    .Y(_02853_));
 sg13g2_a21oi_1 _10708_ (.A1(net3889),
    .A2(\mem.mem[15][1] ),
    .Y(_02854_),
    .B1(_02853_));
 sg13g2_a21oi_1 _10709_ (.A1(net3741),
    .A2(_02854_),
    .Y(_02855_),
    .B1(net3150));
 sg13g2_a221oi_1 _10710_ (.B2(_02855_),
    .C1(net3111),
    .B1(_02852_),
    .A1(net3150),
    .Y(_02856_),
    .A2(_02849_));
 sg13g2_mux4_1 _10711_ (.S0(net3925),
    .A0(\mem.mem[0][1] ),
    .A1(\mem.mem[1][1] ),
    .A2(\mem.mem[2][1] ),
    .A3(\mem.mem[3][1] ),
    .S1(net3752),
    .X(_02857_));
 sg13g2_nand2_1 _10712_ (.Y(_02858_),
    .A(net3884),
    .B(\mem.mem[7][1] ));
 sg13g2_nand2b_1 _10713_ (.Y(_02859_),
    .B(\mem.mem[6][1] ),
    .A_N(net3879));
 sg13g2_nand3_1 _10714_ (.B(_02858_),
    .C(_02859_),
    .A(net3738),
    .Y(_02860_));
 sg13g2_nand2b_1 _10715_ (.Y(_02861_),
    .B(\mem.mem[4][1] ),
    .A_N(net3882));
 sg13g2_a21oi_1 _10716_ (.A1(net3882),
    .A2(\mem.mem[5][1] ),
    .Y(_02862_),
    .B1(net3738));
 sg13g2_a21oi_1 _10717_ (.A1(_02861_),
    .A2(_02862_),
    .Y(_02863_),
    .B1(net3150));
 sg13g2_a221oi_1 _10718_ (.B2(_02863_),
    .C1(net3644),
    .B1(_02860_),
    .A1(net3151),
    .Y(_02864_),
    .A2(_02857_));
 sg13g2_or3_1 _10719_ (.A(net3628),
    .B(_02856_),
    .C(_02864_),
    .X(_02865_));
 sg13g2_mux4_1 _10720_ (.S0(net3943),
    .A0(\mem.mem[24][1] ),
    .A1(\mem.mem[25][1] ),
    .A2(\mem.mem[26][1] ),
    .A3(\mem.mem[27][1] ),
    .S1(net3756),
    .X(_02866_));
 sg13g2_mux4_1 _10721_ (.S0(net3929),
    .A0(\mem.mem[28][1] ),
    .A1(\mem.mem[29][1] ),
    .A2(\mem.mem[30][1] ),
    .A3(\mem.mem[31][1] ),
    .S1(net3754),
    .X(_02867_));
 sg13g2_nand2_1 _10722_ (.Y(_02868_),
    .A(net3682),
    .B(_02867_));
 sg13g2_a21oi_1 _10723_ (.A1(net3164),
    .A2(_02866_),
    .Y(_02869_),
    .B1(net3115));
 sg13g2_mux2_1 _10724_ (.A0(\mem.mem[18][1] ),
    .A1(\mem.mem[19][1] ),
    .S(net3929),
    .X(_02870_));
 sg13g2_mux2_1 _10725_ (.A0(\mem.mem[16][1] ),
    .A1(\mem.mem[17][1] ),
    .S(net3929),
    .X(_02871_));
 sg13g2_nor2_1 _10726_ (.A(net3751),
    .B(_02871_),
    .Y(_02872_));
 sg13g2_o21ai_1 _10727_ (.B1(net3160),
    .Y(_02873_),
    .A1(net3221),
    .A2(_02870_));
 sg13g2_nand2b_1 _10728_ (.Y(_02874_),
    .B(\mem.mem[22][1] ),
    .A_N(net3940));
 sg13g2_a21oi_1 _10729_ (.A1(net3940),
    .A2(\mem.mem[23][1] ),
    .Y(_02875_),
    .B1(net3222));
 sg13g2_nand2b_1 _10730_ (.Y(_02876_),
    .B(net3940),
    .A_N(\mem.mem[21][1] ));
 sg13g2_o21ai_1 _10731_ (.B1(_02876_),
    .Y(_02877_),
    .A1(net3940),
    .A2(\mem.mem[20][1] ));
 sg13g2_a221oi_1 _10732_ (.B2(net3222),
    .C1(net3161),
    .B1(_02877_),
    .A1(_02874_),
    .Y(_02878_),
    .A2(_02875_));
 sg13g2_o21ai_1 _10733_ (.B1(net3117),
    .Y(_02879_),
    .A1(_02872_),
    .A2(_02873_));
 sg13g2_a21oi_1 _10734_ (.A1(_02868_),
    .A2(_02869_),
    .Y(_02880_),
    .B1(net3098));
 sg13g2_o21ai_1 _10735_ (.B1(_02880_),
    .Y(_02881_),
    .A1(_02878_),
    .A2(_02879_));
 sg13g2_mux4_1 _10736_ (.S0(net3950),
    .A0(\mem.mem[40][1] ),
    .A1(\mem.mem[41][1] ),
    .A2(\mem.mem[42][1] ),
    .A3(\mem.mem[43][1] ),
    .S1(net3758),
    .X(_02882_));
 sg13g2_nand2_1 _10737_ (.Y(_02883_),
    .A(net3163),
    .B(_02882_));
 sg13g2_mux4_1 _10738_ (.S0(net3936),
    .A0(\mem.mem[44][1] ),
    .A1(\mem.mem[45][1] ),
    .A2(\mem.mem[46][1] ),
    .A3(\mem.mem[47][1] ),
    .S1(net3753),
    .X(_02884_));
 sg13g2_a21oi_1 _10739_ (.A1(net3684),
    .A2(_02884_),
    .Y(_02885_),
    .B1(net3116));
 sg13g2_nand2b_1 _10740_ (.Y(_02886_),
    .B(\mem.mem[36][1] ),
    .A_N(net3950));
 sg13g2_a21oi_1 _10741_ (.A1(net3950),
    .A2(\mem.mem[37][1] ),
    .Y(_02887_),
    .B1(net3758));
 sg13g2_mux2_1 _10742_ (.A0(\mem.mem[38][1] ),
    .A1(\mem.mem[39][1] ),
    .S(net3946),
    .X(_02888_));
 sg13g2_a21oi_1 _10743_ (.A1(_02886_),
    .A2(_02887_),
    .Y(_02889_),
    .B1(net3163));
 sg13g2_o21ai_1 _10744_ (.B1(_02889_),
    .Y(_02890_),
    .A1(net3225),
    .A2(_02888_));
 sg13g2_mux4_1 _10745_ (.S0(net3932),
    .A0(\mem.mem[32][1] ),
    .A1(\mem.mem[33][1] ),
    .A2(\mem.mem[34][1] ),
    .A3(\mem.mem[35][1] ),
    .S1(net3753),
    .X(_02891_));
 sg13g2_a21oi_1 _10746_ (.A1(net3160),
    .A2(_02891_),
    .Y(_02892_),
    .B1(net3649));
 sg13g2_a221oi_1 _10747_ (.B2(_02892_),
    .C1(net3627),
    .B1(_02890_),
    .A1(_02883_),
    .Y(_02893_),
    .A2(_02885_));
 sg13g2_mux4_1 _10748_ (.S0(net3977),
    .A0(\mem.mem[56][1] ),
    .A1(\mem.mem[57][1] ),
    .A2(\mem.mem[58][1] ),
    .A3(\mem.mem[59][1] ),
    .S1(net3766),
    .X(_02894_));
 sg13g2_mux4_1 _10749_ (.S0(net3983),
    .A0(\mem.mem[60][1] ),
    .A1(\mem.mem[61][1] ),
    .A2(\mem.mem[62][1] ),
    .A3(\mem.mem[63][1] ),
    .S1(net3768),
    .X(_02895_));
 sg13g2_nand2_1 _10750_ (.Y(_02896_),
    .A(net3688),
    .B(_02895_));
 sg13g2_a21oi_1 _10751_ (.A1(net3170),
    .A2(_02894_),
    .Y(_02897_),
    .B1(net3118));
 sg13g2_nand2_1 _10752_ (.Y(_02898_),
    .A(net3958),
    .B(\mem.mem[51][1] ));
 sg13g2_nand2b_1 _10753_ (.Y(_02899_),
    .B(\mem.mem[50][1] ),
    .A_N(net3957));
 sg13g2_nand3_1 _10754_ (.B(_02898_),
    .C(_02899_),
    .A(net3760),
    .Y(_02900_));
 sg13g2_nand2b_1 _10755_ (.Y(_02901_),
    .B(\mem.mem[48][1] ),
    .A_N(net3957));
 sg13g2_a21oi_1 _10756_ (.A1(net3962),
    .A2(\mem.mem[49][1] ),
    .Y(_02902_),
    .B1(net3760));
 sg13g2_a21oi_1 _10757_ (.A1(_02901_),
    .A2(_02902_),
    .Y(_02903_),
    .B1(net3686));
 sg13g2_mux2_1 _10758_ (.A0(\mem.mem[54][1] ),
    .A1(\mem.mem[55][1] ),
    .S(net3976),
    .X(_02904_));
 sg13g2_nand2b_1 _10759_ (.Y(_02905_),
    .B(\mem.mem[52][1] ),
    .A_N(net3976));
 sg13g2_a21oi_1 _10760_ (.A1(net3976),
    .A2(\mem.mem[53][1] ),
    .Y(_02906_),
    .B1(net3766));
 sg13g2_a21oi_1 _10761_ (.A1(_02905_),
    .A2(_02906_),
    .Y(_02907_),
    .B1(net3170));
 sg13g2_o21ai_1 _10762_ (.B1(_02907_),
    .Y(_02908_),
    .A1(net3232),
    .A2(_02904_));
 sg13g2_a21oi_1 _10763_ (.A1(_02900_),
    .A2(_02903_),
    .Y(_02909_),
    .B1(net3652));
 sg13g2_a221oi_1 _10764_ (.B2(_02909_),
    .C1(net3099),
    .B1(_02908_),
    .A1(_02896_),
    .Y(_02910_),
    .A2(_02897_));
 sg13g2_mux2_1 _10765_ (.A0(\mem.mem[74][1] ),
    .A1(\mem.mem[75][1] ),
    .S(net3780),
    .X(_02911_));
 sg13g2_mux2_1 _10766_ (.A0(\mem.mem[72][1] ),
    .A1(\mem.mem[73][1] ),
    .S(net3780),
    .X(_02912_));
 sg13g2_nor2_1 _10767_ (.A(net3695),
    .B(_02912_),
    .Y(_02913_));
 sg13g2_o21ai_1 _10768_ (.B1(net3131),
    .Y(_02914_),
    .A1(net3183),
    .A2(_02911_));
 sg13g2_mux4_1 _10769_ (.S0(net3800),
    .A0(\mem.mem[76][1] ),
    .A1(\mem.mem[77][1] ),
    .A2(\mem.mem[78][1] ),
    .A3(\mem.mem[79][1] ),
    .S1(net3704),
    .X(_02915_));
 sg13g2_a21oi_1 _10770_ (.A1(net3662),
    .A2(_02915_),
    .Y(_02916_),
    .B1(net3103));
 sg13g2_o21ai_1 _10771_ (.B1(_02916_),
    .Y(_02917_),
    .A1(_02913_),
    .A2(_02914_));
 sg13g2_mux4_1 _10772_ (.S0(net3795),
    .A0(\mem.mem[64][1] ),
    .A1(\mem.mem[65][1] ),
    .A2(\mem.mem[66][1] ),
    .A3(\mem.mem[67][1] ),
    .S1(net3699),
    .X(_02918_));
 sg13g2_nand2_1 _10773_ (.Y(_02919_),
    .A(net3127),
    .B(_02918_));
 sg13g2_mux4_1 _10774_ (.S0(net3812),
    .A0(\mem.mem[68][1] ),
    .A1(\mem.mem[69][1] ),
    .A2(\mem.mem[70][1] ),
    .A3(\mem.mem[71][1] ),
    .S1(net3709),
    .X(_02920_));
 sg13g2_a21oi_1 _10775_ (.A1(net3664),
    .A2(_02920_),
    .Y(_02921_),
    .B1(net3635));
 sg13g2_a21oi_1 _10776_ (.A1(_02919_),
    .A2(_02921_),
    .Y(_02922_),
    .B1(net3621));
 sg13g2_and2_1 _10777_ (.A(_02917_),
    .B(_02922_),
    .X(_02923_));
 sg13g2_mux4_1 _10778_ (.S0(net3803),
    .A0(\mem.mem[88][1] ),
    .A1(\mem.mem[89][1] ),
    .A2(\mem.mem[90][1] ),
    .A3(\mem.mem[91][1] ),
    .S1(net3705),
    .X(_02924_));
 sg13g2_nand2b_1 _10779_ (.Y(_02925_),
    .B(\mem.mem[92][1] ),
    .A_N(net3804));
 sg13g2_a21oi_1 _10780_ (.A1(net3804),
    .A2(\mem.mem[93][1] ),
    .Y(_02926_),
    .B1(net3707));
 sg13g2_mux2_1 _10781_ (.A0(\mem.mem[94][1] ),
    .A1(\mem.mem[95][1] ),
    .S(net3804),
    .X(_02927_));
 sg13g2_a21oi_1 _10782_ (.A1(_02925_),
    .A2(_02926_),
    .Y(_02928_),
    .B1(net3129));
 sg13g2_o21ai_1 _10783_ (.B1(_02928_),
    .Y(_02929_),
    .A1(net3183),
    .A2(_02927_));
 sg13g2_a21oi_1 _10784_ (.A1(net3129),
    .A2(_02924_),
    .Y(_02930_),
    .B1(net3104));
 sg13g2_nand2b_1 _10785_ (.Y(_02931_),
    .B(net3814),
    .A_N(\mem.mem[85][1] ));
 sg13g2_o21ai_1 _10786_ (.B1(_02931_),
    .Y(_02932_),
    .A1(net3814),
    .A2(\mem.mem[84][1] ));
 sg13g2_mux2_1 _10787_ (.A0(\mem.mem[86][1] ),
    .A1(\mem.mem[87][1] ),
    .S(net3814),
    .X(_02933_));
 sg13g2_o21ai_1 _10788_ (.B1(net3665),
    .Y(_02934_),
    .A1(net3186),
    .A2(_02933_));
 sg13g2_a21o_1 _10789_ (.A2(_02932_),
    .A1(net3186),
    .B1(_02934_),
    .X(_02935_));
 sg13g2_mux4_1 _10790_ (.S0(net3804),
    .A0(\mem.mem[80][1] ),
    .A1(\mem.mem[81][1] ),
    .A2(\mem.mem[82][1] ),
    .A3(\mem.mem[83][1] ),
    .S1(net3711),
    .X(_02936_));
 sg13g2_a21oi_1 _10791_ (.A1(net3130),
    .A2(_02936_),
    .Y(_02937_),
    .B1(net3635));
 sg13g2_a221oi_1 _10792_ (.B2(_02937_),
    .C1(net3094),
    .B1(_02935_),
    .A1(_02929_),
    .Y(_02938_),
    .A2(_02930_));
 sg13g2_mux4_1 _10793_ (.S0(net3841),
    .A0(\mem.mem[120][1] ),
    .A1(\mem.mem[121][1] ),
    .A2(\mem.mem[122][1] ),
    .A3(\mem.mem[123][1] ),
    .S1(net3721),
    .X(_02939_));
 sg13g2_mux4_1 _10794_ (.S0(net3849),
    .A0(\mem.mem[124][1] ),
    .A1(\mem.mem[125][1] ),
    .A2(\mem.mem[126][1] ),
    .A3(\mem.mem[127][1] ),
    .S1(net3725),
    .X(_02940_));
 sg13g2_nand2_1 _10795_ (.Y(_02941_),
    .A(net3669),
    .B(_02940_));
 sg13g2_a21oi_1 _10796_ (.A1(net3134),
    .A2(_02939_),
    .Y(_02942_),
    .B1(net3108));
 sg13g2_mux4_1 _10797_ (.S0(net3833),
    .A0(\mem.mem[112][1] ),
    .A1(\mem.mem[113][1] ),
    .A2(\mem.mem[114][1] ),
    .A3(\mem.mem[115][1] ),
    .S1(net3719),
    .X(_02943_));
 sg13g2_nor2b_1 _10798_ (.A(net3821),
    .B_N(\mem.mem[118][1] ),
    .Y(_02944_));
 sg13g2_a21oi_1 _10799_ (.A1(net3821),
    .A2(\mem.mem[119][1] ),
    .Y(_02945_),
    .B1(_02944_));
 sg13g2_mux2_1 _10800_ (.A0(\mem.mem[116][1] ),
    .A1(\mem.mem[117][1] ),
    .S(net3822),
    .X(_02946_));
 sg13g2_o21ai_1 _10801_ (.B1(net3670),
    .Y(_02947_),
    .A1(net3714),
    .A2(_02946_));
 sg13g2_a21o_1 _10802_ (.A2(_02945_),
    .A1(net3714),
    .B1(_02947_),
    .X(_02948_));
 sg13g2_a21oi_1 _10803_ (.A1(net3137),
    .A2(_02943_),
    .Y(_02949_),
    .B1(net3639));
 sg13g2_a221oi_1 _10804_ (.B2(_02949_),
    .C1(net3095),
    .B1(_02948_),
    .A1(_02941_),
    .Y(_02950_),
    .A2(_02942_));
 sg13g2_mux4_1 _10805_ (.S0(net3902),
    .A0(\mem.mem[108][1] ),
    .A1(\mem.mem[109][1] ),
    .A2(\mem.mem[110][1] ),
    .A3(\mem.mem[111][1] ),
    .S1(net3743),
    .X(_02951_));
 sg13g2_nand2_1 _10806_ (.Y(_02952_),
    .A(net3678),
    .B(_02951_));
 sg13g2_nand2_1 _10807_ (.Y(_02953_),
    .A(net3917),
    .B(\mem.mem[107][1] ));
 sg13g2_nand2b_1 _10808_ (.Y(_02954_),
    .B(\mem.mem[106][1] ),
    .A_N(net3917));
 sg13g2_nand3_1 _10809_ (.B(_02953_),
    .C(_02954_),
    .A(net3749),
    .Y(_02955_));
 sg13g2_nand2b_1 _10810_ (.Y(_02956_),
    .B(\mem.mem[104][1] ),
    .A_N(net3918));
 sg13g2_a21oi_1 _10811_ (.A1(net3918),
    .A2(\mem.mem[105][1] ),
    .Y(_02957_),
    .B1(net3748));
 sg13g2_a21oi_1 _10812_ (.A1(_02956_),
    .A2(_02957_),
    .Y(_02958_),
    .B1(net3680));
 sg13g2_a21oi_2 _10813_ (.B1(net3113),
    .Y(_02959_),
    .A2(_02958_),
    .A1(_02955_));
 sg13g2_nor2b_1 _10814_ (.A(net3903),
    .B_N(\mem.mem[98][1] ),
    .Y(_02960_));
 sg13g2_a21oi_1 _10815_ (.A1(net3903),
    .A2(\mem.mem[99][1] ),
    .Y(_02961_),
    .B1(_02960_));
 sg13g2_mux2_1 _10816_ (.A0(\mem.mem[96][1] ),
    .A1(\mem.mem[97][1] ),
    .S(net3900),
    .X(_02962_));
 sg13g2_o21ai_1 _10817_ (.B1(net3154),
    .Y(_02963_),
    .A1(net3743),
    .A2(_02962_));
 sg13g2_a21o_1 _10818_ (.A2(_02961_),
    .A1(net3743),
    .B1(_02963_),
    .X(_02964_));
 sg13g2_mux4_1 _10819_ (.S0(net3919),
    .A0(\mem.mem[100][1] ),
    .A1(\mem.mem[101][1] ),
    .A2(\mem.mem[102][1] ),
    .A3(\mem.mem[103][1] ),
    .S1(net3750),
    .X(_02965_));
 sg13g2_a21oi_1 _10820_ (.A1(net3677),
    .A2(_02965_),
    .Y(_02966_),
    .B1(net3646));
 sg13g2_a221oi_1 _10821_ (.B2(_02966_),
    .C1(net3631),
    .B1(_02964_),
    .A1(_02952_),
    .Y(_02967_),
    .A2(_02959_));
 sg13g2_o21ai_1 _10822_ (.B1(net3090),
    .Y(_02968_),
    .A1(_02923_),
    .A2(_02938_));
 sg13g2_o21ai_1 _10823_ (.B1(net3616),
    .Y(_02969_),
    .A1(_02950_),
    .A2(_02967_));
 sg13g2_nand3_1 _10824_ (.B(_02968_),
    .C(_02969_),
    .A(net3612),
    .Y(_02970_));
 sg13g2_a21oi_2 _10825_ (.B1(net3618),
    .Y(_02971_),
    .A2(_02881_),
    .A1(_02865_));
 sg13g2_o21ai_1 _10826_ (.B1(net3618),
    .Y(_02972_),
    .A1(_02893_),
    .A2(_02910_));
 sg13g2_nand2_2 _10827_ (.Y(_02973_),
    .A(_02148_),
    .B(_02972_));
 sg13g2_o21ai_1 _10828_ (.B1(_02970_),
    .Y(_02974_),
    .A1(_02971_),
    .A2(_02973_));
 sg13g2_mux4_1 _10829_ (.S0(net3874),
    .A0(\mem.mem[164][1] ),
    .A1(\mem.mem[165][1] ),
    .A2(\mem.mem[166][1] ),
    .A3(\mem.mem[167][1] ),
    .S1(net3734),
    .X(_02975_));
 sg13g2_mux4_1 _10830_ (.S0(net3838),
    .A0(\mem.mem[160][1] ),
    .A1(\mem.mem[161][1] ),
    .A2(\mem.mem[162][1] ),
    .A3(\mem.mem[163][1] ),
    .S1(net3718),
    .X(_02976_));
 sg13g2_nand2_1 _10831_ (.Y(_02977_),
    .A(net3138),
    .B(_02976_));
 sg13g2_a21oi_1 _10832_ (.A1(net3669),
    .A2(_02975_),
    .Y(_02978_),
    .B1(net3643));
 sg13g2_nand2b_1 _10833_ (.Y(_02979_),
    .B(\mem.mem[172][1] ),
    .A_N(net3835));
 sg13g2_a21oi_1 _10834_ (.A1(net3835),
    .A2(\mem.mem[173][1] ),
    .Y(_02980_),
    .B1(net3719));
 sg13g2_mux2_1 _10835_ (.A0(\mem.mem[174][1] ),
    .A1(\mem.mem[175][1] ),
    .S(net3836),
    .X(_02981_));
 sg13g2_a21oi_1 _10836_ (.A1(_02979_),
    .A2(_02980_),
    .Y(_02982_),
    .B1(net3137));
 sg13g2_o21ai_1 _10837_ (.B1(_02982_),
    .Y(_02983_),
    .A1(net3191),
    .A2(_02981_));
 sg13g2_nand2b_1 _10838_ (.Y(_02984_),
    .B(\mem.mem[168][1] ),
    .A_N(net3894));
 sg13g2_nand2_1 _10839_ (.Y(_02985_),
    .A(net3894),
    .B(\mem.mem[169][1] ));
 sg13g2_nand3_1 _10840_ (.B(_02984_),
    .C(_02985_),
    .A(net3209),
    .Y(_02986_));
 sg13g2_nor2b_1 _10841_ (.A(net3894),
    .B_N(\mem.mem[170][1] ),
    .Y(_02987_));
 sg13g2_a21oi_1 _10842_ (.A1(net3894),
    .A2(\mem.mem[171][1] ),
    .Y(_02988_),
    .B1(_02987_));
 sg13g2_a21oi_1 _10843_ (.A1(net3742),
    .A2(_02988_),
    .Y(_02989_),
    .B1(net3677));
 sg13g2_a21oi_1 _10844_ (.A1(_02986_),
    .A2(_02989_),
    .Y(_02990_),
    .B1(net3111));
 sg13g2_a221oi_1 _10845_ (.B2(_02990_),
    .C1(net3625),
    .B1(_02983_),
    .A1(_02977_),
    .Y(_02991_),
    .A2(_02978_));
 sg13g2_mux4_1 _10846_ (.S0(net3852),
    .A0(\mem.mem[176][1] ),
    .A1(\mem.mem[177][1] ),
    .A2(\mem.mem[178][1] ),
    .A3(\mem.mem[179][1] ),
    .S1(net3726),
    .X(_02992_));
 sg13g2_nand2_1 _10847_ (.Y(_02993_),
    .A(net3859),
    .B(\mem.mem[183][1] ));
 sg13g2_nand2b_1 _10848_ (.Y(_02994_),
    .B(\mem.mem[182][1] ),
    .A_N(net3859));
 sg13g2_nand3_1 _10849_ (.B(_02993_),
    .C(_02994_),
    .A(net3729),
    .Y(_02995_));
 sg13g2_nand2b_1 _10850_ (.Y(_02996_),
    .B(\mem.mem[180][1] ),
    .A_N(net3859));
 sg13g2_a21oi_1 _10851_ (.A1(net3859),
    .A2(\mem.mem[181][1] ),
    .Y(_02997_),
    .B1(net3728));
 sg13g2_a21oi_1 _10852_ (.A1(_02996_),
    .A2(_02997_),
    .Y(_02998_),
    .B1(net3142));
 sg13g2_a221oi_1 _10853_ (.B2(_02998_),
    .C1(net3640),
    .B1(_02995_),
    .A1(net3142),
    .Y(_02999_),
    .A2(_02992_));
 sg13g2_mux2_1 _10854_ (.A0(\mem.mem[184][1] ),
    .A1(\mem.mem[185][1] ),
    .S(net3848),
    .X(_03000_));
 sg13g2_nor2_1 _10855_ (.A(net3724),
    .B(_03000_),
    .Y(_03001_));
 sg13g2_mux2_1 _10856_ (.A0(\mem.mem[186][1] ),
    .A1(\mem.mem[187][1] ),
    .S(net3848),
    .X(_03002_));
 sg13g2_o21ai_1 _10857_ (.B1(net3145),
    .Y(_03003_),
    .A1(net3197),
    .A2(_03002_));
 sg13g2_nand2b_1 _10858_ (.Y(_03004_),
    .B(\mem.mem[188][1] ),
    .A_N(net3846));
 sg13g2_a21oi_1 _10859_ (.A1(net3846),
    .A2(\mem.mem[189][1] ),
    .Y(_03005_),
    .B1(net3723));
 sg13g2_nor2b_1 _10860_ (.A(net3846),
    .B_N(\mem.mem[190][1] ),
    .Y(_03006_));
 sg13g2_a21oi_1 _10861_ (.A1(net3847),
    .A2(\mem.mem[191][1] ),
    .Y(_03007_),
    .B1(_03006_));
 sg13g2_a221oi_1 _10862_ (.B2(net3723),
    .C1(net3140),
    .B1(_03007_),
    .A1(_03004_),
    .Y(_03008_),
    .A2(_03005_));
 sg13g2_o21ai_1 _10863_ (.B1(net3641),
    .Y(_03009_),
    .A1(_03001_),
    .A2(_03003_));
 sg13g2_o21ai_1 _10864_ (.B1(net3622),
    .Y(_03010_),
    .A1(_03008_),
    .A2(_03009_));
 sg13g2_nor2_2 _10865_ (.A(_02999_),
    .B(_03010_),
    .Y(_03011_));
 sg13g2_o21ai_1 _10866_ (.B1(net3617),
    .Y(_03012_),
    .A1(_02991_),
    .A2(_03011_));
 sg13g2_mux4_1 _10867_ (.S0(net3887),
    .A0(\mem.mem[128][1] ),
    .A1(\mem.mem[129][1] ),
    .A2(\mem.mem[130][1] ),
    .A3(\mem.mem[131][1] ),
    .S1(net3740),
    .X(_03013_));
 sg13g2_nand2_1 _10868_ (.Y(_03014_),
    .A(net3890),
    .B(\mem.mem[135][1] ));
 sg13g2_nand2b_1 _10869_ (.Y(_03015_),
    .B(\mem.mem[134][1] ),
    .A_N(net3911));
 sg13g2_nand3_1 _10870_ (.B(_03014_),
    .C(_03015_),
    .A(net3739),
    .Y(_03016_));
 sg13g2_nand2b_1 _10871_ (.Y(_03017_),
    .B(\mem.mem[132][1] ),
    .A_N(net3886));
 sg13g2_a21oi_1 _10872_ (.A1(net3890),
    .A2(\mem.mem[133][1] ),
    .Y(_03018_),
    .B1(net3740));
 sg13g2_a21oi_1 _10873_ (.A1(_03017_),
    .A2(_03018_),
    .Y(_03019_),
    .B1(net3152));
 sg13g2_a221oi_1 _10874_ (.B2(_03019_),
    .C1(net3647),
    .B1(_03016_),
    .A1(net3155),
    .Y(_03020_),
    .A2(_03013_));
 sg13g2_nand2b_1 _10875_ (.Y(_03021_),
    .B(\mem.mem[140][1] ),
    .A_N(net3907));
 sg13g2_a21oi_1 _10876_ (.A1(net3907),
    .A2(\mem.mem[141][1] ),
    .Y(_03022_),
    .B1(net3747));
 sg13g2_nand2_1 _10877_ (.Y(_03023_),
    .A(net3907),
    .B(\mem.mem[143][1] ));
 sg13g2_nand2b_1 _10878_ (.Y(_03024_),
    .B(\mem.mem[142][1] ),
    .A_N(net3910));
 sg13g2_nand3_1 _10879_ (.B(_03023_),
    .C(_03024_),
    .A(net3746),
    .Y(_03025_));
 sg13g2_a21oi_1 _10880_ (.A1(_03021_),
    .A2(_03022_),
    .Y(_03026_),
    .B1(net3155));
 sg13g2_nand2b_1 _10881_ (.Y(_03027_),
    .B(\mem.mem[136][1] ),
    .A_N(net3899));
 sg13g2_nand2_1 _10882_ (.Y(_03028_),
    .A(net3898),
    .B(\mem.mem[137][1] ));
 sg13g2_nand3_1 _10883_ (.B(_03027_),
    .C(_03028_),
    .A(net3213),
    .Y(_03029_));
 sg13g2_nor2b_1 _10884_ (.A(net3897),
    .B_N(\mem.mem[138][1] ),
    .Y(_03030_));
 sg13g2_a21oi_1 _10885_ (.A1(net3897),
    .A2(\mem.mem[139][1] ),
    .Y(_03031_),
    .B1(_03030_));
 sg13g2_a21oi_1 _10886_ (.A1(net3742),
    .A2(_03031_),
    .Y(_03032_),
    .B1(net3679));
 sg13g2_a221oi_1 _10887_ (.B2(_03032_),
    .C1(net3113),
    .B1(_03029_),
    .A1(_03025_),
    .Y(_03033_),
    .A2(_03026_));
 sg13g2_nor3_1 _10888_ (.A(net3625),
    .B(_03020_),
    .C(_03033_),
    .Y(_03034_));
 sg13g2_mux4_1 _10889_ (.S0(net3921),
    .A0(\mem.mem[144][1] ),
    .A1(\mem.mem[145][1] ),
    .A2(\mem.mem[146][1] ),
    .A3(\mem.mem[147][1] ),
    .S1(net3750),
    .X(_03035_));
 sg13g2_nand2_1 _10890_ (.Y(_03036_),
    .A(net3965),
    .B(\mem.mem[151][1] ));
 sg13g2_nand2b_1 _10891_ (.Y(_03037_),
    .B(\mem.mem[150][1] ),
    .A_N(net3965));
 sg13g2_nand3_1 _10892_ (.B(_03036_),
    .C(_03037_),
    .A(net3762),
    .Y(_03038_));
 sg13g2_nand2b_1 _10893_ (.Y(_03039_),
    .B(\mem.mem[148][1] ),
    .A_N(net3981));
 sg13g2_a21oi_1 _10894_ (.A1(net3981),
    .A2(\mem.mem[149][1] ),
    .Y(_03040_),
    .B1(net3768));
 sg13g2_a21oi_2 _10895_ (.B1(net3172),
    .Y(_03041_),
    .A2(_03040_),
    .A1(_03039_));
 sg13g2_a221oi_1 _10896_ (.B2(_03041_),
    .C1(net3651),
    .B1(_03038_),
    .A1(net3168),
    .Y(_03042_),
    .A2(_03035_));
 sg13g2_mux2_1 _10897_ (.A0(\mem.mem[152][1] ),
    .A1(\mem.mem[153][1] ),
    .S(net3986),
    .X(_03043_));
 sg13g2_nor2_1 _10898_ (.A(net3768),
    .B(_03043_),
    .Y(_03044_));
 sg13g2_mux2_1 _10899_ (.A0(\mem.mem[154][1] ),
    .A1(\mem.mem[155][1] ),
    .S(net3986),
    .X(_03045_));
 sg13g2_o21ai_1 _10900_ (.B1(net3173),
    .Y(_03046_),
    .A1(net3235),
    .A2(_03045_));
 sg13g2_nand2b_1 _10901_ (.Y(_03047_),
    .B(\mem.mem[156][1] ),
    .A_N(net3964));
 sg13g2_a21oi_1 _10902_ (.A1(net3966),
    .A2(\mem.mem[157][1] ),
    .Y(_03048_),
    .B1(net3749));
 sg13g2_nor2b_1 _10903_ (.A(net3964),
    .B_N(\mem.mem[158][1] ),
    .Y(_03049_));
 sg13g2_a21oi_1 _10904_ (.A1(net3964),
    .A2(\mem.mem[159][1] ),
    .Y(_03050_),
    .B1(_03049_));
 sg13g2_a221oi_1 _10905_ (.B2(net3749),
    .C1(net3159),
    .B1(_03050_),
    .A1(_03047_),
    .Y(_03051_),
    .A2(_03048_));
 sg13g2_o21ai_1 _10906_ (.B1(net3653),
    .Y(_03052_),
    .A1(_03044_),
    .A2(_03046_));
 sg13g2_o21ai_1 _10907_ (.B1(net3629),
    .Y(_03053_),
    .A1(_03051_),
    .A2(_03052_));
 sg13g2_nor2_2 _10908_ (.A(_03042_),
    .B(_03053_),
    .Y(_03054_));
 sg13g2_o21ai_1 _10909_ (.B1(net3093),
    .Y(_03055_),
    .A1(_03034_),
    .A2(_03054_));
 sg13g2_a21o_1 _10910_ (.A2(_03055_),
    .A1(_03012_),
    .B1(net3613),
    .X(_03056_));
 sg13g2_mux4_1 _10911_ (.S0(net3793),
    .A0(\mem.mem[212][1] ),
    .A1(\mem.mem[213][1] ),
    .A2(\mem.mem[214][1] ),
    .A3(\mem.mem[215][1] ),
    .S1(net3699),
    .X(_03057_));
 sg13g2_nand2_1 _10912_ (.Y(_03058_),
    .A(net3660),
    .B(_03057_));
 sg13g2_mux4_1 _10913_ (.S0(net3785),
    .A0(\mem.mem[208][1] ),
    .A1(\mem.mem[209][1] ),
    .A2(\mem.mem[210][1] ),
    .A3(\mem.mem[211][1] ),
    .S1(net3697),
    .X(_03059_));
 sg13g2_a21oi_1 _10914_ (.A1(net3125),
    .A2(_03059_),
    .Y(_03060_),
    .B1(net3633));
 sg13g2_mux2_1 _10915_ (.A0(\mem.mem[216][1] ),
    .A1(\mem.mem[217][1] ),
    .S(net3787),
    .X(_03061_));
 sg13g2_nor2_1 _10916_ (.A(net3696),
    .B(_03061_),
    .Y(_03062_));
 sg13g2_mux2_1 _10917_ (.A0(\mem.mem[218][1] ),
    .A1(\mem.mem[219][1] ),
    .S(net3788),
    .X(_03063_));
 sg13g2_o21ai_1 _10918_ (.B1(net3125),
    .Y(_03064_),
    .A1(net3178),
    .A2(_03063_));
 sg13g2_nand2b_1 _10919_ (.Y(_03065_),
    .B(\mem.mem[220][1] ),
    .A_N(net3793));
 sg13g2_a21oi_1 _10920_ (.A1(net3793),
    .A2(\mem.mem[221][1] ),
    .Y(_03066_),
    .B1(net3698));
 sg13g2_nor2b_1 _10921_ (.A(net3787),
    .B_N(\mem.mem[222][1] ),
    .Y(_03067_));
 sg13g2_a21oi_1 _10922_ (.A1(net3793),
    .A2(\mem.mem[223][1] ),
    .Y(_03068_),
    .B1(_03067_));
 sg13g2_a221oi_1 _10923_ (.B2(net3698),
    .C1(net3127),
    .B1(_03068_),
    .A1(_03065_),
    .Y(_03069_),
    .A2(_03066_));
 sg13g2_o21ai_1 _10924_ (.B1(net3633),
    .Y(_03070_),
    .A1(_03062_),
    .A2(_03064_));
 sg13g2_a21oi_1 _10925_ (.A1(_03058_),
    .A2(_03060_),
    .Y(_03071_),
    .B1(net3094));
 sg13g2_o21ai_1 _10926_ (.B1(_03071_),
    .Y(_03072_),
    .A1(_03069_),
    .A2(_03070_));
 sg13g2_nand2b_1 _10927_ (.Y(_03073_),
    .B(\mem.mem[198][1] ),
    .A_N(net3776));
 sg13g2_a21oi_1 _10928_ (.A1(net3776),
    .A2(\mem.mem[199][1] ),
    .Y(_03074_),
    .B1(net3176));
 sg13g2_nor2b_1 _10929_ (.A(net3774),
    .B_N(\mem.mem[196][1] ),
    .Y(_03075_));
 sg13g2_a21oi_1 _10930_ (.A1(net3774),
    .A2(\mem.mem[197][1] ),
    .Y(_03076_),
    .B1(_03075_));
 sg13g2_a221oi_1 _10931_ (.B2(net3176),
    .C1(net3122),
    .B1(_03076_),
    .A1(_03073_),
    .Y(_03077_),
    .A2(_03074_));
 sg13g2_mux2_1 _10932_ (.A0(\mem.mem[192][1] ),
    .A1(\mem.mem[193][1] ),
    .S(net3772),
    .X(_03078_));
 sg13g2_nor2_1 _10933_ (.A(net3691),
    .B(_03078_),
    .Y(_03079_));
 sg13g2_mux2_1 _10934_ (.A0(\mem.mem[194][1] ),
    .A1(\mem.mem[195][1] ),
    .S(net3771),
    .X(_03080_));
 sg13g2_o21ai_1 _10935_ (.B1(net3121),
    .Y(_03081_),
    .A1(net3175),
    .A2(_03080_));
 sg13g2_o21ai_1 _10936_ (.B1(net3101),
    .Y(_03082_),
    .A1(_03079_),
    .A2(_03081_));
 sg13g2_nor2_1 _10937_ (.A(_03077_),
    .B(_03082_),
    .Y(_03083_));
 sg13g2_nor2b_1 _10938_ (.A(net3781),
    .B_N(\mem.mem[204][1] ),
    .Y(_03084_));
 sg13g2_a21oi_1 _10939_ (.A1(net3781),
    .A2(\mem.mem[205][1] ),
    .Y(_03085_),
    .B1(_03084_));
 sg13g2_nand2b_1 _10940_ (.Y(_03086_),
    .B(\mem.mem[206][1] ),
    .A_N(net3780));
 sg13g2_a21oi_1 _10941_ (.A1(net3780),
    .A2(\mem.mem[207][1] ),
    .Y(_03087_),
    .B1(net3177));
 sg13g2_a221oi_1 _10942_ (.B2(_03087_),
    .C1(net3124),
    .B1(_03086_),
    .A1(net3177),
    .Y(_03088_),
    .A2(_03085_));
 sg13g2_nor2b_1 _10943_ (.A(net3780),
    .B_N(\mem.mem[200][1] ),
    .Y(_03089_));
 sg13g2_a21oi_1 _10944_ (.A1(net3779),
    .A2(\mem.mem[201][1] ),
    .Y(_03090_),
    .B1(_03089_));
 sg13g2_nand2b_1 _10945_ (.Y(_03091_),
    .B(\mem.mem[202][1] ),
    .A_N(net3779));
 sg13g2_a21oi_1 _10946_ (.A1(net3780),
    .A2(\mem.mem[203][1] ),
    .Y(_03092_),
    .B1(net3177));
 sg13g2_a221oi_1 _10947_ (.B2(_03092_),
    .C1(net3658),
    .B1(_03091_),
    .A1(net3177),
    .Y(_03093_),
    .A2(_03090_));
 sg13g2_nor3_1 _10948_ (.A(net3101),
    .B(_03088_),
    .C(_03093_),
    .Y(_03094_));
 sg13g2_or3_1 _10949_ (.A(net3620),
    .B(_03083_),
    .C(_03094_),
    .X(_03095_));
 sg13g2_nand3_1 _10950_ (.B(_03072_),
    .C(_03095_),
    .A(net3090),
    .Y(_03096_));
 sg13g2_nor2_1 _10951_ (.A(net3868),
    .B(\mem.mem[230][1] ),
    .Y(_03097_));
 sg13g2_nor2b_1 _10952_ (.A(\mem.mem[231][1] ),
    .B_N(net3868),
    .Y(_03098_));
 sg13g2_nor3_1 _10953_ (.A(net3200),
    .B(_03097_),
    .C(_03098_),
    .Y(_03099_));
 sg13g2_nor2_1 _10954_ (.A(net3868),
    .B(\mem.mem[228][1] ),
    .Y(_03100_));
 sg13g2_nor2b_1 _10955_ (.A(\mem.mem[229][1] ),
    .B_N(net3868),
    .Y(_03101_));
 sg13g2_nor3_1 _10956_ (.A(net3736),
    .B(_03100_),
    .C(_03101_),
    .Y(_03102_));
 sg13g2_nor3_1 _10957_ (.A(net3147),
    .B(_03099_),
    .C(_03102_),
    .Y(_03103_));
 sg13g2_mux4_1 _10958_ (.S0(net3866),
    .A0(\mem.mem[224][1] ),
    .A1(\mem.mem[225][1] ),
    .A2(\mem.mem[226][1] ),
    .A3(\mem.mem[227][1] ),
    .S1(net3733),
    .X(_03104_));
 sg13g2_nor2_1 _10959_ (.A(net3674),
    .B(_03104_),
    .Y(_03105_));
 sg13g2_o21ai_1 _10960_ (.B1(net3111),
    .Y(_03106_),
    .A1(_03103_),
    .A2(_03105_));
 sg13g2_mux4_1 _10961_ (.S0(net3832),
    .A0(\mem.mem[232][1] ),
    .A1(\mem.mem[233][1] ),
    .A2(\mem.mem[234][1] ),
    .A3(\mem.mem[235][1] ),
    .S1(net3716),
    .X(_03107_));
 sg13g2_mux2_1 _10962_ (.A0(\mem.mem[238][1] ),
    .A1(\mem.mem[239][1] ),
    .S(net3838),
    .X(_03108_));
 sg13g2_nand2b_1 _10963_ (.Y(_03109_),
    .B(\mem.mem[236][1] ),
    .A_N(net3830));
 sg13g2_a21oi_1 _10964_ (.A1(net3838),
    .A2(\mem.mem[237][1] ),
    .Y(_03110_),
    .B1(net3718));
 sg13g2_a21oi_1 _10965_ (.A1(_03109_),
    .A2(_03110_),
    .Y(_03111_),
    .B1(net3136));
 sg13g2_o21ai_1 _10966_ (.B1(_03111_),
    .Y(_03112_),
    .A1(net3190),
    .A2(_03108_));
 sg13g2_a21oi_1 _10967_ (.A1(net3136),
    .A2(_03107_),
    .Y(_03113_),
    .B1(net3107));
 sg13g2_a21oi_1 _10968_ (.A1(_03112_),
    .A2(_03113_),
    .Y(_03114_),
    .B1(net3623));
 sg13g2_mux4_1 _10969_ (.S0(net3828),
    .A0(\mem.mem[240][1] ),
    .A1(\mem.mem[241][1] ),
    .A2(\mem.mem[242][1] ),
    .A3(\mem.mem[243][1] ),
    .S1(net3715),
    .X(_03115_));
 sg13g2_and2_1 _10970_ (.A(net3135),
    .B(_03115_),
    .X(_03116_));
 sg13g2_nor2b_1 _10971_ (.A(net3819),
    .B_N(\mem.mem[244][1] ),
    .Y(_03117_));
 sg13g2_a21oi_1 _10972_ (.A1(net3828),
    .A2(\mem.mem[245][1] ),
    .Y(_03118_),
    .B1(_03117_));
 sg13g2_nand2b_1 _10973_ (.Y(_03119_),
    .B(\mem.mem[246][1] ),
    .A_N(net3828));
 sg13g2_a21oi_1 _10974_ (.A1(net3828),
    .A2(\mem.mem[247][1] ),
    .Y(_03120_),
    .B1(net3190));
 sg13g2_a221oi_1 _10975_ (.B2(_03120_),
    .C1(net3133),
    .B1(_03119_),
    .A1(net3190),
    .Y(_03121_),
    .A2(_03118_));
 sg13g2_or3_1 _10976_ (.A(net3639),
    .B(_03116_),
    .C(_03121_),
    .X(_03122_));
 sg13g2_mux4_1 _10977_ (.S0(net3829),
    .A0(\mem.mem[248][1] ),
    .A1(\mem.mem[249][1] ),
    .A2(\mem.mem[250][1] ),
    .A3(\mem.mem[251][1] ),
    .S1(net3717),
    .X(_03123_));
 sg13g2_nand2_1 _10978_ (.Y(_03124_),
    .A(net3136),
    .B(_03123_));
 sg13g2_a21oi_1 _10979_ (.A1(net3670),
    .A2(\mem.mem[252][1] ),
    .Y(_03125_),
    .B1(net3107));
 sg13g2_a21oi_1 _10980_ (.A1(_03124_),
    .A2(_03125_),
    .Y(_03126_),
    .B1(net3095));
 sg13g2_a221oi_1 _10981_ (.B2(_03126_),
    .C1(net3091),
    .B1(_03122_),
    .A1(_03106_),
    .Y(_03127_),
    .A2(_03114_));
 sg13g2_nor2_2 _10982_ (.A(net3089),
    .B(_03127_),
    .Y(_03128_));
 sg13g2_a21oi_1 _10983_ (.A1(_03096_),
    .A2(_03128_),
    .Y(_03129_),
    .B1(_02149_));
 sg13g2_a221oi_1 _10984_ (.B2(_03129_),
    .C1(_02258_),
    .B1(_03056_),
    .A1(_02149_),
    .Y(_03130_),
    .A2(_02974_));
 sg13g2_a21oi_2 _10985_ (.B1(_03130_),
    .Y(_03131_),
    .A2(_02536_),
    .A1(net2));
 sg13g2_o21ai_1 _10986_ (.B1(net4006),
    .Y(_03132_),
    .A1(net5194),
    .A2(_02534_));
 sg13g2_a21oi_1 _10987_ (.A1(_02534_),
    .A2(_03131_),
    .Y(_00596_),
    .B1(_03132_));
 sg13g2_nand2_2 _10988_ (.Y(_03133_),
    .A(net3),
    .B(_02536_));
 sg13g2_a21oi_1 _10989_ (.A1(net3879),
    .A2(\mem.mem[5][2] ),
    .Y(_03134_),
    .B1(net3738));
 sg13g2_o21ai_1 _10990_ (.B1(_03134_),
    .Y(_03135_),
    .A1(net3879),
    .A2(_02151_));
 sg13g2_nor2b_1 _10991_ (.A(net3882),
    .B_N(\mem.mem[6][2] ),
    .Y(_03136_));
 sg13g2_a21oi_1 _10992_ (.A1(net3879),
    .A2(\mem.mem[7][2] ),
    .Y(_03137_),
    .B1(_03136_));
 sg13g2_a21oi_1 _10993_ (.A1(net3738),
    .A2(_03137_),
    .Y(_03138_),
    .B1(net3150));
 sg13g2_mux4_1 _10994_ (.S0(net3925),
    .A0(\mem.mem[0][2] ),
    .A1(\mem.mem[1][2] ),
    .A2(\mem.mem[2][2] ),
    .A3(\mem.mem[3][2] ),
    .S1(net3752),
    .X(_03139_));
 sg13g2_a221oi_1 _10995_ (.B2(net3150),
    .C1(net3644),
    .B1(_03139_),
    .A1(_03135_),
    .Y(_03140_),
    .A2(_03138_));
 sg13g2_mux4_1 _10996_ (.S0(net3877),
    .A0(\mem.mem[8][2] ),
    .A1(\mem.mem[9][2] ),
    .A2(\mem.mem[10][2] ),
    .A3(\mem.mem[11][2] ),
    .S1(net3735),
    .X(_03141_));
 sg13g2_a21oi_1 _10997_ (.A1(net3889),
    .A2(\mem.mem[15][2] ),
    .Y(_03142_),
    .B1(net3207));
 sg13g2_o21ai_1 _10998_ (.B1(_03142_),
    .Y(_03143_),
    .A1(net3888),
    .A2(_02152_));
 sg13g2_nand2b_1 _10999_ (.Y(_03144_),
    .B(\mem.mem[12][2] ),
    .A_N(net3888));
 sg13g2_a21oi_1 _11000_ (.A1(net3888),
    .A2(\mem.mem[13][2] ),
    .Y(_03145_),
    .B1(net3739));
 sg13g2_a21oi_1 _11001_ (.A1(_03144_),
    .A2(_03145_),
    .Y(_03146_),
    .B1(net3153));
 sg13g2_a221oi_1 _11002_ (.B2(_03146_),
    .C1(net3111),
    .B1(_03143_),
    .A1(net3152),
    .Y(_03147_),
    .A2(_03141_));
 sg13g2_o21ai_1 _11003_ (.B1(net3098),
    .Y(_03148_),
    .A1(_03140_),
    .A2(_03147_));
 sg13g2_nand2b_1 _11004_ (.Y(_03149_),
    .B(\mem.mem[22][2] ),
    .A_N(net3939));
 sg13g2_a21oi_1 _11005_ (.A1(net3939),
    .A2(\mem.mem[23][2] ),
    .Y(_03150_),
    .B1(net3227));
 sg13g2_nor2b_1 _11006_ (.A(net3942),
    .B_N(\mem.mem[20][2] ),
    .Y(_03151_));
 sg13g2_a21oi_1 _11007_ (.A1(net3942),
    .A2(\mem.mem[21][2] ),
    .Y(_03152_),
    .B1(_03151_));
 sg13g2_a221oi_1 _11008_ (.B2(net3227),
    .C1(net3161),
    .B1(_03152_),
    .A1(_03149_),
    .Y(_03153_),
    .A2(_03150_));
 sg13g2_nor2b_1 _11009_ (.A(net3927),
    .B_N(\mem.mem[16][2] ),
    .Y(_03154_));
 sg13g2_a21oi_1 _11010_ (.A1(net3927),
    .A2(\mem.mem[17][2] ),
    .Y(_03155_),
    .B1(_03154_));
 sg13g2_nand2b_1 _11011_ (.Y(_03156_),
    .B(\mem.mem[18][2] ),
    .A_N(net3927));
 sg13g2_a21oi_1 _11012_ (.A1(net3927),
    .A2(\mem.mem[19][2] ),
    .Y(_03157_),
    .B1(net3219));
 sg13g2_a221oi_1 _11013_ (.B2(_03157_),
    .C1(net3682),
    .B1(_03156_),
    .A1(net3221),
    .Y(_03158_),
    .A2(_03155_));
 sg13g2_nor3_1 _11014_ (.A(net3650),
    .B(_03153_),
    .C(_03158_),
    .Y(_03159_));
 sg13g2_nor2b_1 _11015_ (.A(net3944),
    .B_N(\mem.mem[24][2] ),
    .Y(_03160_));
 sg13g2_a21oi_1 _11016_ (.A1(net3944),
    .A2(\mem.mem[25][2] ),
    .Y(_03161_),
    .B1(_03160_));
 sg13g2_nand2b_1 _11017_ (.Y(_03162_),
    .B(\mem.mem[26][2] ),
    .A_N(net3944));
 sg13g2_a21oi_1 _11018_ (.A1(net3944),
    .A2(\mem.mem[27][2] ),
    .Y(_03163_),
    .B1(net3223));
 sg13g2_a221oi_1 _11019_ (.B2(_03163_),
    .C1(net3684),
    .B1(_03162_),
    .A1(net3223),
    .Y(_03164_),
    .A2(_03161_));
 sg13g2_nand2b_1 _11020_ (.Y(_03165_),
    .B(\mem.mem[28][2] ),
    .A_N(net3929));
 sg13g2_a21oi_1 _11021_ (.A1(net3929),
    .A2(\mem.mem[29][2] ),
    .Y(_03166_),
    .B1(net3751));
 sg13g2_nor2b_1 _11022_ (.A(net3934),
    .B_N(\mem.mem[30][2] ),
    .Y(_03167_));
 sg13g2_a21oi_1 _11023_ (.A1(net3929),
    .A2(\mem.mem[31][2] ),
    .Y(_03168_),
    .B1(_03167_));
 sg13g2_a221oi_1 _11024_ (.B2(net3751),
    .C1(net3160),
    .B1(_03168_),
    .A1(_03165_),
    .Y(_03169_),
    .A2(_03166_));
 sg13g2_nor3_1 _11025_ (.A(net3117),
    .B(_03164_),
    .C(_03169_),
    .Y(_03170_));
 sg13g2_o21ai_1 _11026_ (.B1(net3626),
    .Y(_03171_),
    .A1(_03159_),
    .A2(_03170_));
 sg13g2_nand3_1 _11027_ (.B(_03148_),
    .C(_03171_),
    .A(net3093),
    .Y(_03172_));
 sg13g2_a21oi_1 _11028_ (.A1(net3936),
    .A2(\mem.mem[39][2] ),
    .Y(_03173_),
    .B1(net3226));
 sg13g2_o21ai_1 _11029_ (.B1(_03173_),
    .Y(_03174_),
    .A1(net3936),
    .A2(_02153_));
 sg13g2_nand2b_1 _11030_ (.Y(_03175_),
    .B(\mem.mem[36][2] ),
    .A_N(net3945));
 sg13g2_a21oi_1 _11031_ (.A1(net3945),
    .A2(\mem.mem[37][2] ),
    .Y(_03176_),
    .B1(net3757));
 sg13g2_a21oi_1 _11032_ (.A1(_03175_),
    .A2(_03176_),
    .Y(_03177_),
    .B1(net3162));
 sg13g2_mux4_1 _11033_ (.S0(net3932),
    .A0(\mem.mem[32][2] ),
    .A1(\mem.mem[33][2] ),
    .A2(\mem.mem[34][2] ),
    .A3(\mem.mem[35][2] ),
    .S1(net3753),
    .X(_03178_));
 sg13g2_a221oi_1 _11034_ (.B2(net3160),
    .C1(net3649),
    .B1(_03178_),
    .A1(_03174_),
    .Y(_03179_),
    .A2(_03177_));
 sg13g2_nor2b_1 _11035_ (.A(net3979),
    .B_N(\mem.mem[40][2] ),
    .Y(_03180_));
 sg13g2_a21oi_1 _11036_ (.A1(net3979),
    .A2(\mem.mem[41][2] ),
    .Y(_03181_),
    .B1(_03180_));
 sg13g2_nand2b_1 _11037_ (.Y(_03182_),
    .B(\mem.mem[42][2] ),
    .A_N(net3979));
 sg13g2_a21oi_1 _11038_ (.A1(net3979),
    .A2(\mem.mem[43][2] ),
    .Y(_03183_),
    .B1(net3233));
 sg13g2_a221oi_1 _11039_ (.B2(_03183_),
    .C1(net3689),
    .B1(_03182_),
    .A1(net3233),
    .Y(_03184_),
    .A2(_03181_));
 sg13g2_nand2b_1 _11040_ (.Y(_03185_),
    .B(\mem.mem[44][2] ),
    .A_N(net3959));
 sg13g2_a21oi_1 _11041_ (.A1(net3974),
    .A2(\mem.mem[45][2] ),
    .Y(_03186_),
    .B1(net3760));
 sg13g2_nor2b_1 _11042_ (.A(net3959),
    .B_N(\mem.mem[46][2] ),
    .Y(_03187_));
 sg13g2_a21oi_1 _11043_ (.A1(net3959),
    .A2(\mem.mem[47][2] ),
    .Y(_03188_),
    .B1(_03187_));
 sg13g2_a221oi_1 _11044_ (.B2(net3760),
    .C1(net3169),
    .B1(_03188_),
    .A1(_03185_),
    .Y(_03189_),
    .A2(_03186_));
 sg13g2_nor3_1 _11045_ (.A(net3118),
    .B(_03184_),
    .C(_03189_),
    .Y(_03190_));
 sg13g2_o21ai_1 _11046_ (.B1(net3099),
    .Y(_03191_),
    .A1(_03179_),
    .A2(_03190_));
 sg13g2_nor2b_1 _11047_ (.A(net3968),
    .B_N(\mem.mem[52][2] ),
    .Y(_03192_));
 sg13g2_a21oi_1 _11048_ (.A1(net3962),
    .A2(\mem.mem[53][2] ),
    .Y(_03193_),
    .B1(_03192_));
 sg13g2_nand2b_1 _11049_ (.Y(_03194_),
    .B(\mem.mem[54][2] ),
    .A_N(net3961));
 sg13g2_a21oi_1 _11050_ (.A1(net3961),
    .A2(\mem.mem[55][2] ),
    .Y(_03195_),
    .B1(net3228));
 sg13g2_a221oi_1 _11051_ (.B2(_03195_),
    .C1(net3166),
    .B1(_03194_),
    .A1(net3228),
    .Y(_03196_),
    .A2(_03193_));
 sg13g2_mux2_1 _11052_ (.A0(\mem.mem[48][2] ),
    .A1(\mem.mem[49][2] ),
    .S(net3957),
    .X(_03197_));
 sg13g2_nor2_1 _11053_ (.A(net3760),
    .B(_03197_),
    .Y(_03198_));
 sg13g2_mux2_1 _11054_ (.A0(\mem.mem[50][2] ),
    .A1(\mem.mem[51][2] ),
    .S(net3957),
    .X(_03199_));
 sg13g2_o21ai_1 _11055_ (.B1(net3166),
    .Y(_03200_),
    .A1(net3228),
    .A2(_03199_));
 sg13g2_o21ai_1 _11056_ (.B1(net3119),
    .Y(_03201_),
    .A1(_03198_),
    .A2(_03200_));
 sg13g2_mux4_1 _11057_ (.S0(net3978),
    .A0(\mem.mem[56][2] ),
    .A1(\mem.mem[57][2] ),
    .A2(\mem.mem[58][2] ),
    .A3(\mem.mem[59][2] ),
    .S1(net3765),
    .X(_03202_));
 sg13g2_mux2_1 _11058_ (.A0(\mem.mem[62][2] ),
    .A1(\mem.mem[63][2] ),
    .S(net3984),
    .X(_03203_));
 sg13g2_nor2_1 _11059_ (.A(net3235),
    .B(_03203_),
    .Y(_03204_));
 sg13g2_mux2_1 _11060_ (.A0(\mem.mem[60][2] ),
    .A1(\mem.mem[61][2] ),
    .S(net3984),
    .X(_03205_));
 sg13g2_o21ai_1 _11061_ (.B1(net3688),
    .Y(_03206_),
    .A1(net3767),
    .A2(_03205_));
 sg13g2_a21oi_1 _11062_ (.A1(net3171),
    .A2(_03202_),
    .Y(_03207_),
    .B1(net3118));
 sg13g2_o21ai_1 _11063_ (.B1(_03207_),
    .Y(_03208_),
    .A1(_03204_),
    .A2(_03206_));
 sg13g2_o21ai_1 _11064_ (.B1(_03208_),
    .Y(_03209_),
    .A1(_03196_),
    .A2(_03201_));
 sg13g2_a21oi_1 _11065_ (.A1(net3630),
    .A2(_03209_),
    .Y(_03210_),
    .B1(net3092));
 sg13g2_a21oi_2 _11066_ (.B1(net3614),
    .Y(_03211_),
    .A2(_03210_),
    .A1(_03191_));
 sg13g2_mux4_1 _11067_ (.S0(net3814),
    .A0(\mem.mem[84][2] ),
    .A1(\mem.mem[85][2] ),
    .A2(\mem.mem[86][2] ),
    .A3(\mem.mem[87][2] ),
    .S1(net3710),
    .X(_03212_));
 sg13g2_nand2_1 _11068_ (.Y(_03213_),
    .A(net3663),
    .B(_03212_));
 sg13g2_mux4_1 _11069_ (.S0(net3803),
    .A0(\mem.mem[80][2] ),
    .A1(\mem.mem[81][2] ),
    .A2(\mem.mem[82][2] ),
    .A3(\mem.mem[83][2] ),
    .S1(net3705),
    .X(_03214_));
 sg13g2_mux4_1 _11070_ (.S0(net3806),
    .A0(\mem.mem[92][2] ),
    .A1(\mem.mem[93][2] ),
    .A2(\mem.mem[94][2] ),
    .A3(\mem.mem[95][2] ),
    .S1(net3706),
    .X(_03215_));
 sg13g2_nand2_1 _11071_ (.Y(_03216_),
    .A(net3663),
    .B(_03215_));
 sg13g2_mux4_1 _11072_ (.S0(net3803),
    .A0(\mem.mem[88][2] ),
    .A1(\mem.mem[89][2] ),
    .A2(\mem.mem[90][2] ),
    .A3(\mem.mem[91][2] ),
    .S1(net3705),
    .X(_03217_));
 sg13g2_mux4_1 _11073_ (.S0(net3808),
    .A0(\mem.mem[68][2] ),
    .A1(\mem.mem[69][2] ),
    .A2(\mem.mem[70][2] ),
    .A3(\mem.mem[71][2] ),
    .S1(net3708),
    .X(_03218_));
 sg13g2_mux4_1 _11074_ (.S0(net3791),
    .A0(\mem.mem[64][2] ),
    .A1(\mem.mem[65][2] ),
    .A2(\mem.mem[66][2] ),
    .A3(\mem.mem[67][2] ),
    .S1(net3698),
    .X(_03219_));
 sg13g2_nand2_1 _11075_ (.Y(_03220_),
    .A(net3123),
    .B(_03219_));
 sg13g2_a21oi_1 _11076_ (.A1(net3664),
    .A2(_03218_),
    .Y(_03221_),
    .B1(net3636));
 sg13g2_nor2b_1 _11077_ (.A(net3797),
    .B_N(\mem.mem[78][2] ),
    .Y(_03222_));
 sg13g2_a21oi_1 _11078_ (.A1(net3797),
    .A2(\mem.mem[79][2] ),
    .Y(_03223_),
    .B1(_03222_));
 sg13g2_mux2_1 _11079_ (.A0(\mem.mem[76][2] ),
    .A1(\mem.mem[77][2] ),
    .S(net3797),
    .X(_03224_));
 sg13g2_o21ai_1 _11080_ (.B1(net3661),
    .Y(_03225_),
    .A1(net3702),
    .A2(_03224_));
 sg13g2_a21o_1 _11081_ (.A2(_03223_),
    .A1(net3702),
    .B1(_03225_),
    .X(_03226_));
 sg13g2_mux4_1 _11082_ (.S0(net3781),
    .A0(\mem.mem[72][2] ),
    .A1(\mem.mem[73][2] ),
    .A2(\mem.mem[74][2] ),
    .A3(\mem.mem[75][2] ),
    .S1(net3695),
    .X(_03227_));
 sg13g2_a21oi_2 _11083_ (.B1(net3101),
    .Y(_03228_),
    .A2(_03227_),
    .A1(net3123));
 sg13g2_a221oi_1 _11084_ (.B2(_03228_),
    .C1(net3620),
    .B1(_03226_),
    .A1(_03220_),
    .Y(_03229_),
    .A2(_03221_));
 sg13g2_a21oi_1 _11085_ (.A1(net3129),
    .A2(_03214_),
    .Y(_03230_),
    .B1(net3635));
 sg13g2_a21oi_1 _11086_ (.A1(net3129),
    .A2(_03217_),
    .Y(_03231_),
    .B1(net3104));
 sg13g2_a221oi_1 _11087_ (.B2(_03216_),
    .C1(net3094),
    .B1(_03231_),
    .A1(_03213_),
    .Y(_03232_),
    .A2(_03230_));
 sg13g2_o21ai_1 _11088_ (.B1(net3091),
    .Y(_03233_),
    .A1(_03229_),
    .A2(_03232_));
 sg13g2_a21oi_1 _11089_ (.A1(net3908),
    .A2(\mem.mem[103][2] ),
    .Y(_03234_),
    .B1(net3213));
 sg13g2_o21ai_1 _11090_ (.B1(_03234_),
    .Y(_03235_),
    .A1(net3908),
    .A2(_02154_));
 sg13g2_nand2b_1 _11091_ (.Y(_03236_),
    .B(\mem.mem[100][2] ),
    .A_N(net3916));
 sg13g2_a21oi_1 _11092_ (.A1(net3919),
    .A2(\mem.mem[101][2] ),
    .Y(_03237_),
    .B1(net3748));
 sg13g2_a21oi_1 _11093_ (.A1(_03236_),
    .A2(_03237_),
    .Y(_03238_),
    .B1(net3158));
 sg13g2_mux4_1 _11094_ (.S0(net3915),
    .A0(\mem.mem[96][2] ),
    .A1(\mem.mem[97][2] ),
    .A2(\mem.mem[98][2] ),
    .A3(\mem.mem[99][2] ),
    .S1(net3748),
    .X(_03239_));
 sg13g2_a221oi_1 _11095_ (.B2(net3158),
    .C1(net3647),
    .B1(_03239_),
    .A1(_03235_),
    .Y(_03240_),
    .A2(_03238_));
 sg13g2_nor2b_1 _11096_ (.A(net3905),
    .B_N(\mem.mem[104][2] ),
    .Y(_03241_));
 sg13g2_a21oi_1 _11097_ (.A1(net3905),
    .A2(\mem.mem[105][2] ),
    .Y(_03242_),
    .B1(_03241_));
 sg13g2_nand2b_1 _11098_ (.Y(_03243_),
    .B(\mem.mem[106][2] ),
    .A_N(net3905));
 sg13g2_a21oi_1 _11099_ (.A1(net3905),
    .A2(\mem.mem[107][2] ),
    .Y(_03244_),
    .B1(net3215));
 sg13g2_a221oi_1 _11100_ (.B2(_03244_),
    .C1(net3680),
    .B1(_03243_),
    .A1(net3215),
    .Y(_03245_),
    .A2(_03242_));
 sg13g2_nand2b_1 _11101_ (.Y(_03246_),
    .B(\mem.mem[108][2] ),
    .A_N(net3904));
 sg13g2_a21oi_1 _11102_ (.A1(net3904),
    .A2(\mem.mem[109][2] ),
    .Y(_03247_),
    .B1(net3744));
 sg13g2_nor2b_1 _11103_ (.A(net3904),
    .B_N(\mem.mem[110][2] ),
    .Y(_03248_));
 sg13g2_a21oi_1 _11104_ (.A1(net3904),
    .A2(\mem.mem[111][2] ),
    .Y(_03249_),
    .B1(_03248_));
 sg13g2_a221oi_1 _11105_ (.B2(net3744),
    .C1(net3154),
    .B1(_03249_),
    .A1(_03246_),
    .Y(_03250_),
    .A2(_03247_));
 sg13g2_nor3_2 _11106_ (.A(net3112),
    .B(_03245_),
    .C(_03250_),
    .Y(_03251_));
 sg13g2_o21ai_1 _11107_ (.B1(net3100),
    .Y(_03252_),
    .A1(_03240_),
    .A2(_03251_));
 sg13g2_nor2b_1 _11108_ (.A(net3820),
    .B_N(\mem.mem[116][2] ),
    .Y(_03253_));
 sg13g2_a21oi_1 _11109_ (.A1(net3820),
    .A2(\mem.mem[117][2] ),
    .Y(_03254_),
    .B1(_03253_));
 sg13g2_nand2b_1 _11110_ (.Y(_03255_),
    .B(\mem.mem[118][2] ),
    .A_N(net3820));
 sg13g2_a21oi_1 _11111_ (.A1(net3824),
    .A2(\mem.mem[119][2] ),
    .Y(_03256_),
    .B1(net3187));
 sg13g2_a221oi_1 _11112_ (.B2(_03256_),
    .C1(net3134),
    .B1(_03255_),
    .A1(net3187),
    .Y(_03257_),
    .A2(_03254_));
 sg13g2_nor2b_1 _11113_ (.A(net3834),
    .B_N(\mem.mem[112][2] ),
    .Y(_03258_));
 sg13g2_a21oi_1 _11114_ (.A1(net3834),
    .A2(\mem.mem[113][2] ),
    .Y(_03259_),
    .B1(_03258_));
 sg13g2_nand2b_1 _11115_ (.Y(_03260_),
    .B(\mem.mem[114][2] ),
    .A_N(net3834));
 sg13g2_a21oi_1 _11116_ (.A1(net3834),
    .A2(\mem.mem[115][2] ),
    .Y(_03261_),
    .B1(net3191));
 sg13g2_a221oi_1 _11117_ (.B2(_03261_),
    .C1(net3669),
    .B1(_03260_),
    .A1(net3191),
    .Y(_03262_),
    .A2(_03259_));
 sg13g2_nor3_2 _11118_ (.A(net3639),
    .B(_03257_),
    .C(_03262_),
    .Y(_03263_));
 sg13g2_nor2b_1 _11119_ (.A(net3841),
    .B_N(\mem.mem[120][2] ),
    .Y(_03264_));
 sg13g2_a21oi_1 _11120_ (.A1(net3841),
    .A2(\mem.mem[121][2] ),
    .Y(_03265_),
    .B1(_03264_));
 sg13g2_nand2b_1 _11121_ (.Y(_03266_),
    .B(\mem.mem[122][2] ),
    .A_N(net3841));
 sg13g2_a21oi_1 _11122_ (.A1(net3841),
    .A2(\mem.mem[123][2] ),
    .Y(_03267_),
    .B1(net3192));
 sg13g2_a221oi_1 _11123_ (.B2(_03267_),
    .C1(net3671),
    .B1(_03266_),
    .A1(net3192),
    .Y(_03268_),
    .A2(_03265_));
 sg13g2_nor2b_1 _11124_ (.A(net3849),
    .B_N(\mem.mem[126][2] ),
    .Y(_03269_));
 sg13g2_a21oi_1 _11125_ (.A1(net3849),
    .A2(\mem.mem[127][2] ),
    .Y(_03270_),
    .B1(_03269_));
 sg13g2_nand2b_1 _11126_ (.Y(_03271_),
    .B(\mem.mem[124][2] ),
    .A_N(net3849));
 sg13g2_a21oi_1 _11127_ (.A1(net3849),
    .A2(\mem.mem[125][2] ),
    .Y(_03272_),
    .B1(net3725));
 sg13g2_a221oi_1 _11128_ (.B2(_03272_),
    .C1(net3139),
    .B1(_03271_),
    .A1(net3725),
    .Y(_03273_),
    .A2(_03270_));
 sg13g2_nor3_1 _11129_ (.A(net3109),
    .B(_03268_),
    .C(_03273_),
    .Y(_03274_));
 sg13g2_o21ai_1 _11130_ (.B1(net3624),
    .Y(_03275_),
    .A1(_03263_),
    .A2(_03274_));
 sg13g2_nand3_1 _11131_ (.B(_03252_),
    .C(_03275_),
    .A(net3617),
    .Y(_03276_));
 sg13g2_and2_1 _11132_ (.A(net3613),
    .B(_03233_),
    .X(_03277_));
 sg13g2_a22oi_1 _11133_ (.Y(_03278_),
    .B1(_03276_),
    .B2(_03277_),
    .A2(_03211_),
    .A1(_03172_));
 sg13g2_nand2b_1 _11134_ (.Y(_03279_),
    .B(net3880),
    .A_N(\mem.mem[229][2] ));
 sg13g2_o21ai_1 _11135_ (.B1(_03279_),
    .Y(_03280_),
    .A1(net3880),
    .A2(\mem.mem[228][2] ));
 sg13g2_mux2_1 _11136_ (.A0(\mem.mem[230][2] ),
    .A1(\mem.mem[231][2] ),
    .S(net3868),
    .X(_03281_));
 sg13g2_o21ai_1 _11137_ (.B1(net3675),
    .Y(_03282_),
    .A1(net3204),
    .A2(_03281_));
 sg13g2_a21o_1 _11138_ (.A2(_03280_),
    .A1(net3204),
    .B1(_03282_),
    .X(_03283_));
 sg13g2_mux4_1 _11139_ (.S0(net3865),
    .A0(\mem.mem[224][2] ),
    .A1(\mem.mem[225][2] ),
    .A2(\mem.mem[226][2] ),
    .A3(\mem.mem[227][2] ),
    .S1(net3733),
    .X(_03284_));
 sg13g2_a21oi_1 _11140_ (.A1(net3148),
    .A2(_03284_),
    .Y(_03285_),
    .B1(net3643));
 sg13g2_mux4_1 _11141_ (.S0(net3866),
    .A0(\mem.mem[236][2] ),
    .A1(\mem.mem[237][2] ),
    .A2(\mem.mem[238][2] ),
    .A3(\mem.mem[239][2] ),
    .S1(net3733),
    .X(_03286_));
 sg13g2_nor2b_1 _11142_ (.A(net3864),
    .B_N(\mem.mem[234][2] ),
    .Y(_03287_));
 sg13g2_a21oi_1 _11143_ (.A1(net3864),
    .A2(\mem.mem[235][2] ),
    .Y(_03288_),
    .B1(_03287_));
 sg13g2_nand2_1 _11144_ (.Y(_03289_),
    .A(net3865),
    .B(\mem.mem[233][2] ));
 sg13g2_nand2b_1 _11145_ (.Y(_03290_),
    .B(\mem.mem[232][2] ),
    .A_N(net3864));
 sg13g2_nand3_1 _11146_ (.B(_03289_),
    .C(_03290_),
    .A(net3201),
    .Y(_03291_));
 sg13g2_a21oi_1 _11147_ (.A1(net3733),
    .A2(_03288_),
    .Y(_03292_),
    .B1(net3674));
 sg13g2_a221oi_1 _11148_ (.B2(_03292_),
    .C1(net3111),
    .B1(_03291_),
    .A1(net3674),
    .Y(_03293_),
    .A2(_03286_));
 sg13g2_a21oi_2 _11149_ (.B1(_03293_),
    .Y(_03294_),
    .A2(_03285_),
    .A1(_03283_));
 sg13g2_nand2b_1 _11150_ (.Y(_03295_),
    .B(\mem.mem[246][2] ),
    .A_N(net3817));
 sg13g2_a21oi_1 _11151_ (.A1(net3817),
    .A2(\mem.mem[247][2] ),
    .Y(_03296_),
    .B1(net3189));
 sg13g2_nor2b_1 _11152_ (.A(net3817),
    .B_N(\mem.mem[244][2] ),
    .Y(_03297_));
 sg13g2_a21oi_1 _11153_ (.A1(net3816),
    .A2(\mem.mem[245][2] ),
    .Y(_03298_),
    .B1(_03297_));
 sg13g2_a221oi_1 _11154_ (.B2(net3189),
    .C1(net3133),
    .B1(_03298_),
    .A1(_03295_),
    .Y(_03299_),
    .A2(_03296_));
 sg13g2_mux4_1 _11155_ (.S0(net3817),
    .A0(\mem.mem[240][2] ),
    .A1(\mem.mem[241][2] ),
    .A2(\mem.mem[242][2] ),
    .A3(\mem.mem[243][2] ),
    .S1(net3712),
    .X(_03300_));
 sg13g2_a21oi_1 _11156_ (.A1(net3133),
    .A2(_03300_),
    .Y(_03301_),
    .B1(_03299_));
 sg13g2_mux4_1 _11157_ (.S0(net3823),
    .A0(\mem.mem[248][2] ),
    .A1(\mem.mem[249][2] ),
    .A2(\mem.mem[250][2] ),
    .A3(\mem.mem[251][2] ),
    .S1(net3714),
    .X(_03302_));
 sg13g2_nand2_1 _11158_ (.Y(_03303_),
    .A(net3133),
    .B(_03302_));
 sg13g2_a21oi_1 _11159_ (.A1(net3667),
    .A2(\mem.mem[252][2] ),
    .Y(_03304_),
    .B1(net3106));
 sg13g2_a22oi_1 _11160_ (.Y(_03305_),
    .B1(_03303_),
    .B2(_03304_),
    .A2(_03301_),
    .A1(net3106));
 sg13g2_mux4_1 _11161_ (.S0(net3774),
    .A0(\mem.mem[196][2] ),
    .A1(\mem.mem[197][2] ),
    .A2(\mem.mem[198][2] ),
    .A3(\mem.mem[199][2] ),
    .S1(net3692),
    .X(_03306_));
 sg13g2_mux4_1 _11162_ (.S0(net3772),
    .A0(\mem.mem[192][2] ),
    .A1(\mem.mem[193][2] ),
    .A2(\mem.mem[194][2] ),
    .A3(\mem.mem[195][2] ),
    .S1(net3692),
    .X(_03307_));
 sg13g2_nand2_1 _11163_ (.Y(_03308_),
    .A(net3121),
    .B(_03307_));
 sg13g2_a21oi_1 _11164_ (.A1(net3657),
    .A2(_03306_),
    .Y(_03309_),
    .B1(net3632));
 sg13g2_nor2b_1 _11165_ (.A(net3778),
    .B_N(\mem.mem[206][2] ),
    .Y(_03310_));
 sg13g2_a21oi_1 _11166_ (.A1(net3778),
    .A2(\mem.mem[207][2] ),
    .Y(_03311_),
    .B1(_03310_));
 sg13g2_mux2_1 _11167_ (.A0(\mem.mem[204][2] ),
    .A1(\mem.mem[205][2] ),
    .S(net3777),
    .X(_03312_));
 sg13g2_a21oi_1 _11168_ (.A1(net3693),
    .A2(_03311_),
    .Y(_03313_),
    .B1(net3123));
 sg13g2_o21ai_1 _11169_ (.B1(_03313_),
    .Y(_03314_),
    .A1(net3693),
    .A2(_03312_));
 sg13g2_mux4_1 _11170_ (.S0(net3773),
    .A0(\mem.mem[200][2] ),
    .A1(\mem.mem[201][2] ),
    .A2(\mem.mem[202][2] ),
    .A3(\mem.mem[203][2] ),
    .S1(net3692),
    .X(_03315_));
 sg13g2_a21oi_1 _11171_ (.A1(net3121),
    .A2(_03315_),
    .Y(_03316_),
    .B1(net3101));
 sg13g2_a22oi_1 _11172_ (.Y(_03317_),
    .B1(_03314_),
    .B2(_03316_),
    .A2(_03309_),
    .A1(_03308_));
 sg13g2_nand2b_1 _11173_ (.Y(_03318_),
    .B(\mem.mem[222][2] ),
    .A_N(net3819));
 sg13g2_a21oi_1 _11174_ (.A1(net3818),
    .A2(\mem.mem[223][2] ),
    .Y(_03319_),
    .B1(net3189));
 sg13g2_nor2b_1 _11175_ (.A(net3818),
    .B_N(\mem.mem[220][2] ),
    .Y(_03320_));
 sg13g2_a21oi_1 _11176_ (.A1(net3818),
    .A2(\mem.mem[221][2] ),
    .Y(_03321_),
    .B1(_03320_));
 sg13g2_a221oi_1 _11177_ (.B2(net3189),
    .C1(net3126),
    .B1(_03321_),
    .A1(_03318_),
    .Y(_03322_),
    .A2(_03319_));
 sg13g2_nor2b_1 _11178_ (.A(net3816),
    .B_N(\mem.mem[218][2] ),
    .Y(_03323_));
 sg13g2_a21oi_1 _11179_ (.A1(net3816),
    .A2(\mem.mem[219][2] ),
    .Y(_03324_),
    .B1(_03323_));
 sg13g2_mux2_1 _11180_ (.A0(\mem.mem[216][2] ),
    .A1(\mem.mem[217][2] ),
    .S(net3816),
    .X(_03325_));
 sg13g2_o21ai_1 _11181_ (.B1(net3126),
    .Y(_03326_),
    .A1(net3712),
    .A2(_03325_));
 sg13g2_a21oi_1 _11182_ (.A1(net3712),
    .A2(_03324_),
    .Y(_03327_),
    .B1(_03326_));
 sg13g2_nor3_1 _11183_ (.A(net3102),
    .B(_03322_),
    .C(_03327_),
    .Y(_03328_));
 sg13g2_nor2b_1 _11184_ (.A(net3783),
    .B_N(\mem.mem[210][2] ),
    .Y(_03329_));
 sg13g2_a21oi_1 _11185_ (.A1(net3783),
    .A2(\mem.mem[211][2] ),
    .Y(_03330_),
    .B1(_03329_));
 sg13g2_mux2_1 _11186_ (.A0(\mem.mem[208][2] ),
    .A1(\mem.mem[209][2] ),
    .S(net3786),
    .X(_03331_));
 sg13g2_o21ai_1 _11187_ (.B1(net3125),
    .Y(_03332_),
    .A1(net3697),
    .A2(_03331_));
 sg13g2_a21oi_2 _11188_ (.B1(_03332_),
    .Y(_03333_),
    .A2(_03330_),
    .A1(net3697));
 sg13g2_nand2b_1 _11189_ (.Y(_03334_),
    .B(\mem.mem[214][2] ),
    .A_N(net3793));
 sg13g2_a21oi_1 _11190_ (.A1(net3794),
    .A2(\mem.mem[215][2] ),
    .Y(_03335_),
    .B1(net3180));
 sg13g2_nand2b_1 _11191_ (.Y(_03336_),
    .B(net3793),
    .A_N(\mem.mem[213][2] ));
 sg13g2_o21ai_1 _11192_ (.B1(_03336_),
    .Y(_03337_),
    .A1(net3794),
    .A2(\mem.mem[212][2] ));
 sg13g2_a221oi_1 _11193_ (.B2(net3180),
    .C1(net3127),
    .B1(_03337_),
    .A1(_03334_),
    .Y(_03338_),
    .A2(_03335_));
 sg13g2_nor3_1 _11194_ (.A(net3637),
    .B(_03333_),
    .C(_03338_),
    .Y(_03339_));
 sg13g2_nor2_1 _11195_ (.A(_03328_),
    .B(_03339_),
    .Y(_03340_));
 sg13g2_mux4_1 _11196_ (.S0(net3623),
    .A0(_03294_),
    .A1(_03305_),
    .A2(_03317_),
    .A3(_03340_),
    .S1(net3090),
    .X(_03341_));
 sg13g2_and2_1 _11197_ (.A(net3613),
    .B(_03341_),
    .X(_03342_));
 sg13g2_nor2b_1 _11198_ (.A(\mem.mem[167][2] ),
    .B_N(net3875),
    .Y(_03343_));
 sg13g2_o21ai_1 _11199_ (.B1(net3735),
    .Y(_03344_),
    .A1(net3875),
    .A2(\mem.mem[166][2] ));
 sg13g2_mux2_1 _11200_ (.A0(\mem.mem[164][2] ),
    .A1(\mem.mem[165][2] ),
    .S(net3875),
    .X(_03345_));
 sg13g2_o21ai_1 _11201_ (.B1(net3676),
    .Y(_03346_),
    .A1(_03343_),
    .A2(_03344_));
 sg13g2_a21oi_1 _11202_ (.A1(net3202),
    .A2(_03345_),
    .Y(_03347_),
    .B1(_03346_));
 sg13g2_mux2_1 _11203_ (.A0(\mem.mem[162][2] ),
    .A1(\mem.mem[163][2] ),
    .S(net3872),
    .X(_03348_));
 sg13g2_nand2b_1 _11204_ (.Y(_03349_),
    .B(net3872),
    .A_N(\mem.mem[161][2] ));
 sg13g2_nor2_1 _11205_ (.A(net3872),
    .B(\mem.mem[160][2] ),
    .Y(_03350_));
 sg13g2_nor2_1 _11206_ (.A(net3734),
    .B(_03350_),
    .Y(_03351_));
 sg13g2_a221oi_1 _11207_ (.B2(_03351_),
    .C1(net3675),
    .B1(_03349_),
    .A1(net3734),
    .Y(_03352_),
    .A2(_03348_));
 sg13g2_or3_1 _11208_ (.A(net3643),
    .B(_03347_),
    .C(_03352_),
    .X(_03353_));
 sg13g2_mux4_1 _11209_ (.S0(net3849),
    .A0(\mem.mem[168][2] ),
    .A1(\mem.mem[169][2] ),
    .A2(\mem.mem[170][2] ),
    .A3(\mem.mem[171][2] ),
    .S1(net3725),
    .X(_03354_));
 sg13g2_mux2_1 _11210_ (.A0(\mem.mem[172][2] ),
    .A1(\mem.mem[173][2] ),
    .S(net3834),
    .X(_03355_));
 sg13g2_nand2_1 _11211_ (.Y(_03356_),
    .A(net3191),
    .B(_03355_));
 sg13g2_mux2_1 _11212_ (.A0(\mem.mem[174][2] ),
    .A1(\mem.mem[175][2] ),
    .S(net3833),
    .X(_03357_));
 sg13g2_a21oi_1 _11213_ (.A1(net3719),
    .A2(_03357_),
    .Y(_03358_),
    .B1(net3137));
 sg13g2_a21oi_1 _11214_ (.A1(_03356_),
    .A2(_03358_),
    .Y(_03359_),
    .B1(net3107));
 sg13g2_o21ai_1 _11215_ (.B1(_03359_),
    .Y(_03360_),
    .A1(net3669),
    .A2(_03354_));
 sg13g2_nand3_1 _11216_ (.B(_03353_),
    .C(_03360_),
    .A(net3095),
    .Y(_03361_));
 sg13g2_mux2_1 _11217_ (.A0(\mem.mem[182][2] ),
    .A1(\mem.mem[183][2] ),
    .S(net3854),
    .X(_03362_));
 sg13g2_nand2_1 _11218_ (.Y(_03363_),
    .A(net3727),
    .B(_03362_));
 sg13g2_mux2_1 _11219_ (.A0(\mem.mem[180][2] ),
    .A1(\mem.mem[181][2] ),
    .S(net3860),
    .X(_03364_));
 sg13g2_a21oi_1 _11220_ (.A1(net3194),
    .A2(_03364_),
    .Y(_03365_),
    .B1(net3143));
 sg13g2_mux2_1 _11221_ (.A0(\mem.mem[178][2] ),
    .A1(\mem.mem[179][2] ),
    .S(net3854),
    .X(_03366_));
 sg13g2_nand2_1 _11222_ (.Y(_03367_),
    .A(net3727),
    .B(_03366_));
 sg13g2_mux2_1 _11223_ (.A0(\mem.mem[176][2] ),
    .A1(\mem.mem[177][2] ),
    .S(net3856),
    .X(_03368_));
 sg13g2_a21oi_1 _11224_ (.A1(net3193),
    .A2(_03368_),
    .Y(_03369_),
    .B1(net3672));
 sg13g2_a221oi_1 _11225_ (.B2(_03369_),
    .C1(net3640),
    .B1(_03367_),
    .A1(_03363_),
    .Y(_03370_),
    .A2(_03365_));
 sg13g2_mux4_1 _11226_ (.S0(net3848),
    .A0(\mem.mem[184][2] ),
    .A1(\mem.mem[185][2] ),
    .A2(\mem.mem[186][2] ),
    .A3(\mem.mem[187][2] ),
    .S1(net3724),
    .X(_03371_));
 sg13g2_mux2_1 _11227_ (.A0(\mem.mem[188][2] ),
    .A1(\mem.mem[189][2] ),
    .S(net3846),
    .X(_03372_));
 sg13g2_nand2_1 _11228_ (.Y(_03373_),
    .A(net3197),
    .B(_03372_));
 sg13g2_mux2_1 _11229_ (.A0(\mem.mem[190][2] ),
    .A1(\mem.mem[191][2] ),
    .S(net3846),
    .X(_03374_));
 sg13g2_a21oi_1 _11230_ (.A1(net3723),
    .A2(_03374_),
    .Y(_03375_),
    .B1(net3140));
 sg13g2_a21oi_1 _11231_ (.A1(_03373_),
    .A2(_03375_),
    .Y(_03376_),
    .B1(net3109));
 sg13g2_o21ai_1 _11232_ (.B1(_03376_),
    .Y(_03377_),
    .A1(net3671),
    .A2(_03371_));
 sg13g2_nand3b_1 _11233_ (.B(_03377_),
    .C(net3622),
    .Y(_03378_),
    .A_N(_03370_));
 sg13g2_nand3_1 _11234_ (.B(_03361_),
    .C(_03378_),
    .A(net3616),
    .Y(_03379_));
 sg13g2_a21oi_1 _11235_ (.A1(net3890),
    .A2(\mem.mem[133][2] ),
    .Y(_03380_),
    .B1(net3739));
 sg13g2_o21ai_1 _11236_ (.B1(_03380_),
    .Y(_03381_),
    .A1(net3890),
    .A2(_02155_));
 sg13g2_nor2b_1 _11237_ (.A(net3891),
    .B_N(\mem.mem[134][2] ),
    .Y(_03382_));
 sg13g2_a21oi_1 _11238_ (.A1(net3891),
    .A2(\mem.mem[135][2] ),
    .Y(_03383_),
    .B1(_03382_));
 sg13g2_a21oi_1 _11239_ (.A1(net3740),
    .A2(_03383_),
    .Y(_03384_),
    .B1(net3152));
 sg13g2_mux4_1 _11240_ (.S0(net3886),
    .A0(\mem.mem[128][2] ),
    .A1(\mem.mem[129][2] ),
    .A2(\mem.mem[130][2] ),
    .A3(\mem.mem[131][2] ),
    .S1(net3740),
    .X(_03385_));
 sg13g2_a221oi_1 _11241_ (.B2(net3152),
    .C1(net3644),
    .B1(_03385_),
    .A1(_03381_),
    .Y(_03386_),
    .A2(_03384_));
 sg13g2_nor2b_1 _11242_ (.A(net3896),
    .B_N(\mem.mem[136][2] ),
    .Y(_03387_));
 sg13g2_a21oi_1 _11243_ (.A1(net3896),
    .A2(\mem.mem[137][2] ),
    .Y(_03388_),
    .B1(_03387_));
 sg13g2_nand2b_1 _11244_ (.Y(_03389_),
    .B(\mem.mem[138][2] ),
    .A_N(net3898));
 sg13g2_a21oi_1 _11245_ (.A1(net3898),
    .A2(\mem.mem[139][2] ),
    .Y(_03390_),
    .B1(net3209));
 sg13g2_a221oi_1 _11246_ (.B2(_03390_),
    .C1(net3677),
    .B1(_03389_),
    .A1(net3209),
    .Y(_03391_),
    .A2(_03388_));
 sg13g2_nor2b_1 _11247_ (.A(net3911),
    .B_N(\mem.mem[142][2] ),
    .Y(_03392_));
 sg13g2_a21oi_1 _11248_ (.A1(net3913),
    .A2(\mem.mem[143][2] ),
    .Y(_03393_),
    .B1(_03392_));
 sg13g2_nand2b_1 _11249_ (.Y(_03394_),
    .B(\mem.mem[140][2] ),
    .A_N(net3913));
 sg13g2_a21oi_1 _11250_ (.A1(net3913),
    .A2(\mem.mem[141][2] ),
    .Y(_03395_),
    .B1(net3747));
 sg13g2_a221oi_1 _11251_ (.B2(_03395_),
    .C1(net3155),
    .B1(_03394_),
    .A1(net3746),
    .Y(_03396_),
    .A2(_03393_));
 sg13g2_nor3_1 _11252_ (.A(net3113),
    .B(_03391_),
    .C(_03396_),
    .Y(_03397_));
 sg13g2_o21ai_1 _11253_ (.B1(net3099),
    .Y(_03398_),
    .A1(_03386_),
    .A2(_03397_));
 sg13g2_nand2b_1 _11254_ (.Y(_03399_),
    .B(\mem.mem[150][2] ),
    .A_N(net3971));
 sg13g2_a21oi_1 _11255_ (.A1(net3971),
    .A2(\mem.mem[151][2] ),
    .Y(_03400_),
    .B1(net3234));
 sg13g2_nor2b_1 _11256_ (.A(net3981),
    .B_N(\mem.mem[148][2] ),
    .Y(_03401_));
 sg13g2_a21oi_1 _11257_ (.A1(net3981),
    .A2(\mem.mem[149][2] ),
    .Y(_03402_),
    .B1(_03401_));
 sg13g2_a221oi_1 _11258_ (.B2(net3236),
    .C1(net3167),
    .B1(_03402_),
    .A1(_03399_),
    .Y(_03403_),
    .A2(_03400_));
 sg13g2_nor2b_1 _11259_ (.A(net3920),
    .B_N(\mem.mem[144][2] ),
    .Y(_03404_));
 sg13g2_a21oi_1 _11260_ (.A1(net3920),
    .A2(\mem.mem[145][2] ),
    .Y(_03405_),
    .B1(_03404_));
 sg13g2_nand2b_1 _11261_ (.Y(_03406_),
    .B(\mem.mem[146][2] ),
    .A_N(net3920));
 sg13g2_a21oi_1 _11262_ (.A1(net3920),
    .A2(\mem.mem[147][2] ),
    .Y(_03407_),
    .B1(net3230));
 sg13g2_a221oi_1 _11263_ (.B2(_03407_),
    .C1(net3687),
    .B1(_03406_),
    .A1(net3230),
    .Y(_03408_),
    .A2(_03405_));
 sg13g2_nor3_1 _11264_ (.A(net3652),
    .B(_03403_),
    .C(_03408_),
    .Y(_03409_));
 sg13g2_nor2b_1 _11265_ (.A(net3986),
    .B_N(\mem.mem[152][2] ),
    .Y(_03410_));
 sg13g2_a21oi_1 _11266_ (.A1(net3986),
    .A2(\mem.mem[153][2] ),
    .Y(_03411_),
    .B1(_03410_));
 sg13g2_nand2b_1 _11267_ (.Y(_03412_),
    .B(\mem.mem[154][2] ),
    .A_N(net3982));
 sg13g2_a21oi_1 _11268_ (.A1(net3982),
    .A2(\mem.mem[155][2] ),
    .Y(_03413_),
    .B1(net3235));
 sg13g2_a221oi_1 _11269_ (.B2(_03413_),
    .C1(net3689),
    .B1(_03412_),
    .A1(net3236),
    .Y(_03414_),
    .A2(_03411_));
 sg13g2_nand2b_1 _11270_ (.Y(_03415_),
    .B(\mem.mem[156][2] ),
    .A_N(net3970));
 sg13g2_a21oi_1 _11271_ (.A1(net3970),
    .A2(\mem.mem[157][2] ),
    .Y(_03416_),
    .B1(net3763));
 sg13g2_nor2b_1 _11272_ (.A(net3969),
    .B_N(\mem.mem[158][2] ),
    .Y(_03417_));
 sg13g2_a21oi_1 _11273_ (.A1(net3970),
    .A2(\mem.mem[159][2] ),
    .Y(_03418_),
    .B1(_03417_));
 sg13g2_a221oi_1 _11274_ (.B2(net3763),
    .C1(net3168),
    .B1(_03418_),
    .A1(_03415_),
    .Y(_03419_),
    .A2(_03416_));
 sg13g2_nor3_2 _11275_ (.A(net3119),
    .B(_03414_),
    .C(_03419_),
    .Y(_03420_));
 sg13g2_o21ai_1 _11276_ (.B1(net3630),
    .Y(_03421_),
    .A1(_03409_),
    .A2(_03420_));
 sg13g2_nand3_1 _11277_ (.B(_03398_),
    .C(_03421_),
    .A(net3093),
    .Y(_03422_));
 sg13g2_a21oi_2 _11278_ (.B1(net3612),
    .Y(_03423_),
    .A2(_03422_),
    .A1(_03379_));
 sg13g2_nor3_1 _11279_ (.A(_02149_),
    .B(_03342_),
    .C(_03423_),
    .Y(_03424_));
 sg13g2_o21ai_1 _11280_ (.B1(_02259_),
    .Y(_03425_),
    .A1(net3611),
    .A2(_03278_));
 sg13g2_o21ai_1 _11281_ (.B1(_03133_),
    .Y(_03426_),
    .A1(_03424_),
    .A2(_03425_));
 sg13g2_o21ai_1 _11282_ (.B1(net4002),
    .Y(_03427_),
    .A1(_02535_),
    .A2(_03426_));
 sg13g2_a21oi_1 _11283_ (.A1(_02142_),
    .A2(_02535_),
    .Y(_00597_),
    .B1(_03427_));
 sg13g2_mux4_1 _11284_ (.S0(net3771),
    .A0(\mem.mem[192][3] ),
    .A1(\mem.mem[193][3] ),
    .A2(\mem.mem[194][3] ),
    .A3(\mem.mem[195][3] ),
    .S1(net3691),
    .X(_03428_));
 sg13g2_nand2_1 _11285_ (.Y(_03429_),
    .A(net3121),
    .B(_03428_));
 sg13g2_mux4_1 _11286_ (.S0(net3772),
    .A0(\mem.mem[196][3] ),
    .A1(\mem.mem[197][3] ),
    .A2(\mem.mem[198][3] ),
    .A3(\mem.mem[199][3] ),
    .S1(net3691),
    .X(_03430_));
 sg13g2_a21oi_1 _11287_ (.A1(net3657),
    .A2(_03430_),
    .Y(_03431_),
    .B1(net3632));
 sg13g2_mux4_1 _11288_ (.S0(net3772),
    .A0(\mem.mem[200][3] ),
    .A1(\mem.mem[201][3] ),
    .A2(\mem.mem[202][3] ),
    .A3(\mem.mem[203][3] ),
    .S1(net3691),
    .X(_03432_));
 sg13g2_mux4_1 _11289_ (.S0(net3777),
    .A0(\mem.mem[204][3] ),
    .A1(\mem.mem[205][3] ),
    .A2(\mem.mem[206][3] ),
    .A3(\mem.mem[207][3] ),
    .S1(net3693),
    .X(_03433_));
 sg13g2_nand2_1 _11290_ (.Y(_03434_),
    .A(net3658),
    .B(_03433_));
 sg13g2_a21oi_1 _11291_ (.A1(net3121),
    .A2(_03432_),
    .Y(_03435_),
    .B1(net3101));
 sg13g2_a22oi_1 _11292_ (.Y(_03436_),
    .B1(_03434_),
    .B2(_03435_),
    .A2(_03431_),
    .A1(_03429_));
 sg13g2_nor2b_1 _11293_ (.A(net3816),
    .B_N(\mem.mem[218][3] ),
    .Y(_03437_));
 sg13g2_a21oi_1 _11294_ (.A1(net3816),
    .A2(\mem.mem[219][3] ),
    .Y(_03438_),
    .B1(_03437_));
 sg13g2_nand2_1 _11295_ (.Y(_03439_),
    .A(net3816),
    .B(\mem.mem[217][3] ));
 sg13g2_nand2b_1 _11296_ (.Y(_03440_),
    .B(\mem.mem[216][3] ),
    .A_N(net3816));
 sg13g2_nand3_1 _11297_ (.B(_03439_),
    .C(_03440_),
    .A(net3189),
    .Y(_03441_));
 sg13g2_a21oi_1 _11298_ (.A1(net3712),
    .A2(_03438_),
    .Y(_03442_),
    .B1(net3660));
 sg13g2_mux4_1 _11299_ (.S0(net3818),
    .A0(\mem.mem[220][3] ),
    .A1(\mem.mem[221][3] ),
    .A2(\mem.mem[222][3] ),
    .A3(\mem.mem[223][3] ),
    .S1(net3713),
    .X(_03443_));
 sg13g2_a221oi_1 _11300_ (.B2(net3659),
    .C1(net3102),
    .B1(_03443_),
    .A1(_03441_),
    .Y(_03444_),
    .A2(_03442_));
 sg13g2_mux4_1 _11301_ (.S0(net3793),
    .A0(\mem.mem[212][3] ),
    .A1(\mem.mem[213][3] ),
    .A2(\mem.mem[214][3] ),
    .A3(\mem.mem[215][3] ),
    .S1(net3699),
    .X(_03445_));
 sg13g2_mux4_1 _11302_ (.S0(net3786),
    .A0(\mem.mem[208][3] ),
    .A1(\mem.mem[209][3] ),
    .A2(\mem.mem[210][3] ),
    .A3(\mem.mem[211][3] ),
    .S1(net3697),
    .X(_03446_));
 sg13g2_nand2_1 _11303_ (.Y(_03447_),
    .A(net3125),
    .B(_03446_));
 sg13g2_a21oi_1 _11304_ (.A1(net3660),
    .A2(_03445_),
    .Y(_03448_),
    .B1(net3633));
 sg13g2_a21oi_1 _11305_ (.A1(_03447_),
    .A2(_03448_),
    .Y(_03449_),
    .B1(_03444_));
 sg13g2_nand2b_1 _11306_ (.Y(_03450_),
    .B(\mem.mem[230][3] ),
    .A_N(net3869));
 sg13g2_a21oi_1 _11307_ (.A1(net3869),
    .A2(\mem.mem[231][3] ),
    .Y(_03451_),
    .B1(net3200));
 sg13g2_nor2b_1 _11308_ (.A(net3867),
    .B_N(\mem.mem[228][3] ),
    .Y(_03452_));
 sg13g2_a21oi_1 _11309_ (.A1(net3867),
    .A2(\mem.mem[229][3] ),
    .Y(_03453_),
    .B1(_03452_));
 sg13g2_a221oi_1 _11310_ (.B2(net3200),
    .C1(net3147),
    .B1(_03453_),
    .A1(_03450_),
    .Y(_03454_),
    .A2(_03451_));
 sg13g2_mux4_1 _11311_ (.S0(net3867),
    .A0(\mem.mem[224][3] ),
    .A1(\mem.mem[225][3] ),
    .A2(\mem.mem[226][3] ),
    .A3(\mem.mem[227][3] ),
    .S1(net3732),
    .X(_03455_));
 sg13g2_a21oi_2 _11312_ (.B1(_03454_),
    .Y(_03456_),
    .A2(_03455_),
    .A1(net3147));
 sg13g2_nor2b_1 _11313_ (.A(net3864),
    .B_N(\mem.mem[232][3] ),
    .Y(_03457_));
 sg13g2_a21oi_1 _11314_ (.A1(net3864),
    .A2(\mem.mem[233][3] ),
    .Y(_03458_),
    .B1(_03457_));
 sg13g2_nand2b_1 _11315_ (.Y(_03459_),
    .B(\mem.mem[234][3] ),
    .A_N(net3864));
 sg13g2_a21oi_1 _11316_ (.A1(net3864),
    .A2(\mem.mem[235][3] ),
    .Y(_03460_),
    .B1(net3201));
 sg13g2_a221oi_1 _11317_ (.B2(_03460_),
    .C1(net3674),
    .B1(_03459_),
    .A1(net3201),
    .Y(_03461_),
    .A2(_03458_));
 sg13g2_nand2b_1 _11318_ (.Y(_03462_),
    .B(\mem.mem[236][3] ),
    .A_N(net3831));
 sg13g2_a21oi_1 _11319_ (.A1(net3831),
    .A2(\mem.mem[237][3] ),
    .Y(_03463_),
    .B1(net3716));
 sg13g2_mux2_1 _11320_ (.A0(\mem.mem[238][3] ),
    .A1(\mem.mem[239][3] ),
    .S(net3830),
    .X(_03464_));
 sg13g2_a21oi_1 _11321_ (.A1(_03462_),
    .A2(_03463_),
    .Y(_03465_),
    .B1(net3136));
 sg13g2_o21ai_1 _11322_ (.B1(_03465_),
    .Y(_03466_),
    .A1(net3190),
    .A2(_03464_));
 sg13g2_nor2_1 _11323_ (.A(net3107),
    .B(_03461_),
    .Y(_03467_));
 sg13g2_a22oi_1 _11324_ (.Y(_03468_),
    .B1(_03466_),
    .B2(_03467_),
    .A2(_03456_),
    .A1(net3107));
 sg13g2_mux4_1 _11325_ (.S0(net3819),
    .A0(\mem.mem[248][3] ),
    .A1(\mem.mem[249][3] ),
    .A2(\mem.mem[250][3] ),
    .A3(\mem.mem[251][3] ),
    .S1(net3713),
    .X(_03469_));
 sg13g2_mux4_1 _11326_ (.S0(net3818),
    .A0(\mem.mem[244][3] ),
    .A1(\mem.mem[245][3] ),
    .A2(\mem.mem[246][3] ),
    .A3(\mem.mem[247][3] ),
    .S1(net3712),
    .X(_03470_));
 sg13g2_mux4_1 _11327_ (.S0(net3817),
    .A0(\mem.mem[240][3] ),
    .A1(\mem.mem[241][3] ),
    .A2(\mem.mem[242][3] ),
    .A3(\mem.mem[243][3] ),
    .S1(net3712),
    .X(_03471_));
 sg13g2_mux4_1 _11328_ (.S0(net3133),
    .A0(\mem.mem[252][3] ),
    .A1(_03469_),
    .A2(_03470_),
    .A3(_03471_),
    .S1(net3106),
    .X(_03472_));
 sg13g2_mux4_1 _11329_ (.S0(net3623),
    .A0(_03436_),
    .A1(_03449_),
    .A2(_03468_),
    .A3(_03472_),
    .S1(net3615),
    .X(_03473_));
 sg13g2_nand2_1 _11330_ (.Y(_03474_),
    .A(net3613),
    .B(_03473_));
 sg13g2_nand2b_1 _11331_ (.Y(_03475_),
    .B(\mem.mem[166][3] ),
    .A_N(net3875));
 sg13g2_a21oi_1 _11332_ (.A1(net3876),
    .A2(\mem.mem[167][3] ),
    .Y(_03476_),
    .B1(net3202));
 sg13g2_nor2b_1 _11333_ (.A(net3897),
    .B_N(\mem.mem[164][3] ),
    .Y(_03477_));
 sg13g2_a21oi_1 _11334_ (.A1(net3898),
    .A2(\mem.mem[165][3] ),
    .Y(_03478_),
    .B1(_03477_));
 sg13g2_a221oi_1 _11335_ (.B2(net3203),
    .C1(net3149),
    .B1(_03478_),
    .A1(_03475_),
    .Y(_03479_),
    .A2(_03476_));
 sg13g2_nor2b_1 _11336_ (.A(net3877),
    .B_N(\mem.mem[160][3] ),
    .Y(_03480_));
 sg13g2_a21oi_1 _11337_ (.A1(net3877),
    .A2(\mem.mem[161][3] ),
    .Y(_03481_),
    .B1(_03480_));
 sg13g2_nand2b_1 _11338_ (.Y(_03482_),
    .B(\mem.mem[162][3] ),
    .A_N(net3875));
 sg13g2_a21oi_1 _11339_ (.A1(net3877),
    .A2(\mem.mem[163][3] ),
    .Y(_03483_),
    .B1(net3202));
 sg13g2_a221oi_1 _11340_ (.B2(_03483_),
    .C1(net3675),
    .B1(_03482_),
    .A1(net3202),
    .Y(_03484_),
    .A2(_03481_));
 sg13g2_nor2_2 _11341_ (.A(_03479_),
    .B(_03484_),
    .Y(_03485_));
 sg13g2_nor2b_1 _11342_ (.A(net3899),
    .B_N(\mem.mem[168][3] ),
    .Y(_03486_));
 sg13g2_a21oi_1 _11343_ (.A1(net3894),
    .A2(\mem.mem[169][3] ),
    .Y(_03487_),
    .B1(_03486_));
 sg13g2_nand2b_1 _11344_ (.Y(_03488_),
    .B(\mem.mem[170][3] ),
    .A_N(net3894));
 sg13g2_a21oi_1 _11345_ (.A1(net3896),
    .A2(\mem.mem[171][3] ),
    .Y(_03489_),
    .B1(net3209));
 sg13g2_a221oi_1 _11346_ (.B2(_03489_),
    .C1(net3677),
    .B1(_03488_),
    .A1(net3209),
    .Y(_03490_),
    .A2(_03487_));
 sg13g2_nand2b_1 _11347_ (.Y(_03491_),
    .B(\mem.mem[172][3] ),
    .A_N(net3835));
 sg13g2_a21oi_1 _11348_ (.A1(net3835),
    .A2(\mem.mem[173][3] ),
    .Y(_03492_),
    .B1(net3718));
 sg13g2_mux2_1 _11349_ (.A0(\mem.mem[174][3] ),
    .A1(\mem.mem[175][3] ),
    .S(net3894),
    .X(_03493_));
 sg13g2_a21oi_2 _11350_ (.B1(net3137),
    .Y(_03494_),
    .A2(_03492_),
    .A1(_03491_));
 sg13g2_o21ai_1 _11351_ (.B1(_03494_),
    .Y(_03495_),
    .A1(net3209),
    .A2(_03493_));
 sg13g2_nor2_1 _11352_ (.A(net3112),
    .B(_03490_),
    .Y(_03496_));
 sg13g2_a22oi_1 _11353_ (.Y(_03497_),
    .B1(_03495_),
    .B2(_03496_),
    .A2(_03485_),
    .A1(net3112));
 sg13g2_nor2b_1 _11354_ (.A(net3860),
    .B_N(\mem.mem[180][3] ),
    .Y(_03498_));
 sg13g2_a21oi_1 _11355_ (.A1(net3900),
    .A2(\mem.mem[181][3] ),
    .Y(_03499_),
    .B1(_03498_));
 sg13g2_nand2b_1 _11356_ (.Y(_03500_),
    .B(\mem.mem[182][3] ),
    .A_N(net3900));
 sg13g2_a21oi_1 _11357_ (.A1(net3900),
    .A2(\mem.mem[183][3] ),
    .Y(_03501_),
    .B1(net3210));
 sg13g2_a221oi_1 _11358_ (.B2(_03501_),
    .C1(net3142),
    .B1(_03500_),
    .A1(net3210),
    .Y(_03502_),
    .A2(_03499_));
 sg13g2_mux4_1 _11359_ (.S0(net3852),
    .A0(\mem.mem[176][3] ),
    .A1(\mem.mem[177][3] ),
    .A2(\mem.mem[178][3] ),
    .A3(\mem.mem[179][3] ),
    .S1(net3726),
    .X(_03503_));
 sg13g2_nand2_1 _11360_ (.Y(_03504_),
    .A(net3144),
    .B(_03503_));
 sg13g2_nor2_1 _11361_ (.A(net3646),
    .B(_03502_),
    .Y(_03505_));
 sg13g2_mux4_1 _11362_ (.S0(net3857),
    .A0(\mem.mem[184][3] ),
    .A1(\mem.mem[185][3] ),
    .A2(\mem.mem[186][3] ),
    .A3(\mem.mem[187][3] ),
    .S1(net3727),
    .X(_03506_));
 sg13g2_a21oi_1 _11363_ (.A1(net3855),
    .A2(\mem.mem[191][3] ),
    .Y(_03507_),
    .B1(net3193));
 sg13g2_o21ai_1 _11364_ (.B1(_03507_),
    .Y(_03508_),
    .A1(net3855),
    .A2(_02157_));
 sg13g2_nand2b_1 _11365_ (.Y(_03509_),
    .B(\mem.mem[188][3] ),
    .A_N(net3854));
 sg13g2_a21oi_1 _11366_ (.A1(net3854),
    .A2(\mem.mem[189][3] ),
    .Y(_03510_),
    .B1(net3727));
 sg13g2_a21oi_1 _11367_ (.A1(_03509_),
    .A2(_03510_),
    .Y(_03511_),
    .B1(net3141));
 sg13g2_a221oi_1 _11368_ (.B2(_03511_),
    .C1(net3110),
    .B1(_03508_),
    .A1(net3141),
    .Y(_03512_),
    .A2(_03506_));
 sg13g2_a21oi_2 _11369_ (.B1(_03512_),
    .Y(_03513_),
    .A2(_03505_),
    .A1(_03504_));
 sg13g2_nor2b_1 _11370_ (.A(net3911),
    .B_N(\mem.mem[132][3] ),
    .Y(_03514_));
 sg13g2_a21oi_1 _11371_ (.A1(net3911),
    .A2(\mem.mem[133][3] ),
    .Y(_03515_),
    .B1(_03514_));
 sg13g2_nand2b_1 _11372_ (.Y(_03516_),
    .B(\mem.mem[134][3] ),
    .A_N(net3911));
 sg13g2_a21oi_1 _11373_ (.A1(net3911),
    .A2(\mem.mem[135][3] ),
    .Y(_03517_),
    .B1(net3214));
 sg13g2_a221oi_1 _11374_ (.B2(_03517_),
    .C1(net3157),
    .B1(_03516_),
    .A1(net3214),
    .Y(_03518_),
    .A2(_03515_));
 sg13g2_mux4_1 _11375_ (.S0(net3898),
    .A0(\mem.mem[128][3] ),
    .A1(\mem.mem[129][3] ),
    .A2(\mem.mem[130][3] ),
    .A3(\mem.mem[131][3] ),
    .S1(net3745),
    .X(_03519_));
 sg13g2_nand2_1 _11376_ (.Y(_03520_),
    .A(net3154),
    .B(_03519_));
 sg13g2_nor2_1 _11377_ (.A(net3647),
    .B(_03518_),
    .Y(_03521_));
 sg13g2_nor2b_1 _11378_ (.A(net3895),
    .B_N(\mem.mem[136][3] ),
    .Y(_03522_));
 sg13g2_a21oi_1 _11379_ (.A1(net3895),
    .A2(\mem.mem[137][3] ),
    .Y(_03523_),
    .B1(_03522_));
 sg13g2_nand2b_1 _11380_ (.Y(_03524_),
    .B(\mem.mem[138][3] ),
    .A_N(net3894));
 sg13g2_a21oi_1 _11381_ (.A1(net3895),
    .A2(\mem.mem[139][3] ),
    .Y(_03525_),
    .B1(net3212));
 sg13g2_a221oi_1 _11382_ (.B2(_03525_),
    .C1(net3677),
    .B1(_03524_),
    .A1(net3212),
    .Y(_03526_),
    .A2(_03523_));
 sg13g2_mux2_1 _11383_ (.A0(\mem.mem[142][3] ),
    .A1(\mem.mem[143][3] ),
    .S(net3910),
    .X(_03527_));
 sg13g2_nand2b_1 _11384_ (.Y(_03528_),
    .B(\mem.mem[140][3] ),
    .A_N(net3907));
 sg13g2_a21oi_1 _11385_ (.A1(net3907),
    .A2(\mem.mem[141][3] ),
    .Y(_03529_),
    .B1(net3746));
 sg13g2_a21oi_1 _11386_ (.A1(_03528_),
    .A2(_03529_),
    .Y(_03530_),
    .B1(net3156));
 sg13g2_o21ai_1 _11387_ (.B1(_03530_),
    .Y(_03531_),
    .A1(net3213),
    .A2(_03527_));
 sg13g2_nor2_1 _11388_ (.A(net3112),
    .B(_03526_),
    .Y(_03532_));
 sg13g2_a22oi_1 _11389_ (.Y(_03533_),
    .B1(_03531_),
    .B2(_03532_),
    .A2(_03521_),
    .A1(_03520_));
 sg13g2_nand2b_1 _11390_ (.Y(_03534_),
    .B(\mem.mem[150][3] ),
    .A_N(net3971));
 sg13g2_a21oi_1 _11391_ (.A1(net3972),
    .A2(\mem.mem[151][3] ),
    .Y(_03535_),
    .B1(net3234));
 sg13g2_nor2b_1 _11392_ (.A(net3981),
    .B_N(\mem.mem[148][3] ),
    .Y(_03536_));
 sg13g2_a21oi_1 _11393_ (.A1(net3971),
    .A2(\mem.mem[149][3] ),
    .Y(_03537_),
    .B1(_03536_));
 sg13g2_a221oi_1 _11394_ (.B2(net3234),
    .C1(net3167),
    .B1(_03537_),
    .A1(_03534_),
    .Y(_03538_),
    .A2(_03535_));
 sg13g2_nor2b_1 _11395_ (.A(net3965),
    .B_N(\mem.mem[144][3] ),
    .Y(_03539_));
 sg13g2_a21oi_1 _11396_ (.A1(net3965),
    .A2(\mem.mem[145][3] ),
    .Y(_03540_),
    .B1(_03539_));
 sg13g2_nand2b_1 _11397_ (.Y(_03541_),
    .B(\mem.mem[146][3] ),
    .A_N(net3965));
 sg13g2_a21oi_1 _11398_ (.A1(net3965),
    .A2(\mem.mem[147][3] ),
    .Y(_03542_),
    .B1(net3230));
 sg13g2_a221oi_1 _11399_ (.B2(_03542_),
    .C1(net3687),
    .B1(_03541_),
    .A1(net3230),
    .Y(_03543_),
    .A2(_03540_));
 sg13g2_nor2_1 _11400_ (.A(_03538_),
    .B(_03543_),
    .Y(_03544_));
 sg13g2_nor2b_1 _11401_ (.A(net3986),
    .B_N(\mem.mem[152][3] ),
    .Y(_03545_));
 sg13g2_a21oi_1 _11402_ (.A1(net3987),
    .A2(\mem.mem[153][3] ),
    .Y(_03546_),
    .B1(_03545_));
 sg13g2_nand2b_1 _11403_ (.Y(_03547_),
    .B(\mem.mem[154][3] ),
    .A_N(net3986));
 sg13g2_a21oi_1 _11404_ (.A1(net3987),
    .A2(\mem.mem[155][3] ),
    .Y(_03548_),
    .B1(net3235));
 sg13g2_a221oi_1 _11405_ (.B2(_03548_),
    .C1(net3688),
    .B1(_03547_),
    .A1(net3235),
    .Y(_03549_),
    .A2(_03546_));
 sg13g2_nand2b_1 _11406_ (.Y(_03550_),
    .B(\mem.mem[156][3] ),
    .A_N(net3966));
 sg13g2_a21oi_1 _11407_ (.A1(net3965),
    .A2(\mem.mem[157][3] ),
    .Y(_03551_),
    .B1(net3762));
 sg13g2_mux2_1 _11408_ (.A0(\mem.mem[158][3] ),
    .A1(\mem.mem[159][3] ),
    .S(net3966),
    .X(_03552_));
 sg13g2_a21oi_1 _11409_ (.A1(_03550_),
    .A2(_03551_),
    .Y(_03553_),
    .B1(net3168));
 sg13g2_o21ai_1 _11410_ (.B1(_03553_),
    .Y(_03554_),
    .A1(net3230),
    .A2(_03552_));
 sg13g2_nor2_1 _11411_ (.A(net3119),
    .B(_03549_),
    .Y(_03555_));
 sg13g2_a22oi_1 _11412_ (.Y(_03556_),
    .B1(_03554_),
    .B2(_03555_),
    .A2(_03544_),
    .A1(net3119));
 sg13g2_mux4_1 _11413_ (.S0(net3625),
    .A0(_03497_),
    .A1(_03513_),
    .A2(_03533_),
    .A3(_03556_),
    .S1(net3093),
    .X(_03557_));
 sg13g2_a21oi_1 _11414_ (.A1(net3089),
    .A2(_03557_),
    .Y(_03558_),
    .B1(_02149_));
 sg13g2_mux4_1 _11415_ (.S0(net3945),
    .A0(\mem.mem[44][3] ),
    .A1(\mem.mem[45][3] ),
    .A2(\mem.mem[46][3] ),
    .A3(\mem.mem[47][3] ),
    .S1(net3757),
    .X(_03559_));
 sg13g2_mux4_1 _11416_ (.S0(net3950),
    .A0(\mem.mem[40][3] ),
    .A1(\mem.mem[41][3] ),
    .A2(\mem.mem[42][3] ),
    .A3(\mem.mem[43][3] ),
    .S1(net3758),
    .X(_03560_));
 sg13g2_mux2_1 _11417_ (.A0(_03559_),
    .A1(_03560_),
    .S(net3163),
    .X(_03561_));
 sg13g2_nand2_1 _11418_ (.Y(_03562_),
    .A(net3648),
    .B(_03561_));
 sg13g2_mux4_1 _11419_ (.S0(net3934),
    .A0(\mem.mem[32][3] ),
    .A1(\mem.mem[33][3] ),
    .A2(\mem.mem[34][3] ),
    .A3(\mem.mem[35][3] ),
    .S1(net3753),
    .X(_03563_));
 sg13g2_mux4_1 _11420_ (.S0(net3947),
    .A0(\mem.mem[36][3] ),
    .A1(\mem.mem[37][3] ),
    .A2(\mem.mem[38][3] ),
    .A3(\mem.mem[39][3] ),
    .S1(net3757),
    .X(_03564_));
 sg13g2_mux2_1 _11421_ (.A0(_03563_),
    .A1(_03564_),
    .S(net3684),
    .X(_03565_));
 sg13g2_a21oi_1 _11422_ (.A1(net3116),
    .A2(_03565_),
    .Y(_03566_),
    .B1(net3627));
 sg13g2_mux2_1 _11423_ (.A0(\mem.mem[58][3] ),
    .A1(\mem.mem[59][3] ),
    .S(net3979),
    .X(_03567_));
 sg13g2_mux2_1 _11424_ (.A0(\mem.mem[56][3] ),
    .A1(\mem.mem[57][3] ),
    .S(net3978),
    .X(_03568_));
 sg13g2_nor2_1 _11425_ (.A(net3766),
    .B(_03568_),
    .Y(_03569_));
 sg13g2_o21ai_1 _11426_ (.B1(net3171),
    .Y(_03570_),
    .A1(net3233),
    .A2(_03567_));
 sg13g2_mux4_1 _11427_ (.S0(net3984),
    .A0(\mem.mem[60][3] ),
    .A1(\mem.mem[61][3] ),
    .A2(\mem.mem[62][3] ),
    .A3(\mem.mem[63][3] ),
    .S1(net3767),
    .X(_03571_));
 sg13g2_a21oi_1 _11428_ (.A1(net3688),
    .A2(_03571_),
    .Y(_03572_),
    .B1(net3118));
 sg13g2_o21ai_1 _11429_ (.B1(_03572_),
    .Y(_03573_),
    .A1(_03569_),
    .A2(_03570_));
 sg13g2_nand2b_1 _11430_ (.Y(_03574_),
    .B(net3976),
    .A_N(\mem.mem[53][3] ));
 sg13g2_o21ai_1 _11431_ (.B1(_03574_),
    .Y(_03575_),
    .A1(net3974),
    .A2(\mem.mem[52][3] ));
 sg13g2_nand2b_1 _11432_ (.Y(_03576_),
    .B(\mem.mem[54][3] ),
    .A_N(net3974));
 sg13g2_a21oi_1 _11433_ (.A1(net3974),
    .A2(\mem.mem[55][3] ),
    .Y(_03577_),
    .B1(net3232));
 sg13g2_a221oi_1 _11434_ (.B2(_03577_),
    .C1(net3170),
    .B1(_03576_),
    .A1(net3232),
    .Y(_03578_),
    .A2(_03575_));
 sg13g2_mux2_1 _11435_ (.A0(\mem.mem[50][3] ),
    .A1(\mem.mem[51][3] ),
    .S(net3956),
    .X(_03579_));
 sg13g2_mux2_1 _11436_ (.A0(\mem.mem[48][3] ),
    .A1(\mem.mem[49][3] ),
    .S(net3960),
    .X(_03580_));
 sg13g2_nor2_1 _11437_ (.A(net3761),
    .B(_03580_),
    .Y(_03581_));
 sg13g2_o21ai_1 _11438_ (.B1(net3169),
    .Y(_03582_),
    .A1(net3229),
    .A2(_03579_));
 sg13g2_o21ai_1 _11439_ (.B1(net3119),
    .Y(_03583_),
    .A1(_03581_),
    .A2(_03582_));
 sg13g2_o21ai_1 _11440_ (.B1(_03573_),
    .Y(_03584_),
    .A1(_03578_),
    .A2(_03583_));
 sg13g2_a221oi_1 _11441_ (.B2(net3626),
    .C1(net3092),
    .B1(_03584_),
    .A1(_03562_),
    .Y(_03585_),
    .A2(_03566_));
 sg13g2_mux4_1 _11442_ (.S0(net3926),
    .A0(\mem.mem[12][3] ),
    .A1(\mem.mem[13][3] ),
    .A2(\mem.mem[14][3] ),
    .A3(\mem.mem[15][3] ),
    .S1(net3752),
    .X(_03586_));
 sg13g2_mux4_1 _11443_ (.S0(net3880),
    .A0(\mem.mem[8][3] ),
    .A1(\mem.mem[9][3] ),
    .A2(\mem.mem[10][3] ),
    .A3(\mem.mem[11][3] ),
    .S1(net3738),
    .X(_03587_));
 sg13g2_mux2_1 _11444_ (.A0(_03586_),
    .A1(_03587_),
    .S(net3160),
    .X(_03588_));
 sg13g2_nand2_1 _11445_ (.Y(_03589_),
    .A(net3650),
    .B(_03588_));
 sg13g2_mux4_1 _11446_ (.S0(net3879),
    .A0(\mem.mem[4][3] ),
    .A1(\mem.mem[5][3] ),
    .A2(\mem.mem[6][3] ),
    .A3(\mem.mem[7][3] ),
    .S1(net3738),
    .X(_03590_));
 sg13g2_mux4_1 _11447_ (.S0(net3925),
    .A0(\mem.mem[0][3] ),
    .A1(\mem.mem[1][3] ),
    .A2(\mem.mem[2][3] ),
    .A3(\mem.mem[3][3] ),
    .S1(net3752),
    .X(_03591_));
 sg13g2_mux2_1 _11448_ (.A0(_03590_),
    .A1(_03591_),
    .S(net3160),
    .X(_03592_));
 sg13g2_a21oi_1 _11449_ (.A1(net3117),
    .A2(_03592_),
    .Y(_03593_),
    .B1(net3626));
 sg13g2_mux4_1 _11450_ (.S0(net3944),
    .A0(\mem.mem[24][3] ),
    .A1(\mem.mem[25][3] ),
    .A2(\mem.mem[26][3] ),
    .A3(\mem.mem[27][3] ),
    .S1(net3756),
    .X(_03594_));
 sg13g2_nand2_1 _11451_ (.Y(_03595_),
    .A(net3164),
    .B(_03594_));
 sg13g2_mux4_1 _11452_ (.S0(net3942),
    .A0(\mem.mem[28][3] ),
    .A1(\mem.mem[29][3] ),
    .A2(\mem.mem[30][3] ),
    .A3(\mem.mem[31][3] ),
    .S1(net3755),
    .X(_03596_));
 sg13g2_a21oi_1 _11453_ (.A1(net3684),
    .A2(_03596_),
    .Y(_03597_),
    .B1(net3115));
 sg13g2_nand2_1 _11454_ (.Y(_03598_),
    .A(_03595_),
    .B(_03597_));
 sg13g2_mux4_1 _11455_ (.S0(net3927),
    .A0(\mem.mem[16][3] ),
    .A1(\mem.mem[17][3] ),
    .A2(\mem.mem[18][3] ),
    .A3(\mem.mem[19][3] ),
    .S1(net3751),
    .X(_03599_));
 sg13g2_and2_1 _11456_ (.A(net3161),
    .B(_03599_),
    .X(_03600_));
 sg13g2_mux2_1 _11457_ (.A0(\mem.mem[22][3] ),
    .A1(\mem.mem[23][3] ),
    .S(net3943),
    .X(_03601_));
 sg13g2_mux2_1 _11458_ (.A0(\mem.mem[20][3] ),
    .A1(\mem.mem[21][3] ),
    .S(net3943),
    .X(_03602_));
 sg13g2_nor2_1 _11459_ (.A(net3756),
    .B(_03602_),
    .Y(_03603_));
 sg13g2_o21ai_1 _11460_ (.B1(net3683),
    .Y(_03604_),
    .A1(net3223),
    .A2(_03601_));
 sg13g2_o21ai_1 _11461_ (.B1(net3115),
    .Y(_03605_),
    .A1(_03603_),
    .A2(_03604_));
 sg13g2_o21ai_1 _11462_ (.B1(_03598_),
    .Y(_03606_),
    .A1(_03600_),
    .A2(_03605_));
 sg13g2_a221oi_1 _11463_ (.B2(net3626),
    .C1(net3618),
    .B1(_03606_),
    .A1(_03589_),
    .Y(_03607_),
    .A2(_03593_));
 sg13g2_or3_2 _11464_ (.A(net3614),
    .B(_03585_),
    .C(_03607_),
    .X(_03608_));
 sg13g2_mux4_1 _11465_ (.S0(net3824),
    .A0(\mem.mem[112][3] ),
    .A1(\mem.mem[113][3] ),
    .A2(\mem.mem[114][3] ),
    .A3(\mem.mem[115][3] ),
    .S1(net3714),
    .X(_03609_));
 sg13g2_mux4_1 _11466_ (.S0(net3820),
    .A0(\mem.mem[116][3] ),
    .A1(\mem.mem[117][3] ),
    .A2(\mem.mem[118][3] ),
    .A3(\mem.mem[119][3] ),
    .S1(net3714),
    .X(_03610_));
 sg13g2_and2_1 _11467_ (.A(net3670),
    .B(_03610_),
    .X(_03611_));
 sg13g2_a21oi_2 _11468_ (.B1(_03611_),
    .Y(_03612_),
    .A2(_03609_),
    .A1(net3134));
 sg13g2_mux4_1 _11469_ (.S0(net3850),
    .A0(\mem.mem[124][3] ),
    .A1(\mem.mem[125][3] ),
    .A2(\mem.mem[126][3] ),
    .A3(\mem.mem[127][3] ),
    .S1(net3725),
    .X(_03613_));
 sg13g2_mux4_1 _11470_ (.S0(net3841),
    .A0(\mem.mem[120][3] ),
    .A1(\mem.mem[121][3] ),
    .A2(\mem.mem[122][3] ),
    .A3(\mem.mem[123][3] ),
    .S1(net3721),
    .X(_03614_));
 sg13g2_mux2_1 _11471_ (.A0(_03613_),
    .A1(_03614_),
    .S(net3139),
    .X(_03615_));
 sg13g2_a21oi_1 _11472_ (.A1(net3640),
    .A2(_03615_),
    .Y(_03616_),
    .B1(net3096));
 sg13g2_o21ai_1 _11473_ (.B1(_03616_),
    .Y(_03617_),
    .A1(net3640),
    .A2(_03612_));
 sg13g2_mux4_1 _11474_ (.S0(net3915),
    .A0(\mem.mem[96][3] ),
    .A1(\mem.mem[97][3] ),
    .A2(\mem.mem[98][3] ),
    .A3(\mem.mem[99][3] ),
    .S1(net3748),
    .X(_03618_));
 sg13g2_nor2b_1 _11475_ (.A(net3915),
    .B_N(\mem.mem[102][3] ),
    .Y(_03619_));
 sg13g2_a21oi_1 _11476_ (.A1(net3915),
    .A2(\mem.mem[103][3] ),
    .Y(_03620_),
    .B1(_03619_));
 sg13g2_nand2_1 _11477_ (.Y(_03621_),
    .A(net3919),
    .B(\mem.mem[101][3] ));
 sg13g2_nand2b_1 _11478_ (.Y(_03622_),
    .B(\mem.mem[100][3] ),
    .A_N(net3916));
 sg13g2_nand3_1 _11479_ (.B(_03621_),
    .C(_03622_),
    .A(net3215),
    .Y(_03623_));
 sg13g2_a21oi_1 _11480_ (.A1(net3748),
    .A2(_03620_),
    .Y(_03624_),
    .B1(net3158));
 sg13g2_a221oi_1 _11481_ (.B2(_03624_),
    .C1(net3647),
    .B1(_03623_),
    .A1(net3158),
    .Y(_03625_),
    .A2(_03618_));
 sg13g2_mux4_1 _11482_ (.S0(net3904),
    .A0(\mem.mem[108][3] ),
    .A1(\mem.mem[109][3] ),
    .A2(\mem.mem[110][3] ),
    .A3(\mem.mem[111][3] ),
    .S1(net3744),
    .X(_03626_));
 sg13g2_nor2b_1 _11483_ (.A(net3922),
    .B_N(\mem.mem[106][3] ),
    .Y(_03627_));
 sg13g2_a21oi_1 _11484_ (.A1(net3917),
    .A2(\mem.mem[107][3] ),
    .Y(_03628_),
    .B1(_03627_));
 sg13g2_nand2_1 _11485_ (.Y(_03629_),
    .A(net3918),
    .B(\mem.mem[105][3] ));
 sg13g2_nand2b_1 _11486_ (.Y(_03630_),
    .B(\mem.mem[104][3] ),
    .A_N(net3918));
 sg13g2_nand3_1 _11487_ (.B(_03629_),
    .C(_03630_),
    .A(net3215),
    .Y(_03631_));
 sg13g2_a21oi_1 _11488_ (.A1(net3748),
    .A2(_03628_),
    .Y(_03632_),
    .B1(net3679));
 sg13g2_a221oi_1 _11489_ (.B2(_03632_),
    .C1(net3113),
    .B1(_03631_),
    .A1(net3679),
    .Y(_03633_),
    .A2(_03626_));
 sg13g2_o21ai_1 _11490_ (.B1(net3097),
    .Y(_03634_),
    .A1(_03625_),
    .A2(_03633_));
 sg13g2_and3_1 _11491_ (.X(_03635_),
    .A(net3616),
    .B(_03617_),
    .C(_03634_));
 sg13g2_mux4_1 _11492_ (.S0(net3803),
    .A0(\mem.mem[88][3] ),
    .A1(\mem.mem[89][3] ),
    .A2(\mem.mem[90][3] ),
    .A3(\mem.mem[91][3] ),
    .S1(net3705),
    .X(_03636_));
 sg13g2_nand2_1 _11493_ (.Y(_03637_),
    .A(net3129),
    .B(_03636_));
 sg13g2_mux4_1 _11494_ (.S0(net3802),
    .A0(\mem.mem[92][3] ),
    .A1(\mem.mem[93][3] ),
    .A2(\mem.mem[94][3] ),
    .A3(\mem.mem[95][3] ),
    .S1(net3706),
    .X(_03638_));
 sg13g2_a21oi_1 _11495_ (.A1(net3663),
    .A2(_03638_),
    .Y(_03639_),
    .B1(net3104));
 sg13g2_mux2_1 _11496_ (.A0(\mem.mem[82][3] ),
    .A1(\mem.mem[83][3] ),
    .S(net3798),
    .X(_03640_));
 sg13g2_mux2_1 _11497_ (.A0(\mem.mem[80][3] ),
    .A1(\mem.mem[81][3] ),
    .S(net3798),
    .X(_03641_));
 sg13g2_nor2_1 _11498_ (.A(net3703),
    .B(_03641_),
    .Y(_03642_));
 sg13g2_o21ai_1 _11499_ (.B1(net3128),
    .Y(_03643_),
    .A1(net3182),
    .A2(_03640_));
 sg13g2_mux4_1 _11500_ (.S0(net3809),
    .A0(\mem.mem[84][3] ),
    .A1(\mem.mem[85][3] ),
    .A2(\mem.mem[86][3] ),
    .A3(\mem.mem[87][3] ),
    .S1(net3708),
    .X(_03644_));
 sg13g2_a21oi_1 _11501_ (.A1(net3662),
    .A2(_03644_),
    .Y(_03645_),
    .B1(net3634));
 sg13g2_o21ai_1 _11502_ (.B1(_03645_),
    .Y(_03646_),
    .A1(_03642_),
    .A2(_03643_));
 sg13g2_mux4_1 _11503_ (.S0(net3791),
    .A0(\mem.mem[64][3] ),
    .A1(\mem.mem[65][3] ),
    .A2(\mem.mem[66][3] ),
    .A3(\mem.mem[67][3] ),
    .S1(net3698),
    .X(_03647_));
 sg13g2_mux4_1 _11504_ (.S0(net3808),
    .A0(\mem.mem[68][3] ),
    .A1(\mem.mem[69][3] ),
    .A2(\mem.mem[70][3] ),
    .A3(\mem.mem[71][3] ),
    .S1(net3708),
    .X(_03648_));
 sg13g2_nand2_1 _11505_ (.Y(_03649_),
    .A(net3661),
    .B(_03648_));
 sg13g2_a21oi_1 _11506_ (.A1(net3128),
    .A2(_03647_),
    .Y(_03650_),
    .B1(net3634));
 sg13g2_mux4_1 _11507_ (.S0(net3778),
    .A0(\mem.mem[72][3] ),
    .A1(\mem.mem[73][3] ),
    .A2(\mem.mem[74][3] ),
    .A3(\mem.mem[75][3] ),
    .S1(net3694),
    .X(_03651_));
 sg13g2_nand2_1 _11508_ (.Y(_03652_),
    .A(net3128),
    .B(_03651_));
 sg13g2_mux4_1 _11509_ (.S0(net3798),
    .A0(\mem.mem[76][3] ),
    .A1(\mem.mem[77][3] ),
    .A2(\mem.mem[78][3] ),
    .A3(\mem.mem[79][3] ),
    .S1(net3702),
    .X(_03653_));
 sg13g2_a21oi_1 _11510_ (.A1(net3661),
    .A2(_03653_),
    .Y(_03654_),
    .B1(net3103));
 sg13g2_a221oi_1 _11511_ (.B2(_03654_),
    .C1(net3624),
    .B1(_03652_),
    .A1(_03649_),
    .Y(_03655_),
    .A2(_03650_));
 sg13g2_a21oi_2 _11512_ (.B1(net3094),
    .Y(_03656_),
    .A2(_03639_),
    .A1(_03637_));
 sg13g2_a21oi_2 _11513_ (.B1(_03655_),
    .Y(_03657_),
    .A2(_03656_),
    .A1(_03646_));
 sg13g2_o21ai_1 _11514_ (.B1(net3612),
    .Y(_03658_),
    .A1(net3615),
    .A2(_03657_));
 sg13g2_o21ai_1 _11515_ (.B1(_03608_),
    .Y(_03659_),
    .A1(_03635_),
    .A2(_03658_));
 sg13g2_a22oi_1 _11516_ (.Y(_03660_),
    .B1(_03659_),
    .B2(_02149_),
    .A2(_03558_),
    .A1(_03474_));
 sg13g2_a22oi_1 _11517_ (.Y(_03661_),
    .B1(_03660_),
    .B2(_02259_),
    .A2(_02536_),
    .A1(net4));
 sg13g2_o21ai_1 _11518_ (.B1(net4006),
    .Y(_03662_),
    .A1(net5191),
    .A2(net3055));
 sg13g2_a21oi_1 _11519_ (.A1(net3055),
    .A2(_03661_),
    .Y(_00598_),
    .B1(_03662_));
 sg13g2_mux2_1 _11520_ (.A0(\mem.mem[214][4] ),
    .A1(\mem.mem[215][4] ),
    .S(net3790),
    .X(_03663_));
 sg13g2_nand2_1 _11521_ (.Y(_03664_),
    .A(net3698),
    .B(_03663_));
 sg13g2_mux2_1 _11522_ (.A0(\mem.mem[212][4] ),
    .A1(\mem.mem[213][4] ),
    .S(net3792),
    .X(_03665_));
 sg13g2_a21oi_1 _11523_ (.A1(net3179),
    .A2(_03665_),
    .Y(_03666_),
    .B1(net3127));
 sg13g2_mux2_1 _11524_ (.A0(\mem.mem[210][4] ),
    .A1(\mem.mem[211][4] ),
    .S(net3785),
    .X(_03667_));
 sg13g2_nand2_1 _11525_ (.Y(_03668_),
    .A(net3697),
    .B(_03667_));
 sg13g2_mux2_1 _11526_ (.A0(\mem.mem[208][4] ),
    .A1(\mem.mem[209][4] ),
    .S(net3785),
    .X(_03669_));
 sg13g2_a21oi_1 _11527_ (.A1(net3178),
    .A2(_03669_),
    .Y(_03670_),
    .B1(net3659));
 sg13g2_a22oi_1 _11528_ (.Y(_03671_),
    .B1(_03668_),
    .B2(_03670_),
    .A2(_03666_),
    .A1(_03664_));
 sg13g2_mux4_1 _11529_ (.S0(net3788),
    .A0(\mem.mem[216][4] ),
    .A1(\mem.mem[217][4] ),
    .A2(\mem.mem[218][4] ),
    .A3(\mem.mem[219][4] ),
    .S1(net3696),
    .X(_03672_));
 sg13g2_nand2b_1 _11530_ (.Y(_03673_),
    .B(net3125),
    .A_N(_03672_));
 sg13g2_mux2_1 _11531_ (.A0(\mem.mem[220][4] ),
    .A1(\mem.mem[221][4] ),
    .S(net3793),
    .X(_03674_));
 sg13g2_nand2_1 _11532_ (.Y(_03675_),
    .A(net3179),
    .B(_03674_));
 sg13g2_mux2_1 _11533_ (.A0(\mem.mem[222][4] ),
    .A1(\mem.mem[223][4] ),
    .S(net3787),
    .X(_03676_));
 sg13g2_a21oi_1 _11534_ (.A1(net3696),
    .A2(_03676_),
    .Y(_03677_),
    .B1(net3125));
 sg13g2_a21oi_1 _11535_ (.A1(_03675_),
    .A2(_03677_),
    .Y(_03678_),
    .B1(net3102));
 sg13g2_a221oi_1 _11536_ (.B2(_03678_),
    .C1(net3094),
    .B1(_03673_),
    .A1(net3102),
    .Y(_03679_),
    .A2(_03671_));
 sg13g2_mux2_1 _11537_ (.A0(\mem.mem[198][4] ),
    .A1(\mem.mem[199][4] ),
    .S(net3774),
    .X(_03680_));
 sg13g2_nand2_1 _11538_ (.Y(_03681_),
    .A(net3691),
    .B(_03680_));
 sg13g2_mux2_1 _11539_ (.A0(\mem.mem[196][4] ),
    .A1(\mem.mem[197][4] ),
    .S(net3771),
    .X(_03682_));
 sg13g2_a21oi_1 _11540_ (.A1(net3175),
    .A2(_03682_),
    .Y(_03683_),
    .B1(net3121));
 sg13g2_mux2_1 _11541_ (.A0(\mem.mem[194][4] ),
    .A1(\mem.mem[195][4] ),
    .S(net3771),
    .X(_03684_));
 sg13g2_nand2_1 _11542_ (.Y(_03685_),
    .A(net3691),
    .B(_03684_));
 sg13g2_mux2_1 _11543_ (.A0(\mem.mem[192][4] ),
    .A1(\mem.mem[193][4] ),
    .S(net3771),
    .X(_03686_));
 sg13g2_a21oi_1 _11544_ (.A1(net3175),
    .A2(_03686_),
    .Y(_03687_),
    .B1(net3657));
 sg13g2_a221oi_1 _11545_ (.B2(_03687_),
    .C1(net3632),
    .B1(_03685_),
    .A1(_03681_),
    .Y(_03688_),
    .A2(_03683_));
 sg13g2_mux4_1 _11546_ (.S0(net3781),
    .A0(\mem.mem[204][4] ),
    .A1(\mem.mem[205][4] ),
    .A2(\mem.mem[206][4] ),
    .A3(\mem.mem[207][4] ),
    .S1(net3694),
    .X(_03689_));
 sg13g2_inv_1 _11547_ (.Y(_03690_),
    .A(_03689_));
 sg13g2_mux4_1 _11548_ (.S0(net3777),
    .A0(\mem.mem[200][4] ),
    .A1(\mem.mem[201][4] ),
    .A2(\mem.mem[202][4] ),
    .A3(\mem.mem[203][4] ),
    .S1(net3693),
    .X(_03691_));
 sg13g2_o21ai_1 _11549_ (.B1(net3633),
    .Y(_03692_),
    .A1(net3658),
    .A2(_03691_));
 sg13g2_a21oi_1 _11550_ (.A1(net3658),
    .A2(_03690_),
    .Y(_03693_),
    .B1(_03692_));
 sg13g2_nor3_2 _11551_ (.A(net3620),
    .B(_03688_),
    .C(_03693_),
    .Y(_03694_));
 sg13g2_nor3_2 _11552_ (.A(net3615),
    .B(_03679_),
    .C(_03694_),
    .Y(_03695_));
 sg13g2_mux2_1 _11553_ (.A0(\mem.mem[236][4] ),
    .A1(\mem.mem[237][4] ),
    .S(net3866),
    .X(_03696_));
 sg13g2_nand2_1 _11554_ (.Y(_03697_),
    .A(net3201),
    .B(_03696_));
 sg13g2_mux2_1 _11555_ (.A0(\mem.mem[238][4] ),
    .A1(\mem.mem[239][4] ),
    .S(net3866),
    .X(_03698_));
 sg13g2_a21oi_1 _11556_ (.A1(net3733),
    .A2(_03698_),
    .Y(_03699_),
    .B1(net3148));
 sg13g2_mux4_1 _11557_ (.S0(net3864),
    .A0(\mem.mem[232][4] ),
    .A1(\mem.mem[233][4] ),
    .A2(\mem.mem[234][4] ),
    .A3(\mem.mem[235][4] ),
    .S1(net3733),
    .X(_03700_));
 sg13g2_o21ai_1 _11558_ (.B1(net3643),
    .Y(_03701_),
    .A1(net3674),
    .A2(_03700_));
 sg13g2_a21oi_1 _11559_ (.A1(_03697_),
    .A2(_03699_),
    .Y(_03702_),
    .B1(_03701_));
 sg13g2_mux2_1 _11560_ (.A0(\mem.mem[230][4] ),
    .A1(\mem.mem[231][4] ),
    .S(net3869),
    .X(_03703_));
 sg13g2_mux2_1 _11561_ (.A0(\mem.mem[228][4] ),
    .A1(\mem.mem[229][4] ),
    .S(net3879),
    .X(_03704_));
 sg13g2_nand2_1 _11562_ (.Y(_03705_),
    .A(net3205),
    .B(_03704_));
 sg13g2_a21oi_1 _11563_ (.A1(net3732),
    .A2(_03703_),
    .Y(_03706_),
    .B1(net3147));
 sg13g2_mux2_1 _11564_ (.A0(\mem.mem[226][4] ),
    .A1(\mem.mem[227][4] ),
    .S(net3867),
    .X(_03707_));
 sg13g2_nand2_1 _11565_ (.Y(_03708_),
    .A(net3732),
    .B(_03707_));
 sg13g2_mux2_1 _11566_ (.A0(\mem.mem[224][4] ),
    .A1(\mem.mem[225][4] ),
    .S(net3867),
    .X(_03709_));
 sg13g2_a21oi_1 _11567_ (.A1(net3200),
    .A2(_03709_),
    .Y(_03710_),
    .B1(net3674));
 sg13g2_a221oi_1 _11568_ (.B2(_03710_),
    .C1(net3644),
    .B1(_03708_),
    .A1(_03705_),
    .Y(_03711_),
    .A2(_03706_));
 sg13g2_nor3_2 _11569_ (.A(net3625),
    .B(_03702_),
    .C(_03711_),
    .Y(_03712_));
 sg13g2_mux4_1 _11570_ (.S0(net3819),
    .A0(\mem.mem[244][4] ),
    .A1(\mem.mem[245][4] ),
    .A2(\mem.mem[246][4] ),
    .A3(\mem.mem[247][4] ),
    .S1(net3713),
    .X(_03713_));
 sg13g2_mux4_1 _11571_ (.S0(net3819),
    .A0(\mem.mem[248][4] ),
    .A1(\mem.mem[249][4] ),
    .A2(\mem.mem[250][4] ),
    .A3(\mem.mem[251][4] ),
    .S1(net3713),
    .X(_03714_));
 sg13g2_mux4_1 _11572_ (.S0(net3840),
    .A0(\mem.mem[240][4] ),
    .A1(\mem.mem[241][4] ),
    .A2(\mem.mem[242][4] ),
    .A3(\mem.mem[243][4] ),
    .S1(net3713),
    .X(_03715_));
 sg13g2_mux4_1 _11573_ (.S0(net3106),
    .A0(\mem.mem[252][4] ),
    .A1(_03713_),
    .A2(_03714_),
    .A3(_03715_),
    .S1(net3133),
    .X(_03716_));
 sg13g2_o21ai_1 _11574_ (.B1(net3617),
    .Y(_03717_),
    .A1(net3095),
    .A2(_03716_));
 sg13g2_nor2_1 _11575_ (.A(_03712_),
    .B(_03717_),
    .Y(_03718_));
 sg13g2_mux4_1 _11576_ (.S0(net3873),
    .A0(\mem.mem[160][4] ),
    .A1(\mem.mem[161][4] ),
    .A2(\mem.mem[162][4] ),
    .A3(\mem.mem[163][4] ),
    .S1(net3734),
    .X(_03719_));
 sg13g2_nand2_1 _11577_ (.Y(_03720_),
    .A(net3875),
    .B(\mem.mem[165][4] ));
 sg13g2_nand2b_1 _11578_ (.Y(_03721_),
    .B(\mem.mem[164][4] ),
    .A_N(net3875));
 sg13g2_nand3_1 _11579_ (.B(_03720_),
    .C(_03721_),
    .A(net3202),
    .Y(_03722_));
 sg13g2_nor2b_1 _11580_ (.A(net3874),
    .B_N(\mem.mem[166][4] ),
    .Y(_03723_));
 sg13g2_a21oi_1 _11581_ (.A1(net3874),
    .A2(\mem.mem[167][4] ),
    .Y(_03724_),
    .B1(_03723_));
 sg13g2_a21oi_1 _11582_ (.A1(net3734),
    .A2(_03724_),
    .Y(_03725_),
    .B1(net3149));
 sg13g2_a221oi_1 _11583_ (.B2(_03725_),
    .C1(net3645),
    .B1(_03722_),
    .A1(net3149),
    .Y(_03726_),
    .A2(_03719_));
 sg13g2_nor2b_1 _11584_ (.A(net3835),
    .B_N(\mem.mem[172][4] ),
    .Y(_03727_));
 sg13g2_a21oi_1 _11585_ (.A1(net3835),
    .A2(\mem.mem[173][4] ),
    .Y(_03728_),
    .B1(_03727_));
 sg13g2_nand2b_1 _11586_ (.Y(_03729_),
    .B(\mem.mem[174][4] ),
    .A_N(net3836));
 sg13g2_a21oi_1 _11587_ (.A1(net3852),
    .A2(\mem.mem[175][4] ),
    .Y(_03730_),
    .B1(net3196));
 sg13g2_a221oi_1 _11588_ (.B2(_03730_),
    .C1(net3137),
    .B1(_03729_),
    .A1(net3196),
    .Y(_03731_),
    .A2(_03728_));
 sg13g2_mux2_1 _11589_ (.A0(\mem.mem[168][4] ),
    .A1(\mem.mem[169][4] ),
    .S(net3852),
    .X(_03732_));
 sg13g2_nor2_1 _11590_ (.A(net3726),
    .B(_03732_),
    .Y(_03733_));
 sg13g2_mux2_1 _11591_ (.A0(\mem.mem[170][4] ),
    .A1(\mem.mem[171][4] ),
    .S(net3851),
    .X(_03734_));
 sg13g2_o21ai_1 _11592_ (.B1(net3144),
    .Y(_03735_),
    .A1(net3209),
    .A2(_03734_));
 sg13g2_o21ai_1 _11593_ (.B1(net3646),
    .Y(_03736_),
    .A1(_03733_),
    .A2(_03735_));
 sg13g2_o21ai_1 _11594_ (.B1(net3097),
    .Y(_03737_),
    .A1(_03731_),
    .A2(_03736_));
 sg13g2_nor2_1 _11595_ (.A(_03726_),
    .B(_03737_),
    .Y(_03738_));
 sg13g2_mux4_1 _11596_ (.S0(net3858),
    .A0(\mem.mem[176][4] ),
    .A1(\mem.mem[177][4] ),
    .A2(\mem.mem[178][4] ),
    .A3(\mem.mem[179][4] ),
    .S1(net3728),
    .X(_03739_));
 sg13g2_nand2_1 _11597_ (.Y(_03740_),
    .A(net3900),
    .B(\mem.mem[181][4] ));
 sg13g2_nand2b_1 _11598_ (.Y(_03741_),
    .B(\mem.mem[180][4] ),
    .A_N(net3858));
 sg13g2_nand3_1 _11599_ (.B(_03740_),
    .C(_03741_),
    .A(net3210),
    .Y(_03742_));
 sg13g2_nor2b_1 _11600_ (.A(net3858),
    .B_N(\mem.mem[182][4] ),
    .Y(_03743_));
 sg13g2_a21oi_1 _11601_ (.A1(net3858),
    .A2(\mem.mem[183][4] ),
    .Y(_03744_),
    .B1(_03743_));
 sg13g2_a21oi_1 _11602_ (.A1(net3728),
    .A2(_03744_),
    .Y(_03745_),
    .B1(net3142));
 sg13g2_a221oi_1 _11603_ (.B2(_03745_),
    .C1(net3646),
    .B1(_03742_),
    .A1(net3142),
    .Y(_03746_),
    .A2(_03739_));
 sg13g2_mux2_1 _11604_ (.A0(\mem.mem[184][4] ),
    .A1(\mem.mem[185][4] ),
    .S(net3857),
    .X(_03747_));
 sg13g2_nor2_1 _11605_ (.A(net3727),
    .B(_03747_),
    .Y(_03748_));
 sg13g2_mux2_1 _11606_ (.A0(\mem.mem[186][4] ),
    .A1(\mem.mem[187][4] ),
    .S(net3860),
    .X(_03749_));
 sg13g2_o21ai_1 _11607_ (.B1(net3141),
    .Y(_03750_),
    .A1(net3194),
    .A2(_03749_));
 sg13g2_nor2b_1 _11608_ (.A(net3856),
    .B_N(\mem.mem[188][4] ),
    .Y(_03751_));
 sg13g2_a21oi_1 _11609_ (.A1(net3856),
    .A2(\mem.mem[189][4] ),
    .Y(_03752_),
    .B1(_03751_));
 sg13g2_nand2b_1 _11610_ (.Y(_03753_),
    .B(\mem.mem[190][4] ),
    .A_N(net3857));
 sg13g2_a21oi_1 _11611_ (.A1(net3855),
    .A2(\mem.mem[191][4] ),
    .Y(_03754_),
    .B1(net3194));
 sg13g2_a221oi_1 _11612_ (.B2(_03754_),
    .C1(net3141),
    .B1(_03753_),
    .A1(net3194),
    .Y(_03755_),
    .A2(_03752_));
 sg13g2_o21ai_1 _11613_ (.B1(net3641),
    .Y(_03756_),
    .A1(_03748_),
    .A2(_03750_));
 sg13g2_o21ai_1 _11614_ (.B1(net3622),
    .Y(_03757_),
    .A1(_03755_),
    .A2(_03756_));
 sg13g2_nor2_2 _11615_ (.A(_03746_),
    .B(_03757_),
    .Y(_03758_));
 sg13g2_o21ai_1 _11616_ (.B1(net3616),
    .Y(_03759_),
    .A1(_03738_),
    .A2(_03758_));
 sg13g2_mux4_1 _11617_ (.S0(net3910),
    .A0(\mem.mem[128][4] ),
    .A1(\mem.mem[129][4] ),
    .A2(\mem.mem[130][4] ),
    .A3(\mem.mem[131][4] ),
    .S1(net3746),
    .X(_03760_));
 sg13g2_nand2_1 _11618_ (.Y(_03761_),
    .A(net3155),
    .B(_03760_));
 sg13g2_nand2_1 _11619_ (.Y(_03762_),
    .A(net3955),
    .B(\mem.mem[133][4] ));
 sg13g2_nand2b_1 _11620_ (.Y(_03763_),
    .B(\mem.mem[132][4] ),
    .A_N(net3955));
 sg13g2_nand3_1 _11621_ (.B(_03762_),
    .C(_03763_),
    .A(net3228),
    .Y(_03764_));
 sg13g2_nor2b_1 _11622_ (.A(net3955),
    .B_N(\mem.mem[134][4] ),
    .Y(_03765_));
 sg13g2_a21oi_1 _11623_ (.A1(net3955),
    .A2(\mem.mem[135][4] ),
    .Y(_03766_),
    .B1(_03765_));
 sg13g2_a21oi_1 _11624_ (.A1(net3760),
    .A2(_03766_),
    .Y(_03767_),
    .B1(net3166));
 sg13g2_a21oi_1 _11625_ (.A1(_03764_),
    .A2(_03767_),
    .Y(_03768_),
    .B1(net3652));
 sg13g2_mux4_1 _11626_ (.S0(net3897),
    .A0(\mem.mem[136][4] ),
    .A1(\mem.mem[137][4] ),
    .A2(\mem.mem[138][4] ),
    .A3(\mem.mem[139][4] ),
    .S1(net3742),
    .X(_03769_));
 sg13g2_nand2_1 _11627_ (.Y(_03770_),
    .A(net3155),
    .B(_03769_));
 sg13g2_nand2b_1 _11628_ (.Y(_03771_),
    .B(\mem.mem[142][4] ),
    .A_N(net3912));
 sg13g2_a21oi_1 _11629_ (.A1(net3911),
    .A2(\mem.mem[143][4] ),
    .Y(_03772_),
    .B1(net3214));
 sg13g2_nor2b_1 _11630_ (.A(net3913),
    .B_N(\mem.mem[140][4] ),
    .Y(_03773_));
 sg13g2_a21oi_1 _11631_ (.A1(net3911),
    .A2(\mem.mem[141][4] ),
    .Y(_03774_),
    .B1(_03773_));
 sg13g2_a221oi_1 _11632_ (.B2(net3214),
    .C1(net3157),
    .B1(_03774_),
    .A1(_03771_),
    .Y(_03775_),
    .A2(_03772_));
 sg13g2_nor2_1 _11633_ (.A(net3113),
    .B(_03775_),
    .Y(_03776_));
 sg13g2_a221oi_1 _11634_ (.B2(_03776_),
    .C1(net3629),
    .B1(_03770_),
    .A1(_03761_),
    .Y(_03777_),
    .A2(_03768_));
 sg13g2_mux4_1 _11635_ (.S0(net3967),
    .A0(\mem.mem[144][4] ),
    .A1(\mem.mem[145][4] ),
    .A2(\mem.mem[146][4] ),
    .A3(\mem.mem[147][4] ),
    .S1(net3762),
    .X(_03778_));
 sg13g2_nand2_1 _11636_ (.Y(_03779_),
    .A(net3981),
    .B(\mem.mem[149][4] ));
 sg13g2_nand2b_1 _11637_ (.Y(_03780_),
    .B(\mem.mem[148][4] ),
    .A_N(net3981));
 sg13g2_nand3_1 _11638_ (.B(_03779_),
    .C(_03780_),
    .A(net3234),
    .Y(_03781_));
 sg13g2_nor2b_1 _11639_ (.A(net3972),
    .B_N(\mem.mem[150][4] ),
    .Y(_03782_));
 sg13g2_a21oi_1 _11640_ (.A1(net3972),
    .A2(\mem.mem[151][4] ),
    .Y(_03783_),
    .B1(_03782_));
 sg13g2_a21oi_1 _11641_ (.A1(net3763),
    .A2(_03783_),
    .Y(_03784_),
    .B1(net3167));
 sg13g2_a221oi_1 _11642_ (.B2(_03784_),
    .C1(net3651),
    .B1(_03781_),
    .A1(net3167),
    .Y(_03785_),
    .A2(_03778_));
 sg13g2_mux2_1 _11643_ (.A0(\mem.mem[152][4] ),
    .A1(\mem.mem[153][4] ),
    .S(net3987),
    .X(_03786_));
 sg13g2_nor2_1 _11644_ (.A(net3767),
    .B(_03786_),
    .Y(_03787_));
 sg13g2_mux2_1 _11645_ (.A0(\mem.mem[154][4] ),
    .A1(\mem.mem[155][4] ),
    .S(net3986),
    .X(_03788_));
 sg13g2_o21ai_1 _11646_ (.B1(net3172),
    .Y(_03789_),
    .A1(net3235),
    .A2(_03788_));
 sg13g2_nor2b_1 _11647_ (.A(net3969),
    .B_N(\mem.mem[156][4] ),
    .Y(_03790_));
 sg13g2_a21oi_1 _11648_ (.A1(net3969),
    .A2(\mem.mem[157][4] ),
    .Y(_03791_),
    .B1(_03790_));
 sg13g2_nand2b_1 _11649_ (.Y(_03792_),
    .B(\mem.mem[158][4] ),
    .A_N(net3970));
 sg13g2_a21oi_1 _11650_ (.A1(net3969),
    .A2(\mem.mem[159][4] ),
    .Y(_03793_),
    .B1(net3230));
 sg13g2_a221oi_1 _11651_ (.B2(_03793_),
    .C1(net3168),
    .B1(_03792_),
    .A1(net3230),
    .Y(_03794_),
    .A2(_03791_));
 sg13g2_o21ai_1 _11652_ (.B1(net3654),
    .Y(_03795_),
    .A1(_03787_),
    .A2(_03789_));
 sg13g2_o21ai_1 _11653_ (.B1(net3629),
    .Y(_03796_),
    .A1(_03794_),
    .A2(_03795_));
 sg13g2_nor2_2 _11654_ (.A(_03785_),
    .B(_03796_),
    .Y(_03797_));
 sg13g2_o21ai_1 _11655_ (.B1(net3093),
    .Y(_03798_),
    .A1(_03777_),
    .A2(_03797_));
 sg13g2_o21ai_1 _11656_ (.B1(net3612),
    .Y(_03799_),
    .A1(_03695_),
    .A2(_03718_));
 sg13g2_a21o_1 _11657_ (.A2(_03798_),
    .A1(_03759_),
    .B1(net3613),
    .X(_03800_));
 sg13g2_nand3_1 _11658_ (.B(_03799_),
    .C(_03800_),
    .A(net3611),
    .Y(_03801_));
 sg13g2_mux2_1 _11659_ (.A0(\mem.mem[6][4] ),
    .A1(\mem.mem[7][4] ),
    .S(net3884),
    .X(_03802_));
 sg13g2_nand2_1 _11660_ (.Y(_03803_),
    .A(net3737),
    .B(_03802_));
 sg13g2_mux2_1 _11661_ (.A0(\mem.mem[4][4] ),
    .A1(\mem.mem[5][4] ),
    .S(net3884),
    .X(_03804_));
 sg13g2_a21oi_1 _11662_ (.A1(net3219),
    .A2(_03804_),
    .Y(_03805_),
    .B1(net3151));
 sg13g2_mux2_1 _11663_ (.A0(\mem.mem[2][4] ),
    .A1(\mem.mem[3][4] ),
    .S(net3925),
    .X(_03806_));
 sg13g2_nand2_1 _11664_ (.Y(_03807_),
    .A(net3737),
    .B(_03806_));
 sg13g2_mux2_1 _11665_ (.A0(\mem.mem[0][4] ),
    .A1(\mem.mem[1][4] ),
    .S(net3884),
    .X(_03808_));
 sg13g2_a21oi_1 _11666_ (.A1(net3219),
    .A2(_03808_),
    .Y(_03809_),
    .B1(net3682));
 sg13g2_a221oi_1 _11667_ (.B2(_03809_),
    .C1(net3650),
    .B1(_03807_),
    .A1(_03803_),
    .Y(_03810_),
    .A2(_03805_));
 sg13g2_mux2_1 _11668_ (.A0(\mem.mem[12][4] ),
    .A1(\mem.mem[13][4] ),
    .S(net3926),
    .X(_03811_));
 sg13g2_nand2_1 _11669_ (.Y(_03812_),
    .A(net3219),
    .B(_03811_));
 sg13g2_mux2_1 _11670_ (.A0(\mem.mem[14][4] ),
    .A1(\mem.mem[15][4] ),
    .S(net3931),
    .X(_03813_));
 sg13g2_a21oi_1 _11671_ (.A1(net3737),
    .A2(_03813_),
    .Y(_03814_),
    .B1(net3151));
 sg13g2_mux4_1 _11672_ (.S0(net3883),
    .A0(\mem.mem[8][4] ),
    .A1(\mem.mem[9][4] ),
    .A2(\mem.mem[10][4] ),
    .A3(\mem.mem[11][4] ),
    .S1(net3737),
    .X(_03815_));
 sg13g2_o21ai_1 _11673_ (.B1(net3644),
    .Y(_03816_),
    .A1(net3681),
    .A2(_03815_));
 sg13g2_a21oi_1 _11674_ (.A1(_03812_),
    .A2(_03814_),
    .Y(_03817_),
    .B1(_03816_));
 sg13g2_nor3_1 _11675_ (.A(net3628),
    .B(_03810_),
    .C(_03817_),
    .Y(_03818_));
 sg13g2_mux2_1 _11676_ (.A0(\mem.mem[22][4] ),
    .A1(\mem.mem[23][4] ),
    .S(net3939),
    .X(_03819_));
 sg13g2_nand2_1 _11677_ (.Y(_03820_),
    .A(net3755),
    .B(_03819_));
 sg13g2_mux2_1 _11678_ (.A0(\mem.mem[20][4] ),
    .A1(\mem.mem[21][4] ),
    .S(net3943),
    .X(_03821_));
 sg13g2_a21oi_1 _11679_ (.A1(net3223),
    .A2(_03821_),
    .Y(_03822_),
    .B1(net3161));
 sg13g2_mux2_1 _11680_ (.A0(\mem.mem[18][4] ),
    .A1(\mem.mem[19][4] ),
    .S(net3927),
    .X(_03823_));
 sg13g2_nand2_1 _11681_ (.Y(_03824_),
    .A(net3751),
    .B(_03823_));
 sg13g2_mux2_1 _11682_ (.A0(\mem.mem[16][4] ),
    .A1(\mem.mem[17][4] ),
    .S(net3939),
    .X(_03825_));
 sg13g2_a21oi_1 _11683_ (.A1(net3222),
    .A2(_03825_),
    .Y(_03826_),
    .B1(net3683));
 sg13g2_a221oi_1 _11684_ (.B2(_03826_),
    .C1(net3648),
    .B1(_03824_),
    .A1(_03820_),
    .Y(_03827_),
    .A2(_03822_));
 sg13g2_mux4_1 _11685_ (.S0(net3944),
    .A0(\mem.mem[24][4] ),
    .A1(\mem.mem[25][4] ),
    .A2(\mem.mem[26][4] ),
    .A3(\mem.mem[27][4] ),
    .S1(net3756),
    .X(_03828_));
 sg13g2_nor2_1 _11686_ (.A(net3684),
    .B(_03828_),
    .Y(_03829_));
 sg13g2_nor2b_1 _11687_ (.A(\mem.mem[29][4] ),
    .B_N(net3941),
    .Y(_03830_));
 sg13g2_nor2_1 _11688_ (.A(net3940),
    .B(\mem.mem[28][4] ),
    .Y(_03831_));
 sg13g2_nor3_1 _11689_ (.A(net3755),
    .B(_03830_),
    .C(_03831_),
    .Y(_03832_));
 sg13g2_nor2b_1 _11690_ (.A(\mem.mem[31][4] ),
    .B_N(net3940),
    .Y(_03833_));
 sg13g2_o21ai_1 _11691_ (.B1(net3751),
    .Y(_03834_),
    .A1(net3930),
    .A2(\mem.mem[30][4] ));
 sg13g2_o21ai_1 _11692_ (.B1(net3683),
    .Y(_03835_),
    .A1(_03833_),
    .A2(_03834_));
 sg13g2_o21ai_1 _11693_ (.B1(net3648),
    .Y(_03836_),
    .A1(_03832_),
    .A2(_03835_));
 sg13g2_o21ai_1 _11694_ (.B1(net3626),
    .Y(_03837_),
    .A1(_03829_),
    .A2(_03836_));
 sg13g2_o21ai_1 _11695_ (.B1(net3092),
    .Y(_03838_),
    .A1(_03827_),
    .A2(_03837_));
 sg13g2_nor2_2 _11696_ (.A(_03818_),
    .B(_03838_),
    .Y(_03839_));
 sg13g2_nand2b_1 _11697_ (.Y(_03840_),
    .B(\mem.mem[38][4] ),
    .A_N(net3950));
 sg13g2_a21oi_1 _11698_ (.A1(net3950),
    .A2(\mem.mem[39][4] ),
    .Y(_03841_),
    .B1(net3225));
 sg13g2_nor2b_1 _11699_ (.A(net3951),
    .B_N(\mem.mem[36][4] ),
    .Y(_03842_));
 sg13g2_a21oi_1 _11700_ (.A1(net3951),
    .A2(\mem.mem[37][4] ),
    .Y(_03843_),
    .B1(_03842_));
 sg13g2_a221oi_1 _11701_ (.B2(net3224),
    .C1(net3163),
    .B1(_03843_),
    .A1(_03840_),
    .Y(_03844_),
    .A2(_03841_));
 sg13g2_nor2b_1 _11702_ (.A(net3935),
    .B_N(\mem.mem[32][4] ),
    .Y(_03845_));
 sg13g2_a21oi_1 _11703_ (.A1(net3935),
    .A2(\mem.mem[33][4] ),
    .Y(_03846_),
    .B1(_03845_));
 sg13g2_nand2b_1 _11704_ (.Y(_03847_),
    .B(\mem.mem[34][4] ),
    .A_N(net3932));
 sg13g2_a21oi_1 _11705_ (.A1(net3932),
    .A2(\mem.mem[35][4] ),
    .Y(_03848_),
    .B1(net3221));
 sg13g2_a221oi_1 _11706_ (.B2(_03848_),
    .C1(net3685),
    .B1(_03847_),
    .A1(net3221),
    .Y(_03849_),
    .A2(_03846_));
 sg13g2_o21ai_1 _11707_ (.B1(net3116),
    .Y(_03850_),
    .A1(_03844_),
    .A2(_03849_));
 sg13g2_mux4_1 _11708_ (.S0(net3979),
    .A0(\mem.mem[40][4] ),
    .A1(\mem.mem[41][4] ),
    .A2(\mem.mem[42][4] ),
    .A3(\mem.mem[43][4] ),
    .S1(net3765),
    .X(_03851_));
 sg13g2_nand2b_1 _11709_ (.Y(_03852_),
    .B(\mem.mem[44][4] ),
    .A_N(net3975));
 sg13g2_a21oi_1 _11710_ (.A1(net3975),
    .A2(\mem.mem[45][4] ),
    .Y(_03853_),
    .B1(net3766));
 sg13g2_nor2b_1 _11711_ (.A(net3975),
    .B_N(\mem.mem[46][4] ),
    .Y(_03854_));
 sg13g2_a21oi_1 _11712_ (.A1(net3975),
    .A2(\mem.mem[47][4] ),
    .Y(_03855_),
    .B1(_03854_));
 sg13g2_a221oi_1 _11713_ (.B2(net3766),
    .C1(net3170),
    .B1(_03855_),
    .A1(_03852_),
    .Y(_03856_),
    .A2(_03853_));
 sg13g2_a21o_1 _11714_ (.A2(_03851_),
    .A1(net3170),
    .B1(_03856_),
    .X(_03857_));
 sg13g2_a21oi_1 _11715_ (.A1(net3653),
    .A2(_03857_),
    .Y(_03858_),
    .B1(net3630));
 sg13g2_nor2b_1 _11716_ (.A(net3974),
    .B_N(\mem.mem[52][4] ),
    .Y(_03859_));
 sg13g2_a21oi_1 _11717_ (.A1(net3974),
    .A2(\mem.mem[53][4] ),
    .Y(_03860_),
    .B1(_03859_));
 sg13g2_nand2b_1 _11718_ (.Y(_03861_),
    .B(\mem.mem[54][4] ),
    .A_N(net3960));
 sg13g2_a21oi_1 _11719_ (.A1(net3974),
    .A2(\mem.mem[55][4] ),
    .Y(_03862_),
    .B1(net3232));
 sg13g2_a221oi_1 _11720_ (.B2(_03862_),
    .C1(net3170),
    .B1(_03861_),
    .A1(net3232),
    .Y(_03863_),
    .A2(_03860_));
 sg13g2_nor2b_1 _11721_ (.A(net3955),
    .B_N(\mem.mem[48][4] ),
    .Y(_03864_));
 sg13g2_a21oi_1 _11722_ (.A1(net3955),
    .A2(\mem.mem[49][4] ),
    .Y(_03865_),
    .B1(_03864_));
 sg13g2_nand2b_1 _11723_ (.Y(_03866_),
    .B(\mem.mem[50][4] ),
    .A_N(net3956));
 sg13g2_a21oi_1 _11724_ (.A1(net3956),
    .A2(\mem.mem[51][4] ),
    .Y(_03867_),
    .B1(net3228));
 sg13g2_a221oi_1 _11725_ (.B2(_03867_),
    .C1(net3686),
    .B1(_03866_),
    .A1(net3229),
    .Y(_03868_),
    .A2(_03865_));
 sg13g2_o21ai_1 _11726_ (.B1(net3118),
    .Y(_03869_),
    .A1(_03863_),
    .A2(_03868_));
 sg13g2_mux4_1 _11727_ (.S0(net3980),
    .A0(\mem.mem[56][4] ),
    .A1(\mem.mem[57][4] ),
    .A2(\mem.mem[58][4] ),
    .A3(\mem.mem[59][4] ),
    .S1(net3765),
    .X(_03870_));
 sg13g2_nor2b_1 _11728_ (.A(net3985),
    .B_N(\mem.mem[62][4] ),
    .Y(_03871_));
 sg13g2_a21oi_1 _11729_ (.A1(net3985),
    .A2(\mem.mem[63][4] ),
    .Y(_03872_),
    .B1(_03871_));
 sg13g2_nand2b_1 _11730_ (.Y(_03873_),
    .B(\mem.mem[60][4] ),
    .A_N(net3985));
 sg13g2_a21oi_1 _11731_ (.A1(net3985),
    .A2(\mem.mem[61][4] ),
    .Y(_03874_),
    .B1(net3767));
 sg13g2_a221oi_1 _11732_ (.B2(_03874_),
    .C1(net3172),
    .B1(_03873_),
    .A1(net3767),
    .Y(_03875_),
    .A2(_03872_));
 sg13g2_a21o_1 _11733_ (.A2(_03870_),
    .A1(net3171),
    .B1(_03875_),
    .X(_03876_));
 sg13g2_a21oi_1 _11734_ (.A1(net3653),
    .A2(_03876_),
    .Y(_03877_),
    .B1(net3099));
 sg13g2_a221oi_1 _11735_ (.B2(_03877_),
    .C1(net3092),
    .B1(_03869_),
    .A1(_03850_),
    .Y(_03878_),
    .A2(_03858_));
 sg13g2_mux4_1 _11736_ (.S0(net3798),
    .A0(\mem.mem[80][4] ),
    .A1(\mem.mem[81][4] ),
    .A2(\mem.mem[82][4] ),
    .A3(\mem.mem[83][4] ),
    .S1(net3703),
    .X(_03879_));
 sg13g2_mux2_1 _11737_ (.A0(\mem.mem[84][4] ),
    .A1(\mem.mem[85][4] ),
    .S(net3813),
    .X(_03880_));
 sg13g2_nand2_1 _11738_ (.Y(_03881_),
    .A(net3184),
    .B(_03880_));
 sg13g2_mux2_1 _11739_ (.A0(\mem.mem[86][4] ),
    .A1(\mem.mem[87][4] ),
    .S(net3813),
    .X(_03882_));
 sg13g2_a21oi_1 _11740_ (.A1(net3709),
    .A2(_03882_),
    .Y(_03883_),
    .B1(net3132));
 sg13g2_a21oi_1 _11741_ (.A1(_03881_),
    .A2(_03883_),
    .Y(_03884_),
    .B1(net3636));
 sg13g2_o21ai_1 _11742_ (.B1(_03884_),
    .Y(_03885_),
    .A1(net3664),
    .A2(_03879_));
 sg13g2_mux4_1 _11743_ (.S0(net3802),
    .A0(\mem.mem[88][4] ),
    .A1(\mem.mem[89][4] ),
    .A2(\mem.mem[90][4] ),
    .A3(\mem.mem[91][4] ),
    .S1(net3705),
    .X(_03886_));
 sg13g2_nor2_1 _11744_ (.A(net3663),
    .B(_03886_),
    .Y(_03887_));
 sg13g2_mux2_1 _11745_ (.A0(\mem.mem[92][4] ),
    .A1(\mem.mem[93][4] ),
    .S(net3802),
    .X(_03888_));
 sg13g2_nor2b_1 _11746_ (.A(\mem.mem[95][4] ),
    .B_N(net3802),
    .Y(_03889_));
 sg13g2_o21ai_1 _11747_ (.B1(net3706),
    .Y(_03890_),
    .A1(net3802),
    .A2(\mem.mem[94][4] ));
 sg13g2_o21ai_1 _11748_ (.B1(net3663),
    .Y(_03891_),
    .A1(_03889_),
    .A2(_03890_));
 sg13g2_a21oi_1 _11749_ (.A1(net3183),
    .A2(_03888_),
    .Y(_03892_),
    .B1(_03891_));
 sg13g2_nor3_2 _11750_ (.A(net3103),
    .B(_03887_),
    .C(_03892_),
    .Y(_03893_));
 sg13g2_nor2_1 _11751_ (.A(net3094),
    .B(_03893_),
    .Y(_03894_));
 sg13g2_mux4_1 _11752_ (.S0(net3795),
    .A0(\mem.mem[64][4] ),
    .A1(\mem.mem[65][4] ),
    .A2(\mem.mem[66][4] ),
    .A3(\mem.mem[67][4] ),
    .S1(net3699),
    .X(_03895_));
 sg13g2_nor2_1 _11753_ (.A(net3665),
    .B(_03895_),
    .Y(_03896_));
 sg13g2_mux2_1 _11754_ (.A0(\mem.mem[70][4] ),
    .A1(\mem.mem[71][4] ),
    .S(net3813),
    .X(_03897_));
 sg13g2_nand2b_1 _11755_ (.Y(_03898_),
    .B(net3813),
    .A_N(\mem.mem[69][4] ));
 sg13g2_o21ai_1 _11756_ (.B1(_03898_),
    .Y(_03899_),
    .A1(net3813),
    .A2(\mem.mem[68][4] ));
 sg13g2_o21ai_1 _11757_ (.B1(net3664),
    .Y(_03900_),
    .A1(net3708),
    .A2(_03899_));
 sg13g2_a21oi_1 _11758_ (.A1(net3708),
    .A2(_03897_),
    .Y(_03901_),
    .B1(_03900_));
 sg13g2_or3_1 _11759_ (.A(net3635),
    .B(_03896_),
    .C(_03901_),
    .X(_03902_));
 sg13g2_mux4_1 _11760_ (.S0(net3798),
    .A0(\mem.mem[76][4] ),
    .A1(\mem.mem[77][4] ),
    .A2(\mem.mem[78][4] ),
    .A3(\mem.mem[79][4] ),
    .S1(net3702),
    .X(_03903_));
 sg13g2_inv_1 _11761_ (.Y(_03904_),
    .A(_03903_));
 sg13g2_mux4_1 _11762_ (.S0(net3797),
    .A0(\mem.mem[72][4] ),
    .A1(\mem.mem[73][4] ),
    .A2(\mem.mem[74][4] ),
    .A3(\mem.mem[75][4] ),
    .S1(net3702),
    .X(_03905_));
 sg13g2_o21ai_1 _11763_ (.B1(net3634),
    .Y(_03906_),
    .A1(net3661),
    .A2(_03905_));
 sg13g2_a21oi_2 _11764_ (.B1(_03906_),
    .Y(_03907_),
    .A2(_03904_),
    .A1(net3661));
 sg13g2_nor2_1 _11765_ (.A(net3621),
    .B(_03907_),
    .Y(_03908_));
 sg13g2_a221oi_1 _11766_ (.B2(_03908_),
    .C1(net3615),
    .B1(_03902_),
    .A1(_03885_),
    .Y(_03909_),
    .A2(_03894_));
 sg13g2_nand2b_1 _11767_ (.Y(_03910_),
    .B(\mem.mem[102][4] ),
    .A_N(net3909));
 sg13g2_a21oi_1 _11768_ (.A1(net3909),
    .A2(\mem.mem[103][4] ),
    .Y(_03911_),
    .B1(net3213));
 sg13g2_nor2b_1 _11769_ (.A(net3913),
    .B_N(\mem.mem[100][4] ),
    .Y(_03912_));
 sg13g2_a21oi_1 _11770_ (.A1(net3913),
    .A2(\mem.mem[101][4] ),
    .Y(_03913_),
    .B1(_03912_));
 sg13g2_a221oi_1 _11771_ (.B2(net3213),
    .C1(net3156),
    .B1(_03913_),
    .A1(_03910_),
    .Y(_03914_),
    .A2(_03911_));
 sg13g2_nor2b_1 _11772_ (.A(net3902),
    .B_N(\mem.mem[96][4] ),
    .Y(_03915_));
 sg13g2_a21oi_1 _11773_ (.A1(net3896),
    .A2(\mem.mem[97][4] ),
    .Y(_03916_),
    .B1(_03915_));
 sg13g2_nand2b_1 _11774_ (.Y(_03917_),
    .B(\mem.mem[98][4] ),
    .A_N(net3900));
 sg13g2_a21oi_1 _11775_ (.A1(net3896),
    .A2(\mem.mem[99][4] ),
    .Y(_03918_),
    .B1(net3210));
 sg13g2_a221oi_1 _11776_ (.B2(_03918_),
    .C1(net3678),
    .B1(_03917_),
    .A1(net3210),
    .Y(_03919_),
    .A2(_03916_));
 sg13g2_o21ai_1 _11777_ (.B1(net3112),
    .Y(_03920_),
    .A1(_03914_),
    .A2(_03919_));
 sg13g2_mux4_1 _11778_ (.S0(net3905),
    .A0(\mem.mem[104][4] ),
    .A1(\mem.mem[105][4] ),
    .A2(\mem.mem[106][4] ),
    .A3(\mem.mem[107][4] ),
    .S1(net3744),
    .X(_03921_));
 sg13g2_nand2b_1 _11779_ (.Y(_03922_),
    .B(\mem.mem[108][4] ),
    .A_N(net3861));
 sg13g2_a21oi_1 _11780_ (.A1(net3861),
    .A2(\mem.mem[109][4] ),
    .Y(_03923_),
    .B1(net3728));
 sg13g2_nor2b_1 _11781_ (.A(net3860),
    .B_N(\mem.mem[110][4] ),
    .Y(_03924_));
 sg13g2_a21oi_1 _11782_ (.A1(net3860),
    .A2(\mem.mem[111][4] ),
    .Y(_03925_),
    .B1(_03924_));
 sg13g2_a221oi_1 _11783_ (.B2(net3728),
    .C1(net3142),
    .B1(_03925_),
    .A1(_03922_),
    .Y(_03926_),
    .A2(_03923_));
 sg13g2_a21o_2 _11784_ (.A2(_03921_),
    .A1(net3142),
    .B1(_03926_),
    .X(_03927_));
 sg13g2_a21oi_1 _11785_ (.A1(net3640),
    .A2(_03927_),
    .Y(_03928_),
    .B1(net3624));
 sg13g2_nor2b_1 _11786_ (.A(net3822),
    .B_N(\mem.mem[116][4] ),
    .Y(_03929_));
 sg13g2_a21oi_1 _11787_ (.A1(net3821),
    .A2(\mem.mem[117][4] ),
    .Y(_03930_),
    .B1(_03929_));
 sg13g2_nand2b_1 _11788_ (.Y(_03931_),
    .B(\mem.mem[118][4] ),
    .A_N(net3821));
 sg13g2_a21oi_1 _11789_ (.A1(net3821),
    .A2(\mem.mem[119][4] ),
    .Y(_03932_),
    .B1(net3187));
 sg13g2_a221oi_1 _11790_ (.B2(_03932_),
    .C1(net3134),
    .B1(_03931_),
    .A1(net3187),
    .Y(_03933_),
    .A2(_03930_));
 sg13g2_nor2b_1 _11791_ (.A(net3833),
    .B_N(\mem.mem[112][4] ),
    .Y(_03934_));
 sg13g2_a21oi_1 _11792_ (.A1(net3833),
    .A2(\mem.mem[113][4] ),
    .Y(_03935_),
    .B1(_03934_));
 sg13g2_nand2b_1 _11793_ (.Y(_03936_),
    .B(\mem.mem[114][4] ),
    .A_N(net3833));
 sg13g2_a21oi_1 _11794_ (.A1(net3833),
    .A2(\mem.mem[115][4] ),
    .Y(_03937_),
    .B1(net3191));
 sg13g2_a221oi_1 _11795_ (.B2(_03937_),
    .C1(net3670),
    .B1(_03936_),
    .A1(net3191),
    .Y(_03938_),
    .A2(_03935_));
 sg13g2_mux4_1 _11796_ (.S0(net3841),
    .A0(\mem.mem[120][4] ),
    .A1(\mem.mem[121][4] ),
    .A2(\mem.mem[122][4] ),
    .A3(\mem.mem[123][4] ),
    .S1(net3721),
    .X(_03939_));
 sg13g2_a21oi_1 _11797_ (.A1(net3844),
    .A2(\mem.mem[127][4] ),
    .Y(_03940_),
    .B1(net3192));
 sg13g2_o21ai_1 _11798_ (.B1(_03940_),
    .Y(_03941_),
    .A1(net3844),
    .A2(_02159_));
 sg13g2_nand2b_1 _11799_ (.Y(_03942_),
    .B(\mem.mem[124][4] ),
    .A_N(net3843));
 sg13g2_a21oi_1 _11800_ (.A1(net3842),
    .A2(\mem.mem[125][4] ),
    .Y(_03943_),
    .B1(net3722));
 sg13g2_a21oi_1 _11801_ (.A1(_03942_),
    .A2(_03943_),
    .Y(_03944_),
    .B1(net3140));
 sg13g2_nor3_2 _11802_ (.A(net3638),
    .B(_03933_),
    .C(_03938_),
    .Y(_03945_));
 sg13g2_a221oi_1 _11803_ (.B2(_03944_),
    .C1(net3109),
    .B1(_03941_),
    .A1(net3139),
    .Y(_03946_),
    .A2(_03939_));
 sg13g2_or2_1 _11804_ (.X(_03947_),
    .B(_03946_),
    .A(_03945_));
 sg13g2_a221oi_1 _11805_ (.B2(net3624),
    .C1(net3091),
    .B1(_03947_),
    .A1(_03920_),
    .Y(_03948_),
    .A2(_03928_));
 sg13g2_o21ai_1 _11806_ (.B1(net3612),
    .Y(_03949_),
    .A1(_03909_),
    .A2(_03948_));
 sg13g2_o21ai_1 _11807_ (.B1(_02148_),
    .Y(_03950_),
    .A1(_03839_),
    .A2(_03878_));
 sg13g2_nand3_1 _11808_ (.B(_03949_),
    .C(_03950_),
    .A(_02149_),
    .Y(_03951_));
 sg13g2_and2_1 _11809_ (.A(_03801_),
    .B(_03951_),
    .X(_03952_));
 sg13g2_a22oi_1 _11810_ (.Y(_03953_),
    .B1(_03952_),
    .B2(_02259_),
    .A2(_02536_),
    .A1(net5));
 sg13g2_o21ai_1 _11811_ (.B1(net4006),
    .Y(_03954_),
    .A1(net5193),
    .A2(net3055));
 sg13g2_a21oi_1 _11812_ (.A1(net3055),
    .A2(_03953_),
    .Y(_00599_),
    .B1(_03954_));
 sg13g2_mux2_1 _11813_ (.A0(\mem.mem[140][5] ),
    .A1(\mem.mem[141][5] ),
    .S(net3913),
    .X(_03955_));
 sg13g2_nand2_1 _11814_ (.Y(_03956_),
    .A(net3214),
    .B(_03955_));
 sg13g2_mux2_1 _11815_ (.A0(\mem.mem[142][5] ),
    .A1(\mem.mem[143][5] ),
    .S(net3912),
    .X(_03957_));
 sg13g2_a21oi_1 _11816_ (.A1(net3747),
    .A2(_03957_),
    .Y(_03958_),
    .B1(net3157));
 sg13g2_mux4_1 _11817_ (.S0(net3898),
    .A0(\mem.mem[136][5] ),
    .A1(\mem.mem[137][5] ),
    .A2(\mem.mem[138][5] ),
    .A3(\mem.mem[139][5] ),
    .S1(net3742),
    .X(_03959_));
 sg13g2_o21ai_1 _11818_ (.B1(net3647),
    .Y(_03960_),
    .A1(net3679),
    .A2(_03959_));
 sg13g2_a21oi_1 _11819_ (.A1(_03956_),
    .A2(_03958_),
    .Y(_03961_),
    .B1(_03960_));
 sg13g2_mux2_1 _11820_ (.A0(\mem.mem[134][5] ),
    .A1(\mem.mem[135][5] ),
    .S(net3891),
    .X(_03962_));
 sg13g2_mux2_1 _11821_ (.A0(\mem.mem[132][5] ),
    .A1(\mem.mem[133][5] ),
    .S(net3891),
    .X(_03963_));
 sg13g2_nand2_1 _11822_ (.Y(_03964_),
    .A(net3207),
    .B(_03963_));
 sg13g2_a21oi_1 _11823_ (.A1(net3739),
    .A2(_03962_),
    .Y(_03965_),
    .B1(net3152));
 sg13g2_mux2_1 _11824_ (.A0(\mem.mem[130][5] ),
    .A1(\mem.mem[131][5] ),
    .S(net3890),
    .X(_03966_));
 sg13g2_nand2_1 _11825_ (.Y(_03967_),
    .A(net3739),
    .B(_03966_));
 sg13g2_mux2_1 _11826_ (.A0(\mem.mem[128][5] ),
    .A1(\mem.mem[129][5] ),
    .S(net3886),
    .X(_03968_));
 sg13g2_a21oi_1 _11827_ (.A1(net3207),
    .A2(_03968_),
    .Y(_03969_),
    .B1(net3676));
 sg13g2_a221oi_1 _11828_ (.B2(_03969_),
    .C1(net3644),
    .B1(_03967_),
    .A1(_03964_),
    .Y(_03970_),
    .A2(_03965_));
 sg13g2_nor3_1 _11829_ (.A(net3629),
    .B(_03961_),
    .C(_03970_),
    .Y(_03971_));
 sg13g2_mux4_1 _11830_ (.S0(net3967),
    .A0(\mem.mem[144][5] ),
    .A1(\mem.mem[145][5] ),
    .A2(\mem.mem[146][5] ),
    .A3(\mem.mem[147][5] ),
    .S1(net3762),
    .X(_03972_));
 sg13g2_nor2_1 _11831_ (.A(net3687),
    .B(_03972_),
    .Y(_03973_));
 sg13g2_mux2_1 _11832_ (.A0(\mem.mem[150][5] ),
    .A1(\mem.mem[151][5] ),
    .S(net3972),
    .X(_03974_));
 sg13g2_nand2b_1 _11833_ (.Y(_03975_),
    .B(net3983),
    .A_N(\mem.mem[149][5] ));
 sg13g2_o21ai_1 _11834_ (.B1(_03975_),
    .Y(_03976_),
    .A1(net3983),
    .A2(\mem.mem[148][5] ));
 sg13g2_o21ai_1 _11835_ (.B1(net3688),
    .Y(_03977_),
    .A1(net3763),
    .A2(_03976_));
 sg13g2_a21oi_1 _11836_ (.A1(net3763),
    .A2(_03974_),
    .Y(_03978_),
    .B1(_03977_));
 sg13g2_nor3_1 _11837_ (.A(net3651),
    .B(_03973_),
    .C(_03978_),
    .Y(_03979_));
 sg13g2_mux4_1 _11838_ (.S0(net3982),
    .A0(\mem.mem[152][5] ),
    .A1(\mem.mem[153][5] ),
    .A2(\mem.mem[154][5] ),
    .A3(\mem.mem[155][5] ),
    .S1(net3768),
    .X(_03980_));
 sg13g2_nor2_2 _11839_ (.A(net3688),
    .B(_03980_),
    .Y(_03981_));
 sg13g2_nor2b_1 _11840_ (.A(\mem.mem[157][5] ),
    .B_N(net3921),
    .Y(_03982_));
 sg13g2_nor2_1 _11841_ (.A(net3921),
    .B(\mem.mem[156][5] ),
    .Y(_03983_));
 sg13g2_nor3_1 _11842_ (.A(net3749),
    .B(_03982_),
    .C(_03983_),
    .Y(_03984_));
 sg13g2_nor2b_1 _11843_ (.A(\mem.mem[159][5] ),
    .B_N(net3921),
    .Y(_03985_));
 sg13g2_o21ai_1 _11844_ (.B1(net3749),
    .Y(_03986_),
    .A1(net3921),
    .A2(\mem.mem[158][5] ));
 sg13g2_o21ai_1 _11845_ (.B1(net3679),
    .Y(_03987_),
    .A1(_03985_),
    .A2(_03986_));
 sg13g2_o21ai_1 _11846_ (.B1(net3651),
    .Y(_03988_),
    .A1(_03984_),
    .A2(_03987_));
 sg13g2_o21ai_1 _11847_ (.B1(net3629),
    .Y(_03989_),
    .A1(_03981_),
    .A2(_03988_));
 sg13g2_o21ai_1 _11848_ (.B1(net3092),
    .Y(_03990_),
    .A1(_03979_),
    .A2(_03989_));
 sg13g2_nand2b_1 _11849_ (.Y(_03991_),
    .B(\mem.mem[166][5] ),
    .A_N(net3874));
 sg13g2_a21oi_1 _11850_ (.A1(net3874),
    .A2(\mem.mem[167][5] ),
    .Y(_03992_),
    .B1(net3203));
 sg13g2_nor2b_1 _11851_ (.A(net3895),
    .B_N(\mem.mem[164][5] ),
    .Y(_03993_));
 sg13g2_a21oi_1 _11852_ (.A1(net3895),
    .A2(\mem.mem[165][5] ),
    .Y(_03994_),
    .B1(_03993_));
 sg13g2_a221oi_1 _11853_ (.B2(net3203),
    .C1(net3149),
    .B1(_03994_),
    .A1(_03991_),
    .Y(_03995_),
    .A2(_03992_));
 sg13g2_nor2b_1 _11854_ (.A(net3877),
    .B_N(\mem.mem[160][5] ),
    .Y(_03996_));
 sg13g2_a21oi_1 _11855_ (.A1(net3877),
    .A2(\mem.mem[161][5] ),
    .Y(_03997_),
    .B1(_03996_));
 sg13g2_nand2b_1 _11856_ (.Y(_03998_),
    .B(\mem.mem[162][5] ),
    .A_N(net3872));
 sg13g2_a21oi_1 _11857_ (.A1(net3873),
    .A2(\mem.mem[163][5] ),
    .Y(_03999_),
    .B1(net3203));
 sg13g2_a221oi_1 _11858_ (.B2(_03999_),
    .C1(net3675),
    .B1(_03998_),
    .A1(net3203),
    .Y(_04000_),
    .A2(_03997_));
 sg13g2_nor3_2 _11859_ (.A(net3643),
    .B(_03995_),
    .C(_04000_),
    .Y(_04001_));
 sg13g2_mux4_1 _11860_ (.S0(net3849),
    .A0(\mem.mem[168][5] ),
    .A1(\mem.mem[169][5] ),
    .A2(\mem.mem[170][5] ),
    .A3(\mem.mem[171][5] ),
    .S1(net3725),
    .X(_04002_));
 sg13g2_mux2_1 _11861_ (.A0(\mem.mem[172][5] ),
    .A1(\mem.mem[173][5] ),
    .S(net3833),
    .X(_04003_));
 sg13g2_o21ai_1 _11862_ (.B1(net3726),
    .Y(_04004_),
    .A1(net3851),
    .A2(_02162_));
 sg13g2_a21oi_1 _11863_ (.A1(net3851),
    .A2(\mem.mem[175][5] ),
    .Y(_04005_),
    .B1(_04004_));
 sg13g2_o21ai_1 _11864_ (.B1(net3669),
    .Y(_04006_),
    .A1(net3719),
    .A2(_04003_));
 sg13g2_o21ai_1 _11865_ (.B1(net3640),
    .Y(_04007_),
    .A1(_04005_),
    .A2(_04006_));
 sg13g2_a21oi_1 _11866_ (.A1(net3144),
    .A2(_04002_),
    .Y(_04008_),
    .B1(_04007_));
 sg13g2_o21ai_1 _11867_ (.B1(net3095),
    .Y(_04009_),
    .A1(_04001_),
    .A2(_04008_));
 sg13g2_nor2b_1 _11868_ (.A(net3860),
    .B_N(\mem.mem[180][5] ),
    .Y(_04010_));
 sg13g2_a21oi_1 _11869_ (.A1(net3860),
    .A2(\mem.mem[181][5] ),
    .Y(_04011_),
    .B1(_04010_));
 sg13g2_nand2b_1 _11870_ (.Y(_04012_),
    .B(\mem.mem[182][5] ),
    .A_N(net3859));
 sg13g2_a21oi_1 _11871_ (.A1(net3855),
    .A2(\mem.mem[183][5] ),
    .Y(_04013_),
    .B1(net3193));
 sg13g2_a221oi_1 _11872_ (.B2(_04013_),
    .C1(net3141),
    .B1(_04012_),
    .A1(net3193),
    .Y(_04014_),
    .A2(_04011_));
 sg13g2_nor2b_1 _11873_ (.A(net3850),
    .B_N(\mem.mem[176][5] ),
    .Y(_04015_));
 sg13g2_a21oi_1 _11874_ (.A1(net3850),
    .A2(\mem.mem[177][5] ),
    .Y(_04016_),
    .B1(_04015_));
 sg13g2_nand2b_1 _11875_ (.Y(_04017_),
    .B(\mem.mem[178][5] ),
    .A_N(net3854));
 sg13g2_a21oi_1 _11876_ (.A1(net3854),
    .A2(\mem.mem[179][5] ),
    .Y(_04018_),
    .B1(net3193));
 sg13g2_a221oi_1 _11877_ (.B2(_04018_),
    .C1(net3672),
    .B1(_04017_),
    .A1(net3193),
    .Y(_04019_),
    .A2(_04016_));
 sg13g2_nor3_1 _11878_ (.A(net3640),
    .B(_04014_),
    .C(_04019_),
    .Y(_04020_));
 sg13g2_mux4_1 _11879_ (.S0(net3848),
    .A0(\mem.mem[184][5] ),
    .A1(\mem.mem[185][5] ),
    .A2(\mem.mem[186][5] ),
    .A3(\mem.mem[187][5] ),
    .S1(net3724),
    .X(_04021_));
 sg13g2_a21oi_1 _11880_ (.A1(net3847),
    .A2(\mem.mem[191][5] ),
    .Y(_04022_),
    .B1(net3192));
 sg13g2_o21ai_1 _11881_ (.B1(_04022_),
    .Y(_04023_),
    .A1(net3847),
    .A2(_02163_));
 sg13g2_nand2b_1 _11882_ (.Y(_04024_),
    .B(\mem.mem[188][5] ),
    .A_N(net3847));
 sg13g2_a21oi_1 _11883_ (.A1(net3847),
    .A2(\mem.mem[189][5] ),
    .Y(_04025_),
    .B1(net3723));
 sg13g2_a21oi_1 _11884_ (.A1(_04024_),
    .A2(_04025_),
    .Y(_04026_),
    .B1(net3140));
 sg13g2_a221oi_1 _11885_ (.B2(_04026_),
    .C1(net3109),
    .B1(_04023_),
    .A1(net3140),
    .Y(_04027_),
    .A2(_04021_));
 sg13g2_o21ai_1 _11886_ (.B1(net3622),
    .Y(_04028_),
    .A1(_04020_),
    .A2(_04027_));
 sg13g2_nand3_1 _11887_ (.B(_04009_),
    .C(_04028_),
    .A(net3616),
    .Y(_04029_));
 sg13g2_o21ai_1 _11888_ (.B1(_02148_),
    .Y(_04030_),
    .A1(_03971_),
    .A2(_03990_));
 sg13g2_nor2b_1 _11889_ (.A(_04030_),
    .B_N(_04029_),
    .Y(_04031_));
 sg13g2_mux2_1 _11890_ (.A0(\mem.mem[214][5] ),
    .A1(\mem.mem[215][5] ),
    .S(net3790),
    .X(_04032_));
 sg13g2_nand2_1 _11891_ (.Y(_04033_),
    .A(net3698),
    .B(_04032_));
 sg13g2_mux2_1 _11892_ (.A0(\mem.mem[212][5] ),
    .A1(\mem.mem[213][5] ),
    .S(net3790),
    .X(_04034_));
 sg13g2_a21oi_1 _11893_ (.A1(net3178),
    .A2(_04034_),
    .Y(_04035_),
    .B1(net3125));
 sg13g2_mux2_1 _11894_ (.A0(\mem.mem[210][5] ),
    .A1(\mem.mem[211][5] ),
    .S(net3784),
    .X(_04036_));
 sg13g2_nand2_1 _11895_ (.Y(_04037_),
    .A(net3697),
    .B(_04036_));
 sg13g2_mux2_1 _11896_ (.A0(\mem.mem[208][5] ),
    .A1(\mem.mem[209][5] ),
    .S(net3784),
    .X(_04038_));
 sg13g2_a21oi_1 _11897_ (.A1(net3178),
    .A2(_04038_),
    .Y(_04039_),
    .B1(net3659));
 sg13g2_a221oi_1 _11898_ (.B2(_04039_),
    .C1(net3632),
    .B1(_04037_),
    .A1(_04033_),
    .Y(_04040_),
    .A2(_04035_));
 sg13g2_mux4_1 _11899_ (.S0(net3788),
    .A0(\mem.mem[216][5] ),
    .A1(\mem.mem[217][5] ),
    .A2(\mem.mem[218][5] ),
    .A3(\mem.mem[219][5] ),
    .S1(net3696),
    .X(_04041_));
 sg13g2_nor2_1 _11900_ (.A(net3659),
    .B(_04041_),
    .Y(_04042_));
 sg13g2_nor2b_1 _11901_ (.A(\mem.mem[221][5] ),
    .B_N(net3787),
    .Y(_04043_));
 sg13g2_nor2_1 _11902_ (.A(net3787),
    .B(\mem.mem[220][5] ),
    .Y(_04044_));
 sg13g2_nor3_1 _11903_ (.A(net3696),
    .B(_04043_),
    .C(_04044_),
    .Y(_04045_));
 sg13g2_nor2b_1 _11904_ (.A(\mem.mem[223][5] ),
    .B_N(net3787),
    .Y(_04046_));
 sg13g2_o21ai_1 _11905_ (.B1(net3697),
    .Y(_04047_),
    .A1(net3787),
    .A2(\mem.mem[222][5] ));
 sg13g2_o21ai_1 _11906_ (.B1(net3659),
    .Y(_04048_),
    .A1(_04046_),
    .A2(_04047_));
 sg13g2_o21ai_1 _11907_ (.B1(net3637),
    .Y(_04049_),
    .A1(_04045_),
    .A2(_04048_));
 sg13g2_o21ai_1 _11908_ (.B1(net3621),
    .Y(_04050_),
    .A1(_04042_),
    .A2(_04049_));
 sg13g2_mux2_1 _11909_ (.A0(\mem.mem[204][5] ),
    .A1(\mem.mem[205][5] ),
    .S(net3777),
    .X(_04051_));
 sg13g2_nand2_1 _11910_ (.Y(_04052_),
    .A(net3177),
    .B(_04051_));
 sg13g2_mux2_1 _11911_ (.A0(\mem.mem[206][5] ),
    .A1(\mem.mem[207][5] ),
    .S(net3781),
    .X(_04053_));
 sg13g2_a21oi_1 _11912_ (.A1(net3693),
    .A2(_04053_),
    .Y(_04054_),
    .B1(net3123));
 sg13g2_mux4_1 _11913_ (.S0(net3777),
    .A0(\mem.mem[200][5] ),
    .A1(\mem.mem[201][5] ),
    .A2(\mem.mem[202][5] ),
    .A3(\mem.mem[203][5] ),
    .S1(net3693),
    .X(_04055_));
 sg13g2_o21ai_1 _11914_ (.B1(net3633),
    .Y(_04056_),
    .A1(net3658),
    .A2(_04055_));
 sg13g2_a21oi_1 _11915_ (.A1(_04052_),
    .A2(_04054_),
    .Y(_04057_),
    .B1(_04056_));
 sg13g2_mux2_1 _11916_ (.A0(\mem.mem[198][5] ),
    .A1(\mem.mem[199][5] ),
    .S(net3771),
    .X(_04058_));
 sg13g2_mux2_1 _11917_ (.A0(\mem.mem[196][5] ),
    .A1(\mem.mem[197][5] ),
    .S(net3771),
    .X(_04059_));
 sg13g2_nand2_1 _11918_ (.Y(_04060_),
    .A(net3175),
    .B(_04059_));
 sg13g2_a21oi_1 _11919_ (.A1(net3691),
    .A2(_04058_),
    .Y(_04061_),
    .B1(net3121));
 sg13g2_mux2_1 _11920_ (.A0(\mem.mem[194][5] ),
    .A1(\mem.mem[195][5] ),
    .S(net3771),
    .X(_04062_));
 sg13g2_nand2_1 _11921_ (.Y(_04063_),
    .A(net3691),
    .B(_04062_));
 sg13g2_mux2_1 _11922_ (.A0(\mem.mem[192][5] ),
    .A1(\mem.mem[193][5] ),
    .S(net3773),
    .X(_04064_));
 sg13g2_a21oi_1 _11923_ (.A1(net3175),
    .A2(_04064_),
    .Y(_04065_),
    .B1(net3657));
 sg13g2_a221oi_1 _11924_ (.B2(_04065_),
    .C1(net3632),
    .B1(_04063_),
    .A1(_04060_),
    .Y(_04066_),
    .A2(_04061_));
 sg13g2_nor3_2 _11925_ (.A(net3620),
    .B(_04057_),
    .C(_04066_),
    .Y(_04067_));
 sg13g2_o21ai_1 _11926_ (.B1(net3090),
    .Y(_04068_),
    .A1(_04040_),
    .A2(_04050_));
 sg13g2_nor2_2 _11927_ (.A(_04067_),
    .B(_04068_),
    .Y(_04069_));
 sg13g2_mux2_1 _11928_ (.A0(\mem.mem[236][5] ),
    .A1(\mem.mem[237][5] ),
    .S(net3831),
    .X(_04070_));
 sg13g2_nand2_1 _11929_ (.Y(_04071_),
    .A(net3190),
    .B(_04070_));
 sg13g2_mux2_1 _11930_ (.A0(\mem.mem[238][5] ),
    .A1(\mem.mem[239][5] ),
    .S(net3830),
    .X(_04072_));
 sg13g2_a21oi_1 _11931_ (.A1(net3716),
    .A2(_04072_),
    .Y(_04073_),
    .B1(net3136));
 sg13g2_mux4_1 _11932_ (.S0(net3832),
    .A0(\mem.mem[232][5] ),
    .A1(\mem.mem[233][5] ),
    .A2(\mem.mem[234][5] ),
    .A3(\mem.mem[235][5] ),
    .S1(net3716),
    .X(_04074_));
 sg13g2_o21ai_1 _11933_ (.B1(net3638),
    .Y(_04075_),
    .A1(net3668),
    .A2(_04074_));
 sg13g2_a21oi_1 _11934_ (.A1(_04071_),
    .A2(_04073_),
    .Y(_04076_),
    .B1(_04075_));
 sg13g2_mux2_1 _11935_ (.A0(\mem.mem[230][5] ),
    .A1(\mem.mem[231][5] ),
    .S(net3868),
    .X(_04077_));
 sg13g2_mux2_1 _11936_ (.A0(\mem.mem[228][5] ),
    .A1(\mem.mem[229][5] ),
    .S(net3879),
    .X(_04078_));
 sg13g2_nand2_1 _11937_ (.Y(_04079_),
    .A(net3205),
    .B(_04078_));
 sg13g2_a21oi_1 _11938_ (.A1(net3732),
    .A2(_04077_),
    .Y(_04080_),
    .B1(net3147));
 sg13g2_mux2_1 _11939_ (.A0(\mem.mem[226][5] ),
    .A1(\mem.mem[227][5] ),
    .S(net3867),
    .X(_04081_));
 sg13g2_nand2_1 _11940_ (.Y(_04082_),
    .A(net3732),
    .B(_04081_));
 sg13g2_mux2_1 _11941_ (.A0(\mem.mem[224][5] ),
    .A1(\mem.mem[225][5] ),
    .S(net3867),
    .X(_04083_));
 sg13g2_a21oi_1 _11942_ (.A1(net3200),
    .A2(_04083_),
    .Y(_04084_),
    .B1(net3674));
 sg13g2_a221oi_1 _11943_ (.B2(_04084_),
    .C1(net3643),
    .B1(_04082_),
    .A1(_04079_),
    .Y(_04085_),
    .A2(_04080_));
 sg13g2_nor3_2 _11944_ (.A(net3625),
    .B(_04076_),
    .C(_04085_),
    .Y(_04086_));
 sg13g2_mux4_1 _11945_ (.S0(net3829),
    .A0(\mem.mem[244][5] ),
    .A1(\mem.mem[245][5] ),
    .A2(\mem.mem[246][5] ),
    .A3(\mem.mem[247][5] ),
    .S1(net3715),
    .X(_04087_));
 sg13g2_inv_1 _11946_ (.Y(_04088_),
    .A(_04087_));
 sg13g2_mux4_1 _11947_ (.S0(net3827),
    .A0(\mem.mem[240][5] ),
    .A1(\mem.mem[241][5] ),
    .A2(\mem.mem[242][5] ),
    .A3(\mem.mem[243][5] ),
    .S1(net3715),
    .X(_04089_));
 sg13g2_o21ai_1 _11948_ (.B1(net3107),
    .Y(_04090_),
    .A1(net3668),
    .A2(_04089_));
 sg13g2_a21oi_1 _11949_ (.A1(net3668),
    .A2(_04088_),
    .Y(_04091_),
    .B1(_04090_));
 sg13g2_nand2b_1 _11950_ (.Y(_04092_),
    .B(net3668),
    .A_N(\mem.mem[252][5] ));
 sg13g2_mux4_1 _11951_ (.S0(net3825),
    .A0(\mem.mem[248][5] ),
    .A1(\mem.mem[249][5] ),
    .A2(\mem.mem[250][5] ),
    .A3(\mem.mem[251][5] ),
    .S1(net3720),
    .X(_04093_));
 sg13g2_o21ai_1 _11952_ (.B1(_04092_),
    .Y(_04094_),
    .A1(net3667),
    .A2(_04093_));
 sg13g2_o21ai_1 _11953_ (.B1(net3623),
    .Y(_04095_),
    .A1(net3106),
    .A2(_04094_));
 sg13g2_o21ai_1 _11954_ (.B1(net3617),
    .Y(_04096_),
    .A1(_04091_),
    .A2(_04095_));
 sg13g2_o21ai_1 _11955_ (.B1(net3612),
    .Y(_04097_),
    .A1(_04086_),
    .A2(_04096_));
 sg13g2_nor2_2 _11956_ (.A(_04069_),
    .B(_04097_),
    .Y(_04098_));
 sg13g2_o21ai_1 _11957_ (.B1(net3611),
    .Y(_04099_),
    .A1(_04031_),
    .A2(_04098_));
 sg13g2_nand2b_1 _11958_ (.Y(_04100_),
    .B(\mem.mem[38][5] ),
    .A_N(net3948));
 sg13g2_a21oi_1 _11959_ (.A1(net3948),
    .A2(\mem.mem[39][5] ),
    .Y(_04101_),
    .B1(net3224));
 sg13g2_nor2b_1 _11960_ (.A(net3948),
    .B_N(\mem.mem[36][5] ),
    .Y(_04102_));
 sg13g2_a21oi_1 _11961_ (.A1(net3949),
    .A2(\mem.mem[37][5] ),
    .Y(_04103_),
    .B1(_04102_));
 sg13g2_a221oi_1 _11962_ (.B2(net3224),
    .C1(net3163),
    .B1(_04103_),
    .A1(_04100_),
    .Y(_04104_),
    .A2(_04101_));
 sg13g2_nor2b_1 _11963_ (.A(net3935),
    .B_N(\mem.mem[32][5] ),
    .Y(_04105_));
 sg13g2_a21oi_1 _11964_ (.A1(net3935),
    .A2(\mem.mem[33][5] ),
    .Y(_04106_),
    .B1(_04105_));
 sg13g2_nand2b_1 _11965_ (.Y(_04107_),
    .B(\mem.mem[34][5] ),
    .A_N(net3936));
 sg13g2_a21oi_1 _11966_ (.A1(net3936),
    .A2(\mem.mem[35][5] ),
    .Y(_04108_),
    .B1(net3220));
 sg13g2_a221oi_1 _11967_ (.B2(_04108_),
    .C1(net3685),
    .B1(_04107_),
    .A1(net3220),
    .Y(_04109_),
    .A2(_04106_));
 sg13g2_o21ai_1 _11968_ (.B1(net3115),
    .Y(_04110_),
    .A1(_04104_),
    .A2(_04109_));
 sg13g2_mux4_1 _11969_ (.S0(net3979),
    .A0(\mem.mem[40][5] ),
    .A1(\mem.mem[41][5] ),
    .A2(\mem.mem[42][5] ),
    .A3(\mem.mem[43][5] ),
    .S1(net3765),
    .X(_04111_));
 sg13g2_nand2_1 _11970_ (.Y(_04112_),
    .A(net3171),
    .B(_04111_));
 sg13g2_mux2_1 _11971_ (.A0(\mem.mem[44][5] ),
    .A1(\mem.mem[45][5] ),
    .S(net3975),
    .X(_04113_));
 sg13g2_mux2_1 _11972_ (.A0(\mem.mem[46][5] ),
    .A1(\mem.mem[47][5] ),
    .S(net3974),
    .X(_04114_));
 sg13g2_nor2_1 _11973_ (.A(net3233),
    .B(_04114_),
    .Y(_04115_));
 sg13g2_o21ai_1 _11974_ (.B1(net3689),
    .Y(_04116_),
    .A1(net3766),
    .A2(_04113_));
 sg13g2_o21ai_1 _11975_ (.B1(_04112_),
    .Y(_04117_),
    .A1(_04115_),
    .A2(_04116_));
 sg13g2_a21oi_1 _11976_ (.A1(net3653),
    .A2(_04117_),
    .Y(_04118_),
    .B1(net3627));
 sg13g2_nor2b_1 _11977_ (.A(net3962),
    .B_N(\mem.mem[52][5] ),
    .Y(_04119_));
 sg13g2_a21oi_1 _11978_ (.A1(net3962),
    .A2(\mem.mem[53][5] ),
    .Y(_04120_),
    .B1(_04119_));
 sg13g2_nand2b_1 _11979_ (.Y(_04121_),
    .B(\mem.mem[54][5] ),
    .A_N(net3962));
 sg13g2_a21oi_1 _11980_ (.A1(net3962),
    .A2(\mem.mem[55][5] ),
    .Y(_04122_),
    .B1(net3233));
 sg13g2_a221oi_1 _11981_ (.B2(_04122_),
    .C1(net3166),
    .B1(_04121_),
    .A1(net3232),
    .Y(_04123_),
    .A2(_04120_));
 sg13g2_nor2b_1 _11982_ (.A(net3961),
    .B_N(\mem.mem[48][5] ),
    .Y(_04124_));
 sg13g2_a21oi_1 _11983_ (.A1(net3961),
    .A2(\mem.mem[49][5] ),
    .Y(_04125_),
    .B1(_04124_));
 sg13g2_nand2b_1 _11984_ (.Y(_04126_),
    .B(\mem.mem[50][5] ),
    .A_N(net3961));
 sg13g2_a21oi_1 _11985_ (.A1(net3961),
    .A2(\mem.mem[51][5] ),
    .Y(_04127_),
    .B1(net3229));
 sg13g2_a221oi_1 _11986_ (.B2(_04127_),
    .C1(net3686),
    .B1(_04126_),
    .A1(net3229),
    .Y(_04128_),
    .A2(_04125_));
 sg13g2_mux4_1 _11987_ (.S0(net3980),
    .A0(\mem.mem[56][5] ),
    .A1(\mem.mem[57][5] ),
    .A2(\mem.mem[58][5] ),
    .A3(\mem.mem[59][5] ),
    .S1(net3765),
    .X(_04129_));
 sg13g2_a21oi_1 _11988_ (.A1(net3978),
    .A2(\mem.mem[63][5] ),
    .Y(_04130_),
    .B1(net3235));
 sg13g2_o21ai_1 _11989_ (.B1(_04130_),
    .Y(_04131_),
    .A1(net3978),
    .A2(_02161_));
 sg13g2_nand2b_1 _11990_ (.Y(_04132_),
    .B(\mem.mem[60][5] ),
    .A_N(net3978));
 sg13g2_a21oi_1 _11991_ (.A1(net3978),
    .A2(\mem.mem[61][5] ),
    .Y(_04133_),
    .B1(net3765));
 sg13g2_a21oi_1 _11992_ (.A1(_04132_),
    .A2(_04133_),
    .Y(_04134_),
    .B1(net3171));
 sg13g2_nor3_1 _11993_ (.A(net3653),
    .B(_04123_),
    .C(_04128_),
    .Y(_04135_));
 sg13g2_a221oi_1 _11994_ (.B2(_04134_),
    .C1(net3118),
    .B1(_04131_),
    .A1(net3171),
    .Y(_04136_),
    .A2(_04129_));
 sg13g2_o21ai_1 _11995_ (.B1(net3630),
    .Y(_04137_),
    .A1(_04135_),
    .A2(_04136_));
 sg13g2_a21oi_1 _11996_ (.A1(_04110_),
    .A2(_04118_),
    .Y(_04138_),
    .B1(net3092));
 sg13g2_nand2_2 _11997_ (.Y(_04139_),
    .A(_04137_),
    .B(_04138_));
 sg13g2_mux4_1 _11998_ (.S0(net3947),
    .A0(\mem.mem[28][5] ),
    .A1(\mem.mem[29][5] ),
    .A2(\mem.mem[30][5] ),
    .A3(\mem.mem[31][5] ),
    .S1(net3757),
    .X(_04140_));
 sg13g2_mux4_1 _11999_ (.S0(net3944),
    .A0(\mem.mem[24][5] ),
    .A1(\mem.mem[25][5] ),
    .A2(\mem.mem[26][5] ),
    .A3(\mem.mem[27][5] ),
    .S1(net3756),
    .X(_04141_));
 sg13g2_nor2_1 _12000_ (.A(net3683),
    .B(_04141_),
    .Y(_04142_));
 sg13g2_nor2_1 _12001_ (.A(net3115),
    .B(_04142_),
    .Y(_04143_));
 sg13g2_o21ai_1 _12002_ (.B1(_04143_),
    .Y(_04144_),
    .A1(net3161),
    .A2(_04140_));
 sg13g2_mux4_1 _12003_ (.S0(net3943),
    .A0(\mem.mem[20][5] ),
    .A1(\mem.mem[21][5] ),
    .A2(\mem.mem[22][5] ),
    .A3(\mem.mem[23][5] ),
    .S1(net3756),
    .X(_04145_));
 sg13g2_mux4_1 _12004_ (.S0(net3928),
    .A0(\mem.mem[16][5] ),
    .A1(\mem.mem[17][5] ),
    .A2(\mem.mem[18][5] ),
    .A3(\mem.mem[19][5] ),
    .S1(net3751),
    .X(_04146_));
 sg13g2_mux2_1 _12005_ (.A0(_04145_),
    .A1(_04146_),
    .S(net3161),
    .X(_04147_));
 sg13g2_a21oi_1 _12006_ (.A1(net3115),
    .A2(_04147_),
    .Y(_04148_),
    .B1(net3098));
 sg13g2_mux2_1 _12007_ (.A0(\mem.mem[6][5] ),
    .A1(\mem.mem[7][5] ),
    .S(net3883),
    .X(_04149_));
 sg13g2_nand2_1 _12008_ (.Y(_04150_),
    .A(net3737),
    .B(_04149_));
 sg13g2_mux2_1 _12009_ (.A0(\mem.mem[4][5] ),
    .A1(\mem.mem[5][5] ),
    .S(net3885),
    .X(_04151_));
 sg13g2_a21oi_1 _12010_ (.A1(net3205),
    .A2(_04151_),
    .Y(_04152_),
    .B1(net3150));
 sg13g2_mux2_1 _12011_ (.A0(\mem.mem[2][5] ),
    .A1(\mem.mem[3][5] ),
    .S(net3883),
    .X(_04153_));
 sg13g2_nand2_1 _12012_ (.Y(_04154_),
    .A(net3737),
    .B(_04153_));
 sg13g2_mux2_1 _12013_ (.A0(\mem.mem[0][5] ),
    .A1(\mem.mem[1][5] ),
    .S(net3885),
    .X(_04155_));
 sg13g2_a21oi_1 _12014_ (.A1(net3219),
    .A2(_04155_),
    .Y(_04156_),
    .B1(net3682));
 sg13g2_a221oi_1 _12015_ (.B2(_04156_),
    .C1(net3650),
    .B1(_04154_),
    .A1(_04150_),
    .Y(_04157_),
    .A2(_04152_));
 sg13g2_mux2_1 _12016_ (.A0(\mem.mem[12][5] ),
    .A1(\mem.mem[13][5] ),
    .S(net3931),
    .X(_04158_));
 sg13g2_nor2b_1 _12017_ (.A(\mem.mem[15][5] ),
    .B_N(net3931),
    .Y(_04159_));
 sg13g2_o21ai_1 _12018_ (.B1(net3753),
    .Y(_04160_),
    .A1(net3931),
    .A2(\mem.mem[14][5] ));
 sg13g2_o21ai_1 _12019_ (.B1(net3682),
    .Y(_04161_),
    .A1(_04159_),
    .A2(_04160_));
 sg13g2_a21oi_1 _12020_ (.A1(net3220),
    .A2(_04158_),
    .Y(_04162_),
    .B1(_04161_));
 sg13g2_mux4_1 _12021_ (.S0(net3887),
    .A0(\mem.mem[8][5] ),
    .A1(\mem.mem[9][5] ),
    .A2(\mem.mem[10][5] ),
    .A3(\mem.mem[11][5] ),
    .S1(net3739),
    .X(_04163_));
 sg13g2_o21ai_1 _12022_ (.B1(net3650),
    .Y(_04164_),
    .A1(net3681),
    .A2(_04163_));
 sg13g2_o21ai_1 _12023_ (.B1(net3098),
    .Y(_04165_),
    .A1(_04162_),
    .A2(_04164_));
 sg13g2_a21oi_2 _12024_ (.B1(net3618),
    .Y(_04166_),
    .A2(_04148_),
    .A1(_04144_));
 sg13g2_o21ai_1 _12025_ (.B1(_04166_),
    .Y(_04167_),
    .A1(_04157_),
    .A2(_04165_));
 sg13g2_mux4_1 _12026_ (.S0(net3778),
    .A0(\mem.mem[72][5] ),
    .A1(\mem.mem[73][5] ),
    .A2(\mem.mem[74][5] ),
    .A3(\mem.mem[75][5] ),
    .S1(net3694),
    .X(_04168_));
 sg13g2_mux4_1 _12027_ (.S0(net3797),
    .A0(\mem.mem[76][5] ),
    .A1(\mem.mem[77][5] ),
    .A2(\mem.mem[78][5] ),
    .A3(\mem.mem[79][5] ),
    .S1(net3702),
    .X(_04169_));
 sg13g2_inv_1 _12028_ (.Y(_04170_),
    .A(_04169_));
 sg13g2_o21ai_1 _12029_ (.B1(net3634),
    .Y(_04171_),
    .A1(net3661),
    .A2(_04168_));
 sg13g2_a21oi_2 _12030_ (.B1(_04171_),
    .Y(_04172_),
    .A2(_04170_),
    .A1(net3661));
 sg13g2_mux2_1 _12031_ (.A0(\mem.mem[70][5] ),
    .A1(\mem.mem[71][5] ),
    .S(net3812),
    .X(_04173_));
 sg13g2_nand2_1 _12032_ (.Y(_04174_),
    .A(net3708),
    .B(_04173_));
 sg13g2_mux2_1 _12033_ (.A0(\mem.mem[68][5] ),
    .A1(\mem.mem[69][5] ),
    .S(net3812),
    .X(_04175_));
 sg13g2_a21oi_1 _12034_ (.A1(net3185),
    .A2(_04175_),
    .Y(_04176_),
    .B1(net3132));
 sg13g2_mux2_1 _12035_ (.A0(\mem.mem[66][5] ),
    .A1(\mem.mem[67][5] ),
    .S(net3812),
    .X(_04177_));
 sg13g2_nand2_1 _12036_ (.Y(_04178_),
    .A(net3709),
    .B(_04177_));
 sg13g2_mux2_1 _12037_ (.A0(\mem.mem[64][5] ),
    .A1(\mem.mem[65][5] ),
    .S(net3795),
    .X(_04179_));
 sg13g2_a21oi_1 _12038_ (.A1(net3185),
    .A2(_04179_),
    .Y(_04180_),
    .B1(net3664));
 sg13g2_a221oi_1 _12039_ (.B2(_04180_),
    .C1(net3636),
    .B1(_04178_),
    .A1(_04174_),
    .Y(_04181_),
    .A2(_04176_));
 sg13g2_nor3_1 _12040_ (.A(net3621),
    .B(_04172_),
    .C(_04181_),
    .Y(_04182_));
 sg13g2_mux4_1 _12041_ (.S0(net3815),
    .A0(\mem.mem[84][5] ),
    .A1(\mem.mem[85][5] ),
    .A2(\mem.mem[86][5] ),
    .A3(\mem.mem[87][5] ),
    .S1(net3710),
    .X(_04183_));
 sg13g2_mux4_1 _12042_ (.S0(net3803),
    .A0(\mem.mem[80][5] ),
    .A1(\mem.mem[81][5] ),
    .A2(\mem.mem[82][5] ),
    .A3(\mem.mem[83][5] ),
    .S1(net3705),
    .X(_04184_));
 sg13g2_mux2_1 _12043_ (.A0(_04183_),
    .A1(_04184_),
    .S(net3130),
    .X(_04185_));
 sg13g2_mux4_1 _12044_ (.S0(net3803),
    .A0(\mem.mem[88][5] ),
    .A1(\mem.mem[89][5] ),
    .A2(\mem.mem[90][5] ),
    .A3(\mem.mem[91][5] ),
    .S1(net3705),
    .X(_04186_));
 sg13g2_nand2b_1 _12045_ (.Y(_04187_),
    .B(net3130),
    .A_N(_04186_));
 sg13g2_mux2_1 _12046_ (.A0(\mem.mem[92][5] ),
    .A1(\mem.mem[93][5] ),
    .S(net3814),
    .X(_04188_));
 sg13g2_nand2_1 _12047_ (.Y(_04189_),
    .A(net3183),
    .B(_04188_));
 sg13g2_mux2_1 _12048_ (.A0(\mem.mem[94][5] ),
    .A1(\mem.mem[95][5] ),
    .S(net3804),
    .X(_04190_));
 sg13g2_a21oi_1 _12049_ (.A1(net3707),
    .A2(_04190_),
    .Y(_04191_),
    .B1(net3129));
 sg13g2_a21oi_1 _12050_ (.A1(_04189_),
    .A2(_04191_),
    .Y(_04192_),
    .B1(net3103));
 sg13g2_a221oi_1 _12051_ (.B2(_04192_),
    .C1(net3094),
    .B1(_04187_),
    .A1(net3103),
    .Y(_04193_),
    .A2(_04185_));
 sg13g2_nor3_2 _12052_ (.A(net3615),
    .B(_04182_),
    .C(_04193_),
    .Y(_04194_));
 sg13g2_nand2b_1 _12053_ (.Y(_04195_),
    .B(net3915),
    .A_N(\mem.mem[103][5] ));
 sg13g2_o21ai_1 _12054_ (.B1(_04195_),
    .Y(_04196_),
    .A1(net3915),
    .A2(\mem.mem[102][5] ));
 sg13g2_mux2_1 _12055_ (.A0(\mem.mem[100][5] ),
    .A1(\mem.mem[101][5] ),
    .S(net3922),
    .X(_04197_));
 sg13g2_a21oi_1 _12056_ (.A1(net3216),
    .A2(_04197_),
    .Y(_04198_),
    .B1(net3158));
 sg13g2_o21ai_1 _12057_ (.B1(_04198_),
    .Y(_04199_),
    .A1(net3215),
    .A2(_04196_));
 sg13g2_mux2_1 _12058_ (.A0(\mem.mem[98][5] ),
    .A1(\mem.mem[99][5] ),
    .S(net3900),
    .X(_04200_));
 sg13g2_nand2_1 _12059_ (.Y(_04201_),
    .A(net3743),
    .B(_04200_));
 sg13g2_mux2_1 _12060_ (.A0(\mem.mem[96][5] ),
    .A1(\mem.mem[97][5] ),
    .S(net3902),
    .X(_04202_));
 sg13g2_a21oi_1 _12061_ (.A1(net3210),
    .A2(_04202_),
    .Y(_04203_),
    .B1(net3677));
 sg13g2_a21oi_1 _12062_ (.A1(_04201_),
    .A2(_04203_),
    .Y(_04204_),
    .B1(net3646));
 sg13g2_mux2_1 _12063_ (.A0(\mem.mem[106][5] ),
    .A1(\mem.mem[107][5] ),
    .S(net3917),
    .X(_04205_));
 sg13g2_nand2_1 _12064_ (.Y(_04206_),
    .A(net3748),
    .B(_04205_));
 sg13g2_mux2_1 _12065_ (.A0(\mem.mem[104][5] ),
    .A1(\mem.mem[105][5] ),
    .S(net3918),
    .X(_04207_));
 sg13g2_a21oi_1 _12066_ (.A1(net3215),
    .A2(_04207_),
    .Y(_04208_),
    .B1(net3679));
 sg13g2_nand2b_1 _12067_ (.Y(_04209_),
    .B(net3902),
    .A_N(\mem.mem[109][5] ));
 sg13g2_o21ai_1 _12068_ (.B1(_04209_),
    .Y(_04210_),
    .A1(net3902),
    .A2(\mem.mem[108][5] ));
 sg13g2_mux2_1 _12069_ (.A0(\mem.mem[110][5] ),
    .A1(\mem.mem[111][5] ),
    .S(net3901),
    .X(_04211_));
 sg13g2_a21oi_1 _12070_ (.A1(net3743),
    .A2(_04211_),
    .Y(_04212_),
    .B1(net3154));
 sg13g2_o21ai_1 _12071_ (.B1(_04212_),
    .Y(_04213_),
    .A1(net3744),
    .A2(_04210_));
 sg13g2_a21oi_2 _12072_ (.B1(net3113),
    .Y(_04214_),
    .A2(_04208_),
    .A1(_04206_));
 sg13g2_a22oi_1 _12073_ (.Y(_04215_),
    .B1(_04213_),
    .B2(_04214_),
    .A2(_04204_),
    .A1(_04199_));
 sg13g2_mux4_1 _12074_ (.S0(net3825),
    .A0(\mem.mem[112][5] ),
    .A1(\mem.mem[113][5] ),
    .A2(\mem.mem[114][5] ),
    .A3(\mem.mem[115][5] ),
    .S1(net3714),
    .X(_04216_));
 sg13g2_mux2_1 _12075_ (.A0(\mem.mem[116][5] ),
    .A1(\mem.mem[117][5] ),
    .S(net3822),
    .X(_04217_));
 sg13g2_nor2b_1 _12076_ (.A(\mem.mem[119][5] ),
    .B_N(net3821),
    .Y(_04218_));
 sg13g2_o21ai_1 _12077_ (.B1(net3714),
    .Y(_04219_),
    .A1(net3821),
    .A2(\mem.mem[118][5] ));
 sg13g2_o21ai_1 _12078_ (.B1(net3667),
    .Y(_04220_),
    .A1(_04218_),
    .A2(_04219_));
 sg13g2_a21oi_1 _12079_ (.A1(net3187),
    .A2(_04217_),
    .Y(_04221_),
    .B1(_04220_));
 sg13g2_nor2_1 _12080_ (.A(net3638),
    .B(_04221_),
    .Y(_04222_));
 sg13g2_o21ai_1 _12081_ (.B1(_04222_),
    .Y(_04223_),
    .A1(net3670),
    .A2(_04216_));
 sg13g2_mux4_1 _12082_ (.S0(net3845),
    .A0(\mem.mem[120][5] ),
    .A1(\mem.mem[121][5] ),
    .A2(\mem.mem[122][5] ),
    .A3(\mem.mem[123][5] ),
    .S1(net3721),
    .X(_04224_));
 sg13g2_nand2b_1 _12083_ (.Y(_04225_),
    .B(net3139),
    .A_N(_04224_));
 sg13g2_mux2_1 _12084_ (.A0(\mem.mem[124][5] ),
    .A1(\mem.mem[125][5] ),
    .S(net3844),
    .X(_04226_));
 sg13g2_nor2b_1 _12085_ (.A(\mem.mem[127][5] ),
    .B_N(net3844),
    .Y(_04227_));
 sg13g2_o21ai_1 _12086_ (.B1(net3721),
    .Y(_04228_),
    .A1(net3844),
    .A2(\mem.mem[126][5] ));
 sg13g2_o21ai_1 _12087_ (.B1(net3671),
    .Y(_04229_),
    .A1(_04227_),
    .A2(_04228_));
 sg13g2_a21oi_1 _12088_ (.A1(net3192),
    .A2(_04226_),
    .Y(_04230_),
    .B1(_04229_));
 sg13g2_nor2_1 _12089_ (.A(net3109),
    .B(_04230_),
    .Y(_04231_));
 sg13g2_a21oi_1 _12090_ (.A1(_04225_),
    .A2(_04231_),
    .Y(_04232_),
    .B1(net3096));
 sg13g2_a221oi_1 _12091_ (.B2(_04232_),
    .C1(net3091),
    .B1(_04223_),
    .A1(net3096),
    .Y(_04233_),
    .A2(_04215_));
 sg13g2_o21ai_1 _12092_ (.B1(net3612),
    .Y(_04234_),
    .A1(_04194_),
    .A2(_04233_));
 sg13g2_a21oi_2 _12093_ (.B1(net3614),
    .Y(_04235_),
    .A2(_04167_),
    .A1(_04139_));
 sg13g2_nor2_1 _12094_ (.A(net3611),
    .B(_04235_),
    .Y(_04236_));
 sg13g2_a21oi_2 _12095_ (.B1(_02258_),
    .Y(_04237_),
    .A2(_04236_),
    .A1(_04234_));
 sg13g2_a22oi_1 _12096_ (.Y(_04238_),
    .B1(_04099_),
    .B2(_04237_),
    .A2(_02536_),
    .A1(net6));
 sg13g2_o21ai_1 _12097_ (.B1(net4004),
    .Y(_04239_),
    .A1(net5197),
    .A2(net3055));
 sg13g2_a21oi_1 _12098_ (.A1(net3055),
    .A2(_04238_),
    .Y(_00600_),
    .B1(_04239_));
 sg13g2_mux4_1 _12099_ (.S0(net3878),
    .A0(\mem.mem[160][6] ),
    .A1(\mem.mem[161][6] ),
    .A2(\mem.mem[162][6] ),
    .A3(\mem.mem[163][6] ),
    .S1(net3734),
    .X(_04240_));
 sg13g2_mux2_1 _12100_ (.A0(\mem.mem[166][6] ),
    .A1(\mem.mem[167][6] ),
    .S(net3876),
    .X(_04241_));
 sg13g2_nand2b_1 _12101_ (.Y(_04242_),
    .B(net3876),
    .A_N(\mem.mem[165][6] ));
 sg13g2_o21ai_1 _12102_ (.B1(_04242_),
    .Y(_04243_),
    .A1(net3876),
    .A2(\mem.mem[164][6] ));
 sg13g2_o21ai_1 _12103_ (.B1(net3676),
    .Y(_04244_),
    .A1(net3735),
    .A2(_04243_));
 sg13g2_a21oi_1 _12104_ (.A1(net3735),
    .A2(_04241_),
    .Y(_04245_),
    .B1(_04244_));
 sg13g2_nor2_1 _12105_ (.A(net3645),
    .B(_04245_),
    .Y(_04246_));
 sg13g2_o21ai_1 _12106_ (.B1(_04246_),
    .Y(_04247_),
    .A1(net3675),
    .A2(_04240_));
 sg13g2_mux2_1 _12107_ (.A0(\mem.mem[172][6] ),
    .A1(\mem.mem[173][6] ),
    .S(net3837),
    .X(_04248_));
 sg13g2_nor2b_1 _12108_ (.A(\mem.mem[175][6] ),
    .B_N(net3833),
    .Y(_04249_));
 sg13g2_o21ai_1 _12109_ (.B1(net3718),
    .Y(_04250_),
    .A1(net3837),
    .A2(\mem.mem[174][6] ));
 sg13g2_o21ai_1 _12110_ (.B1(net3669),
    .Y(_04251_),
    .A1(_04249_),
    .A2(_04250_));
 sg13g2_a21oi_1 _12111_ (.A1(net3191),
    .A2(_04248_),
    .Y(_04252_),
    .B1(_04251_));
 sg13g2_mux4_1 _12112_ (.S0(net3851),
    .A0(\mem.mem[168][6] ),
    .A1(\mem.mem[169][6] ),
    .A2(\mem.mem[170][6] ),
    .A3(\mem.mem[171][6] ),
    .S1(net3725),
    .X(_04253_));
 sg13g2_nor2_1 _12113_ (.A(net3108),
    .B(_04252_),
    .Y(_04254_));
 sg13g2_o21ai_1 _12114_ (.B1(_04254_),
    .Y(_04255_),
    .A1(net3671),
    .A2(_04253_));
 sg13g2_nand3_1 _12115_ (.B(_04247_),
    .C(_04255_),
    .A(net3097),
    .Y(_04256_));
 sg13g2_mux4_1 _12116_ (.S0(net3853),
    .A0(\mem.mem[176][6] ),
    .A1(\mem.mem[177][6] ),
    .A2(\mem.mem[178][6] ),
    .A3(\mem.mem[179][6] ),
    .S1(net3726),
    .X(_04257_));
 sg13g2_mux2_1 _12117_ (.A0(\mem.mem[182][6] ),
    .A1(\mem.mem[183][6] ),
    .S(net3900),
    .X(_04258_));
 sg13g2_nand2_1 _12118_ (.Y(_04259_),
    .A(net3728),
    .B(_04258_));
 sg13g2_mux2_1 _12119_ (.A0(\mem.mem[180][6] ),
    .A1(\mem.mem[181][6] ),
    .S(net3861),
    .X(_04260_));
 sg13g2_a21oi_1 _12120_ (.A1(net3210),
    .A2(_04260_),
    .Y(_04261_),
    .B1(net3143));
 sg13g2_a21oi_1 _12121_ (.A1(_04259_),
    .A2(_04261_),
    .Y(_04262_),
    .B1(net3646));
 sg13g2_o21ai_1 _12122_ (.B1(_04262_),
    .Y(_04263_),
    .A1(net3678),
    .A2(_04257_));
 sg13g2_mux4_1 _12123_ (.S0(net3848),
    .A0(\mem.mem[184][6] ),
    .A1(\mem.mem[185][6] ),
    .A2(\mem.mem[186][6] ),
    .A3(\mem.mem[187][6] ),
    .S1(net3723),
    .X(_04264_));
 sg13g2_nor2_1 _12124_ (.A(net3671),
    .B(_04264_),
    .Y(_04265_));
 sg13g2_mux2_1 _12125_ (.A0(\mem.mem[188][6] ),
    .A1(\mem.mem[189][6] ),
    .S(net3846),
    .X(_04266_));
 sg13g2_nor2b_1 _12126_ (.A(\mem.mem[191][6] ),
    .B_N(net3846),
    .Y(_04267_));
 sg13g2_o21ai_1 _12127_ (.B1(net3723),
    .Y(_04268_),
    .A1(net3846),
    .A2(\mem.mem[190][6] ));
 sg13g2_o21ai_1 _12128_ (.B1(net3671),
    .Y(_04269_),
    .A1(_04267_),
    .A2(_04268_));
 sg13g2_a21oi_1 _12129_ (.A1(net3197),
    .A2(_04266_),
    .Y(_04270_),
    .B1(_04269_));
 sg13g2_or3_2 _12130_ (.A(net3109),
    .B(_04265_),
    .C(_04270_),
    .X(_04271_));
 sg13g2_nand3_1 _12131_ (.B(_04263_),
    .C(_04271_),
    .A(net3625),
    .Y(_04272_));
 sg13g2_nand3_1 _12132_ (.B(_04256_),
    .C(_04272_),
    .A(net3616),
    .Y(_04273_));
 sg13g2_mux4_1 _12133_ (.S0(net3919),
    .A0(\mem.mem[144][6] ),
    .A1(\mem.mem[145][6] ),
    .A2(\mem.mem[146][6] ),
    .A3(\mem.mem[147][6] ),
    .S1(net3749),
    .X(_04274_));
 sg13g2_nor2_1 _12134_ (.A(net3686),
    .B(_04274_),
    .Y(_04275_));
 sg13g2_mux2_1 _12135_ (.A0(\mem.mem[148][6] ),
    .A1(\mem.mem[149][6] ),
    .S(net3968),
    .X(_04276_));
 sg13g2_nor2b_1 _12136_ (.A(\mem.mem[151][6] ),
    .B_N(net3968),
    .Y(_04277_));
 sg13g2_o21ai_1 _12137_ (.B1(net3763),
    .Y(_04278_),
    .A1(net3968),
    .A2(\mem.mem[150][6] ));
 sg13g2_o21ai_1 _12138_ (.B1(net3686),
    .Y(_04279_),
    .A1(_04277_),
    .A2(_04278_));
 sg13g2_a21oi_2 _12139_ (.B1(_04279_),
    .Y(_04280_),
    .A2(_04276_),
    .A1(net3230));
 sg13g2_nor3_2 _12140_ (.A(net3651),
    .B(_04275_),
    .C(_04280_),
    .Y(_04281_));
 sg13g2_mux4_1 _12141_ (.S0(net3982),
    .A0(\mem.mem[152][6] ),
    .A1(\mem.mem[153][6] ),
    .A2(\mem.mem[154][6] ),
    .A3(\mem.mem[155][6] ),
    .S1(net3768),
    .X(_04282_));
 sg13g2_nor2_2 _12142_ (.A(net3688),
    .B(_04282_),
    .Y(_04283_));
 sg13g2_mux4_1 _12143_ (.S0(net3921),
    .A0(\mem.mem[156][6] ),
    .A1(\mem.mem[157][6] ),
    .A2(\mem.mem[158][6] ),
    .A3(\mem.mem[159][6] ),
    .S1(net3749),
    .X(_04284_));
 sg13g2_o21ai_1 _12144_ (.B1(net3651),
    .Y(_04285_),
    .A1(net3158),
    .A2(_04284_));
 sg13g2_o21ai_1 _12145_ (.B1(net3629),
    .Y(_04286_),
    .A1(_04283_),
    .A2(_04285_));
 sg13g2_mux4_1 _12146_ (.S0(net3932),
    .A0(\mem.mem[132][6] ),
    .A1(\mem.mem[133][6] ),
    .A2(\mem.mem[134][6] ),
    .A3(\mem.mem[135][6] ),
    .S1(net3753),
    .X(_04287_));
 sg13g2_nor2_1 _12147_ (.A(net3152),
    .B(_04287_),
    .Y(_04288_));
 sg13g2_mux4_1 _12148_ (.S0(net3886),
    .A0(\mem.mem[128][6] ),
    .A1(\mem.mem[129][6] ),
    .A2(\mem.mem[130][6] ),
    .A3(\mem.mem[131][6] ),
    .S1(net3740),
    .X(_04289_));
 sg13g2_o21ai_1 _12149_ (.B1(net3111),
    .Y(_04290_),
    .A1(net3676),
    .A2(_04289_));
 sg13g2_mux2_1 _12150_ (.A0(\mem.mem[140][6] ),
    .A1(\mem.mem[141][6] ),
    .S(net3914),
    .X(_04291_));
 sg13g2_nand2_1 _12151_ (.Y(_04292_),
    .A(net3214),
    .B(_04291_));
 sg13g2_mux2_1 _12152_ (.A0(\mem.mem[142][6] ),
    .A1(\mem.mem[143][6] ),
    .S(net3914),
    .X(_04293_));
 sg13g2_a21oi_1 _12153_ (.A1(net3747),
    .A2(_04293_),
    .Y(_04294_),
    .B1(net3157));
 sg13g2_mux4_1 _12154_ (.S0(net3898),
    .A0(\mem.mem[136][6] ),
    .A1(\mem.mem[137][6] ),
    .A2(\mem.mem[138][6] ),
    .A3(\mem.mem[139][6] ),
    .S1(net3742),
    .X(_04295_));
 sg13g2_o21ai_1 _12155_ (.B1(net3647),
    .Y(_04296_),
    .A1(net3679),
    .A2(_04295_));
 sg13g2_a21oi_1 _12156_ (.A1(_04292_),
    .A2(_04294_),
    .Y(_04297_),
    .B1(_04296_));
 sg13g2_o21ai_1 _12157_ (.B1(net3098),
    .Y(_04298_),
    .A1(_04288_),
    .A2(_04290_));
 sg13g2_nor2_1 _12158_ (.A(_04297_),
    .B(_04298_),
    .Y(_04299_));
 sg13g2_nor2_1 _12159_ (.A(net3618),
    .B(_04299_),
    .Y(_04300_));
 sg13g2_o21ai_1 _12160_ (.B1(_04300_),
    .Y(_04301_),
    .A1(_04281_),
    .A2(_04286_));
 sg13g2_mux2_1 _12161_ (.A0(\mem.mem[204][6] ),
    .A1(\mem.mem[205][6] ),
    .S(net3779),
    .X(_04302_));
 sg13g2_nand2_1 _12162_ (.Y(_04303_),
    .A(net3181),
    .B(_04302_));
 sg13g2_mux2_1 _12163_ (.A0(\mem.mem[206][6] ),
    .A1(\mem.mem[207][6] ),
    .S(net3780),
    .X(_04304_));
 sg13g2_a21oi_1 _12164_ (.A1(net3695),
    .A2(_04304_),
    .Y(_04305_),
    .B1(net3124));
 sg13g2_mux4_1 _12165_ (.S0(net3779),
    .A0(\mem.mem[200][6] ),
    .A1(\mem.mem[201][6] ),
    .A2(\mem.mem[202][6] ),
    .A3(\mem.mem[203][6] ),
    .S1(net3695),
    .X(_04306_));
 sg13g2_o21ai_1 _12166_ (.B1(net3632),
    .Y(_04307_),
    .A1(net3658),
    .A2(_04306_));
 sg13g2_a21oi_1 _12167_ (.A1(_04303_),
    .A2(_04305_),
    .Y(_04308_),
    .B1(_04307_));
 sg13g2_mux4_1 _12168_ (.S0(net3774),
    .A0(\mem.mem[192][6] ),
    .A1(\mem.mem[193][6] ),
    .A2(\mem.mem[194][6] ),
    .A3(\mem.mem[195][6] ),
    .S1(net3692),
    .X(_04309_));
 sg13g2_nor2_1 _12169_ (.A(net3657),
    .B(_04309_),
    .Y(_04310_));
 sg13g2_mux2_1 _12170_ (.A0(\mem.mem[198][6] ),
    .A1(\mem.mem[199][6] ),
    .S(net3775),
    .X(_04311_));
 sg13g2_nand2b_1 _12171_ (.Y(_04312_),
    .B(net3774),
    .A_N(\mem.mem[197][6] ));
 sg13g2_o21ai_1 _12172_ (.B1(_04312_),
    .Y(_04313_),
    .A1(net3774),
    .A2(\mem.mem[196][6] ));
 sg13g2_o21ai_1 _12173_ (.B1(net3657),
    .Y(_04314_),
    .A1(net3692),
    .A2(_04313_));
 sg13g2_a21oi_1 _12174_ (.A1(net3692),
    .A2(_04311_),
    .Y(_04315_),
    .B1(_04314_));
 sg13g2_nor3_2 _12175_ (.A(net3632),
    .B(_04310_),
    .C(_04315_),
    .Y(_04316_));
 sg13g2_nor3_2 _12176_ (.A(net3620),
    .B(_04308_),
    .C(_04316_),
    .Y(_04317_));
 sg13g2_mux4_1 _12177_ (.S0(net3820),
    .A0(\mem.mem[220][6] ),
    .A1(\mem.mem[221][6] ),
    .A2(\mem.mem[222][6] ),
    .A3(\mem.mem[223][6] ),
    .S1(net3712),
    .X(_04318_));
 sg13g2_nor2_1 _12178_ (.A(net3133),
    .B(_04318_),
    .Y(_04319_));
 sg13g2_mux4_1 _12179_ (.S0(net3788),
    .A0(\mem.mem[216][6] ),
    .A1(\mem.mem[217][6] ),
    .A2(\mem.mem[218][6] ),
    .A3(\mem.mem[219][6] ),
    .S1(net3696),
    .X(_04320_));
 sg13g2_o21ai_1 _12180_ (.B1(net3638),
    .Y(_04321_),
    .A1(net3667),
    .A2(_04320_));
 sg13g2_nand2b_1 _12181_ (.Y(_04322_),
    .B(\mem.mem[210][6] ),
    .A_N(net3783));
 sg13g2_a21oi_1 _12182_ (.A1(net3783),
    .A2(\mem.mem[211][6] ),
    .Y(_04323_),
    .B1(net3178));
 sg13g2_nor2b_1 _12183_ (.A(net3783),
    .B_N(\mem.mem[208][6] ),
    .Y(_04324_));
 sg13g2_a21oi_1 _12184_ (.A1(net3783),
    .A2(\mem.mem[209][6] ),
    .Y(_04325_),
    .B1(_04324_));
 sg13g2_a221oi_1 _12185_ (.B2(net3178),
    .C1(net3659),
    .B1(_04325_),
    .A1(_04322_),
    .Y(_04326_),
    .A2(_04323_));
 sg13g2_nor2b_1 _12186_ (.A(net3791),
    .B_N(\mem.mem[212][6] ),
    .Y(_04327_));
 sg13g2_a21oi_1 _12187_ (.A1(net3791),
    .A2(\mem.mem[213][6] ),
    .Y(_04328_),
    .B1(_04327_));
 sg13g2_nand2b_1 _12188_ (.Y(_04329_),
    .B(\mem.mem[214][6] ),
    .A_N(net3790));
 sg13g2_a21oi_1 _12189_ (.A1(net3790),
    .A2(\mem.mem[215][6] ),
    .Y(_04330_),
    .B1(net3179));
 sg13g2_a221oi_1 _12190_ (.B2(_04330_),
    .C1(net3123),
    .B1(_04329_),
    .A1(net3179),
    .Y(_04331_),
    .A2(_04328_));
 sg13g2_o21ai_1 _12191_ (.B1(net3102),
    .Y(_04332_),
    .A1(_04326_),
    .A2(_04331_));
 sg13g2_o21ai_1 _12192_ (.B1(net3623),
    .Y(_04333_),
    .A1(_04319_),
    .A2(_04321_));
 sg13g2_nor2b_1 _12193_ (.A(_04333_),
    .B_N(_04332_),
    .Y(_04334_));
 sg13g2_nor3_2 _12194_ (.A(net3615),
    .B(_04317_),
    .C(_04334_),
    .Y(_04335_));
 sg13g2_nand2b_1 _12195_ (.Y(_04336_),
    .B(\mem.mem[230][6] ),
    .A_N(net3868));
 sg13g2_a21oi_1 _12196_ (.A1(net3868),
    .A2(\mem.mem[231][6] ),
    .Y(_04337_),
    .B1(net3200));
 sg13g2_nor2b_1 _12197_ (.A(net3880),
    .B_N(\mem.mem[228][6] ),
    .Y(_04338_));
 sg13g2_a21oi_1 _12198_ (.A1(net3880),
    .A2(\mem.mem[229][6] ),
    .Y(_04339_),
    .B1(_04338_));
 sg13g2_a221oi_1 _12199_ (.B2(net3200),
    .C1(net3148),
    .B1(_04339_),
    .A1(_04336_),
    .Y(_04340_),
    .A2(_04337_));
 sg13g2_nor2b_1 _12200_ (.A(net3865),
    .B_N(\mem.mem[224][6] ),
    .Y(_04341_));
 sg13g2_a21oi_1 _12201_ (.A1(net3865),
    .A2(\mem.mem[225][6] ),
    .Y(_04342_),
    .B1(_04341_));
 sg13g2_nand2b_1 _12202_ (.Y(_04343_),
    .B(\mem.mem[226][6] ),
    .A_N(net3865));
 sg13g2_a21oi_1 _12203_ (.A1(net3865),
    .A2(\mem.mem[227][6] ),
    .Y(_04344_),
    .B1(net3201));
 sg13g2_a221oi_1 _12204_ (.B2(_04344_),
    .C1(net3675),
    .B1(_04343_),
    .A1(net3200),
    .Y(_04345_),
    .A2(_04342_));
 sg13g2_o21ai_1 _12205_ (.B1(net3111),
    .Y(_04346_),
    .A1(_04340_),
    .A2(_04345_));
 sg13g2_mux4_1 _12206_ (.S0(net3832),
    .A0(\mem.mem[232][6] ),
    .A1(\mem.mem[233][6] ),
    .A2(\mem.mem[234][6] ),
    .A3(\mem.mem[235][6] ),
    .S1(net3716),
    .X(_04347_));
 sg13g2_nand2b_1 _12207_ (.Y(_04348_),
    .B(\mem.mem[236][6] ),
    .A_N(net3830));
 sg13g2_a21oi_1 _12208_ (.A1(net3830),
    .A2(\mem.mem[237][6] ),
    .Y(_04349_),
    .B1(net3717));
 sg13g2_nor2b_1 _12209_ (.A(net3830),
    .B_N(\mem.mem[238][6] ),
    .Y(_04350_));
 sg13g2_a21oi_1 _12210_ (.A1(net3830),
    .A2(\mem.mem[239][6] ),
    .Y(_04351_),
    .B1(_04350_));
 sg13g2_a221oi_1 _12211_ (.B2(net3716),
    .C1(net3135),
    .B1(_04351_),
    .A1(_04348_),
    .Y(_04352_),
    .A2(_04349_));
 sg13g2_a21o_1 _12212_ (.A2(_04347_),
    .A1(net3135),
    .B1(_04352_),
    .X(_04353_));
 sg13g2_a21oi_1 _12213_ (.A1(net3638),
    .A2(_04353_),
    .Y(_04354_),
    .B1(net3623));
 sg13g2_nor2b_1 _12214_ (.A(net3828),
    .B_N(\mem.mem[246][6] ),
    .Y(_04355_));
 sg13g2_a21oi_1 _12215_ (.A1(net3827),
    .A2(\mem.mem[247][6] ),
    .Y(_04356_),
    .B1(_04355_));
 sg13g2_nand2b_1 _12216_ (.Y(_04357_),
    .B(\mem.mem[244][6] ),
    .A_N(net3827));
 sg13g2_a21oi_1 _12217_ (.A1(net3827),
    .A2(\mem.mem[245][6] ),
    .Y(_04358_),
    .B1(net3715));
 sg13g2_a221oi_1 _12218_ (.B2(_04358_),
    .C1(net3135),
    .B1(_04357_),
    .A1(net3715),
    .Y(_04359_),
    .A2(_04356_));
 sg13g2_nor2b_1 _12219_ (.A(net3827),
    .B_N(\mem.mem[240][6] ),
    .Y(_04360_));
 sg13g2_a21oi_1 _12220_ (.A1(net3827),
    .A2(\mem.mem[241][6] ),
    .Y(_04361_),
    .B1(_04360_));
 sg13g2_nand2b_1 _12221_ (.Y(_04362_),
    .B(\mem.mem[242][6] ),
    .A_N(net3827));
 sg13g2_a21oi_1 _12222_ (.A1(net3827),
    .A2(\mem.mem[243][6] ),
    .Y(_04363_),
    .B1(net3190));
 sg13g2_a221oi_1 _12223_ (.B2(_04363_),
    .C1(net3668),
    .B1(_04362_),
    .A1(net3190),
    .Y(_04364_),
    .A2(_04361_));
 sg13g2_o21ai_1 _12224_ (.B1(net3107),
    .Y(_04365_),
    .A1(_04359_),
    .A2(_04364_));
 sg13g2_mux4_1 _12225_ (.S0(net3834),
    .A0(\mem.mem[248][6] ),
    .A1(\mem.mem[249][6] ),
    .A2(\mem.mem[250][6] ),
    .A3(\mem.mem[251][6] ),
    .S1(net3715),
    .X(_04366_));
 sg13g2_inv_1 _12226_ (.Y(_04367_),
    .A(_04366_));
 sg13g2_o21ai_1 _12227_ (.B1(net3639),
    .Y(_04368_),
    .A1(net3135),
    .A2(\mem.mem[252][6] ));
 sg13g2_a21oi_1 _12228_ (.A1(net3135),
    .A2(_04367_),
    .Y(_04369_),
    .B1(_04368_));
 sg13g2_nor2_1 _12229_ (.A(net3095),
    .B(_04369_),
    .Y(_04370_));
 sg13g2_a221oi_1 _12230_ (.B2(_04370_),
    .C1(net3091),
    .B1(_04365_),
    .A1(_04346_),
    .Y(_04371_),
    .A2(_04354_));
 sg13g2_a21oi_2 _12231_ (.B1(net3613),
    .Y(_04372_),
    .A2(_04301_),
    .A1(_04273_));
 sg13g2_o21ai_1 _12232_ (.B1(net3612),
    .Y(_04373_),
    .A1(_04335_),
    .A2(_04371_));
 sg13g2_nand2_1 _12233_ (.Y(_04374_),
    .A(net3611),
    .B(_04373_));
 sg13g2_nor2_1 _12234_ (.A(_04372_),
    .B(_04374_),
    .Y(_04375_));
 sg13g2_mux2_1 _12235_ (.A0(\mem.mem[76][6] ),
    .A1(\mem.mem[77][6] ),
    .S(net3800),
    .X(_04376_));
 sg13g2_nand2_1 _12236_ (.Y(_04377_),
    .A(net3182),
    .B(_04376_));
 sg13g2_mux2_1 _12237_ (.A0(\mem.mem[78][6] ),
    .A1(\mem.mem[79][6] ),
    .S(net3800),
    .X(_04378_));
 sg13g2_a21oi_1 _12238_ (.A1(net3704),
    .A2(_04378_),
    .Y(_04379_),
    .B1(net3128));
 sg13g2_mux4_1 _12239_ (.S0(net3797),
    .A0(\mem.mem[72][6] ),
    .A1(\mem.mem[73][6] ),
    .A2(\mem.mem[74][6] ),
    .A3(\mem.mem[75][6] ),
    .S1(net3702),
    .X(_04380_));
 sg13g2_o21ai_1 _12240_ (.B1(net3634),
    .Y(_04381_),
    .A1(net3661),
    .A2(_04380_));
 sg13g2_a21oi_2 _12241_ (.B1(_04381_),
    .Y(_04382_),
    .A2(_04379_),
    .A1(_04377_));
 sg13g2_mux2_1 _12242_ (.A0(\mem.mem[70][6] ),
    .A1(\mem.mem[71][6] ),
    .S(net3812),
    .X(_04383_));
 sg13g2_mux2_1 _12243_ (.A0(\mem.mem[68][6] ),
    .A1(\mem.mem[69][6] ),
    .S(net3812),
    .X(_04384_));
 sg13g2_nand2_1 _12244_ (.Y(_04385_),
    .A(net3185),
    .B(_04384_));
 sg13g2_a21oi_1 _12245_ (.A1(net3709),
    .A2(_04383_),
    .Y(_04386_),
    .B1(net3132));
 sg13g2_mux2_1 _12246_ (.A0(\mem.mem[66][6] ),
    .A1(\mem.mem[67][6] ),
    .S(net3812),
    .X(_04387_));
 sg13g2_nand2_1 _12247_ (.Y(_04388_),
    .A(net3709),
    .B(_04387_));
 sg13g2_mux2_1 _12248_ (.A0(\mem.mem[64][6] ),
    .A1(\mem.mem[65][6] ),
    .S(net3812),
    .X(_04389_));
 sg13g2_a21oi_1 _12249_ (.A1(net3185),
    .A2(_04389_),
    .Y(_04390_),
    .B1(net3664));
 sg13g2_a221oi_1 _12250_ (.B2(_04390_),
    .C1(net3635),
    .B1(_04388_),
    .A1(_04385_),
    .Y(_04391_),
    .A2(_04386_));
 sg13g2_nor3_2 _12251_ (.A(net3621),
    .B(_04382_),
    .C(_04391_),
    .Y(_04392_));
 sg13g2_mux4_1 _12252_ (.S0(net3800),
    .A0(\mem.mem[80][6] ),
    .A1(\mem.mem[81][6] ),
    .A2(\mem.mem[82][6] ),
    .A3(\mem.mem[83][6] ),
    .S1(net3704),
    .X(_04393_));
 sg13g2_nor2_1 _12253_ (.A(net3662),
    .B(_04393_),
    .Y(_04394_));
 sg13g2_mux2_1 _12254_ (.A0(\mem.mem[84][6] ),
    .A1(\mem.mem[85][6] ),
    .S(net3813),
    .X(_04395_));
 sg13g2_nor2b_1 _12255_ (.A(\mem.mem[87][6] ),
    .B_N(net3813),
    .Y(_04396_));
 sg13g2_o21ai_1 _12256_ (.B1(net3708),
    .Y(_04397_),
    .A1(net3813),
    .A2(\mem.mem[86][6] ));
 sg13g2_o21ai_1 _12257_ (.B1(net3664),
    .Y(_04398_),
    .A1(_04396_),
    .A2(_04397_));
 sg13g2_a21oi_1 _12258_ (.A1(net3184),
    .A2(_04395_),
    .Y(_04399_),
    .B1(_04398_));
 sg13g2_nor3_1 _12259_ (.A(net3635),
    .B(_04394_),
    .C(_04399_),
    .Y(_04400_));
 sg13g2_mux2_1 _12260_ (.A0(\mem.mem[92][6] ),
    .A1(\mem.mem[93][6] ),
    .S(net3805),
    .X(_04401_));
 sg13g2_mux2_1 _12261_ (.A0(\mem.mem[94][6] ),
    .A1(\mem.mem[95][6] ),
    .S(net3804),
    .X(_04402_));
 sg13g2_nand2_1 _12262_ (.Y(_04403_),
    .A(net3707),
    .B(_04402_));
 sg13g2_a21oi_1 _12263_ (.A1(net3183),
    .A2(_04401_),
    .Y(_04404_),
    .B1(net3129));
 sg13g2_mux2_1 _12264_ (.A0(\mem.mem[90][6] ),
    .A1(\mem.mem[91][6] ),
    .S(net3804),
    .X(_04405_));
 sg13g2_nand2_1 _12265_ (.Y(_04406_),
    .A(net3707),
    .B(_04405_));
 sg13g2_mux2_1 _12266_ (.A0(\mem.mem[88][6] ),
    .A1(\mem.mem[89][6] ),
    .S(net3805),
    .X(_04407_));
 sg13g2_a21oi_1 _12267_ (.A1(net3183),
    .A2(_04407_),
    .Y(_04408_),
    .B1(net3663));
 sg13g2_a221oi_1 _12268_ (.B2(_04408_),
    .C1(net3103),
    .B1(_04406_),
    .A1(_04403_),
    .Y(_04409_),
    .A2(_04404_));
 sg13g2_nand2b_1 _12269_ (.Y(_04410_),
    .B(net3621),
    .A_N(_04409_));
 sg13g2_o21ai_1 _12270_ (.B1(net3091),
    .Y(_04411_),
    .A1(_04400_),
    .A2(_04410_));
 sg13g2_nand2b_1 _12271_ (.Y(_04412_),
    .B(\mem.mem[102][6] ),
    .A_N(net3909));
 sg13g2_a21oi_1 _12272_ (.A1(net3909),
    .A2(\mem.mem[103][6] ),
    .Y(_04413_),
    .B1(net3213));
 sg13g2_nor2b_1 _12273_ (.A(net3914),
    .B_N(\mem.mem[100][6] ),
    .Y(_04414_));
 sg13g2_a21oi_1 _12274_ (.A1(net3913),
    .A2(\mem.mem[101][6] ),
    .Y(_04415_),
    .B1(_04414_));
 sg13g2_a221oi_1 _12275_ (.B2(net3213),
    .C1(net3156),
    .B1(_04415_),
    .A1(_04412_),
    .Y(_04416_),
    .A2(_04413_));
 sg13g2_nor2b_1 _12276_ (.A(net3899),
    .B_N(\mem.mem[96][6] ),
    .Y(_04417_));
 sg13g2_a21oi_1 _12277_ (.A1(net3903),
    .A2(\mem.mem[97][6] ),
    .Y(_04418_),
    .B1(_04417_));
 sg13g2_nand2b_1 _12278_ (.Y(_04419_),
    .B(\mem.mem[98][6] ),
    .A_N(net3903));
 sg13g2_a21oi_1 _12279_ (.A1(net3903),
    .A2(\mem.mem[99][6] ),
    .Y(_04420_),
    .B1(net3211));
 sg13g2_a221oi_1 _12280_ (.B2(_04420_),
    .C1(net3678),
    .B1(_04419_),
    .A1(net3211),
    .Y(_04421_),
    .A2(_04418_));
 sg13g2_nor3_1 _12281_ (.A(net3646),
    .B(_04416_),
    .C(_04421_),
    .Y(_04422_));
 sg13g2_mux4_1 _12282_ (.S0(net3905),
    .A0(\mem.mem[104][6] ),
    .A1(\mem.mem[105][6] ),
    .A2(\mem.mem[106][6] ),
    .A3(\mem.mem[107][6] ),
    .S1(net3744),
    .X(_04423_));
 sg13g2_mux2_1 _12283_ (.A0(\mem.mem[108][6] ),
    .A1(\mem.mem[109][6] ),
    .S(net3901),
    .X(_04424_));
 sg13g2_o21ai_1 _12284_ (.B1(net3743),
    .Y(_04425_),
    .A1(net3901),
    .A2(_02166_));
 sg13g2_a21oi_1 _12285_ (.A1(net3901),
    .A2(\mem.mem[111][6] ),
    .Y(_04426_),
    .B1(_04425_));
 sg13g2_o21ai_1 _12286_ (.B1(net3678),
    .Y(_04427_),
    .A1(net3743),
    .A2(_04424_));
 sg13g2_o21ai_1 _12287_ (.B1(net3646),
    .Y(_04428_),
    .A1(_04426_),
    .A2(_04427_));
 sg13g2_a21oi_2 _12288_ (.B1(_04428_),
    .Y(_04429_),
    .A2(_04423_),
    .A1(net3154));
 sg13g2_o21ai_1 _12289_ (.B1(net3097),
    .Y(_04430_),
    .A1(_04422_),
    .A2(_04429_));
 sg13g2_nor2b_1 _12290_ (.A(net3822),
    .B_N(\mem.mem[116][6] ),
    .Y(_04431_));
 sg13g2_a21oi_1 _12291_ (.A1(net3822),
    .A2(\mem.mem[117][6] ),
    .Y(_04432_),
    .B1(_04431_));
 sg13g2_nand2b_1 _12292_ (.Y(_04433_),
    .B(\mem.mem[118][6] ),
    .A_N(net3821));
 sg13g2_a21oi_1 _12293_ (.A1(net3826),
    .A2(\mem.mem[119][6] ),
    .Y(_04434_),
    .B1(net3187));
 sg13g2_a221oi_1 _12294_ (.B2(_04434_),
    .C1(net3134),
    .B1(_04433_),
    .A1(net3187),
    .Y(_04435_),
    .A2(_04432_));
 sg13g2_nor2b_1 _12295_ (.A(net3825),
    .B_N(\mem.mem[112][6] ),
    .Y(_04436_));
 sg13g2_a21oi_1 _12296_ (.A1(net3825),
    .A2(\mem.mem[113][6] ),
    .Y(_04437_),
    .B1(_04436_));
 sg13g2_nand2b_1 _12297_ (.Y(_04438_),
    .B(\mem.mem[114][6] ),
    .A_N(net3826));
 sg13g2_a21oi_1 _12298_ (.A1(net3825),
    .A2(\mem.mem[115][6] ),
    .Y(_04439_),
    .B1(net3188));
 sg13g2_a221oi_1 _12299_ (.B2(_04439_),
    .C1(net3667),
    .B1(_04438_),
    .A1(net3188),
    .Y(_04440_),
    .A2(_04437_));
 sg13g2_nor3_2 _12300_ (.A(net3638),
    .B(_04435_),
    .C(_04440_),
    .Y(_04441_));
 sg13g2_mux4_1 _12301_ (.S0(net3841),
    .A0(\mem.mem[120][6] ),
    .A1(\mem.mem[121][6] ),
    .A2(\mem.mem[122][6] ),
    .A3(\mem.mem[123][6] ),
    .S1(net3721),
    .X(_04442_));
 sg13g2_a21oi_1 _12302_ (.A1(net3842),
    .A2(\mem.mem[127][6] ),
    .Y(_04443_),
    .B1(net3192));
 sg13g2_o21ai_1 _12303_ (.B1(_04443_),
    .Y(_04444_),
    .A1(net3842),
    .A2(_02167_));
 sg13g2_nand2b_1 _12304_ (.Y(_04445_),
    .B(\mem.mem[124][6] ),
    .A_N(net3843));
 sg13g2_a21oi_1 _12305_ (.A1(net3843),
    .A2(\mem.mem[125][6] ),
    .Y(_04446_),
    .B1(net3722));
 sg13g2_a21oi_1 _12306_ (.A1(_04445_),
    .A2(_04446_),
    .Y(_04447_),
    .B1(net3139));
 sg13g2_a221oi_1 _12307_ (.B2(_04447_),
    .C1(net3109),
    .B1(_04444_),
    .A1(net3139),
    .Y(_04448_),
    .A2(_04442_));
 sg13g2_o21ai_1 _12308_ (.B1(net3622),
    .Y(_04449_),
    .A1(_04441_),
    .A2(_04448_));
 sg13g2_and2_1 _12309_ (.A(net3615),
    .B(_04449_),
    .X(_04450_));
 sg13g2_nand2b_1 _12310_ (.Y(_04451_),
    .B(\mem.mem[38][6] ),
    .A_N(net3946));
 sg13g2_a21oi_1 _12311_ (.A1(net3946),
    .A2(\mem.mem[39][6] ),
    .Y(_04452_),
    .B1(net3224));
 sg13g2_nor2b_1 _12312_ (.A(net3949),
    .B_N(\mem.mem[36][6] ),
    .Y(_04453_));
 sg13g2_a21oi_1 _12313_ (.A1(net3949),
    .A2(\mem.mem[37][6] ),
    .Y(_04454_),
    .B1(_04453_));
 sg13g2_a221oi_1 _12314_ (.B2(net3224),
    .C1(net3163),
    .B1(_04454_),
    .A1(_04451_),
    .Y(_04455_),
    .A2(_04452_));
 sg13g2_nor2b_1 _12315_ (.A(net3935),
    .B_N(\mem.mem[32][6] ),
    .Y(_04456_));
 sg13g2_a21oi_1 _12316_ (.A1(net3935),
    .A2(\mem.mem[33][6] ),
    .Y(_04457_),
    .B1(_04456_));
 sg13g2_nand2b_1 _12317_ (.Y(_04458_),
    .B(\mem.mem[34][6] ),
    .A_N(net3935));
 sg13g2_a21oi_1 _12318_ (.A1(net3935),
    .A2(\mem.mem[35][6] ),
    .Y(_04459_),
    .B1(net3221));
 sg13g2_a221oi_1 _12319_ (.B2(_04459_),
    .C1(net3685),
    .B1(_04458_),
    .A1(net3220),
    .Y(_04460_),
    .A2(_04457_));
 sg13g2_nor3_2 _12320_ (.A(net3649),
    .B(_04455_),
    .C(_04460_),
    .Y(_04461_));
 sg13g2_mux4_1 _12321_ (.S0(net3979),
    .A0(\mem.mem[40][6] ),
    .A1(\mem.mem[41][6] ),
    .A2(\mem.mem[42][6] ),
    .A3(\mem.mem[43][6] ),
    .S1(net3765),
    .X(_04462_));
 sg13g2_mux2_1 _12322_ (.A0(\mem.mem[44][6] ),
    .A1(\mem.mem[45][6] ),
    .S(net3960),
    .X(_04463_));
 sg13g2_o21ai_1 _12323_ (.B1(net3761),
    .Y(_04464_),
    .A1(net3959),
    .A2(_02164_));
 sg13g2_a21oi_1 _12324_ (.A1(net3959),
    .A2(\mem.mem[47][6] ),
    .Y(_04465_),
    .B1(_04464_));
 sg13g2_o21ai_1 _12325_ (.B1(net3689),
    .Y(_04466_),
    .A1(net3761),
    .A2(_04463_));
 sg13g2_o21ai_1 _12326_ (.B1(net3653),
    .Y(_04467_),
    .A1(_04465_),
    .A2(_04466_));
 sg13g2_a21oi_1 _12327_ (.A1(net3166),
    .A2(_04462_),
    .Y(_04468_),
    .B1(_04467_));
 sg13g2_o21ai_1 _12328_ (.B1(net3098),
    .Y(_04469_),
    .A1(_04461_),
    .A2(_04468_));
 sg13g2_nor2b_1 _12329_ (.A(net3961),
    .B_N(\mem.mem[52][6] ),
    .Y(_04470_));
 sg13g2_a21oi_1 _12330_ (.A1(net3963),
    .A2(\mem.mem[53][6] ),
    .Y(_04471_),
    .B1(_04470_));
 sg13g2_nand2b_1 _12331_ (.Y(_04472_),
    .B(\mem.mem[54][6] ),
    .A_N(net3963));
 sg13g2_a21oi_1 _12332_ (.A1(net3961),
    .A2(\mem.mem[55][6] ),
    .Y(_04473_),
    .B1(net3229));
 sg13g2_a221oi_1 _12333_ (.B2(_04473_),
    .C1(net3166),
    .B1(_04472_),
    .A1(net3229),
    .Y(_04474_),
    .A2(_04471_));
 sg13g2_nor2b_1 _12334_ (.A(net3957),
    .B_N(\mem.mem[48][6] ),
    .Y(_04475_));
 sg13g2_a21oi_1 _12335_ (.A1(net3958),
    .A2(\mem.mem[49][6] ),
    .Y(_04476_),
    .B1(_04475_));
 sg13g2_nand2b_1 _12336_ (.Y(_04477_),
    .B(\mem.mem[50][6] ),
    .A_N(net3957));
 sg13g2_a21oi_1 _12337_ (.A1(net3957),
    .A2(\mem.mem[51][6] ),
    .Y(_04478_),
    .B1(net3228));
 sg13g2_a221oi_1 _12338_ (.B2(_04478_),
    .C1(net3686),
    .B1(_04477_),
    .A1(net3228),
    .Y(_04479_),
    .A2(_04476_));
 sg13g2_nor3_1 _12339_ (.A(net3652),
    .B(_04474_),
    .C(_04479_),
    .Y(_04480_));
 sg13g2_mux4_1 _12340_ (.S0(net3977),
    .A0(\mem.mem[56][6] ),
    .A1(\mem.mem[57][6] ),
    .A2(\mem.mem[58][6] ),
    .A3(\mem.mem[59][6] ),
    .S1(net3766),
    .X(_04481_));
 sg13g2_a21oi_1 _12341_ (.A1(net3984),
    .A2(\mem.mem[63][6] ),
    .Y(_04482_),
    .B1(net3235));
 sg13g2_o21ai_1 _12342_ (.B1(_04482_),
    .Y(_04483_),
    .A1(net3984),
    .A2(_02165_));
 sg13g2_nand2b_1 _12343_ (.Y(_04484_),
    .B(\mem.mem[60][6] ),
    .A_N(net3983));
 sg13g2_a21oi_1 _12344_ (.A1(net3983),
    .A2(\mem.mem[61][6] ),
    .Y(_04485_),
    .B1(net3768));
 sg13g2_a21oi_1 _12345_ (.A1(_04484_),
    .A2(_04485_),
    .Y(_04486_),
    .B1(net3172));
 sg13g2_a221oi_1 _12346_ (.B2(_04486_),
    .C1(net3118),
    .B1(_04483_),
    .A1(net3170),
    .Y(_04487_),
    .A2(_04481_));
 sg13g2_o21ai_1 _12347_ (.B1(net3630),
    .Y(_04488_),
    .A1(_04480_),
    .A2(_04487_));
 sg13g2_nand3_1 _12348_ (.B(_04469_),
    .C(_04488_),
    .A(net3618),
    .Y(_04489_));
 sg13g2_mux2_1 _12349_ (.A0(\mem.mem[12][6] ),
    .A1(\mem.mem[13][6] ),
    .S(net3889),
    .X(_04490_));
 sg13g2_nand2_1 _12350_ (.Y(_04491_),
    .A(net3220),
    .B(_04490_));
 sg13g2_mux2_1 _12351_ (.A0(\mem.mem[14][6] ),
    .A1(\mem.mem[15][6] ),
    .S(net3888),
    .X(_04492_));
 sg13g2_a21oi_1 _12352_ (.A1(net3739),
    .A2(_04492_),
    .Y(_04493_),
    .B1(net3152));
 sg13g2_mux4_1 _12353_ (.S0(net3887),
    .A0(\mem.mem[8][6] ),
    .A1(\mem.mem[9][6] ),
    .A2(\mem.mem[10][6] ),
    .A3(\mem.mem[11][6] ),
    .S1(net3740),
    .X(_04494_));
 sg13g2_o21ai_1 _12354_ (.B1(net3645),
    .Y(_04495_),
    .A1(net3676),
    .A2(_04494_));
 sg13g2_a21oi_1 _12355_ (.A1(_04491_),
    .A2(_04493_),
    .Y(_04496_),
    .B1(_04495_));
 sg13g2_mux2_1 _12356_ (.A0(\mem.mem[6][6] ),
    .A1(\mem.mem[7][6] ),
    .S(net3884),
    .X(_04497_));
 sg13g2_mux2_1 _12357_ (.A0(\mem.mem[4][6] ),
    .A1(\mem.mem[5][6] ),
    .S(net3884),
    .X(_04498_));
 sg13g2_nand2_1 _12358_ (.Y(_04499_),
    .A(net3206),
    .B(_04498_));
 sg13g2_a21oi_1 _12359_ (.A1(net3737),
    .A2(_04497_),
    .Y(_04500_),
    .B1(net3151));
 sg13g2_mux2_1 _12360_ (.A0(\mem.mem[2][6] ),
    .A1(\mem.mem[3][6] ),
    .S(net3925),
    .X(_04501_));
 sg13g2_nand2_1 _12361_ (.Y(_04502_),
    .A(net3737),
    .B(_04501_));
 sg13g2_mux2_1 _12362_ (.A0(\mem.mem[0][6] ),
    .A1(\mem.mem[1][6] ),
    .S(net3884),
    .X(_04503_));
 sg13g2_a21oi_1 _12363_ (.A1(net3219),
    .A2(_04503_),
    .Y(_04504_),
    .B1(net3682));
 sg13g2_a221oi_1 _12364_ (.B2(_04504_),
    .C1(net3650),
    .B1(_04502_),
    .A1(_04499_),
    .Y(_04505_),
    .A2(_04500_));
 sg13g2_nor3_1 _12365_ (.A(net3628),
    .B(_04496_),
    .C(_04505_),
    .Y(_04506_));
 sg13g2_mux2_1 _12366_ (.A0(\mem.mem[22][6] ),
    .A1(\mem.mem[23][6] ),
    .S(net3939),
    .X(_04507_));
 sg13g2_nand2_1 _12367_ (.Y(_04508_),
    .A(net3755),
    .B(_04507_));
 sg13g2_mux2_1 _12368_ (.A0(\mem.mem[20][6] ),
    .A1(\mem.mem[21][6] ),
    .S(net3939),
    .X(_04509_));
 sg13g2_a21oi_1 _12369_ (.A1(net3222),
    .A2(_04509_),
    .Y(_04510_),
    .B1(net3161));
 sg13g2_mux2_1 _12370_ (.A0(\mem.mem[18][6] ),
    .A1(\mem.mem[19][6] ),
    .S(net3927),
    .X(_04511_));
 sg13g2_nand2_1 _12371_ (.Y(_04512_),
    .A(net3751),
    .B(_04511_));
 sg13g2_mux2_1 _12372_ (.A0(\mem.mem[16][6] ),
    .A1(\mem.mem[17][6] ),
    .S(net3939),
    .X(_04513_));
 sg13g2_a21oi_1 _12373_ (.A1(net3222),
    .A2(_04513_),
    .Y(_04514_),
    .B1(net3683));
 sg13g2_a221oi_1 _12374_ (.B2(_04514_),
    .C1(net3648),
    .B1(_04512_),
    .A1(_04508_),
    .Y(_04515_),
    .A2(_04510_));
 sg13g2_mux4_1 _12375_ (.S0(net3949),
    .A0(\mem.mem[24][6] ),
    .A1(\mem.mem[25][6] ),
    .A2(\mem.mem[26][6] ),
    .A3(\mem.mem[27][6] ),
    .S1(net3757),
    .X(_04516_));
 sg13g2_nor2_1 _12376_ (.A(net3684),
    .B(_04516_),
    .Y(_04517_));
 sg13g2_nor2b_1 _12377_ (.A(\mem.mem[29][6] ),
    .B_N(net3933),
    .Y(_04518_));
 sg13g2_nor2_1 _12378_ (.A(net3933),
    .B(\mem.mem[28][6] ),
    .Y(_04519_));
 sg13g2_nor3_1 _12379_ (.A(net3754),
    .B(_04518_),
    .C(_04519_),
    .Y(_04520_));
 sg13g2_nor2b_1 _12380_ (.A(\mem.mem[31][6] ),
    .B_N(net3933),
    .Y(_04521_));
 sg13g2_o21ai_1 _12381_ (.B1(net3753),
    .Y(_04522_),
    .A1(net3933),
    .A2(\mem.mem[30][6] ));
 sg13g2_o21ai_1 _12382_ (.B1(net3685),
    .Y(_04523_),
    .A1(_04521_),
    .A2(_04522_));
 sg13g2_o21ai_1 _12383_ (.B1(net3649),
    .Y(_04524_),
    .A1(_04520_),
    .A2(_04523_));
 sg13g2_o21ai_1 _12384_ (.B1(net3626),
    .Y(_04525_),
    .A1(_04517_),
    .A2(_04524_));
 sg13g2_o21ai_1 _12385_ (.B1(net3092),
    .Y(_04526_),
    .A1(_04515_),
    .A2(_04525_));
 sg13g2_o21ai_1 _12386_ (.B1(net3089),
    .Y(_04527_),
    .A1(_04506_),
    .A2(_04526_));
 sg13g2_nand2b_2 _12387_ (.Y(_04528_),
    .B(_04489_),
    .A_N(_04527_));
 sg13g2_a21oi_1 _12388_ (.A1(_04430_),
    .A2(_04450_),
    .Y(_04529_),
    .B1(net3089));
 sg13g2_o21ai_1 _12389_ (.B1(_04529_),
    .Y(_04530_),
    .A1(_04392_),
    .A2(_04411_));
 sg13g2_a21oi_1 _12390_ (.A1(_04528_),
    .A2(_04530_),
    .Y(_04531_),
    .B1(net3611));
 sg13g2_nor3_2 _12391_ (.A(_02258_),
    .B(_04375_),
    .C(_04531_),
    .Y(_04532_));
 sg13g2_a21o_2 _12392_ (.A2(_02536_),
    .A1(net7),
    .B1(_04532_),
    .X(_04533_));
 sg13g2_o21ai_1 _12393_ (.B1(net4005),
    .Y(_04534_),
    .A1(_02535_),
    .A2(_04533_));
 sg13g2_a21oi_1 _12394_ (.A1(_02141_),
    .A2(_02535_),
    .Y(_00601_),
    .B1(_04534_));
 sg13g2_nor2b_1 _12395_ (.A(net3808),
    .B_N(\mem.mem[68][7] ),
    .Y(_04535_));
 sg13g2_a21oi_1 _12396_ (.A1(net3808),
    .A2(\mem.mem[69][7] ),
    .Y(_04536_),
    .B1(_04535_));
 sg13g2_nand2b_1 _12397_ (.Y(_04537_),
    .B(\mem.mem[70][7] ),
    .A_N(net3808));
 sg13g2_a21oi_1 _12398_ (.A1(net3808),
    .A2(\mem.mem[71][7] ),
    .Y(_04538_),
    .B1(net3182));
 sg13g2_a221oi_1 _12399_ (.B2(_04538_),
    .C1(net3128),
    .B1(_04537_),
    .A1(net3182),
    .Y(_04539_),
    .A2(_04536_));
 sg13g2_nor2b_1 _12400_ (.A(net3792),
    .B_N(\mem.mem[64][7] ),
    .Y(_04540_));
 sg13g2_a21oi_1 _12401_ (.A1(net3791),
    .A2(\mem.mem[65][7] ),
    .Y(_04541_),
    .B1(_04540_));
 sg13g2_nand2b_1 _12402_ (.Y(_04542_),
    .B(\mem.mem[66][7] ),
    .A_N(net3791));
 sg13g2_a21oi_1 _12403_ (.A1(net3791),
    .A2(\mem.mem[67][7] ),
    .Y(_04543_),
    .B1(net3179));
 sg13g2_a221oi_1 _12404_ (.B2(_04543_),
    .C1(net3660),
    .B1(_04542_),
    .A1(net3179),
    .Y(_04544_),
    .A2(_04541_));
 sg13g2_nor3_1 _12405_ (.A(net3634),
    .B(_04539_),
    .C(_04544_),
    .Y(_04545_));
 sg13g2_mux4_1 _12406_ (.S0(net3778),
    .A0(\mem.mem[72][7] ),
    .A1(\mem.mem[73][7] ),
    .A2(\mem.mem[74][7] ),
    .A3(\mem.mem[75][7] ),
    .S1(net3694),
    .X(_04546_));
 sg13g2_a21oi_1 _12407_ (.A1(net3799),
    .A2(\mem.mem[79][7] ),
    .Y(_04547_),
    .B1(net3182));
 sg13g2_o21ai_1 _12408_ (.B1(_04547_),
    .Y(_04548_),
    .A1(net3799),
    .A2(_02172_));
 sg13g2_nand2b_1 _12409_ (.Y(_04549_),
    .B(\mem.mem[76][7] ),
    .A_N(net3797));
 sg13g2_a21oi_1 _12410_ (.A1(net3797),
    .A2(\mem.mem[77][7] ),
    .Y(_04550_),
    .B1(net3702));
 sg13g2_a21oi_1 _12411_ (.A1(_04549_),
    .A2(_04550_),
    .Y(_04551_),
    .B1(net3128));
 sg13g2_a221oi_1 _12412_ (.B2(_04551_),
    .C1(net3103),
    .B1(_04548_),
    .A1(net3128),
    .Y(_04552_),
    .A2(_04546_));
 sg13g2_o21ai_1 _12413_ (.B1(net3096),
    .Y(_04553_),
    .A1(_04545_),
    .A2(_04552_));
 sg13g2_nand2b_1 _12414_ (.Y(_04554_),
    .B(\mem.mem[84][7] ),
    .A_N(net3809));
 sg13g2_a21oi_1 _12415_ (.A1(net3809),
    .A2(\mem.mem[85][7] ),
    .Y(_04555_),
    .B1(net3708));
 sg13g2_nor2b_1 _12416_ (.A(net3809),
    .B_N(\mem.mem[86][7] ),
    .Y(_04556_));
 sg13g2_a21oi_1 _12417_ (.A1(net3809),
    .A2(\mem.mem[87][7] ),
    .Y(_04557_),
    .B1(_04556_));
 sg13g2_a221oi_1 _12418_ (.B2(net3704),
    .C1(net3128),
    .B1(_04557_),
    .A1(_04554_),
    .Y(_04558_),
    .A2(_04555_));
 sg13g2_nand2b_1 _12419_ (.Y(_04559_),
    .B(\mem.mem[80][7] ),
    .A_N(net3798));
 sg13g2_a21oi_1 _12420_ (.A1(net3798),
    .A2(\mem.mem[81][7] ),
    .Y(_04560_),
    .B1(net3703));
 sg13g2_nor2b_1 _12421_ (.A(net3798),
    .B_N(\mem.mem[82][7] ),
    .Y(_04561_));
 sg13g2_a21oi_1 _12422_ (.A1(net3799),
    .A2(\mem.mem[83][7] ),
    .Y(_04562_),
    .B1(_04561_));
 sg13g2_a221oi_1 _12423_ (.B2(net3703),
    .C1(net3662),
    .B1(_04562_),
    .A1(_04559_),
    .Y(_04563_),
    .A2(_04560_));
 sg13g2_nor3_1 _12424_ (.A(net3634),
    .B(_04558_),
    .C(_04563_),
    .Y(_04564_));
 sg13g2_mux4_1 _12425_ (.S0(net3803),
    .A0(\mem.mem[88][7] ),
    .A1(\mem.mem[89][7] ),
    .A2(\mem.mem[90][7] ),
    .A3(\mem.mem[91][7] ),
    .S1(net3705),
    .X(_04565_));
 sg13g2_o21ai_1 _12426_ (.B1(net3706),
    .Y(_04566_),
    .A1(net3802),
    .A2(_02173_));
 sg13g2_a21oi_1 _12427_ (.A1(net3802),
    .A2(\mem.mem[95][7] ),
    .Y(_04567_),
    .B1(_04566_));
 sg13g2_mux2_1 _12428_ (.A0(\mem.mem[92][7] ),
    .A1(\mem.mem[93][7] ),
    .S(net3802),
    .X(_04568_));
 sg13g2_o21ai_1 _12429_ (.B1(net3663),
    .Y(_04569_),
    .A1(net3706),
    .A2(_04568_));
 sg13g2_o21ai_1 _12430_ (.B1(net3635),
    .Y(_04570_),
    .A1(_04567_),
    .A2(_04569_));
 sg13g2_a21oi_2 _12431_ (.B1(_04570_),
    .Y(_04571_),
    .A2(_04565_),
    .A1(net3129));
 sg13g2_o21ai_1 _12432_ (.B1(net3621),
    .Y(_04572_),
    .A1(_04564_),
    .A2(_04571_));
 sg13g2_nand3_1 _12433_ (.B(_04553_),
    .C(_04572_),
    .A(net3090),
    .Y(_04573_));
 sg13g2_nor2b_1 _12434_ (.A(net3919),
    .B_N(\mem.mem[100][7] ),
    .Y(_04574_));
 sg13g2_a21oi_1 _12435_ (.A1(net3919),
    .A2(\mem.mem[101][7] ),
    .Y(_04575_),
    .B1(_04574_));
 sg13g2_nand2b_1 _12436_ (.Y(_04576_),
    .B(\mem.mem[102][7] ),
    .A_N(net3916));
 sg13g2_a21oi_1 _12437_ (.A1(net3916),
    .A2(\mem.mem[103][7] ),
    .Y(_04577_),
    .B1(net3216));
 sg13g2_a221oi_1 _12438_ (.B2(_04577_),
    .C1(net3158),
    .B1(_04576_),
    .A1(net3216),
    .Y(_04578_),
    .A2(_04575_));
 sg13g2_nor2b_1 _12439_ (.A(net3899),
    .B_N(\mem.mem[96][7] ),
    .Y(_04579_));
 sg13g2_a21oi_1 _12440_ (.A1(net3906),
    .A2(\mem.mem[97][7] ),
    .Y(_04580_),
    .B1(_04579_));
 sg13g2_nand2b_1 _12441_ (.Y(_04581_),
    .B(\mem.mem[98][7] ),
    .A_N(net3903));
 sg13g2_a21oi_1 _12442_ (.A1(net3903),
    .A2(\mem.mem[99][7] ),
    .Y(_04582_),
    .B1(net3211));
 sg13g2_a221oi_1 _12443_ (.B2(_04582_),
    .C1(net3677),
    .B1(_04581_),
    .A1(net3211),
    .Y(_04583_),
    .A2(_04580_));
 sg13g2_nor3_1 _12444_ (.A(net3647),
    .B(_04578_),
    .C(_04583_),
    .Y(_04584_));
 sg13g2_mux4_1 _12445_ (.S0(net3917),
    .A0(\mem.mem[104][7] ),
    .A1(\mem.mem[105][7] ),
    .A2(\mem.mem[106][7] ),
    .A3(\mem.mem[107][7] ),
    .S1(net3748),
    .X(_04585_));
 sg13g2_a21oi_1 _12446_ (.A1(net3901),
    .A2(\mem.mem[111][7] ),
    .Y(_04586_),
    .B1(net3210));
 sg13g2_o21ai_1 _12447_ (.B1(_04586_),
    .Y(_04587_),
    .A1(net3901),
    .A2(_02174_));
 sg13g2_nand2b_1 _12448_ (.Y(_04588_),
    .B(\mem.mem[108][7] ),
    .A_N(net3901));
 sg13g2_a21oi_1 _12449_ (.A1(net3901),
    .A2(\mem.mem[109][7] ),
    .Y(_04589_),
    .B1(net3743));
 sg13g2_a21oi_1 _12450_ (.A1(_04588_),
    .A2(_04589_),
    .Y(_04590_),
    .B1(net3154));
 sg13g2_a221oi_1 _12451_ (.B2(_04590_),
    .C1(net3112),
    .B1(_04587_),
    .A1(net3154),
    .Y(_04591_),
    .A2(_04585_));
 sg13g2_o21ai_1 _12452_ (.B1(net3097),
    .Y(_04592_),
    .A1(_04584_),
    .A2(_04591_));
 sg13g2_nor2b_1 _12453_ (.A(net3820),
    .B_N(\mem.mem[116][7] ),
    .Y(_04593_));
 sg13g2_a21oi_1 _12454_ (.A1(net3820),
    .A2(\mem.mem[117][7] ),
    .Y(_04594_),
    .B1(_04593_));
 sg13g2_nand2b_1 _12455_ (.Y(_04595_),
    .B(\mem.mem[118][7] ),
    .A_N(net3824));
 sg13g2_a21oi_1 _12456_ (.A1(net3824),
    .A2(\mem.mem[119][7] ),
    .Y(_04596_),
    .B1(net3187));
 sg13g2_a221oi_1 _12457_ (.B2(_04596_),
    .C1(net3134),
    .B1(_04595_),
    .A1(net3189),
    .Y(_04597_),
    .A2(_04594_));
 sg13g2_nor2b_1 _12458_ (.A(net3824),
    .B_N(\mem.mem[112][7] ),
    .Y(_04598_));
 sg13g2_a21oi_1 _12459_ (.A1(net3824),
    .A2(\mem.mem[113][7] ),
    .Y(_04599_),
    .B1(_04598_));
 sg13g2_nand2b_1 _12460_ (.Y(_04600_),
    .B(\mem.mem[114][7] ),
    .A_N(net3824));
 sg13g2_a21oi_1 _12461_ (.A1(net3824),
    .A2(\mem.mem[115][7] ),
    .Y(_04601_),
    .B1(net3188));
 sg13g2_a221oi_1 _12462_ (.B2(_04601_),
    .C1(net3667),
    .B1(_04600_),
    .A1(net3188),
    .Y(_04602_),
    .A2(_04599_));
 sg13g2_nor3_2 _12463_ (.A(net3638),
    .B(_04597_),
    .C(_04602_),
    .Y(_04603_));
 sg13g2_mux4_1 _12464_ (.S0(net3842),
    .A0(\mem.mem[120][7] ),
    .A1(\mem.mem[121][7] ),
    .A2(\mem.mem[122][7] ),
    .A3(\mem.mem[123][7] ),
    .S1(net3722),
    .X(_04604_));
 sg13g2_a21oi_1 _12465_ (.A1(net3842),
    .A2(\mem.mem[127][7] ),
    .Y(_04605_),
    .B1(net3192));
 sg13g2_o21ai_1 _12466_ (.B1(_04605_),
    .Y(_04606_),
    .A1(net3842),
    .A2(_02175_));
 sg13g2_nand2b_1 _12467_ (.Y(_04607_),
    .B(\mem.mem[124][7] ),
    .A_N(net3843));
 sg13g2_a21oi_1 _12468_ (.A1(net3842),
    .A2(\mem.mem[125][7] ),
    .Y(_04608_),
    .B1(net3722));
 sg13g2_a21oi_1 _12469_ (.A1(_04607_),
    .A2(_04608_),
    .Y(_04609_),
    .B1(net3140));
 sg13g2_a221oi_1 _12470_ (.B2(_04609_),
    .C1(net3106),
    .B1(_04606_),
    .A1(net3139),
    .Y(_04610_),
    .A2(_04604_));
 sg13g2_o21ai_1 _12471_ (.B1(net3623),
    .Y(_04611_),
    .A1(_04603_),
    .A2(_04610_));
 sg13g2_nand3_1 _12472_ (.B(_04592_),
    .C(_04611_),
    .A(net3619),
    .Y(_04612_));
 sg13g2_a21oi_1 _12473_ (.A1(_04573_),
    .A2(_04612_),
    .Y(_04613_),
    .B1(net3089));
 sg13g2_nor2b_1 _12474_ (.A(net3948),
    .B_N(\mem.mem[36][7] ),
    .Y(_04614_));
 sg13g2_a21oi_1 _12475_ (.A1(net3948),
    .A2(\mem.mem[37][7] ),
    .Y(_04615_),
    .B1(_04614_));
 sg13g2_nand2b_1 _12476_ (.Y(_04616_),
    .B(\mem.mem[38][7] ),
    .A_N(net3948));
 sg13g2_a21oi_1 _12477_ (.A1(net3948),
    .A2(\mem.mem[39][7] ),
    .Y(_04617_),
    .B1(net3224));
 sg13g2_a221oi_1 _12478_ (.B2(_04617_),
    .C1(net3163),
    .B1(_04616_),
    .A1(net3224),
    .Y(_04618_),
    .A2(_04615_));
 sg13g2_nor2b_1 _12479_ (.A(net3934),
    .B_N(\mem.mem[32][7] ),
    .Y(_04619_));
 sg13g2_a21oi_1 _12480_ (.A1(net3934),
    .A2(\mem.mem[33][7] ),
    .Y(_04620_),
    .B1(_04619_));
 sg13g2_nand2b_1 _12481_ (.Y(_04621_),
    .B(\mem.mem[34][7] ),
    .A_N(net3933));
 sg13g2_a21oi_1 _12482_ (.A1(net3933),
    .A2(\mem.mem[35][7] ),
    .Y(_04622_),
    .B1(net3220));
 sg13g2_a221oi_1 _12483_ (.B2(_04622_),
    .C1(net3682),
    .B1(_04621_),
    .A1(net3220),
    .Y(_04623_),
    .A2(_04620_));
 sg13g2_nor3_1 _12484_ (.A(net3648),
    .B(_04618_),
    .C(_04623_),
    .Y(_04624_));
 sg13g2_mux4_1 _12485_ (.S0(net3951),
    .A0(\mem.mem[40][7] ),
    .A1(\mem.mem[41][7] ),
    .A2(\mem.mem[42][7] ),
    .A3(\mem.mem[43][7] ),
    .S1(net3758),
    .X(_04625_));
 sg13g2_a21oi_1 _12486_ (.A1(net3945),
    .A2(\mem.mem[47][7] ),
    .Y(_04626_),
    .B1(net3226));
 sg13g2_o21ai_1 _12487_ (.B1(_04626_),
    .Y(_04627_),
    .A1(net3945),
    .A2(_02170_));
 sg13g2_nand2b_1 _12488_ (.Y(_04628_),
    .B(\mem.mem[44][7] ),
    .A_N(net3946));
 sg13g2_a21oi_1 _12489_ (.A1(net3945),
    .A2(\mem.mem[45][7] ),
    .Y(_04629_),
    .B1(net3757));
 sg13g2_a21oi_1 _12490_ (.A1(_04628_),
    .A2(_04629_),
    .Y(_04630_),
    .B1(net3162));
 sg13g2_a221oi_1 _12491_ (.B2(_04630_),
    .C1(net3116),
    .B1(_04627_),
    .A1(net3162),
    .Y(_04631_),
    .A2(_04625_));
 sg13g2_o21ai_1 _12492_ (.B1(net3098),
    .Y(_04632_),
    .A1(_04624_),
    .A2(_04631_));
 sg13g2_nand2b_1 _12493_ (.Y(_04633_),
    .B(\mem.mem[52][7] ),
    .A_N(net3962));
 sg13g2_a21oi_1 _12494_ (.A1(net3959),
    .A2(\mem.mem[53][7] ),
    .Y(_04634_),
    .B1(net3761));
 sg13g2_nor2b_1 _12495_ (.A(net3959),
    .B_N(\mem.mem[54][7] ),
    .Y(_04635_));
 sg13g2_a21oi_1 _12496_ (.A1(net3959),
    .A2(\mem.mem[55][7] ),
    .Y(_04636_),
    .B1(_04635_));
 sg13g2_a221oi_1 _12497_ (.B2(net3761),
    .C1(net3166),
    .B1(_04636_),
    .A1(_04633_),
    .Y(_04637_),
    .A2(_04634_));
 sg13g2_nand2b_1 _12498_ (.Y(_04638_),
    .B(\mem.mem[48][7] ),
    .A_N(net3955));
 sg13g2_a21oi_1 _12499_ (.A1(net3960),
    .A2(\mem.mem[49][7] ),
    .Y(_04639_),
    .B1(net3761));
 sg13g2_nor2b_1 _12500_ (.A(net3956),
    .B_N(\mem.mem[50][7] ),
    .Y(_04640_));
 sg13g2_a21oi_1 _12501_ (.A1(net3955),
    .A2(\mem.mem[51][7] ),
    .Y(_04641_),
    .B1(_04640_));
 sg13g2_a221oi_1 _12502_ (.B2(net3760),
    .C1(net3686),
    .B1(_04641_),
    .A1(_04638_),
    .Y(_04642_),
    .A2(_04639_));
 sg13g2_nor3_1 _12503_ (.A(net3653),
    .B(_04637_),
    .C(_04642_),
    .Y(_04643_));
 sg13g2_mux4_1 _12504_ (.S0(net3980),
    .A0(\mem.mem[56][7] ),
    .A1(\mem.mem[57][7] ),
    .A2(\mem.mem[58][7] ),
    .A3(\mem.mem[59][7] ),
    .S1(net3765),
    .X(_04644_));
 sg13g2_o21ai_1 _12505_ (.B1(net3767),
    .Y(_04645_),
    .A1(net3984),
    .A2(_02171_));
 sg13g2_a21oi_1 _12506_ (.A1(net3984),
    .A2(\mem.mem[63][7] ),
    .Y(_04646_),
    .B1(_04645_));
 sg13g2_mux2_1 _12507_ (.A0(\mem.mem[60][7] ),
    .A1(\mem.mem[61][7] ),
    .S(net3984),
    .X(_04647_));
 sg13g2_o21ai_1 _12508_ (.B1(net3688),
    .Y(_04648_),
    .A1(net3767),
    .A2(_04647_));
 sg13g2_o21ai_1 _12509_ (.B1(net3654),
    .Y(_04649_),
    .A1(_04646_),
    .A2(_04648_));
 sg13g2_a21oi_2 _12510_ (.B1(_04649_),
    .Y(_04650_),
    .A2(_04644_),
    .A1(net3171));
 sg13g2_o21ai_1 _12511_ (.B1(net3630),
    .Y(_04651_),
    .A1(_04643_),
    .A2(_04650_));
 sg13g2_nand3_1 _12512_ (.B(_04632_),
    .C(_04651_),
    .A(net3618),
    .Y(_04652_));
 sg13g2_nor2b_1 _12513_ (.A(net3881),
    .B_N(\mem.mem[4][7] ),
    .Y(_04653_));
 sg13g2_a21oi_1 _12514_ (.A1(net3881),
    .A2(\mem.mem[5][7] ),
    .Y(_04654_),
    .B1(_04653_));
 sg13g2_nand2b_1 _12515_ (.Y(_04655_),
    .B(\mem.mem[6][7] ),
    .A_N(net3881));
 sg13g2_a21oi_1 _12516_ (.A1(net3881),
    .A2(\mem.mem[7][7] ),
    .Y(_04656_),
    .B1(net3206));
 sg13g2_a221oi_1 _12517_ (.B2(_04656_),
    .C1(net3150),
    .B1(_04655_),
    .A1(net3206),
    .Y(_04657_),
    .A2(_04654_));
 sg13g2_nor2b_1 _12518_ (.A(net3925),
    .B_N(\mem.mem[0][7] ),
    .Y(_04658_));
 sg13g2_a21oi_1 _12519_ (.A1(net3926),
    .A2(\mem.mem[1][7] ),
    .Y(_04659_),
    .B1(_04658_));
 sg13g2_nand2b_1 _12520_ (.Y(_04660_),
    .B(\mem.mem[2][7] ),
    .A_N(net3926));
 sg13g2_a21oi_1 _12521_ (.A1(net3926),
    .A2(\mem.mem[3][7] ),
    .Y(_04661_),
    .B1(net3219));
 sg13g2_a221oi_1 _12522_ (.B2(_04661_),
    .C1(net3682),
    .B1(_04660_),
    .A1(net3219),
    .Y(_04662_),
    .A2(_04659_));
 sg13g2_nor3_1 _12523_ (.A(net3650),
    .B(_04657_),
    .C(_04662_),
    .Y(_04663_));
 sg13g2_mux4_1 _12524_ (.S0(net3888),
    .A0(\mem.mem[8][7] ),
    .A1(\mem.mem[9][7] ),
    .A2(\mem.mem[10][7] ),
    .A3(\mem.mem[11][7] ),
    .S1(net3739),
    .X(_04664_));
 sg13g2_a21oi_1 _12525_ (.A1(net3931),
    .A2(\mem.mem[15][7] ),
    .Y(_04665_),
    .B1(net3220));
 sg13g2_o21ai_1 _12526_ (.B1(_04665_),
    .Y(_04666_),
    .A1(net3931),
    .A2(_02168_));
 sg13g2_nand2b_1 _12527_ (.Y(_04667_),
    .B(\mem.mem[12][7] ),
    .A_N(net3931));
 sg13g2_a21oi_1 _12528_ (.A1(net3931),
    .A2(\mem.mem[13][7] ),
    .Y(_04668_),
    .B1(net3752));
 sg13g2_a21oi_1 _12529_ (.A1(_04667_),
    .A2(_04668_),
    .Y(_04669_),
    .B1(net3165));
 sg13g2_a221oi_1 _12530_ (.B2(_04669_),
    .C1(net3117),
    .B1(_04666_),
    .A1(net3165),
    .Y(_04670_),
    .A2(_04664_));
 sg13g2_o21ai_1 _12531_ (.B1(net3098),
    .Y(_04671_),
    .A1(_04663_),
    .A2(_04670_));
 sg13g2_mux2_1 _12532_ (.A0(\mem.mem[20][7] ),
    .A1(\mem.mem[21][7] ),
    .S(net3941),
    .X(_04672_));
 sg13g2_o21ai_1 _12533_ (.B1(net3755),
    .Y(_04673_),
    .A1(net3941),
    .A2(_02169_));
 sg13g2_a21oi_1 _12534_ (.A1(net3941),
    .A2(\mem.mem[23][7] ),
    .Y(_04674_),
    .B1(_04673_));
 sg13g2_o21ai_1 _12535_ (.B1(net3683),
    .Y(_04675_),
    .A1(net3755),
    .A2(_04672_));
 sg13g2_nor2b_1 _12536_ (.A(net3940),
    .B_N(\mem.mem[16][7] ),
    .Y(_04676_));
 sg13g2_a21oi_1 _12537_ (.A1(net3940),
    .A2(\mem.mem[17][7] ),
    .Y(_04677_),
    .B1(_04676_));
 sg13g2_nand2b_1 _12538_ (.Y(_04678_),
    .B(\mem.mem[18][7] ),
    .A_N(net3929));
 sg13g2_a21oi_1 _12539_ (.A1(net3929),
    .A2(\mem.mem[19][7] ),
    .Y(_04679_),
    .B1(net3222));
 sg13g2_a221oi_1 _12540_ (.B2(_04679_),
    .C1(net3683),
    .B1(_04678_),
    .A1(net3223),
    .Y(_04680_),
    .A2(_04677_));
 sg13g2_nor2_1 _12541_ (.A(net3648),
    .B(_04680_),
    .Y(_04681_));
 sg13g2_o21ai_1 _12542_ (.B1(_04681_),
    .Y(_04682_),
    .A1(_04674_),
    .A2(_04675_));
 sg13g2_mux4_1 _12543_ (.S0(net3949),
    .A0(\mem.mem[24][7] ),
    .A1(\mem.mem[25][7] ),
    .A2(\mem.mem[26][7] ),
    .A3(\mem.mem[27][7] ),
    .S1(net3758),
    .X(_04683_));
 sg13g2_nor2b_1 _12544_ (.A(net3942),
    .B_N(\mem.mem[30][7] ),
    .Y(_04684_));
 sg13g2_a21oi_1 _12545_ (.A1(net3941),
    .A2(\mem.mem[31][7] ),
    .Y(_04685_),
    .B1(_04684_));
 sg13g2_nand2b_1 _12546_ (.Y(_04686_),
    .B(\mem.mem[28][7] ),
    .A_N(net3941));
 sg13g2_a21oi_1 _12547_ (.A1(net3941),
    .A2(\mem.mem[29][7] ),
    .Y(_04687_),
    .B1(net3755));
 sg13g2_a221oi_1 _12548_ (.B2(_04687_),
    .C1(net3161),
    .B1(_04686_),
    .A1(net3755),
    .Y(_04688_),
    .A2(_04685_));
 sg13g2_a21o_1 _12549_ (.A2(_04683_),
    .A1(net3164),
    .B1(net3115),
    .X(_04689_));
 sg13g2_o21ai_1 _12550_ (.B1(_04682_),
    .Y(_04690_),
    .A1(_04688_),
    .A2(_04689_));
 sg13g2_a21oi_1 _12551_ (.A1(net3626),
    .A2(_04690_),
    .Y(_04691_),
    .B1(net3618));
 sg13g2_nand2_2 _12552_ (.Y(_04692_),
    .A(_04671_),
    .B(_04691_));
 sg13g2_a21oi_2 _12553_ (.B1(net3614),
    .Y(_04693_),
    .A2(_04692_),
    .A1(_04652_));
 sg13g2_nor3_1 _12554_ (.A(net3611),
    .B(_04613_),
    .C(_04693_),
    .Y(_04694_));
 sg13g2_nor2b_1 _12555_ (.A(net3776),
    .B_N(\mem.mem[196][7] ),
    .Y(_04695_));
 sg13g2_a21oi_1 _12556_ (.A1(net3776),
    .A2(\mem.mem[197][7] ),
    .Y(_04696_),
    .B1(_04695_));
 sg13g2_nand2b_1 _12557_ (.Y(_04697_),
    .B(\mem.mem[198][7] ),
    .A_N(net3776));
 sg13g2_a21oi_1 _12558_ (.A1(net3776),
    .A2(\mem.mem[199][7] ),
    .Y(_04698_),
    .B1(net3175));
 sg13g2_a221oi_1 _12559_ (.B2(_04698_),
    .C1(net3121),
    .B1(_04697_),
    .A1(net3175),
    .Y(_04699_),
    .A2(_04696_));
 sg13g2_nor2b_1 _12560_ (.A(net3772),
    .B_N(\mem.mem[192][7] ),
    .Y(_04700_));
 sg13g2_a21oi_1 _12561_ (.A1(net3772),
    .A2(\mem.mem[193][7] ),
    .Y(_04701_),
    .B1(_04700_));
 sg13g2_nand2b_1 _12562_ (.Y(_04702_),
    .B(\mem.mem[194][7] ),
    .A_N(net3772));
 sg13g2_a21oi_1 _12563_ (.A1(net3772),
    .A2(\mem.mem[195][7] ),
    .Y(_04703_),
    .B1(net3176));
 sg13g2_a221oi_1 _12564_ (.B2(_04703_),
    .C1(net3657),
    .B1(_04702_),
    .A1(net3175),
    .Y(_04704_),
    .A2(_04701_));
 sg13g2_nor3_1 _12565_ (.A(net3632),
    .B(_04699_),
    .C(_04704_),
    .Y(_04705_));
 sg13g2_mux4_1 _12566_ (.S0(net3777),
    .A0(\mem.mem[200][7] ),
    .A1(\mem.mem[201][7] ),
    .A2(\mem.mem[202][7] ),
    .A3(\mem.mem[203][7] ),
    .S1(net3693),
    .X(_04706_));
 sg13g2_a21oi_1 _12567_ (.A1(net3777),
    .A2(\mem.mem[207][7] ),
    .Y(_04707_),
    .B1(net3177));
 sg13g2_o21ai_1 _12568_ (.B1(_04707_),
    .Y(_04708_),
    .A1(net3777),
    .A2(_02179_));
 sg13g2_nand2b_1 _12569_ (.Y(_04709_),
    .B(\mem.mem[204][7] ),
    .A_N(net3778));
 sg13g2_a21oi_1 _12570_ (.A1(net3778),
    .A2(\mem.mem[205][7] ),
    .Y(_04710_),
    .B1(net3693));
 sg13g2_a21oi_1 _12571_ (.A1(_04709_),
    .A2(_04710_),
    .Y(_04711_),
    .B1(net3123));
 sg13g2_a221oi_1 _12572_ (.B2(_04711_),
    .C1(net3101),
    .B1(_04708_),
    .A1(net3123),
    .Y(_04712_),
    .A2(_04706_));
 sg13g2_o21ai_1 _12573_ (.B1(net3094),
    .Y(_04713_),
    .A1(_04705_),
    .A2(_04712_));
 sg13g2_nand2b_1 _12574_ (.Y(_04714_),
    .B(\mem.mem[214][7] ),
    .A_N(net3790));
 sg13g2_a21oi_1 _12575_ (.A1(net3790),
    .A2(\mem.mem[215][7] ),
    .Y(_04715_),
    .B1(net3179));
 sg13g2_nor2b_1 _12576_ (.A(net3791),
    .B_N(\mem.mem[212][7] ),
    .Y(_04716_));
 sg13g2_a21oi_1 _12577_ (.A1(net3792),
    .A2(\mem.mem[213][7] ),
    .Y(_04717_),
    .B1(_04716_));
 sg13g2_a221oi_1 _12578_ (.B2(net3179),
    .C1(net3127),
    .B1(_04717_),
    .A1(_04714_),
    .Y(_04718_),
    .A2(_04715_));
 sg13g2_nor2b_1 _12579_ (.A(net3784),
    .B_N(\mem.mem[208][7] ),
    .Y(_04719_));
 sg13g2_a21oi_1 _12580_ (.A1(net3784),
    .A2(\mem.mem[209][7] ),
    .Y(_04720_),
    .B1(_04719_));
 sg13g2_nand2b_1 _12581_ (.Y(_04721_),
    .B(\mem.mem[210][7] ),
    .A_N(net3784));
 sg13g2_a21oi_1 _12582_ (.A1(net3784),
    .A2(\mem.mem[211][7] ),
    .Y(_04722_),
    .B1(net3176));
 sg13g2_a221oi_1 _12583_ (.B2(_04722_),
    .C1(net3657),
    .B1(_04721_),
    .A1(net3178),
    .Y(_04723_),
    .A2(_04720_));
 sg13g2_nor3_1 _12584_ (.A(net3633),
    .B(_04718_),
    .C(_04723_),
    .Y(_04724_));
 sg13g2_mux4_1 _12585_ (.S0(net3788),
    .A0(\mem.mem[216][7] ),
    .A1(\mem.mem[217][7] ),
    .A2(\mem.mem[218][7] ),
    .A3(\mem.mem[219][7] ),
    .S1(net3696),
    .X(_04725_));
 sg13g2_mux2_1 _12586_ (.A0(\mem.mem[220][7] ),
    .A1(\mem.mem[221][7] ),
    .S(net3820),
    .X(_04726_));
 sg13g2_o21ai_1 _12587_ (.B1(net3700),
    .Y(_04727_),
    .A1(net3794),
    .A2(_02180_));
 sg13g2_a21oi_1 _12588_ (.A1(net3794),
    .A2(\mem.mem[223][7] ),
    .Y(_04728_),
    .B1(_04727_));
 sg13g2_o21ai_1 _12589_ (.B1(net3660),
    .Y(_04729_),
    .A1(net3698),
    .A2(_04726_));
 sg13g2_o21ai_1 _12590_ (.B1(net3633),
    .Y(_04730_),
    .A1(_04728_),
    .A2(_04729_));
 sg13g2_a21oi_1 _12591_ (.A1(net3125),
    .A2(_04725_),
    .Y(_04731_),
    .B1(_04730_));
 sg13g2_o21ai_1 _12592_ (.B1(net3620),
    .Y(_04732_),
    .A1(_04724_),
    .A2(_04731_));
 sg13g2_nand3_1 _12593_ (.B(_04713_),
    .C(_04732_),
    .A(net3090),
    .Y(_04733_));
 sg13g2_nand2b_1 _12594_ (.Y(_04734_),
    .B(\mem.mem[228][7] ),
    .A_N(net3880));
 sg13g2_a21oi_1 _12595_ (.A1(net3880),
    .A2(\mem.mem[229][7] ),
    .Y(_04735_),
    .B1(net3738));
 sg13g2_nand2_1 _12596_ (.Y(_04736_),
    .A(net3877),
    .B(\mem.mem[231][7] ));
 sg13g2_nand2b_1 _12597_ (.Y(_04737_),
    .B(\mem.mem[230][7] ),
    .A_N(net3877));
 sg13g2_nand3_1 _12598_ (.B(_04736_),
    .C(_04737_),
    .A(net3732),
    .Y(_04738_));
 sg13g2_a21oi_1 _12599_ (.A1(_04734_),
    .A2(_04735_),
    .Y(_04739_),
    .B1(net3147));
 sg13g2_mux4_1 _12600_ (.S0(net3867),
    .A0(\mem.mem[224][7] ),
    .A1(\mem.mem[225][7] ),
    .A2(\mem.mem[226][7] ),
    .A3(\mem.mem[227][7] ),
    .S1(net3732),
    .X(_04740_));
 sg13g2_a221oi_1 _12601_ (.B2(net3147),
    .C1(net3643),
    .B1(_04740_),
    .A1(_04738_),
    .Y(_04741_),
    .A2(_04739_));
 sg13g2_nor2b_1 _12602_ (.A(net3871),
    .B_N(\mem.mem[232][7] ),
    .Y(_04742_));
 sg13g2_a21oi_1 _12603_ (.A1(net3866),
    .A2(\mem.mem[233][7] ),
    .Y(_04743_),
    .B1(_04742_));
 sg13g2_nand2b_1 _12604_ (.Y(_04744_),
    .B(\mem.mem[234][7] ),
    .A_N(net3871));
 sg13g2_a21oi_1 _12605_ (.A1(net3866),
    .A2(\mem.mem[235][7] ),
    .Y(_04745_),
    .B1(net3201));
 sg13g2_a221oi_1 _12606_ (.B2(_04745_),
    .C1(net3674),
    .B1(_04744_),
    .A1(net3201),
    .Y(_04746_),
    .A2(_04743_));
 sg13g2_nor2b_1 _12607_ (.A(net3872),
    .B_N(\mem.mem[238][7] ),
    .Y(_04747_));
 sg13g2_a21oi_1 _12608_ (.A1(net3872),
    .A2(\mem.mem[239][7] ),
    .Y(_04748_),
    .B1(_04747_));
 sg13g2_nand2b_1 _12609_ (.Y(_04749_),
    .B(\mem.mem[236][7] ),
    .A_N(net3872));
 sg13g2_a21oi_1 _12610_ (.A1(net3872),
    .A2(\mem.mem[237][7] ),
    .Y(_04750_),
    .B1(net3734));
 sg13g2_a221oi_1 _12611_ (.B2(_04750_),
    .C1(net3148),
    .B1(_04749_),
    .A1(net3733),
    .Y(_04751_),
    .A2(_04748_));
 sg13g2_nor3_1 _12612_ (.A(net3111),
    .B(_04746_),
    .C(_04751_),
    .Y(_04752_));
 sg13g2_o21ai_1 _12613_ (.B1(net3097),
    .Y(_04753_),
    .A1(_04741_),
    .A2(_04752_));
 sg13g2_mux4_1 _12614_ (.S0(net3829),
    .A0(\mem.mem[244][7] ),
    .A1(\mem.mem[245][7] ),
    .A2(\mem.mem[246][7] ),
    .A3(\mem.mem[247][7] ),
    .S1(net3715),
    .X(_04754_));
 sg13g2_nand2_1 _12615_ (.Y(_04755_),
    .A(net3668),
    .B(_04754_));
 sg13g2_mux4_1 _12616_ (.S0(net3828),
    .A0(\mem.mem[240][7] ),
    .A1(\mem.mem[241][7] ),
    .A2(\mem.mem[242][7] ),
    .A3(\mem.mem[243][7] ),
    .S1(net3715),
    .X(_04756_));
 sg13g2_a21oi_1 _12617_ (.A1(net3135),
    .A2(_04756_),
    .Y(_04757_),
    .B1(net3639));
 sg13g2_mux4_1 _12618_ (.S0(net3834),
    .A0(\mem.mem[248][7] ),
    .A1(\mem.mem[249][7] ),
    .A2(\mem.mem[250][7] ),
    .A3(\mem.mem[251][7] ),
    .S1(net3719),
    .X(_04758_));
 sg13g2_nand2_1 _12619_ (.Y(_04759_),
    .A(net3135),
    .B(_04758_));
 sg13g2_a21oi_1 _12620_ (.A1(net3668),
    .A2(\mem.mem[252][7] ),
    .Y(_04760_),
    .B1(net3107));
 sg13g2_a22oi_1 _12621_ (.Y(_04761_),
    .B1(_04759_),
    .B2(_04760_),
    .A2(_04757_),
    .A1(_04755_));
 sg13g2_nor2_1 _12622_ (.A(net3095),
    .B(_04761_),
    .Y(_04762_));
 sg13g2_nor2_1 _12623_ (.A(net3091),
    .B(_04762_),
    .Y(_04763_));
 sg13g2_nor2b_1 _12624_ (.A(net3890),
    .B_N(\mem.mem[132][7] ),
    .Y(_04764_));
 sg13g2_a21oi_1 _12625_ (.A1(net3890),
    .A2(\mem.mem[133][7] ),
    .Y(_04765_),
    .B1(_04764_));
 sg13g2_nand2b_1 _12626_ (.Y(_04766_),
    .B(\mem.mem[134][7] ),
    .A_N(net3890));
 sg13g2_a21oi_1 _12627_ (.A1(net3891),
    .A2(\mem.mem[135][7] ),
    .Y(_04767_),
    .B1(net3207));
 sg13g2_a221oi_1 _12628_ (.B2(_04767_),
    .C1(net3152),
    .B1(_04766_),
    .A1(net3207),
    .Y(_04768_),
    .A2(_04765_));
 sg13g2_nor2b_1 _12629_ (.A(net3886),
    .B_N(\mem.mem[128][7] ),
    .Y(_04769_));
 sg13g2_a21oi_1 _12630_ (.A1(net3886),
    .A2(\mem.mem[129][7] ),
    .Y(_04770_),
    .B1(_04769_));
 sg13g2_nand2b_1 _12631_ (.Y(_04771_),
    .B(\mem.mem[130][7] ),
    .A_N(net3886));
 sg13g2_a21oi_1 _12632_ (.A1(net3886),
    .A2(\mem.mem[131][7] ),
    .Y(_04772_),
    .B1(net3207));
 sg13g2_a221oi_1 _12633_ (.B2(_04772_),
    .C1(net3676),
    .B1(_04771_),
    .A1(net3207),
    .Y(_04773_),
    .A2(_04770_));
 sg13g2_nor3_2 _12634_ (.A(net3644),
    .B(_04768_),
    .C(_04773_),
    .Y(_04774_));
 sg13g2_mux4_1 _12635_ (.S0(net3896),
    .A0(\mem.mem[136][7] ),
    .A1(\mem.mem[137][7] ),
    .A2(\mem.mem[138][7] ),
    .A3(\mem.mem[139][7] ),
    .S1(net3742),
    .X(_04775_));
 sg13g2_a21oi_1 _12636_ (.A1(net3908),
    .A2(\mem.mem[143][7] ),
    .Y(_04776_),
    .B1(net3213));
 sg13g2_o21ai_1 _12637_ (.B1(_04776_),
    .Y(_04777_),
    .A1(net3907),
    .A2(_02176_));
 sg13g2_nand2b_1 _12638_ (.Y(_04778_),
    .B(\mem.mem[140][7] ),
    .A_N(net3907));
 sg13g2_a21oi_1 _12639_ (.A1(net3907),
    .A2(\mem.mem[141][7] ),
    .Y(_04779_),
    .B1(net3746));
 sg13g2_a21oi_1 _12640_ (.A1(_04778_),
    .A2(_04779_),
    .Y(_04780_),
    .B1(net3155));
 sg13g2_a221oi_1 _12641_ (.B2(_04780_),
    .C1(net3113),
    .B1(_04777_),
    .A1(net3156),
    .Y(_04781_),
    .A2(_04775_));
 sg13g2_o21ai_1 _12642_ (.B1(net3097),
    .Y(_04782_),
    .A1(_04774_),
    .A2(_04781_));
 sg13g2_nand2b_1 _12643_ (.Y(_04783_),
    .B(\mem.mem[150][7] ),
    .A_N(net3972));
 sg13g2_a21oi_1 _12644_ (.A1(net3971),
    .A2(\mem.mem[151][7] ),
    .Y(_04784_),
    .B1(net3234));
 sg13g2_nor2b_1 _12645_ (.A(net3981),
    .B_N(\mem.mem[148][7] ),
    .Y(_04785_));
 sg13g2_a21oi_1 _12646_ (.A1(net3971),
    .A2(\mem.mem[149][7] ),
    .Y(_04786_),
    .B1(_04785_));
 sg13g2_a221oi_1 _12647_ (.B2(net3234),
    .C1(net3167),
    .B1(_04786_),
    .A1(_04783_),
    .Y(_04787_),
    .A2(_04784_));
 sg13g2_nand2b_1 _12648_ (.Y(_04788_),
    .B(\mem.mem[144][7] ),
    .A_N(net3964));
 sg13g2_a21oi_1 _12649_ (.A1(net3964),
    .A2(\mem.mem[145][7] ),
    .Y(_04789_),
    .B1(net3763));
 sg13g2_nor2b_1 _12650_ (.A(net3967),
    .B_N(\mem.mem[146][7] ),
    .Y(_04790_));
 sg13g2_a21oi_1 _12651_ (.A1(net3967),
    .A2(\mem.mem[147][7] ),
    .Y(_04791_),
    .B1(_04790_));
 sg13g2_a221oi_1 _12652_ (.B2(net3762),
    .C1(net3687),
    .B1(_04791_),
    .A1(_04788_),
    .Y(_04792_),
    .A2(_04789_));
 sg13g2_nor3_1 _12653_ (.A(net3651),
    .B(_04787_),
    .C(_04792_),
    .Y(_04793_));
 sg13g2_mux4_1 _12654_ (.S0(net3987),
    .A0(\mem.mem[152][7] ),
    .A1(\mem.mem[153][7] ),
    .A2(\mem.mem[154][7] ),
    .A3(\mem.mem[155][7] ),
    .S1(net3767),
    .X(_04794_));
 sg13g2_and2_2 _12655_ (.A(net3172),
    .B(_04794_),
    .X(_04795_));
 sg13g2_nand2b_1 _12656_ (.Y(_04796_),
    .B(\mem.mem[156][7] ),
    .A_N(net3964));
 sg13g2_a21oi_1 _12657_ (.A1(net3965),
    .A2(\mem.mem[157][7] ),
    .Y(_04797_),
    .B1(net3762));
 sg13g2_nor2b_1 _12658_ (.A(net3964),
    .B_N(\mem.mem[158][7] ),
    .Y(_04798_));
 sg13g2_a21oi_1 _12659_ (.A1(net3964),
    .A2(\mem.mem[159][7] ),
    .Y(_04799_),
    .B1(_04798_));
 sg13g2_a221oi_1 _12660_ (.B2(net3762),
    .C1(net3168),
    .B1(_04799_),
    .A1(_04796_),
    .Y(_04800_),
    .A2(_04797_));
 sg13g2_nor3_1 _12661_ (.A(net3119),
    .B(_04795_),
    .C(_04800_),
    .Y(_04801_));
 sg13g2_o21ai_1 _12662_ (.B1(net3629),
    .Y(_04802_),
    .A1(_04793_),
    .A2(_04801_));
 sg13g2_nand3_1 _12663_ (.B(_04782_),
    .C(_04802_),
    .A(net3093),
    .Y(_04803_));
 sg13g2_nor2b_1 _12664_ (.A(net3875),
    .B_N(\mem.mem[164][7] ),
    .Y(_04804_));
 sg13g2_a21oi_1 _12665_ (.A1(net3876),
    .A2(\mem.mem[165][7] ),
    .Y(_04805_),
    .B1(_04804_));
 sg13g2_nand2b_1 _12666_ (.Y(_04806_),
    .B(\mem.mem[166][7] ),
    .A_N(net3876));
 sg13g2_a21oi_1 _12667_ (.A1(net3876),
    .A2(\mem.mem[167][7] ),
    .Y(_04807_),
    .B1(net3203));
 sg13g2_a221oi_1 _12668_ (.B2(_04807_),
    .C1(net3149),
    .B1(_04806_),
    .A1(net3202),
    .Y(_04808_),
    .A2(_04805_));
 sg13g2_nor2b_1 _12669_ (.A(net3873),
    .B_N(\mem.mem[160][7] ),
    .Y(_04809_));
 sg13g2_a21oi_1 _12670_ (.A1(net3873),
    .A2(\mem.mem[161][7] ),
    .Y(_04810_),
    .B1(_04809_));
 sg13g2_nand2b_1 _12671_ (.Y(_04811_),
    .B(\mem.mem[162][7] ),
    .A_N(net3873));
 sg13g2_a21oi_1 _12672_ (.A1(net3873),
    .A2(\mem.mem[163][7] ),
    .Y(_04812_),
    .B1(net3202));
 sg13g2_a221oi_1 _12673_ (.B2(_04812_),
    .C1(net3675),
    .B1(_04811_),
    .A1(net3202),
    .Y(_04813_),
    .A2(_04810_));
 sg13g2_nor3_2 _12674_ (.A(net3645),
    .B(_04808_),
    .C(_04813_),
    .Y(_04814_));
 sg13g2_mux4_1 _12675_ (.S0(net3851),
    .A0(\mem.mem[168][7] ),
    .A1(\mem.mem[169][7] ),
    .A2(\mem.mem[170][7] ),
    .A3(\mem.mem[171][7] ),
    .S1(net3726),
    .X(_04815_));
 sg13g2_a21oi_1 _12676_ (.A1(net3851),
    .A2(\mem.mem[175][7] ),
    .Y(_04816_),
    .B1(net3196));
 sg13g2_o21ai_1 _12677_ (.B1(_04816_),
    .Y(_04817_),
    .A1(net3852),
    .A2(_02177_));
 sg13g2_nand2b_1 _12678_ (.Y(_04818_),
    .B(\mem.mem[172][7] ),
    .A_N(net3837));
 sg13g2_a21oi_1 _12679_ (.A1(net3836),
    .A2(\mem.mem[173][7] ),
    .Y(_04819_),
    .B1(net3718));
 sg13g2_a21oi_1 _12680_ (.A1(_04818_),
    .A2(_04819_),
    .Y(_04820_),
    .B1(net3137));
 sg13g2_a221oi_1 _12681_ (.B2(_04820_),
    .C1(net3110),
    .B1(_04817_),
    .A1(net3144),
    .Y(_04821_),
    .A2(_04815_));
 sg13g2_o21ai_1 _12682_ (.B1(net3097),
    .Y(_04822_),
    .A1(_04814_),
    .A2(_04821_));
 sg13g2_nand2b_1 _12683_ (.Y(_04823_),
    .B(\mem.mem[182][7] ),
    .A_N(net3859));
 sg13g2_a21oi_1 _12684_ (.A1(net3858),
    .A2(\mem.mem[183][7] ),
    .Y(_04824_),
    .B1(net3195));
 sg13g2_nor2b_1 _12685_ (.A(net3861),
    .B_N(\mem.mem[180][7] ),
    .Y(_04825_));
 sg13g2_a21oi_1 _12686_ (.A1(net3861),
    .A2(\mem.mem[181][7] ),
    .Y(_04826_),
    .B1(_04825_));
 sg13g2_a221oi_1 _12687_ (.B2(net3195),
    .C1(net3142),
    .B1(_04826_),
    .A1(_04823_),
    .Y(_04827_),
    .A2(_04824_));
 sg13g2_nor2b_1 _12688_ (.A(net3858),
    .B_N(\mem.mem[176][7] ),
    .Y(_04828_));
 sg13g2_a21oi_1 _12689_ (.A1(net3858),
    .A2(\mem.mem[177][7] ),
    .Y(_04829_),
    .B1(_04828_));
 sg13g2_nand2b_1 _12690_ (.Y(_04830_),
    .B(\mem.mem[178][7] ),
    .A_N(net3859));
 sg13g2_a21oi_1 _12691_ (.A1(net3858),
    .A2(\mem.mem[179][7] ),
    .Y(_04831_),
    .B1(net3195));
 sg13g2_a221oi_1 _12692_ (.B2(_04831_),
    .C1(net3672),
    .B1(_04830_),
    .A1(net3195),
    .Y(_04832_),
    .A2(_04829_));
 sg13g2_nor3_1 _12693_ (.A(net3641),
    .B(_04827_),
    .C(_04832_),
    .Y(_04833_));
 sg13g2_mux4_1 _12694_ (.S0(net3857),
    .A0(\mem.mem[184][7] ),
    .A1(\mem.mem[185][7] ),
    .A2(\mem.mem[186][7] ),
    .A3(\mem.mem[187][7] ),
    .S1(net3728),
    .X(_04834_));
 sg13g2_mux2_1 _12695_ (.A0(\mem.mem[188][7] ),
    .A1(\mem.mem[189][7] ),
    .S(net3848),
    .X(_04835_));
 sg13g2_o21ai_1 _12696_ (.B1(net3723),
    .Y(_04836_),
    .A1(net3847),
    .A2(_02178_));
 sg13g2_a21oi_1 _12697_ (.A1(net3847),
    .A2(\mem.mem[191][7] ),
    .Y(_04837_),
    .B1(_04836_));
 sg13g2_o21ai_1 _12698_ (.B1(net3671),
    .Y(_04838_),
    .A1(net3723),
    .A2(_04835_));
 sg13g2_o21ai_1 _12699_ (.B1(net3641),
    .Y(_04839_),
    .A1(_04837_),
    .A2(_04838_));
 sg13g2_a21oi_1 _12700_ (.A1(net3141),
    .A2(_04834_),
    .Y(_04840_),
    .B1(_04839_));
 sg13g2_o21ai_1 _12701_ (.B1(net3631),
    .Y(_04841_),
    .A1(_04833_),
    .A2(_04840_));
 sg13g2_nand3_1 _12702_ (.B(_04822_),
    .C(_04841_),
    .A(net3616),
    .Y(_04842_));
 sg13g2_nand3_1 _12703_ (.B(_04803_),
    .C(_04842_),
    .A(net3089),
    .Y(_04843_));
 sg13g2_a21oi_1 _12704_ (.A1(_04753_),
    .A2(_04763_),
    .Y(_04844_),
    .B1(net3089));
 sg13g2_nand2_2 _12705_ (.Y(_04845_),
    .A(_04733_),
    .B(_04844_));
 sg13g2_a21oi_1 _12706_ (.A1(_04843_),
    .A2(_04845_),
    .Y(_04846_),
    .B1(_02149_));
 sg13g2_nor3_2 _12707_ (.A(_02258_),
    .B(_04694_),
    .C(_04846_),
    .Y(_04847_));
 sg13g2_a21o_2 _12708_ (.A2(_02536_),
    .A1(net8),
    .B1(_04847_),
    .X(_04848_));
 sg13g2_o21ai_1 _12709_ (.B1(net4003),
    .Y(_04849_),
    .A1(_02535_),
    .A2(_04848_));
 sg13g2_a21oi_1 _12710_ (.A1(_02140_),
    .A2(_02535_),
    .Y(_00602_),
    .B1(_04849_));
 sg13g2_nor2_1 _12711_ (.A(net3610),
    .B(_02409_),
    .Y(_04850_));
 sg13g2_o21ai_1 _12712_ (.B1(net4006),
    .Y(_04851_),
    .A1(net5196),
    .A2(net3052));
 sg13g2_a21oi_1 _12713_ (.A1(_02847_),
    .A2(net3052),
    .Y(_00603_),
    .B1(_04851_));
 sg13g2_o21ai_1 _12714_ (.B1(net4006),
    .Y(_04852_),
    .A1(net5199),
    .A2(net3052));
 sg13g2_a21oi_1 _12715_ (.A1(_03131_),
    .A2(net3052),
    .Y(_00604_),
    .B1(_04852_));
 sg13g2_nor2b_1 _12716_ (.A(_03426_),
    .B_N(net3054),
    .Y(_04853_));
 sg13g2_o21ai_1 _12717_ (.B1(net4004),
    .Y(_04854_),
    .A1(net5205),
    .A2(net3054));
 sg13g2_nor2_1 _12718_ (.A(_04853_),
    .B(_04854_),
    .Y(_00605_));
 sg13g2_o21ai_1 _12719_ (.B1(net4006),
    .Y(_04855_),
    .A1(net5186),
    .A2(net3052));
 sg13g2_a21oi_1 _12720_ (.A1(_03661_),
    .A2(net3052),
    .Y(_00606_),
    .B1(_04855_));
 sg13g2_o21ai_1 _12721_ (.B1(net4006),
    .Y(_04856_),
    .A1(net5184),
    .A2(net3052));
 sg13g2_a21oi_1 _12722_ (.A1(_03953_),
    .A2(net3052),
    .Y(_00607_),
    .B1(_04856_));
 sg13g2_o21ai_1 _12723_ (.B1(net4004),
    .Y(_04857_),
    .A1(net5185),
    .A2(net3053));
 sg13g2_a21oi_1 _12724_ (.A1(_04238_),
    .A2(net3053),
    .Y(_00608_),
    .B1(_04857_));
 sg13g2_nor2b_1 _12725_ (.A(_04533_),
    .B_N(net3054),
    .Y(_04858_));
 sg13g2_o21ai_1 _12726_ (.B1(net4003),
    .Y(_04859_),
    .A1(net5204),
    .A2(net3054));
 sg13g2_nor2_1 _12727_ (.A(_04858_),
    .B(_04859_),
    .Y(_00609_));
 sg13g2_nor2b_1 _12728_ (.A(_04848_),
    .B_N(net3054),
    .Y(_04860_));
 sg13g2_o21ai_1 _12729_ (.B1(net4004),
    .Y(_04861_),
    .A1(net5192),
    .A2(net3054));
 sg13g2_nor2_1 _12730_ (.A(_04860_),
    .B(_04861_),
    .Y(_00610_));
 sg13g2_o21ai_1 _12731_ (.B1(net4007),
    .Y(_04862_),
    .A1(net5200),
    .A2(net3086));
 sg13g2_a21oi_1 _12732_ (.A1(net3086),
    .A2(_02847_),
    .Y(_00611_),
    .B1(_04862_));
 sg13g2_o21ai_1 _12733_ (.B1(net4007),
    .Y(_04863_),
    .A1(net5198),
    .A2(_02410_));
 sg13g2_a21oi_1 _12734_ (.A1(_02410_),
    .A2(_03131_),
    .Y(_00612_),
    .B1(_04863_));
 sg13g2_o21ai_1 _12735_ (.B1(net4004),
    .Y(_04864_),
    .A1(_02411_),
    .A2(_03426_));
 sg13g2_a21oi_1 _12736_ (.A1(_02139_),
    .A2(_02411_),
    .Y(_00613_),
    .B1(_04864_));
 sg13g2_o21ai_1 _12737_ (.B1(net4004),
    .Y(_04865_),
    .A1(net5181),
    .A2(net3086));
 sg13g2_a21oi_1 _12738_ (.A1(net3086),
    .A2(_03661_),
    .Y(_00614_),
    .B1(_04865_));
 sg13g2_o21ai_1 _12739_ (.B1(net4007),
    .Y(_04866_),
    .A1(net5172),
    .A2(net3086));
 sg13g2_a21oi_1 _12740_ (.A1(net3086),
    .A2(_03953_),
    .Y(_00615_),
    .B1(_04866_));
 sg13g2_o21ai_1 _12741_ (.B1(net4004),
    .Y(_04867_),
    .A1(net5190),
    .A2(net3086));
 sg13g2_a21oi_1 _12742_ (.A1(net3086),
    .A2(_04238_),
    .Y(_00616_),
    .B1(_04867_));
 sg13g2_o21ai_1 _12743_ (.B1(net4005),
    .Y(_04868_),
    .A1(_02411_),
    .A2(_04533_));
 sg13g2_a21oi_1 _12744_ (.A1(_02138_),
    .A2(_02411_),
    .Y(_00617_),
    .B1(_04868_));
 sg13g2_o21ai_1 _12745_ (.B1(net4005),
    .Y(_04869_),
    .A1(_02411_),
    .A2(_04848_));
 sg13g2_a21oi_1 _12746_ (.A1(_02137_),
    .A2(_02411_),
    .Y(_00618_),
    .B1(_04869_));
 sg13g2_nor3_1 _12747_ (.A(_02437_),
    .B(_02449_),
    .C(_02458_),
    .Y(_04870_));
 sg13g2_o21ai_1 _12748_ (.B1(_04870_),
    .Y(_04871_),
    .A1(_02404_),
    .A2(_02426_));
 sg13g2_or4_1 _12749_ (.A(_02468_),
    .B(_02482_),
    .C(_02490_),
    .D(_04871_),
    .X(_04872_));
 sg13g2_nand3_1 _12750_ (.B(_02399_),
    .C(_04872_),
    .A(net9),
    .Y(_04873_));
 sg13g2_nor2_1 _12751_ (.A(_02189_),
    .B(net3053),
    .Y(_04874_));
 sg13g2_a221oi_1 _12752_ (.B2(_04874_),
    .C1(net3994),
    .B1(_04873_),
    .A1(halted),
    .Y(_00619_),
    .A2(net5211));
 sg13g2_o21ai_1 _12753_ (.B1(net4009),
    .Y(_04875_),
    .A1(net3060),
    .A2(_02416_));
 sg13g2_inv_1 _12754_ (.Y(_00620_),
    .A(_04875_));
 sg13g2_nand2_1 _12755_ (.Y(_04876_),
    .A(net4007),
    .B(_02398_));
 sg13g2_a21oi_1 _12756_ (.A1(_02136_),
    .A2(net5188),
    .Y(_00621_),
    .B1(_04876_));
 sg13g2_nor2_1 _12757_ (.A(net4001),
    .B(net10),
    .Y(_04877_));
 sg13g2_nor2_2 _12758_ (.A(_02191_),
    .B(_04877_),
    .Y(_04878_));
 sg13g2_nand2b_2 _12759_ (.Y(_04879_),
    .B(halted),
    .A_N(_04877_));
 sg13g2_nor2_2 _12760_ (.A(_02399_),
    .B(_04878_),
    .Y(_04880_));
 sg13g2_nand2_1 _12761_ (.Y(_04881_),
    .A(_02400_),
    .B(_04879_));
 sg13g2_mux2_1 _12762_ (.A0(_00010_),
    .A1(net1),
    .S(net4001),
    .X(_04882_));
 sg13g2_a22oi_1 _12763_ (.Y(_04883_),
    .B1(_04882_),
    .B2(_04878_),
    .A2(_04880_),
    .A1(net5212));
 sg13g2_a21oi_1 _12764_ (.A1(_02405_),
    .A2(net5213),
    .Y(_00622_),
    .B1(net3994));
 sg13g2_mux2_1 _12765_ (.A0(_02425_),
    .A1(_02150_),
    .S(net4001),
    .X(_04884_));
 sg13g2_a21oi_1 _12766_ (.A1(_04878_),
    .A2(_04884_),
    .Y(_04885_),
    .B1(_02399_));
 sg13g2_o21ai_1 _12767_ (.B1(_04885_),
    .Y(_04886_),
    .A1(net5216),
    .A2(_04881_));
 sg13g2_a21oi_1 _12768_ (.A1(_02427_),
    .A2(_04886_),
    .Y(_00623_),
    .B1(net3995));
 sg13g2_o21ai_1 _12769_ (.B1(_04881_),
    .Y(_04887_),
    .A1(net4000),
    .A2(_02424_));
 sg13g2_a21oi_1 _12770_ (.A1(\PC[2] ),
    .A2(_02424_),
    .Y(_04888_),
    .B1(net4000));
 sg13g2_nor2_1 _12771_ (.A(_04879_),
    .B(_04888_),
    .Y(_04889_));
 sg13g2_nand2_1 _12772_ (.Y(_04890_),
    .A(net3),
    .B(net4001));
 sg13g2_a22oi_1 _12773_ (.Y(_04891_),
    .B1(_04889_),
    .B2(_04890_),
    .A2(_04887_),
    .A1(_02133_));
 sg13g2_nand2_1 _12774_ (.Y(_04892_),
    .A(_02400_),
    .B(_04891_));
 sg13g2_a21oi_1 _12775_ (.A1(_02438_),
    .A2(_04892_),
    .Y(_00624_),
    .B1(net3994));
 sg13g2_and3_1 _12776_ (.X(_04893_),
    .A(\PC[3] ),
    .B(\PC[2] ),
    .C(_02424_));
 sg13g2_a21oi_1 _12777_ (.A1(net4),
    .A2(net4000),
    .Y(_04894_),
    .B1(_04879_));
 sg13g2_o21ai_1 _12778_ (.B1(_04894_),
    .Y(_04895_),
    .A1(net4000),
    .A2(_04893_));
 sg13g2_o21ai_1 _12779_ (.B1(_04895_),
    .Y(_04896_),
    .A1(\PC[3] ),
    .A2(_04889_));
 sg13g2_nor2_1 _12780_ (.A(_02399_),
    .B(_04896_),
    .Y(_04897_));
 sg13g2_o21ai_1 _12781_ (.B1(net4007),
    .Y(_04898_),
    .A1(_02450_),
    .A2(_04897_));
 sg13g2_inv_1 _12782_ (.Y(_00625_),
    .A(_04898_));
 sg13g2_and2_1 _12783_ (.A(\PC[4] ),
    .B(_04893_),
    .X(_04899_));
 sg13g2_xor2_1 _12784_ (.B(_04893_),
    .A(\PC[4] ),
    .X(_04900_));
 sg13g2_nor2_1 _12785_ (.A(net4000),
    .B(_04900_),
    .Y(_04901_));
 sg13g2_a21oi_1 _12786_ (.A1(_02158_),
    .A2(net4000),
    .Y(_04902_),
    .B1(_04901_));
 sg13g2_a221oi_1 _12787_ (.B2(_04878_),
    .C1(_02459_),
    .B1(_04902_),
    .A1(net5221),
    .Y(_04903_),
    .A2(_04880_));
 sg13g2_nor2_1 _12788_ (.A(net3994),
    .B(_04903_),
    .Y(_00626_));
 sg13g2_and2_1 _12789_ (.A(\PC[5] ),
    .B(_04899_),
    .X(_04904_));
 sg13g2_xor2_1 _12790_ (.B(_04899_),
    .A(\PC[5] ),
    .X(_04905_));
 sg13g2_nor2_1 _12791_ (.A(net4000),
    .B(_04905_),
    .Y(_04906_));
 sg13g2_a21oi_1 _12792_ (.A1(_02160_),
    .A2(net4000),
    .Y(_04907_),
    .B1(_04906_));
 sg13g2_a221oi_1 _12793_ (.B2(_04878_),
    .C1(_02469_),
    .B1(_04907_),
    .A1(net5223),
    .Y(_04908_),
    .A2(_04880_));
 sg13g2_nor2_1 _12794_ (.A(net3994),
    .B(_04908_),
    .Y(_00627_));
 sg13g2_nand2_1 _12795_ (.Y(_04909_),
    .A(net7),
    .B(net4001));
 sg13g2_a21o_1 _12796_ (.A2(_04904_),
    .A1(\PC[6] ),
    .B1(net4001),
    .X(_04910_));
 sg13g2_nor2_1 _12797_ (.A(\PC[6] ),
    .B(_04904_),
    .Y(_04911_));
 sg13g2_o21ai_1 _12798_ (.B1(_04909_),
    .Y(_04912_),
    .A1(_04910_),
    .A2(_04911_));
 sg13g2_a221oi_1 _12799_ (.B2(_04878_),
    .C1(_02483_),
    .B1(_04912_),
    .A1(net5217),
    .Y(_04913_),
    .A2(_04880_));
 sg13g2_nor2_1 _12800_ (.A(net3994),
    .B(_04913_),
    .Y(_00628_));
 sg13g2_nand2_1 _12801_ (.Y(_04914_),
    .A(_04881_),
    .B(_04910_));
 sg13g2_mux2_1 _12802_ (.A0(_02131_),
    .A1(net8),
    .S(net4001),
    .X(_04915_));
 sg13g2_nor2_1 _12803_ (.A(_04879_),
    .B(_04915_),
    .Y(_04916_));
 sg13g2_a22oi_1 _12804_ (.Y(_04917_),
    .B1(_04916_),
    .B2(_04910_),
    .A2(_04914_),
    .A1(_02131_));
 sg13g2_nand2_1 _12805_ (.Y(_04918_),
    .A(_02400_),
    .B(_04917_));
 sg13g2_a21oi_1 _12806_ (.A1(_02491_),
    .A2(_04918_),
    .Y(_00629_),
    .B1(net3994));
 sg13g2_a21oi_2 _12807_ (.B1(_02390_),
    .Y(_04919_),
    .A2(net3059),
    .A1(_02191_));
 sg13g2_a21o_1 _12808_ (.A2(net3059),
    .A1(_02191_),
    .B1(_02390_),
    .X(_04920_));
 sg13g2_or2_1 _12809_ (.X(_04921_),
    .B(_02847_),
    .A(\mem_A[0] ));
 sg13g2_a21oi_1 _12810_ (.A1(net5203),
    .A2(_02847_),
    .Y(_04922_),
    .B1(net3059));
 sg13g2_o21ai_1 _12811_ (.B1(_04919_),
    .Y(_04923_),
    .A1(net1),
    .A2(_02407_));
 sg13g2_a21oi_1 _12812_ (.A1(_04921_),
    .A2(_04922_),
    .Y(_04924_),
    .B1(_04923_));
 sg13g2_a21oi_1 _12813_ (.A1(net3570),
    .A2(net3047),
    .Y(_04925_),
    .B1(_04924_));
 sg13g2_nor2_1 _12814_ (.A(net3997),
    .B(_04925_),
    .Y(_00638_));
 sg13g2_nor2b_1 _12815_ (.A(_00009_),
    .B_N(_03131_),
    .Y(_04926_));
 sg13g2_xnor2_1 _12816_ (.Y(_04927_),
    .A(_00009_),
    .B(_03131_));
 sg13g2_xnor2_1 _12817_ (.Y(_04928_),
    .A(_04921_),
    .B(_04927_));
 sg13g2_nand2_1 _12818_ (.Y(_04929_),
    .A(net3060),
    .B(_04928_));
 sg13g2_a21oi_1 _12819_ (.A1(_02150_),
    .A2(_02408_),
    .Y(_04930_),
    .B1(net3048));
 sg13g2_a22oi_1 _12820_ (.Y(_04931_),
    .B1(_04929_),
    .B2(_04930_),
    .A2(net3047),
    .A1(net3530));
 sg13g2_nor2_1 _12821_ (.A(net3998),
    .B(_04931_),
    .Y(_00639_));
 sg13g2_a21oi_1 _12822_ (.A1(_04921_),
    .A2(_04927_),
    .Y(_04932_),
    .B1(_04926_));
 sg13g2_a21o_1 _12823_ (.A2(_04927_),
    .A1(_04921_),
    .B1(_04926_),
    .X(_04933_));
 sg13g2_or2_1 _12824_ (.X(_04934_),
    .B(_03426_),
    .A(_02130_));
 sg13g2_xnor2_1 _12825_ (.Y(_04935_),
    .A(_02130_),
    .B(_03426_));
 sg13g2_xnor2_1 _12826_ (.Y(_04936_),
    .A(_04932_),
    .B(_04935_));
 sg13g2_o21ai_1 _12827_ (.B1(_04919_),
    .Y(_04937_),
    .A1(net3),
    .A2(net3060));
 sg13g2_a21oi_1 _12828_ (.A1(net3060),
    .A2(_04936_),
    .Y(_04938_),
    .B1(_04937_));
 sg13g2_a21oi_1 _12829_ (.A1(net3483),
    .A2(net3048),
    .Y(_04939_),
    .B1(_04938_));
 sg13g2_nor2_1 _12830_ (.A(net3997),
    .B(_04939_),
    .Y(_00640_));
 sg13g2_nor2_1 _12831_ (.A(\mem_A[3] ),
    .B(_03661_),
    .Y(_04940_));
 sg13g2_xnor2_1 _12832_ (.Y(_04941_),
    .A(\mem_A[3] ),
    .B(_03661_));
 sg13g2_o21ai_1 _12833_ (.B1(_04934_),
    .Y(_04942_),
    .A1(_04932_),
    .A2(_04935_));
 sg13g2_a21oi_1 _12834_ (.A1(_04941_),
    .A2(_04942_),
    .Y(_04943_),
    .B1(net3059));
 sg13g2_o21ai_1 _12835_ (.B1(_04943_),
    .Y(_04944_),
    .A1(_04941_),
    .A2(_04942_));
 sg13g2_a21oi_1 _12836_ (.A1(_02156_),
    .A2(_02408_),
    .Y(_04945_),
    .B1(net3047));
 sg13g2_a22oi_1 _12837_ (.Y(_04946_),
    .B1(_04944_),
    .B2(_04945_),
    .A2(net3047),
    .A1(net3441));
 sg13g2_nor2_1 _12838_ (.A(net3997),
    .B(_04946_),
    .Y(_00641_));
 sg13g2_nor2_1 _12839_ (.A(_04935_),
    .B(_04941_),
    .Y(_04947_));
 sg13g2_nor2_1 _12840_ (.A(_04934_),
    .B(_04940_),
    .Y(_04948_));
 sg13g2_a221oi_1 _12841_ (.B2(_04947_),
    .C1(_04948_),
    .B1(_04933_),
    .A1(\mem_A[3] ),
    .Y(_04949_),
    .A2(_03661_));
 sg13g2_and2_1 _12842_ (.A(\mem_A[4] ),
    .B(_03953_),
    .X(_04950_));
 sg13g2_nand2_1 _12843_ (.Y(_04951_),
    .A(\mem_A[4] ),
    .B(_03953_));
 sg13g2_xnor2_1 _12844_ (.Y(_04952_),
    .A(\mem_A[4] ),
    .B(_03953_));
 sg13g2_xnor2_1 _12845_ (.Y(_04953_),
    .A(_04949_),
    .B(_04952_));
 sg13g2_nand2_1 _12846_ (.Y(_04954_),
    .A(net3060),
    .B(_04953_));
 sg13g2_a21oi_1 _12847_ (.A1(_02158_),
    .A2(_02408_),
    .Y(_04955_),
    .B1(net3048));
 sg13g2_a22oi_1 _12848_ (.Y(_04956_),
    .B1(_04954_),
    .B2(_04955_),
    .A2(net3048),
    .A1(net3396));
 sg13g2_nor2_1 _12849_ (.A(net3997),
    .B(_04956_),
    .Y(_00642_));
 sg13g2_and2_1 _12850_ (.A(\mem_A[5] ),
    .B(_04238_),
    .X(_04957_));
 sg13g2_or2_1 _12851_ (.X(_04958_),
    .B(_04238_),
    .A(\mem_A[5] ));
 sg13g2_xnor2_1 _12852_ (.Y(_04959_),
    .A(\mem_A[5] ),
    .B(_04238_));
 sg13g2_o21ai_1 _12853_ (.B1(_04951_),
    .Y(_04960_),
    .A1(_04949_),
    .A2(_04952_));
 sg13g2_a21oi_1 _12854_ (.A1(_04959_),
    .A2(_04960_),
    .Y(_04961_),
    .B1(net3059));
 sg13g2_o21ai_1 _12855_ (.B1(_04961_),
    .Y(_04962_),
    .A1(_04959_),
    .A2(_04960_));
 sg13g2_a21oi_1 _12856_ (.A1(_02160_),
    .A2(net3059),
    .Y(_04963_),
    .B1(net3048));
 sg13g2_a22oi_1 _12857_ (.Y(_04964_),
    .B1(_04962_),
    .B2(_04963_),
    .A2(net3047),
    .A1(net3347));
 sg13g2_nor2_1 _12858_ (.A(net3997),
    .B(_04964_),
    .Y(_00643_));
 sg13g2_or2_1 _12859_ (.X(_04965_),
    .B(_04959_),
    .A(_04952_));
 sg13g2_a21oi_1 _12860_ (.A1(_04950_),
    .A2(_04958_),
    .Y(_04966_),
    .B1(_04957_));
 sg13g2_o21ai_1 _12861_ (.B1(_04966_),
    .Y(_04967_),
    .A1(_04949_),
    .A2(_04965_));
 sg13g2_nor2_1 _12862_ (.A(_02129_),
    .B(_04533_),
    .Y(_04968_));
 sg13g2_xnor2_1 _12863_ (.Y(_04969_),
    .A(\mem_A[6] ),
    .B(_04533_));
 sg13g2_xnor2_1 _12864_ (.Y(_04970_),
    .A(_04967_),
    .B(_04969_));
 sg13g2_o21ai_1 _12865_ (.B1(_04919_),
    .Y(_04971_),
    .A1(net7),
    .A2(net3060));
 sg13g2_a21oi_1 _12866_ (.A1(net3060),
    .A2(_04970_),
    .Y(_04972_),
    .B1(_04971_));
 sg13g2_a21oi_1 _12867_ (.A1(net3296),
    .A2(net3047),
    .Y(_04973_),
    .B1(_04972_));
 sg13g2_nor2_1 _12868_ (.A(net3997),
    .B(_04973_),
    .Y(_00644_));
 sg13g2_a21oi_1 _12869_ (.A1(_04967_),
    .A2(_04969_),
    .Y(_04974_),
    .B1(_04968_));
 sg13g2_xnor2_1 _12870_ (.Y(_04975_),
    .A(\mem_A[7] ),
    .B(_04848_));
 sg13g2_or2_1 _12871_ (.X(_04976_),
    .B(_04975_),
    .A(_04974_));
 sg13g2_a21oi_1 _12872_ (.A1(_04974_),
    .A2(_04975_),
    .Y(_04977_),
    .B1(net3059));
 sg13g2_o21ai_1 _12873_ (.B1(_04919_),
    .Y(_04978_),
    .A1(net8),
    .A2(net3060));
 sg13g2_a21o_1 _12874_ (.A2(_04977_),
    .A1(_04976_),
    .B1(_04978_),
    .X(_04979_));
 sg13g2_nand2_1 _12875_ (.Y(_04980_),
    .A(net3256),
    .B(net3047));
 sg13g2_a21oi_1 _12876_ (.A1(_04979_),
    .A2(_04980_),
    .Y(_00645_),
    .B1(net3997));
 sg13g2_o21ai_1 _12877_ (.B1(net4009),
    .Y(_04981_),
    .A1(net5203),
    .A2(net3056));
 sg13g2_a21oi_1 _12878_ (.A1(net3056),
    .A2(_02847_),
    .Y(_00646_),
    .B1(_04981_));
 sg13g2_o21ai_1 _12879_ (.B1(net4008),
    .Y(_04982_),
    .A1(net5167),
    .A2(net3057));
 sg13g2_a21oi_1 _12880_ (.A1(net3056),
    .A2(_03131_),
    .Y(_00647_),
    .B1(_04982_));
 sg13g2_o21ai_1 _12881_ (.B1(net4003),
    .Y(_04983_),
    .A1(_02414_),
    .A2(_03426_));
 sg13g2_a21oi_1 _12882_ (.A1(_02130_),
    .A2(_02414_),
    .Y(_00648_),
    .B1(_04983_));
 sg13g2_o21ai_1 _12883_ (.B1(net4009),
    .Y(_04984_),
    .A1(net5208),
    .A2(net3056));
 sg13g2_a21oi_1 _12884_ (.A1(net3056),
    .A2(_03661_),
    .Y(_00649_),
    .B1(_04984_));
 sg13g2_o21ai_1 _12885_ (.B1(net4008),
    .Y(_04985_),
    .A1(net5207),
    .A2(net3056));
 sg13g2_a21oi_1 _12886_ (.A1(net3056),
    .A2(_03953_),
    .Y(_00650_),
    .B1(_04985_));
 sg13g2_o21ai_1 _12887_ (.B1(net4008),
    .Y(_04986_),
    .A1(net5209),
    .A2(net3057));
 sg13g2_a21oi_1 _12888_ (.A1(net3056),
    .A2(_04238_),
    .Y(_00651_),
    .B1(_04986_));
 sg13g2_o21ai_1 _12889_ (.B1(net4004),
    .Y(_04987_),
    .A1(_02414_),
    .A2(_04533_));
 sg13g2_a21oi_1 _12890_ (.A1(_02129_),
    .A2(_02414_),
    .Y(_00652_),
    .B1(_04987_));
 sg13g2_o21ai_1 _12891_ (.B1(net4003),
    .Y(_04988_),
    .A1(_02414_),
    .A2(_04848_));
 sg13g2_a21oi_1 _12892_ (.A1(_02128_),
    .A2(_02414_),
    .Y(_00653_),
    .B1(_04988_));
 sg13g2_nand2_2 _12893_ (.Y(_04989_),
    .A(net3083),
    .B(net3036));
 sg13g2_mux2_1 _12894_ (.A0(net3565),
    .A1(net4096),
    .S(_04989_),
    .X(_00654_));
 sg13g2_mux2_1 _12895_ (.A0(net3521),
    .A1(net4106),
    .S(_04989_),
    .X(_00655_));
 sg13g2_mux2_1 _12896_ (.A0(net3473),
    .A1(net5020),
    .S(_04989_),
    .X(_00656_));
 sg13g2_mux2_1 _12897_ (.A0(net3429),
    .A1(net2885),
    .S(_04989_),
    .X(_00657_));
 sg13g2_mux2_1 _12898_ (.A0(net3381),
    .A1(net5045),
    .S(_04989_),
    .X(_00658_));
 sg13g2_mux2_1 _12899_ (.A0(net3336),
    .A1(net4661),
    .S(_04989_),
    .X(_00659_));
 sg13g2_mux2_1 _12900_ (.A0(net3291),
    .A1(net4890),
    .S(_04989_),
    .X(_00660_));
 sg13g2_mux2_1 _12901_ (.A0(net3245),
    .A1(net4071),
    .S(_04989_),
    .X(_00661_));
 sg13g2_nor2_2 _12902_ (.A(_02268_),
    .B(_02298_),
    .Y(_04990_));
 sg13g2_mux2_1 _12903_ (.A0(net2503),
    .A1(net3569),
    .S(_04990_),
    .X(_00662_));
 sg13g2_mux2_1 _12904_ (.A0(net2671),
    .A1(net3521),
    .S(_04990_),
    .X(_00663_));
 sg13g2_mux2_1 _12905_ (.A0(net2770),
    .A1(net3473),
    .S(_04990_),
    .X(_00664_));
 sg13g2_mux2_1 _12906_ (.A0(net2576),
    .A1(net3429),
    .S(_04990_),
    .X(_00665_));
 sg13g2_mux2_1 _12907_ (.A0(net2444),
    .A1(net3381),
    .S(_04990_),
    .X(_00666_));
 sg13g2_mux2_1 _12908_ (.A0(net2662),
    .A1(net3336),
    .S(_04990_),
    .X(_00667_));
 sg13g2_mux2_1 _12909_ (.A0(net2651),
    .A1(net3291),
    .S(_04990_),
    .X(_00668_));
 sg13g2_mux2_1 _12910_ (.A0(net2244),
    .A1(net3245),
    .S(_04990_),
    .X(_00669_));
 sg13g2_nand2_2 _12911_ (.Y(_04991_),
    .A(net3037),
    .B(_02297_));
 sg13g2_mux2_1 _12912_ (.A0(net3591),
    .A1(net4066),
    .S(_04991_),
    .X(_00670_));
 sg13g2_mux2_1 _12913_ (.A0(net3547),
    .A1(net4810),
    .S(_04991_),
    .X(_00671_));
 sg13g2_mux2_1 _12914_ (.A0(net3501),
    .A1(net2960),
    .S(_04991_),
    .X(_00672_));
 sg13g2_mux2_1 _12915_ (.A0(net3455),
    .A1(net4551),
    .S(_04991_),
    .X(_00673_));
 sg13g2_mux2_1 _12916_ (.A0(net3409),
    .A1(net2913),
    .S(_04991_),
    .X(_00674_));
 sg13g2_mux2_1 _12917_ (.A0(net3365),
    .A1(net4315),
    .S(_04991_),
    .X(_00675_));
 sg13g2_mux2_1 _12918_ (.A0(net3319),
    .A1(net4388),
    .S(_04991_),
    .X(_00676_));
 sg13g2_mux2_1 _12919_ (.A0(net3270),
    .A1(net4982),
    .S(_04991_),
    .X(_00677_));
 sg13g2_nand2_2 _12920_ (.Y(_04992_),
    .A(net3080),
    .B(net3037));
 sg13g2_mux2_1 _12921_ (.A0(net3601),
    .A1(net4405),
    .S(_04992_),
    .X(_00678_));
 sg13g2_mux2_1 _12922_ (.A0(net3547),
    .A1(net4358),
    .S(_04992_),
    .X(_00679_));
 sg13g2_mux2_1 _12923_ (.A0(net3500),
    .A1(net4739),
    .S(_04992_),
    .X(_00680_));
 sg13g2_mux2_1 _12924_ (.A0(net3455),
    .A1(net4753),
    .S(_04992_),
    .X(_00681_));
 sg13g2_mux2_1 _12925_ (.A0(net3409),
    .A1(net4100),
    .S(_04992_),
    .X(_00682_));
 sg13g2_mux2_1 _12926_ (.A0(net3365),
    .A1(net3009),
    .S(_04992_),
    .X(_00683_));
 sg13g2_mux2_1 _12927_ (.A0(net3319),
    .A1(net4045),
    .S(_04992_),
    .X(_00684_));
 sg13g2_mux2_1 _12928_ (.A0(net3270),
    .A1(net4552),
    .S(_04992_),
    .X(_00685_));
 sg13g2_nand2_2 _12929_ (.Y(_04993_),
    .A(net3077),
    .B(net3034));
 sg13g2_mux2_1 _12930_ (.A0(net3593),
    .A1(net4113),
    .S(_04993_),
    .X(_00686_));
 sg13g2_mux2_1 _12931_ (.A0(net3546),
    .A1(net4735),
    .S(_04993_),
    .X(_00687_));
 sg13g2_mux2_1 _12932_ (.A0(net3501),
    .A1(net4234),
    .S(_04993_),
    .X(_00688_));
 sg13g2_mux2_1 _12933_ (.A0(net3456),
    .A1(net4168),
    .S(_04993_),
    .X(_00689_));
 sg13g2_mux2_1 _12934_ (.A0(net3408),
    .A1(net4076),
    .S(_04993_),
    .X(_00690_));
 sg13g2_mux2_1 _12935_ (.A0(net3368),
    .A1(net4844),
    .S(_04993_),
    .X(_00691_));
 sg13g2_mux2_1 _12936_ (.A0(net3320),
    .A1(net4027),
    .S(_04993_),
    .X(_00692_));
 sg13g2_mux2_1 _12937_ (.A0(net3271),
    .A1(net4986),
    .S(_04993_),
    .X(_00693_));
 sg13g2_nand2_2 _12938_ (.Y(_04994_),
    .A(net3085),
    .B(net3034));
 sg13g2_mux2_1 _12939_ (.A0(net3592),
    .A1(net5059),
    .S(_04994_),
    .X(_00694_));
 sg13g2_mux2_1 _12940_ (.A0(net3546),
    .A1(net5049),
    .S(_04994_),
    .X(_00695_));
 sg13g2_mux2_1 _12941_ (.A0(net3501),
    .A1(net2910),
    .S(_04994_),
    .X(_00696_));
 sg13g2_mux2_1 _12942_ (.A0(net3456),
    .A1(net5082),
    .S(_04994_),
    .X(_00697_));
 sg13g2_mux2_1 _12943_ (.A0(net3408),
    .A1(net4309),
    .S(_04994_),
    .X(_00698_));
 sg13g2_mux2_1 _12944_ (.A0(net3368),
    .A1(net4586),
    .S(_04994_),
    .X(_00699_));
 sg13g2_mux2_1 _12945_ (.A0(net3320),
    .A1(net4241),
    .S(_04994_),
    .X(_00700_));
 sg13g2_mux2_1 _12946_ (.A0(net3271),
    .A1(net4166),
    .S(_04994_),
    .X(_00701_));
 sg13g2_nand2_2 _12947_ (.Y(_04995_),
    .A(_02274_),
    .B(_02293_));
 sg13g2_mux2_1 _12948_ (.A0(net3590),
    .A1(net4459),
    .S(_04995_),
    .X(_00702_));
 sg13g2_mux2_1 _12949_ (.A0(net3545),
    .A1(net4490),
    .S(_04995_),
    .X(_00703_));
 sg13g2_mux2_1 _12950_ (.A0(net3499),
    .A1(net4518),
    .S(_04995_),
    .X(_00704_));
 sg13g2_mux2_1 _12951_ (.A0(net3454),
    .A1(net4245),
    .S(_04995_),
    .X(_00705_));
 sg13g2_mux2_1 _12952_ (.A0(net3408),
    .A1(net2834),
    .S(_04995_),
    .X(_00706_));
 sg13g2_mux2_1 _12953_ (.A0(net3355),
    .A1(net2701),
    .S(_04995_),
    .X(_00707_));
 sg13g2_mux2_1 _12954_ (.A0(net3320),
    .A1(net2800),
    .S(_04995_),
    .X(_00708_));
 sg13g2_mux2_1 _12955_ (.A0(net3269),
    .A1(net4854),
    .S(_04995_),
    .X(_00709_));
 sg13g2_nor2_2 _12956_ (.A(_02322_),
    .B(_02350_),
    .Y(_04996_));
 sg13g2_mux2_1 _12957_ (.A0(net2465),
    .A1(net3592),
    .S(_04996_),
    .X(_00710_));
 sg13g2_mux2_1 _12958_ (.A0(net2483),
    .A1(net3546),
    .S(_04996_),
    .X(_00711_));
 sg13g2_mux2_1 _12959_ (.A0(net2406),
    .A1(net3501),
    .S(_04996_),
    .X(_00712_));
 sg13g2_mux2_1 _12960_ (.A0(net2461),
    .A1(net3456),
    .S(_04996_),
    .X(_00713_));
 sg13g2_mux2_1 _12961_ (.A0(net2422),
    .A1(net3410),
    .S(_04996_),
    .X(_00714_));
 sg13g2_mux2_1 _12962_ (.A0(net2328),
    .A1(net3366),
    .S(_04996_),
    .X(_00715_));
 sg13g2_mux2_1 _12963_ (.A0(net2245),
    .A1(net3320),
    .S(_04996_),
    .X(_00716_));
 sg13g2_mux2_1 _12964_ (.A0(net2264),
    .A1(net3271),
    .S(_04996_),
    .X(_00717_));
 sg13g2_nand2_2 _12965_ (.Y(_04997_),
    .A(net3071),
    .B(net3035));
 sg13g2_mux2_1 _12966_ (.A0(net3593),
    .A1(net4367),
    .S(_04997_),
    .X(_00718_));
 sg13g2_mux2_1 _12967_ (.A0(net3549),
    .A1(net4964),
    .S(_04997_),
    .X(_00719_));
 sg13g2_mux2_1 _12968_ (.A0(net3502),
    .A1(net4461),
    .S(_04997_),
    .X(_00720_));
 sg13g2_mux2_1 _12969_ (.A0(net3457),
    .A1(net4730),
    .S(_04997_),
    .X(_00721_));
 sg13g2_mux2_1 _12970_ (.A0(net3411),
    .A1(net5107),
    .S(_04997_),
    .X(_00722_));
 sg13g2_mux2_1 _12971_ (.A0(net3367),
    .A1(net2992),
    .S(_04997_),
    .X(_00723_));
 sg13g2_mux2_1 _12972_ (.A0(net3321),
    .A1(net2943),
    .S(_04997_),
    .X(_00724_));
 sg13g2_mux2_1 _12973_ (.A0(net3272),
    .A1(net4935),
    .S(_04997_),
    .X(_00725_));
 sg13g2_nand2_2 _12974_ (.Y(_04998_),
    .A(_02330_),
    .B(net3035));
 sg13g2_mux2_1 _12975_ (.A0(net3593),
    .A1(net4654),
    .S(_04998_),
    .X(_00726_));
 sg13g2_mux2_1 _12976_ (.A0(net3549),
    .A1(net4222),
    .S(_04998_),
    .X(_00727_));
 sg13g2_mux2_1 _12977_ (.A0(net3502),
    .A1(net4190),
    .S(_04998_),
    .X(_00728_));
 sg13g2_mux2_1 _12978_ (.A0(net3457),
    .A1(net4685),
    .S(_04998_),
    .X(_00729_));
 sg13g2_mux2_1 _12979_ (.A0(net3411),
    .A1(net4626),
    .S(_04998_),
    .X(_00730_));
 sg13g2_mux2_1 _12980_ (.A0(net3367),
    .A1(net4891),
    .S(_04998_),
    .X(_00731_));
 sg13g2_mux2_1 _12981_ (.A0(net3322),
    .A1(net4959),
    .S(_04998_),
    .X(_00732_));
 sg13g2_mux2_1 _12982_ (.A0(net3272),
    .A1(net4726),
    .S(_04998_),
    .X(_00733_));
 sg13g2_nand2_2 _12983_ (.Y(_04999_),
    .A(net3070),
    .B(net3035));
 sg13g2_mux2_1 _12984_ (.A0(net3593),
    .A1(net5096),
    .S(_04999_),
    .X(_00734_));
 sg13g2_mux2_1 _12985_ (.A0(net3549),
    .A1(net4729),
    .S(_04999_),
    .X(_00735_));
 sg13g2_mux2_1 _12986_ (.A0(net3502),
    .A1(net4853),
    .S(_04999_),
    .X(_00736_));
 sg13g2_mux2_1 _12987_ (.A0(net3457),
    .A1(net5130),
    .S(_04999_),
    .X(_00737_));
 sg13g2_mux2_1 _12988_ (.A0(net3411),
    .A1(net2918),
    .S(_04999_),
    .X(_00738_));
 sg13g2_mux2_1 _12989_ (.A0(net3367),
    .A1(net5151),
    .S(_04999_),
    .X(_00739_));
 sg13g2_mux2_1 _12990_ (.A0(net3322),
    .A1(net2974),
    .S(_04999_),
    .X(_00740_));
 sg13g2_mux2_1 _12991_ (.A0(net3272),
    .A1(net2934),
    .S(_04999_),
    .X(_00741_));
 sg13g2_nor2_2 _12992_ (.A(_02255_),
    .B(_02322_),
    .Y(_05000_));
 sg13g2_mux2_1 _12993_ (.A0(net2332),
    .A1(net3573),
    .S(_05000_),
    .X(_00742_));
 sg13g2_mux2_1 _12994_ (.A0(net2253),
    .A1(net3528),
    .S(_05000_),
    .X(_00743_));
 sg13g2_mux2_1 _12995_ (.A0(net2322),
    .A1(net3480),
    .S(_05000_),
    .X(_00744_));
 sg13g2_mux2_1 _12996_ (.A0(net2540),
    .A1(net3434),
    .S(_05000_),
    .X(_00745_));
 sg13g2_mux2_1 _12997_ (.A0(net2269),
    .A1(net3387),
    .S(_05000_),
    .X(_00746_));
 sg13g2_mux2_1 _12998_ (.A0(net2558),
    .A1(net3346),
    .S(_05000_),
    .X(_00747_));
 sg13g2_mux2_1 _12999_ (.A0(net2598),
    .A1(net3299),
    .S(_05000_),
    .X(_00748_));
 sg13g2_mux2_1 _13000_ (.A0(net2231),
    .A1(net3251),
    .S(_05000_),
    .X(_00749_));
 sg13g2_nor2_2 _13001_ (.A(_02255_),
    .B(net3039),
    .Y(_05001_));
 sg13g2_nand2_2 _13002_ (.Y(_05002_),
    .A(_02254_),
    .B(net3042));
 sg13g2_nor2_2 _13003_ (.A(_02335_),
    .B(_05002_),
    .Y(_05003_));
 sg13g2_mux2_1 _13004_ (.A0(net2256),
    .A1(net3574),
    .S(_05003_),
    .X(_00750_));
 sg13g2_mux2_1 _13005_ (.A0(net2450),
    .A1(net3526),
    .S(_05003_),
    .X(_00751_));
 sg13g2_mux2_1 _13006_ (.A0(net2197),
    .A1(net3481),
    .S(_05003_),
    .X(_00752_));
 sg13g2_mux2_1 _13007_ (.A0(net2419),
    .A1(net3434),
    .S(_05003_),
    .X(_00753_));
 sg13g2_mux2_1 _13008_ (.A0(net2398),
    .A1(net3388),
    .S(_05003_),
    .X(_00754_));
 sg13g2_mux2_1 _13009_ (.A0(net2241),
    .A1(net3343),
    .S(_05003_),
    .X(_00755_));
 sg13g2_mux2_1 _13010_ (.A0(net2443),
    .A1(net3297),
    .S(_05003_),
    .X(_00756_));
 sg13g2_mux2_1 _13011_ (.A0(net2428),
    .A1(net3252),
    .S(_05003_),
    .X(_00757_));
 sg13g2_nand2_2 _13012_ (.Y(_05004_),
    .A(_02297_),
    .B(_02375_));
 sg13g2_mux2_1 _13013_ (.A0(net3597),
    .A1(net4533),
    .S(_05004_),
    .X(_00758_));
 sg13g2_mux2_1 _13014_ (.A0(net3552),
    .A1(net4176),
    .S(_05004_),
    .X(_00759_));
 sg13g2_mux2_1 _13015_ (.A0(net3505),
    .A1(net4622),
    .S(_05004_),
    .X(_00760_));
 sg13g2_mux2_1 _13016_ (.A0(net3461),
    .A1(net5038),
    .S(_05004_),
    .X(_00761_));
 sg13g2_mux2_1 _13017_ (.A0(net3413),
    .A1(net4141),
    .S(_05004_),
    .X(_00762_));
 sg13g2_mux2_1 _13018_ (.A0(net3369),
    .A1(net4205),
    .S(_05004_),
    .X(_00763_));
 sg13g2_mux2_1 _13019_ (.A0(net3323),
    .A1(net4780),
    .S(_05004_),
    .X(_00764_));
 sg13g2_mux2_1 _13020_ (.A0(net3277),
    .A1(net4246),
    .S(_05004_),
    .X(_00765_));
 sg13g2_nand2_2 _13021_ (.Y(_05005_),
    .A(net3038),
    .B(_02309_));
 sg13g2_mux2_1 _13022_ (.A0(net3592),
    .A1(net4110),
    .S(_05005_),
    .X(_00766_));
 sg13g2_mux2_1 _13023_ (.A0(net3548),
    .A1(net5062),
    .S(_05005_),
    .X(_00767_));
 sg13g2_mux2_1 _13024_ (.A0(net3503),
    .A1(net4111),
    .S(_05005_),
    .X(_00768_));
 sg13g2_mux2_1 _13025_ (.A0(net3458),
    .A1(net4454),
    .S(_05005_),
    .X(_00769_));
 sg13g2_mux2_1 _13026_ (.A0(net3412),
    .A1(net4978),
    .S(_05005_),
    .X(_00770_));
 sg13g2_mux2_1 _13027_ (.A0(net3368),
    .A1(net4624),
    .S(_05005_),
    .X(_00771_));
 sg13g2_mux2_1 _13028_ (.A0(net3322),
    .A1(net2961),
    .S(_05005_),
    .X(_00772_));
 sg13g2_mux2_1 _13029_ (.A0(net3273),
    .A1(net4333),
    .S(_05005_),
    .X(_00773_));
 sg13g2_nor2_2 _13030_ (.A(_02253_),
    .B(_02290_),
    .Y(_05006_));
 sg13g2_and2_2 _13031_ (.A(net3043),
    .B(net3051),
    .X(_05007_));
 sg13g2_nand2_2 _13032_ (.Y(_05008_),
    .A(net3043),
    .B(_05006_));
 sg13g2_nor2_2 _13033_ (.A(_02307_),
    .B(_05008_),
    .Y(_05009_));
 sg13g2_mux2_1 _13034_ (.A0(net2220),
    .A1(net3575),
    .S(_05009_),
    .X(_00774_));
 sg13g2_mux2_1 _13035_ (.A0(net2415),
    .A1(net3527),
    .S(_05009_),
    .X(_00775_));
 sg13g2_mux2_1 _13036_ (.A0(net2686),
    .A1(net3489),
    .S(_05009_),
    .X(_00776_));
 sg13g2_mux2_1 _13037_ (.A0(net2815),
    .A1(net3436),
    .S(_05009_),
    .X(_00777_));
 sg13g2_mux2_1 _13038_ (.A0(net2474),
    .A1(net3397),
    .S(_05009_),
    .X(_00778_));
 sg13g2_mux2_1 _13039_ (.A0(net2589),
    .A1(net3345),
    .S(_05009_),
    .X(_00779_));
 sg13g2_mux2_1 _13040_ (.A0(net2275),
    .A1(net3299),
    .S(_05009_),
    .X(_00780_));
 sg13g2_mux2_1 _13041_ (.A0(net2390),
    .A1(net3258),
    .S(_05009_),
    .X(_00781_));
 sg13g2_nand2_2 _13042_ (.Y(_05010_),
    .A(_02346_),
    .B(net3051));
 sg13g2_mux2_1 _13043_ (.A0(net3582),
    .A1(net4597),
    .S(_05010_),
    .X(_00782_));
 sg13g2_mux2_1 _13044_ (.A0(net3536),
    .A1(net5001),
    .S(_05010_),
    .X(_00783_));
 sg13g2_mux2_1 _13045_ (.A0(net3493),
    .A1(net4406),
    .S(_05010_),
    .X(_00784_));
 sg13g2_mux2_1 _13046_ (.A0(net3443),
    .A1(net5064),
    .S(_05010_),
    .X(_00785_));
 sg13g2_mux2_1 _13047_ (.A0(net3401),
    .A1(net5118),
    .S(_05010_),
    .X(_00786_));
 sg13g2_mux2_1 _13048_ (.A0(net3355),
    .A1(net4998),
    .S(_05010_),
    .X(_00787_));
 sg13g2_mux2_1 _13049_ (.A0(net3310),
    .A1(net4540),
    .S(_05010_),
    .X(_00788_));
 sg13g2_mux2_1 _13050_ (.A0(net3262),
    .A1(net4084),
    .S(_05010_),
    .X(_00789_));
 sg13g2_nand2_2 _13051_ (.Y(_05011_),
    .A(net3074),
    .B(net3034));
 sg13g2_mux2_1 _13052_ (.A0(net3593),
    .A1(net4605),
    .S(_05011_),
    .X(_00790_));
 sg13g2_mux2_1 _13053_ (.A0(net3546),
    .A1(net4121),
    .S(_05011_),
    .X(_00791_));
 sg13g2_mux2_1 _13054_ (.A0(net3502),
    .A1(net4833),
    .S(_05011_),
    .X(_00792_));
 sg13g2_mux2_1 _13055_ (.A0(net3456),
    .A1(net4442),
    .S(_05011_),
    .X(_00793_));
 sg13g2_mux2_1 _13056_ (.A0(net3410),
    .A1(net4278),
    .S(_05011_),
    .X(_00794_));
 sg13g2_mux2_1 _13057_ (.A0(net3368),
    .A1(net4709),
    .S(_05011_),
    .X(_00795_));
 sg13g2_mux2_1 _13058_ (.A0(net3319),
    .A1(net4156),
    .S(_05011_),
    .X(_00796_));
 sg13g2_mux2_1 _13059_ (.A0(net3271),
    .A1(net4274),
    .S(_05011_),
    .X(_00797_));
 sg13g2_nand2_2 _13060_ (.Y(_05012_),
    .A(net3078),
    .B(_02328_));
 sg13g2_mux2_1 _13061_ (.A0(net3562),
    .A1(net4869),
    .S(_05012_),
    .X(_00798_));
 sg13g2_mux2_1 _13062_ (.A0(net3516),
    .A1(net4777),
    .S(_05012_),
    .X(_00799_));
 sg13g2_mux2_1 _13063_ (.A0(net3478),
    .A1(net4073),
    .S(_05012_),
    .X(_00800_));
 sg13g2_mux2_1 _13064_ (.A0(net3432),
    .A1(net4488),
    .S(_05012_),
    .X(_00801_));
 sg13g2_mux2_1 _13065_ (.A0(net3379),
    .A1(net4148),
    .S(_05012_),
    .X(_00802_));
 sg13g2_mux2_1 _13066_ (.A0(net3333),
    .A1(net5136),
    .S(_05012_),
    .X(_00803_));
 sg13g2_mux2_1 _13067_ (.A0(net3288),
    .A1(net4147),
    .S(_05012_),
    .X(_00804_));
 sg13g2_mux2_1 _13068_ (.A0(net3241),
    .A1(net4480),
    .S(_05012_),
    .X(_00805_));
 sg13g2_nor3_1 _13069_ (.A(net3039),
    .B(_02265_),
    .C(_02290_),
    .Y(_05013_));
 sg13g2_and2_2 _13070_ (.A(_02297_),
    .B(net3024),
    .X(_05014_));
 sg13g2_mux2_1 _13071_ (.A0(net2527),
    .A1(net3585),
    .S(_05014_),
    .X(_00806_));
 sg13g2_mux2_1 _13072_ (.A0(net2700),
    .A1(net3541),
    .S(_05014_),
    .X(_00807_));
 sg13g2_mux2_1 _13073_ (.A0(net2575),
    .A1(net3495),
    .S(_05014_),
    .X(_00808_));
 sg13g2_mux2_1 _13074_ (.A0(net2531),
    .A1(net3453),
    .S(_05014_),
    .X(_00809_));
 sg13g2_mux2_1 _13075_ (.A0(net2363),
    .A1(net3403),
    .S(_05014_),
    .X(_00810_));
 sg13g2_mux2_1 _13076_ (.A0(net2412),
    .A1(net3360),
    .S(_05014_),
    .X(_00811_));
 sg13g2_mux2_1 _13077_ (.A0(net2525),
    .A1(net3314),
    .S(_05014_),
    .X(_00812_));
 sg13g2_mux2_1 _13078_ (.A0(net2306),
    .A1(net3264),
    .S(_05014_),
    .X(_00813_));
 sg13g2_nand2_2 _13079_ (.Y(_05015_),
    .A(net3080),
    .B(net3024));
 sg13g2_mux2_1 _13080_ (.A0(net3585),
    .A1(net4602),
    .S(_05015_),
    .X(_00814_));
 sg13g2_mux2_1 _13081_ (.A0(net3541),
    .A1(net2693),
    .S(_05015_),
    .X(_00815_));
 sg13g2_mux2_1 _13082_ (.A0(net3495),
    .A1(net4638),
    .S(_05015_),
    .X(_00816_));
 sg13g2_mux2_1 _13083_ (.A0(net3449),
    .A1(net2962),
    .S(_05015_),
    .X(_00817_));
 sg13g2_mux2_1 _13084_ (.A0(net3404),
    .A1(net2970),
    .S(_05015_),
    .X(_00818_));
 sg13g2_mux2_1 _13085_ (.A0(net3360),
    .A1(net2811),
    .S(_05015_),
    .X(_00819_));
 sg13g2_mux2_1 _13086_ (.A0(net3315),
    .A1(net2971),
    .S(_05015_),
    .X(_00820_));
 sg13g2_mux2_1 _13087_ (.A0(net3264),
    .A1(net2920),
    .S(_05015_),
    .X(_00821_));
 sg13g2_nor2_2 _13088_ (.A(_02268_),
    .B(net3076),
    .Y(_05016_));
 sg13g2_mux2_1 _13089_ (.A0(net2217),
    .A1(net3568),
    .S(_05016_),
    .X(_00822_));
 sg13g2_mux2_1 _13090_ (.A0(net2374),
    .A1(net3520),
    .S(_05016_),
    .X(_00823_));
 sg13g2_mux2_1 _13091_ (.A0(net2592),
    .A1(net3474),
    .S(_05016_),
    .X(_00824_));
 sg13g2_mux2_1 _13092_ (.A0(net2358),
    .A1(net3428),
    .S(_05016_),
    .X(_00825_));
 sg13g2_mux2_1 _13093_ (.A0(net2317),
    .A1(net3382),
    .S(_05016_),
    .X(_00826_));
 sg13g2_mux2_1 _13094_ (.A0(net2514),
    .A1(net3337),
    .S(_05016_),
    .X(_00827_));
 sg13g2_mux2_1 _13095_ (.A0(net2706),
    .A1(net3292),
    .S(_05016_),
    .X(_00828_));
 sg13g2_mux2_1 _13096_ (.A0(net2480),
    .A1(net3244),
    .S(_05016_),
    .X(_00829_));
 sg13g2_nand2_2 _13097_ (.Y(_05017_),
    .A(_02284_),
    .B(net3036));
 sg13g2_mux2_1 _13098_ (.A0(net3597),
    .A1(net4611),
    .S(_05017_),
    .X(_00830_));
 sg13g2_mux2_1 _13099_ (.A0(net3552),
    .A1(net4760),
    .S(_05017_),
    .X(_00831_));
 sg13g2_mux2_1 _13100_ (.A0(net3505),
    .A1(net2846),
    .S(_05017_),
    .X(_00832_));
 sg13g2_mux2_1 _13101_ (.A0(net3461),
    .A1(net2816),
    .S(_05017_),
    .X(_00833_));
 sg13g2_mux2_1 _13102_ (.A0(net3413),
    .A1(net4723),
    .S(_05017_),
    .X(_00834_));
 sg13g2_mux2_1 _13103_ (.A0(net3369),
    .A1(net4775),
    .S(_05017_),
    .X(_00835_));
 sg13g2_mux2_1 _13104_ (.A0(net3323),
    .A1(net4855),
    .S(_05017_),
    .X(_00836_));
 sg13g2_mux2_1 _13105_ (.A0(net3277),
    .A1(net2904),
    .S(_05017_),
    .X(_00837_));
 sg13g2_nand2_1 _13106_ (.Y(_05018_),
    .A(net3084),
    .B(_02254_));
 sg13g2_o21ai_1 _13107_ (.B1(net4009),
    .Y(_05019_),
    .A1(\mem.out_strobe ),
    .A2(net2130));
 sg13g2_a21oi_1 _13108_ (.A1(net2130),
    .A2(_05018_),
    .Y(_00838_),
    .B1(_05019_));
 sg13g2_or3_2 _13109_ (.A(_00008_),
    .B(_02247_),
    .C(_02257_),
    .X(_05020_));
 sg13g2_o21ai_1 _13110_ (.B1(net4002),
    .Y(_05021_),
    .A1(net3568),
    .A2(net3046));
 sg13g2_a21oi_1 _13111_ (.A1(_02127_),
    .A2(_05020_),
    .Y(_00839_),
    .B1(_05021_));
 sg13g2_o21ai_1 _13112_ (.B1(net4003),
    .Y(_05022_),
    .A1(net3522),
    .A2(net3046));
 sg13g2_a21oi_1 _13113_ (.A1(_02126_),
    .A2(net3046),
    .Y(_00840_),
    .B1(_05022_));
 sg13g2_o21ai_1 _13114_ (.B1(net4002),
    .Y(_05023_),
    .A1(net3475),
    .A2(net3045));
 sg13g2_a21oi_1 _13115_ (.A1(_02125_),
    .A2(net3045),
    .Y(_00841_),
    .B1(_05023_));
 sg13g2_o21ai_1 _13116_ (.B1(net4002),
    .Y(_05024_),
    .A1(net3431),
    .A2(net3045));
 sg13g2_a21oi_1 _13117_ (.A1(_02124_),
    .A2(net3045),
    .Y(_00842_),
    .B1(_05024_));
 sg13g2_o21ai_1 _13118_ (.B1(net4002),
    .Y(_05025_),
    .A1(net3383),
    .A2(net3045));
 sg13g2_a21oi_1 _13119_ (.A1(_02123_),
    .A2(net3046),
    .Y(_00843_),
    .B1(_05025_));
 sg13g2_o21ai_1 _13120_ (.B1(net4002),
    .Y(_05026_),
    .A1(net3337),
    .A2(net3045));
 sg13g2_a21oi_1 _13121_ (.A1(_02122_),
    .A2(net3045),
    .Y(_00844_),
    .B1(_05026_));
 sg13g2_o21ai_1 _13122_ (.B1(net4002),
    .Y(_05027_),
    .A1(net3292),
    .A2(net3045));
 sg13g2_a21oi_1 _13123_ (.A1(_02121_),
    .A2(net3046),
    .Y(_00845_),
    .B1(_05027_));
 sg13g2_o21ai_1 _13124_ (.B1(net4002),
    .Y(_05028_),
    .A1(net3247),
    .A2(net3046));
 sg13g2_a21oi_1 _13125_ (.A1(_02120_),
    .A2(net3046),
    .Y(_00846_),
    .B1(_05028_));
 sg13g2_nand2_2 _13126_ (.Y(_05029_),
    .A(net3074),
    .B(net3026));
 sg13g2_mux2_1 _13127_ (.A0(net3585),
    .A1(net2914),
    .S(_05029_),
    .X(_00847_));
 sg13g2_mux2_1 _13128_ (.A0(net3541),
    .A1(net4678),
    .S(_05029_),
    .X(_00848_));
 sg13g2_mux2_1 _13129_ (.A0(net3498),
    .A1(net4292),
    .S(_05029_),
    .X(_00849_));
 sg13g2_mux2_1 _13130_ (.A0(net3449),
    .A1(net4641),
    .S(_05029_),
    .X(_00850_));
 sg13g2_mux2_1 _13131_ (.A0(net3393),
    .A1(net4108),
    .S(_05029_),
    .X(_00851_));
 sg13g2_mux2_1 _13132_ (.A0(net3360),
    .A1(net4617),
    .S(_05029_),
    .X(_00852_));
 sg13g2_mux2_1 _13133_ (.A0(net3314),
    .A1(net4283),
    .S(_05029_),
    .X(_00853_));
 sg13g2_mux2_1 _13134_ (.A0(net3265),
    .A1(net4821),
    .S(_05029_),
    .X(_00854_));
 sg13g2_nand2_2 _13135_ (.Y(_05030_),
    .A(_02349_),
    .B(net3025));
 sg13g2_mux2_1 _13136_ (.A0(net3585),
    .A1(net4257),
    .S(_05030_),
    .X(_00855_));
 sg13g2_mux2_1 _13137_ (.A0(net3540),
    .A1(net4970),
    .S(_05030_),
    .X(_00856_));
 sg13g2_mux2_1 _13138_ (.A0(net3495),
    .A1(net4593),
    .S(_05030_),
    .X(_00857_));
 sg13g2_mux2_1 _13139_ (.A0(net3451),
    .A1(net4064),
    .S(_05030_),
    .X(_00858_));
 sg13g2_mux2_1 _13140_ (.A0(net3403),
    .A1(net4545),
    .S(_05030_),
    .X(_00859_));
 sg13g2_mux2_1 _13141_ (.A0(net3359),
    .A1(net5127),
    .S(_05030_),
    .X(_00860_));
 sg13g2_mux2_1 _13142_ (.A0(net3314),
    .A1(net4085),
    .S(_05030_),
    .X(_00861_));
 sg13g2_mux2_1 _13143_ (.A0(net3265),
    .A1(net4879),
    .S(_05030_),
    .X(_00862_));
 sg13g2_nor2_2 _13144_ (.A(_02268_),
    .B(_02335_),
    .Y(_05031_));
 sg13g2_mux2_1 _13145_ (.A0(net2468),
    .A1(net3568),
    .S(_05031_),
    .X(_00863_));
 sg13g2_mux2_1 _13146_ (.A0(net2752),
    .A1(net3520),
    .S(_05031_),
    .X(_00864_));
 sg13g2_mux2_1 _13147_ (.A0(net2681),
    .A1(net3473),
    .S(_05031_),
    .X(_00865_));
 sg13g2_mux2_1 _13148_ (.A0(net2559),
    .A1(net3428),
    .S(_05031_),
    .X(_00866_));
 sg13g2_mux2_1 _13149_ (.A0(net2615),
    .A1(net3382),
    .S(_05031_),
    .X(_00867_));
 sg13g2_mux2_1 _13150_ (.A0(net2688),
    .A1(net3336),
    .S(_05031_),
    .X(_00868_));
 sg13g2_mux2_1 _13151_ (.A0(net2486),
    .A1(net3292),
    .S(_05031_),
    .X(_00869_));
 sg13g2_mux2_1 _13152_ (.A0(net2316),
    .A1(net3244),
    .S(_05031_),
    .X(_00870_));
 sg13g2_nand2_2 _13153_ (.Y(_05032_),
    .A(net3071),
    .B(_02370_));
 sg13g2_mux2_1 _13154_ (.A0(net3584),
    .A1(net4493),
    .S(_05032_),
    .X(_00871_));
 sg13g2_mux2_1 _13155_ (.A0(net3540),
    .A1(net4385),
    .S(_05032_),
    .X(_00872_));
 sg13g2_mux2_1 _13156_ (.A0(net3498),
    .A1(net4122),
    .S(_05032_),
    .X(_00873_));
 sg13g2_mux2_1 _13157_ (.A0(net3447),
    .A1(net5086),
    .S(_05032_),
    .X(_00874_));
 sg13g2_mux2_1 _13158_ (.A0(net3403),
    .A1(net4873),
    .S(_05032_),
    .X(_00875_));
 sg13g2_mux2_1 _13159_ (.A0(net3359),
    .A1(net4252),
    .S(_05032_),
    .X(_00876_));
 sg13g2_mux2_1 _13160_ (.A0(net3315),
    .A1(net5094),
    .S(_05032_),
    .X(_00877_));
 sg13g2_mux2_1 _13161_ (.A0(net3264),
    .A1(net4317),
    .S(_05032_),
    .X(_00878_));
 sg13g2_and2_2 _13162_ (.A(_02288_),
    .B(net3024),
    .X(_05033_));
 sg13g2_mux2_1 _13163_ (.A0(net2715),
    .A1(net3585),
    .S(_05033_),
    .X(_00879_));
 sg13g2_mux2_1 _13164_ (.A0(net2189),
    .A1(net3541),
    .S(_05033_),
    .X(_00880_));
 sg13g2_mux2_1 _13165_ (.A0(net2387),
    .A1(net3495),
    .S(_05033_),
    .X(_00881_));
 sg13g2_mux2_1 _13166_ (.A0(net2378),
    .A1(net3449),
    .S(_05033_),
    .X(_00882_));
 sg13g2_mux2_1 _13167_ (.A0(net2305),
    .A1(net3403),
    .S(_05033_),
    .X(_00883_));
 sg13g2_mux2_1 _13168_ (.A0(net2138),
    .A1(net3360),
    .S(_05033_),
    .X(_00884_));
 sg13g2_mux2_1 _13169_ (.A0(net2724),
    .A1(net3314),
    .S(_05033_),
    .X(_00885_));
 sg13g2_mux2_1 _13170_ (.A0(net2209),
    .A1(net3265),
    .S(_05033_),
    .X(_00886_));
 sg13g2_nand2_2 _13171_ (.Y(_05034_),
    .A(net3082),
    .B(_02283_));
 sg13g2_mux2_1 _13172_ (.A0(net3590),
    .A1(net2897),
    .S(_05034_),
    .X(_00887_));
 sg13g2_mux2_1 _13173_ (.A0(net3545),
    .A1(net4364),
    .S(_05034_),
    .X(_00888_));
 sg13g2_mux2_1 _13174_ (.A0(net3499),
    .A1(net4880),
    .S(_05034_),
    .X(_00889_));
 sg13g2_mux2_1 _13175_ (.A0(net3454),
    .A1(net4348),
    .S(_05034_),
    .X(_00890_));
 sg13g2_mux2_1 _13176_ (.A0(net3400),
    .A1(net2788),
    .S(_05034_),
    .X(_00891_));
 sg13g2_mux2_1 _13177_ (.A0(net3355),
    .A1(net2825),
    .S(_05034_),
    .X(_00892_));
 sg13g2_mux2_1 _13178_ (.A0(net3310),
    .A1(net2721),
    .S(_05034_),
    .X(_00893_));
 sg13g2_mux2_1 _13179_ (.A0(net3269),
    .A1(net4194),
    .S(_05034_),
    .X(_00894_));
 sg13g2_nand2_2 _13180_ (.Y(_05035_),
    .A(_02277_),
    .B(net3025));
 sg13g2_mux2_1 _13181_ (.A0(net3587),
    .A1(net2990),
    .S(_05035_),
    .X(_00895_));
 sg13g2_mux2_1 _13182_ (.A0(net3543),
    .A1(net4804),
    .S(_05035_),
    .X(_00896_));
 sg13g2_mux2_1 _13183_ (.A0(net3496),
    .A1(net4764),
    .S(_05035_),
    .X(_00897_));
 sg13g2_mux2_1 _13184_ (.A0(net3451),
    .A1(net4065),
    .S(_05035_),
    .X(_00898_));
 sg13g2_mux2_1 _13185_ (.A0(net3405),
    .A1(net2941),
    .S(_05035_),
    .X(_00899_));
 sg13g2_mux2_1 _13186_ (.A0(net3362),
    .A1(net2807),
    .S(_05035_),
    .X(_00900_));
 sg13g2_mux2_1 _13187_ (.A0(net3316),
    .A1(net2969),
    .S(_05035_),
    .X(_00901_));
 sg13g2_mux2_1 _13188_ (.A0(net3266),
    .A1(net4613),
    .S(_05035_),
    .X(_00902_));
 sg13g2_nand2_2 _13189_ (.Y(_05036_),
    .A(net3069),
    .B(net3025));
 sg13g2_mux2_1 _13190_ (.A0(net3588),
    .A1(net4325),
    .S(_05036_),
    .X(_00903_));
 sg13g2_mux2_1 _13191_ (.A0(net3543),
    .A1(net4811),
    .S(_05036_),
    .X(_00904_));
 sg13g2_mux2_1 _13192_ (.A0(net3496),
    .A1(net4965),
    .S(_05036_),
    .X(_00905_));
 sg13g2_mux2_1 _13193_ (.A0(net3451),
    .A1(net4789),
    .S(_05036_),
    .X(_00906_));
 sg13g2_mux2_1 _13194_ (.A0(net3405),
    .A1(net4990),
    .S(_05036_),
    .X(_00907_));
 sg13g2_mux2_1 _13195_ (.A0(net3362),
    .A1(net4532),
    .S(_05036_),
    .X(_00908_));
 sg13g2_mux2_1 _13196_ (.A0(net3316),
    .A1(net4095),
    .S(_05036_),
    .X(_00909_));
 sg13g2_mux2_1 _13197_ (.A0(net3266),
    .A1(net4057),
    .S(_05036_),
    .X(_00910_));
 sg13g2_nand2_2 _13198_ (.Y(_05037_),
    .A(_02383_),
    .B(net3025));
 sg13g2_mux2_1 _13199_ (.A0(net3588),
    .A1(net4042),
    .S(_05037_),
    .X(_00911_));
 sg13g2_mux2_1 _13200_ (.A0(net3543),
    .A1(net4203),
    .S(_05037_),
    .X(_00912_));
 sg13g2_mux2_1 _13201_ (.A0(net3495),
    .A1(net4633),
    .S(_05037_),
    .X(_00913_));
 sg13g2_mux2_1 _13202_ (.A0(net3451),
    .A1(net2889),
    .S(_05037_),
    .X(_00914_));
 sg13g2_mux2_1 _13203_ (.A0(net3405),
    .A1(net4182),
    .S(_05037_),
    .X(_00915_));
 sg13g2_mux2_1 _13204_ (.A0(net3361),
    .A1(net4671),
    .S(_05037_),
    .X(_00916_));
 sg13g2_mux2_1 _13205_ (.A0(net3316),
    .A1(net5010),
    .S(_05037_),
    .X(_00917_));
 sg13g2_mux2_1 _13206_ (.A0(net3267),
    .A1(net5177),
    .S(_05037_),
    .X(_00918_));
 sg13g2_nand2_2 _13207_ (.Y(_05038_),
    .A(_02309_),
    .B(net3025));
 sg13g2_mux2_1 _13208_ (.A0(net3588),
    .A1(net2909),
    .S(_05038_),
    .X(_00919_));
 sg13g2_mux2_1 _13209_ (.A0(net3543),
    .A1(net4179),
    .S(_05038_),
    .X(_00920_));
 sg13g2_mux2_1 _13210_ (.A0(net3497),
    .A1(net4498),
    .S(_05038_),
    .X(_00921_));
 sg13g2_mux2_1 _13211_ (.A0(net3451),
    .A1(net4189),
    .S(_05038_),
    .X(_00922_));
 sg13g2_mux2_1 _13212_ (.A0(net3405),
    .A1(net5023),
    .S(_05038_),
    .X(_00923_));
 sg13g2_mux2_1 _13213_ (.A0(net3361),
    .A1(net2946),
    .S(_05038_),
    .X(_00924_));
 sg13g2_mux2_1 _13214_ (.A0(net3316),
    .A1(net4542),
    .S(_05038_),
    .X(_00925_));
 sg13g2_mux2_1 _13215_ (.A0(net3266),
    .A1(net4632),
    .S(_05038_),
    .X(_00926_));
 sg13g2_and2_2 _13216_ (.A(_02337_),
    .B(net3024),
    .X(_05039_));
 sg13g2_mux2_1 _13217_ (.A0(net2456),
    .A1(net3587),
    .S(_05039_),
    .X(_00927_));
 sg13g2_mux2_1 _13218_ (.A0(net2266),
    .A1(net3543),
    .S(_05039_),
    .X(_00928_));
 sg13g2_mux2_1 _13219_ (.A0(net2309),
    .A1(net3496),
    .S(_05039_),
    .X(_00929_));
 sg13g2_mux2_1 _13220_ (.A0(net2485),
    .A1(net3451),
    .S(_05039_),
    .X(_00930_));
 sg13g2_mux2_1 _13221_ (.A0(net2657),
    .A1(net3404),
    .S(_05039_),
    .X(_00931_));
 sg13g2_mux2_1 _13222_ (.A0(net2196),
    .A1(net3361),
    .S(_05039_),
    .X(_00932_));
 sg13g2_mux2_1 _13223_ (.A0(net2537),
    .A1(net3314),
    .S(_05039_),
    .X(_00933_));
 sg13g2_mux2_1 _13224_ (.A0(net2665),
    .A1(net3267),
    .S(_05039_),
    .X(_00934_));
 sg13g2_nand2_2 _13225_ (.Y(_05040_),
    .A(_02334_),
    .B(net3024));
 sg13g2_mux2_1 _13226_ (.A0(net3587),
    .A1(net4082),
    .S(_05040_),
    .X(_00935_));
 sg13g2_mux2_1 _13227_ (.A0(net3543),
    .A1(net2958),
    .S(_05040_),
    .X(_00936_));
 sg13g2_mux2_1 _13228_ (.A0(net3495),
    .A1(net5121),
    .S(_05040_),
    .X(_00937_));
 sg13g2_mux2_1 _13229_ (.A0(net3451),
    .A1(net4748),
    .S(_05040_),
    .X(_00938_));
 sg13g2_mux2_1 _13230_ (.A0(net3404),
    .A1(net4705),
    .S(_05040_),
    .X(_00939_));
 sg13g2_mux2_1 _13231_ (.A0(net3361),
    .A1(net4762),
    .S(_05040_),
    .X(_00940_));
 sg13g2_mux2_1 _13232_ (.A0(net3315),
    .A1(net4791),
    .S(_05040_),
    .X(_00941_));
 sg13g2_mux2_1 _13233_ (.A0(net3267),
    .A1(net4417),
    .S(_05040_),
    .X(_00942_));
 sg13g2_nand2_2 _13234_ (.Y(_05041_),
    .A(_02330_),
    .B(net3025));
 sg13g2_mux2_1 _13235_ (.A0(net3587),
    .A1(net2931),
    .S(_05041_),
    .X(_00943_));
 sg13g2_mux2_1 _13236_ (.A0(net3542),
    .A1(net4401),
    .S(_05041_),
    .X(_00944_));
 sg13g2_mux2_1 _13237_ (.A0(net3495),
    .A1(net4884),
    .S(_05041_),
    .X(_00945_));
 sg13g2_mux2_1 _13238_ (.A0(net3451),
    .A1(net2944),
    .S(_05041_),
    .X(_00946_));
 sg13g2_mux2_1 _13239_ (.A0(net3403),
    .A1(net4619),
    .S(_05041_),
    .X(_00947_));
 sg13g2_mux2_1 _13240_ (.A0(net3361),
    .A1(net2812),
    .S(_05041_),
    .X(_00948_));
 sg13g2_mux2_1 _13241_ (.A0(net3314),
    .A1(net4966),
    .S(_05041_),
    .X(_00949_));
 sg13g2_mux2_1 _13242_ (.A0(net3267),
    .A1(net4174),
    .S(_05041_),
    .X(_00950_));
 sg13g2_nand2_2 _13243_ (.Y(_05042_),
    .A(_02327_),
    .B(net3024));
 sg13g2_mux2_1 _13244_ (.A0(net3587),
    .A1(net2978),
    .S(_05042_),
    .X(_00951_));
 sg13g2_mux2_1 _13245_ (.A0(net3542),
    .A1(net2994),
    .S(_05042_),
    .X(_00952_));
 sg13g2_mux2_1 _13246_ (.A0(net3495),
    .A1(net5076),
    .S(_05042_),
    .X(_00953_));
 sg13g2_mux2_1 _13247_ (.A0(net3452),
    .A1(net4118),
    .S(_05042_),
    .X(_00954_));
 sg13g2_mux2_1 _13248_ (.A0(net3407),
    .A1(net4272),
    .S(_05042_),
    .X(_00955_));
 sg13g2_mux2_1 _13249_ (.A0(net3362),
    .A1(net5046),
    .S(_05042_),
    .X(_00956_));
 sg13g2_mux2_1 _13250_ (.A0(net3314),
    .A1(net4328),
    .S(_05042_),
    .X(_00957_));
 sg13g2_mux2_1 _13251_ (.A0(net3266),
    .A1(net4669),
    .S(_05042_),
    .X(_00958_));
 sg13g2_nand3_1 _13252_ (.B(net3087),
    .C(net3026),
    .A(_02244_),
    .Y(_05043_));
 sg13g2_mux2_1 _13253_ (.A0(net3585),
    .A1(net4549),
    .S(_05043_),
    .X(_00959_));
 sg13g2_mux2_1 _13254_ (.A0(net3541),
    .A1(net5126),
    .S(_05043_),
    .X(_00960_));
 sg13g2_mux2_1 _13255_ (.A0(net3498),
    .A1(net4356),
    .S(_05043_),
    .X(_00961_));
 sg13g2_mux2_1 _13256_ (.A0(net3449),
    .A1(net5168),
    .S(_05043_),
    .X(_00962_));
 sg13g2_mux2_1 _13257_ (.A0(net3392),
    .A1(net5163),
    .S(_05043_),
    .X(_00963_));
 sg13g2_mux2_1 _13258_ (.A0(net3360),
    .A1(net4701),
    .S(_05043_),
    .X(_00964_));
 sg13g2_mux2_1 _13259_ (.A0(net3314),
    .A1(net2633),
    .S(_05043_),
    .X(_00965_));
 sg13g2_mux2_1 _13260_ (.A0(net3265),
    .A1(net4332),
    .S(_05043_),
    .X(_00966_));
 sg13g2_nand2_2 _13261_ (.Y(_05044_),
    .A(net3082),
    .B(_02332_));
 sg13g2_mux2_1 _13262_ (.A0(net3589),
    .A1(net4339),
    .S(_05044_),
    .X(_00967_));
 sg13g2_mux2_1 _13263_ (.A0(net3537),
    .A1(net4765),
    .S(_05044_),
    .X(_00968_));
 sg13g2_mux2_1 _13264_ (.A0(net3492),
    .A1(net4629),
    .S(_05044_),
    .X(_00969_));
 sg13g2_mux2_1 _13265_ (.A0(net3445),
    .A1(net4812),
    .S(_05044_),
    .X(_00970_));
 sg13g2_mux2_1 _13266_ (.A0(net3401),
    .A1(net4923),
    .S(_05044_),
    .X(_00971_));
 sg13g2_mux2_1 _13267_ (.A0(net3356),
    .A1(net4793),
    .S(_05044_),
    .X(_00972_));
 sg13g2_mux2_1 _13268_ (.A0(net3311),
    .A1(net4132),
    .S(_05044_),
    .X(_00973_));
 sg13g2_mux2_1 _13269_ (.A0(net3263),
    .A1(net4606),
    .S(_05044_),
    .X(_00974_));
 sg13g2_nand2_1 _13270_ (.Y(_05045_),
    .A(net3084),
    .B(net3024));
 sg13g2_mux2_1 _13271_ (.A0(net3585),
    .A1(net2786),
    .S(net3014),
    .X(_00975_));
 sg13g2_mux2_1 _13272_ (.A0(net3541),
    .A1(net4989),
    .S(_05045_),
    .X(_00976_));
 sg13g2_mux2_1 _13273_ (.A0(net3498),
    .A1(net2856),
    .S(net3014),
    .X(_00977_));
 sg13g2_mux2_1 _13274_ (.A0(net3449),
    .A1(net5135),
    .S(net3014),
    .X(_00978_));
 sg13g2_mux2_1 _13275_ (.A0(net3392),
    .A1(net2872),
    .S(net3014),
    .X(_00979_));
 sg13g2_mux2_1 _13276_ (.A0(net3360),
    .A1(net2870),
    .S(net3014),
    .X(_00980_));
 sg13g2_nor2_1 _13277_ (.A(net3306),
    .B(net3014),
    .Y(_05046_));
 sg13g2_a21oi_1 _13278_ (.A1(_02166_),
    .A2(net3014),
    .Y(_00981_),
    .B1(_05046_));
 sg13g2_mux2_1 _13279_ (.A0(net3264),
    .A1(net2925),
    .S(net3014),
    .X(_00982_));
 sg13g2_and2_2 _13280_ (.A(net3077),
    .B(net3024),
    .X(_05047_));
 sg13g2_mux2_1 _13281_ (.A0(net2697),
    .A1(net3585),
    .S(_05047_),
    .X(_00983_));
 sg13g2_mux2_1 _13282_ (.A0(net2463),
    .A1(net3541),
    .S(_05047_),
    .X(_00984_));
 sg13g2_mux2_1 _13283_ (.A0(net2347),
    .A1(net3498),
    .S(_05047_),
    .X(_00985_));
 sg13g2_mux2_1 _13284_ (.A0(net2734),
    .A1(net3449),
    .S(_05047_),
    .X(_00986_));
 sg13g2_mux2_1 _13285_ (.A0(net2630),
    .A1(net3392),
    .S(_05047_),
    .X(_00987_));
 sg13g2_mux2_1 _13286_ (.A0(net2583),
    .A1(net3359),
    .S(_05047_),
    .X(_00988_));
 sg13g2_mux2_1 _13287_ (.A0(net2346),
    .A1(net3306),
    .S(_05047_),
    .X(_00989_));
 sg13g2_mux2_1 _13288_ (.A0(net2298),
    .A1(net3265),
    .S(_05047_),
    .X(_00990_));
 sg13g2_nand2_2 _13289_ (.Y(_05048_),
    .A(_02283_),
    .B(net3068));
 sg13g2_mux2_1 _13290_ (.A0(net3574),
    .A1(net2647),
    .S(_05048_),
    .X(_00991_));
 sg13g2_mux2_1 _13291_ (.A0(net3525),
    .A1(net4992),
    .S(_05048_),
    .X(_00992_));
 sg13g2_mux2_1 _13292_ (.A0(net3482),
    .A1(net4225),
    .S(_05048_),
    .X(_00993_));
 sg13g2_mux2_1 _13293_ (.A0(net3435),
    .A1(net4583),
    .S(_05048_),
    .X(_00994_));
 sg13g2_mux2_1 _13294_ (.A0(net3390),
    .A1(net2999),
    .S(_05048_),
    .X(_00995_));
 sg13g2_mux2_1 _13295_ (.A0(net3342),
    .A1(net4530),
    .S(_05048_),
    .X(_00996_));
 sg13g2_mux2_1 _13296_ (.A0(net3297),
    .A1(net2997),
    .S(_05048_),
    .X(_00997_));
 sg13g2_mux2_1 _13297_ (.A0(net3249),
    .A1(net4250),
    .S(_05048_),
    .X(_00998_));
 sg13g2_nor2_2 _13298_ (.A(_02298_),
    .B(_02359_),
    .Y(_05049_));
 sg13g2_mux2_1 _13299_ (.A0(net2819),
    .A1(net3574),
    .S(_05049_),
    .X(_00999_));
 sg13g2_mux2_1 _13300_ (.A0(net2239),
    .A1(net3528),
    .S(_05049_),
    .X(_01000_));
 sg13g2_mux2_1 _13301_ (.A0(net2523),
    .A1(net3482),
    .S(_05049_),
    .X(_01001_));
 sg13g2_mux2_1 _13302_ (.A0(net2301),
    .A1(net3435),
    .S(_05049_),
    .X(_01002_));
 sg13g2_mux2_1 _13303_ (.A0(net2383),
    .A1(net3390),
    .S(_05049_),
    .X(_01003_));
 sg13g2_mux2_1 _13304_ (.A0(net2384),
    .A1(net3342),
    .S(_05049_),
    .X(_01004_));
 sg13g2_mux2_1 _13305_ (.A0(net2661),
    .A1(net3297),
    .S(_05049_),
    .X(_01005_));
 sg13g2_mux2_1 _13306_ (.A0(net2512),
    .A1(net3248),
    .S(_05049_),
    .X(_01006_));
 sg13g2_nand2_2 _13307_ (.Y(_05050_),
    .A(net3036),
    .B(net3068));
 sg13g2_mux2_1 _13308_ (.A0(net3574),
    .A1(net2709),
    .S(_05050_),
    .X(_01007_));
 sg13g2_mux2_1 _13309_ (.A0(net3528),
    .A1(net4301),
    .S(_05050_),
    .X(_01008_));
 sg13g2_mux2_1 _13310_ (.A0(net3482),
    .A1(net4220),
    .S(_05050_),
    .X(_01009_));
 sg13g2_mux2_1 _13311_ (.A0(net3435),
    .A1(net4187),
    .S(_05050_),
    .X(_01010_));
 sg13g2_mux2_1 _13312_ (.A0(net3390),
    .A1(net4218),
    .S(_05050_),
    .X(_01011_));
 sg13g2_mux2_1 _13313_ (.A0(net3342),
    .A1(net4056),
    .S(_05050_),
    .X(_01012_));
 sg13g2_mux2_1 _13314_ (.A0(net3297),
    .A1(net4214),
    .S(_05050_),
    .X(_01013_));
 sg13g2_mux2_1 _13315_ (.A0(net3249),
    .A1(net4188),
    .S(_05050_),
    .X(_01014_));
 sg13g2_nand2_2 _13316_ (.Y(_05051_),
    .A(net3033),
    .B(net3067));
 sg13g2_mux2_1 _13317_ (.A0(net3574),
    .A1(net4374),
    .S(_05051_),
    .X(_01015_));
 sg13g2_mux2_1 _13318_ (.A0(net3528),
    .A1(net4539),
    .S(_05051_),
    .X(_01016_));
 sg13g2_mux2_1 _13319_ (.A0(net3482),
    .A1(net4749),
    .S(_05051_),
    .X(_01017_));
 sg13g2_mux2_1 _13320_ (.A0(net3437),
    .A1(net4487),
    .S(_05051_),
    .X(_01018_));
 sg13g2_mux2_1 _13321_ (.A0(net3390),
    .A1(net4422),
    .S(_05051_),
    .X(_01019_));
 sg13g2_mux2_1 _13322_ (.A0(net3342),
    .A1(net4645),
    .S(_05051_),
    .X(_01020_));
 sg13g2_mux2_1 _13323_ (.A0(net3297),
    .A1(net4915),
    .S(_05051_),
    .X(_01021_));
 sg13g2_mux2_1 _13324_ (.A0(net3248),
    .A1(net4192),
    .S(_05051_),
    .X(_01022_));
 sg13g2_nor2_2 _13325_ (.A(net3081),
    .B(_02359_),
    .Y(_05052_));
 sg13g2_mux2_1 _13326_ (.A0(net2228),
    .A1(net3563),
    .S(_05052_),
    .X(_01023_));
 sg13g2_mux2_1 _13327_ (.A0(net2176),
    .A1(net3518),
    .S(_05052_),
    .X(_01024_));
 sg13g2_mux2_1 _13328_ (.A0(net2181),
    .A1(net3481),
    .S(_05052_),
    .X(_01025_));
 sg13g2_mux2_1 _13329_ (.A0(net2747),
    .A1(net3437),
    .S(_05052_),
    .X(_01026_));
 sg13g2_mux2_1 _13330_ (.A0(net2193),
    .A1(net3389),
    .S(_05052_),
    .X(_01027_));
 sg13g2_mux2_1 _13331_ (.A0(net2163),
    .A1(net3334),
    .S(_05052_),
    .X(_01028_));
 sg13g2_mux2_1 _13332_ (.A0(net2172),
    .A1(net3289),
    .S(_05052_),
    .X(_01029_));
 sg13g2_mux2_1 _13333_ (.A0(net2234),
    .A1(net3248),
    .S(_05052_),
    .X(_01030_));
 sg13g2_nand2_2 _13334_ (.Y(_05053_),
    .A(_02346_),
    .B(net3067));
 sg13g2_mux2_1 _13335_ (.A0(net3563),
    .A1(net4711),
    .S(_05053_),
    .X(_01031_));
 sg13g2_mux2_1 _13336_ (.A0(net3518),
    .A1(net4664),
    .S(_05053_),
    .X(_01032_));
 sg13g2_mux2_1 _13337_ (.A0(net3481),
    .A1(net4692),
    .S(_05053_),
    .X(_01033_));
 sg13g2_mux2_1 _13338_ (.A0(net3435),
    .A1(net4489),
    .S(_05053_),
    .X(_01034_));
 sg13g2_mux2_1 _13339_ (.A0(net3389),
    .A1(net4662),
    .S(_05053_),
    .X(_01035_));
 sg13g2_mux2_1 _13340_ (.A0(net3342),
    .A1(net4983),
    .S(_05053_),
    .X(_01036_));
 sg13g2_mux2_1 _13341_ (.A0(net3289),
    .A1(net4167),
    .S(_05053_),
    .X(_01037_));
 sg13g2_mux2_1 _13342_ (.A0(net3248),
    .A1(net4370),
    .S(_05053_),
    .X(_01038_));
 sg13g2_nand2_2 _13343_ (.Y(_05054_),
    .A(net3067),
    .B(_02385_));
 sg13g2_mux2_1 _13344_ (.A0(net3563),
    .A1(net4718),
    .S(_05054_),
    .X(_01039_));
 sg13g2_mux2_1 _13345_ (.A0(net3534),
    .A1(net2928),
    .S(_05054_),
    .X(_01040_));
 sg13g2_mux2_1 _13346_ (.A0(net3481),
    .A1(net4248),
    .S(_05054_),
    .X(_01041_));
 sg13g2_mux2_1 _13347_ (.A0(net3435),
    .A1(net4728),
    .S(_05054_),
    .X(_01042_));
 sg13g2_mux2_1 _13348_ (.A0(net3389),
    .A1(net4243),
    .S(_05054_),
    .X(_01043_));
 sg13g2_mux2_1 _13349_ (.A0(net3342),
    .A1(net4905),
    .S(_05054_),
    .X(_01044_));
 sg13g2_mux2_1 _13350_ (.A0(net3302),
    .A1(net4254),
    .S(_05054_),
    .X(_01045_));
 sg13g2_mux2_1 _13351_ (.A0(net3248),
    .A1(net4698),
    .S(_05054_),
    .X(_01046_));
 sg13g2_nand2_2 _13352_ (.Y(_05055_),
    .A(net3082),
    .B(_02328_));
 sg13g2_mux2_1 _13353_ (.A0(net3582),
    .A1(net5024),
    .S(_05055_),
    .X(_01047_));
 sg13g2_mux2_1 _13354_ (.A0(net3537),
    .A1(net5002),
    .S(_05055_),
    .X(_01048_));
 sg13g2_mux2_1 _13355_ (.A0(net3492),
    .A1(net4431),
    .S(_05055_),
    .X(_01049_));
 sg13g2_mux2_1 _13356_ (.A0(net3445),
    .A1(net4116),
    .S(_05055_),
    .X(_01050_));
 sg13g2_mux2_1 _13357_ (.A0(net3400),
    .A1(net4319),
    .S(_05055_),
    .X(_01051_));
 sg13g2_mux2_1 _13358_ (.A0(net3357),
    .A1(net4238),
    .S(_05055_),
    .X(_01052_));
 sg13g2_mux2_1 _13359_ (.A0(net3311),
    .A1(net4781),
    .S(_05055_),
    .X(_01053_));
 sg13g2_mux2_1 _13360_ (.A0(net3262),
    .A1(net4993),
    .S(_05055_),
    .X(_01054_));
 sg13g2_nor2_2 _13361_ (.A(_02338_),
    .B(_02359_),
    .Y(_05056_));
 sg13g2_mux2_1 _13362_ (.A0(net2571),
    .A1(net3571),
    .S(_05056_),
    .X(_01055_));
 sg13g2_mux2_1 _13363_ (.A0(net2459),
    .A1(net3531),
    .S(_05056_),
    .X(_01056_));
 sg13g2_mux2_1 _13364_ (.A0(net2354),
    .A1(net3484),
    .S(_05056_),
    .X(_01057_));
 sg13g2_mux2_1 _13365_ (.A0(net2568),
    .A1(net3441),
    .S(_05056_),
    .X(_01058_));
 sg13g2_mux2_1 _13366_ (.A0(net2235),
    .A1(net3391),
    .S(_05056_),
    .X(_01059_));
 sg13g2_mux2_1 _13367_ (.A0(net2403),
    .A1(net3348),
    .S(_05056_),
    .X(_01060_));
 sg13g2_mux2_1 _13368_ (.A0(net2603),
    .A1(net3295),
    .S(_05056_),
    .X(_01061_));
 sg13g2_mux2_1 _13369_ (.A0(net2869),
    .A1(net3248),
    .S(_05056_),
    .X(_01062_));
 sg13g2_nor2_2 _13370_ (.A(_02335_),
    .B(_02359_),
    .Y(_05057_));
 sg13g2_mux2_1 _13371_ (.A0(net2554),
    .A1(net3571),
    .S(_05057_),
    .X(_01063_));
 sg13g2_mux2_1 _13372_ (.A0(net2338),
    .A1(net3531),
    .S(_05057_),
    .X(_01064_));
 sg13g2_mux2_1 _13373_ (.A0(net2356),
    .A1(net3484),
    .S(_05057_),
    .X(_01065_));
 sg13g2_mux2_1 _13374_ (.A0(net2381),
    .A1(net3441),
    .S(_05057_),
    .X(_01066_));
 sg13g2_mux2_1 _13375_ (.A0(net2606),
    .A1(net3391),
    .S(_05057_),
    .X(_01067_));
 sg13g2_mux2_1 _13376_ (.A0(net2279),
    .A1(net3348),
    .S(_05057_),
    .X(_01068_));
 sg13g2_mux2_1 _13377_ (.A0(net2490),
    .A1(net3295),
    .S(_05057_),
    .X(_01069_));
 sg13g2_mux2_1 _13378_ (.A0(net2642),
    .A1(net3249),
    .S(_05057_),
    .X(_01070_));
 sg13g2_nand2_2 _13379_ (.Y(_05058_),
    .A(_02332_),
    .B(net3067));
 sg13g2_mux2_1 _13380_ (.A0(net3570),
    .A1(net5081),
    .S(_05058_),
    .X(_01071_));
 sg13g2_mux2_1 _13381_ (.A0(net3531),
    .A1(net4038),
    .S(_05058_),
    .X(_01072_));
 sg13g2_mux2_1 _13382_ (.A0(net3484),
    .A1(net2899),
    .S(_05058_),
    .X(_01073_));
 sg13g2_mux2_1 _13383_ (.A0(net3441),
    .A1(net4895),
    .S(_05058_),
    .X(_01074_));
 sg13g2_mux2_1 _13384_ (.A0(net3391),
    .A1(net4279),
    .S(_05058_),
    .X(_01075_));
 sg13g2_mux2_1 _13385_ (.A0(net3348),
    .A1(net4437),
    .S(_05058_),
    .X(_01076_));
 sg13g2_mux2_1 _13386_ (.A0(net3295),
    .A1(net4273),
    .S(_05058_),
    .X(_01077_));
 sg13g2_mux2_1 _13387_ (.A0(net3248),
    .A1(net5160),
    .S(_05058_),
    .X(_01078_));
 sg13g2_nand2_2 _13388_ (.Y(_05059_),
    .A(_02328_),
    .B(net3067));
 sg13g2_mux2_1 _13389_ (.A0(net3570),
    .A1(net4927),
    .S(_05059_),
    .X(_01079_));
 sg13g2_mux2_1 _13390_ (.A0(net3531),
    .A1(net4910),
    .S(_05059_),
    .X(_01080_));
 sg13g2_mux2_1 _13391_ (.A0(net3484),
    .A1(net2998),
    .S(_05059_),
    .X(_01081_));
 sg13g2_mux2_1 _13392_ (.A0(net3441),
    .A1(net4807),
    .S(_05059_),
    .X(_01082_));
 sg13g2_mux2_1 _13393_ (.A0(net3391),
    .A1(net4971),
    .S(_05059_),
    .X(_01083_));
 sg13g2_mux2_1 _13394_ (.A0(net3348),
    .A1(net4049),
    .S(_05059_),
    .X(_01084_));
 sg13g2_mux2_1 _13395_ (.A0(net3295),
    .A1(net4050),
    .S(_05059_),
    .X(_01085_));
 sg13g2_mux2_1 _13396_ (.A0(net3249),
    .A1(net4227),
    .S(_05059_),
    .X(_01086_));
 sg13g2_nand2_2 _13397_ (.Y(_05060_),
    .A(net3072),
    .B(net3067));
 sg13g2_mux2_1 _13398_ (.A0(net3578),
    .A1(net2827),
    .S(_05060_),
    .X(_01087_));
 sg13g2_mux2_1 _13399_ (.A0(net3531),
    .A1(net5117),
    .S(_05060_),
    .X(_01088_));
 sg13g2_mux2_1 _13400_ (.A0(net3485),
    .A1(net4362),
    .S(_05060_),
    .X(_01089_));
 sg13g2_mux2_1 _13401_ (.A0(net3438),
    .A1(net5078),
    .S(_05060_),
    .X(_01090_));
 sg13g2_mux2_1 _13402_ (.A0(net3391),
    .A1(net4713),
    .S(_05060_),
    .X(_01091_));
 sg13g2_mux2_1 _13403_ (.A0(net3348),
    .A1(net2824),
    .S(_05060_),
    .X(_01092_));
 sg13g2_mux2_1 _13404_ (.A0(net3303),
    .A1(net4256),
    .S(_05060_),
    .X(_01093_));
 sg13g2_mux2_1 _13405_ (.A0(net3249),
    .A1(net5058),
    .S(_05060_),
    .X(_01094_));
 sg13g2_nand3_1 _13406_ (.B(net3073),
    .C(net3067),
    .A(net3042),
    .Y(_05061_));
 sg13g2_mux2_1 _13407_ (.A0(net3578),
    .A1(net5148),
    .S(_05061_),
    .X(_01095_));
 sg13g2_mux2_1 _13408_ (.A0(net3528),
    .A1(net4562),
    .S(_05061_),
    .X(_01096_));
 sg13g2_mux2_1 _13409_ (.A0(net3485),
    .A1(net4402),
    .S(_05061_),
    .X(_01097_));
 sg13g2_mux2_1 _13410_ (.A0(net3438),
    .A1(net4799),
    .S(_05061_),
    .X(_01098_));
 sg13g2_mux2_1 _13411_ (.A0(net3391),
    .A1(net4550),
    .S(_05061_),
    .X(_01099_));
 sg13g2_mux2_1 _13412_ (.A0(net3349),
    .A1(net5179),
    .S(_05061_),
    .X(_01100_));
 sg13g2_mux2_1 _13413_ (.A0(net3303),
    .A1(net4198),
    .S(_05061_),
    .X(_01101_));
 sg13g2_mux2_1 _13414_ (.A0(net3249),
    .A1(net4967),
    .S(_05061_),
    .X(_01102_));
 sg13g2_nand3_1 _13415_ (.B(net3042),
    .C(net3068),
    .A(net3084),
    .Y(_05062_));
 sg13g2_mux2_1 _13416_ (.A0(net3578),
    .A1(net2750),
    .S(_05062_),
    .X(_01103_));
 sg13g2_mux2_1 _13417_ (.A0(net3531),
    .A1(net4635),
    .S(_05062_),
    .X(_01104_));
 sg13g2_mux2_1 _13418_ (.A0(net3485),
    .A1(net4628),
    .S(_05062_),
    .X(_01105_));
 sg13g2_mux2_1 _13419_ (.A0(net3438),
    .A1(net4721),
    .S(_05062_),
    .X(_01106_));
 sg13g2_mux2_1 _13420_ (.A0(net3391),
    .A1(net4756),
    .S(_05062_),
    .X(_01107_));
 sg13g2_mux2_1 _13421_ (.A0(net3348),
    .A1(net4786),
    .S(_05062_),
    .X(_01108_));
 sg13g2_mux2_1 _13422_ (.A0(net3303),
    .A1(net3007),
    .S(_05062_),
    .X(_01109_));
 sg13g2_mux2_1 _13423_ (.A0(net3256),
    .A1(net4674),
    .S(_05062_),
    .X(_01110_));
 sg13g2_nor2_2 _13424_ (.A(net3039),
    .B(_02477_),
    .Y(_05063_));
 sg13g2_mux2_1 _13425_ (.A0(net2808),
    .A1(net3578),
    .S(_05063_),
    .X(_01111_));
 sg13g2_mux2_1 _13426_ (.A0(net2302),
    .A1(net3532),
    .S(_05063_),
    .X(_01112_));
 sg13g2_mux2_1 _13427_ (.A0(net2336),
    .A1(net3485),
    .S(_05063_),
    .X(_01113_));
 sg13g2_mux2_1 _13428_ (.A0(net2607),
    .A1(net3438),
    .S(_05063_),
    .X(_01114_));
 sg13g2_mux2_1 _13429_ (.A0(net2417),
    .A1(net3391),
    .S(_05063_),
    .X(_01115_));
 sg13g2_mux2_1 _13430_ (.A0(net2499),
    .A1(net3348),
    .S(_05063_),
    .X(_01116_));
 sg13g2_mux2_1 _13431_ (.A0(net2365),
    .A1(net3303),
    .S(_05063_),
    .X(_01117_));
 sg13g2_mux2_1 _13432_ (.A0(net2429),
    .A1(net3256),
    .S(_05063_),
    .X(_01118_));
 sg13g2_nand2_2 _13433_ (.Y(_05064_),
    .A(net3080),
    .B(_02370_));
 sg13g2_mux2_1 _13434_ (.A0(net3584),
    .A1(net4477),
    .S(_05064_),
    .X(_01119_));
 sg13g2_mux2_1 _13435_ (.A0(net3542),
    .A1(net4822),
    .S(_05064_),
    .X(_01120_));
 sg13g2_mux2_1 _13436_ (.A0(net3492),
    .A1(net4580),
    .S(_05064_),
    .X(_01121_));
 sg13g2_mux2_1 _13437_ (.A0(net3446),
    .A1(net4829),
    .S(_05064_),
    .X(_01122_));
 sg13g2_mux2_1 _13438_ (.A0(net3405),
    .A1(net4672),
    .S(_05064_),
    .X(_01123_));
 sg13g2_mux2_1 _13439_ (.A0(net3356),
    .A1(net2831),
    .S(_05064_),
    .X(_01124_));
 sg13g2_mux2_1 _13440_ (.A0(net3311),
    .A1(net4037),
    .S(_05064_),
    .X(_01125_));
 sg13g2_mux2_1 _13441_ (.A0(net3261),
    .A1(net4704),
    .S(_05064_),
    .X(_01126_));
 sg13g2_nand2_2 _13442_ (.Y(_05065_),
    .A(net3082),
    .B(_02321_));
 sg13g2_mux2_1 _13443_ (.A0(net3590),
    .A1(net4544),
    .S(_05065_),
    .X(_01127_));
 sg13g2_mux2_1 _13444_ (.A0(net3536),
    .A1(net4346),
    .S(_05065_),
    .X(_01128_));
 sg13g2_mux2_1 _13445_ (.A0(net3500),
    .A1(net4916),
    .S(_05065_),
    .X(_01129_));
 sg13g2_mux2_1 _13446_ (.A0(net3454),
    .A1(net4820),
    .S(_05065_),
    .X(_01130_));
 sg13g2_mux2_1 _13447_ (.A0(net3408),
    .A1(net2794),
    .S(_05065_),
    .X(_01131_));
 sg13g2_mux2_1 _13448_ (.A0(net3365),
    .A1(net2730),
    .S(_05065_),
    .X(_01132_));
 sg13g2_mux2_1 _13449_ (.A0(net3310),
    .A1(net2844),
    .S(_05065_),
    .X(_01133_));
 sg13g2_mux2_1 _13450_ (.A0(net3269),
    .A1(net4178),
    .S(_05065_),
    .X(_01134_));
 sg13g2_nor2_2 _13451_ (.A(_02289_),
    .B(_02371_),
    .Y(_05066_));
 sg13g2_mux2_1 _13452_ (.A0(net2529),
    .A1(net3586),
    .S(_05066_),
    .X(_01135_));
 sg13g2_mux2_1 _13453_ (.A0(net2479),
    .A1(net3542),
    .S(_05066_),
    .X(_01136_));
 sg13g2_mux2_1 _13454_ (.A0(net2753),
    .A1(net3492),
    .S(_05066_),
    .X(_01137_));
 sg13g2_mux2_1 _13455_ (.A0(net2487),
    .A1(net3448),
    .S(_05066_),
    .X(_01138_));
 sg13g2_mux2_1 _13456_ (.A0(net2605),
    .A1(net3405),
    .S(_05066_),
    .X(_01139_));
 sg13g2_mux2_1 _13457_ (.A0(net2157),
    .A1(net3357),
    .S(_05066_),
    .X(_01140_));
 sg13g2_mux2_1 _13458_ (.A0(net2449),
    .A1(net3311),
    .S(_05066_),
    .X(_01141_));
 sg13g2_mux2_1 _13459_ (.A0(net2330),
    .A1(net3261),
    .S(_05066_),
    .X(_01142_));
 sg13g2_and2_2 _13460_ (.A(_02349_),
    .B(_02370_),
    .X(_05067_));
 sg13g2_mux2_1 _13461_ (.A0(net2663),
    .A1(net3586),
    .S(_05067_),
    .X(_01143_));
 sg13g2_mux2_1 _13462_ (.A0(net2522),
    .A1(net3537),
    .S(_05067_),
    .X(_01144_));
 sg13g2_mux2_1 _13463_ (.A0(net2362),
    .A1(net3492),
    .S(_05067_),
    .X(_01145_));
 sg13g2_mux2_1 _13464_ (.A0(net2278),
    .A1(net3450),
    .S(_05067_),
    .X(_01146_));
 sg13g2_mux2_1 _13465_ (.A0(net2430),
    .A1(net3405),
    .S(_05067_),
    .X(_01147_));
 sg13g2_mux2_1 _13466_ (.A0(net2638),
    .A1(net3357),
    .S(_05067_),
    .X(_01148_));
 sg13g2_mux2_1 _13467_ (.A0(net2258),
    .A1(net3311),
    .S(_05067_),
    .X(_01149_));
 sg13g2_mux2_1 _13468_ (.A0(net2311),
    .A1(net3261),
    .S(_05067_),
    .X(_01150_));
 sg13g2_nor2_2 _13469_ (.A(net3081),
    .B(_02371_),
    .Y(_05068_));
 sg13g2_mux2_1 _13470_ (.A0(net2218),
    .A1(net3587),
    .S(_05068_),
    .X(_01151_));
 sg13g2_mux2_1 _13471_ (.A0(net2400),
    .A1(net3537),
    .S(_05068_),
    .X(_01152_));
 sg13g2_mux2_1 _13472_ (.A0(net2427),
    .A1(net3494),
    .S(_05068_),
    .X(_01153_));
 sg13g2_mux2_1 _13473_ (.A0(net2355),
    .A1(net3452),
    .S(_05068_),
    .X(_01154_));
 sg13g2_mux2_1 _13474_ (.A0(net2247),
    .A1(net3406),
    .S(_05068_),
    .X(_01155_));
 sg13g2_mux2_1 _13475_ (.A0(net2146),
    .A1(net3357),
    .S(_05068_),
    .X(_01156_));
 sg13g2_mux2_1 _13476_ (.A0(net2445),
    .A1(net3311),
    .S(_05068_),
    .X(_01157_));
 sg13g2_mux2_1 _13477_ (.A0(net2169),
    .A1(net3261),
    .S(_05068_),
    .X(_01158_));
 sg13g2_and2_2 _13478_ (.A(net3069),
    .B(_02370_),
    .X(_05069_));
 sg13g2_mux2_1 _13479_ (.A0(net2749),
    .A1(net3587),
    .S(_05069_),
    .X(_01159_));
 sg13g2_mux2_1 _13480_ (.A0(net2214),
    .A1(net3537),
    .S(_05069_),
    .X(_01160_));
 sg13g2_mux2_1 _13481_ (.A0(net2670),
    .A1(net3500),
    .S(_05069_),
    .X(_01161_));
 sg13g2_mux2_1 _13482_ (.A0(net2416),
    .A1(net3450),
    .S(_05069_),
    .X(_01162_));
 sg13g2_mux2_1 _13483_ (.A0(net2516),
    .A1(net3413),
    .S(_05069_),
    .X(_01163_));
 sg13g2_mux2_1 _13484_ (.A0(net2669),
    .A1(net3356),
    .S(_05069_),
    .X(_01164_));
 sg13g2_mux2_1 _13485_ (.A0(net2313),
    .A1(net3319),
    .S(_05069_),
    .X(_01165_));
 sg13g2_mux2_1 _13486_ (.A0(net2335),
    .A1(net3263),
    .S(_05069_),
    .X(_01166_));
 sg13g2_and2_2 _13487_ (.A(_02370_),
    .B(net3065),
    .X(_05070_));
 sg13g2_mux2_1 _13488_ (.A0(net2312),
    .A1(net3586),
    .S(_05070_),
    .X(_01167_));
 sg13g2_mux2_1 _13489_ (.A0(net2513),
    .A1(net3538),
    .S(_05070_),
    .X(_01168_));
 sg13g2_mux2_1 _13490_ (.A0(net2382),
    .A1(net3500),
    .S(_05070_),
    .X(_01169_));
 sg13g2_mux2_1 _13491_ (.A0(net2357),
    .A1(net3450),
    .S(_05070_),
    .X(_01170_));
 sg13g2_mux2_1 _13492_ (.A0(net2401),
    .A1(net3413),
    .S(_05070_),
    .X(_01171_));
 sg13g2_mux2_1 _13493_ (.A0(net2139),
    .A1(net3356),
    .S(_05070_),
    .X(_01172_));
 sg13g2_mux2_1 _13494_ (.A0(net2352),
    .A1(net3319),
    .S(_05070_),
    .X(_01173_));
 sg13g2_mux2_1 _13495_ (.A0(net2587),
    .A1(net3261),
    .S(_05070_),
    .X(_01174_));
 sg13g2_nand2_2 _13496_ (.Y(_05071_),
    .A(_02309_),
    .B(_02370_));
 sg13g2_mux2_1 _13497_ (.A0(net3586),
    .A1(net2906),
    .S(_05071_),
    .X(_01175_));
 sg13g2_mux2_1 _13498_ (.A0(net3537),
    .A1(net4304),
    .S(_05071_),
    .X(_01176_));
 sg13g2_mux2_1 _13499_ (.A0(net3500),
    .A1(net4119),
    .S(_05071_),
    .X(_01177_));
 sg13g2_mux2_1 _13500_ (.A0(net3450),
    .A1(net5103),
    .S(_05071_),
    .X(_01178_));
 sg13g2_mux2_1 _13501_ (.A0(net3413),
    .A1(net4772),
    .S(_05071_),
    .X(_01179_));
 sg13g2_mux2_1 _13502_ (.A0(net3356),
    .A1(net4963),
    .S(_05071_),
    .X(_01180_));
 sg13g2_mux2_1 _13503_ (.A0(net3319),
    .A1(net4302),
    .S(_05071_),
    .X(_01181_));
 sg13g2_mux2_1 _13504_ (.A0(net3261),
    .A1(net4165),
    .S(_05071_),
    .X(_01182_));
 sg13g2_nor2_2 _13505_ (.A(_02338_),
    .B(_02371_),
    .Y(_05072_));
 sg13g2_mux2_1 _13506_ (.A0(net2274),
    .A1(net3584),
    .S(_05072_),
    .X(_01183_));
 sg13g2_mux2_1 _13507_ (.A0(net2212),
    .A1(net3540),
    .S(_05072_),
    .X(_01184_));
 sg13g2_mux2_1 _13508_ (.A0(net2190),
    .A1(net3498),
    .S(_05072_),
    .X(_01185_));
 sg13g2_mux2_1 _13509_ (.A0(net2195),
    .A1(net3447),
    .S(_05072_),
    .X(_01186_));
 sg13g2_mux2_1 _13510_ (.A0(net2284),
    .A1(net3403),
    .S(_05072_),
    .X(_01187_));
 sg13g2_mux2_1 _13511_ (.A0(net2549),
    .A1(net3359),
    .S(_05072_),
    .X(_01188_));
 sg13g2_mux2_1 _13512_ (.A0(net2646),
    .A1(net3315),
    .S(_05072_),
    .X(_01189_));
 sg13g2_mux2_1 _13513_ (.A0(net2751),
    .A1(net3264),
    .S(_05072_),
    .X(_01190_));
 sg13g2_nor2_2 _13514_ (.A(_02335_),
    .B(_02371_),
    .Y(_05073_));
 sg13g2_mux2_1 _13515_ (.A0(net2424),
    .A1(net3584),
    .S(_05073_),
    .X(_01191_));
 sg13g2_mux2_1 _13516_ (.A0(net2388),
    .A1(net3540),
    .S(_05073_),
    .X(_01192_));
 sg13g2_mux2_1 _13517_ (.A0(net2310),
    .A1(net3498),
    .S(_05073_),
    .X(_01193_));
 sg13g2_mux2_1 _13518_ (.A0(net2654),
    .A1(net3447),
    .S(_05073_),
    .X(_01194_));
 sg13g2_mux2_1 _13519_ (.A0(net2526),
    .A1(net3403),
    .S(_05073_),
    .X(_01195_));
 sg13g2_mux2_1 _13520_ (.A0(net2545),
    .A1(net3359),
    .S(_05073_),
    .X(_01196_));
 sg13g2_mux2_1 _13521_ (.A0(net2343),
    .A1(net3315),
    .S(_05073_),
    .X(_01197_));
 sg13g2_mux2_1 _13522_ (.A0(net2737),
    .A1(net3264),
    .S(_05073_),
    .X(_01198_));
 sg13g2_nor2_2 _13523_ (.A(_02331_),
    .B(_02371_),
    .Y(_05074_));
 sg13g2_mux2_1 _13524_ (.A0(net2254),
    .A1(net3584),
    .S(_05074_),
    .X(_01199_));
 sg13g2_mux2_1 _13525_ (.A0(net2281),
    .A1(net3540),
    .S(_05074_),
    .X(_01200_));
 sg13g2_mux2_1 _13526_ (.A0(net2473),
    .A1(net3498),
    .S(_05074_),
    .X(_01201_));
 sg13g2_mux2_1 _13527_ (.A0(net2577),
    .A1(net3447),
    .S(_05074_),
    .X(_01202_));
 sg13g2_mux2_1 _13528_ (.A0(net2432),
    .A1(net3403),
    .S(_05074_),
    .X(_01203_));
 sg13g2_mux2_1 _13529_ (.A0(net2341),
    .A1(net3359),
    .S(_05074_),
    .X(_01204_));
 sg13g2_mux2_1 _13530_ (.A0(net2548),
    .A1(net3315),
    .S(_05074_),
    .X(_01205_));
 sg13g2_mux2_1 _13531_ (.A0(net2438),
    .A1(net3264),
    .S(_05074_),
    .X(_01206_));
 sg13g2_nand2_2 _13532_ (.Y(_05075_),
    .A(_02311_),
    .B(net3074));
 sg13g2_mux2_1 _13533_ (.A0(net3590),
    .A1(net4312),
    .S(_05075_),
    .X(_01207_));
 sg13g2_mux2_1 _13534_ (.A0(net3536),
    .A1(net4128),
    .S(_05075_),
    .X(_01208_));
 sg13g2_mux2_1 _13535_ (.A0(net3499),
    .A1(net5183),
    .S(_05075_),
    .X(_01209_));
 sg13g2_mux2_1 _13536_ (.A0(net3454),
    .A1(net4691),
    .S(_05075_),
    .X(_01210_));
 sg13g2_mux2_1 _13537_ (.A0(net3408),
    .A1(net4885),
    .S(_05075_),
    .X(_01211_));
 sg13g2_mux2_1 _13538_ (.A0(net3365),
    .A1(net5109),
    .S(_05075_),
    .X(_01212_));
 sg13g2_mux2_1 _13539_ (.A0(net3310),
    .A1(net4994),
    .S(_05075_),
    .X(_01213_));
 sg13g2_mux2_1 _13540_ (.A0(net3269),
    .A1(net4734),
    .S(_05075_),
    .X(_01214_));
 sg13g2_nor2_2 _13541_ (.A(_02322_),
    .B(_02369_),
    .Y(_05076_));
 sg13g2_mux2_1 _13542_ (.A0(net2178),
    .A1(net3586),
    .S(_05076_),
    .X(_01215_));
 sg13g2_mux2_1 _13543_ (.A0(net2612),
    .A1(net3542),
    .S(_05076_),
    .X(_01216_));
 sg13g2_mux2_1 _13544_ (.A0(net2506),
    .A1(net3497),
    .S(_05076_),
    .X(_01217_));
 sg13g2_mux2_1 _13545_ (.A0(net2530),
    .A1(net3450),
    .S(_05076_),
    .X(_01218_));
 sg13g2_mux2_1 _13546_ (.A0(net2186),
    .A1(net3406),
    .S(_05076_),
    .X(_01219_));
 sg13g2_mux2_1 _13547_ (.A0(net2134),
    .A1(net3363),
    .S(_05076_),
    .X(_01220_));
 sg13g2_mux2_1 _13548_ (.A0(net2287),
    .A1(net3316),
    .S(_05076_),
    .X(_01221_));
 sg13g2_mux2_1 _13549_ (.A0(net2564),
    .A1(net3266),
    .S(_05076_),
    .X(_01222_));
 sg13g2_nand2_2 _13550_ (.Y(_05077_),
    .A(net3074),
    .B(_02370_));
 sg13g2_mux2_1 _13551_ (.A0(net3586),
    .A1(net4642),
    .S(_05077_),
    .X(_01223_));
 sg13g2_mux2_1 _13552_ (.A0(net3542),
    .A1(net4275),
    .S(_05077_),
    .X(_01224_));
 sg13g2_mux2_1 _13553_ (.A0(net3497),
    .A1(net4508),
    .S(_05077_),
    .X(_01225_));
 sg13g2_mux2_1 _13554_ (.A0(net3450),
    .A1(net4649),
    .S(_05077_),
    .X(_01226_));
 sg13g2_mux2_1 _13555_ (.A0(net3406),
    .A1(net4204),
    .S(_05077_),
    .X(_01227_));
 sg13g2_mux2_1 _13556_ (.A0(net3363),
    .A1(net4382),
    .S(_05077_),
    .X(_01228_));
 sg13g2_mux2_1 _13557_ (.A0(net3316),
    .A1(net4263),
    .S(_05077_),
    .X(_01229_));
 sg13g2_mux2_1 _13558_ (.A0(net3266),
    .A1(net4504),
    .S(_05077_),
    .X(_01230_));
 sg13g2_nand2_2 _13559_ (.Y(_05078_),
    .A(net3085),
    .B(_02370_));
 sg13g2_mux2_1 _13560_ (.A0(net3586),
    .A1(net4021),
    .S(_05078_),
    .X(_01231_));
 sg13g2_mux2_1 _13561_ (.A0(net3542),
    .A1(net3004),
    .S(_05078_),
    .X(_01232_));
 sg13g2_mux2_1 _13562_ (.A0(net3497),
    .A1(net4630),
    .S(_05078_),
    .X(_01233_));
 sg13g2_mux2_1 _13563_ (.A0(net3450),
    .A1(net2880),
    .S(_05078_),
    .X(_01234_));
 sg13g2_mux2_1 _13564_ (.A0(net3406),
    .A1(net3000),
    .S(_05078_),
    .X(_01235_));
 sg13g2_mux2_1 _13565_ (.A0(net3363),
    .A1(net2850),
    .S(_05078_),
    .X(_01236_));
 sg13g2_mux2_1 _13566_ (.A0(net3316),
    .A1(net2849),
    .S(_05078_),
    .X(_01237_));
 sg13g2_mux2_1 _13567_ (.A0(net3266),
    .A1(net4209),
    .S(_05078_),
    .X(_01238_));
 sg13g2_nor2_2 _13568_ (.A(_02307_),
    .B(_02371_),
    .Y(_05079_));
 sg13g2_mux2_1 _13569_ (.A0(net2405),
    .A1(net3586),
    .S(_05079_),
    .X(_01239_));
 sg13g2_mux2_1 _13570_ (.A0(net2376),
    .A1(net3542),
    .S(_05079_),
    .X(_01240_));
 sg13g2_mux2_1 _13571_ (.A0(net2249),
    .A1(net3497),
    .S(_05079_),
    .X(_01241_));
 sg13g2_mux2_1 _13572_ (.A0(net2515),
    .A1(net3450),
    .S(_05079_),
    .X(_01242_));
 sg13g2_mux2_1 _13573_ (.A0(net2360),
    .A1(net3406),
    .S(_05079_),
    .X(_01243_));
 sg13g2_mux2_1 _13574_ (.A0(net2550),
    .A1(net3363),
    .S(_05079_),
    .X(_01244_));
 sg13g2_mux2_1 _13575_ (.A0(net2769),
    .A1(net3316),
    .S(_05079_),
    .X(_01245_));
 sg13g2_mux2_1 _13576_ (.A0(net2372),
    .A1(net3266),
    .S(_05079_),
    .X(_01246_));
 sg13g2_and2_2 _13577_ (.A(net3080),
    .B(net3027),
    .X(_05080_));
 sg13g2_mux2_1 _13578_ (.A0(net2502),
    .A1(net3596),
    .S(_05080_),
    .X(_01247_));
 sg13g2_mux2_1 _13579_ (.A0(net2685),
    .A1(net3551),
    .S(_05080_),
    .X(_01248_));
 sg13g2_mux2_1 _13580_ (.A0(net2170),
    .A1(net3504),
    .S(_05080_),
    .X(_01249_));
 sg13g2_mux2_1 _13581_ (.A0(net2216),
    .A1(net3460),
    .S(_05080_),
    .X(_01250_));
 sg13g2_mux2_1 _13582_ (.A0(net2689),
    .A1(net3414),
    .S(_05080_),
    .X(_01251_));
 sg13g2_mux2_1 _13583_ (.A0(net2493),
    .A1(net3370),
    .S(_05080_),
    .X(_01252_));
 sg13g2_mux2_1 _13584_ (.A0(net2676),
    .A1(net3317),
    .S(_05080_),
    .X(_01253_));
 sg13g2_mux2_1 _13585_ (.A0(net2691),
    .A1(net3276),
    .S(_05080_),
    .X(_01254_));
 sg13g2_nand2_2 _13586_ (.Y(_05081_),
    .A(_02297_),
    .B(net3027));
 sg13g2_mux2_1 _13587_ (.A0(net3596),
    .A1(net4517),
    .S(_05081_),
    .X(_01255_));
 sg13g2_mux2_1 _13588_ (.A0(net3551),
    .A1(net4149),
    .S(_05081_),
    .X(_01256_));
 sg13g2_mux2_1 _13589_ (.A0(net3504),
    .A1(net4259),
    .S(_05081_),
    .X(_01257_));
 sg13g2_mux2_1 _13590_ (.A0(net3460),
    .A1(net4264),
    .S(_05081_),
    .X(_01258_));
 sg13g2_mux2_1 _13591_ (.A0(net3414),
    .A1(net4594),
    .S(_05081_),
    .X(_01259_));
 sg13g2_mux2_1 _13592_ (.A0(net3370),
    .A1(net4247),
    .S(_05081_),
    .X(_01260_));
 sg13g2_mux2_1 _13593_ (.A0(net3317),
    .A1(net4506),
    .S(_05081_),
    .X(_01261_));
 sg13g2_mux2_1 _13594_ (.A0(net3276),
    .A1(net4492),
    .S(_05081_),
    .X(_01262_));
 sg13g2_nand2_2 _13595_ (.Y(_05082_),
    .A(net3036),
    .B(_02365_));
 sg13g2_mux2_1 _13596_ (.A0(net3596),
    .A1(net4610),
    .S(_05082_),
    .X(_01263_));
 sg13g2_mux2_1 _13597_ (.A0(net3551),
    .A1(net4747),
    .S(_05082_),
    .X(_01264_));
 sg13g2_mux2_1 _13598_ (.A0(net3504),
    .A1(net4670),
    .S(_05082_),
    .X(_01265_));
 sg13g2_mux2_1 _13599_ (.A0(net3460),
    .A1(net4828),
    .S(_05082_),
    .X(_01266_));
 sg13g2_mux2_1 _13600_ (.A0(net3414),
    .A1(net4696),
    .S(_05082_),
    .X(_01267_));
 sg13g2_mux2_1 _13601_ (.A0(net3370),
    .A1(net5069),
    .S(_05082_),
    .X(_01268_));
 sg13g2_mux2_1 _13602_ (.A0(net3317),
    .A1(net4114),
    .S(_05082_),
    .X(_01269_));
 sg13g2_mux2_1 _13603_ (.A0(net3276),
    .A1(net4079),
    .S(_05082_),
    .X(_01270_));
 sg13g2_nand2_2 _13604_ (.Y(_05083_),
    .A(net3033),
    .B(_02365_));
 sg13g2_mux2_1 _13605_ (.A0(net3596),
    .A1(net5101),
    .S(_05083_),
    .X(_01271_));
 sg13g2_mux2_1 _13606_ (.A0(net3552),
    .A1(net4763),
    .S(_05083_),
    .X(_01272_));
 sg13g2_mux2_1 _13607_ (.A0(net3504),
    .A1(net4616),
    .S(_05083_),
    .X(_01273_));
 sg13g2_mux2_1 _13608_ (.A0(net3460),
    .A1(net4541),
    .S(_05083_),
    .X(_01274_));
 sg13g2_mux2_1 _13609_ (.A0(net3414),
    .A1(net5031),
    .S(_05083_),
    .X(_01275_));
 sg13g2_mux2_1 _13610_ (.A0(net3370),
    .A1(net4197),
    .S(_05083_),
    .X(_01276_));
 sg13g2_mux2_1 _13611_ (.A0(net3317),
    .A1(net4957),
    .S(_05083_),
    .X(_01277_));
 sg13g2_mux2_1 _13612_ (.A0(net3276),
    .A1(net5061),
    .S(_05083_),
    .X(_01278_));
 sg13g2_nand2_2 _13613_ (.Y(_05084_),
    .A(_02277_),
    .B(net3028));
 sg13g2_mux2_1 _13614_ (.A0(net3598),
    .A1(net4298),
    .S(_05084_),
    .X(_01279_));
 sg13g2_mux2_1 _13615_ (.A0(net3553),
    .A1(net4083),
    .S(_05084_),
    .X(_01280_));
 sg13g2_mux2_1 _13616_ (.A0(net3508),
    .A1(net2955),
    .S(_05084_),
    .X(_01281_));
 sg13g2_mux2_1 _13617_ (.A0(net3463),
    .A1(net4016),
    .S(_05084_),
    .X(_01282_));
 sg13g2_mux2_1 _13618_ (.A0(net3414),
    .A1(net4796),
    .S(_05084_),
    .X(_01283_));
 sg13g2_mux2_1 _13619_ (.A0(net3372),
    .A1(net4693),
    .S(_05084_),
    .X(_01284_));
 sg13g2_mux2_1 _13620_ (.A0(net3326),
    .A1(net2684),
    .S(_05084_),
    .X(_01285_));
 sg13g2_mux2_1 _13621_ (.A0(net3279),
    .A1(net2929),
    .S(_05084_),
    .X(_01286_));
 sg13g2_nand2_2 _13622_ (.Y(_05085_),
    .A(net3085),
    .B(_02311_));
 sg13g2_mux2_1 _13623_ (.A0(net3591),
    .A1(net2762),
    .S(_05085_),
    .X(_01287_));
 sg13g2_mux2_1 _13624_ (.A0(net3538),
    .A1(net2947),
    .S(_05085_),
    .X(_01288_));
 sg13g2_mux2_1 _13625_ (.A0(net3493),
    .A1(net4815),
    .S(_05085_),
    .X(_01289_));
 sg13g2_mux2_1 _13626_ (.A0(net3455),
    .A1(net4683),
    .S(_05085_),
    .X(_01290_));
 sg13g2_mux2_1 _13627_ (.A0(net3409),
    .A1(net2790),
    .S(_05085_),
    .X(_01291_));
 sg13g2_mux2_1 _13628_ (.A0(net3365),
    .A1(net4520),
    .S(_05085_),
    .X(_01292_));
 sg13g2_mux2_1 _13629_ (.A0(net3312),
    .A1(net2842),
    .S(_05085_),
    .X(_01293_));
 sg13g2_mux2_1 _13630_ (.A0(net3270),
    .A1(net4232),
    .S(_05085_),
    .X(_01294_));
 sg13g2_nand2_2 _13631_ (.Y(_05086_),
    .A(net3028),
    .B(net3065));
 sg13g2_mux2_1 _13632_ (.A0(net3596),
    .A1(net2975),
    .S(_05086_),
    .X(_01295_));
 sg13g2_mux2_1 _13633_ (.A0(net3552),
    .A1(net5142),
    .S(_05086_),
    .X(_01296_));
 sg13g2_mux2_1 _13634_ (.A0(net3508),
    .A1(net5021),
    .S(_05086_),
    .X(_01297_));
 sg13g2_mux2_1 _13635_ (.A0(net3461),
    .A1(net4538),
    .S(_05086_),
    .X(_01298_));
 sg13g2_mux2_1 _13636_ (.A0(net3414),
    .A1(net2908),
    .S(_05086_),
    .X(_01299_));
 sg13g2_mux2_1 _13637_ (.A0(net3370),
    .A1(net2726),
    .S(_05086_),
    .X(_01300_));
 sg13g2_mux2_1 _13638_ (.A0(net3324),
    .A1(net4135),
    .S(_05086_),
    .X(_01301_));
 sg13g2_mux2_1 _13639_ (.A0(net3278),
    .A1(net4072),
    .S(_05086_),
    .X(_01302_));
 sg13g2_nand2_2 _13640_ (.Y(_05087_),
    .A(net3049),
    .B(_02365_));
 sg13g2_mux2_1 _13641_ (.A0(net3596),
    .A1(net4835),
    .S(_05087_),
    .X(_01303_));
 sg13g2_mux2_1 _13642_ (.A0(net3551),
    .A1(net2912),
    .S(_05087_),
    .X(_01304_));
 sg13g2_mux2_1 _13643_ (.A0(net3508),
    .A1(net4447),
    .S(_05087_),
    .X(_01305_));
 sg13g2_mux2_1 _13644_ (.A0(net3461),
    .A1(net4379),
    .S(_05087_),
    .X(_01306_));
 sg13g2_mux2_1 _13645_ (.A0(net3414),
    .A1(net4034),
    .S(_05087_),
    .X(_01307_));
 sg13g2_mux2_1 _13646_ (.A0(net3370),
    .A1(net4647),
    .S(_05087_),
    .X(_01308_));
 sg13g2_mux2_1 _13647_ (.A0(net3324),
    .A1(net2986),
    .S(_05087_),
    .X(_01309_));
 sg13g2_mux2_1 _13648_ (.A0(net3278),
    .A1(net4115),
    .S(_05087_),
    .X(_01310_));
 sg13g2_nand2_2 _13649_ (.Y(_05088_),
    .A(_02337_),
    .B(net3027));
 sg13g2_mux2_1 _13650_ (.A0(net3600),
    .A1(net4897),
    .S(_05088_),
    .X(_01311_));
 sg13g2_mux2_1 _13651_ (.A0(net3555),
    .A1(net2793),
    .S(_05088_),
    .X(_01312_));
 sg13g2_mux2_1 _13652_ (.A0(net3509),
    .A1(net4410),
    .S(_05088_),
    .X(_01313_));
 sg13g2_mux2_1 _13653_ (.A0(net3463),
    .A1(net2855),
    .S(_05088_),
    .X(_01314_));
 sg13g2_mux2_1 _13654_ (.A0(net3418),
    .A1(net4061),
    .S(_05088_),
    .X(_01315_));
 sg13g2_mux2_1 _13655_ (.A0(net3372),
    .A1(net4868),
    .S(_05088_),
    .X(_01316_));
 sg13g2_mux2_1 _13656_ (.A0(net3326),
    .A1(net4411),
    .S(_05088_),
    .X(_01317_));
 sg13g2_mux2_1 _13657_ (.A0(net3279),
    .A1(net4327),
    .S(_05088_),
    .X(_01318_));
 sg13g2_nand2_2 _13658_ (.Y(_05089_),
    .A(net3070),
    .B(net3028));
 sg13g2_mux2_1 _13659_ (.A0(net3598),
    .A1(net4028),
    .S(_05089_),
    .X(_01319_));
 sg13g2_mux2_1 _13660_ (.A0(net3553),
    .A1(net4801),
    .S(_05089_),
    .X(_01320_));
 sg13g2_mux2_1 _13661_ (.A0(net3509),
    .A1(net2945),
    .S(_05089_),
    .X(_01321_));
 sg13g2_mux2_1 _13662_ (.A0(net3463),
    .A1(net5072),
    .S(_05089_),
    .X(_01322_));
 sg13g2_mux2_1 _13663_ (.A0(net3418),
    .A1(net4643),
    .S(_05089_),
    .X(_01323_));
 sg13g2_mux2_1 _13664_ (.A0(net3372),
    .A1(net4688),
    .S(_05089_),
    .X(_01324_));
 sg13g2_mux2_1 _13665_ (.A0(net3326),
    .A1(net4702),
    .S(_05089_),
    .X(_01325_));
 sg13g2_mux2_1 _13666_ (.A0(net3279),
    .A1(net4565),
    .S(_05089_),
    .X(_01326_));
 sg13g2_nand2_2 _13667_ (.Y(_05090_),
    .A(_02330_),
    .B(net3027));
 sg13g2_mux2_1 _13668_ (.A0(net3598),
    .A1(net4805),
    .S(_05090_),
    .X(_01327_));
 sg13g2_mux2_1 _13669_ (.A0(net3555),
    .A1(net2871),
    .S(_05090_),
    .X(_01328_));
 sg13g2_mux2_1 _13670_ (.A0(net3509),
    .A1(net4290),
    .S(_05090_),
    .X(_01329_));
 sg13g2_mux2_1 _13671_ (.A0(net3463),
    .A1(net4485),
    .S(_05090_),
    .X(_01330_));
 sg13g2_mux2_1 _13672_ (.A0(net3418),
    .A1(net2756),
    .S(_05090_),
    .X(_01331_));
 sg13g2_mux2_1 _13673_ (.A0(net3372),
    .A1(net4725),
    .S(_05090_),
    .X(_01332_));
 sg13g2_mux2_1 _13674_ (.A0(net3326),
    .A1(net4788),
    .S(_05090_),
    .X(_01333_));
 sg13g2_mux2_1 _13675_ (.A0(net3279),
    .A1(net4987),
    .S(_05090_),
    .X(_01334_));
 sg13g2_nand2_2 _13676_ (.Y(_05091_),
    .A(net3071),
    .B(net3027));
 sg13g2_mux2_1 _13677_ (.A0(net3598),
    .A1(net4778),
    .S(_05091_),
    .X(_01335_));
 sg13g2_mux2_1 _13678_ (.A0(net3555),
    .A1(net4962),
    .S(_05091_),
    .X(_01336_));
 sg13g2_mux2_1 _13679_ (.A0(net3509),
    .A1(net2996),
    .S(_05091_),
    .X(_01337_));
 sg13g2_mux2_1 _13680_ (.A0(net3463),
    .A1(net4087),
    .S(_05091_),
    .X(_01338_));
 sg13g2_mux2_1 _13681_ (.A0(net3418),
    .A1(net4320),
    .S(_05091_),
    .X(_01339_));
 sg13g2_mux2_1 _13682_ (.A0(net3372),
    .A1(net4219),
    .S(_05091_),
    .X(_01340_));
 sg13g2_mux2_1 _13683_ (.A0(net3326),
    .A1(net5112),
    .S(_05091_),
    .X(_01341_));
 sg13g2_mux2_1 _13684_ (.A0(net3279),
    .A1(net4046),
    .S(_05091_),
    .X(_01342_));
 sg13g2_nand2_2 _13685_ (.Y(_05092_),
    .A(net3072),
    .B(_02365_));
 sg13g2_mux2_1 _13686_ (.A0(net3597),
    .A1(net4570),
    .S(_05092_),
    .X(_01343_));
 sg13g2_mux2_1 _13687_ (.A0(net3551),
    .A1(net4848),
    .S(_05092_),
    .X(_01344_));
 sg13g2_mux2_1 _13688_ (.A0(net3504),
    .A1(net2938),
    .S(_05092_),
    .X(_01345_));
 sg13g2_mux2_1 _13689_ (.A0(net3460),
    .A1(net4300),
    .S(_05092_),
    .X(_01346_));
 sg13g2_mux2_1 _13690_ (.A0(net3414),
    .A1(net2896),
    .S(_05092_),
    .X(_01347_));
 sg13g2_mux2_1 _13691_ (.A0(net3361),
    .A1(net4075),
    .S(_05092_),
    .X(_01348_));
 sg13g2_mux2_1 _13692_ (.A0(net3317),
    .A1(net4746),
    .S(_05092_),
    .X(_01349_));
 sg13g2_mux2_1 _13693_ (.A0(net3276),
    .A1(net4997),
    .S(_05092_),
    .X(_01350_));
 sg13g2_nand2_2 _13694_ (.Y(_05093_),
    .A(net3073),
    .B(net3027));
 sg13g2_mux2_1 _13695_ (.A0(net3596),
    .A1(net2982),
    .S(_05093_),
    .X(_01351_));
 sg13g2_mux2_1 _13696_ (.A0(net3551),
    .A1(net4825),
    .S(_05093_),
    .X(_01352_));
 sg13g2_mux2_1 _13697_ (.A0(net3504),
    .A1(net2881),
    .S(_05093_),
    .X(_01353_));
 sg13g2_mux2_1 _13698_ (.A0(net3460),
    .A1(net4600),
    .S(_05093_),
    .X(_01354_));
 sg13g2_mux2_1 _13699_ (.A0(net3415),
    .A1(net4985),
    .S(_05093_),
    .X(_01355_));
 sg13g2_mux2_1 _13700_ (.A0(net3361),
    .A1(net2902),
    .S(_05093_),
    .X(_01356_));
 sg13g2_mux2_1 _13701_ (.A0(net3317),
    .A1(net4012),
    .S(_05093_),
    .X(_01357_));
 sg13g2_mux2_1 _13702_ (.A0(net3276),
    .A1(net4559),
    .S(_05093_),
    .X(_01358_));
 sg13g2_nand2_2 _13703_ (.Y(_05094_),
    .A(net3084),
    .B(net3027));
 sg13g2_mux2_1 _13704_ (.A0(net3596),
    .A1(net4051),
    .S(_05094_),
    .X(_01359_));
 sg13g2_mux2_1 _13705_ (.A0(net3551),
    .A1(net2919),
    .S(_05094_),
    .X(_01360_));
 sg13g2_mux2_1 _13706_ (.A0(net3505),
    .A1(net4560),
    .S(_05094_),
    .X(_01361_));
 sg13g2_mux2_1 _13707_ (.A0(net3460),
    .A1(net2882),
    .S(_05094_),
    .X(_01362_));
 sg13g2_mux2_1 _13708_ (.A0(net3415),
    .A1(net4133),
    .S(_05094_),
    .X(_01363_));
 sg13g2_mux2_1 _13709_ (.A0(net3361),
    .A1(net4306),
    .S(_05094_),
    .X(_01364_));
 sg13g2_mux2_1 _13710_ (.A0(net3317),
    .A1(net4438),
    .S(_05094_),
    .X(_01365_));
 sg13g2_mux2_1 _13711_ (.A0(net3276),
    .A1(net4191),
    .S(_05094_),
    .X(_01366_));
 sg13g2_and2_2 _13712_ (.A(net3077),
    .B(_02311_),
    .X(_05095_));
 sg13g2_mux2_1 _13713_ (.A0(net2711),
    .A1(net3591),
    .S(_05095_),
    .X(_01367_));
 sg13g2_mux2_1 _13714_ (.A0(net2572),
    .A1(net3538),
    .S(_05095_),
    .X(_01368_));
 sg13g2_mux2_1 _13715_ (.A0(net2837),
    .A1(net3500),
    .S(_05095_),
    .X(_01369_));
 sg13g2_mux2_1 _13716_ (.A0(net2695),
    .A1(net3455),
    .S(_05095_),
    .X(_01370_));
 sg13g2_mux2_1 _13717_ (.A0(net2740),
    .A1(net3409),
    .S(_05095_),
    .X(_01371_));
 sg13g2_mux2_1 _13718_ (.A0(net2277),
    .A1(net3365),
    .S(_05095_),
    .X(_01372_));
 sg13g2_mux2_1 _13719_ (.A0(net2742),
    .A1(net3312),
    .S(_05095_),
    .X(_01373_));
 sg13g2_mux2_1 _13720_ (.A0(net2409),
    .A1(net3281),
    .S(_05095_),
    .X(_01374_));
 sg13g2_and2_2 _13721_ (.A(net3079),
    .B(net3029),
    .X(_05096_));
 sg13g2_mux2_1 _13722_ (.A0(net2553),
    .A1(net3575),
    .S(_05096_),
    .X(_01375_));
 sg13g2_mux2_1 _13723_ (.A0(net2484),
    .A1(net3527),
    .S(_05096_),
    .X(_01376_));
 sg13g2_mux2_1 _13724_ (.A0(net2319),
    .A1(net3491),
    .S(_05096_),
    .X(_01377_));
 sg13g2_mux2_1 _13725_ (.A0(net2207),
    .A1(net3444),
    .S(_05096_),
    .X(_01378_));
 sg13g2_mux2_1 _13726_ (.A0(net2457),
    .A1(net3399),
    .S(_05096_),
    .X(_01379_));
 sg13g2_mux2_1 _13727_ (.A0(net2199),
    .A1(net3353),
    .S(_05096_),
    .X(_01380_));
 sg13g2_mux2_1 _13728_ (.A0(net2806),
    .A1(net3301),
    .S(_05096_),
    .X(_01381_));
 sg13g2_mux2_1 _13729_ (.A0(net2542),
    .A1(net3258),
    .S(_05096_),
    .X(_01382_));
 sg13g2_nand2_2 _13730_ (.Y(_05097_),
    .A(_02297_),
    .B(net3029));
 sg13g2_mux2_1 _13731_ (.A0(net3575),
    .A1(net4615),
    .S(_05097_),
    .X(_01383_));
 sg13g2_mux2_1 _13732_ (.A0(net3527),
    .A1(net4445),
    .S(_05097_),
    .X(_01384_));
 sg13g2_mux2_1 _13733_ (.A0(net3491),
    .A1(net3005),
    .S(_05097_),
    .X(_01385_));
 sg13g2_mux2_1 _13734_ (.A0(net3446),
    .A1(net4803),
    .S(_05097_),
    .X(_01386_));
 sg13g2_mux2_1 _13735_ (.A0(net3399),
    .A1(net4483),
    .S(_05097_),
    .X(_01387_));
 sg13g2_mux2_1 _13736_ (.A0(net3354),
    .A1(net4180),
    .S(_05097_),
    .X(_01388_));
 sg13g2_mux2_1 _13737_ (.A0(net3300),
    .A1(net5089),
    .S(_05097_),
    .X(_01389_));
 sg13g2_mux2_1 _13738_ (.A0(net3258),
    .A1(net2942),
    .S(_05097_),
    .X(_01390_));
 sg13g2_nand2_2 _13739_ (.Y(_05098_),
    .A(_02293_),
    .B(_02362_));
 sg13g2_mux2_1 _13740_ (.A0(net3575),
    .A1(net4686),
    .S(_05098_),
    .X(_01391_));
 sg13g2_mux2_1 _13741_ (.A0(net3527),
    .A1(net4677),
    .S(_05098_),
    .X(_01392_));
 sg13g2_mux2_1 _13742_ (.A0(net3491),
    .A1(net2672),
    .S(_05098_),
    .X(_01393_));
 sg13g2_mux2_1 _13743_ (.A0(net3444),
    .A1(net4862),
    .S(_05098_),
    .X(_01394_));
 sg13g2_mux2_1 _13744_ (.A0(net3399),
    .A1(net4458),
    .S(_05098_),
    .X(_01395_));
 sg13g2_mux2_1 _13745_ (.A0(net3354),
    .A1(net4196),
    .S(_05098_),
    .X(_01396_));
 sg13g2_mux2_1 _13746_ (.A0(net3300),
    .A1(net4130),
    .S(_05098_),
    .X(_01397_));
 sg13g2_mux2_1 _13747_ (.A0(net3260),
    .A1(net4134),
    .S(_05098_),
    .X(_01398_));
 sg13g2_nand2_2 _13748_ (.Y(_05099_),
    .A(_02349_),
    .B(net3029));
 sg13g2_mux2_1 _13749_ (.A0(net3575),
    .A1(net2916),
    .S(_05099_),
    .X(_01399_));
 sg13g2_mux2_1 _13750_ (.A0(net3527),
    .A1(net4047),
    .S(_05099_),
    .X(_01400_));
 sg13g2_mux2_1 _13751_ (.A0(net3491),
    .A1(net5028),
    .S(_05099_),
    .X(_01401_));
 sg13g2_mux2_1 _13752_ (.A0(net3444),
    .A1(net4907),
    .S(_05099_),
    .X(_01402_));
 sg13g2_mux2_1 _13753_ (.A0(net3399),
    .A1(net4463),
    .S(_05099_),
    .X(_01403_));
 sg13g2_mux2_1 _13754_ (.A0(net3354),
    .A1(net3006),
    .S(_05099_),
    .X(_01404_));
 sg13g2_mux2_1 _13755_ (.A0(net3300),
    .A1(net4903),
    .S(_05099_),
    .X(_01405_));
 sg13g2_mux2_1 _13756_ (.A0(net3260),
    .A1(net5123),
    .S(_05099_),
    .X(_01406_));
 sg13g2_nand2_2 _13757_ (.Y(_05100_),
    .A(_02277_),
    .B(net3029));
 sg13g2_mux2_1 _13758_ (.A0(net3584),
    .A1(net4863),
    .S(_05100_),
    .X(_01407_));
 sg13g2_mux2_1 _13759_ (.A0(net3535),
    .A1(net5128),
    .S(_05100_),
    .X(_01408_));
 sg13g2_mux2_1 _13760_ (.A0(net3494),
    .A1(net2666),
    .S(_05100_),
    .X(_01409_));
 sg13g2_mux2_1 _13761_ (.A0(net3448),
    .A1(net2883),
    .S(_05100_),
    .X(_01410_));
 sg13g2_mux2_1 _13762_ (.A0(net3399),
    .A1(net4603),
    .S(_05100_),
    .X(_01411_));
 sg13g2_mux2_1 _13763_ (.A0(net3359),
    .A1(net2903),
    .S(_05100_),
    .X(_01412_));
 sg13g2_mux2_1 _13764_ (.A0(net3309),
    .A1(net4543),
    .S(_05100_),
    .X(_01413_));
 sg13g2_mux2_1 _13765_ (.A0(net3260),
    .A1(net4351),
    .S(_05100_),
    .X(_01414_));
 sg13g2_nand2_2 _13766_ (.Y(_05101_),
    .A(net3069),
    .B(net3029));
 sg13g2_mux2_1 _13767_ (.A0(net3584),
    .A1(net4359),
    .S(_05101_),
    .X(_01415_));
 sg13g2_mux2_1 _13768_ (.A0(net3535),
    .A1(net4719),
    .S(_05101_),
    .X(_01416_));
 sg13g2_mux2_1 _13769_ (.A0(net3494),
    .A1(net5035),
    .S(_05101_),
    .X(_01417_));
 sg13g2_mux2_1 _13770_ (.A0(net3448),
    .A1(net4666),
    .S(_05101_),
    .X(_01418_));
 sg13g2_mux2_1 _13771_ (.A0(net3399),
    .A1(net2981),
    .S(_05101_),
    .X(_01419_));
 sg13g2_mux2_1 _13772_ (.A0(net3359),
    .A1(net4070),
    .S(_05101_),
    .X(_01420_));
 sg13g2_mux2_1 _13773_ (.A0(net3313),
    .A1(net4557),
    .S(_05101_),
    .X(_01421_));
 sg13g2_mux2_1 _13774_ (.A0(net3260),
    .A1(net4797),
    .S(_05101_),
    .X(_01422_));
 sg13g2_nand2_2 _13775_ (.Y(_05102_),
    .A(net3029),
    .B(net3065));
 sg13g2_mux2_1 _13776_ (.A0(net3583),
    .A1(net2877),
    .S(_05102_),
    .X(_01423_));
 sg13g2_mux2_1 _13777_ (.A0(net3539),
    .A1(net4099),
    .S(_05102_),
    .X(_01424_));
 sg13g2_mux2_1 _13778_ (.A0(net3491),
    .A1(net4841),
    .S(_05102_),
    .X(_01425_));
 sg13g2_mux2_1 _13779_ (.A0(net3444),
    .A1(net4827),
    .S(_05102_),
    .X(_01426_));
 sg13g2_mux2_1 _13780_ (.A0(net3402),
    .A1(net2907),
    .S(_05102_),
    .X(_01427_));
 sg13g2_mux2_1 _13781_ (.A0(net3354),
    .A1(net4400),
    .S(_05102_),
    .X(_01428_));
 sg13g2_mux2_1 _13782_ (.A0(net3313),
    .A1(net2748),
    .S(_05102_),
    .X(_01429_));
 sg13g2_mux2_1 _13783_ (.A0(net3260),
    .A1(net4707),
    .S(_05102_),
    .X(_01430_));
 sg13g2_nand2_2 _13784_ (.Y(_05103_),
    .A(net3049),
    .B(_02362_));
 sg13g2_mux2_1 _13785_ (.A0(net3575),
    .A1(net4288),
    .S(_05103_),
    .X(_01431_));
 sg13g2_mux2_1 _13786_ (.A0(net3539),
    .A1(net4771),
    .S(_05103_),
    .X(_01432_));
 sg13g2_mux2_1 _13787_ (.A0(net3491),
    .A1(net4230),
    .S(_05103_),
    .X(_01433_));
 sg13g2_mux2_1 _13788_ (.A0(net3444),
    .A1(net4953),
    .S(_05103_),
    .X(_01434_));
 sg13g2_mux2_1 _13789_ (.A0(net3402),
    .A1(net2917),
    .S(_05103_),
    .X(_01435_));
 sg13g2_mux2_1 _13790_ (.A0(net3353),
    .A1(net4479),
    .S(_05103_),
    .X(_01436_));
 sg13g2_mux2_1 _13791_ (.A0(net3313),
    .A1(net4436),
    .S(_05103_),
    .X(_01437_));
 sg13g2_mux2_1 _13792_ (.A0(net3260),
    .A1(net4157),
    .S(_05103_),
    .X(_01438_));
 sg13g2_nand2_2 _13793_ (.Y(_05104_),
    .A(_02337_),
    .B(net3030));
 sg13g2_mux2_1 _13794_ (.A0(net3579),
    .A1(net4253),
    .S(_05104_),
    .X(_01439_));
 sg13g2_mux2_1 _13795_ (.A0(net3532),
    .A1(net4845),
    .S(_05104_),
    .X(_01440_));
 sg13g2_mux2_1 _13796_ (.A0(net3485),
    .A1(net4655),
    .S(_05104_),
    .X(_01441_));
 sg13g2_mux2_1 _13797_ (.A0(net3438),
    .A1(net4212),
    .S(_05104_),
    .X(_01442_));
 sg13g2_mux2_1 _13798_ (.A0(net3395),
    .A1(net2702),
    .S(_05104_),
    .X(_01443_));
 sg13g2_mux2_1 _13799_ (.A0(net3349),
    .A1(net5083),
    .S(_05104_),
    .X(_01444_));
 sg13g2_mux2_1 _13800_ (.A0(net3305),
    .A1(net5088),
    .S(_05104_),
    .X(_01445_));
 sg13g2_mux2_1 _13801_ (.A0(net3254),
    .A1(net4625),
    .S(_05104_),
    .X(_01446_));
 sg13g2_nand2_2 _13802_ (.Y(_05105_),
    .A(net3079),
    .B(net3034));
 sg13g2_mux2_1 _13803_ (.A0(net3591),
    .A1(net2976),
    .S(_05105_),
    .X(_01447_));
 sg13g2_mux2_1 _13804_ (.A0(net3545),
    .A1(net2582),
    .S(_05105_),
    .X(_01448_));
 sg13g2_mux2_1 _13805_ (.A0(net3499),
    .A1(net4525),
    .S(_05105_),
    .X(_01449_));
 sg13g2_mux2_1 _13806_ (.A0(net3455),
    .A1(net4391),
    .S(_05105_),
    .X(_01450_));
 sg13g2_mux2_1 _13807_ (.A0(net3410),
    .A1(net2713),
    .S(_05105_),
    .X(_01451_));
 sg13g2_mux2_1 _13808_ (.A0(net3366),
    .A1(net2967),
    .S(_05105_),
    .X(_01452_));
 sg13g2_mux2_1 _13809_ (.A0(net3321),
    .A1(net2705),
    .S(_05105_),
    .X(_01453_));
 sg13g2_mux2_1 _13810_ (.A0(net3270),
    .A1(net2965),
    .S(_05105_),
    .X(_01454_));
 sg13g2_nand2_2 _13811_ (.Y(_05106_),
    .A(_02330_),
    .B(net3030));
 sg13g2_mux2_1 _13812_ (.A0(net3579),
    .A1(net4720),
    .S(_05106_),
    .X(_01455_));
 sg13g2_mux2_1 _13813_ (.A0(net3540),
    .A1(net2924),
    .S(_05106_),
    .X(_01456_));
 sg13g2_mux2_1 _13814_ (.A0(net3485),
    .A1(net4952),
    .S(_05106_),
    .X(_01457_));
 sg13g2_mux2_1 _13815_ (.A0(net3447),
    .A1(net2922),
    .S(_05106_),
    .X(_01458_));
 sg13g2_mux2_1 _13816_ (.A0(net3395),
    .A1(net2795),
    .S(_05106_),
    .X(_01459_));
 sg13g2_mux2_1 _13817_ (.A0(net3349),
    .A1(net4039),
    .S(_05106_),
    .X(_01460_));
 sg13g2_mux2_1 _13818_ (.A0(net3305),
    .A1(net4601),
    .S(_05106_),
    .X(_01461_));
 sg13g2_mux2_1 _13819_ (.A0(net3254),
    .A1(net4177),
    .S(_05106_),
    .X(_01462_));
 sg13g2_nand2_2 _13820_ (.Y(_05107_),
    .A(net3071),
    .B(net3029));
 sg13g2_mux2_1 _13821_ (.A0(net3579),
    .A1(net4703),
    .S(_05107_),
    .X(_01463_));
 sg13g2_mux2_1 _13822_ (.A0(net3540),
    .A1(net4700),
    .S(_05107_),
    .X(_01464_));
 sg13g2_mux2_1 _13823_ (.A0(net3485),
    .A1(net4942),
    .S(_05107_),
    .X(_01465_));
 sg13g2_mux2_1 _13824_ (.A0(net3447),
    .A1(net4409),
    .S(_05107_),
    .X(_01466_));
 sg13g2_mux2_1 _13825_ (.A0(net3395),
    .A1(net4924),
    .S(_05107_),
    .X(_01467_));
 sg13g2_mux2_1 _13826_ (.A0(net3349),
    .A1(net4722),
    .S(_05107_),
    .X(_01468_));
 sg13g2_mux2_1 _13827_ (.A0(net3305),
    .A1(net4120),
    .S(_05107_),
    .X(_01469_));
 sg13g2_mux2_1 _13828_ (.A0(net3254),
    .A1(net4011),
    .S(_05107_),
    .X(_01470_));
 sg13g2_nand2_2 _13829_ (.Y(_05108_),
    .A(net3072),
    .B(_02362_));
 sg13g2_mux2_1 _13830_ (.A0(net3575),
    .A1(net2845),
    .S(_05108_),
    .X(_01471_));
 sg13g2_mux2_1 _13831_ (.A0(net3528),
    .A1(net4486),
    .S(_05108_),
    .X(_01472_));
 sg13g2_mux2_1 _13832_ (.A0(net3488),
    .A1(net2860),
    .S(_05108_),
    .X(_01473_));
 sg13g2_mux2_1 _13833_ (.A0(net3436),
    .A1(net4322),
    .S(_05108_),
    .X(_01474_));
 sg13g2_mux2_1 _13834_ (.A0(net3390),
    .A1(net2898),
    .S(_05108_),
    .X(_01475_));
 sg13g2_mux2_1 _13835_ (.A0(net3346),
    .A1(net2708),
    .S(_05108_),
    .X(_01476_));
 sg13g2_mux2_1 _13836_ (.A0(net3300),
    .A1(net2766),
    .S(_05108_),
    .X(_01477_));
 sg13g2_mux2_1 _13837_ (.A0(net3253),
    .A1(net4124),
    .S(_05108_),
    .X(_01478_));
 sg13g2_nand2_2 _13838_ (.Y(_05109_),
    .A(net3073),
    .B(net3029));
 sg13g2_mux2_1 _13839_ (.A0(net3576),
    .A1(net4229),
    .S(_05109_),
    .X(_01479_));
 sg13g2_mux2_1 _13840_ (.A0(net3528),
    .A1(net4270),
    .S(_05109_),
    .X(_01480_));
 sg13g2_mux2_1 _13841_ (.A0(net3482),
    .A1(net4383),
    .S(_05109_),
    .X(_01481_));
 sg13g2_mux2_1 _13842_ (.A0(net3436),
    .A1(net4774),
    .S(_05109_),
    .X(_01482_));
 sg13g2_mux2_1 _13843_ (.A0(net3390),
    .A1(net5033),
    .S(_05109_),
    .X(_01483_));
 sg13g2_mux2_1 _13844_ (.A0(net3346),
    .A1(net5006),
    .S(_05109_),
    .X(_01484_));
 sg13g2_mux2_1 _13845_ (.A0(net3300),
    .A1(net4276),
    .S(_05109_),
    .X(_01485_));
 sg13g2_mux2_1 _13846_ (.A0(net3253),
    .A1(net4553),
    .S(_05109_),
    .X(_01486_));
 sg13g2_nand2_1 _13847_ (.Y(_05110_),
    .A(net3084),
    .B(net3030));
 sg13g2_mux2_1 _13848_ (.A0(net3577),
    .A1(net4596),
    .S(net3013),
    .X(_01487_));
 sg13g2_mux2_1 _13849_ (.A0(net3529),
    .A1(net2771),
    .S(net3013),
    .X(_01488_));
 sg13g2_mux2_1 _13850_ (.A0(net3486),
    .A1(net2866),
    .S(net3013),
    .X(_01489_));
 sg13g2_mux2_1 _13851_ (.A0(net3438),
    .A1(net2698),
    .S(net3013),
    .X(_01490_));
 sg13g2_mux2_1 _13852_ (.A0(net3390),
    .A1(net4639),
    .S(_05110_),
    .X(_01491_));
 sg13g2_nor2_1 _13853_ (.A(net3349),
    .B(net3013),
    .Y(_05111_));
 sg13g2_a21oi_1 _13854_ (.A1(_02162_),
    .A2(net3013),
    .Y(_01492_),
    .B1(_05111_));
 sg13g2_mux2_1 _13855_ (.A0(net3300),
    .A1(net4369),
    .S(net3013),
    .X(_01493_));
 sg13g2_mux2_1 _13856_ (.A0(net3253),
    .A1(net4305),
    .S(net3013),
    .X(_01494_));
 sg13g2_and2_2 _13857_ (.A(net3077),
    .B(net3030),
    .X(_05112_));
 sg13g2_mux2_1 _13858_ (.A0(net2307),
    .A1(net3577),
    .S(_05112_),
    .X(_01495_));
 sg13g2_mux2_1 _13859_ (.A0(net2757),
    .A1(net3527),
    .S(_05112_),
    .X(_01496_));
 sg13g2_mux2_1 _13860_ (.A0(net2610),
    .A1(net3482),
    .S(_05112_),
    .X(_01497_));
 sg13g2_mux2_1 _13861_ (.A0(net2764),
    .A1(net3447),
    .S(_05112_),
    .X(_01498_));
 sg13g2_mux2_1 _13862_ (.A0(net2270),
    .A1(net3395),
    .S(_05112_),
    .X(_01499_));
 sg13g2_mux2_1 _13863_ (.A0(net2694),
    .A1(net3349),
    .S(_05112_),
    .X(_01500_));
 sg13g2_mux2_1 _13864_ (.A0(net2259),
    .A1(net3300),
    .S(_05112_),
    .X(_01501_));
 sg13g2_mux2_1 _13865_ (.A0(net2294),
    .A1(net3253),
    .S(_05112_),
    .X(_01502_));
 sg13g2_and2_2 _13866_ (.A(net3079),
    .B(net3031),
    .X(_05113_));
 sg13g2_mux2_1 _13867_ (.A0(net2491),
    .A1(net3579),
    .S(_05113_),
    .X(_01503_));
 sg13g2_mux2_1 _13868_ (.A0(net2205),
    .A1(net3532),
    .S(_05113_),
    .X(_01504_));
 sg13g2_mux2_1 _13869_ (.A0(net2154),
    .A1(net3486),
    .S(_05113_),
    .X(_01505_));
 sg13g2_mux2_1 _13870_ (.A0(net2555),
    .A1(net3440),
    .S(_05113_),
    .X(_01506_));
 sg13g2_mux2_1 _13871_ (.A0(net2371),
    .A1(net3392),
    .S(_05113_),
    .X(_01507_));
 sg13g2_mux2_1 _13872_ (.A0(net2208),
    .A1(net3350),
    .S(_05113_),
    .X(_01508_));
 sg13g2_mux2_1 _13873_ (.A0(net2379),
    .A1(net3305),
    .S(_05113_),
    .X(_01509_));
 sg13g2_mux2_1 _13874_ (.A0(net2394),
    .A1(net3254),
    .S(_05113_),
    .X(_01510_));
 sg13g2_nand2_2 _13875_ (.Y(_05114_),
    .A(_02297_),
    .B(net3031));
 sg13g2_mux2_1 _13876_ (.A0(net3578),
    .A1(net4103),
    .S(_05114_),
    .X(_01511_));
 sg13g2_mux2_1 _13877_ (.A0(net3532),
    .A1(net4846),
    .S(_05114_),
    .X(_01512_));
 sg13g2_mux2_1 _13878_ (.A0(net3486),
    .A1(net5011),
    .S(_05114_),
    .X(_01513_));
 sg13g2_mux2_1 _13879_ (.A0(net3438),
    .A1(net4441),
    .S(_05114_),
    .X(_01514_));
 sg13g2_mux2_1 _13880_ (.A0(net3392),
    .A1(net5137),
    .S(_05114_),
    .X(_01515_));
 sg13g2_mux2_1 _13881_ (.A0(net3350),
    .A1(net4484),
    .S(_05114_),
    .X(_01516_));
 sg13g2_mux2_1 _13882_ (.A0(net3305),
    .A1(net2988),
    .S(_05114_),
    .X(_01517_));
 sg13g2_mux2_1 _13883_ (.A0(net3254),
    .A1(net4104),
    .S(_05114_),
    .X(_01518_));
 sg13g2_nand2_2 _13884_ (.Y(_05115_),
    .A(_02288_),
    .B(net3031));
 sg13g2_mux2_1 _13885_ (.A0(net3579),
    .A1(net4407),
    .S(_05115_),
    .X(_01519_));
 sg13g2_mux2_1 _13886_ (.A0(net3532),
    .A1(net4663),
    .S(_05115_),
    .X(_01520_));
 sg13g2_mux2_1 _13887_ (.A0(net3486),
    .A1(net2743),
    .S(_05115_),
    .X(_01521_));
 sg13g2_mux2_1 _13888_ (.A0(net3438),
    .A1(net5106),
    .S(_05115_),
    .X(_01522_));
 sg13g2_mux2_1 _13889_ (.A0(net3392),
    .A1(net4316),
    .S(_05115_),
    .X(_01523_));
 sg13g2_mux2_1 _13890_ (.A0(net3350),
    .A1(net4776),
    .S(_05115_),
    .X(_01524_));
 sg13g2_mux2_1 _13891_ (.A0(net3305),
    .A1(net5015),
    .S(_05115_),
    .X(_01525_));
 sg13g2_mux2_1 _13892_ (.A0(net3254),
    .A1(net4945),
    .S(_05115_),
    .X(_01526_));
 sg13g2_nand2_2 _13893_ (.Y(_05116_),
    .A(_02297_),
    .B(net3034));
 sg13g2_mux2_1 _13894_ (.A0(net3590),
    .A1(net4800),
    .S(_05116_),
    .X(_01527_));
 sg13g2_mux2_1 _13895_ (.A0(net3545),
    .A1(net5152),
    .S(_05116_),
    .X(_01528_));
 sg13g2_mux2_1 _13896_ (.A0(net3499),
    .A1(net4929),
    .S(_05116_),
    .X(_01529_));
 sg13g2_mux2_1 _13897_ (.A0(net3454),
    .A1(net5063),
    .S(_05116_),
    .X(_01530_));
 sg13g2_mux2_1 _13898_ (.A0(net3410),
    .A1(net5174),
    .S(_05116_),
    .X(_01531_));
 sg13g2_mux2_1 _13899_ (.A0(net3366),
    .A1(net4896),
    .S(_05116_),
    .X(_01532_));
 sg13g2_mux2_1 _13900_ (.A0(net3321),
    .A1(net5143),
    .S(_05116_),
    .X(_01533_));
 sg13g2_mux2_1 _13901_ (.A0(net3269),
    .A1(net4294),
    .S(_05116_),
    .X(_01534_));
 sg13g2_nand2_2 _13902_ (.Y(_05117_),
    .A(_02277_),
    .B(net3031));
 sg13g2_mux2_1 _13903_ (.A0(net3580),
    .A1(net2804),
    .S(_05117_),
    .X(_01535_));
 sg13g2_mux2_1 _13904_ (.A0(net3533),
    .A1(net4660),
    .S(_05117_),
    .X(_01536_));
 sg13g2_mux2_1 _13905_ (.A0(net3487),
    .A1(net2833),
    .S(_05117_),
    .X(_01537_));
 sg13g2_mux2_1 _13906_ (.A0(net3440),
    .A1(net4806),
    .S(_05117_),
    .X(_01538_));
 sg13g2_mux2_1 _13907_ (.A0(net3393),
    .A1(net5178),
    .S(_05117_),
    .X(_01539_));
 sg13g2_mux2_1 _13908_ (.A0(net3349),
    .A1(net4314),
    .S(_05117_),
    .X(_01540_));
 sg13g2_mux2_1 _13909_ (.A0(net3306),
    .A1(net2626),
    .S(_05117_),
    .X(_01541_));
 sg13g2_mux2_1 _13910_ (.A0(net3255),
    .A1(net2954),
    .S(_05117_),
    .X(_01542_));
 sg13g2_nand2_2 _13911_ (.Y(_05118_),
    .A(net3069),
    .B(net3032));
 sg13g2_mux2_1 _13912_ (.A0(net3579),
    .A1(net4564),
    .S(_05118_),
    .X(_01543_));
 sg13g2_mux2_1 _13913_ (.A0(net3533),
    .A1(net3003),
    .S(_05118_),
    .X(_01544_));
 sg13g2_mux2_1 _13914_ (.A0(net3487),
    .A1(net5084),
    .S(_05118_),
    .X(_01545_));
 sg13g2_mux2_1 _13915_ (.A0(net3440),
    .A1(net4412),
    .S(_05118_),
    .X(_01546_));
 sg13g2_mux2_1 _13916_ (.A0(net3404),
    .A1(net5050),
    .S(_05118_),
    .X(_01547_));
 sg13g2_mux2_1 _13917_ (.A0(net3350),
    .A1(net4146),
    .S(_05118_),
    .X(_01548_));
 sg13g2_mux2_1 _13918_ (.A0(net3306),
    .A1(net4481),
    .S(_05118_),
    .X(_01549_));
 sg13g2_mux2_1 _13919_ (.A0(net3255),
    .A1(net4109),
    .S(_05118_),
    .X(_01550_));
 sg13g2_nand2_2 _13920_ (.Y(_05119_),
    .A(net3031),
    .B(net3065));
 sg13g2_mux2_1 _13921_ (.A0(net3580),
    .A1(net4284),
    .S(_05119_),
    .X(_01551_));
 sg13g2_mux2_1 _13922_ (.A0(net3532),
    .A1(net5133),
    .S(_05119_),
    .X(_01552_));
 sg13g2_mux2_1 _13923_ (.A0(net3486),
    .A1(net2703),
    .S(_05119_),
    .X(_01553_));
 sg13g2_mux2_1 _13924_ (.A0(net3449),
    .A1(net4199),
    .S(_05119_),
    .X(_01554_));
 sg13g2_mux2_1 _13925_ (.A0(net3392),
    .A1(net2952),
    .S(_05119_),
    .X(_01555_));
 sg13g2_mux2_1 _13926_ (.A0(net3350),
    .A1(net4416),
    .S(_05119_),
    .X(_01556_));
 sg13g2_mux2_1 _13927_ (.A0(net3306),
    .A1(net2875),
    .S(_05119_),
    .X(_01557_));
 sg13g2_mux2_1 _13928_ (.A0(net3254),
    .A1(net4837),
    .S(_05119_),
    .X(_01558_));
 sg13g2_nand2_2 _13929_ (.Y(_05120_),
    .A(_02309_),
    .B(net3031));
 sg13g2_mux2_1 _13930_ (.A0(net3580),
    .A1(net4474),
    .S(_05120_),
    .X(_01559_));
 sg13g2_mux2_1 _13931_ (.A0(net3532),
    .A1(net2933),
    .S(_05120_),
    .X(_01560_));
 sg13g2_mux2_1 _13932_ (.A0(net3486),
    .A1(net4421),
    .S(_05120_),
    .X(_01561_));
 sg13g2_mux2_1 _13933_ (.A0(net3449),
    .A1(net4554),
    .S(_05120_),
    .X(_01562_));
 sg13g2_mux2_1 _13934_ (.A0(net3392),
    .A1(net4102),
    .S(_05120_),
    .X(_01563_));
 sg13g2_mux2_1 _13935_ (.A0(net3350),
    .A1(net4651),
    .S(_05120_),
    .X(_01564_));
 sg13g2_mux2_1 _13936_ (.A0(net3306),
    .A1(net4267),
    .S(_05120_),
    .X(_01565_));
 sg13g2_mux2_1 _13937_ (.A0(net3255),
    .A1(net5144),
    .S(_05120_),
    .X(_01566_));
 sg13g2_nand2_2 _13938_ (.Y(_05121_),
    .A(_02337_),
    .B(net3032));
 sg13g2_mux2_1 _13939_ (.A0(net3581),
    .A1(net2784),
    .S(_05121_),
    .X(_01567_));
 sg13g2_mux2_1 _13940_ (.A0(net3531),
    .A1(net2803),
    .S(_05121_),
    .X(_01568_));
 sg13g2_mux2_1 _13941_ (.A0(net3483),
    .A1(net4067),
    .S(_05121_),
    .X(_01569_));
 sg13g2_mux2_1 _13942_ (.A0(net3439),
    .A1(net5051),
    .S(_05121_),
    .X(_01570_));
 sg13g2_mux2_1 _13943_ (.A0(net3394),
    .A1(net2873),
    .S(_05121_),
    .X(_01571_));
 sg13g2_mux2_1 _13944_ (.A0(net3351),
    .A1(net5166),
    .S(_05121_),
    .X(_01572_));
 sg13g2_mux2_1 _13945_ (.A0(net3304),
    .A1(net4163),
    .S(_05121_),
    .X(_01573_));
 sg13g2_mux2_1 _13946_ (.A0(net3255),
    .A1(net2900),
    .S(_05121_),
    .X(_01574_));
 sg13g2_nand2_2 _13947_ (.Y(_05122_),
    .A(net3070),
    .B(net3032));
 sg13g2_mux2_1 _13948_ (.A0(net3581),
    .A1(net5110),
    .S(_05122_),
    .X(_01575_));
 sg13g2_mux2_1 _13949_ (.A0(net3530),
    .A1(net4824),
    .S(_05122_),
    .X(_01576_));
 sg13g2_mux2_1 _13950_ (.A0(net3483),
    .A1(net4139),
    .S(_05122_),
    .X(_01577_));
 sg13g2_mux2_1 _13951_ (.A0(net3439),
    .A1(net4925),
    .S(_05122_),
    .X(_01578_));
 sg13g2_mux2_1 _13952_ (.A0(net3394),
    .A1(net4955),
    .S(_05122_),
    .X(_01579_));
 sg13g2_mux2_1 _13953_ (.A0(net3347),
    .A1(net4017),
    .S(_05122_),
    .X(_01580_));
 sg13g2_mux2_1 _13954_ (.A0(net3304),
    .A1(net4773),
    .S(_05122_),
    .X(_01581_));
 sg13g2_mux2_1 _13955_ (.A0(net3255),
    .A1(net4690),
    .S(_05122_),
    .X(_01582_));
 sg13g2_nand2_2 _13956_ (.Y(_05123_),
    .A(_02330_),
    .B(net3032));
 sg13g2_mux2_1 _13957_ (.A0(net3580),
    .A1(net2864),
    .S(_05123_),
    .X(_01583_));
 sg13g2_mux2_1 _13958_ (.A0(net3530),
    .A1(net2608),
    .S(_05123_),
    .X(_01584_));
 sg13g2_mux2_1 _13959_ (.A0(net3483),
    .A1(net4631),
    .S(_05123_),
    .X(_01585_));
 sg13g2_mux2_1 _13960_ (.A0(net3439),
    .A1(net2940),
    .S(_05123_),
    .X(_01586_));
 sg13g2_mux2_1 _13961_ (.A0(net3393),
    .A1(net2775),
    .S(_05123_),
    .X(_01587_));
 sg13g2_mux2_1 _13962_ (.A0(net3347),
    .A1(net4768),
    .S(_05123_),
    .X(_01588_));
 sg13g2_mux2_1 _13963_ (.A0(net3303),
    .A1(net5043),
    .S(_05123_),
    .X(_01589_));
 sg13g2_mux2_1 _13964_ (.A0(net3255),
    .A1(net4575),
    .S(_05123_),
    .X(_01590_));
 sg13g2_nand2_2 _13965_ (.Y(_05124_),
    .A(net3071),
    .B(net3032));
 sg13g2_mux2_1 _13966_ (.A0(net3580),
    .A1(net5116),
    .S(_05124_),
    .X(_01591_));
 sg13g2_mux2_1 _13967_ (.A0(net3530),
    .A1(net4882),
    .S(_05124_),
    .X(_01592_));
 sg13g2_mux2_1 _13968_ (.A0(net3483),
    .A1(net5079),
    .S(_05124_),
    .X(_01593_));
 sg13g2_mux2_1 _13969_ (.A0(net3439),
    .A1(net2993),
    .S(_05124_),
    .X(_01594_));
 sg13g2_mux2_1 _13970_ (.A0(net3393),
    .A1(net5019),
    .S(_05124_),
    .X(_01595_));
 sg13g2_mux2_1 _13971_ (.A0(net3347),
    .A1(net4448),
    .S(_05124_),
    .X(_01596_));
 sg13g2_mux2_1 _13972_ (.A0(net3303),
    .A1(net4125),
    .S(_05124_),
    .X(_01597_));
 sg13g2_mux2_1 _13973_ (.A0(net3255),
    .A1(net2977),
    .S(_05124_),
    .X(_01598_));
 sg13g2_or3_2 _13974_ (.A(net3088),
    .B(_02322_),
    .C(_02354_),
    .X(_05125_));
 sg13g2_mux2_1 _13975_ (.A0(net3578),
    .A1(net4342),
    .S(_05125_),
    .X(_01599_));
 sg13g2_mux2_1 _13976_ (.A0(net3530),
    .A1(net4921),
    .S(_05125_),
    .X(_01600_));
 sg13g2_mux2_1 _13977_ (.A0(net3483),
    .A1(net2836),
    .S(_05125_),
    .X(_01601_));
 sg13g2_mux2_1 _13978_ (.A0(net3439),
    .A1(net4153),
    .S(_05125_),
    .X(_01602_));
 sg13g2_mux2_1 _13979_ (.A0(net3394),
    .A1(net4293),
    .S(_05125_),
    .X(_01603_));
 sg13g2_mux2_1 _13980_ (.A0(net3347),
    .A1(net5000),
    .S(_05125_),
    .X(_01604_));
 sg13g2_mux2_1 _13981_ (.A0(net3304),
    .A1(net2761),
    .S(_05125_),
    .X(_01605_));
 sg13g2_mux2_1 _13982_ (.A0(net3256),
    .A1(net4030),
    .S(_05125_),
    .X(_01606_));
 sg13g2_nand2_2 _13983_ (.Y(_05126_),
    .A(_02288_),
    .B(net3034));
 sg13g2_mux2_1 _13984_ (.A0(net3590),
    .A1(net4766),
    .S(_05126_),
    .X(_01607_));
 sg13g2_mux2_1 _13985_ (.A0(net3545),
    .A1(net2659),
    .S(_05126_),
    .X(_01608_));
 sg13g2_mux2_1 _13986_ (.A0(net3499),
    .A1(net4430),
    .S(_05126_),
    .X(_01609_));
 sg13g2_mux2_1 _13987_ (.A0(net3455),
    .A1(net4022),
    .S(_05126_),
    .X(_01610_));
 sg13g2_mux2_1 _13988_ (.A0(net3408),
    .A1(net2759),
    .S(_05126_),
    .X(_01611_));
 sg13g2_mux2_1 _13989_ (.A0(net3366),
    .A1(net4195),
    .S(_05126_),
    .X(_01612_));
 sg13g2_mux2_1 _13990_ (.A0(net3320),
    .A1(net2854),
    .S(_05126_),
    .X(_01613_));
 sg13g2_mux2_1 _13991_ (.A0(net3269),
    .A1(net4413),
    .S(_05126_),
    .X(_01614_));
 sg13g2_nand2_1 _13992_ (.Y(_05127_),
    .A(net3084),
    .B(net3032));
 sg13g2_mux2_1 _13993_ (.A0(net3581),
    .A1(net4418),
    .S(_05127_),
    .X(_01615_));
 sg13g2_mux2_1 _13994_ (.A0(net3530),
    .A1(net4255),
    .S(net3012),
    .X(_01616_));
 sg13g2_mux2_1 _13995_ (.A0(net3483),
    .A1(net4371),
    .S(net3012),
    .X(_01617_));
 sg13g2_mux2_1 _13996_ (.A0(net3439),
    .A1(net4604),
    .S(net3012),
    .X(_01618_));
 sg13g2_mux2_1 _13997_ (.A0(net3394),
    .A1(net5056),
    .S(net3012),
    .X(_01619_));
 sg13g2_mux2_1 _13998_ (.A0(net3347),
    .A1(net4048),
    .S(net3012),
    .X(_01620_));
 sg13g2_mux2_1 _13999_ (.A0(net3303),
    .A1(net5115),
    .S(net3012),
    .X(_01621_));
 sg13g2_nor2_1 _14000_ (.A(net3256),
    .B(net3012),
    .Y(_05128_));
 sg13g2_a21oi_1 _14001_ (.A1(_02178_),
    .A2(net3012),
    .Y(_01622_),
    .B1(_05128_));
 sg13g2_and2_2 _14002_ (.A(net3077),
    .B(net3032),
    .X(_05129_));
 sg13g2_mux2_1 _14003_ (.A0(net2460),
    .A1(net3578),
    .S(_05129_),
    .X(_01623_));
 sg13g2_mux2_1 _14004_ (.A0(net2472),
    .A1(net3530),
    .S(_05129_),
    .X(_01624_));
 sg13g2_mux2_1 _14005_ (.A0(net2767),
    .A1(net3483),
    .S(_05129_),
    .X(_01625_));
 sg13g2_mux2_1 _14006_ (.A0(net2591),
    .A1(net3439),
    .S(_05129_),
    .X(_01626_));
 sg13g2_mux2_1 _14007_ (.A0(net2280),
    .A1(net3394),
    .S(_05129_),
    .X(_01627_));
 sg13g2_mux2_1 _14008_ (.A0(net2561),
    .A1(net3347),
    .S(_05129_),
    .X(_01628_));
 sg13g2_mux2_1 _14009_ (.A0(net2198),
    .A1(net3303),
    .S(_05129_),
    .X(_01629_));
 sg13g2_mux2_1 _14010_ (.A0(net2643),
    .A1(net3256),
    .S(_05129_),
    .X(_01630_));
 sg13g2_nand2_2 _14011_ (.Y(_05130_),
    .A(_02283_),
    .B(net3066));
 sg13g2_mux2_1 _14012_ (.A0(net3558),
    .A1(net4297),
    .S(_05130_),
    .X(_01631_));
 sg13g2_mux2_1 _14013_ (.A0(net3513),
    .A1(net2878),
    .S(_05130_),
    .X(_01632_));
 sg13g2_mux2_1 _14014_ (.A0(net3468),
    .A1(net4170),
    .S(_05130_),
    .X(_01633_));
 sg13g2_mux2_1 _14015_ (.A0(net3422),
    .A1(net4334),
    .S(_05130_),
    .X(_01634_));
 sg13g2_mux2_1 _14016_ (.A0(net3375),
    .A1(net2829),
    .S(_05130_),
    .X(_01635_));
 sg13g2_mux2_1 _14017_ (.A0(net3331),
    .A1(net2692),
    .S(_05130_),
    .X(_01636_));
 sg13g2_mux2_1 _14018_ (.A0(net3283),
    .A1(net2935),
    .S(_05130_),
    .X(_01637_));
 sg13g2_mux2_1 _14019_ (.A0(net3238),
    .A1(net2857),
    .S(_05130_),
    .X(_01638_));
 sg13g2_nor2_2 _14020_ (.A(_02298_),
    .B(_02381_),
    .Y(_05131_));
 sg13g2_mux2_1 _14021_ (.A0(net2396),
    .A1(net3558),
    .S(_05131_),
    .X(_01639_));
 sg13g2_mux2_1 _14022_ (.A0(net2664),
    .A1(net3513),
    .S(_05131_),
    .X(_01640_));
 sg13g2_mux2_1 _14023_ (.A0(net2431),
    .A1(net3467),
    .S(_05131_),
    .X(_01641_));
 sg13g2_mux2_1 _14024_ (.A0(net2237),
    .A1(net3422),
    .S(_05131_),
    .X(_01642_));
 sg13g2_mux2_1 _14025_ (.A0(net2653),
    .A1(net3375),
    .S(_05131_),
    .X(_01643_));
 sg13g2_mux2_1 _14026_ (.A0(net2618),
    .A1(net3331),
    .S(_05131_),
    .X(_01644_));
 sg13g2_mux2_1 _14027_ (.A0(net2263),
    .A1(net3283),
    .S(_05131_),
    .X(_01645_));
 sg13g2_mux2_1 _14028_ (.A0(net2423),
    .A1(net3238),
    .S(_05131_),
    .X(_01646_));
 sg13g2_nand2_2 _14029_ (.Y(_05132_),
    .A(net3036),
    .B(net3066));
 sg13g2_mux2_1 _14030_ (.A0(net3558),
    .A1(net5119),
    .S(_05132_),
    .X(_01647_));
 sg13g2_mux2_1 _14031_ (.A0(net3513),
    .A1(net2797),
    .S(_05132_),
    .X(_01648_));
 sg13g2_mux2_1 _14032_ (.A0(net3467),
    .A1(net5102),
    .S(_05132_),
    .X(_01649_));
 sg13g2_mux2_1 _14033_ (.A0(net3422),
    .A1(net4338),
    .S(_05132_),
    .X(_01650_));
 sg13g2_mux2_1 _14034_ (.A0(net3375),
    .A1(net2768),
    .S(_05132_),
    .X(_01651_));
 sg13g2_mux2_1 _14035_ (.A0(net3331),
    .A1(net2789),
    .S(_05132_),
    .X(_01652_));
 sg13g2_mux2_1 _14036_ (.A0(net3283),
    .A1(net5055),
    .S(_05132_),
    .X(_01653_));
 sg13g2_mux2_1 _14037_ (.A0(net3238),
    .A1(net4465),
    .S(_05132_),
    .X(_01654_));
 sg13g2_nand2_2 _14038_ (.Y(_05133_),
    .A(net3033),
    .B(net3066));
 sg13g2_mux2_1 _14039_ (.A0(net3558),
    .A1(net4875),
    .S(_05133_),
    .X(_01655_));
 sg13g2_mux2_1 _14040_ (.A0(net3513),
    .A1(net4311),
    .S(_05133_),
    .X(_01656_));
 sg13g2_mux2_1 _14041_ (.A0(net3467),
    .A1(net4609),
    .S(_05133_),
    .X(_01657_));
 sg13g2_mux2_1 _14042_ (.A0(net3422),
    .A1(net4206),
    .S(_05133_),
    .X(_01658_));
 sg13g2_mux2_1 _14043_ (.A0(net3375),
    .A1(net5129),
    .S(_05133_),
    .X(_01659_));
 sg13g2_mux2_1 _14044_ (.A0(net3331),
    .A1(net4381),
    .S(_05133_),
    .X(_01660_));
 sg13g2_mux2_1 _14045_ (.A0(net3283),
    .A1(net4759),
    .S(_05133_),
    .X(_01661_));
 sg13g2_mux2_1 _14046_ (.A0(net3238),
    .A1(net4961),
    .S(_05133_),
    .X(_01662_));
 sg13g2_nor2_2 _14047_ (.A(net3081),
    .B(_02381_),
    .Y(_05134_));
 sg13g2_mux2_1 _14048_ (.A0(net2649),
    .A1(net3558),
    .S(_05134_),
    .X(_01663_));
 sg13g2_mux2_1 _14049_ (.A0(net2268),
    .A1(net3515),
    .S(_05134_),
    .X(_01664_));
 sg13g2_mux2_1 _14050_ (.A0(net2246),
    .A1(net3467),
    .S(_05134_),
    .X(_01665_));
 sg13g2_mux2_1 _14051_ (.A0(net2369),
    .A1(net3422),
    .S(_05134_),
    .X(_01666_));
 sg13g2_mux2_1 _14052_ (.A0(net2132),
    .A1(net3375),
    .S(_05134_),
    .X(_01667_));
 sg13g2_mux2_1 _14053_ (.A0(net2159),
    .A1(net3331),
    .S(_05134_),
    .X(_01668_));
 sg13g2_mux2_1 _14054_ (.A0(net2492),
    .A1(net3283),
    .S(_05134_),
    .X(_01669_));
 sg13g2_mux2_1 _14055_ (.A0(net2230),
    .A1(net3238),
    .S(_05134_),
    .X(_01670_));
 sg13g2_nand2_2 _14056_ (.Y(_05135_),
    .A(_02346_),
    .B(net3066));
 sg13g2_mux2_1 _14057_ (.A0(net3558),
    .A1(net4186),
    .S(_05135_),
    .X(_01671_));
 sg13g2_mux2_1 _14058_ (.A0(net3513),
    .A1(net4673),
    .S(_05135_),
    .X(_01672_));
 sg13g2_mux2_1 _14059_ (.A0(net3468),
    .A1(net4069),
    .S(_05135_),
    .X(_01673_));
 sg13g2_mux2_1 _14060_ (.A0(net3422),
    .A1(net4667),
    .S(_05135_),
    .X(_01674_));
 sg13g2_mux2_1 _14061_ (.A0(net3375),
    .A1(net4491),
    .S(_05135_),
    .X(_01675_));
 sg13g2_mux2_1 _14062_ (.A0(net3331),
    .A1(net4834),
    .S(_05135_),
    .X(_01676_));
 sg13g2_mux2_1 _14063_ (.A0(net3283),
    .A1(net2949),
    .S(_05135_),
    .X(_01677_));
 sg13g2_mux2_1 _14064_ (.A0(net3239),
    .A1(net4695),
    .S(_05135_),
    .X(_01678_));
 sg13g2_nand2_2 _14065_ (.Y(_05136_),
    .A(net3066),
    .B(_02385_));
 sg13g2_mux2_1 _14066_ (.A0(net3558),
    .A1(net4101),
    .S(_05136_),
    .X(_01679_));
 sg13g2_mux2_1 _14067_ (.A0(net3513),
    .A1(net4818),
    .S(_05136_),
    .X(_01680_));
 sg13g2_mux2_1 _14068_ (.A0(net3468),
    .A1(net4462),
    .S(_05136_),
    .X(_01681_));
 sg13g2_mux2_1 _14069_ (.A0(net3423),
    .A1(net4592),
    .S(_05136_),
    .X(_01682_));
 sg13g2_mux2_1 _14070_ (.A0(net3375),
    .A1(net2763),
    .S(_05136_),
    .X(_01683_));
 sg13g2_mux2_1 _14071_ (.A0(net3331),
    .A1(net2863),
    .S(_05136_),
    .X(_01684_));
 sg13g2_mux2_1 _14072_ (.A0(net3283),
    .A1(net2798),
    .S(_05136_),
    .X(_01685_));
 sg13g2_mux2_1 _14073_ (.A0(net3239),
    .A1(net4036),
    .S(_05136_),
    .X(_01686_));
 sg13g2_nand2_2 _14074_ (.Y(_05137_),
    .A(_02297_),
    .B(_02311_));
 sg13g2_mux2_1 _14075_ (.A0(net3590),
    .A1(net4809),
    .S(_05137_),
    .X(_01687_));
 sg13g2_mux2_1 _14076_ (.A0(net3545),
    .A1(net4675),
    .S(_05137_),
    .X(_01688_));
 sg13g2_mux2_1 _14077_ (.A0(net3499),
    .A1(net4510),
    .S(_05137_),
    .X(_01689_));
 sg13g2_mux2_1 _14078_ (.A0(net3454),
    .A1(net4386),
    .S(_05137_),
    .X(_01690_));
 sg13g2_mux2_1 _14079_ (.A0(net3400),
    .A1(net4954),
    .S(_05137_),
    .X(_01691_));
 sg13g2_mux2_1 _14080_ (.A0(net3355),
    .A1(net4494),
    .S(_05137_),
    .X(_01692_));
 sg13g2_mux2_1 _14081_ (.A0(net3310),
    .A1(net5170),
    .S(_05137_),
    .X(_01693_));
 sg13g2_mux2_1 _14082_ (.A0(net3269),
    .A1(net5147),
    .S(_05137_),
    .X(_01694_));
 sg13g2_nor2_2 _14083_ (.A(_02338_),
    .B(_02381_),
    .Y(_05138_));
 sg13g2_mux2_1 _14084_ (.A0(net2368),
    .A1(net3559),
    .S(_05138_),
    .X(_01695_));
 sg13g2_mux2_1 _14085_ (.A0(net2321),
    .A1(net3515),
    .S(_05138_),
    .X(_01696_));
 sg13g2_mux2_1 _14086_ (.A0(net2320),
    .A1(net3467),
    .S(_05138_),
    .X(_01697_));
 sg13g2_mux2_1 _14087_ (.A0(net2690),
    .A1(net3423),
    .S(_05138_),
    .X(_01698_));
 sg13g2_mux2_1 _14088_ (.A0(net2573),
    .A1(net3376),
    .S(_05138_),
    .X(_01699_));
 sg13g2_mux2_1 _14089_ (.A0(net2847),
    .A1(net3329),
    .S(_05138_),
    .X(_01700_));
 sg13g2_mux2_1 _14090_ (.A0(net2411),
    .A1(net3285),
    .S(_05138_),
    .X(_01701_));
 sg13g2_mux2_1 _14091_ (.A0(net2533),
    .A1(net3239),
    .S(_05138_),
    .X(_01702_));
 sg13g2_nor2_2 _14092_ (.A(_02335_),
    .B(_02381_),
    .Y(_05139_));
 sg13g2_mux2_1 _14093_ (.A0(net2538),
    .A1(net3559),
    .S(_05139_),
    .X(_01703_));
 sg13g2_mux2_1 _14094_ (.A0(net2334),
    .A1(net3515),
    .S(_05139_),
    .X(_01704_));
 sg13g2_mux2_1 _14095_ (.A0(net2510),
    .A1(net3467),
    .S(_05139_),
    .X(_01705_));
 sg13g2_mux2_1 _14096_ (.A0(net2619),
    .A1(net3423),
    .S(_05139_),
    .X(_01706_));
 sg13g2_mux2_1 _14097_ (.A0(net2462),
    .A1(net3376),
    .S(_05139_),
    .X(_01707_));
 sg13g2_mux2_1 _14098_ (.A0(net2602),
    .A1(net3329),
    .S(_05139_),
    .X(_01708_));
 sg13g2_mux2_1 _14099_ (.A0(net2380),
    .A1(net3285),
    .S(_05139_),
    .X(_01709_));
 sg13g2_mux2_1 _14100_ (.A0(net2622),
    .A1(net3238),
    .S(_05139_),
    .X(_01710_));
 sg13g2_nand2_2 _14101_ (.Y(_05140_),
    .A(_02332_),
    .B(net3066));
 sg13g2_mux2_1 _14102_ (.A0(net3559),
    .A1(net4475),
    .S(_05140_),
    .X(_01711_));
 sg13g2_mux2_1 _14103_ (.A0(net3513),
    .A1(net5154),
    .S(_05140_),
    .X(_01712_));
 sg13g2_mux2_1 _14104_ (.A0(net3467),
    .A1(net4377),
    .S(_05140_),
    .X(_01713_));
 sg13g2_mux2_1 _14105_ (.A0(net3422),
    .A1(net4043),
    .S(_05140_),
    .X(_01714_));
 sg13g2_mux2_1 _14106_ (.A0(net3376),
    .A1(net4614),
    .S(_05140_),
    .X(_01715_));
 sg13g2_mux2_1 _14107_ (.A0(net3329),
    .A1(net4644),
    .S(_05140_),
    .X(_01716_));
 sg13g2_mux2_1 _14108_ (.A0(net3285),
    .A1(net4694),
    .S(_05140_),
    .X(_01717_));
 sg13g2_mux2_1 _14109_ (.A0(net3238),
    .A1(net4015),
    .S(_05140_),
    .X(_01718_));
 sg13g2_nand2_2 _14110_ (.Y(_05141_),
    .A(_02328_),
    .B(net3066));
 sg13g2_mux2_1 _14111_ (.A0(net3559),
    .A1(net4318),
    .S(_05141_),
    .X(_01719_));
 sg13g2_mux2_1 _14112_ (.A0(net3514),
    .A1(net3008),
    .S(_05141_),
    .X(_01720_));
 sg13g2_mux2_1 _14113_ (.A0(net3467),
    .A1(net4904),
    .S(_05141_),
    .X(_01721_));
 sg13g2_mux2_1 _14114_ (.A0(net3422),
    .A1(net4876),
    .S(_05141_),
    .X(_01722_));
 sg13g2_mux2_1 _14115_ (.A0(net3376),
    .A1(net4940),
    .S(_05141_),
    .X(_01723_));
 sg13g2_mux2_1 _14116_ (.A0(net3329),
    .A1(net4086),
    .S(_05141_),
    .X(_01724_));
 sg13g2_mux2_1 _14117_ (.A0(net3285),
    .A1(net4782),
    .S(_05141_),
    .X(_01725_));
 sg13g2_mux2_1 _14118_ (.A0(net3238),
    .A1(net4816),
    .S(_05141_),
    .X(_01726_));
 sg13g2_nand2_2 _14119_ (.Y(_05142_),
    .A(net3072),
    .B(_02379_));
 sg13g2_mux2_1 _14120_ (.A0(net3561),
    .A1(net4059),
    .S(_05142_),
    .X(_01727_));
 sg13g2_mux2_1 _14121_ (.A0(net3514),
    .A1(net4126),
    .S(_05142_),
    .X(_01728_));
 sg13g2_mux2_1 _14122_ (.A0(net3469),
    .A1(net2774),
    .S(_05142_),
    .X(_01729_));
 sg13g2_mux2_1 _14123_ (.A0(net3427),
    .A1(net4856),
    .S(_05142_),
    .X(_01730_));
 sg13g2_mux2_1 _14124_ (.A0(net3376),
    .A1(net5111),
    .S(_05142_),
    .X(_01731_));
 sg13g2_mux2_1 _14125_ (.A0(net3329),
    .A1(net2597),
    .S(_05142_),
    .X(_01732_));
 sg13g2_mux2_1 _14126_ (.A0(net3285),
    .A1(net2823),
    .S(_05142_),
    .X(_01733_));
 sg13g2_mux2_1 _14127_ (.A0(net3243),
    .A1(net4738),
    .S(_05142_),
    .X(_01734_));
 sg13g2_and3_2 _14128_ (.X(_05143_),
    .A(net3041),
    .B(net3073),
    .C(_02379_));
 sg13g2_mux2_1 _14129_ (.A0(net2802),
    .A1(net3564),
    .S(_05143_),
    .X(_01735_));
 sg13g2_mux2_1 _14130_ (.A0(net2285),
    .A1(net3514),
    .S(_05143_),
    .X(_01736_));
 sg13g2_mux2_1 _14131_ (.A0(net2544),
    .A1(net3472),
    .S(_05143_),
    .X(_01737_));
 sg13g2_mux2_1 _14132_ (.A0(net2801),
    .A1(net3424),
    .S(_05143_),
    .X(_01738_));
 sg13g2_mux2_1 _14133_ (.A0(net2518),
    .A1(net3376),
    .S(_05143_),
    .X(_01739_));
 sg13g2_mux2_1 _14134_ (.A0(net2840),
    .A1(net3329),
    .S(_05143_),
    .X(_01740_));
 sg13g2_mux2_1 _14135_ (.A0(net2723),
    .A1(net3285),
    .S(_05143_),
    .X(_01741_));
 sg13g2_mux2_1 _14136_ (.A0(net2541),
    .A1(net3240),
    .S(_05143_),
    .X(_01742_));
 sg13g2_nor2_2 _14137_ (.A(_02249_),
    .B(_02381_),
    .Y(_05144_));
 sg13g2_mux2_1 _14138_ (.A0(net2509),
    .A1(net3561),
    .S(_05144_),
    .X(_01743_));
 sg13g2_mux2_1 _14139_ (.A0(net2318),
    .A1(net3514),
    .S(_05144_),
    .X(_01744_));
 sg13g2_mux2_1 _14140_ (.A0(net2200),
    .A1(net3469),
    .S(_05144_),
    .X(_01745_));
 sg13g2_mux2_1 _14141_ (.A0(net2679),
    .A1(net3424),
    .S(_05144_),
    .X(_01746_));
 sg13g2_mux2_1 _14142_ (.A0(net2377),
    .A1(net3376),
    .S(_05144_),
    .X(_01747_));
 sg13g2_mux2_1 _14143_ (.A0(net2150),
    .A1(net3329),
    .S(_05144_),
    .X(_01748_));
 sg13g2_mux2_1 _14144_ (.A0(net2145),
    .A1(net3285),
    .S(_05144_),
    .X(_01749_));
 sg13g2_mux2_1 _14145_ (.A0(net2471),
    .A1(net3240),
    .S(_05144_),
    .X(_01750_));
 sg13g2_nor2_2 _14146_ (.A(net3076),
    .B(_02381_),
    .Y(_05145_));
 sg13g2_mux2_1 _14147_ (.A0(net2447),
    .A1(net3561),
    .S(_05145_),
    .X(_01751_));
 sg13g2_mux2_1 _14148_ (.A0(net2325),
    .A1(net3514),
    .S(_05145_),
    .X(_01752_));
 sg13g2_mux2_1 _14149_ (.A0(net2507),
    .A1(net3469),
    .S(_05145_),
    .X(_01753_));
 sg13g2_mux2_1 _14150_ (.A0(net2640),
    .A1(net3424),
    .S(_05145_),
    .X(_01754_));
 sg13g2_mux2_1 _14151_ (.A0(net2719),
    .A1(net3376),
    .S(_05145_),
    .X(_01755_));
 sg13g2_mux2_1 _14152_ (.A0(net2677),
    .A1(net3329),
    .S(_05145_),
    .X(_01756_));
 sg13g2_mux2_1 _14153_ (.A0(net2505),
    .A1(net3285),
    .S(_05145_),
    .X(_01757_));
 sg13g2_mux2_1 _14154_ (.A0(net2265),
    .A1(net3240),
    .S(_05145_),
    .X(_01758_));
 sg13g2_nand2_2 _14155_ (.Y(_05146_),
    .A(net3079),
    .B(_02300_));
 sg13g2_mux2_1 _14156_ (.A0(net3560),
    .A1(net4469),
    .S(_05146_),
    .X(_01759_));
 sg13g2_mux2_1 _14157_ (.A0(net3516),
    .A1(net4523),
    .S(_05146_),
    .X(_01760_));
 sg13g2_mux2_1 _14158_ (.A0(net3470),
    .A1(net2820),
    .S(_05146_),
    .X(_01761_));
 sg13g2_mux2_1 _14159_ (.A0(net3425),
    .A1(net4808),
    .S(_05146_),
    .X(_01762_));
 sg13g2_mux2_1 _14160_ (.A0(net3377),
    .A1(net2725),
    .S(_05146_),
    .X(_01763_));
 sg13g2_mux2_1 _14161_ (.A0(net3332),
    .A1(net2830),
    .S(_05146_),
    .X(_01764_));
 sg13g2_mux2_1 _14162_ (.A0(net3284),
    .A1(net4340),
    .S(_05146_),
    .X(_01765_));
 sg13g2_mux2_1 _14163_ (.A0(net3241),
    .A1(net2890),
    .S(_05146_),
    .X(_01766_));
 sg13g2_nand2_2 _14164_ (.Y(_05147_),
    .A(_02277_),
    .B(net3034));
 sg13g2_mux2_1 _14165_ (.A0(net3595),
    .A1(net4802),
    .S(_05147_),
    .X(_01767_));
 sg13g2_mux2_1 _14166_ (.A0(net3549),
    .A1(net4859),
    .S(_05147_),
    .X(_01768_));
 sg13g2_mux2_1 _14167_ (.A0(net3503),
    .A1(net2887),
    .S(_05147_),
    .X(_01769_));
 sg13g2_mux2_1 _14168_ (.A0(net3456),
    .A1(net2839),
    .S(_05147_),
    .X(_01770_));
 sg13g2_mux2_1 _14169_ (.A0(net3410),
    .A1(net2604),
    .S(_05147_),
    .X(_01771_));
 sg13g2_mux2_1 _14170_ (.A0(net3367),
    .A1(net2973),
    .S(_05147_),
    .X(_01772_));
 sg13g2_mux2_1 _14171_ (.A0(net3321),
    .A1(net2637),
    .S(_05147_),
    .X(_01773_));
 sg13g2_mux2_1 _14172_ (.A0(net3271),
    .A1(net2760),
    .S(_05147_),
    .X(_01774_));
 sg13g2_nand2_2 _14173_ (.Y(_05148_),
    .A(net3036),
    .B(net3078));
 sg13g2_mux2_1 _14174_ (.A0(net3560),
    .A1(net4372),
    .S(_05148_),
    .X(_01775_));
 sg13g2_mux2_1 _14175_ (.A0(net3516),
    .A1(net4794),
    .S(_05148_),
    .X(_01776_));
 sg13g2_mux2_1 _14176_ (.A0(net3470),
    .A1(net2968),
    .S(_05148_),
    .X(_01777_));
 sg13g2_mux2_1 _14177_ (.A0(net3425),
    .A1(net3001),
    .S(_05148_),
    .X(_01778_));
 sg13g2_mux2_1 _14178_ (.A0(net3377),
    .A1(net2888),
    .S(_05148_),
    .X(_01779_));
 sg13g2_mux2_1 _14179_ (.A0(net3332),
    .A1(net2817),
    .S(_05148_),
    .X(_01780_));
 sg13g2_mux2_1 _14180_ (.A0(net3284),
    .A1(net4573),
    .S(_05148_),
    .X(_01781_));
 sg13g2_mux2_1 _14181_ (.A0(net3241),
    .A1(net4077),
    .S(_05148_),
    .X(_01782_));
 sg13g2_nand2_2 _14182_ (.Y(_05149_),
    .A(net3078),
    .B(net3033));
 sg13g2_mux2_1 _14183_ (.A0(net3560),
    .A1(net4155),
    .S(_05149_),
    .X(_01783_));
 sg13g2_mux2_1 _14184_ (.A0(net3516),
    .A1(net4024),
    .S(_05149_),
    .X(_01784_));
 sg13g2_mux2_1 _14185_ (.A0(net3470),
    .A1(net4344),
    .S(_05149_),
    .X(_01785_));
 sg13g2_mux2_1 _14186_ (.A0(net3425),
    .A1(net4871),
    .S(_05149_),
    .X(_01786_));
 sg13g2_mux2_1 _14187_ (.A0(net3377),
    .A1(net4591),
    .S(_05149_),
    .X(_01787_));
 sg13g2_mux2_1 _14188_ (.A0(net3332),
    .A1(net4426),
    .S(_05149_),
    .X(_01788_));
 sg13g2_mux2_1 _14189_ (.A0(net3284),
    .A1(net4744),
    .S(_05149_),
    .X(_01789_));
 sg13g2_mux2_1 _14190_ (.A0(net3241),
    .A1(net4277),
    .S(_05149_),
    .X(_01790_));
 sg13g2_nor2_2 _14191_ (.A(net3081),
    .B(_02301_),
    .Y(_05150_));
 sg13g2_mux2_1 _14192_ (.A0(net2353),
    .A1(net3561),
    .S(_05150_),
    .X(_01791_));
 sg13g2_mux2_1 _14193_ (.A0(net2308),
    .A1(net3517),
    .S(_05150_),
    .X(_01792_));
 sg13g2_mux2_1 _14194_ (.A0(net2614),
    .A1(net3471),
    .S(_05150_),
    .X(_01793_));
 sg13g2_mux2_1 _14195_ (.A0(net2504),
    .A1(net3426),
    .S(_05150_),
    .X(_01794_));
 sg13g2_mux2_1 _14196_ (.A0(net2143),
    .A1(net3378),
    .S(_05150_),
    .X(_01795_));
 sg13g2_mux2_1 _14197_ (.A0(net2149),
    .A1(net3335),
    .S(_05150_),
    .X(_01796_));
 sg13g2_mux2_1 _14198_ (.A0(net2229),
    .A1(net3286),
    .S(_05150_),
    .X(_01797_));
 sg13g2_mux2_1 _14199_ (.A0(net2210),
    .A1(net3242),
    .S(_05150_),
    .X(_01798_));
 sg13g2_nand2_2 _14200_ (.Y(_05151_),
    .A(net3078),
    .B(_02346_));
 sg13g2_mux2_1 _14201_ (.A0(net3561),
    .A1(net4515),
    .S(_05151_),
    .X(_01799_));
 sg13g2_mux2_1 _14202_ (.A0(net3517),
    .A1(net4973),
    .S(_05151_),
    .X(_01800_));
 sg13g2_mux2_1 _14203_ (.A0(net3471),
    .A1(net2893),
    .S(_05151_),
    .X(_01801_));
 sg13g2_mux2_1 _14204_ (.A0(net3426),
    .A1(net4434),
    .S(_05151_),
    .X(_01802_));
 sg13g2_mux2_1 _14205_ (.A0(net3378),
    .A1(net4864),
    .S(_05151_),
    .X(_01803_));
 sg13g2_mux2_1 _14206_ (.A0(net3334),
    .A1(net4390),
    .S(_05151_),
    .X(_01804_));
 sg13g2_mux2_1 _14207_ (.A0(net3286),
    .A1(net4193),
    .S(_05151_),
    .X(_01805_));
 sg13g2_mux2_1 _14208_ (.A0(net3242),
    .A1(net4956),
    .S(_05151_),
    .X(_01806_));
 sg13g2_nand2_2 _14209_ (.Y(_05152_),
    .A(net3078),
    .B(_02385_));
 sg13g2_mux2_1 _14210_ (.A0(net3561),
    .A1(net5060),
    .S(_05152_),
    .X(_01807_));
 sg13g2_mux2_1 _14211_ (.A0(net3517),
    .A1(net4736),
    .S(_05152_),
    .X(_01808_));
 sg13g2_mux2_1 _14212_ (.A0(net3471),
    .A1(net5034),
    .S(_05152_),
    .X(_01809_));
 sg13g2_mux2_1 _14213_ (.A0(net3425),
    .A1(net4798),
    .S(_05152_),
    .X(_01810_));
 sg13g2_mux2_1 _14214_ (.A0(net3378),
    .A1(net2859),
    .S(_05152_),
    .X(_01811_));
 sg13g2_mux2_1 _14215_ (.A0(net3334),
    .A1(net2746),
    .S(_05152_),
    .X(_01812_));
 sg13g2_mux2_1 _14216_ (.A0(net3286),
    .A1(net4724),
    .S(_05152_),
    .X(_01813_));
 sg13g2_mux2_1 _14217_ (.A0(net3242),
    .A1(net4682),
    .S(_05152_),
    .X(_01814_));
 sg13g2_nand2_2 _14218_ (.Y(_05153_),
    .A(net3078),
    .B(net3049));
 sg13g2_mux2_1 _14219_ (.A0(net3561),
    .A1(net2991),
    .S(_05153_),
    .X(_01815_));
 sg13g2_mux2_1 _14220_ (.A0(net3517),
    .A1(net4528),
    .S(_05153_),
    .X(_01816_));
 sg13g2_mux2_1 _14221_ (.A0(net3471),
    .A1(net4501),
    .S(_05153_),
    .X(_01817_));
 sg13g2_mux2_1 _14222_ (.A0(net3425),
    .A1(net5047),
    .S(_05153_),
    .X(_01818_));
 sg13g2_mux2_1 _14223_ (.A0(net3378),
    .A1(net5054),
    .S(_05153_),
    .X(_01819_));
 sg13g2_mux2_1 _14224_ (.A0(net3334),
    .A1(net4866),
    .S(_05153_),
    .X(_01820_));
 sg13g2_mux2_1 _14225_ (.A0(net3286),
    .A1(net4098),
    .S(_05153_),
    .X(_01821_));
 sg13g2_mux2_1 _14226_ (.A0(net3242),
    .A1(net4787),
    .S(_05153_),
    .X(_01822_));
 sg13g2_nand2_2 _14227_ (.Y(_05154_),
    .A(_02299_),
    .B(_02339_));
 sg13g2_mux2_1 _14228_ (.A0(net3562),
    .A1(net4497),
    .S(_05154_),
    .X(_01823_));
 sg13g2_mux2_1 _14229_ (.A0(net3516),
    .A1(net2728),
    .S(_05154_),
    .X(_01824_));
 sg13g2_mux2_1 _14230_ (.A0(net3478),
    .A1(net2773),
    .S(_05154_),
    .X(_01825_));
 sg13g2_mux2_1 _14231_ (.A0(net3432),
    .A1(net4144),
    .S(_05154_),
    .X(_01826_));
 sg13g2_mux2_1 _14232_ (.A0(net3377),
    .A1(net4976),
    .S(_05154_),
    .X(_01827_));
 sg13g2_mux2_1 _14233_ (.A0(net3333),
    .A1(net2963),
    .S(_05154_),
    .X(_01828_));
 sg13g2_mux2_1 _14234_ (.A0(net3288),
    .A1(net4097),
    .S(_05154_),
    .X(_01829_));
 sg13g2_mux2_1 _14235_ (.A0(net3241),
    .A1(net5105),
    .S(_05154_),
    .X(_01830_));
 sg13g2_nand2_2 _14236_ (.Y(_05155_),
    .A(_02300_),
    .B(net3070));
 sg13g2_mux2_1 _14237_ (.A0(net3562),
    .A1(net4223),
    .S(_05155_),
    .X(_01831_));
 sg13g2_mux2_1 _14238_ (.A0(net3516),
    .A1(net4922),
    .S(_05155_),
    .X(_01832_));
 sg13g2_mux2_1 _14239_ (.A0(net3478),
    .A1(net4582),
    .S(_05155_),
    .X(_01833_));
 sg13g2_mux2_1 _14240_ (.A0(net3432),
    .A1(net4295),
    .S(_05155_),
    .X(_01834_));
 sg13g2_mux2_1 _14241_ (.A0(net3379),
    .A1(net5074),
    .S(_05155_),
    .X(_01835_));
 sg13g2_mux2_1 _14242_ (.A0(net3333),
    .A1(net4428),
    .S(_05155_),
    .X(_01836_));
 sg13g2_mux2_1 _14243_ (.A0(net3288),
    .A1(net4519),
    .S(_05155_),
    .X(_01837_));
 sg13g2_mux2_1 _14244_ (.A0(net3241),
    .A1(net4425),
    .S(_05155_),
    .X(_01838_));
 sg13g2_nand2_2 _14245_ (.Y(_05156_),
    .A(net3078),
    .B(_02332_));
 sg13g2_mux2_1 _14246_ (.A0(net3562),
    .A1(net2951),
    .S(_05156_),
    .X(_01839_));
 sg13g2_mux2_1 _14247_ (.A0(net3516),
    .A1(net2745),
    .S(_05156_),
    .X(_01840_));
 sg13g2_mux2_1 _14248_ (.A0(net3478),
    .A1(net4235),
    .S(_05156_),
    .X(_01841_));
 sg13g2_mux2_1 _14249_ (.A0(net3432),
    .A1(net4080),
    .S(_05156_),
    .X(_01842_));
 sg13g2_mux2_1 _14250_ (.A0(net3377),
    .A1(net4972),
    .S(_05156_),
    .X(_01843_));
 sg13g2_mux2_1 _14251_ (.A0(net3333),
    .A1(net2936),
    .S(_05156_),
    .X(_01844_));
 sg13g2_mux2_1 _14252_ (.A0(net3288),
    .A1(net4657),
    .S(_05156_),
    .X(_01845_));
 sg13g2_mux2_1 _14253_ (.A0(net3241),
    .A1(net4040),
    .S(_05156_),
    .X(_01846_));
 sg13g2_nand2_2 _14254_ (.Y(_05157_),
    .A(net3069),
    .B(net3035));
 sg13g2_mux2_1 _14255_ (.A0(net3595),
    .A1(net4033),
    .S(_05157_),
    .X(_01847_));
 sg13g2_mux2_1 _14256_ (.A0(net3549),
    .A1(net4014),
    .S(_05157_),
    .X(_01848_));
 sg13g2_mux2_1 _14257_ (.A0(net3502),
    .A1(net4918),
    .S(_05157_),
    .X(_01849_));
 sg13g2_mux2_1 _14258_ (.A0(net3456),
    .A1(net5171),
    .S(_05157_),
    .X(_01850_));
 sg13g2_mux2_1 _14259_ (.A0(net3410),
    .A1(net4889),
    .S(_05157_),
    .X(_01851_));
 sg13g2_mux2_1 _14260_ (.A0(net3367),
    .A1(net4107),
    .S(_05157_),
    .X(_01852_));
 sg13g2_mux2_1 _14261_ (.A0(net3321),
    .A1(net5027),
    .S(_05157_),
    .X(_01853_));
 sg13g2_mux2_1 _14262_ (.A0(net3271),
    .A1(net5156),
    .S(_05157_),
    .X(_01854_));
 sg13g2_nand2_2 _14263_ (.Y(_05158_),
    .A(_02299_),
    .B(net3072));
 sg13g2_mux2_1 _14264_ (.A0(net3562),
    .A1(net4423),
    .S(_05158_),
    .X(_01855_));
 sg13g2_mux2_1 _14265_ (.A0(net3517),
    .A1(net4931),
    .S(_05158_),
    .X(_01856_));
 sg13g2_mux2_1 _14266_ (.A0(net3479),
    .A1(net4154),
    .S(_05158_),
    .X(_01857_));
 sg13g2_mux2_1 _14267_ (.A0(net3433),
    .A1(net5132),
    .S(_05158_),
    .X(_01858_));
 sg13g2_mux2_1 _14268_ (.A0(net3378),
    .A1(net2865),
    .S(_05158_),
    .X(_01859_));
 sg13g2_mux2_1 _14269_ (.A0(net3332),
    .A1(net2980),
    .S(_05158_),
    .X(_01860_));
 sg13g2_mux2_1 _14270_ (.A0(net3288),
    .A1(net4936),
    .S(_05158_),
    .X(_01861_));
 sg13g2_mux2_1 _14271_ (.A0(net3250),
    .A1(net2799),
    .S(_05158_),
    .X(_01862_));
 sg13g2_nand2_2 _14272_ (.Y(_05159_),
    .A(_02300_),
    .B(net3073));
 sg13g2_mux2_1 _14273_ (.A0(net3562),
    .A1(net4052),
    .S(_05159_),
    .X(_01863_));
 sg13g2_mux2_1 _14274_ (.A0(net3518),
    .A1(net5149),
    .S(_05159_),
    .X(_01864_));
 sg13g2_mux2_1 _14275_ (.A0(net3479),
    .A1(net4068),
    .S(_05159_),
    .X(_01865_));
 sg13g2_mux2_1 _14276_ (.A0(net3433),
    .A1(net4457),
    .S(_05159_),
    .X(_01866_));
 sg13g2_mux2_1 _14277_ (.A0(net3378),
    .A1(net4658),
    .S(_05159_),
    .X(_01867_));
 sg13g2_mux2_1 _14278_ (.A0(net3332),
    .A1(net5012),
    .S(_05159_),
    .X(_01868_));
 sg13g2_mux2_1 _14279_ (.A0(net3288),
    .A1(net4947),
    .S(_05159_),
    .X(_01869_));
 sg13g2_mux2_1 _14280_ (.A0(net3250),
    .A1(net5104),
    .S(_05159_),
    .X(_01870_));
 sg13g2_nand2_1 _14281_ (.Y(_05160_),
    .A(net3084),
    .B(_02300_));
 sg13g2_mux2_1 _14282_ (.A0(net3562),
    .A1(net2950),
    .S(net3011),
    .X(_01871_));
 sg13g2_mux2_1 _14283_ (.A0(net3519),
    .A1(net2901),
    .S(net3011),
    .X(_01872_));
 sg13g2_mux2_1 _14284_ (.A0(net3479),
    .A1(net4499),
    .S(net3011),
    .X(_01873_));
 sg13g2_mux2_1 _14285_ (.A0(net3433),
    .A1(net4117),
    .S(_05160_),
    .X(_01874_));
 sg13g2_mux2_1 _14286_ (.A0(net3377),
    .A1(net2738),
    .S(net3011),
    .X(_01875_));
 sg13g2_mux2_1 _14287_ (.A0(net3332),
    .A1(net4757),
    .S(net3011),
    .X(_01876_));
 sg13g2_mux2_1 _14288_ (.A0(net3288),
    .A1(net5032),
    .S(net3011),
    .X(_01877_));
 sg13g2_nor2_1 _14289_ (.A(net3242),
    .B(net3011),
    .Y(_05161_));
 sg13g2_a21oi_1 _14290_ (.A1(_02180_),
    .A2(net3011),
    .Y(_01878_),
    .B1(_05161_));
 sg13g2_nor2_2 _14291_ (.A(_02301_),
    .B(net3076),
    .Y(_05162_));
 sg13g2_mux2_1 _14292_ (.A0(net2567),
    .A1(net3562),
    .S(_05162_),
    .X(_01879_));
 sg13g2_mux2_1 _14293_ (.A0(net2448),
    .A1(net3517),
    .S(_05162_),
    .X(_01880_));
 sg13g2_mux2_1 _14294_ (.A0(net2425),
    .A1(net3479),
    .S(_05162_),
    .X(_01881_));
 sg13g2_mux2_1 _14295_ (.A0(net2304),
    .A1(net3433),
    .S(_05162_),
    .X(_01882_));
 sg13g2_mux2_1 _14296_ (.A0(net2613),
    .A1(net3377),
    .S(_05162_),
    .X(_01883_));
 sg13g2_mux2_1 _14297_ (.A0(net2224),
    .A1(net3332),
    .S(_05162_),
    .X(_01884_));
 sg13g2_mux2_1 _14298_ (.A0(net2342),
    .A1(net3288),
    .S(_05162_),
    .X(_01885_));
 sg13g2_mux2_1 _14299_ (.A0(net2261),
    .A1(net3242),
    .S(_05162_),
    .X(_01886_));
 sg13g2_nand2_2 _14300_ (.Y(_05163_),
    .A(net3079),
    .B(_05007_));
 sg13g2_mux2_1 _14301_ (.A0(net3583),
    .A1(net2785),
    .S(_05163_),
    .X(_01887_));
 sg13g2_mux2_1 _14302_ (.A0(net3535),
    .A1(net4414),
    .S(_05163_),
    .X(_01888_));
 sg13g2_mux2_1 _14303_ (.A0(net3490),
    .A1(net4216),
    .S(_05163_),
    .X(_01889_));
 sg13g2_mux2_1 _14304_ (.A0(net3444),
    .A1(net4013),
    .S(_05163_),
    .X(_01890_));
 sg13g2_mux2_1 _14305_ (.A0(net3398),
    .A1(net2838),
    .S(_05163_),
    .X(_01891_));
 sg13g2_mux2_1 _14306_ (.A0(net3353),
    .A1(net4032),
    .S(_05163_),
    .X(_01892_));
 sg13g2_mux2_1 _14307_ (.A0(net3309),
    .A1(net2979),
    .S(_05163_),
    .X(_01893_));
 sg13g2_mux2_1 _14308_ (.A0(net3259),
    .A1(net4689),
    .S(_05163_),
    .X(_01894_));
 sg13g2_nor2_2 _14309_ (.A(_02298_),
    .B(_05008_),
    .Y(_05164_));
 sg13g2_mux2_1 _14310_ (.A0(net2566),
    .A1(net3583),
    .S(_05164_),
    .X(_01895_));
 sg13g2_mux2_1 _14311_ (.A0(net2326),
    .A1(net3535),
    .S(_05164_),
    .X(_01896_));
 sg13g2_mux2_1 _14312_ (.A0(net2451),
    .A1(net3490),
    .S(_05164_),
    .X(_01897_));
 sg13g2_mux2_1 _14313_ (.A0(net2593),
    .A1(net3444),
    .S(_05164_),
    .X(_01898_));
 sg13g2_mux2_1 _14314_ (.A0(net2652),
    .A1(net3398),
    .S(_05164_),
    .X(_01899_));
 sg13g2_mux2_1 _14315_ (.A0(net2627),
    .A1(net3353),
    .S(_05164_),
    .X(_01900_));
 sg13g2_mux2_1 _14316_ (.A0(net2466),
    .A1(net3309),
    .S(_05164_),
    .X(_01901_));
 sg13g2_mux2_1 _14317_ (.A0(net2532),
    .A1(net3259),
    .S(_05164_),
    .X(_01902_));
 sg13g2_nand2_2 _14318_ (.Y(_05165_),
    .A(net3036),
    .B(net3051));
 sg13g2_mux2_1 _14319_ (.A0(net3583),
    .A1(net2858),
    .S(_05165_),
    .X(_01903_));
 sg13g2_mux2_1 _14320_ (.A0(net3535),
    .A1(net4460),
    .S(_05165_),
    .X(_01904_));
 sg13g2_mux2_1 _14321_ (.A0(net3490),
    .A1(net4899),
    .S(_05165_),
    .X(_01905_));
 sg13g2_mux2_1 _14322_ (.A0(net3443),
    .A1(net4239),
    .S(_05165_),
    .X(_01906_));
 sg13g2_mux2_1 _14323_ (.A0(net3401),
    .A1(net2822),
    .S(_05165_),
    .X(_01907_));
 sg13g2_mux2_1 _14324_ (.A0(net3353),
    .A1(net2853),
    .S(_05165_),
    .X(_01908_));
 sg13g2_mux2_1 _14325_ (.A0(net3309),
    .A1(net4637),
    .S(_05165_),
    .X(_01909_));
 sg13g2_mux2_1 _14326_ (.A0(net3259),
    .A1(net5018),
    .S(_05165_),
    .X(_01910_));
 sg13g2_nand2_2 _14327_ (.Y(_05166_),
    .A(_02349_),
    .B(_05007_));
 sg13g2_mux2_1 _14328_ (.A0(net3583),
    .A1(net5029),
    .S(_05166_),
    .X(_01911_));
 sg13g2_mux2_1 _14329_ (.A0(net3535),
    .A1(net4620),
    .S(_05166_),
    .X(_01912_));
 sg13g2_mux2_1 _14330_ (.A0(net3490),
    .A1(net5145),
    .S(_05166_),
    .X(_01913_));
 sg13g2_mux2_1 _14331_ (.A0(net3443),
    .A1(net4732),
    .S(_05166_),
    .X(_01914_));
 sg13g2_mux2_1 _14332_ (.A0(net3398),
    .A1(net4830),
    .S(_05166_),
    .X(_01915_));
 sg13g2_mux2_1 _14333_ (.A0(net3353),
    .A1(net5041),
    .S(_05166_),
    .X(_01916_));
 sg13g2_mux2_1 _14334_ (.A0(net3309),
    .A1(net4152),
    .S(_05166_),
    .X(_01917_));
 sg13g2_mux2_1 _14335_ (.A0(net3259),
    .A1(net5077),
    .S(_05166_),
    .X(_01918_));
 sg13g2_nor2_2 _14336_ (.A(net3081),
    .B(_05008_),
    .Y(_05167_));
 sg13g2_mux2_1 _14337_ (.A0(net2188),
    .A1(net3582),
    .S(_05167_),
    .X(_01919_));
 sg13g2_mux2_1 _14338_ (.A0(net2250),
    .A1(net3536),
    .S(_05167_),
    .X(_01920_));
 sg13g2_mux2_1 _14339_ (.A0(net2623),
    .A1(net3493),
    .S(_05167_),
    .X(_01921_));
 sg13g2_mux2_1 _14340_ (.A0(net2165),
    .A1(net3443),
    .S(_05167_),
    .X(_01922_));
 sg13g2_mux2_1 _14341_ (.A0(net2142),
    .A1(net3401),
    .S(_05167_),
    .X(_01923_));
 sg13g2_mux2_1 _14342_ (.A0(net2151),
    .A1(net3355),
    .S(_05167_),
    .X(_01924_));
 sg13g2_mux2_1 _14343_ (.A0(net2202),
    .A1(net3310),
    .S(_05167_),
    .X(_01925_));
 sg13g2_mux2_1 _14344_ (.A0(net2329),
    .A1(net3262),
    .S(_05167_),
    .X(_01926_));
 sg13g2_nand2_1 _14345_ (.Y(_05168_),
    .A(net3035),
    .B(net3065));
 sg13g2_mux2_1 _14346_ (.A0(net3595),
    .A1(net4496),
    .S(net3010),
    .X(_01927_));
 sg13g2_mux2_1 _14347_ (.A0(net3549),
    .A1(net4215),
    .S(_05168_),
    .X(_01928_));
 sg13g2_mux2_1 _14348_ (.A0(net3502),
    .A1(net4435),
    .S(net3010),
    .X(_01929_));
 sg13g2_mux2_1 _14349_ (.A0(net3456),
    .A1(net2632),
    .S(net3010),
    .X(_01930_));
 sg13g2_mux2_1 _14350_ (.A0(net3410),
    .A1(net2699),
    .S(net3010),
    .X(_01931_));
 sg13g2_mux2_1 _14351_ (.A0(net3367),
    .A1(net4137),
    .S(net3010),
    .X(_01932_));
 sg13g2_mux2_1 _14352_ (.A0(net3321),
    .A1(net2848),
    .S(net3010),
    .X(_01933_));
 sg13g2_nor2_1 _14353_ (.A(net3271),
    .B(net3010),
    .Y(_05169_));
 sg13g2_a21oi_1 _14354_ (.A1(_02169_),
    .A2(net3010),
    .Y(_01934_),
    .B1(_05169_));
 sg13g2_nand2_2 _14355_ (.Y(_05170_),
    .A(net3065),
    .B(_05007_));
 sg13g2_mux2_1 _14356_ (.A0(net3583),
    .A1(net4548),
    .S(_05170_),
    .X(_01935_));
 sg13g2_mux2_1 _14357_ (.A0(net3535),
    .A1(net2948),
    .S(_05170_),
    .X(_01936_));
 sg13g2_mux2_1 _14358_ (.A0(net3490),
    .A1(net2644),
    .S(_05170_),
    .X(_01937_));
 sg13g2_mux2_1 _14359_ (.A0(net3443),
    .A1(net4343),
    .S(_05170_),
    .X(_01938_));
 sg13g2_mux2_1 _14360_ (.A0(net3398),
    .A1(net2821),
    .S(_05170_),
    .X(_01939_));
 sg13g2_mux2_1 _14361_ (.A0(net3353),
    .A1(net2716),
    .S(_05170_),
    .X(_01940_));
 sg13g2_mux2_1 _14362_ (.A0(net3309),
    .A1(net4621),
    .S(_05170_),
    .X(_01941_));
 sg13g2_mux2_1 _14363_ (.A0(net3259),
    .A1(net4060),
    .S(_05170_),
    .X(_01942_));
 sg13g2_nand2_2 _14364_ (.Y(_05171_),
    .A(net3049),
    .B(net3051));
 sg13g2_mux2_1 _14365_ (.A0(net3583),
    .A1(net2937),
    .S(_05171_),
    .X(_01943_));
 sg13g2_mux2_1 _14366_ (.A0(net3535),
    .A1(net2989),
    .S(_05171_),
    .X(_01944_));
 sg13g2_mux2_1 _14367_ (.A0(net3490),
    .A1(net4608),
    .S(_05171_),
    .X(_01945_));
 sg13g2_mux2_1 _14368_ (.A0(net3443),
    .A1(net4395),
    .S(_05171_),
    .X(_01946_));
 sg13g2_mux2_1 _14369_ (.A0(net3398),
    .A1(net4883),
    .S(_05171_),
    .X(_01947_));
 sg13g2_mux2_1 _14370_ (.A0(net3353),
    .A1(net4286),
    .S(_05171_),
    .X(_01948_));
 sg13g2_mux2_1 _14371_ (.A0(net3309),
    .A1(net4262),
    .S(_05171_),
    .X(_01949_));
 sg13g2_mux2_1 _14372_ (.A0(net3259),
    .A1(net4031),
    .S(_05171_),
    .X(_01950_));
 sg13g2_nor2_2 _14373_ (.A(_02338_),
    .B(_05008_),
    .Y(_05172_));
 sg13g2_mux2_1 _14374_ (.A0(net2260),
    .A1(net3576),
    .S(_05172_),
    .X(_01951_));
 sg13g2_mux2_1 _14375_ (.A0(net2364),
    .A1(net3529),
    .S(_05172_),
    .X(_01952_));
 sg13g2_mux2_1 _14376_ (.A0(net2629),
    .A1(net3489),
    .S(_05172_),
    .X(_01953_));
 sg13g2_mux2_1 _14377_ (.A0(net2370),
    .A1(net3436),
    .S(_05172_),
    .X(_01954_));
 sg13g2_mux2_1 _14378_ (.A0(net2722),
    .A1(net3397),
    .S(_05172_),
    .X(_01955_));
 sg13g2_mux2_1 _14379_ (.A0(net2569),
    .A1(net3345),
    .S(_05172_),
    .X(_01956_));
 sg13g2_mux2_1 _14380_ (.A0(net2796),
    .A1(net3299),
    .S(_05172_),
    .X(_01957_));
 sg13g2_mux2_1 _14381_ (.A0(net2236),
    .A1(net3258),
    .S(_05172_),
    .X(_01958_));
 sg13g2_nand2_2 _14382_ (.Y(_05173_),
    .A(net3070),
    .B(_05007_));
 sg13g2_mux2_1 _14383_ (.A0(net3576),
    .A1(net4143),
    .S(_05173_),
    .X(_01959_));
 sg13g2_mux2_1 _14384_ (.A0(net3529),
    .A1(net4237),
    .S(_05173_),
    .X(_01960_));
 sg13g2_mux2_1 _14385_ (.A0(net3489),
    .A1(net4380),
    .S(_05173_),
    .X(_01961_));
 sg13g2_mux2_1 _14386_ (.A0(net3436),
    .A1(net4653),
    .S(_05173_),
    .X(_01962_));
 sg13g2_mux2_1 _14387_ (.A0(net3397),
    .A1(net4743),
    .S(_05173_),
    .X(_01963_));
 sg13g2_mux2_1 _14388_ (.A0(net3345),
    .A1(net4981),
    .S(_05173_),
    .X(_01964_));
 sg13g2_mux2_1 _14389_ (.A0(net3299),
    .A1(net4522),
    .S(_05173_),
    .X(_01965_));
 sg13g2_mux2_1 _14390_ (.A0(net3258),
    .A1(net4337),
    .S(_05173_),
    .X(_01966_));
 sg13g2_nand2_2 _14391_ (.Y(_05174_),
    .A(_02332_),
    .B(net3051));
 sg13g2_mux2_1 _14392_ (.A0(net3576),
    .A1(net4574),
    .S(_05174_),
    .X(_01967_));
 sg13g2_mux2_1 _14393_ (.A0(net3526),
    .A1(net4368),
    .S(_05174_),
    .X(_01968_));
 sg13g2_mux2_1 _14394_ (.A0(net3489),
    .A1(net2966),
    .S(_05174_),
    .X(_01969_));
 sg13g2_mux2_1 _14395_ (.A0(net3443),
    .A1(net4521),
    .S(_05174_),
    .X(_01970_));
 sg13g2_mux2_1 _14396_ (.A0(net3397),
    .A1(net3002),
    .S(_05174_),
    .X(_01971_));
 sg13g2_mux2_1 _14397_ (.A0(net3345),
    .A1(net4451),
    .S(_05174_),
    .X(_01972_));
 sg13g2_mux2_1 _14398_ (.A0(net3298),
    .A1(net4507),
    .S(_05174_),
    .X(_01973_));
 sg13g2_mux2_1 _14399_ (.A0(net3252),
    .A1(net5146),
    .S(_05174_),
    .X(_01974_));
 sg13g2_nand2_2 _14400_ (.Y(_05175_),
    .A(_02328_),
    .B(net3051));
 sg13g2_mux2_1 _14401_ (.A0(net3576),
    .A1(net4058),
    .S(_05175_),
    .X(_01975_));
 sg13g2_mux2_1 _14402_ (.A0(net3526),
    .A1(net4974),
    .S(_05175_),
    .X(_01976_));
 sg13g2_mux2_1 _14403_ (.A0(net3489),
    .A1(net4341),
    .S(_05175_),
    .X(_01977_));
 sg13g2_mux2_1 _14404_ (.A0(net3443),
    .A1(net4183),
    .S(_05175_),
    .X(_01978_));
 sg13g2_mux2_1 _14405_ (.A0(net3397),
    .A1(net4112),
    .S(_05175_),
    .X(_01979_));
 sg13g2_mux2_1 _14406_ (.A0(net3345),
    .A1(net4534),
    .S(_05175_),
    .X(_01980_));
 sg13g2_mux2_1 _14407_ (.A0(net3301),
    .A1(net4849),
    .S(_05175_),
    .X(_01981_));
 sg13g2_mux2_1 _14408_ (.A0(net3258),
    .A1(net5155),
    .S(_05175_),
    .X(_01982_));
 sg13g2_nand2_2 _14409_ (.Y(_05176_),
    .A(net3072),
    .B(net3051));
 sg13g2_mux2_1 _14410_ (.A0(net3576),
    .A1(net2805),
    .S(_05176_),
    .X(_01983_));
 sg13g2_mux2_1 _14411_ (.A0(net3529),
    .A1(net4717),
    .S(_05176_),
    .X(_01984_));
 sg13g2_mux2_1 _14412_ (.A0(net3489),
    .A1(net4715),
    .S(_05176_),
    .X(_01985_));
 sg13g2_mux2_1 _14413_ (.A0(net3436),
    .A1(net4727),
    .S(_05176_),
    .X(_01986_));
 sg13g2_mux2_1 _14414_ (.A0(net3397),
    .A1(net2639),
    .S(_05176_),
    .X(_01987_));
 sg13g2_mux2_1 _14415_ (.A0(net3345),
    .A1(net2841),
    .S(_05176_),
    .X(_01988_));
 sg13g2_mux2_1 _14416_ (.A0(net3299),
    .A1(net4151),
    .S(_05176_),
    .X(_01989_));
 sg13g2_mux2_1 _14417_ (.A0(net3258),
    .A1(net5048),
    .S(_05176_),
    .X(_01990_));
 sg13g2_nand3_1 _14418_ (.B(net3073),
    .C(net3051),
    .A(net3043),
    .Y(_05177_));
 sg13g2_mux2_1 _14419_ (.A0(net3576),
    .A1(net4502),
    .S(_05177_),
    .X(_01991_));
 sg13g2_mux2_1 _14420_ (.A0(net3527),
    .A1(net4470),
    .S(_05177_),
    .X(_01992_));
 sg13g2_mux2_1 _14421_ (.A0(net3489),
    .A1(net4424),
    .S(_05177_),
    .X(_01993_));
 sg13g2_mux2_1 _14422_ (.A0(net3436),
    .A1(net2964),
    .S(_05177_),
    .X(_01994_));
 sg13g2_mux2_1 _14423_ (.A0(net3397),
    .A1(net5141),
    .S(_05177_),
    .X(_01995_));
 sg13g2_mux2_1 _14424_ (.A0(net3345),
    .A1(net4464),
    .S(_05177_),
    .X(_01996_));
 sg13g2_mux2_1 _14425_ (.A0(net3299),
    .A1(net5070),
    .S(_05177_),
    .X(_01997_));
 sg13g2_mux2_1 _14426_ (.A0(net3258),
    .A1(net4513),
    .S(_05177_),
    .X(_01998_));
 sg13g2_nand2_2 _14427_ (.Y(_05178_),
    .A(net3084),
    .B(_05007_));
 sg13g2_mux2_1 _14428_ (.A0(net3575),
    .A1(net5158),
    .S(_05178_),
    .X(_01999_));
 sg13g2_mux2_1 _14429_ (.A0(net3527),
    .A1(net2772),
    .S(_05178_),
    .X(_02000_));
 sg13g2_mux2_1 _14430_ (.A0(net3489),
    .A1(net4920),
    .S(_05178_),
    .X(_02001_));
 sg13g2_mux2_1 _14431_ (.A0(net3436),
    .A1(net2832),
    .S(_05178_),
    .X(_02002_));
 sg13g2_mux2_1 _14432_ (.A0(net3397),
    .A1(net2894),
    .S(_05178_),
    .X(_02003_));
 sg13g2_mux2_1 _14433_ (.A0(net3345),
    .A1(net2879),
    .S(_05178_),
    .X(_02004_));
 sg13g2_mux2_1 _14434_ (.A0(net3299),
    .A1(net4640),
    .S(_05178_),
    .X(_02005_));
 sg13g2_mux2_1 _14435_ (.A0(net3259),
    .A1(net4025),
    .S(_05178_),
    .X(_02006_));
 sg13g2_nand2_2 _14436_ (.Y(_05179_),
    .A(_02309_),
    .B(net3035));
 sg13g2_mux2_1 _14437_ (.A0(net3595),
    .A1(net4020),
    .S(_05179_),
    .X(_02007_));
 sg13g2_mux2_1 _14438_ (.A0(net3549),
    .A1(net4285),
    .S(_05179_),
    .X(_02008_));
 sg13g2_mux2_1 _14439_ (.A0(net3502),
    .A1(net4943),
    .S(_05179_),
    .X(_02009_));
 sg13g2_mux2_1 _14440_ (.A0(net3456),
    .A1(net4731),
    .S(_05179_),
    .X(_02010_));
 sg13g2_mux2_1 _14441_ (.A0(net3410),
    .A1(net4612),
    .S(_05179_),
    .X(_02011_));
 sg13g2_mux2_1 _14442_ (.A0(net3367),
    .A1(net4878),
    .S(_05179_),
    .X(_02012_));
 sg13g2_mux2_1 _14443_ (.A0(net3321),
    .A1(net5162),
    .S(_05179_),
    .X(_02013_));
 sg13g2_mux2_1 _14444_ (.A0(net3271),
    .A1(net4265),
    .S(_05179_),
    .X(_02014_));
 sg13g2_nand2_2 _14445_ (.Y(_05180_),
    .A(net3079),
    .B(_05001_));
 sg13g2_mux2_1 _14446_ (.A0(net3572),
    .A1(net4053),
    .S(_05180_),
    .X(_02015_));
 sg13g2_mux2_1 _14447_ (.A0(net3525),
    .A1(net4712),
    .S(_05180_),
    .X(_02016_));
 sg13g2_mux2_1 _14448_ (.A0(net3479),
    .A1(net4287),
    .S(_05180_),
    .X(_02017_));
 sg13g2_mux2_1 _14449_ (.A0(net3432),
    .A1(net5026),
    .S(_05180_),
    .X(_02018_));
 sg13g2_mux2_1 _14450_ (.A0(net3388),
    .A1(net4281),
    .S(_05180_),
    .X(_02019_));
 sg13g2_mux2_1 _14451_ (.A0(net3344),
    .A1(net4210),
    .S(_05180_),
    .X(_02020_));
 sg13g2_mux2_1 _14452_ (.A0(net3297),
    .A1(net4361),
    .S(_05180_),
    .X(_02021_));
 sg13g2_mux2_1 _14453_ (.A0(net3250),
    .A1(net4932),
    .S(_05180_),
    .X(_02022_));
 sg13g2_nor2_2 _14454_ (.A(_02298_),
    .B(_05002_),
    .Y(_05181_));
 sg13g2_mux2_1 _14455_ (.A0(net2755),
    .A1(net3572),
    .S(_05181_),
    .X(_02023_));
 sg13g2_mux2_1 _14456_ (.A0(net2599),
    .A1(net3525),
    .S(_05181_),
    .X(_02024_));
 sg13g2_mux2_1 _14457_ (.A0(net2223),
    .A1(net3479),
    .S(_05181_),
    .X(_02025_));
 sg13g2_mux2_1 _14458_ (.A0(net2273),
    .A1(net3432),
    .S(_05181_),
    .X(_02026_));
 sg13g2_mux2_1 _14459_ (.A0(net2668),
    .A1(net3388),
    .S(_05181_),
    .X(_02027_));
 sg13g2_mux2_1 _14460_ (.A0(net2391),
    .A1(net3344),
    .S(_05181_),
    .X(_02028_));
 sg13g2_mux2_1 _14461_ (.A0(net2233),
    .A1(net3298),
    .S(_05181_),
    .X(_02029_));
 sg13g2_mux2_1 _14462_ (.A0(net2574),
    .A1(net3251),
    .S(_05181_),
    .X(_02030_));
 sg13g2_nand2_2 _14463_ (.Y(_05182_),
    .A(_02288_),
    .B(_05001_));
 sg13g2_mux2_1 _14464_ (.A0(net3572),
    .A1(net5139),
    .S(_05182_),
    .X(_02031_));
 sg13g2_mux2_1 _14465_ (.A0(net3525),
    .A1(net4928),
    .S(_05182_),
    .X(_02032_));
 sg13g2_mux2_1 _14466_ (.A0(net3478),
    .A1(net4914),
    .S(_05182_),
    .X(_02033_));
 sg13g2_mux2_1 _14467_ (.A0(net3435),
    .A1(net2932),
    .S(_05182_),
    .X(_02034_));
 sg13g2_mux2_1 _14468_ (.A0(net3388),
    .A1(net4975),
    .S(_05182_),
    .X(_02035_));
 sg13g2_mux2_1 _14469_ (.A0(net3344),
    .A1(net4710),
    .S(_05182_),
    .X(_02036_));
 sg13g2_mux2_1 _14470_ (.A0(net3298),
    .A1(net4740),
    .S(_05182_),
    .X(_02037_));
 sg13g2_mux2_1 _14471_ (.A0(net3250),
    .A1(net4567),
    .S(_05182_),
    .X(_02038_));
 sg13g2_nand2_2 _14472_ (.Y(_05183_),
    .A(_02254_),
    .B(net3033));
 sg13g2_mux2_1 _14473_ (.A0(net3572),
    .A1(net4941),
    .S(_05183_),
    .X(_02039_));
 sg13g2_mux2_1 _14474_ (.A0(net3526),
    .A1(net4750),
    .S(_05183_),
    .X(_02040_));
 sg13g2_mux2_1 _14475_ (.A0(net3480),
    .A1(net4164),
    .S(_05183_),
    .X(_02041_));
 sg13g2_mux2_1 _14476_ (.A0(net3434),
    .A1(net4129),
    .S(_05183_),
    .X(_02042_));
 sg13g2_mux2_1 _14477_ (.A0(net3388),
    .A1(net5161),
    .S(_05183_),
    .X(_02043_));
 sg13g2_mux2_1 _14478_ (.A0(net3344),
    .A1(net4926),
    .S(_05183_),
    .X(_02044_));
 sg13g2_mux2_1 _14479_ (.A0(net3298),
    .A1(net4607),
    .S(_05183_),
    .X(_02045_));
 sg13g2_mux2_1 _14480_ (.A0(net3251),
    .A1(net4427),
    .S(_05183_),
    .X(_02046_));
 sg13g2_nor2_2 _14481_ (.A(net3081),
    .B(_05002_),
    .Y(_05184_));
 sg13g2_mux2_1 _14482_ (.A0(net2286),
    .A1(net3572),
    .S(_05184_),
    .X(_02047_));
 sg13g2_mux2_1 _14483_ (.A0(net2168),
    .A1(net3525),
    .S(_05184_),
    .X(_02048_));
 sg13g2_mux2_1 _14484_ (.A0(net2712),
    .A1(net3478),
    .S(_05184_),
    .X(_02049_));
 sg13g2_mux2_1 _14485_ (.A0(net2580),
    .A1(net3433),
    .S(_05184_),
    .X(_02050_));
 sg13g2_mux2_1 _14486_ (.A0(net2407),
    .A1(net3387),
    .S(_05184_),
    .X(_02051_));
 sg13g2_mux2_1 _14487_ (.A0(net2192),
    .A1(net3344),
    .S(_05184_),
    .X(_02052_));
 sg13g2_mux2_1 _14488_ (.A0(net2348),
    .A1(net3298),
    .S(_05184_),
    .X(_02053_));
 sg13g2_mux2_1 _14489_ (.A0(net2609),
    .A1(net3251),
    .S(_05184_),
    .X(_02054_));
 sg13g2_and2_2 _14490_ (.A(_02254_),
    .B(_02346_),
    .X(_05185_));
 sg13g2_mux2_1 _14491_ (.A0(net2563),
    .A1(net3572),
    .S(_05185_),
    .X(_02055_));
 sg13g2_mux2_1 _14492_ (.A0(net2232),
    .A1(net3525),
    .S(_05185_),
    .X(_02056_));
 sg13g2_mux2_1 _14493_ (.A0(net2225),
    .A1(net3478),
    .S(_05185_),
    .X(_02057_));
 sg13g2_mux2_1 _14494_ (.A0(net2300),
    .A1(net3433),
    .S(_05185_),
    .X(_02058_));
 sg13g2_mux2_1 _14495_ (.A0(net2497),
    .A1(net3387),
    .S(_05185_),
    .X(_02059_));
 sg13g2_mux2_1 _14496_ (.A0(net2238),
    .A1(net3344),
    .S(_05185_),
    .X(_02060_));
 sg13g2_mux2_1 _14497_ (.A0(net2476),
    .A1(net3298),
    .S(_05185_),
    .X(_02061_));
 sg13g2_mux2_1 _14498_ (.A0(net2392),
    .A1(net3251),
    .S(_05185_),
    .X(_02062_));
 sg13g2_and2_2 _14499_ (.A(_02254_),
    .B(_02385_),
    .X(_05186_));
 sg13g2_mux2_1 _14500_ (.A0(net2243),
    .A1(net3572),
    .S(_05186_),
    .X(_02063_));
 sg13g2_mux2_1 _14501_ (.A0(net2345),
    .A1(net3525),
    .S(_05186_),
    .X(_02064_));
 sg13g2_mux2_1 _14502_ (.A0(net2421),
    .A1(net3478),
    .S(_05186_),
    .X(_02065_));
 sg13g2_mux2_1 _14503_ (.A0(net2452),
    .A1(net3432),
    .S(_05186_),
    .X(_02066_));
 sg13g2_mux2_1 _14504_ (.A0(net2441),
    .A1(net3387),
    .S(_05186_),
    .X(_02067_));
 sg13g2_mux2_1 _14505_ (.A0(net2552),
    .A1(net3344),
    .S(_05186_),
    .X(_02068_));
 sg13g2_mux2_1 _14506_ (.A0(net2206),
    .A1(net3298),
    .S(_05186_),
    .X(_02069_));
 sg13g2_mux2_1 _14507_ (.A0(net2634),
    .A1(net3251),
    .S(_05186_),
    .X(_02070_));
 sg13g2_nand2_2 _14508_ (.Y(_05187_),
    .A(_02309_),
    .B(_05001_));
 sg13g2_mux2_1 _14509_ (.A0(net3572),
    .A1(net4888),
    .S(_05187_),
    .X(_02071_));
 sg13g2_mux2_1 _14510_ (.A0(net3526),
    .A1(net4310),
    .S(_05187_),
    .X(_02072_));
 sg13g2_mux2_1 _14511_ (.A0(net3480),
    .A1(net4268),
    .S(_05187_),
    .X(_02073_));
 sg13g2_mux2_1 _14512_ (.A0(net3432),
    .A1(net4326),
    .S(_05187_),
    .X(_02074_));
 sg13g2_mux2_1 _14513_ (.A0(net3387),
    .A1(net4576),
    .S(_05187_),
    .X(_02075_));
 sg13g2_mux2_1 _14514_ (.A0(net3344),
    .A1(net4378),
    .S(_05187_),
    .X(_02076_));
 sg13g2_mux2_1 _14515_ (.A0(net3298),
    .A1(net4213),
    .S(_05187_),
    .X(_02077_));
 sg13g2_mux2_1 _14516_ (.A0(net3251),
    .A1(net4026),
    .S(_05187_),
    .X(_02078_));
 sg13g2_nor2_2 _14517_ (.A(_02338_),
    .B(_05002_),
    .Y(_05188_));
 sg13g2_mux2_1 _14518_ (.A0(net2586),
    .A1(net3573),
    .S(_05188_),
    .X(_02079_));
 sg13g2_mux2_1 _14519_ (.A0(net2570),
    .A1(net3526),
    .S(_05188_),
    .X(_02080_));
 sg13g2_mux2_1 _14520_ (.A0(net2557),
    .A1(net3482),
    .S(_05188_),
    .X(_02081_));
 sg13g2_mux2_1 _14521_ (.A0(net2488),
    .A1(net3434),
    .S(_05188_),
    .X(_02082_));
 sg13g2_mux2_1 _14522_ (.A0(net2272),
    .A1(net3387),
    .S(_05188_),
    .X(_02083_));
 sg13g2_mux2_1 _14523_ (.A0(net2687),
    .A1(net3343),
    .S(_05188_),
    .X(_02084_));
 sg13g2_mux2_1 _14524_ (.A0(net2778),
    .A1(net3297),
    .S(_05188_),
    .X(_02085_));
 sg13g2_mux2_1 _14525_ (.A0(net2517),
    .A1(net3251),
    .S(_05188_),
    .X(_02086_));
 sg13g2_nand2_2 _14526_ (.Y(_05189_),
    .A(_02337_),
    .B(net3035));
 sg13g2_mux2_1 _14527_ (.A0(net3593),
    .A1(net4933),
    .S(_05189_),
    .X(_02087_));
 sg13g2_mux2_1 _14528_ (.A0(net3549),
    .A1(net4995),
    .S(_05189_),
    .X(_02088_));
 sg13g2_mux2_1 _14529_ (.A0(net3502),
    .A1(net4161),
    .S(_05189_),
    .X(_02089_));
 sg13g2_mux2_1 _14530_ (.A0(net3457),
    .A1(net4453),
    .S(_05189_),
    .X(_02090_));
 sg13g2_mux2_1 _14531_ (.A0(net3411),
    .A1(net4473),
    .S(_05189_),
    .X(_02091_));
 sg13g2_mux2_1 _14532_ (.A0(net3367),
    .A1(net4901),
    .S(_05189_),
    .X(_02092_));
 sg13g2_mux2_1 _14533_ (.A0(net3321),
    .A1(net4089),
    .S(_05189_),
    .X(_02093_));
 sg13g2_mux2_1 _14534_ (.A0(net3272),
    .A1(net5008),
    .S(_05189_),
    .X(_02094_));
 sg13g2_nor2_2 _14535_ (.A(_02331_),
    .B(_05002_),
    .Y(_05190_));
 sg13g2_mux2_1 _14536_ (.A0(net2331),
    .A1(net3573),
    .S(_05190_),
    .X(_02095_));
 sg13g2_mux2_1 _14537_ (.A0(net2482),
    .A1(net3526),
    .S(_05190_),
    .X(_02096_));
 sg13g2_mux2_1 _14538_ (.A0(net2464),
    .A1(net3481),
    .S(_05190_),
    .X(_02097_));
 sg13g2_mux2_1 _14539_ (.A0(net2562),
    .A1(net3434),
    .S(_05190_),
    .X(_02098_));
 sg13g2_mux2_1 _14540_ (.A0(net2565),
    .A1(net3387),
    .S(_05190_),
    .X(_02099_));
 sg13g2_mux2_1 _14541_ (.A0(net2215),
    .A1(net3343),
    .S(_05190_),
    .X(_02100_));
 sg13g2_mux2_1 _14542_ (.A0(net2467),
    .A1(net3297),
    .S(_05190_),
    .X(_02101_));
 sg13g2_mux2_1 _14543_ (.A0(net2402),
    .A1(net3252),
    .S(_05190_),
    .X(_02102_));
 sg13g2_and2_2 _14544_ (.A(_02254_),
    .B(_02328_),
    .X(_05191_));
 sg13g2_mux2_1 _14545_ (.A0(net2276),
    .A1(net3573),
    .S(_05191_),
    .X(_02103_));
 sg13g2_mux2_1 _14546_ (.A0(net2420),
    .A1(net3526),
    .S(_05191_),
    .X(_02104_));
 sg13g2_mux2_1 _14547_ (.A0(net2397),
    .A1(net3481),
    .S(_05191_),
    .X(_02105_));
 sg13g2_mux2_1 _14548_ (.A0(net2350),
    .A1(net3434),
    .S(_05191_),
    .X(_02106_));
 sg13g2_mux2_1 _14549_ (.A0(net2255),
    .A1(net3387),
    .S(_05191_),
    .X(_02107_));
 sg13g2_mux2_1 _14550_ (.A0(net2404),
    .A1(net3342),
    .S(_05191_),
    .X(_02108_));
 sg13g2_mux2_1 _14551_ (.A0(net2240),
    .A1(net3300),
    .S(_05191_),
    .X(_02109_));
 sg13g2_mux2_1 _14552_ (.A0(net2648),
    .A1(net3252),
    .S(_05191_),
    .X(_02110_));
 sg13g2_nand2_2 _14553_ (.Y(_05192_),
    .A(_02311_),
    .B(net3070));
 sg13g2_mux2_1 _14554_ (.A0(net3582),
    .A1(net5091),
    .S(_05192_),
    .X(_02111_));
 sg13g2_mux2_1 _14555_ (.A0(net3536),
    .A1(net4443),
    .S(_05192_),
    .X(_02112_));
 sg13g2_mux2_1 _14556_ (.A0(net3492),
    .A1(net4387),
    .S(_05192_),
    .X(_02113_));
 sg13g2_mux2_1 _14557_ (.A0(net3445),
    .A1(net4282),
    .S(_05192_),
    .X(_02114_));
 sg13g2_mux2_1 _14558_ (.A0(net3400),
    .A1(net4699),
    .S(_05192_),
    .X(_02115_));
 sg13g2_mux2_1 _14559_ (.A0(net3356),
    .A1(net4886),
    .S(_05192_),
    .X(_02116_));
 sg13g2_mux2_1 _14560_ (.A0(net3311),
    .A1(net4181),
    .S(_05192_),
    .X(_02117_));
 sg13g2_mux2_1 _14561_ (.A0(net3263),
    .A1(net4537),
    .S(_05192_),
    .X(_02118_));
 sg13g2_nor2_1 _14562_ (.A(net3997),
    .B(net3047),
    .Y(_02119_));
 sg13g2_nor3_1 _14563_ (.A(net3998),
    .B(_02421_),
    .C(_02422_),
    .Y(_00630_));
 sg13g2_a21oi_1 _14564_ (.A1(_02432_),
    .A2(_02433_),
    .Y(_00631_),
    .B1(net3996));
 sg13g2_a21oi_1 _14565_ (.A1(_02444_),
    .A2(_02445_),
    .Y(_00632_),
    .B1(net3995));
 sg13g2_a21oi_1 _14566_ (.A1(net3017),
    .A2(_02454_),
    .Y(_00633_),
    .B1(_02455_));
 sg13g2_a21oi_1 _14567_ (.A1(net3019),
    .A2(_02464_),
    .Y(_00634_),
    .B1(_02465_));
 sg13g2_a21oi_1 _14568_ (.A1(net3017),
    .A2(_02475_),
    .Y(_00635_),
    .B1(_02476_));
 sg13g2_nor2_1 _14569_ (.A(net3996),
    .B(_02488_),
    .Y(_00636_));
 sg13g2_nor2_1 _14570_ (.A(net3996),
    .B(_02497_),
    .Y(_00637_));
 sg13g2_dfrbp_1 _14571_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net343),
    .D(_00018_),
    .Q_N(_07284_),
    .Q(\mem.mem[94][0] ));
 sg13g2_dfrbp_1 _14572_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1238),
    .D(_00019_),
    .Q_N(_07283_),
    .Q(\mem.mem[94][1] ));
 sg13g2_dfrbp_1 _14573_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1237),
    .D(_00020_),
    .Q_N(_07282_),
    .Q(\mem.mem[94][2] ));
 sg13g2_dfrbp_1 _14574_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1236),
    .D(_00021_),
    .Q_N(_07281_),
    .Q(\mem.mem[94][3] ));
 sg13g2_dfrbp_1 _14575_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1235),
    .D(_00022_),
    .Q_N(_07280_),
    .Q(\mem.mem[94][4] ));
 sg13g2_dfrbp_1 _14576_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1234),
    .D(_00023_),
    .Q_N(_07279_),
    .Q(\mem.mem[94][5] ));
 sg13g2_dfrbp_1 _14577_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1233),
    .D(_00024_),
    .Q_N(_07278_),
    .Q(\mem.mem[94][6] ));
 sg13g2_dfrbp_1 _14578_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1232),
    .D(_00025_),
    .Q_N(_07277_),
    .Q(\mem.mem[94][7] ));
 sg13g2_dfrbp_1 _14579_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1231),
    .D(_00026_),
    .Q_N(_07276_),
    .Q(\mem.mem[4][0] ));
 sg13g2_dfrbp_1 _14580_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1230),
    .D(_00027_),
    .Q_N(_07275_),
    .Q(\mem.mem[4][1] ));
 sg13g2_dfrbp_1 _14581_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1229),
    .D(_00028_),
    .Q_N(_07274_),
    .Q(\mem.mem[4][2] ));
 sg13g2_dfrbp_1 _14582_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1228),
    .D(_00029_),
    .Q_N(_07273_),
    .Q(\mem.mem[4][3] ));
 sg13g2_dfrbp_1 _14583_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1227),
    .D(_00030_),
    .Q_N(_07272_),
    .Q(\mem.mem[4][4] ));
 sg13g2_dfrbp_1 _14584_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1226),
    .D(_00031_),
    .Q_N(_07271_),
    .Q(\mem.mem[4][5] ));
 sg13g2_dfrbp_1 _14585_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1225),
    .D(_00032_),
    .Q_N(_07270_),
    .Q(\mem.mem[4][6] ));
 sg13g2_dfrbp_1 _14586_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1224),
    .D(_00033_),
    .Q_N(_07269_),
    .Q(\mem.mem[4][7] ));
 sg13g2_dfrbp_1 _14587_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1223),
    .D(_00034_),
    .Q_N(_07268_),
    .Q(\mem.mem[48][0] ));
 sg13g2_dfrbp_1 _14588_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1222),
    .D(_00035_),
    .Q_N(_07267_),
    .Q(\mem.mem[48][1] ));
 sg13g2_dfrbp_1 _14589_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1221),
    .D(_00036_),
    .Q_N(_07266_),
    .Q(\mem.mem[48][2] ));
 sg13g2_dfrbp_1 _14590_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1220),
    .D(_00037_),
    .Q_N(_07265_),
    .Q(\mem.mem[48][3] ));
 sg13g2_dfrbp_1 _14591_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1219),
    .D(_00038_),
    .Q_N(_07264_),
    .Q(\mem.mem[48][4] ));
 sg13g2_dfrbp_1 _14592_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1218),
    .D(_00039_),
    .Q_N(_07263_),
    .Q(\mem.mem[48][5] ));
 sg13g2_dfrbp_1 _14593_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1217),
    .D(_00040_),
    .Q_N(_07262_),
    .Q(\mem.mem[48][6] ));
 sg13g2_dfrbp_1 _14594_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1216),
    .D(_00041_),
    .Q_N(_07261_),
    .Q(\mem.mem[48][7] ));
 sg13g2_dfrbp_1 _14595_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1215),
    .D(_00042_),
    .Q_N(_07260_),
    .Q(\mem.mem[80][0] ));
 sg13g2_dfrbp_1 _14596_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1214),
    .D(_00043_),
    .Q_N(_07259_),
    .Q(\mem.mem[80][1] ));
 sg13g2_dfrbp_1 _14597_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1213),
    .D(_00044_),
    .Q_N(_07258_),
    .Q(\mem.mem[80][2] ));
 sg13g2_dfrbp_1 _14598_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1212),
    .D(_00045_),
    .Q_N(_07257_),
    .Q(\mem.mem[80][3] ));
 sg13g2_dfrbp_1 _14599_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1211),
    .D(_00046_),
    .Q_N(_07256_),
    .Q(\mem.mem[80][4] ));
 sg13g2_dfrbp_1 _14600_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1210),
    .D(_00047_),
    .Q_N(_07255_),
    .Q(\mem.mem[80][5] ));
 sg13g2_dfrbp_1 _14601_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1209),
    .D(_00048_),
    .Q_N(_07254_),
    .Q(\mem.mem[80][6] ));
 sg13g2_dfrbp_1 _14602_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1208),
    .D(_00049_),
    .Q_N(_07253_),
    .Q(\mem.mem[80][7] ));
 sg13g2_dfrbp_1 _14603_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1207),
    .D(_00050_),
    .Q_N(_07252_),
    .Q(\mem.mem[34][0] ));
 sg13g2_dfrbp_1 _14604_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1206),
    .D(_00051_),
    .Q_N(_07251_),
    .Q(\mem.mem[34][1] ));
 sg13g2_dfrbp_1 _14605_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1205),
    .D(_00052_),
    .Q_N(_07250_),
    .Q(\mem.mem[34][2] ));
 sg13g2_dfrbp_1 _14606_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1204),
    .D(_00053_),
    .Q_N(_07249_),
    .Q(\mem.mem[34][3] ));
 sg13g2_dfrbp_1 _14607_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1203),
    .D(_00054_),
    .Q_N(_07248_),
    .Q(\mem.mem[34][4] ));
 sg13g2_dfrbp_1 _14608_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1202),
    .D(_00055_),
    .Q_N(_07247_),
    .Q(\mem.mem[34][5] ));
 sg13g2_dfrbp_1 _14609_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1201),
    .D(_00056_),
    .Q_N(_07246_),
    .Q(\mem.mem[34][6] ));
 sg13g2_dfrbp_1 _14610_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1200),
    .D(_00057_),
    .Q_N(_07245_),
    .Q(\mem.mem[34][7] ));
 sg13g2_dfrbp_1 _14611_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1199),
    .D(_00058_),
    .Q_N(_07244_),
    .Q(\mem.mem[209][0] ));
 sg13g2_dfrbp_1 _14612_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1198),
    .D(_00059_),
    .Q_N(_07243_),
    .Q(\mem.mem[209][1] ));
 sg13g2_dfrbp_1 _14613_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1197),
    .D(_00060_),
    .Q_N(_07242_),
    .Q(\mem.mem[209][2] ));
 sg13g2_dfrbp_1 _14614_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1196),
    .D(_00061_),
    .Q_N(_07241_),
    .Q(\mem.mem[209][3] ));
 sg13g2_dfrbp_1 _14615_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1195),
    .D(_00062_),
    .Q_N(_07240_),
    .Q(\mem.mem[209][4] ));
 sg13g2_dfrbp_1 _14616_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1194),
    .D(_00063_),
    .Q_N(_07239_),
    .Q(\mem.mem[209][5] ));
 sg13g2_dfrbp_1 _14617_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1193),
    .D(_00064_),
    .Q_N(_07238_),
    .Q(\mem.mem[209][6] ));
 sg13g2_dfrbp_1 _14618_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1192),
    .D(_00065_),
    .Q_N(_07237_),
    .Q(\mem.mem[209][7] ));
 sg13g2_dfrbp_1 _14619_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1191),
    .D(_00066_),
    .Q_N(_07236_),
    .Q(prev_run));
 sg13g2_dfrbp_1 _14620_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1190),
    .D(_00067_),
    .Q_N(_07235_),
    .Q(\mem.mem[47][0] ));
 sg13g2_dfrbp_1 _14621_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1189),
    .D(_00068_),
    .Q_N(_07234_),
    .Q(\mem.mem[47][1] ));
 sg13g2_dfrbp_1 _14622_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1188),
    .D(_00069_),
    .Q_N(_07233_),
    .Q(\mem.mem[47][2] ));
 sg13g2_dfrbp_1 _14623_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1187),
    .D(_00070_),
    .Q_N(_07232_),
    .Q(\mem.mem[47][3] ));
 sg13g2_dfrbp_1 _14624_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1186),
    .D(_00071_),
    .Q_N(_07231_),
    .Q(\mem.mem[47][4] ));
 sg13g2_dfrbp_1 _14625_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1185),
    .D(_00072_),
    .Q_N(_07230_),
    .Q(\mem.mem[47][5] ));
 sg13g2_dfrbp_1 _14626_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1184),
    .D(_00073_),
    .Q_N(_07229_),
    .Q(\mem.mem[47][6] ));
 sg13g2_dfrbp_1 _14627_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1183),
    .D(_00074_),
    .Q_N(_07228_),
    .Q(\mem.mem[47][7] ));
 sg13g2_dfrbp_1 _14628_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1182),
    .D(_00075_),
    .Q_N(_07227_),
    .Q(\mem.mem[7][0] ));
 sg13g2_dfrbp_1 _14629_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1181),
    .D(_00076_),
    .Q_N(_07226_),
    .Q(\mem.mem[7][1] ));
 sg13g2_dfrbp_1 _14630_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1180),
    .D(_00077_),
    .Q_N(_07225_),
    .Q(\mem.mem[7][2] ));
 sg13g2_dfrbp_1 _14631_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1179),
    .D(_00078_),
    .Q_N(_07224_),
    .Q(\mem.mem[7][3] ));
 sg13g2_dfrbp_1 _14632_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1178),
    .D(_00079_),
    .Q_N(_07223_),
    .Q(\mem.mem[7][4] ));
 sg13g2_dfrbp_1 _14633_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1177),
    .D(_00080_),
    .Q_N(_07222_),
    .Q(\mem.mem[7][5] ));
 sg13g2_dfrbp_1 _14634_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1176),
    .D(_00081_),
    .Q_N(_07221_),
    .Q(\mem.mem[7][6] ));
 sg13g2_dfrbp_1 _14635_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1175),
    .D(_00082_),
    .Q_N(_07220_),
    .Q(\mem.mem[7][7] ));
 sg13g2_dfrbp_1 _14636_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1174),
    .D(_00083_),
    .Q_N(_07219_),
    .Q(\mem.mem[78][0] ));
 sg13g2_dfrbp_1 _14637_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1173),
    .D(_00084_),
    .Q_N(_07218_),
    .Q(\mem.mem[78][1] ));
 sg13g2_dfrbp_1 _14638_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1172),
    .D(_00085_),
    .Q_N(_07217_),
    .Q(\mem.mem[78][2] ));
 sg13g2_dfrbp_1 _14639_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1171),
    .D(_00086_),
    .Q_N(_07216_),
    .Q(\mem.mem[78][3] ));
 sg13g2_dfrbp_1 _14640_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1170),
    .D(_00087_),
    .Q_N(_07215_),
    .Q(\mem.mem[78][4] ));
 sg13g2_dfrbp_1 _14641_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1169),
    .D(_00088_),
    .Q_N(_07214_),
    .Q(\mem.mem[78][5] ));
 sg13g2_dfrbp_1 _14642_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1168),
    .D(_00089_),
    .Q_N(_07213_),
    .Q(\mem.mem[78][6] ));
 sg13g2_dfrbp_1 _14643_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1167),
    .D(_00090_),
    .Q_N(_07212_),
    .Q(\mem.mem[78][7] ));
 sg13g2_dfrbp_1 _14644_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1166),
    .D(_00091_),
    .Q_N(_07211_),
    .Q(\mem.mem[93][0] ));
 sg13g2_dfrbp_1 _14645_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1165),
    .D(_00092_),
    .Q_N(_07210_),
    .Q(\mem.mem[93][1] ));
 sg13g2_dfrbp_1 _14646_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1164),
    .D(_00093_),
    .Q_N(_07209_),
    .Q(\mem.mem[93][2] ));
 sg13g2_dfrbp_1 _14647_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1163),
    .D(_00094_),
    .Q_N(_07208_),
    .Q(\mem.mem[93][3] ));
 sg13g2_dfrbp_1 _14648_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1162),
    .D(_00095_),
    .Q_N(_07207_),
    .Q(\mem.mem[93][4] ));
 sg13g2_dfrbp_1 _14649_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1161),
    .D(_00096_),
    .Q_N(_07206_),
    .Q(\mem.mem[93][5] ));
 sg13g2_dfrbp_1 _14650_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1160),
    .D(_00097_),
    .Q_N(_07205_),
    .Q(\mem.mem[93][6] ));
 sg13g2_dfrbp_1 _14651_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1159),
    .D(_00098_),
    .Q_N(_07204_),
    .Q(\mem.mem[93][7] ));
 sg13g2_dfrbp_1 _14652_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1158),
    .D(_00099_),
    .Q_N(_07203_),
    .Q(\mem.mem[77][0] ));
 sg13g2_dfrbp_1 _14653_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1157),
    .D(_00100_),
    .Q_N(_07202_),
    .Q(\mem.mem[77][1] ));
 sg13g2_dfrbp_1 _14654_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1156),
    .D(_00101_),
    .Q_N(_07201_),
    .Q(\mem.mem[77][2] ));
 sg13g2_dfrbp_1 _14655_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1155),
    .D(_00102_),
    .Q_N(_07200_),
    .Q(\mem.mem[77][3] ));
 sg13g2_dfrbp_1 _14656_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1154),
    .D(_00103_),
    .Q_N(_07199_),
    .Q(\mem.mem[77][4] ));
 sg13g2_dfrbp_1 _14657_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1153),
    .D(_00104_),
    .Q_N(_07198_),
    .Q(\mem.mem[77][5] ));
 sg13g2_dfrbp_1 _14658_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1152),
    .D(_00105_),
    .Q_N(_07197_),
    .Q(\mem.mem[77][6] ));
 sg13g2_dfrbp_1 _14659_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1151),
    .D(_00106_),
    .Q_N(_07196_),
    .Q(\mem.mem[77][7] ));
 sg13g2_dfrbp_1 _14660_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1150),
    .D(_00107_),
    .Q_N(_07195_),
    .Q(\mem.mem[92][0] ));
 sg13g2_dfrbp_1 _14661_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1149),
    .D(_00108_),
    .Q_N(_07194_),
    .Q(\mem.mem[92][1] ));
 sg13g2_dfrbp_1 _14662_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1148),
    .D(_00109_),
    .Q_N(_07193_),
    .Q(\mem.mem[92][2] ));
 sg13g2_dfrbp_1 _14663_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1147),
    .D(_00110_),
    .Q_N(_07192_),
    .Q(\mem.mem[92][3] ));
 sg13g2_dfrbp_1 _14664_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1146),
    .D(_00111_),
    .Q_N(_07191_),
    .Q(\mem.mem[92][4] ));
 sg13g2_dfrbp_1 _14665_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1145),
    .D(_00112_),
    .Q_N(_07190_),
    .Q(\mem.mem[92][5] ));
 sg13g2_dfrbp_1 _14666_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1144),
    .D(_00113_),
    .Q_N(_07189_),
    .Q(\mem.mem[92][6] ));
 sg13g2_dfrbp_1 _14667_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1143),
    .D(_00114_),
    .Q_N(_07188_),
    .Q(\mem.mem[92][7] ));
 sg13g2_dfrbp_1 _14668_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1142),
    .D(_00115_),
    .Q_N(_07187_),
    .Q(\mem.mem[76][0] ));
 sg13g2_dfrbp_1 _14669_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1141),
    .D(_00116_),
    .Q_N(_07186_),
    .Q(\mem.mem[76][1] ));
 sg13g2_dfrbp_1 _14670_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1140),
    .D(_00117_),
    .Q_N(_07185_),
    .Q(\mem.mem[76][2] ));
 sg13g2_dfrbp_1 _14671_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1139),
    .D(_00118_),
    .Q_N(_07184_),
    .Q(\mem.mem[76][3] ));
 sg13g2_dfrbp_1 _14672_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1138),
    .D(_00119_),
    .Q_N(_07183_),
    .Q(\mem.mem[76][4] ));
 sg13g2_dfrbp_1 _14673_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1137),
    .D(_00120_),
    .Q_N(_07182_),
    .Q(\mem.mem[76][5] ));
 sg13g2_dfrbp_1 _14674_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1136),
    .D(_00121_),
    .Q_N(_07181_),
    .Q(\mem.mem[76][6] ));
 sg13g2_dfrbp_1 _14675_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1135),
    .D(_00122_),
    .Q_N(_07180_),
    .Q(\mem.mem[76][7] ));
 sg13g2_dfrbp_1 _14676_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1134),
    .D(_00123_),
    .Q_N(_07179_),
    .Q(\mem.mem[75][0] ));
 sg13g2_dfrbp_1 _14677_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1133),
    .D(_00124_),
    .Q_N(_07178_),
    .Q(\mem.mem[75][1] ));
 sg13g2_dfrbp_1 _14678_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1132),
    .D(_00125_),
    .Q_N(_07177_),
    .Q(\mem.mem[75][2] ));
 sg13g2_dfrbp_1 _14679_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1131),
    .D(_00126_),
    .Q_N(_07176_),
    .Q(\mem.mem[75][3] ));
 sg13g2_dfrbp_1 _14680_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1130),
    .D(_00127_),
    .Q_N(_07175_),
    .Q(\mem.mem[75][4] ));
 sg13g2_dfrbp_1 _14681_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1129),
    .D(_00128_),
    .Q_N(_07174_),
    .Q(\mem.mem[75][5] ));
 sg13g2_dfrbp_1 _14682_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1128),
    .D(_00129_),
    .Q_N(_07173_),
    .Q(\mem.mem[75][6] ));
 sg13g2_dfrbp_1 _14683_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1127),
    .D(_00130_),
    .Q_N(_07172_),
    .Q(\mem.mem[75][7] ));
 sg13g2_dfrbp_1 _14684_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1126),
    .D(_00131_),
    .Q_N(_07171_),
    .Q(\mem.mem[74][0] ));
 sg13g2_dfrbp_1 _14685_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1125),
    .D(_00132_),
    .Q_N(_07170_),
    .Q(\mem.mem[74][1] ));
 sg13g2_dfrbp_1 _14686_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1124),
    .D(_00133_),
    .Q_N(_07169_),
    .Q(\mem.mem[74][2] ));
 sg13g2_dfrbp_1 _14687_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1123),
    .D(_00134_),
    .Q_N(_07168_),
    .Q(\mem.mem[74][3] ));
 sg13g2_dfrbp_1 _14688_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1122),
    .D(_00135_),
    .Q_N(_07167_),
    .Q(\mem.mem[74][4] ));
 sg13g2_dfrbp_1 _14689_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1121),
    .D(_00136_),
    .Q_N(_07166_),
    .Q(\mem.mem[74][5] ));
 sg13g2_dfrbp_1 _14690_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1120),
    .D(_00137_),
    .Q_N(_07165_),
    .Q(\mem.mem[74][6] ));
 sg13g2_dfrbp_1 _14691_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1119),
    .D(_00138_),
    .Q_N(_07164_),
    .Q(\mem.mem[74][7] ));
 sg13g2_dfrbp_1 _14692_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1118),
    .D(_00139_),
    .Q_N(_07163_),
    .Q(\mem.mem[73][0] ));
 sg13g2_dfrbp_1 _14693_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1117),
    .D(_00140_),
    .Q_N(_07162_),
    .Q(\mem.mem[73][1] ));
 sg13g2_dfrbp_1 _14694_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1116),
    .D(_00141_),
    .Q_N(_07161_),
    .Q(\mem.mem[73][2] ));
 sg13g2_dfrbp_1 _14695_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1115),
    .D(_00142_),
    .Q_N(_07160_),
    .Q(\mem.mem[73][3] ));
 sg13g2_dfrbp_1 _14696_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1114),
    .D(_00143_),
    .Q_N(_07159_),
    .Q(\mem.mem[73][4] ));
 sg13g2_dfrbp_1 _14697_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1113),
    .D(_00144_),
    .Q_N(_07158_),
    .Q(\mem.mem[73][5] ));
 sg13g2_dfrbp_1 _14698_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1112),
    .D(_00145_),
    .Q_N(_07157_),
    .Q(\mem.mem[73][6] ));
 sg13g2_dfrbp_1 _14699_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1111),
    .D(_00146_),
    .Q_N(_07156_),
    .Q(\mem.mem[73][7] ));
 sg13g2_dfrbp_1 _14700_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1110),
    .D(_00147_),
    .Q_N(_07155_),
    .Q(\mem.mem[72][0] ));
 sg13g2_dfrbp_1 _14701_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1109),
    .D(_00148_),
    .Q_N(_07154_),
    .Q(\mem.mem[72][1] ));
 sg13g2_dfrbp_1 _14702_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1108),
    .D(_00149_),
    .Q_N(_07153_),
    .Q(\mem.mem[72][2] ));
 sg13g2_dfrbp_1 _14703_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1107),
    .D(_00150_),
    .Q_N(_07152_),
    .Q(\mem.mem[72][3] ));
 sg13g2_dfrbp_1 _14704_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1106),
    .D(_00151_),
    .Q_N(_07151_),
    .Q(\mem.mem[72][4] ));
 sg13g2_dfrbp_1 _14705_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1105),
    .D(_00152_),
    .Q_N(_07150_),
    .Q(\mem.mem[72][5] ));
 sg13g2_dfrbp_1 _14706_ (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1104),
    .D(_00153_),
    .Q_N(_07149_),
    .Q(\mem.mem[72][6] ));
 sg13g2_dfrbp_1 _14707_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1103),
    .D(_00154_),
    .Q_N(_07148_),
    .Q(\mem.mem[72][7] ));
 sg13g2_dfrbp_1 _14708_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1102),
    .D(_00155_),
    .Q_N(_07147_),
    .Q(\mem.mem[46][0] ));
 sg13g2_dfrbp_1 _14709_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1101),
    .D(_00156_),
    .Q_N(_07146_),
    .Q(\mem.mem[46][1] ));
 sg13g2_dfrbp_1 _14710_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1100),
    .D(_00157_),
    .Q_N(_07145_),
    .Q(\mem.mem[46][2] ));
 sg13g2_dfrbp_1 _14711_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1099),
    .D(_00158_),
    .Q_N(_07144_),
    .Q(\mem.mem[46][3] ));
 sg13g2_dfrbp_1 _14712_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1098),
    .D(_00159_),
    .Q_N(_07143_),
    .Q(\mem.mem[46][4] ));
 sg13g2_dfrbp_1 _14713_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1097),
    .D(_00160_),
    .Q_N(_07142_),
    .Q(\mem.mem[46][5] ));
 sg13g2_dfrbp_1 _14714_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1096),
    .D(_00161_),
    .Q_N(_07141_),
    .Q(\mem.mem[46][6] ));
 sg13g2_dfrbp_1 _14715_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1095),
    .D(_00162_),
    .Q_N(_07140_),
    .Q(\mem.mem[46][7] ));
 sg13g2_dfrbp_1 _14716_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1094),
    .D(_00163_),
    .Q_N(_07139_),
    .Q(\mem.mem[69][0] ));
 sg13g2_dfrbp_1 _14717_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1093),
    .D(_00164_),
    .Q_N(_07138_),
    .Q(\mem.mem[69][1] ));
 sg13g2_dfrbp_1 _14718_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1092),
    .D(_00165_),
    .Q_N(_07137_),
    .Q(\mem.mem[69][2] ));
 sg13g2_dfrbp_1 _14719_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1091),
    .D(_00166_),
    .Q_N(_07136_),
    .Q(\mem.mem[69][3] ));
 sg13g2_dfrbp_1 _14720_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1090),
    .D(_00167_),
    .Q_N(_07135_),
    .Q(\mem.mem[69][4] ));
 sg13g2_dfrbp_1 _14721_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1089),
    .D(_00168_),
    .Q_N(_07134_),
    .Q(\mem.mem[69][5] ));
 sg13g2_dfrbp_1 _14722_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1088),
    .D(_00169_),
    .Q_N(_07133_),
    .Q(\mem.mem[69][6] ));
 sg13g2_dfrbp_1 _14723_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1087),
    .D(_00170_),
    .Q_N(_07132_),
    .Q(\mem.mem[69][7] ));
 sg13g2_dfrbp_1 _14724_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1086),
    .D(_00171_),
    .Q_N(_07131_),
    .Q(\mem.mem[45][0] ));
 sg13g2_dfrbp_1 _14725_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1085),
    .D(_00172_),
    .Q_N(_07130_),
    .Q(\mem.mem[45][1] ));
 sg13g2_dfrbp_1 _14726_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1084),
    .D(_00173_),
    .Q_N(_07129_),
    .Q(\mem.mem[45][2] ));
 sg13g2_dfrbp_1 _14727_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1083),
    .D(_00174_),
    .Q_N(_07128_),
    .Q(\mem.mem[45][3] ));
 sg13g2_dfrbp_1 _14728_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1082),
    .D(_00175_),
    .Q_N(_07127_),
    .Q(\mem.mem[45][4] ));
 sg13g2_dfrbp_1 _14729_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1081),
    .D(_00176_),
    .Q_N(_07126_),
    .Q(\mem.mem[45][5] ));
 sg13g2_dfrbp_1 _14730_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1080),
    .D(_00177_),
    .Q_N(_07125_),
    .Q(\mem.mem[45][6] ));
 sg13g2_dfrbp_1 _14731_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1079),
    .D(_00178_),
    .Q_N(_07124_),
    .Q(\mem.mem[45][7] ));
 sg13g2_dfrbp_1 _14732_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1078),
    .D(_00179_),
    .Q_N(_07123_),
    .Q(\mem.mem[19][0] ));
 sg13g2_dfrbp_1 _14733_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1077),
    .D(_00180_),
    .Q_N(_07122_),
    .Q(\mem.mem[19][1] ));
 sg13g2_dfrbp_1 _14734_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1076),
    .D(_00181_),
    .Q_N(_07121_),
    .Q(\mem.mem[19][2] ));
 sg13g2_dfrbp_1 _14735_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1075),
    .D(_00182_),
    .Q_N(_07120_),
    .Q(\mem.mem[19][3] ));
 sg13g2_dfrbp_1 _14736_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1074),
    .D(_00183_),
    .Q_N(_07119_),
    .Q(\mem.mem[19][4] ));
 sg13g2_dfrbp_1 _14737_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1073),
    .D(_00184_),
    .Q_N(_07118_),
    .Q(\mem.mem[19][5] ));
 sg13g2_dfrbp_1 _14738_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1072),
    .D(_00185_),
    .Q_N(_07117_),
    .Q(\mem.mem[19][6] ));
 sg13g2_dfrbp_1 _14739_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1071),
    .D(_00186_),
    .Q_N(_07116_),
    .Q(\mem.mem[19][7] ));
 sg13g2_dfrbp_1 _14740_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1070),
    .D(_00187_),
    .Q_N(_07115_),
    .Q(\mem.mem[179][0] ));
 sg13g2_dfrbp_1 _14741_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1069),
    .D(_00188_),
    .Q_N(_07114_),
    .Q(\mem.mem[179][1] ));
 sg13g2_dfrbp_1 _14742_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1068),
    .D(_00189_),
    .Q_N(_07113_),
    .Q(\mem.mem[179][2] ));
 sg13g2_dfrbp_1 _14743_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1067),
    .D(_00190_),
    .Q_N(_07112_),
    .Q(\mem.mem[179][3] ));
 sg13g2_dfrbp_1 _14744_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1066),
    .D(_00191_),
    .Q_N(_07111_),
    .Q(\mem.mem[179][4] ));
 sg13g2_dfrbp_1 _14745_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1065),
    .D(_00192_),
    .Q_N(_07110_),
    .Q(\mem.mem[179][5] ));
 sg13g2_dfrbp_1 _14746_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1064),
    .D(_00193_),
    .Q_N(_07109_),
    .Q(\mem.mem[179][6] ));
 sg13g2_dfrbp_1 _14747_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1063),
    .D(_00194_),
    .Q_N(_07108_),
    .Q(\mem.mem[179][7] ));
 sg13g2_dfrbp_1 _14748_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1062),
    .D(_00195_),
    .Q_N(_07107_),
    .Q(\mem.mem[44][0] ));
 sg13g2_dfrbp_1 _14749_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1061),
    .D(_00196_),
    .Q_N(_07106_),
    .Q(\mem.mem[44][1] ));
 sg13g2_dfrbp_1 _14750_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1060),
    .D(_00197_),
    .Q_N(_07105_),
    .Q(\mem.mem[44][2] ));
 sg13g2_dfrbp_1 _14751_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1059),
    .D(_00198_),
    .Q_N(_07104_),
    .Q(\mem.mem[44][3] ));
 sg13g2_dfrbp_1 _14752_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1058),
    .D(_00199_),
    .Q_N(_07103_),
    .Q(\mem.mem[44][4] ));
 sg13g2_dfrbp_1 _14753_ (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1057),
    .D(_00200_),
    .Q_N(_07102_),
    .Q(\mem.mem[44][5] ));
 sg13g2_dfrbp_1 _14754_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1056),
    .D(_00201_),
    .Q_N(_07101_),
    .Q(\mem.mem[44][6] ));
 sg13g2_dfrbp_1 _14755_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1055),
    .D(_00202_),
    .Q_N(_07100_),
    .Q(\mem.mem[44][7] ));
 sg13g2_dfrbp_1 _14756_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1054),
    .D(_00203_),
    .Q_N(_07099_),
    .Q(\mem.mem[119][0] ));
 sg13g2_dfrbp_1 _14757_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1053),
    .D(_00204_),
    .Q_N(_07098_),
    .Q(\mem.mem[119][1] ));
 sg13g2_dfrbp_1 _14758_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1052),
    .D(_00205_),
    .Q_N(_07097_),
    .Q(\mem.mem[119][2] ));
 sg13g2_dfrbp_1 _14759_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1051),
    .D(_00206_),
    .Q_N(_07096_),
    .Q(\mem.mem[119][3] ));
 sg13g2_dfrbp_1 _14760_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1050),
    .D(_00207_),
    .Q_N(_07095_),
    .Q(\mem.mem[119][4] ));
 sg13g2_dfrbp_1 _14761_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1049),
    .D(_00208_),
    .Q_N(_07094_),
    .Q(\mem.mem[119][5] ));
 sg13g2_dfrbp_1 _14762_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1048),
    .D(_00209_),
    .Q_N(_07093_),
    .Q(\mem.mem[119][6] ));
 sg13g2_dfrbp_1 _14763_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1047),
    .D(_00210_),
    .Q_N(_07092_),
    .Q(\mem.mem[119][7] ));
 sg13g2_dfrbp_1 _14764_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1046),
    .D(_00211_),
    .Q_N(_07091_),
    .Q(\mem.mem[43][0] ));
 sg13g2_dfrbp_1 _14765_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1045),
    .D(_00212_),
    .Q_N(_07090_),
    .Q(\mem.mem[43][1] ));
 sg13g2_dfrbp_1 _14766_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1044),
    .D(_00213_),
    .Q_N(_07089_),
    .Q(\mem.mem[43][2] ));
 sg13g2_dfrbp_1 _14767_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1043),
    .D(_00214_),
    .Q_N(_07088_),
    .Q(\mem.mem[43][3] ));
 sg13g2_dfrbp_1 _14768_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1042),
    .D(_00215_),
    .Q_N(_07087_),
    .Q(\mem.mem[43][4] ));
 sg13g2_dfrbp_1 _14769_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1041),
    .D(_00216_),
    .Q_N(_07086_),
    .Q(\mem.mem[43][5] ));
 sg13g2_dfrbp_1 _14770_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1040),
    .D(_00217_),
    .Q_N(_07085_),
    .Q(\mem.mem[43][6] ));
 sg13g2_dfrbp_1 _14771_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1039),
    .D(_00218_),
    .Q_N(_07084_),
    .Q(\mem.mem[43][7] ));
 sg13g2_dfrbp_1 _14772_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1038),
    .D(_00219_),
    .Q_N(_07083_),
    .Q(\mem.mem[169][0] ));
 sg13g2_dfrbp_1 _14773_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1037),
    .D(_00220_),
    .Q_N(_07082_),
    .Q(\mem.mem[169][1] ));
 sg13g2_dfrbp_1 _14774_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1036),
    .D(_00221_),
    .Q_N(_07081_),
    .Q(\mem.mem[169][2] ));
 sg13g2_dfrbp_1 _14775_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1035),
    .D(_00222_),
    .Q_N(_07080_),
    .Q(\mem.mem[169][3] ));
 sg13g2_dfrbp_1 _14776_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1034),
    .D(_00223_),
    .Q_N(_07079_),
    .Q(\mem.mem[169][4] ));
 sg13g2_dfrbp_1 _14777_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1033),
    .D(_00224_),
    .Q_N(_07078_),
    .Q(\mem.mem[169][5] ));
 sg13g2_dfrbp_1 _14778_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1032),
    .D(_00225_),
    .Q_N(_07077_),
    .Q(\mem.mem[169][6] ));
 sg13g2_dfrbp_1 _14779_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1031),
    .D(_00226_),
    .Q_N(_07076_),
    .Q(\mem.mem[169][7] ));
 sg13g2_dfrbp_1 _14780_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1030),
    .D(_00227_),
    .Q_N(_07075_),
    .Q(\mem.mem[159][0] ));
 sg13g2_dfrbp_1 _14781_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1029),
    .D(_00228_),
    .Q_N(_07074_),
    .Q(\mem.mem[159][1] ));
 sg13g2_dfrbp_1 _14782_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1028),
    .D(_00229_),
    .Q_N(_07073_),
    .Q(\mem.mem[159][2] ));
 sg13g2_dfrbp_1 _14783_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1027),
    .D(_00230_),
    .Q_N(_07072_),
    .Q(\mem.mem[159][3] ));
 sg13g2_dfrbp_1 _14784_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1026),
    .D(_00231_),
    .Q_N(_07071_),
    .Q(\mem.mem[159][4] ));
 sg13g2_dfrbp_1 _14785_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1025),
    .D(_00232_),
    .Q_N(_07070_),
    .Q(\mem.mem[159][5] ));
 sg13g2_dfrbp_1 _14786_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1024),
    .D(_00233_),
    .Q_N(_07069_),
    .Q(\mem.mem[159][6] ));
 sg13g2_dfrbp_1 _14787_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1023),
    .D(_00234_),
    .Q_N(_07068_),
    .Q(\mem.mem[159][7] ));
 sg13g2_dfrbp_1 _14788_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1022),
    .D(_00235_),
    .Q_N(_07067_),
    .Q(\mem.mem[79][0] ));
 sg13g2_dfrbp_1 _14789_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1021),
    .D(_00236_),
    .Q_N(_07066_),
    .Q(\mem.mem[79][1] ));
 sg13g2_dfrbp_1 _14790_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1020),
    .D(_00237_),
    .Q_N(_07065_),
    .Q(\mem.mem[79][2] ));
 sg13g2_dfrbp_1 _14791_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1019),
    .D(_00238_),
    .Q_N(_07064_),
    .Q(\mem.mem[79][3] ));
 sg13g2_dfrbp_1 _14792_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1018),
    .D(_00239_),
    .Q_N(_07063_),
    .Q(\mem.mem[79][4] ));
 sg13g2_dfrbp_1 _14793_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1017),
    .D(_00240_),
    .Q_N(_07062_),
    .Q(\mem.mem[79][5] ));
 sg13g2_dfrbp_1 _14794_ (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1016),
    .D(_00241_),
    .Q_N(_07061_),
    .Q(\mem.mem[79][6] ));
 sg13g2_dfrbp_1 _14795_ (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1015),
    .D(_00242_),
    .Q_N(_07060_),
    .Q(\mem.mem[79][7] ));
 sg13g2_dfrbp_1 _14796_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1014),
    .D(_00243_),
    .Q_N(_07059_),
    .Q(\mem.mem[129][0] ));
 sg13g2_dfrbp_1 _14797_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1013),
    .D(_00244_),
    .Q_N(_07058_),
    .Q(\mem.mem[129][1] ));
 sg13g2_dfrbp_1 _14798_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1012),
    .D(_00245_),
    .Q_N(_07057_),
    .Q(\mem.mem[129][2] ));
 sg13g2_dfrbp_1 _14799_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1011),
    .D(_00246_),
    .Q_N(_07056_),
    .Q(\mem.mem[129][3] ));
 sg13g2_dfrbp_1 _14800_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1010),
    .D(_00247_),
    .Q_N(_07055_),
    .Q(\mem.mem[129][4] ));
 sg13g2_dfrbp_1 _14801_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1009),
    .D(_00248_),
    .Q_N(_07054_),
    .Q(\mem.mem[129][5] ));
 sg13g2_dfrbp_1 _14802_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1008),
    .D(_00249_),
    .Q_N(_07053_),
    .Q(\mem.mem[129][6] ));
 sg13g2_dfrbp_1 _14803_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1007),
    .D(_00250_),
    .Q_N(_07052_),
    .Q(\mem.mem[129][7] ));
 sg13g2_dfrbp_1 _14804_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1006),
    .D(_00251_),
    .Q_N(_07051_),
    .Q(\mem.mem[149][0] ));
 sg13g2_dfrbp_1 _14805_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1005),
    .D(_00252_),
    .Q_N(_07050_),
    .Q(\mem.mem[149][1] ));
 sg13g2_dfrbp_1 _14806_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1004),
    .D(_00253_),
    .Q_N(_07049_),
    .Q(\mem.mem[149][2] ));
 sg13g2_dfrbp_1 _14807_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1003),
    .D(_00254_),
    .Q_N(_07048_),
    .Q(\mem.mem[149][3] ));
 sg13g2_dfrbp_1 _14808_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1002),
    .D(_00255_),
    .Q_N(_07047_),
    .Q(\mem.mem[149][4] ));
 sg13g2_dfrbp_1 _14809_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1001),
    .D(_00256_),
    .Q_N(_07046_),
    .Q(\mem.mem[149][5] ));
 sg13g2_dfrbp_1 _14810_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1000),
    .D(_00257_),
    .Q_N(_07045_),
    .Q(\mem.mem[149][6] ));
 sg13g2_dfrbp_1 _14811_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net999),
    .D(_00258_),
    .Q_N(_07044_),
    .Q(\mem.mem[149][7] ));
 sg13g2_dfrbp_1 _14812_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net998),
    .D(_00259_),
    .Q_N(_07043_),
    .Q(\mem.mem[42][0] ));
 sg13g2_dfrbp_1 _14813_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net997),
    .D(_00260_),
    .Q_N(_07042_),
    .Q(\mem.mem[42][1] ));
 sg13g2_dfrbp_1 _14814_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net996),
    .D(_00261_),
    .Q_N(_07041_),
    .Q(\mem.mem[42][2] ));
 sg13g2_dfrbp_1 _14815_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net995),
    .D(_00262_),
    .Q_N(_07040_),
    .Q(\mem.mem[42][3] ));
 sg13g2_dfrbp_1 _14816_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net994),
    .D(_00263_),
    .Q_N(_07039_),
    .Q(\mem.mem[42][4] ));
 sg13g2_dfrbp_1 _14817_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net993),
    .D(_00264_),
    .Q_N(_07038_),
    .Q(\mem.mem[42][5] ));
 sg13g2_dfrbp_1 _14818_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net992),
    .D(_00265_),
    .Q_N(_07037_),
    .Q(\mem.mem[42][6] ));
 sg13g2_dfrbp_1 _14819_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net991),
    .D(_00266_),
    .Q_N(_07036_),
    .Q(\mem.mem[42][7] ));
 sg13g2_dfrbp_1 _14820_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net990),
    .D(_00267_),
    .Q_N(_07035_),
    .Q(\mem.mem[59][0] ));
 sg13g2_dfrbp_1 _14821_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net989),
    .D(_00268_),
    .Q_N(_07034_),
    .Q(\mem.mem[59][1] ));
 sg13g2_dfrbp_1 _14822_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net988),
    .D(_00269_),
    .Q_N(_07033_),
    .Q(\mem.mem[59][2] ));
 sg13g2_dfrbp_1 _14823_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net987),
    .D(_00270_),
    .Q_N(_07032_),
    .Q(\mem.mem[59][3] ));
 sg13g2_dfrbp_1 _14824_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net986),
    .D(_00271_),
    .Q_N(_07031_),
    .Q(\mem.mem[59][4] ));
 sg13g2_dfrbp_1 _14825_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net985),
    .D(_00272_),
    .Q_N(_07030_),
    .Q(\mem.mem[59][5] ));
 sg13g2_dfrbp_1 _14826_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net984),
    .D(_00273_),
    .Q_N(_07029_),
    .Q(\mem.mem[59][6] ));
 sg13g2_dfrbp_1 _14827_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net983),
    .D(_00274_),
    .Q_N(_07028_),
    .Q(\mem.mem[59][7] ));
 sg13g2_dfrbp_1 _14828_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net982),
    .D(_00275_),
    .Q_N(_07027_),
    .Q(\mem.mem[41][0] ));
 sg13g2_dfrbp_1 _14829_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net981),
    .D(_00276_),
    .Q_N(_07026_),
    .Q(\mem.mem[41][1] ));
 sg13g2_dfrbp_1 _14830_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net980),
    .D(_00277_),
    .Q_N(_07025_),
    .Q(\mem.mem[41][2] ));
 sg13g2_dfrbp_1 _14831_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net979),
    .D(_00278_),
    .Q_N(_07024_),
    .Q(\mem.mem[41][3] ));
 sg13g2_dfrbp_1 _14832_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net978),
    .D(_00279_),
    .Q_N(_07023_),
    .Q(\mem.mem[41][4] ));
 sg13g2_dfrbp_1 _14833_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net977),
    .D(_00280_),
    .Q_N(_07022_),
    .Q(\mem.mem[41][5] ));
 sg13g2_dfrbp_1 _14834_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net976),
    .D(_00281_),
    .Q_N(_07021_),
    .Q(\mem.mem[41][6] ));
 sg13g2_dfrbp_1 _14835_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net975),
    .D(_00282_),
    .Q_N(_07020_),
    .Q(\mem.mem[41][7] ));
 sg13g2_dfrbp_1 _14836_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net974),
    .D(_00283_),
    .Q_N(_07019_),
    .Q(\mem.mem[40][0] ));
 sg13g2_dfrbp_1 _14837_ (.CLK(clknet_leaf_176_clk),
    .RESET_B(net973),
    .D(_00284_),
    .Q_N(_07018_),
    .Q(\mem.mem[40][1] ));
 sg13g2_dfrbp_1 _14838_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net972),
    .D(_00285_),
    .Q_N(_07017_),
    .Q(\mem.mem[40][2] ));
 sg13g2_dfrbp_1 _14839_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net971),
    .D(_00286_),
    .Q_N(_07016_),
    .Q(\mem.mem[40][3] ));
 sg13g2_dfrbp_1 _14840_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net970),
    .D(_00287_),
    .Q_N(_07015_),
    .Q(\mem.mem[40][4] ));
 sg13g2_dfrbp_1 _14841_ (.CLK(clknet_leaf_144_clk),
    .RESET_B(net969),
    .D(_00288_),
    .Q_N(_07014_),
    .Q(\mem.mem[40][5] ));
 sg13g2_dfrbp_1 _14842_ (.CLK(clknet_leaf_145_clk),
    .RESET_B(net968),
    .D(_00289_),
    .Q_N(_07013_),
    .Q(\mem.mem[40][6] ));
 sg13g2_dfrbp_1 _14843_ (.CLK(clknet_leaf_177_clk),
    .RESET_B(net967),
    .D(_00290_),
    .Q_N(_07012_),
    .Q(\mem.mem[40][7] ));
 sg13g2_dfrbp_1 _14844_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net966),
    .D(_00291_),
    .Q_N(_07011_),
    .Q(\mem.mem[199][0] ));
 sg13g2_dfrbp_1 _14845_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net965),
    .D(_00292_),
    .Q_N(_07010_),
    .Q(\mem.mem[199][1] ));
 sg13g2_dfrbp_1 _14846_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net964),
    .D(_00293_),
    .Q_N(_07009_),
    .Q(\mem.mem[199][2] ));
 sg13g2_dfrbp_1 _14847_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net963),
    .D(_00294_),
    .Q_N(_07008_),
    .Q(\mem.mem[199][3] ));
 sg13g2_dfrbp_1 _14848_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net962),
    .D(_00295_),
    .Q_N(_07007_),
    .Q(\mem.mem[199][4] ));
 sg13g2_dfrbp_1 _14849_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net961),
    .D(_00296_),
    .Q_N(_07006_),
    .Q(\mem.mem[199][5] ));
 sg13g2_dfrbp_1 _14850_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net960),
    .D(_00297_),
    .Q_N(_07005_),
    .Q(\mem.mem[199][6] ));
 sg13g2_dfrbp_1 _14851_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net959),
    .D(_00298_),
    .Q_N(_07004_),
    .Q(\mem.mem[199][7] ));
 sg13g2_dfrbp_1 _14852_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net958),
    .D(_00299_),
    .Q_N(_07003_),
    .Q(\mem.mem[3][0] ));
 sg13g2_dfrbp_1 _14853_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net957),
    .D(_00300_),
    .Q_N(_07002_),
    .Q(\mem.mem[3][1] ));
 sg13g2_dfrbp_1 _14854_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net956),
    .D(_00301_),
    .Q_N(_07001_),
    .Q(\mem.mem[3][2] ));
 sg13g2_dfrbp_1 _14855_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net955),
    .D(_00302_),
    .Q_N(_07000_),
    .Q(\mem.mem[3][3] ));
 sg13g2_dfrbp_1 _14856_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net954),
    .D(_00303_),
    .Q_N(_06999_),
    .Q(\mem.mem[3][4] ));
 sg13g2_dfrbp_1 _14857_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net953),
    .D(_00304_),
    .Q_N(_06998_),
    .Q(\mem.mem[3][5] ));
 sg13g2_dfrbp_1 _14858_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net952),
    .D(_00305_),
    .Q_N(_06997_),
    .Q(\mem.mem[3][6] ));
 sg13g2_dfrbp_1 _14859_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net951),
    .D(_00306_),
    .Q_N(_06996_),
    .Q(\mem.mem[3][7] ));
 sg13g2_dfrbp_1 _14860_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net950),
    .D(_00307_),
    .Q_N(_06995_),
    .Q(\mem.mem[38][0] ));
 sg13g2_dfrbp_1 _14861_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net949),
    .D(_00308_),
    .Q_N(_06994_),
    .Q(\mem.mem[38][1] ));
 sg13g2_dfrbp_1 _14862_ (.CLK(clknet_leaf_174_clk),
    .RESET_B(net948),
    .D(_00309_),
    .Q_N(_06993_),
    .Q(\mem.mem[38][2] ));
 sg13g2_dfrbp_1 _14863_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net947),
    .D(_00310_),
    .Q_N(_06992_),
    .Q(\mem.mem[38][3] ));
 sg13g2_dfrbp_1 _14864_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net946),
    .D(_00311_),
    .Q_N(_06991_),
    .Q(\mem.mem[38][4] ));
 sg13g2_dfrbp_1 _14865_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net945),
    .D(_00312_),
    .Q_N(_06990_),
    .Q(\mem.mem[38][5] ));
 sg13g2_dfrbp_1 _14866_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net944),
    .D(_00313_),
    .Q_N(_06989_),
    .Q(\mem.mem[38][6] ));
 sg13g2_dfrbp_1 _14867_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net943),
    .D(_00314_),
    .Q_N(_06988_),
    .Q(\mem.mem[38][7] ));
 sg13g2_dfrbp_1 _14868_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net942),
    .D(_00315_),
    .Q_N(_06987_),
    .Q(\mem.mem[189][0] ));
 sg13g2_dfrbp_1 _14869_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net941),
    .D(_00316_),
    .Q_N(_06986_),
    .Q(\mem.mem[189][1] ));
 sg13g2_dfrbp_1 _14870_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net940),
    .D(_00317_),
    .Q_N(_06985_),
    .Q(\mem.mem[189][2] ));
 sg13g2_dfrbp_1 _14871_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net939),
    .D(_00318_),
    .Q_N(_06984_),
    .Q(\mem.mem[189][3] ));
 sg13g2_dfrbp_1 _14872_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net938),
    .D(_00319_),
    .Q_N(_06983_),
    .Q(\mem.mem[189][4] ));
 sg13g2_dfrbp_1 _14873_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net937),
    .D(_00320_),
    .Q_N(_06982_),
    .Q(\mem.mem[189][5] ));
 sg13g2_dfrbp_1 _14874_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net936),
    .D(_00321_),
    .Q_N(_06981_),
    .Q(\mem.mem[189][6] ));
 sg13g2_dfrbp_1 _14875_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net935),
    .D(_00322_),
    .Q_N(_06980_),
    .Q(\mem.mem[189][7] ));
 sg13g2_dfrbp_1 _14876_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net934),
    .D(_00323_),
    .Q_N(_06979_),
    .Q(_00000_));
 sg13g2_dfrbp_1 _14877_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net933),
    .D(_00324_),
    .Q_N(_06978_),
    .Q(_00001_));
 sg13g2_dfrbp_1 _14878_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net932),
    .D(_00325_),
    .Q_N(_06977_),
    .Q(_00002_));
 sg13g2_dfrbp_1 _14879_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net931),
    .D(_00326_),
    .Q_N(_06976_),
    .Q(_00003_));
 sg13g2_dfrbp_1 _14880_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net930),
    .D(_00327_),
    .Q_N(_06975_),
    .Q(_00004_));
 sg13g2_dfrbp_1 _14881_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net929),
    .D(_00328_),
    .Q_N(_06974_),
    .Q(_00005_));
 sg13g2_dfrbp_1 _14882_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net928),
    .D(_00329_),
    .Q_N(_06973_),
    .Q(_00006_));
 sg13g2_dfrbp_1 _14883_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net927),
    .D(_00330_),
    .Q_N(_06972_),
    .Q(_00007_));
 sg13g2_dfrbp_1 _14884_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net926),
    .D(_00331_),
    .Q_N(_06971_),
    .Q(\mem.mem[37][0] ));
 sg13g2_dfrbp_1 _14885_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net925),
    .D(_00332_),
    .Q_N(_06970_),
    .Q(\mem.mem[37][1] ));
 sg13g2_dfrbp_1 _14886_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net924),
    .D(_00333_),
    .Q_N(_06969_),
    .Q(\mem.mem[37][2] ));
 sg13g2_dfrbp_1 _14887_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net923),
    .D(_00334_),
    .Q_N(_06968_),
    .Q(\mem.mem[37][3] ));
 sg13g2_dfrbp_1 _14888_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net922),
    .D(_00335_),
    .Q_N(_06967_),
    .Q(\mem.mem[37][4] ));
 sg13g2_dfrbp_1 _14889_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net921),
    .D(_00336_),
    .Q_N(_06966_),
    .Q(\mem.mem[37][5] ));
 sg13g2_dfrbp_1 _14890_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net920),
    .D(_00337_),
    .Q_N(_06965_),
    .Q(\mem.mem[37][6] ));
 sg13g2_dfrbp_1 _14891_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net919),
    .D(_00338_),
    .Q_N(_06964_),
    .Q(\mem.mem[37][7] ));
 sg13g2_dfrbp_1 _14892_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net918),
    .D(_00339_),
    .Q_N(_06963_),
    .Q(\mem.mem[53][0] ));
 sg13g2_dfrbp_1 _14893_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net917),
    .D(_00340_),
    .Q_N(_06962_),
    .Q(\mem.mem[53][1] ));
 sg13g2_dfrbp_1 _14894_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net916),
    .D(_00341_),
    .Q_N(_06961_),
    .Q(\mem.mem[53][2] ));
 sg13g2_dfrbp_1 _14895_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net915),
    .D(_00342_),
    .Q_N(_06960_),
    .Q(\mem.mem[53][3] ));
 sg13g2_dfrbp_1 _14896_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net914),
    .D(_00343_),
    .Q_N(_06959_),
    .Q(\mem.mem[53][4] ));
 sg13g2_dfrbp_1 _14897_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net913),
    .D(_00344_),
    .Q_N(_06958_),
    .Q(\mem.mem[53][5] ));
 sg13g2_dfrbp_1 _14898_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net912),
    .D(_00345_),
    .Q_N(_06957_),
    .Q(\mem.mem[53][6] ));
 sg13g2_dfrbp_1 _14899_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net911),
    .D(_00346_),
    .Q_N(_06956_),
    .Q(\mem.mem[53][7] ));
 sg13g2_dfrbp_1 _14900_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net910),
    .D(_00347_),
    .Q_N(_06955_),
    .Q(\mem.mem[36][0] ));
 sg13g2_dfrbp_1 _14901_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net909),
    .D(_00348_),
    .Q_N(_06954_),
    .Q(\mem.mem[36][1] ));
 sg13g2_dfrbp_1 _14902_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net908),
    .D(_00349_),
    .Q_N(_06953_),
    .Q(\mem.mem[36][2] ));
 sg13g2_dfrbp_1 _14903_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net907),
    .D(_00350_),
    .Q_N(_06952_),
    .Q(\mem.mem[36][3] ));
 sg13g2_dfrbp_1 _14904_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net906),
    .D(_00351_),
    .Q_N(_06951_),
    .Q(\mem.mem[36][4] ));
 sg13g2_dfrbp_1 _14905_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net905),
    .D(_00352_),
    .Q_N(_06950_),
    .Q(\mem.mem[36][5] ));
 sg13g2_dfrbp_1 _14906_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net904),
    .D(_00353_),
    .Q_N(_06949_),
    .Q(\mem.mem[36][6] ));
 sg13g2_dfrbp_1 _14907_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net903),
    .D(_00354_),
    .Q_N(_06948_),
    .Q(\mem.mem[36][7] ));
 sg13g2_dfrbp_1 _14908_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net902),
    .D(_00355_),
    .Q_N(_06947_),
    .Q(\mem.mem[52][0] ));
 sg13g2_dfrbp_1 _14909_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net901),
    .D(_00356_),
    .Q_N(_06946_),
    .Q(\mem.mem[52][1] ));
 sg13g2_dfrbp_1 _14910_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net900),
    .D(_00357_),
    .Q_N(_06945_),
    .Q(\mem.mem[52][2] ));
 sg13g2_dfrbp_1 _14911_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net899),
    .D(_00358_),
    .Q_N(_06944_),
    .Q(\mem.mem[52][3] ));
 sg13g2_dfrbp_1 _14912_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net898),
    .D(_00359_),
    .Q_N(_06943_),
    .Q(\mem.mem[52][4] ));
 sg13g2_dfrbp_1 _14913_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net897),
    .D(_00360_),
    .Q_N(_06942_),
    .Q(\mem.mem[52][5] ));
 sg13g2_dfrbp_1 _14914_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net896),
    .D(_00361_),
    .Q_N(_06941_),
    .Q(\mem.mem[52][6] ));
 sg13g2_dfrbp_1 _14915_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net895),
    .D(_00362_),
    .Q_N(_06940_),
    .Q(\mem.mem[52][7] ));
 sg13g2_dfrbp_1 _14916_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net894),
    .D(_00363_),
    .Q_N(_06939_),
    .Q(\mem.mem[35][0] ));
 sg13g2_dfrbp_1 _14917_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net893),
    .D(_00364_),
    .Q_N(_06938_),
    .Q(\mem.mem[35][1] ));
 sg13g2_dfrbp_1 _14918_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net892),
    .D(_00365_),
    .Q_N(_06937_),
    .Q(\mem.mem[35][2] ));
 sg13g2_dfrbp_1 _14919_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net891),
    .D(_00366_),
    .Q_N(_06936_),
    .Q(\mem.mem[35][3] ));
 sg13g2_dfrbp_1 _14920_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net890),
    .D(_00367_),
    .Q_N(_06935_),
    .Q(\mem.mem[35][4] ));
 sg13g2_dfrbp_1 _14921_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net889),
    .D(_00368_),
    .Q_N(_06934_),
    .Q(\mem.mem[35][5] ));
 sg13g2_dfrbp_1 _14922_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net888),
    .D(_00369_),
    .Q_N(_06933_),
    .Q(\mem.mem[35][6] ));
 sg13g2_dfrbp_1 _14923_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net887),
    .D(_00370_),
    .Q_N(_06932_),
    .Q(\mem.mem[35][7] ));
 sg13g2_dfrbp_1 _14924_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net886),
    .D(_00371_),
    .Q_N(_06931_),
    .Q(\mem.mem[51][0] ));
 sg13g2_dfrbp_1 _14925_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net885),
    .D(_00372_),
    .Q_N(_06930_),
    .Q(\mem.mem[51][1] ));
 sg13g2_dfrbp_1 _14926_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net884),
    .D(_00373_),
    .Q_N(_06929_),
    .Q(\mem.mem[51][2] ));
 sg13g2_dfrbp_1 _14927_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net883),
    .D(_00374_),
    .Q_N(_06928_),
    .Q(\mem.mem[51][3] ));
 sg13g2_dfrbp_1 _14928_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net882),
    .D(_00375_),
    .Q_N(_06927_),
    .Q(\mem.mem[51][4] ));
 sg13g2_dfrbp_1 _14929_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net881),
    .D(_00376_),
    .Q_N(_06926_),
    .Q(\mem.mem[51][5] ));
 sg13g2_dfrbp_1 _14930_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net880),
    .D(_00377_),
    .Q_N(_06925_),
    .Q(\mem.mem[51][6] ));
 sg13g2_dfrbp_1 _14931_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net879),
    .D(_00378_),
    .Q_N(_06924_),
    .Q(\mem.mem[51][7] ));
 sg13g2_dfrbp_1 _14932_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net878),
    .D(_00379_),
    .Q_N(_06923_),
    .Q(\mem.mem[71][0] ));
 sg13g2_dfrbp_1 _14933_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net877),
    .D(_00380_),
    .Q_N(_06922_),
    .Q(\mem.mem[71][1] ));
 sg13g2_dfrbp_1 _14934_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net876),
    .D(_00381_),
    .Q_N(_06921_),
    .Q(\mem.mem[71][2] ));
 sg13g2_dfrbp_1 _14935_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net875),
    .D(_00382_),
    .Q_N(_06920_),
    .Q(\mem.mem[71][3] ));
 sg13g2_dfrbp_1 _14936_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net874),
    .D(_00383_),
    .Q_N(_06919_),
    .Q(\mem.mem[71][4] ));
 sg13g2_dfrbp_1 _14937_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net873),
    .D(_00384_),
    .Q_N(_06918_),
    .Q(\mem.mem[71][5] ));
 sg13g2_dfrbp_1 _14938_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net872),
    .D(_00385_),
    .Q_N(_06917_),
    .Q(\mem.mem[71][6] ));
 sg13g2_dfrbp_1 _14939_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net871),
    .D(_00386_),
    .Q_N(_06916_),
    .Q(\mem.mem[71][7] ));
 sg13g2_dfrbp_1 _14940_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net870),
    .D(_00387_),
    .Q_N(_06915_),
    .Q(\mem.mem[91][0] ));
 sg13g2_dfrbp_1 _14941_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net869),
    .D(_00388_),
    .Q_N(_06914_),
    .Q(\mem.mem[91][1] ));
 sg13g2_dfrbp_1 _14942_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net868),
    .D(_00389_),
    .Q_N(_06913_),
    .Q(\mem.mem[91][2] ));
 sg13g2_dfrbp_1 _14943_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net867),
    .D(_00390_),
    .Q_N(_06912_),
    .Q(\mem.mem[91][3] ));
 sg13g2_dfrbp_1 _14944_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net866),
    .D(_00391_),
    .Q_N(_06911_),
    .Q(\mem.mem[91][4] ));
 sg13g2_dfrbp_1 _14945_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net865),
    .D(_00392_),
    .Q_N(_06910_),
    .Q(\mem.mem[91][5] ));
 sg13g2_dfrbp_1 _14946_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net864),
    .D(_00393_),
    .Q_N(_06909_),
    .Q(\mem.mem[91][6] ));
 sg13g2_dfrbp_1 _14947_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net863),
    .D(_00394_),
    .Q_N(_06908_),
    .Q(\mem.mem[91][7] ));
 sg13g2_dfrbp_1 _14948_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net862),
    .D(_00395_),
    .Q_N(_06907_),
    .Q(\mem.mem[70][0] ));
 sg13g2_dfrbp_1 _14949_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net861),
    .D(_00396_),
    .Q_N(_06906_),
    .Q(\mem.mem[70][1] ));
 sg13g2_dfrbp_1 _14950_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net860),
    .D(_00397_),
    .Q_N(_06905_),
    .Q(\mem.mem[70][2] ));
 sg13g2_dfrbp_1 _14951_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net859),
    .D(_00398_),
    .Q_N(_06904_),
    .Q(\mem.mem[70][3] ));
 sg13g2_dfrbp_1 _14952_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net858),
    .D(_00399_),
    .Q_N(_06903_),
    .Q(\mem.mem[70][4] ));
 sg13g2_dfrbp_1 _14953_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net857),
    .D(_00400_),
    .Q_N(_06902_),
    .Q(\mem.mem[70][5] ));
 sg13g2_dfrbp_1 _14954_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net856),
    .D(_00401_),
    .Q_N(_06901_),
    .Q(\mem.mem[70][6] ));
 sg13g2_dfrbp_1 _14955_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net855),
    .D(_00402_),
    .Q_N(_06900_),
    .Q(\mem.mem[70][7] ));
 sg13g2_dfrbp_1 _14956_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net854),
    .D(_00403_),
    .Q_N(_06899_),
    .Q(\mem.mem[6][0] ));
 sg13g2_dfrbp_1 _14957_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net853),
    .D(_00404_),
    .Q_N(_06898_),
    .Q(\mem.mem[6][1] ));
 sg13g2_dfrbp_1 _14958_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net852),
    .D(_00405_),
    .Q_N(_06897_),
    .Q(\mem.mem[6][2] ));
 sg13g2_dfrbp_1 _14959_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net851),
    .D(_00406_),
    .Q_N(_06896_),
    .Q(\mem.mem[6][3] ));
 sg13g2_dfrbp_1 _14960_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net850),
    .D(_00407_),
    .Q_N(_06895_),
    .Q(\mem.mem[6][4] ));
 sg13g2_dfrbp_1 _14961_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net849),
    .D(_00408_),
    .Q_N(_06894_),
    .Q(\mem.mem[6][5] ));
 sg13g2_dfrbp_1 _14962_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net848),
    .D(_00409_),
    .Q_N(_06893_),
    .Q(\mem.mem[6][6] ));
 sg13g2_dfrbp_1 _14963_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net847),
    .D(_00410_),
    .Q_N(_06892_),
    .Q(\mem.mem[6][7] ));
 sg13g2_dfrbp_1 _14964_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net846),
    .D(_00411_),
    .Q_N(_06891_),
    .Q(\mem.mem[90][0] ));
 sg13g2_dfrbp_1 _14965_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net845),
    .D(_00412_),
    .Q_N(_06890_),
    .Q(\mem.mem[90][1] ));
 sg13g2_dfrbp_1 _14966_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net844),
    .D(_00413_),
    .Q_N(_06889_),
    .Q(\mem.mem[90][2] ));
 sg13g2_dfrbp_1 _14967_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net843),
    .D(_00414_),
    .Q_N(_06888_),
    .Q(\mem.mem[90][3] ));
 sg13g2_dfrbp_1 _14968_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net842),
    .D(_00415_),
    .Q_N(_06887_),
    .Q(\mem.mem[90][4] ));
 sg13g2_dfrbp_1 _14969_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net841),
    .D(_00416_),
    .Q_N(_06886_),
    .Q(\mem.mem[90][5] ));
 sg13g2_dfrbp_1 _14970_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net840),
    .D(_00417_),
    .Q_N(_06885_),
    .Q(\mem.mem[90][6] ));
 sg13g2_dfrbp_1 _14971_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net839),
    .D(_00418_),
    .Q_N(_06884_),
    .Q(\mem.mem[90][7] ));
 sg13g2_dfrbp_1 _14972_ (.CLK(clknet_leaf_43_clk),
    .RESET_B(net838),
    .D(_00419_),
    .Q_N(_06883_),
    .Q(\mem.mem[68][0] ));
 sg13g2_dfrbp_1 _14973_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net837),
    .D(_00420_),
    .Q_N(_06882_),
    .Q(\mem.mem[68][1] ));
 sg13g2_dfrbp_1 _14974_ (.CLK(clknet_leaf_47_clk),
    .RESET_B(net836),
    .D(_00421_),
    .Q_N(_06881_),
    .Q(\mem.mem[68][2] ));
 sg13g2_dfrbp_1 _14975_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net835),
    .D(_00422_),
    .Q_N(_06880_),
    .Q(\mem.mem[68][3] ));
 sg13g2_dfrbp_1 _14976_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net834),
    .D(_00423_),
    .Q_N(_06879_),
    .Q(\mem.mem[68][4] ));
 sg13g2_dfrbp_1 _14977_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net833),
    .D(_00424_),
    .Q_N(_06878_),
    .Q(\mem.mem[68][5] ));
 sg13g2_dfrbp_1 _14978_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net832),
    .D(_00425_),
    .Q_N(_06877_),
    .Q(\mem.mem[68][6] ));
 sg13g2_dfrbp_1 _14979_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net831),
    .D(_00426_),
    .Q_N(_06876_),
    .Q(\mem.mem[68][7] ));
 sg13g2_dfrbp_1 _14980_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net830),
    .D(_00427_),
    .Q_N(_06875_),
    .Q(\mem.mem[67][0] ));
 sg13g2_dfrbp_1 _14981_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net829),
    .D(_00428_),
    .Q_N(_06874_),
    .Q(\mem.mem[67][1] ));
 sg13g2_dfrbp_1 _14982_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net828),
    .D(_00429_),
    .Q_N(_06873_),
    .Q(\mem.mem[67][2] ));
 sg13g2_dfrbp_1 _14983_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net827),
    .D(_00430_),
    .Q_N(_06872_),
    .Q(\mem.mem[67][3] ));
 sg13g2_dfrbp_1 _14984_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net826),
    .D(_00431_),
    .Q_N(_06871_),
    .Q(\mem.mem[67][4] ));
 sg13g2_dfrbp_1 _14985_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net825),
    .D(_00432_),
    .Q_N(_06870_),
    .Q(\mem.mem[67][5] ));
 sg13g2_dfrbp_1 _14986_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net824),
    .D(_00433_),
    .Q_N(_06869_),
    .Q(\mem.mem[67][6] ));
 sg13g2_dfrbp_1 _14987_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net823),
    .D(_00434_),
    .Q_N(_06868_),
    .Q(\mem.mem[67][7] ));
 sg13g2_dfrbp_1 _14988_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net822),
    .D(_00435_),
    .Q_N(_06867_),
    .Q(\mem.mem[8][0] ));
 sg13g2_dfrbp_1 _14989_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net821),
    .D(_00436_),
    .Q_N(_06866_),
    .Q(\mem.mem[8][1] ));
 sg13g2_dfrbp_1 _14990_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net820),
    .D(_00437_),
    .Q_N(_06865_),
    .Q(\mem.mem[8][2] ));
 sg13g2_dfrbp_1 _14991_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net819),
    .D(_00438_),
    .Q_N(_06864_),
    .Q(\mem.mem[8][3] ));
 sg13g2_dfrbp_1 _14992_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net818),
    .D(_00439_),
    .Q_N(_06863_),
    .Q(\mem.mem[8][4] ));
 sg13g2_dfrbp_1 _14993_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net817),
    .D(_00440_),
    .Q_N(_06862_),
    .Q(\mem.mem[8][5] ));
 sg13g2_dfrbp_1 _14994_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net816),
    .D(_00441_),
    .Q_N(_06861_),
    .Q(\mem.mem[8][6] ));
 sg13g2_dfrbp_1 _14995_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net815),
    .D(_00442_),
    .Q_N(_06860_),
    .Q(\mem.mem[8][7] ));
 sg13g2_dfrbp_1 _14996_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net814),
    .D(_00443_),
    .Q_N(_06859_),
    .Q(\mem.mem[66][0] ));
 sg13g2_dfrbp_1 _14997_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net813),
    .D(_00444_),
    .Q_N(_06858_),
    .Q(\mem.mem[66][1] ));
 sg13g2_dfrbp_1 _14998_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net812),
    .D(_00445_),
    .Q_N(_06857_),
    .Q(\mem.mem[66][2] ));
 sg13g2_dfrbp_1 _14999_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net811),
    .D(_00446_),
    .Q_N(_06856_),
    .Q(\mem.mem[66][3] ));
 sg13g2_dfrbp_1 _15000_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net810),
    .D(_00447_),
    .Q_N(_06855_),
    .Q(\mem.mem[66][4] ));
 sg13g2_dfrbp_1 _15001_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net809),
    .D(_00448_),
    .Q_N(_06854_),
    .Q(\mem.mem[66][5] ));
 sg13g2_dfrbp_1 _15002_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net808),
    .D(_00449_),
    .Q_N(_06853_),
    .Q(\mem.mem[66][6] ));
 sg13g2_dfrbp_1 _15003_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net807),
    .D(_00450_),
    .Q_N(_06852_),
    .Q(\mem.mem[66][7] ));
 sg13g2_dfrbp_1 _15004_ (.CLK(clknet_leaf_48_clk),
    .RESET_B(net806),
    .D(_00451_),
    .Q_N(_06851_),
    .Q(\mem.mem[65][0] ));
 sg13g2_dfrbp_1 _15005_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net805),
    .D(_00452_),
    .Q_N(_06850_),
    .Q(\mem.mem[65][1] ));
 sg13g2_dfrbp_1 _15006_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net804),
    .D(_00453_),
    .Q_N(_06849_),
    .Q(\mem.mem[65][2] ));
 sg13g2_dfrbp_1 _15007_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net803),
    .D(_00454_),
    .Q_N(_06848_),
    .Q(\mem.mem[65][3] ));
 sg13g2_dfrbp_1 _15008_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net802),
    .D(_00455_),
    .Q_N(_06847_),
    .Q(\mem.mem[65][4] ));
 sg13g2_dfrbp_1 _15009_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net801),
    .D(_00456_),
    .Q_N(_06846_),
    .Q(\mem.mem[65][5] ));
 sg13g2_dfrbp_1 _15010_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net800),
    .D(_00457_),
    .Q_N(_06845_),
    .Q(\mem.mem[65][6] ));
 sg13g2_dfrbp_1 _15011_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net799),
    .D(_00458_),
    .Q_N(_06844_),
    .Q(\mem.mem[65][7] ));
 sg13g2_dfrbp_1 _15012_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net798),
    .D(_00459_),
    .Q_N(_06843_),
    .Q(\mem.mem[88][0] ));
 sg13g2_dfrbp_1 _15013_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net797),
    .D(_00460_),
    .Q_N(_06842_),
    .Q(\mem.mem[88][1] ));
 sg13g2_dfrbp_1 _15014_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net796),
    .D(_00461_),
    .Q_N(_06841_),
    .Q(\mem.mem[88][2] ));
 sg13g2_dfrbp_1 _15015_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net795),
    .D(_00462_),
    .Q_N(_06840_),
    .Q(\mem.mem[88][3] ));
 sg13g2_dfrbp_1 _15016_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net794),
    .D(_00463_),
    .Q_N(_06839_),
    .Q(\mem.mem[88][4] ));
 sg13g2_dfrbp_1 _15017_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net793),
    .D(_00464_),
    .Q_N(_06838_),
    .Q(\mem.mem[88][5] ));
 sg13g2_dfrbp_1 _15018_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net792),
    .D(_00465_),
    .Q_N(_06837_),
    .Q(\mem.mem[88][6] ));
 sg13g2_dfrbp_1 _15019_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net791),
    .D(_00466_),
    .Q_N(_06836_),
    .Q(\mem.mem[88][7] ));
 sg13g2_dfrbp_1 _15020_ (.CLK(clknet_leaf_46_clk),
    .RESET_B(net790),
    .D(_00467_),
    .Q_N(_06835_),
    .Q(\mem.mem[64][0] ));
 sg13g2_dfrbp_1 _15021_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net789),
    .D(_00468_),
    .Q_N(_06834_),
    .Q(\mem.mem[64][1] ));
 sg13g2_dfrbp_1 _15022_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net788),
    .D(_00469_),
    .Q_N(_06833_),
    .Q(\mem.mem[64][2] ));
 sg13g2_dfrbp_1 _15023_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net787),
    .D(_00470_),
    .Q_N(_06832_),
    .Q(\mem.mem[64][3] ));
 sg13g2_dfrbp_1 _15024_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net786),
    .D(_00471_),
    .Q_N(_06831_),
    .Q(\mem.mem[64][4] ));
 sg13g2_dfrbp_1 _15025_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net785),
    .D(_00472_),
    .Q_N(_06830_),
    .Q(\mem.mem[64][5] ));
 sg13g2_dfrbp_1 _15026_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net784),
    .D(_00473_),
    .Q_N(_06829_),
    .Q(\mem.mem[64][6] ));
 sg13g2_dfrbp_1 _15027_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net783),
    .D(_00474_),
    .Q_N(_06828_),
    .Q(\mem.mem[64][7] ));
 sg13g2_dfrbp_1 _15028_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net782),
    .D(_00475_),
    .Q_N(_06827_),
    .Q(\mem.mem[63][0] ));
 sg13g2_dfrbp_1 _15029_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net781),
    .D(_00476_),
    .Q_N(_06826_),
    .Q(\mem.mem[63][1] ));
 sg13g2_dfrbp_1 _15030_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net780),
    .D(_00477_),
    .Q_N(_06825_),
    .Q(\mem.mem[63][2] ));
 sg13g2_dfrbp_1 _15031_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net779),
    .D(_00478_),
    .Q_N(_06824_),
    .Q(\mem.mem[63][3] ));
 sg13g2_dfrbp_1 _15032_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net778),
    .D(_00479_),
    .Q_N(_06823_),
    .Q(\mem.mem[63][4] ));
 sg13g2_dfrbp_1 _15033_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net777),
    .D(_00480_),
    .Q_N(_06822_),
    .Q(\mem.mem[63][5] ));
 sg13g2_dfrbp_1 _15034_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net776),
    .D(_00481_),
    .Q_N(_06821_),
    .Q(\mem.mem[63][6] ));
 sg13g2_dfrbp_1 _15035_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net775),
    .D(_00482_),
    .Q_N(_06820_),
    .Q(\mem.mem[63][7] ));
 sg13g2_dfrbp_1 _15036_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net774),
    .D(_00483_),
    .Q_N(_06819_),
    .Q(\mem.mem[87][0] ));
 sg13g2_dfrbp_1 _15037_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net773),
    .D(_00484_),
    .Q_N(_06818_),
    .Q(\mem.mem[87][1] ));
 sg13g2_dfrbp_1 _15038_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net772),
    .D(_00485_),
    .Q_N(_06817_),
    .Q(\mem.mem[87][2] ));
 sg13g2_dfrbp_1 _15039_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net771),
    .D(_00486_),
    .Q_N(_06816_),
    .Q(\mem.mem[87][3] ));
 sg13g2_dfrbp_1 _15040_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net770),
    .D(_00487_),
    .Q_N(_06815_),
    .Q(\mem.mem[87][4] ));
 sg13g2_dfrbp_1 _15041_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net769),
    .D(_00488_),
    .Q_N(_06814_),
    .Q(\mem.mem[87][5] ));
 sg13g2_dfrbp_1 _15042_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net768),
    .D(_00489_),
    .Q_N(_06813_),
    .Q(\mem.mem[87][6] ));
 sg13g2_dfrbp_1 _15043_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net767),
    .D(_00490_),
    .Q_N(_06812_),
    .Q(\mem.mem[87][7] ));
 sg13g2_dfrbp_1 _15044_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net766),
    .D(_00491_),
    .Q_N(_06811_),
    .Q(\mem.mem[62][0] ));
 sg13g2_dfrbp_1 _15045_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net765),
    .D(_00492_),
    .Q_N(_06810_),
    .Q(\mem.mem[62][1] ));
 sg13g2_dfrbp_1 _15046_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net764),
    .D(_00493_),
    .Q_N(_06809_),
    .Q(\mem.mem[62][2] ));
 sg13g2_dfrbp_1 _15047_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net763),
    .D(_00494_),
    .Q_N(_06808_),
    .Q(\mem.mem[62][3] ));
 sg13g2_dfrbp_1 _15048_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net762),
    .D(_00495_),
    .Q_N(_06807_),
    .Q(\mem.mem[62][4] ));
 sg13g2_dfrbp_1 _15049_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net761),
    .D(_00496_),
    .Q_N(_06806_),
    .Q(\mem.mem[62][5] ));
 sg13g2_dfrbp_1 _15050_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net760),
    .D(_00497_),
    .Q_N(_06805_),
    .Q(\mem.mem[62][6] ));
 sg13g2_dfrbp_1 _15051_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net759),
    .D(_00498_),
    .Q_N(_06804_),
    .Q(\mem.mem[62][7] ));
 sg13g2_dfrbp_1 _15052_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net758),
    .D(_00499_),
    .Q_N(_06803_),
    .Q(\mem.mem[61][0] ));
 sg13g2_dfrbp_1 _15053_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net757),
    .D(_00500_),
    .Q_N(_06802_),
    .Q(\mem.mem[61][1] ));
 sg13g2_dfrbp_1 _15054_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net756),
    .D(_00501_),
    .Q_N(_06801_),
    .Q(\mem.mem[61][2] ));
 sg13g2_dfrbp_1 _15055_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net755),
    .D(_00502_),
    .Q_N(_06800_),
    .Q(\mem.mem[61][3] ));
 sg13g2_dfrbp_1 _15056_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net754),
    .D(_00503_),
    .Q_N(_06799_),
    .Q(\mem.mem[61][4] ));
 sg13g2_dfrbp_1 _15057_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net753),
    .D(_00504_),
    .Q_N(_06798_),
    .Q(\mem.mem[61][5] ));
 sg13g2_dfrbp_1 _15058_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net752),
    .D(_00505_),
    .Q_N(_06797_),
    .Q(\mem.mem[61][6] ));
 sg13g2_dfrbp_1 _15059_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net751),
    .D(_00506_),
    .Q_N(_06796_),
    .Q(\mem.mem[61][7] ));
 sg13g2_dfrbp_1 _15060_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net750),
    .D(_00507_),
    .Q_N(_06795_),
    .Q(\mem.mem[86][0] ));
 sg13g2_dfrbp_1 _15061_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net749),
    .D(_00508_),
    .Q_N(_06794_),
    .Q(\mem.mem[86][1] ));
 sg13g2_dfrbp_1 _15062_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net748),
    .D(_00509_),
    .Q_N(_06793_),
    .Q(\mem.mem[86][2] ));
 sg13g2_dfrbp_1 _15063_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net747),
    .D(_00510_),
    .Q_N(_06792_),
    .Q(\mem.mem[86][3] ));
 sg13g2_dfrbp_1 _15064_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net746),
    .D(_00511_),
    .Q_N(_06791_),
    .Q(\mem.mem[86][4] ));
 sg13g2_dfrbp_1 _15065_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net745),
    .D(_00512_),
    .Q_N(_06790_),
    .Q(\mem.mem[86][5] ));
 sg13g2_dfrbp_1 _15066_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net744),
    .D(_00513_),
    .Q_N(_06789_),
    .Q(\mem.mem[86][6] ));
 sg13g2_dfrbp_1 _15067_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net743),
    .D(_00514_),
    .Q_N(_06788_),
    .Q(\mem.mem[86][7] ));
 sg13g2_dfrbp_1 _15068_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net742),
    .D(_00515_),
    .Q_N(_06787_),
    .Q(\mem.mem[60][0] ));
 sg13g2_dfrbp_1 _15069_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net741),
    .D(_00516_),
    .Q_N(_06786_),
    .Q(\mem.mem[60][1] ));
 sg13g2_dfrbp_1 _15070_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net740),
    .D(_00517_),
    .Q_N(_06785_),
    .Q(\mem.mem[60][2] ));
 sg13g2_dfrbp_1 _15071_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net739),
    .D(_00518_),
    .Q_N(_06784_),
    .Q(\mem.mem[60][3] ));
 sg13g2_dfrbp_1 _15072_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net738),
    .D(_00519_),
    .Q_N(_06783_),
    .Q(\mem.mem[60][4] ));
 sg13g2_dfrbp_1 _15073_ (.CLK(clknet_leaf_132_clk),
    .RESET_B(net737),
    .D(_00520_),
    .Q_N(_06782_),
    .Q(\mem.mem[60][5] ));
 sg13g2_dfrbp_1 _15074_ (.CLK(clknet_leaf_133_clk),
    .RESET_B(net736),
    .D(_00521_),
    .Q_N(_06781_),
    .Q(\mem.mem[60][6] ));
 sg13g2_dfrbp_1 _15075_ (.CLK(clknet_leaf_131_clk),
    .RESET_B(net735),
    .D(_00522_),
    .Q_N(_06780_),
    .Q(\mem.mem[60][7] ));
 sg13g2_dfrbp_1 _15076_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net734),
    .D(_00523_),
    .Q_N(_06779_),
    .Q(\mem.mem[5][0] ));
 sg13g2_dfrbp_1 _15077_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net733),
    .D(_00524_),
    .Q_N(_06778_),
    .Q(\mem.mem[5][1] ));
 sg13g2_dfrbp_1 _15078_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net732),
    .D(_00525_),
    .Q_N(_06777_),
    .Q(\mem.mem[5][2] ));
 sg13g2_dfrbp_1 _15079_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net731),
    .D(_00526_),
    .Q_N(_06776_),
    .Q(\mem.mem[5][3] ));
 sg13g2_dfrbp_1 _15080_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net730),
    .D(_00527_),
    .Q_N(_06775_),
    .Q(\mem.mem[5][4] ));
 sg13g2_dfrbp_1 _15081_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net729),
    .D(_00528_),
    .Q_N(_06774_),
    .Q(\mem.mem[5][5] ));
 sg13g2_dfrbp_1 _15082_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net728),
    .D(_00529_),
    .Q_N(_06773_),
    .Q(\mem.mem[5][6] ));
 sg13g2_dfrbp_1 _15083_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net727),
    .D(_00530_),
    .Q_N(_06772_),
    .Q(\mem.mem[5][7] ));
 sg13g2_dfrbp_1 _15084_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net726),
    .D(_00531_),
    .Q_N(_06771_),
    .Q(\mem.mem[85][0] ));
 sg13g2_dfrbp_1 _15085_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net725),
    .D(_00532_),
    .Q_N(_06770_),
    .Q(\mem.mem[85][1] ));
 sg13g2_dfrbp_1 _15086_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net724),
    .D(_00533_),
    .Q_N(_06769_),
    .Q(\mem.mem[85][2] ));
 sg13g2_dfrbp_1 _15087_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net723),
    .D(_00534_),
    .Q_N(_06768_),
    .Q(\mem.mem[85][3] ));
 sg13g2_dfrbp_1 _15088_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net722),
    .D(_00535_),
    .Q_N(_06767_),
    .Q(\mem.mem[85][4] ));
 sg13g2_dfrbp_1 _15089_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net721),
    .D(_00536_),
    .Q_N(_06766_),
    .Q(\mem.mem[85][5] ));
 sg13g2_dfrbp_1 _15090_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net720),
    .D(_00537_),
    .Q_N(_06765_),
    .Q(\mem.mem[85][6] ));
 sg13g2_dfrbp_1 _15091_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net719),
    .D(_00538_),
    .Q_N(_06764_),
    .Q(\mem.mem[85][7] ));
 sg13g2_dfrbp_1 _15092_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net718),
    .D(_00539_),
    .Q_N(_06763_),
    .Q(\mem.mem[58][0] ));
 sg13g2_dfrbp_1 _15093_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net717),
    .D(_00540_),
    .Q_N(_06762_),
    .Q(\mem.mem[58][1] ));
 sg13g2_dfrbp_1 _15094_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net716),
    .D(_00541_),
    .Q_N(_06761_),
    .Q(\mem.mem[58][2] ));
 sg13g2_dfrbp_1 _15095_ (.CLK(clknet_leaf_143_clk),
    .RESET_B(net715),
    .D(_00542_),
    .Q_N(_06760_),
    .Q(\mem.mem[58][3] ));
 sg13g2_dfrbp_1 _15096_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net714),
    .D(_00543_),
    .Q_N(_06759_),
    .Q(\mem.mem[58][4] ));
 sg13g2_dfrbp_1 _15097_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net713),
    .D(_00544_),
    .Q_N(_06758_),
    .Q(\mem.mem[58][5] ));
 sg13g2_dfrbp_1 _15098_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net712),
    .D(_00545_),
    .Q_N(_06757_),
    .Q(\mem.mem[58][6] ));
 sg13g2_dfrbp_1 _15099_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net711),
    .D(_00546_),
    .Q_N(_06756_),
    .Q(\mem.mem[58][7] ));
 sg13g2_dfrbp_1 _15100_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net710),
    .D(_00547_),
    .Q_N(_06755_),
    .Q(\mem.mem[57][0] ));
 sg13g2_dfrbp_1 _15101_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net709),
    .D(_00548_),
    .Q_N(_06754_),
    .Q(\mem.mem[57][1] ));
 sg13g2_dfrbp_1 _15102_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net708),
    .D(_00549_),
    .Q_N(_06753_),
    .Q(\mem.mem[57][2] ));
 sg13g2_dfrbp_1 _15103_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net707),
    .D(_00550_),
    .Q_N(_06752_),
    .Q(\mem.mem[57][3] ));
 sg13g2_dfrbp_1 _15104_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net706),
    .D(_00551_),
    .Q_N(_06751_),
    .Q(\mem.mem[57][4] ));
 sg13g2_dfrbp_1 _15105_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net705),
    .D(_00552_),
    .Q_N(_06750_),
    .Q(\mem.mem[57][5] ));
 sg13g2_dfrbp_1 _15106_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net704),
    .D(_00553_),
    .Q_N(_06749_),
    .Q(\mem.mem[57][6] ));
 sg13g2_dfrbp_1 _15107_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net703),
    .D(_00554_),
    .Q_N(_06748_),
    .Q(\mem.mem[57][7] ));
 sg13g2_dfrbp_1 _15108_ (.CLK(clknet_leaf_56_clk),
    .RESET_B(net702),
    .D(_00555_),
    .Q_N(_06747_),
    .Q(\mem.mem[84][0] ));
 sg13g2_dfrbp_1 _15109_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net701),
    .D(_00556_),
    .Q_N(_06746_),
    .Q(\mem.mem[84][1] ));
 sg13g2_dfrbp_1 _15110_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net700),
    .D(_00557_),
    .Q_N(_06745_),
    .Q(\mem.mem[84][2] ));
 sg13g2_dfrbp_1 _15111_ (.CLK(clknet_leaf_55_clk),
    .RESET_B(net699),
    .D(_00558_),
    .Q_N(_06744_),
    .Q(\mem.mem[84][3] ));
 sg13g2_dfrbp_1 _15112_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net698),
    .D(_00559_),
    .Q_N(_06743_),
    .Q(\mem.mem[84][4] ));
 sg13g2_dfrbp_1 _15113_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net697),
    .D(_00560_),
    .Q_N(_06742_),
    .Q(\mem.mem[84][5] ));
 sg13g2_dfrbp_1 _15114_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net696),
    .D(_00561_),
    .Q_N(_06741_),
    .Q(\mem.mem[84][6] ));
 sg13g2_dfrbp_1 _15115_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net695),
    .D(_00562_),
    .Q_N(_06740_),
    .Q(\mem.mem[84][7] ));
 sg13g2_dfrbp_1 _15116_ (.CLK(clknet_leaf_142_clk),
    .RESET_B(net694),
    .D(_00563_),
    .Q_N(_06739_),
    .Q(\mem.mem[56][0] ));
 sg13g2_dfrbp_1 _15117_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net693),
    .D(_00564_),
    .Q_N(_06738_),
    .Q(\mem.mem[56][1] ));
 sg13g2_dfrbp_1 _15118_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net692),
    .D(_00565_),
    .Q_N(_06737_),
    .Q(\mem.mem[56][2] ));
 sg13g2_dfrbp_1 _15119_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net691),
    .D(_00566_),
    .Q_N(_06736_),
    .Q(\mem.mem[56][3] ));
 sg13g2_dfrbp_1 _15120_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net690),
    .D(_00567_),
    .Q_N(_06735_),
    .Q(\mem.mem[56][4] ));
 sg13g2_dfrbp_1 _15121_ (.CLK(clknet_leaf_140_clk),
    .RESET_B(net689),
    .D(_00568_),
    .Q_N(_06734_),
    .Q(\mem.mem[56][5] ));
 sg13g2_dfrbp_1 _15122_ (.CLK(clknet_leaf_139_clk),
    .RESET_B(net688),
    .D(_00569_),
    .Q_N(_06733_),
    .Q(\mem.mem[56][6] ));
 sg13g2_dfrbp_1 _15123_ (.CLK(clknet_leaf_141_clk),
    .RESET_B(net687),
    .D(_00570_),
    .Q_N(_06732_),
    .Q(\mem.mem[56][7] ));
 sg13g2_dfrbp_1 _15124_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net686),
    .D(_00571_),
    .Q_N(_06731_),
    .Q(\mem.mem[55][0] ));
 sg13g2_dfrbp_1 _15125_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net685),
    .D(_00572_),
    .Q_N(_06730_),
    .Q(\mem.mem[55][1] ));
 sg13g2_dfrbp_1 _15126_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net684),
    .D(_00573_),
    .Q_N(_06729_),
    .Q(\mem.mem[55][2] ));
 sg13g2_dfrbp_1 _15127_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net683),
    .D(_00574_),
    .Q_N(_06728_),
    .Q(\mem.mem[55][3] ));
 sg13g2_dfrbp_1 _15128_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net682),
    .D(_00575_),
    .Q_N(_06727_),
    .Q(\mem.mem[55][4] ));
 sg13g2_dfrbp_1 _15129_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net681),
    .D(_00576_),
    .Q_N(_06726_),
    .Q(\mem.mem[55][5] ));
 sg13g2_dfrbp_1 _15130_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net680),
    .D(_00577_),
    .Q_N(_06725_),
    .Q(\mem.mem[55][6] ));
 sg13g2_dfrbp_1 _15131_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net679),
    .D(_00578_),
    .Q_N(_06724_),
    .Q(\mem.mem[55][7] ));
 sg13g2_dfrbp_1 _15132_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net678),
    .D(_00579_),
    .Q_N(_06723_),
    .Q(\mem.mem[83][0] ));
 sg13g2_dfrbp_1 _15133_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net677),
    .D(_00580_),
    .Q_N(_06722_),
    .Q(\mem.mem[83][1] ));
 sg13g2_dfrbp_1 _15134_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net676),
    .D(_00581_),
    .Q_N(_06721_),
    .Q(\mem.mem[83][2] ));
 sg13g2_dfrbp_1 _15135_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net675),
    .D(_00582_),
    .Q_N(_06720_),
    .Q(\mem.mem[83][3] ));
 sg13g2_dfrbp_1 _15136_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net674),
    .D(_00583_),
    .Q_N(_06719_),
    .Q(\mem.mem[83][4] ));
 sg13g2_dfrbp_1 _15137_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net673),
    .D(_00584_),
    .Q_N(_06718_),
    .Q(\mem.mem[83][5] ));
 sg13g2_dfrbp_1 _15138_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net672),
    .D(_00585_),
    .Q_N(_06717_),
    .Q(\mem.mem[83][6] ));
 sg13g2_dfrbp_1 _15139_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net671),
    .D(_00586_),
    .Q_N(_06716_),
    .Q(\mem.mem[83][7] ));
 sg13g2_dfrbp_1 _15140_ (.CLK(clknet_leaf_138_clk),
    .RESET_B(net670),
    .D(_00587_),
    .Q_N(_06715_),
    .Q(\mem.mem[54][0] ));
 sg13g2_dfrbp_1 _15141_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net669),
    .D(_00588_),
    .Q_N(_06714_),
    .Q(\mem.mem[54][1] ));
 sg13g2_dfrbp_1 _15142_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net668),
    .D(_00589_),
    .Q_N(_06713_),
    .Q(\mem.mem[54][2] ));
 sg13g2_dfrbp_1 _15143_ (.CLK(clknet_leaf_147_clk),
    .RESET_B(net667),
    .D(_00590_),
    .Q_N(_06712_),
    .Q(\mem.mem[54][3] ));
 sg13g2_dfrbp_1 _15144_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net666),
    .D(_00591_),
    .Q_N(_06711_),
    .Q(\mem.mem[54][4] ));
 sg13g2_dfrbp_1 _15145_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net665),
    .D(_00592_),
    .Q_N(_06710_),
    .Q(\mem.mem[54][5] ));
 sg13g2_dfrbp_1 _15146_ (.CLK(clknet_leaf_137_clk),
    .RESET_B(net664),
    .D(_00593_),
    .Q_N(_06709_),
    .Q(\mem.mem[54][6] ));
 sg13g2_dfrbp_1 _15147_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net663),
    .D(_00594_),
    .Q_N(_06708_),
    .Q(\mem.mem[54][7] ));
 sg13g2_dfrbp_1 _15148_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net662),
    .D(_00595_),
    .Q_N(_06707_),
    .Q(\A[0] ));
 sg13g2_dfrbp_1 _15149_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net660),
    .D(net5195),
    .Q_N(_06706_),
    .Q(\A[1] ));
 sg13g2_dfrbp_1 _15150_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net658),
    .D(net2674),
    .Q_N(_06705_),
    .Q(\A[2] ));
 sg13g2_dfrbp_1 _15151_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net656),
    .D(_00598_),
    .Q_N(_06704_),
    .Q(\A[3] ));
 sg13g2_dfrbp_1 _15152_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net654),
    .D(_00599_),
    .Q_N(_06703_),
    .Q(\A[4] ));
 sg13g2_dfrbp_1 _15153_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net652),
    .D(_00600_),
    .Q_N(_06702_),
    .Q(\A[5] ));
 sg13g2_dfrbp_1 _15154_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net650),
    .D(net2783),
    .Q_N(_06701_),
    .Q(\A[6] ));
 sg13g2_dfrbp_1 _15155_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net648),
    .D(net2656),
    .Q_N(_06700_),
    .Q(\A[7] ));
 sg13g2_dfrbp_1 _15156_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net646),
    .D(_00603_),
    .Q_N(_06699_),
    .Q(\B[0] ));
 sg13g2_dfrbp_1 _15157_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net644),
    .D(_00604_),
    .Q_N(_06698_),
    .Q(\B[1] ));
 sg13g2_dfrbp_1 _15158_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net642),
    .D(_00605_),
    .Q_N(_06697_),
    .Q(\B[2] ));
 sg13g2_dfrbp_1 _15159_ (.CLK(clknet_leaf_57_clk),
    .RESET_B(net640),
    .D(_00606_),
    .Q_N(_06696_),
    .Q(\B[3] ));
 sg13g2_dfrbp_1 _15160_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net638),
    .D(_00607_),
    .Q_N(_06695_),
    .Q(\B[4] ));
 sg13g2_dfrbp_1 _15161_ (.CLK(clknet_leaf_58_clk),
    .RESET_B(net636),
    .D(_00608_),
    .Q_N(_06694_),
    .Q(\B[5] ));
 sg13g2_dfrbp_1 _15162_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net634),
    .D(_00609_),
    .Q_N(_06693_),
    .Q(\B[6] ));
 sg13g2_dfrbp_1 _15163_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net632),
    .D(_00610_),
    .Q_N(_06692_),
    .Q(\B[7] ));
 sg13g2_dfrbp_1 _15164_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net630),
    .D(_00611_),
    .Q_N(_06691_),
    .Q(\C[0] ));
 sg13g2_dfrbp_1 _15165_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net628),
    .D(_00612_),
    .Q_N(_06690_),
    .Q(\C[1] ));
 sg13g2_dfrbp_1 _15166_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net626),
    .D(_00613_),
    .Q_N(_00017_),
    .Q(\C[2] ));
 sg13g2_dfrbp_1 _15167_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net624),
    .D(_00614_),
    .Q_N(_00016_),
    .Q(\C[3] ));
 sg13g2_dfrbp_1 _15168_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net622),
    .D(_00615_),
    .Q_N(_00015_),
    .Q(\C[4] ));
 sg13g2_dfrbp_1 _15169_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net620),
    .D(_00616_),
    .Q_N(_00014_),
    .Q(\C[5] ));
 sg13g2_dfrbp_1 _15170_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net618),
    .D(_00617_),
    .Q_N(_00013_),
    .Q(\C[6] ));
 sg13g2_dfrbp_1 _15171_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net616),
    .D(_00618_),
    .Q_N(_00012_),
    .Q(\C[7] ));
 sg13g2_dfrbp_1 _15172_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net614),
    .D(_00619_),
    .Q_N(_06689_),
    .Q(\state[0] ));
 sg13g2_dfrbp_1 _15173_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net612),
    .D(_00620_),
    .Q_N(_06688_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 _15174_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net610),
    .D(net5189),
    .Q_N(_00011_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 _15175_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net608),
    .D(net5214),
    .Q_N(_00010_),
    .Q(\PC[0] ));
 sg13g2_dfrbp_1 _15176_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net606),
    .D(_00623_),
    .Q_N(_06687_),
    .Q(\PC[1] ));
 sg13g2_dfrbp_1 _15177_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net604),
    .D(_00624_),
    .Q_N(_06686_),
    .Q(\PC[2] ));
 sg13g2_dfrbp_1 _15178_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net602),
    .D(_00625_),
    .Q_N(_06685_),
    .Q(\PC[3] ));
 sg13g2_dfrbp_1 _15179_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net600),
    .D(_00626_),
    .Q_N(_06684_),
    .Q(\PC[4] ));
 sg13g2_dfrbp_1 _15180_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net598),
    .D(_00627_),
    .Q_N(_06683_),
    .Q(\PC[5] ));
 sg13g2_dfrbp_1 _15181_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net596),
    .D(_00628_),
    .Q_N(_06682_),
    .Q(\PC[6] ));
 sg13g2_dfrbp_1 _15182_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net594),
    .D(_00629_),
    .Q_N(_06681_),
    .Q(\PC[7] ));
 sg13g2_dfrbp_1 _15183_ (.CLK(clknet_leaf_41_clk),
    .RESET_B(net592),
    .D(_00630_),
    .Q_N(_06680_),
    .Q(\mem.addr[0] ));
 sg13g2_dfrbp_1 _15184_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net590),
    .D(_00631_),
    .Q_N(_06679_),
    .Q(\mem.addr[1] ));
 sg13g2_dfrbp_1 _15185_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net588),
    .D(_00632_),
    .Q_N(_06678_),
    .Q(\mem.addr[2] ));
 sg13g2_dfrbp_1 _15186_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net586),
    .D(_00633_),
    .Q_N(_06677_),
    .Q(\mem.addr[3] ));
 sg13g2_dfrbp_1 _15187_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net584),
    .D(_00634_),
    .Q_N(_06676_),
    .Q(\mem.addr[4] ));
 sg13g2_dfrbp_1 _15188_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net582),
    .D(_00635_),
    .Q_N(_06675_),
    .Q(\mem.addr[5] ));
 sg13g2_dfrbp_1 _15189_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net580),
    .D(_00636_),
    .Q_N(_06674_),
    .Q(\mem.addr[6] ));
 sg13g2_dfrbp_1 _15190_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net578),
    .D(_00637_),
    .Q_N(_06673_),
    .Q(\mem.addr[7] ));
 sg13g2_dfrbp_1 _15191_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net576),
    .D(_00638_),
    .Q_N(_06672_),
    .Q(\mem.data_in[0] ));
 sg13g2_dfrbp_1 _15192_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net574),
    .D(_00639_),
    .Q_N(_06671_),
    .Q(\mem.data_in[1] ));
 sg13g2_dfrbp_1 _15193_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net572),
    .D(_00640_),
    .Q_N(_06670_),
    .Q(\mem.data_in[2] ));
 sg13g2_dfrbp_1 _15194_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net570),
    .D(_00641_),
    .Q_N(_06669_),
    .Q(\mem.data_in[3] ));
 sg13g2_dfrbp_1 _15195_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net568),
    .D(_00642_),
    .Q_N(_06668_),
    .Q(\mem.data_in[4] ));
 sg13g2_dfrbp_1 _15196_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net566),
    .D(_00643_),
    .Q_N(_06667_),
    .Q(\mem.data_in[5] ));
 sg13g2_dfrbp_1 _15197_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net564),
    .D(_00644_),
    .Q_N(_06666_),
    .Q(\mem.data_in[6] ));
 sg13g2_dfrbp_1 _15198_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net562),
    .D(_00645_),
    .Q_N(_06665_),
    .Q(\mem.data_in[7] ));
 sg13g2_dfrbp_1 _15199_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net560),
    .D(_00646_),
    .Q_N(_06664_),
    .Q(\mem_A[0] ));
 sg13g2_dfrbp_1 _15200_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net558),
    .D(_00647_),
    .Q_N(_00009_),
    .Q(\mem_A[1] ));
 sg13g2_dfrbp_1 _15201_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net556),
    .D(net4851),
    .Q_N(_06663_),
    .Q(\mem_A[2] ));
 sg13g2_dfrbp_1 _15202_ (.CLK(clknet_leaf_74_clk),
    .RESET_B(net554),
    .D(_00649_),
    .Q_N(_06662_),
    .Q(\mem_A[3] ));
 sg13g2_dfrbp_1 _15203_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net552),
    .D(_00650_),
    .Q_N(_06661_),
    .Q(\mem_A[4] ));
 sg13g2_dfrbp_1 _15204_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net550),
    .D(_00651_),
    .Q_N(_06660_),
    .Q(\mem_A[5] ));
 sg13g2_dfrbp_1 _15205_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net548),
    .D(net5202),
    .Q_N(_06659_),
    .Q(\mem_A[6] ));
 sg13g2_dfrbp_1 _15206_ (.CLK(clknet_leaf_71_clk),
    .RESET_B(net546),
    .D(net5099),
    .Q_N(_06658_),
    .Q(\mem_A[7] ));
 sg13g2_dfrbp_1 _15207_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net544),
    .D(_00654_),
    .Q_N(_06657_),
    .Q(\mem.mem[82][0] ));
 sg13g2_dfrbp_1 _15208_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net543),
    .D(_00655_),
    .Q_N(_06656_),
    .Q(\mem.mem[82][1] ));
 sg13g2_dfrbp_1 _15209_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net542),
    .D(_00656_),
    .Q_N(_06655_),
    .Q(\mem.mem[82][2] ));
 sg13g2_dfrbp_1 _15210_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net541),
    .D(_00657_),
    .Q_N(_06654_),
    .Q(\mem.mem[82][3] ));
 sg13g2_dfrbp_1 _15211_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net540),
    .D(_00658_),
    .Q_N(_06653_),
    .Q(\mem.mem[82][4] ));
 sg13g2_dfrbp_1 _15212_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net539),
    .D(_00659_),
    .Q_N(_06652_),
    .Q(\mem.mem[82][5] ));
 sg13g2_dfrbp_1 _15213_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net538),
    .D(_00660_),
    .Q_N(_06651_),
    .Q(\mem.mem[82][6] ));
 sg13g2_dfrbp_1 _15214_ (.CLK(clknet_leaf_53_clk),
    .RESET_B(net537),
    .D(_00661_),
    .Q_N(_06650_),
    .Q(\mem.mem[82][7] ));
 sg13g2_dfrbp_1 _15215_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net536),
    .D(_00662_),
    .Q_N(_06649_),
    .Q(\mem.mem[81][0] ));
 sg13g2_dfrbp_1 _15216_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net535),
    .D(_00663_),
    .Q_N(_06648_),
    .Q(\mem.mem[81][1] ));
 sg13g2_dfrbp_1 _15217_ (.CLK(clknet_leaf_63_clk),
    .RESET_B(net534),
    .D(_00664_),
    .Q_N(_06647_),
    .Q(\mem.mem[81][2] ));
 sg13g2_dfrbp_1 _15218_ (.CLK(clknet_leaf_60_clk),
    .RESET_B(net533),
    .D(_00665_),
    .Q_N(_06646_),
    .Q(\mem.mem[81][3] ));
 sg13g2_dfrbp_1 _15219_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net532),
    .D(_00666_),
    .Q_N(_06645_),
    .Q(\mem.mem[81][4] ));
 sg13g2_dfrbp_1 _15220_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net531),
    .D(_00667_),
    .Q_N(_06644_),
    .Q(\mem.mem[81][5] ));
 sg13g2_dfrbp_1 _15221_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net530),
    .D(_00668_),
    .Q_N(_06643_),
    .Q(\mem.mem[81][6] ));
 sg13g2_dfrbp_1 _15222_ (.CLK(clknet_leaf_61_clk),
    .RESET_B(net529),
    .D(_00669_),
    .Q_N(_06642_),
    .Q(\mem.mem[81][7] ));
 sg13g2_dfrbp_1 _15223_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net528),
    .D(_00670_),
    .Q_N(_06641_),
    .Q(\mem.mem[33][0] ));
 sg13g2_dfrbp_1 _15224_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net527),
    .D(_00671_),
    .Q_N(_06640_),
    .Q(\mem.mem[33][1] ));
 sg13g2_dfrbp_1 _15225_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net526),
    .D(_00672_),
    .Q_N(_06639_),
    .Q(\mem.mem[33][2] ));
 sg13g2_dfrbp_1 _15226_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net525),
    .D(_00673_),
    .Q_N(_06638_),
    .Q(\mem.mem[33][3] ));
 sg13g2_dfrbp_1 _15227_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net524),
    .D(_00674_),
    .Q_N(_06637_),
    .Q(\mem.mem[33][4] ));
 sg13g2_dfrbp_1 _15228_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net523),
    .D(_00675_),
    .Q_N(_06636_),
    .Q(\mem.mem[33][5] ));
 sg13g2_dfrbp_1 _15229_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net522),
    .D(_00676_),
    .Q_N(_06635_),
    .Q(\mem.mem[33][6] ));
 sg13g2_dfrbp_1 _15230_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net521),
    .D(_00677_),
    .Q_N(_06634_),
    .Q(\mem.mem[33][7] ));
 sg13g2_dfrbp_1 _15231_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net520),
    .D(_00678_),
    .Q_N(_06633_),
    .Q(\mem.mem[32][0] ));
 sg13g2_dfrbp_1 _15232_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net519),
    .D(_00679_),
    .Q_N(_06632_),
    .Q(\mem.mem[32][1] ));
 sg13g2_dfrbp_1 _15233_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net518),
    .D(_00680_),
    .Q_N(_06631_),
    .Q(\mem.mem[32][2] ));
 sg13g2_dfrbp_1 _15234_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net517),
    .D(_00681_),
    .Q_N(_06630_),
    .Q(\mem.mem[32][3] ));
 sg13g2_dfrbp_1 _15235_ (.CLK(clknet_leaf_171_clk),
    .RESET_B(net516),
    .D(_00682_),
    .Q_N(_06629_),
    .Q(\mem.mem[32][4] ));
 sg13g2_dfrbp_1 _15236_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net515),
    .D(_00683_),
    .Q_N(_06628_),
    .Q(\mem.mem[32][5] ));
 sg13g2_dfrbp_1 _15237_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net514),
    .D(_00684_),
    .Q_N(_06627_),
    .Q(\mem.mem[32][6] ));
 sg13g2_dfrbp_1 _15238_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net513),
    .D(_00685_),
    .Q_N(_06626_),
    .Q(\mem.mem[32][7] ));
 sg13g2_dfrbp_1 _15239_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net512),
    .D(_00686_),
    .Q_N(_06625_),
    .Q(\mem.mem[31][0] ));
 sg13g2_dfrbp_1 _15240_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net511),
    .D(_00687_),
    .Q_N(_06624_),
    .Q(\mem.mem[31][1] ));
 sg13g2_dfrbp_1 _15241_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net510),
    .D(_00688_),
    .Q_N(_06623_),
    .Q(\mem.mem[31][2] ));
 sg13g2_dfrbp_1 _15242_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net509),
    .D(_00689_),
    .Q_N(_06622_),
    .Q(\mem.mem[31][3] ));
 sg13g2_dfrbp_1 _15243_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net508),
    .D(_00690_),
    .Q_N(_06621_),
    .Q(\mem.mem[31][4] ));
 sg13g2_dfrbp_1 _15244_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net507),
    .D(_00691_),
    .Q_N(_06620_),
    .Q(\mem.mem[31][5] ));
 sg13g2_dfrbp_1 _15245_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net506),
    .D(_00692_),
    .Q_N(_06619_),
    .Q(\mem.mem[31][6] ));
 sg13g2_dfrbp_1 _15246_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net505),
    .D(_00693_),
    .Q_N(_06618_),
    .Q(\mem.mem[31][7] ));
 sg13g2_dfrbp_1 _15247_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net504),
    .D(_00694_),
    .Q_N(_06617_),
    .Q(\mem.mem[30][0] ));
 sg13g2_dfrbp_1 _15248_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net503),
    .D(_00695_),
    .Q_N(_06616_),
    .Q(\mem.mem[30][1] ));
 sg13g2_dfrbp_1 _15249_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net502),
    .D(_00696_),
    .Q_N(_06615_),
    .Q(\mem.mem[30][2] ));
 sg13g2_dfrbp_1 _15250_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net501),
    .D(_00697_),
    .Q_N(_06614_),
    .Q(\mem.mem[30][3] ));
 sg13g2_dfrbp_1 _15251_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net500),
    .D(_00698_),
    .Q_N(_06613_),
    .Q(\mem.mem[30][4] ));
 sg13g2_dfrbp_1 _15252_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net499),
    .D(_00699_),
    .Q_N(_06612_),
    .Q(\mem.mem[30][5] ));
 sg13g2_dfrbp_1 _15253_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net498),
    .D(_00700_),
    .Q_N(_06611_),
    .Q(\mem.mem[30][6] ));
 sg13g2_dfrbp_1 _15254_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net497),
    .D(_00701_),
    .Q_N(_06610_),
    .Q(\mem.mem[30][7] ));
 sg13g2_dfrbp_1 _15255_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net496),
    .D(_00702_),
    .Q_N(_06609_),
    .Q(\mem.mem[2][0] ));
 sg13g2_dfrbp_1 _15256_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net495),
    .D(_00703_),
    .Q_N(_06608_),
    .Q(\mem.mem[2][1] ));
 sg13g2_dfrbp_1 _15257_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net494),
    .D(_00704_),
    .Q_N(_06607_),
    .Q(\mem.mem[2][2] ));
 sg13g2_dfrbp_1 _15258_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net493),
    .D(_00705_),
    .Q_N(_06606_),
    .Q(\mem.mem[2][3] ));
 sg13g2_dfrbp_1 _15259_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net492),
    .D(_00706_),
    .Q_N(_06605_),
    .Q(\mem.mem[2][4] ));
 sg13g2_dfrbp_1 _15260_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net491),
    .D(_00707_),
    .Q_N(_06604_),
    .Q(\mem.mem[2][5] ));
 sg13g2_dfrbp_1 _15261_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net490),
    .D(_00708_),
    .Q_N(_06603_),
    .Q(\mem.mem[2][6] ));
 sg13g2_dfrbp_1 _15262_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net489),
    .D(_00709_),
    .Q_N(_06602_),
    .Q(\mem.mem[2][7] ));
 sg13g2_dfrbp_1 _15263_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net488),
    .D(_00710_),
    .Q_N(_06601_),
    .Q(\mem.mem[28][0] ));
 sg13g2_dfrbp_1 _15264_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net487),
    .D(_00711_),
    .Q_N(_06600_),
    .Q(\mem.mem[28][1] ));
 sg13g2_dfrbp_1 _15265_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net486),
    .D(_00712_),
    .Q_N(_06599_),
    .Q(\mem.mem[28][2] ));
 sg13g2_dfrbp_1 _15266_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net485),
    .D(_00713_),
    .Q_N(_06598_),
    .Q(\mem.mem[28][3] ));
 sg13g2_dfrbp_1 _15267_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net484),
    .D(_00714_),
    .Q_N(_06597_),
    .Q(\mem.mem[28][4] ));
 sg13g2_dfrbp_1 _15268_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net483),
    .D(_00715_),
    .Q_N(_06596_),
    .Q(\mem.mem[28][5] ));
 sg13g2_dfrbp_1 _15269_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net482),
    .D(_00716_),
    .Q_N(_06595_),
    .Q(\mem.mem[28][6] ));
 sg13g2_dfrbp_1 _15270_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net481),
    .D(_00717_),
    .Q_N(_06594_),
    .Q(\mem.mem[28][7] ));
 sg13g2_dfrbp_1 _15271_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net480),
    .D(_00718_),
    .Q_N(_06593_),
    .Q(\mem.mem[27][0] ));
 sg13g2_dfrbp_1 _15272_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net479),
    .D(_00719_),
    .Q_N(_06592_),
    .Q(\mem.mem[27][1] ));
 sg13g2_dfrbp_1 _15273_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net478),
    .D(_00720_),
    .Q_N(_06591_),
    .Q(\mem.mem[27][2] ));
 sg13g2_dfrbp_1 _15274_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net477),
    .D(_00721_),
    .Q_N(_06590_),
    .Q(\mem.mem[27][3] ));
 sg13g2_dfrbp_1 _15275_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net476),
    .D(_00722_),
    .Q_N(_06589_),
    .Q(\mem.mem[27][4] ));
 sg13g2_dfrbp_1 _15276_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net475),
    .D(_00723_),
    .Q_N(_06588_),
    .Q(\mem.mem[27][5] ));
 sg13g2_dfrbp_1 _15277_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net474),
    .D(_00724_),
    .Q_N(_06587_),
    .Q(\mem.mem[27][6] ));
 sg13g2_dfrbp_1 _15278_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net473),
    .D(_00725_),
    .Q_N(_06586_),
    .Q(\mem.mem[27][7] ));
 sg13g2_dfrbp_1 _15279_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net472),
    .D(_00726_),
    .Q_N(_06585_),
    .Q(\mem.mem[26][0] ));
 sg13g2_dfrbp_1 _15280_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net471),
    .D(_00727_),
    .Q_N(_06584_),
    .Q(\mem.mem[26][1] ));
 sg13g2_dfrbp_1 _15281_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net470),
    .D(_00728_),
    .Q_N(_06583_),
    .Q(\mem.mem[26][2] ));
 sg13g2_dfrbp_1 _15282_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net469),
    .D(_00729_),
    .Q_N(_06582_),
    .Q(\mem.mem[26][3] ));
 sg13g2_dfrbp_1 _15283_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net468),
    .D(_00730_),
    .Q_N(_06581_),
    .Q(\mem.mem[26][4] ));
 sg13g2_dfrbp_1 _15284_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net467),
    .D(_00731_),
    .Q_N(_06580_),
    .Q(\mem.mem[26][5] ));
 sg13g2_dfrbp_1 _15285_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net466),
    .D(_00732_),
    .Q_N(_06579_),
    .Q(\mem.mem[26][6] ));
 sg13g2_dfrbp_1 _15286_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net465),
    .D(_00733_),
    .Q_N(_06578_),
    .Q(\mem.mem[26][7] ));
 sg13g2_dfrbp_1 _15287_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net464),
    .D(_00734_),
    .Q_N(_06577_),
    .Q(\mem.mem[25][0] ));
 sg13g2_dfrbp_1 _15288_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net463),
    .D(_00735_),
    .Q_N(_06576_),
    .Q(\mem.mem[25][1] ));
 sg13g2_dfrbp_1 _15289_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net462),
    .D(_00736_),
    .Q_N(_06575_),
    .Q(\mem.mem[25][2] ));
 sg13g2_dfrbp_1 _15290_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net461),
    .D(_00737_),
    .Q_N(_06574_),
    .Q(\mem.mem[25][3] ));
 sg13g2_dfrbp_1 _15291_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net460),
    .D(_00738_),
    .Q_N(_06573_),
    .Q(\mem.mem[25][4] ));
 sg13g2_dfrbp_1 _15292_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net459),
    .D(_00739_),
    .Q_N(_06572_),
    .Q(\mem.mem[25][5] ));
 sg13g2_dfrbp_1 _15293_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net458),
    .D(_00740_),
    .Q_N(_06571_),
    .Q(\mem.mem[25][6] ));
 sg13g2_dfrbp_1 _15294_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net457),
    .D(_00741_),
    .Q_N(_06570_),
    .Q(\mem.mem[25][7] ));
 sg13g2_dfrbp_1 _15295_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net456),
    .D(_00742_),
    .Q_N(_06569_),
    .Q(\mem.mem[252][0] ));
 sg13g2_dfrbp_1 _15296_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net455),
    .D(_00743_),
    .Q_N(_06568_),
    .Q(\mem.mem[252][1] ));
 sg13g2_dfrbp_1 _15297_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net454),
    .D(_00744_),
    .Q_N(_06567_),
    .Q(\mem.mem[252][2] ));
 sg13g2_dfrbp_1 _15298_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net453),
    .D(_00745_),
    .Q_N(_06566_),
    .Q(\mem.mem[252][3] ));
 sg13g2_dfrbp_1 _15299_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net452),
    .D(_00746_),
    .Q_N(_06565_),
    .Q(\mem.mem[252][4] ));
 sg13g2_dfrbp_1 _15300_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net451),
    .D(_00747_),
    .Q_N(_06564_),
    .Q(\mem.mem[252][5] ));
 sg13g2_dfrbp_1 _15301_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net450),
    .D(_00748_),
    .Q_N(_06563_),
    .Q(\mem.mem[252][6] ));
 sg13g2_dfrbp_1 _15302_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net449),
    .D(_00749_),
    .Q_N(_06562_),
    .Q(\mem.mem[252][7] ));
 sg13g2_dfrbp_1 _15303_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net448),
    .D(_00750_),
    .Q_N(_06561_),
    .Q(\mem.mem[249][0] ));
 sg13g2_dfrbp_1 _15304_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net447),
    .D(_00751_),
    .Q_N(_06560_),
    .Q(\mem.mem[249][1] ));
 sg13g2_dfrbp_1 _15305_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net446),
    .D(_00752_),
    .Q_N(_06559_),
    .Q(\mem.mem[249][2] ));
 sg13g2_dfrbp_1 _15306_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net445),
    .D(_00753_),
    .Q_N(_06558_),
    .Q(\mem.mem[249][3] ));
 sg13g2_dfrbp_1 _15307_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net444),
    .D(_00754_),
    .Q_N(_06557_),
    .Q(\mem.mem[249][4] ));
 sg13g2_dfrbp_1 _15308_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net443),
    .D(_00755_),
    .Q_N(_06556_),
    .Q(\mem.mem[249][5] ));
 sg13g2_dfrbp_1 _15309_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net442),
    .D(_00756_),
    .Q_N(_06555_),
    .Q(\mem.mem[249][6] ));
 sg13g2_dfrbp_1 _15310_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net441),
    .D(_00757_),
    .Q_N(_06554_),
    .Q(\mem.mem[249][7] ));
 sg13g2_dfrbp_1 _15311_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net440),
    .D(_00758_),
    .Q_N(_06553_),
    .Q(\mem.mem[49][0] ));
 sg13g2_dfrbp_1 _15312_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net439),
    .D(_00759_),
    .Q_N(_06552_),
    .Q(\mem.mem[49][1] ));
 sg13g2_dfrbp_1 _15313_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net438),
    .D(_00760_),
    .Q_N(_06551_),
    .Q(\mem.mem[49][2] ));
 sg13g2_dfrbp_1 _15314_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net437),
    .D(_00761_),
    .Q_N(_06550_),
    .Q(\mem.mem[49][3] ));
 sg13g2_dfrbp_1 _15315_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net436),
    .D(_00762_),
    .Q_N(_06549_),
    .Q(\mem.mem[49][4] ));
 sg13g2_dfrbp_1 _15316_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net435),
    .D(_00763_),
    .Q_N(_06548_),
    .Q(\mem.mem[49][5] ));
 sg13g2_dfrbp_1 _15317_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net434),
    .D(_00764_),
    .Q_N(_06547_),
    .Q(\mem.mem[49][6] ));
 sg13g2_dfrbp_1 _15318_ (.CLK(clknet_leaf_150_clk),
    .RESET_B(net433),
    .D(_00765_),
    .Q_N(_06546_),
    .Q(\mem.mem[49][7] ));
 sg13g2_dfrbp_1 _15319_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net432),
    .D(_00766_),
    .Q_N(_06545_),
    .Q(\mem.mem[39][0] ));
 sg13g2_dfrbp_1 _15320_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net431),
    .D(_00767_),
    .Q_N(_06544_),
    .Q(\mem.mem[39][1] ));
 sg13g2_dfrbp_1 _15321_ (.CLK(clknet_leaf_175_clk),
    .RESET_B(net430),
    .D(_00768_),
    .Q_N(_06543_),
    .Q(\mem.mem[39][2] ));
 sg13g2_dfrbp_1 _15322_ (.CLK(clknet_leaf_183_clk),
    .RESET_B(net429),
    .D(_00769_),
    .Q_N(_06542_),
    .Q(\mem.mem[39][3] ));
 sg13g2_dfrbp_1 _15323_ (.CLK(clknet_leaf_178_clk),
    .RESET_B(net428),
    .D(_00770_),
    .Q_N(_06541_),
    .Q(\mem.mem[39][4] ));
 sg13g2_dfrbp_1 _15324_ (.CLK(clknet_leaf_180_clk),
    .RESET_B(net427),
    .D(_00771_),
    .Q_N(_06540_),
    .Q(\mem.mem[39][5] ));
 sg13g2_dfrbp_1 _15325_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net426),
    .D(_00772_),
    .Q_N(_06539_),
    .Q(\mem.mem[39][6] ));
 sg13g2_dfrbp_1 _15326_ (.CLK(clknet_leaf_179_clk),
    .RESET_B(net425),
    .D(_00773_),
    .Q_N(_06538_),
    .Q(\mem.mem[39][7] ));
 sg13g2_dfrbp_1 _15327_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net424),
    .D(_00774_),
    .Q_N(_06537_),
    .Q(\mem.mem[239][0] ));
 sg13g2_dfrbp_1 _15328_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net423),
    .D(_00775_),
    .Q_N(_06536_),
    .Q(\mem.mem[239][1] ));
 sg13g2_dfrbp_1 _15329_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net422),
    .D(_00776_),
    .Q_N(_06535_),
    .Q(\mem.mem[239][2] ));
 sg13g2_dfrbp_1 _15330_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net421),
    .D(_00777_),
    .Q_N(_06534_),
    .Q(\mem.mem[239][3] ));
 sg13g2_dfrbp_1 _15331_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net420),
    .D(_00778_),
    .Q_N(_06533_),
    .Q(\mem.mem[239][4] ));
 sg13g2_dfrbp_1 _15332_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net419),
    .D(_00779_),
    .Q_N(_06532_),
    .Q(\mem.mem[239][5] ));
 sg13g2_dfrbp_1 _15333_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net418),
    .D(_00780_),
    .Q_N(_06531_),
    .Q(\mem.mem[239][6] ));
 sg13g2_dfrbp_1 _15334_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net417),
    .D(_00781_),
    .Q_N(_06530_),
    .Q(\mem.mem[239][7] ));
 sg13g2_dfrbp_1 _15335_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net416),
    .D(_00782_),
    .Q_N(_06529_),
    .Q(\mem.mem[229][0] ));
 sg13g2_dfrbp_1 _15336_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net415),
    .D(_00783_),
    .Q_N(_06528_),
    .Q(\mem.mem[229][1] ));
 sg13g2_dfrbp_1 _15337_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net414),
    .D(_00784_),
    .Q_N(_06527_),
    .Q(\mem.mem[229][2] ));
 sg13g2_dfrbp_1 _15338_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net413),
    .D(_00785_),
    .Q_N(_06526_),
    .Q(\mem.mem[229][3] ));
 sg13g2_dfrbp_1 _15339_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net412),
    .D(_00786_),
    .Q_N(_06525_),
    .Q(\mem.mem[229][4] ));
 sg13g2_dfrbp_1 _15340_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net411),
    .D(_00787_),
    .Q_N(_06524_),
    .Q(\mem.mem[229][5] ));
 sg13g2_dfrbp_1 _15341_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net410),
    .D(_00788_),
    .Q_N(_06523_),
    .Q(\mem.mem[229][6] ));
 sg13g2_dfrbp_1 _15342_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net409),
    .D(_00789_),
    .Q_N(_06522_),
    .Q(\mem.mem[229][7] ));
 sg13g2_dfrbp_1 _15343_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net408),
    .D(_00790_),
    .Q_N(_06521_),
    .Q(\mem.mem[29][0] ));
 sg13g2_dfrbp_1 _15344_ (.CLK(clknet_leaf_186_clk),
    .RESET_B(net407),
    .D(_00791_),
    .Q_N(_06520_),
    .Q(\mem.mem[29][1] ));
 sg13g2_dfrbp_1 _15345_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net406),
    .D(_00792_),
    .Q_N(_06519_),
    .Q(\mem.mem[29][2] ));
 sg13g2_dfrbp_1 _15346_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net405),
    .D(_00793_),
    .Q_N(_06518_),
    .Q(\mem.mem[29][3] ));
 sg13g2_dfrbp_1 _15347_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net404),
    .D(_00794_),
    .Q_N(_06517_),
    .Q(\mem.mem[29][4] ));
 sg13g2_dfrbp_1 _15348_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net403),
    .D(_00795_),
    .Q_N(_06516_),
    .Q(\mem.mem[29][5] ));
 sg13g2_dfrbp_1 _15349_ (.CLK(clknet_leaf_184_clk),
    .RESET_B(net402),
    .D(_00796_),
    .Q_N(_06515_),
    .Q(\mem.mem[29][6] ));
 sg13g2_dfrbp_1 _15350_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net401),
    .D(_00797_),
    .Q_N(_06514_),
    .Q(\mem.mem[29][7] ));
 sg13g2_dfrbp_1 _15351_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net400),
    .D(_00798_),
    .Q_N(_06513_),
    .Q(\mem.mem[219][0] ));
 sg13g2_dfrbp_1 _15352_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net399),
    .D(_00799_),
    .Q_N(_06512_),
    .Q(\mem.mem[219][1] ));
 sg13g2_dfrbp_1 _15353_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net398),
    .D(_00800_),
    .Q_N(_06511_),
    .Q(\mem.mem[219][2] ));
 sg13g2_dfrbp_1 _15354_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net397),
    .D(_00801_),
    .Q_N(_06510_),
    .Q(\mem.mem[219][3] ));
 sg13g2_dfrbp_1 _15355_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net396),
    .D(_00802_),
    .Q_N(_06509_),
    .Q(\mem.mem[219][4] ));
 sg13g2_dfrbp_1 _15356_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net395),
    .D(_00803_),
    .Q_N(_06508_),
    .Q(\mem.mem[219][5] ));
 sg13g2_dfrbp_1 _15357_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net394),
    .D(_00804_),
    .Q_N(_06507_),
    .Q(\mem.mem[219][6] ));
 sg13g2_dfrbp_1 _15358_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net393),
    .D(_00805_),
    .Q_N(_06506_),
    .Q(\mem.mem[219][7] ));
 sg13g2_dfrbp_1 _15359_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net392),
    .D(_00806_),
    .Q_N(_06505_),
    .Q(\mem.mem[97][0] ));
 sg13g2_dfrbp_1 _15360_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net391),
    .D(_00807_),
    .Q_N(_06504_),
    .Q(\mem.mem[97][1] ));
 sg13g2_dfrbp_1 _15361_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net390),
    .D(_00808_),
    .Q_N(_06503_),
    .Q(\mem.mem[97][2] ));
 sg13g2_dfrbp_1 _15362_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net389),
    .D(_00809_),
    .Q_N(_06502_),
    .Q(\mem.mem[97][3] ));
 sg13g2_dfrbp_1 _15363_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net388),
    .D(_00810_),
    .Q_N(_06501_),
    .Q(\mem.mem[97][4] ));
 sg13g2_dfrbp_1 _15364_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net387),
    .D(_00811_),
    .Q_N(_06500_),
    .Q(\mem.mem[97][5] ));
 sg13g2_dfrbp_1 _15365_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net386),
    .D(_00812_),
    .Q_N(_06499_),
    .Q(\mem.mem[97][6] ));
 sg13g2_dfrbp_1 _15366_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net385),
    .D(_00813_),
    .Q_N(_06498_),
    .Q(\mem.mem[97][7] ));
 sg13g2_dfrbp_1 _15367_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net384),
    .D(_00814_),
    .Q_N(_06497_),
    .Q(\mem.mem[96][0] ));
 sg13g2_dfrbp_1 _15368_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net383),
    .D(_00815_),
    .Q_N(_06496_),
    .Q(\mem.mem[96][1] ));
 sg13g2_dfrbp_1 _15369_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net382),
    .D(_00816_),
    .Q_N(_06495_),
    .Q(\mem.mem[96][2] ));
 sg13g2_dfrbp_1 _15370_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net381),
    .D(_00817_),
    .Q_N(_06494_),
    .Q(\mem.mem[96][3] ));
 sg13g2_dfrbp_1 _15371_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net380),
    .D(_00818_),
    .Q_N(_06493_),
    .Q(\mem.mem[96][4] ));
 sg13g2_dfrbp_1 _15372_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net379),
    .D(_00819_),
    .Q_N(_06492_),
    .Q(\mem.mem[96][5] ));
 sg13g2_dfrbp_1 _15373_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net378),
    .D(_00820_),
    .Q_N(_06491_),
    .Q(\mem.mem[96][6] ));
 sg13g2_dfrbp_1 _15374_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net377),
    .D(_00821_),
    .Q_N(_06490_),
    .Q(\mem.mem[96][7] ));
 sg13g2_dfrbp_1 _15375_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net376),
    .D(_00822_),
    .Q_N(_06489_),
    .Q(\mem.mem[95][0] ));
 sg13g2_dfrbp_1 _15376_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net375),
    .D(_00823_),
    .Q_N(_06488_),
    .Q(\mem.mem[95][1] ));
 sg13g2_dfrbp_1 _15377_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net374),
    .D(_00824_),
    .Q_N(_06487_),
    .Q(\mem.mem[95][2] ));
 sg13g2_dfrbp_1 _15378_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net373),
    .D(_00825_),
    .Q_N(_06486_),
    .Q(\mem.mem[95][3] ));
 sg13g2_dfrbp_1 _15379_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net372),
    .D(_00826_),
    .Q_N(_06485_),
    .Q(\mem.mem[95][4] ));
 sg13g2_dfrbp_1 _15380_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net371),
    .D(_00827_),
    .Q_N(_06484_),
    .Q(\mem.mem[95][5] ));
 sg13g2_dfrbp_1 _15381_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net370),
    .D(_00828_),
    .Q_N(_06483_),
    .Q(\mem.mem[95][6] ));
 sg13g2_dfrbp_1 _15382_ (.CLK(clknet_leaf_67_clk),
    .RESET_B(net369),
    .D(_00829_),
    .Q_N(_06482_),
    .Q(\mem.mem[95][7] ));
 sg13g2_dfrbp_1 _15383_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net368),
    .D(_00830_),
    .Q_N(_06481_),
    .Q(\mem.mem[50][0] ));
 sg13g2_dfrbp_1 _15384_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net367),
    .D(_00831_),
    .Q_N(_06480_),
    .Q(\mem.mem[50][1] ));
 sg13g2_dfrbp_1 _15385_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net366),
    .D(_00832_),
    .Q_N(_06479_),
    .Q(\mem.mem[50][2] ));
 sg13g2_dfrbp_1 _15386_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net365),
    .D(_00833_),
    .Q_N(_06478_),
    .Q(\mem.mem[50][3] ));
 sg13g2_dfrbp_1 _15387_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net364),
    .D(_00834_),
    .Q_N(_06477_),
    .Q(\mem.mem[50][4] ));
 sg13g2_dfrbp_1 _15388_ (.CLK(clknet_leaf_151_clk),
    .RESET_B(net363),
    .D(_00835_),
    .Q_N(_06476_),
    .Q(\mem.mem[50][5] ));
 sg13g2_dfrbp_1 _15389_ (.CLK(clknet_leaf_152_clk),
    .RESET_B(net362),
    .D(_00836_),
    .Q_N(_06475_),
    .Q(\mem.mem[50][6] ));
 sg13g2_dfrbp_1 _15390_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net361),
    .D(_00837_),
    .Q_N(_06474_),
    .Q(\mem.mem[50][7] ));
 sg13g2_dfrbp_1 _15391_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net360),
    .D(net2131),
    .Q_N(_06473_),
    .Q(\mem.out_strobe ));
 sg13g2_dfrbp_1 _15392_ (.CLK(clknet_leaf_73_clk),
    .RESET_B(net358),
    .D(net2204),
    .Q_N(_06472_),
    .Q(\mem.uo_out[0] ));
 sg13g2_dfrbp_1 _15393_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net356),
    .D(_00840_),
    .Q_N(_06471_),
    .Q(\mem.uo_out[1] ));
 sg13g2_dfrbp_1 _15394_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net354),
    .D(_00841_),
    .Q_N(_06470_),
    .Q(\mem.uo_out[2] ));
 sg13g2_dfrbp_1 _15395_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net352),
    .D(_00842_),
    .Q_N(_06469_),
    .Q(\mem.uo_out[3] ));
 sg13g2_dfrbp_1 _15396_ (.CLK(clknet_leaf_59_clk),
    .RESET_B(net350),
    .D(_00843_),
    .Q_N(_06468_),
    .Q(\mem.uo_out[4] ));
 sg13g2_dfrbp_1 _15397_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net348),
    .D(_00844_),
    .Q_N(_06467_),
    .Q(\mem.uo_out[5] ));
 sg13g2_dfrbp_1 _15398_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net346),
    .D(_00845_),
    .Q_N(_06466_),
    .Q(\mem.uo_out[6] ));
 sg13g2_dfrbp_1 _15399_ (.CLK(clknet_leaf_70_clk),
    .RESET_B(net344),
    .D(_00846_),
    .Q_N(_06465_),
    .Q(\mem.uo_out[7] ));
 sg13g2_dfrbp_1 _15400_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net342),
    .D(_00847_),
    .Q_N(_06464_),
    .Q(\mem.mem[109][0] ));
 sg13g2_dfrbp_1 _15401_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net341),
    .D(_00848_),
    .Q_N(_06463_),
    .Q(\mem.mem[109][1] ));
 sg13g2_dfrbp_1 _15402_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net340),
    .D(_00849_),
    .Q_N(_06462_),
    .Q(\mem.mem[109][2] ));
 sg13g2_dfrbp_1 _15403_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net339),
    .D(_00850_),
    .Q_N(_06461_),
    .Q(\mem.mem[109][3] ));
 sg13g2_dfrbp_1 _15404_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net338),
    .D(_00851_),
    .Q_N(_06460_),
    .Q(\mem.mem[109][4] ));
 sg13g2_dfrbp_1 _15405_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net337),
    .D(_00852_),
    .Q_N(_06459_),
    .Q(\mem.mem[109][5] ));
 sg13g2_dfrbp_1 _15406_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net336),
    .D(_00853_),
    .Q_N(_06458_),
    .Q(\mem.mem[109][6] ));
 sg13g2_dfrbp_1 _15407_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net335),
    .D(_00854_),
    .Q_N(_06457_),
    .Q(\mem.mem[109][7] ));
 sg13g2_dfrbp_1 _15408_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net334),
    .D(_00855_),
    .Q_N(_06456_),
    .Q(\mem.mem[99][0] ));
 sg13g2_dfrbp_1 _15409_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net333),
    .D(_00856_),
    .Q_N(_06455_),
    .Q(\mem.mem[99][1] ));
 sg13g2_dfrbp_1 _15410_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net332),
    .D(_00857_),
    .Q_N(_06454_),
    .Q(\mem.mem[99][2] ));
 sg13g2_dfrbp_1 _15411_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net331),
    .D(_00858_),
    .Q_N(_06453_),
    .Q(\mem.mem[99][3] ));
 sg13g2_dfrbp_1 _15412_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net330),
    .D(_00859_),
    .Q_N(_06452_),
    .Q(\mem.mem[99][4] ));
 sg13g2_dfrbp_1 _15413_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net329),
    .D(_00860_),
    .Q_N(_06451_),
    .Q(\mem.mem[99][5] ));
 sg13g2_dfrbp_1 _15414_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net328),
    .D(_00861_),
    .Q_N(_06450_),
    .Q(\mem.mem[99][6] ));
 sg13g2_dfrbp_1 _15415_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net327),
    .D(_00862_),
    .Q_N(_06449_),
    .Q(\mem.mem[99][7] ));
 sg13g2_dfrbp_1 _15416_ (.CLK(clknet_leaf_72_clk),
    .RESET_B(net326),
    .D(_00863_),
    .Q_N(_06448_),
    .Q(\mem.mem[89][0] ));
 sg13g2_dfrbp_1 _15417_ (.CLK(clknet_leaf_62_clk),
    .RESET_B(net325),
    .D(_00864_),
    .Q_N(_06447_),
    .Q(\mem.mem[89][1] ));
 sg13g2_dfrbp_1 _15418_ (.CLK(clknet_leaf_64_clk),
    .RESET_B(net324),
    .D(_00865_),
    .Q_N(_06446_),
    .Q(\mem.mem[89][2] ));
 sg13g2_dfrbp_1 _15419_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net323),
    .D(_00866_),
    .Q_N(_06445_),
    .Q(\mem.mem[89][3] ));
 sg13g2_dfrbp_1 _15420_ (.CLK(clknet_leaf_66_clk),
    .RESET_B(net322),
    .D(_00867_),
    .Q_N(_06444_),
    .Q(\mem.mem[89][4] ));
 sg13g2_dfrbp_1 _15421_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net321),
    .D(_00868_),
    .Q_N(_06443_),
    .Q(\mem.mem[89][5] ));
 sg13g2_dfrbp_1 _15422_ (.CLK(clknet_leaf_68_clk),
    .RESET_B(net320),
    .D(_00869_),
    .Q_N(_06442_),
    .Q(\mem.mem[89][6] ));
 sg13g2_dfrbp_1 _15423_ (.CLK(clknet_leaf_65_clk),
    .RESET_B(net319),
    .D(_00870_),
    .Q_N(_06441_),
    .Q(\mem.mem[89][7] ));
 sg13g2_dfrbp_1 _15424_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net318),
    .D(_00871_),
    .Q_N(_06440_),
    .Q(\mem.mem[139][0] ));
 sg13g2_dfrbp_1 _15425_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net317),
    .D(_00872_),
    .Q_N(_06439_),
    .Q(\mem.mem[139][1] ));
 sg13g2_dfrbp_1 _15426_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net316),
    .D(_00873_),
    .Q_N(_06438_),
    .Q(\mem.mem[139][2] ));
 sg13g2_dfrbp_1 _15427_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net315),
    .D(_00874_),
    .Q_N(_06437_),
    .Q(\mem.mem[139][3] ));
 sg13g2_dfrbp_1 _15428_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net314),
    .D(_00875_),
    .Q_N(_06436_),
    .Q(\mem.mem[139][4] ));
 sg13g2_dfrbp_1 _15429_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net313),
    .D(_00876_),
    .Q_N(_06435_),
    .Q(\mem.mem[139][5] ));
 sg13g2_dfrbp_1 _15430_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net312),
    .D(_00877_),
    .Q_N(_06434_),
    .Q(\mem.mem[139][6] ));
 sg13g2_dfrbp_1 _15431_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net311),
    .D(_00878_),
    .Q_N(_06433_),
    .Q(\mem.mem[139][7] ));
 sg13g2_dfrbp_1 _15432_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net310),
    .D(_00879_),
    .Q_N(_06432_),
    .Q(\mem.mem[98][0] ));
 sg13g2_dfrbp_1 _15433_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net309),
    .D(_00880_),
    .Q_N(_06431_),
    .Q(\mem.mem[98][1] ));
 sg13g2_dfrbp_1 _15434_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net308),
    .D(_00881_),
    .Q_N(_06430_),
    .Q(\mem.mem[98][2] ));
 sg13g2_dfrbp_1 _15435_ (.CLK(clknet_leaf_105_clk),
    .RESET_B(net307),
    .D(_00882_),
    .Q_N(_06429_),
    .Q(\mem.mem[98][3] ));
 sg13g2_dfrbp_1 _15436_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net306),
    .D(_00883_),
    .Q_N(_06428_),
    .Q(\mem.mem[98][4] ));
 sg13g2_dfrbp_1 _15437_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net305),
    .D(_00884_),
    .Q_N(_06427_),
    .Q(\mem.mem[98][5] ));
 sg13g2_dfrbp_1 _15438_ (.CLK(clknet_leaf_99_clk),
    .RESET_B(net304),
    .D(_00885_),
    .Q_N(_06426_),
    .Q(\mem.mem[98][6] ));
 sg13g2_dfrbp_1 _15439_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net303),
    .D(_00886_),
    .Q_N(_06425_),
    .Q(\mem.mem[98][7] ));
 sg13g2_dfrbp_1 _15440_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net302),
    .D(_00887_),
    .Q_N(_06424_),
    .Q(\mem.mem[0][0] ));
 sg13g2_dfrbp_1 _15441_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net301),
    .D(_00888_),
    .Q_N(_06423_),
    .Q(\mem.mem[0][1] ));
 sg13g2_dfrbp_1 _15442_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net300),
    .D(_00889_),
    .Q_N(_06422_),
    .Q(\mem.mem[0][2] ));
 sg13g2_dfrbp_1 _15443_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net299),
    .D(_00890_),
    .Q_N(_06421_),
    .Q(\mem.mem[0][3] ));
 sg13g2_dfrbp_1 _15444_ (.CLK(clknet_leaf_206_clk),
    .RESET_B(net298),
    .D(_00891_),
    .Q_N(_06420_),
    .Q(\mem.mem[0][4] ));
 sg13g2_dfrbp_1 _15445_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net297),
    .D(_00892_),
    .Q_N(_06419_),
    .Q(\mem.mem[0][5] ));
 sg13g2_dfrbp_1 _15446_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net296),
    .D(_00893_),
    .Q_N(_06418_),
    .Q(\mem.mem[0][6] ));
 sg13g2_dfrbp_1 _15447_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net295),
    .D(_00894_),
    .Q_N(_06417_),
    .Q(\mem.mem[0][7] ));
 sg13g2_dfrbp_1 _15448_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net294),
    .D(_00895_),
    .Q_N(_06416_),
    .Q(\mem.mem[100][0] ));
 sg13g2_dfrbp_1 _15449_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net293),
    .D(_00896_),
    .Q_N(_06415_),
    .Q(\mem.mem[100][1] ));
 sg13g2_dfrbp_1 _15450_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net292),
    .D(_00897_),
    .Q_N(_06414_),
    .Q(\mem.mem[100][2] ));
 sg13g2_dfrbp_1 _15451_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net291),
    .D(_00898_),
    .Q_N(_06413_),
    .Q(\mem.mem[100][3] ));
 sg13g2_dfrbp_1 _15452_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net290),
    .D(_00899_),
    .Q_N(_06412_),
    .Q(\mem.mem[100][4] ));
 sg13g2_dfrbp_1 _15453_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net289),
    .D(_00900_),
    .Q_N(_06411_),
    .Q(\mem.mem[100][5] ));
 sg13g2_dfrbp_1 _15454_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net288),
    .D(_00901_),
    .Q_N(_06410_),
    .Q(\mem.mem[100][6] ));
 sg13g2_dfrbp_1 _15455_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net287),
    .D(_00902_),
    .Q_N(_06409_),
    .Q(\mem.mem[100][7] ));
 sg13g2_dfrbp_1 _15456_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net286),
    .D(_00903_),
    .Q_N(_06408_),
    .Q(\mem.mem[101][0] ));
 sg13g2_dfrbp_1 _15457_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net285),
    .D(_00904_),
    .Q_N(_06407_),
    .Q(\mem.mem[101][1] ));
 sg13g2_dfrbp_1 _15458_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net284),
    .D(_00905_),
    .Q_N(_06406_),
    .Q(\mem.mem[101][2] ));
 sg13g2_dfrbp_1 _15459_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net283),
    .D(_00906_),
    .Q_N(_06405_),
    .Q(\mem.mem[101][3] ));
 sg13g2_dfrbp_1 _15460_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net282),
    .D(_00907_),
    .Q_N(_06404_),
    .Q(\mem.mem[101][4] ));
 sg13g2_dfrbp_1 _15461_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net281),
    .D(_00908_),
    .Q_N(_06403_),
    .Q(\mem.mem[101][5] ));
 sg13g2_dfrbp_1 _15462_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net280),
    .D(_00909_),
    .Q_N(_06402_),
    .Q(\mem.mem[101][6] ));
 sg13g2_dfrbp_1 _15463_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net279),
    .D(_00910_),
    .Q_N(_06401_),
    .Q(\mem.mem[101][7] ));
 sg13g2_dfrbp_1 _15464_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net278),
    .D(_00911_),
    .Q_N(_06400_),
    .Q(\mem.mem[102][0] ));
 sg13g2_dfrbp_1 _15465_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net277),
    .D(_00912_),
    .Q_N(_06399_),
    .Q(\mem.mem[102][1] ));
 sg13g2_dfrbp_1 _15466_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net276),
    .D(_00913_),
    .Q_N(_06398_),
    .Q(\mem.mem[102][2] ));
 sg13g2_dfrbp_1 _15467_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net275),
    .D(_00914_),
    .Q_N(_06397_),
    .Q(\mem.mem[102][3] ));
 sg13g2_dfrbp_1 _15468_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net274),
    .D(_00915_),
    .Q_N(_06396_),
    .Q(\mem.mem[102][4] ));
 sg13g2_dfrbp_1 _15469_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net273),
    .D(_00916_),
    .Q_N(_06395_),
    .Q(\mem.mem[102][5] ));
 sg13g2_dfrbp_1 _15470_ (.CLK(clknet_leaf_102_clk),
    .RESET_B(net272),
    .D(_00917_),
    .Q_N(_06394_),
    .Q(\mem.mem[102][6] ));
 sg13g2_dfrbp_1 _15471_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net271),
    .D(_00918_),
    .Q_N(_06393_),
    .Q(\mem.mem[102][7] ));
 sg13g2_dfrbp_1 _15472_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net270),
    .D(_00919_),
    .Q_N(_06392_),
    .Q(\mem.mem[103][0] ));
 sg13g2_dfrbp_1 _15473_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net269),
    .D(_00920_),
    .Q_N(_06391_),
    .Q(\mem.mem[103][1] ));
 sg13g2_dfrbp_1 _15474_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net268),
    .D(_00921_),
    .Q_N(_06390_),
    .Q(\mem.mem[103][2] ));
 sg13g2_dfrbp_1 _15475_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net267),
    .D(_00922_),
    .Q_N(_06389_),
    .Q(\mem.mem[103][3] ));
 sg13g2_dfrbp_1 _15476_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net266),
    .D(_00923_),
    .Q_N(_06388_),
    .Q(\mem.mem[103][4] ));
 sg13g2_dfrbp_1 _15477_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net265),
    .D(_00924_),
    .Q_N(_06387_),
    .Q(\mem.mem[103][5] ));
 sg13g2_dfrbp_1 _15478_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net264),
    .D(_00925_),
    .Q_N(_06386_),
    .Q(\mem.mem[103][6] ));
 sg13g2_dfrbp_1 _15479_ (.CLK(clknet_leaf_103_clk),
    .RESET_B(net263),
    .D(_00926_),
    .Q_N(_06385_),
    .Q(\mem.mem[103][7] ));
 sg13g2_dfrbp_1 _15480_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net262),
    .D(_00927_),
    .Q_N(_06384_),
    .Q(\mem.mem[104][0] ));
 sg13g2_dfrbp_1 _15481_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net261),
    .D(_00928_),
    .Q_N(_06383_),
    .Q(\mem.mem[104][1] ));
 sg13g2_dfrbp_1 _15482_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net260),
    .D(_00929_),
    .Q_N(_06382_),
    .Q(\mem.mem[104][2] ));
 sg13g2_dfrbp_1 _15483_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net259),
    .D(_00930_),
    .Q_N(_06381_),
    .Q(\mem.mem[104][3] ));
 sg13g2_dfrbp_1 _15484_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net258),
    .D(_00931_),
    .Q_N(_06380_),
    .Q(\mem.mem[104][4] ));
 sg13g2_dfrbp_1 _15485_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net257),
    .D(_00932_),
    .Q_N(_06379_),
    .Q(\mem.mem[104][5] ));
 sg13g2_dfrbp_1 _15486_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net256),
    .D(_00933_),
    .Q_N(_06378_),
    .Q(\mem.mem[104][6] ));
 sg13g2_dfrbp_1 _15487_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net255),
    .D(_00934_),
    .Q_N(_06377_),
    .Q(\mem.mem[104][7] ));
 sg13g2_dfrbp_1 _15488_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net254),
    .D(_00935_),
    .Q_N(_06376_),
    .Q(\mem.mem[105][0] ));
 sg13g2_dfrbp_1 _15489_ (.CLK(clknet_leaf_104_clk),
    .RESET_B(net253),
    .D(_00936_),
    .Q_N(_06375_),
    .Q(\mem.mem[105][1] ));
 sg13g2_dfrbp_1 _15490_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net252),
    .D(_00937_),
    .Q_N(_06374_),
    .Q(\mem.mem[105][2] ));
 sg13g2_dfrbp_1 _15491_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net251),
    .D(_00938_),
    .Q_N(_06373_),
    .Q(\mem.mem[105][3] ));
 sg13g2_dfrbp_1 _15492_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net250),
    .D(_00939_),
    .Q_N(_06372_),
    .Q(\mem.mem[105][4] ));
 sg13g2_dfrbp_1 _15493_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net249),
    .D(_00940_),
    .Q_N(_06371_),
    .Q(\mem.mem[105][5] ));
 sg13g2_dfrbp_1 _15494_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net248),
    .D(_00941_),
    .Q_N(_06370_),
    .Q(\mem.mem[105][6] ));
 sg13g2_dfrbp_1 _15495_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net247),
    .D(_00942_),
    .Q_N(_06369_),
    .Q(\mem.mem[105][7] ));
 sg13g2_dfrbp_1 _15496_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net246),
    .D(_00943_),
    .Q_N(_06368_),
    .Q(\mem.mem[106][0] ));
 sg13g2_dfrbp_1 _15497_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net245),
    .D(_00944_),
    .Q_N(_06367_),
    .Q(\mem.mem[106][1] ));
 sg13g2_dfrbp_1 _15498_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net244),
    .D(_00945_),
    .Q_N(_06366_),
    .Q(\mem.mem[106][2] ));
 sg13g2_dfrbp_1 _15499_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net243),
    .D(_00946_),
    .Q_N(_06365_),
    .Q(\mem.mem[106][3] ));
 sg13g2_dfrbp_1 _15500_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net242),
    .D(_00947_),
    .Q_N(_06364_),
    .Q(\mem.mem[106][4] ));
 sg13g2_dfrbp_1 _15501_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net241),
    .D(_00948_),
    .Q_N(_06363_),
    .Q(\mem.mem[106][5] ));
 sg13g2_dfrbp_1 _15502_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net240),
    .D(_00949_),
    .Q_N(_06362_),
    .Q(\mem.mem[106][6] ));
 sg13g2_dfrbp_1 _15503_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net239),
    .D(_00950_),
    .Q_N(_06361_),
    .Q(\mem.mem[106][7] ));
 sg13g2_dfrbp_1 _15504_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net238),
    .D(_00951_),
    .Q_N(_06360_),
    .Q(\mem.mem[107][0] ));
 sg13g2_dfrbp_1 _15505_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net237),
    .D(_00952_),
    .Q_N(_06359_),
    .Q(\mem.mem[107][1] ));
 sg13g2_dfrbp_1 _15506_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net236),
    .D(_00953_),
    .Q_N(_06358_),
    .Q(\mem.mem[107][2] ));
 sg13g2_dfrbp_1 _15507_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net235),
    .D(_00954_),
    .Q_N(_06357_),
    .Q(\mem.mem[107][3] ));
 sg13g2_dfrbp_1 _15508_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net234),
    .D(_00955_),
    .Q_N(_06356_),
    .Q(\mem.mem[107][4] ));
 sg13g2_dfrbp_1 _15509_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net233),
    .D(_00956_),
    .Q_N(_06355_),
    .Q(\mem.mem[107][5] ));
 sg13g2_dfrbp_1 _15510_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net232),
    .D(_00957_),
    .Q_N(_06354_),
    .Q(\mem.mem[107][6] ));
 sg13g2_dfrbp_1 _15511_ (.CLK(clknet_leaf_113_clk),
    .RESET_B(net231),
    .D(_00958_),
    .Q_N(_06353_),
    .Q(\mem.mem[107][7] ));
 sg13g2_dfrbp_1 _15512_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net230),
    .D(_00959_),
    .Q_N(_06352_),
    .Q(\mem.mem[108][0] ));
 sg13g2_dfrbp_1 _15513_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net229),
    .D(_00960_),
    .Q_N(_06351_),
    .Q(\mem.mem[108][1] ));
 sg13g2_dfrbp_1 _15514_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net228),
    .D(_00961_),
    .Q_N(_06350_),
    .Q(\mem.mem[108][2] ));
 sg13g2_dfrbp_1 _15515_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net227),
    .D(_00962_),
    .Q_N(_06349_),
    .Q(\mem.mem[108][3] ));
 sg13g2_dfrbp_1 _15516_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net226),
    .D(_00963_),
    .Q_N(_06348_),
    .Q(\mem.mem[108][4] ));
 sg13g2_dfrbp_1 _15517_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net225),
    .D(_00964_),
    .Q_N(_06347_),
    .Q(\mem.mem[108][5] ));
 sg13g2_dfrbp_1 _15518_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net224),
    .D(_00965_),
    .Q_N(_06346_),
    .Q(\mem.mem[108][6] ));
 sg13g2_dfrbp_1 _15519_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net223),
    .D(_00966_),
    .Q_N(_06345_),
    .Q(\mem.mem[108][7] ));
 sg13g2_dfrbp_1 _15520_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net222),
    .D(_00967_),
    .Q_N(_06344_),
    .Q(\mem.mem[10][0] ));
 sg13g2_dfrbp_1 _15521_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net221),
    .D(_00968_),
    .Q_N(_06343_),
    .Q(\mem.mem[10][1] ));
 sg13g2_dfrbp_1 _15522_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net220),
    .D(_00969_),
    .Q_N(_06342_),
    .Q(\mem.mem[10][2] ));
 sg13g2_dfrbp_1 _15523_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net219),
    .D(_00970_),
    .Q_N(_06341_),
    .Q(\mem.mem[10][3] ));
 sg13g2_dfrbp_1 _15524_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net218),
    .D(_00971_),
    .Q_N(_06340_),
    .Q(\mem.mem[10][4] ));
 sg13g2_dfrbp_1 _15525_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net217),
    .D(_00972_),
    .Q_N(_06339_),
    .Q(\mem.mem[10][5] ));
 sg13g2_dfrbp_1 _15526_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net216),
    .D(_00973_),
    .Q_N(_06338_),
    .Q(\mem.mem[10][6] ));
 sg13g2_dfrbp_1 _15527_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net215),
    .D(_00974_),
    .Q_N(_06337_),
    .Q(\mem.mem[10][7] ));
 sg13g2_dfrbp_1 _15528_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net214),
    .D(_00975_),
    .Q_N(_06336_),
    .Q(\mem.mem[110][0] ));
 sg13g2_dfrbp_1 _15529_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net213),
    .D(_00976_),
    .Q_N(_06335_),
    .Q(\mem.mem[110][1] ));
 sg13g2_dfrbp_1 _15530_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net212),
    .D(_00977_),
    .Q_N(_06334_),
    .Q(\mem.mem[110][2] ));
 sg13g2_dfrbp_1 _15531_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net211),
    .D(_00978_),
    .Q_N(_06333_),
    .Q(\mem.mem[110][3] ));
 sg13g2_dfrbp_1 _15532_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net210),
    .D(_00979_),
    .Q_N(_06332_),
    .Q(\mem.mem[110][4] ));
 sg13g2_dfrbp_1 _15533_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net209),
    .D(_00980_),
    .Q_N(_06331_),
    .Q(\mem.mem[110][5] ));
 sg13g2_dfrbp_1 _15534_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net208),
    .D(_00981_),
    .Q_N(_06330_),
    .Q(\mem.mem[110][6] ));
 sg13g2_dfrbp_1 _15535_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net207),
    .D(_00982_),
    .Q_N(_06329_),
    .Q(\mem.mem[110][7] ));
 sg13g2_dfrbp_1 _15536_ (.CLK(clknet_leaf_112_clk),
    .RESET_B(net206),
    .D(_00983_),
    .Q_N(_06328_),
    .Q(\mem.mem[111][0] ));
 sg13g2_dfrbp_1 _15537_ (.CLK(clknet_leaf_108_clk),
    .RESET_B(net205),
    .D(_00984_),
    .Q_N(_06327_),
    .Q(\mem.mem[111][1] ));
 sg13g2_dfrbp_1 _15538_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net204),
    .D(_00985_),
    .Q_N(_06326_),
    .Q(\mem.mem[111][2] ));
 sg13g2_dfrbp_1 _15539_ (.CLK(clknet_leaf_111_clk),
    .RESET_B(net203),
    .D(_00986_),
    .Q_N(_06325_),
    .Q(\mem.mem[111][3] ));
 sg13g2_dfrbp_1 _15540_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net202),
    .D(_00987_),
    .Q_N(_06324_),
    .Q(\mem.mem[111][4] ));
 sg13g2_dfrbp_1 _15541_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net201),
    .D(_00988_),
    .Q_N(_06323_),
    .Q(\mem.mem[111][5] ));
 sg13g2_dfrbp_1 _15542_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net200),
    .D(_00989_),
    .Q_N(_06322_),
    .Q(\mem.mem[111][6] ));
 sg13g2_dfrbp_1 _15543_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net199),
    .D(_00990_),
    .Q_N(_06321_),
    .Q(\mem.mem[111][7] ));
 sg13g2_dfrbp_1 _15544_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net198),
    .D(_00991_),
    .Q_N(_06320_),
    .Q(\mem.mem[112][0] ));
 sg13g2_dfrbp_1 _15545_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net197),
    .D(_00992_),
    .Q_N(_06319_),
    .Q(\mem.mem[112][1] ));
 sg13g2_dfrbp_1 _15546_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net196),
    .D(_00993_),
    .Q_N(_06318_),
    .Q(\mem.mem[112][2] ));
 sg13g2_dfrbp_1 _15547_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net195),
    .D(_00994_),
    .Q_N(_06317_),
    .Q(\mem.mem[112][3] ));
 sg13g2_dfrbp_1 _15548_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net194),
    .D(_00995_),
    .Q_N(_06316_),
    .Q(\mem.mem[112][4] ));
 sg13g2_dfrbp_1 _15549_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net193),
    .D(_00996_),
    .Q_N(_06315_),
    .Q(\mem.mem[112][5] ));
 sg13g2_dfrbp_1 _15550_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net192),
    .D(_00997_),
    .Q_N(_06314_),
    .Q(\mem.mem[112][6] ));
 sg13g2_dfrbp_1 _15551_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net191),
    .D(_00998_),
    .Q_N(_06313_),
    .Q(\mem.mem[112][7] ));
 sg13g2_dfrbp_1 _15552_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net190),
    .D(_00999_),
    .Q_N(_06312_),
    .Q(\mem.mem[113][0] ));
 sg13g2_dfrbp_1 _15553_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net189),
    .D(_01000_),
    .Q_N(_06311_),
    .Q(\mem.mem[113][1] ));
 sg13g2_dfrbp_1 _15554_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net188),
    .D(_01001_),
    .Q_N(_06310_),
    .Q(\mem.mem[113][2] ));
 sg13g2_dfrbp_1 _15555_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net187),
    .D(_01002_),
    .Q_N(_06309_),
    .Q(\mem.mem[113][3] ));
 sg13g2_dfrbp_1 _15556_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net186),
    .D(_01003_),
    .Q_N(_06308_),
    .Q(\mem.mem[113][4] ));
 sg13g2_dfrbp_1 _15557_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net185),
    .D(_01004_),
    .Q_N(_06307_),
    .Q(\mem.mem[113][5] ));
 sg13g2_dfrbp_1 _15558_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net184),
    .D(_01005_),
    .Q_N(_06306_),
    .Q(\mem.mem[113][6] ));
 sg13g2_dfrbp_1 _15559_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net183),
    .D(_01006_),
    .Q_N(_06305_),
    .Q(\mem.mem[113][7] ));
 sg13g2_dfrbp_1 _15560_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net182),
    .D(_01007_),
    .Q_N(_06304_),
    .Q(\mem.mem[114][0] ));
 sg13g2_dfrbp_1 _15561_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net181),
    .D(_01008_),
    .Q_N(_06303_),
    .Q(\mem.mem[114][1] ));
 sg13g2_dfrbp_1 _15562_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net180),
    .D(_01009_),
    .Q_N(_06302_),
    .Q(\mem.mem[114][2] ));
 sg13g2_dfrbp_1 _15563_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net179),
    .D(_01010_),
    .Q_N(_06301_),
    .Q(\mem.mem[114][3] ));
 sg13g2_dfrbp_1 _15564_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net178),
    .D(_01011_),
    .Q_N(_06300_),
    .Q(\mem.mem[114][4] ));
 sg13g2_dfrbp_1 _15565_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net177),
    .D(_01012_),
    .Q_N(_06299_),
    .Q(\mem.mem[114][5] ));
 sg13g2_dfrbp_1 _15566_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net176),
    .D(_01013_),
    .Q_N(_06298_),
    .Q(\mem.mem[114][6] ));
 sg13g2_dfrbp_1 _15567_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net175),
    .D(_01014_),
    .Q_N(_06297_),
    .Q(\mem.mem[114][7] ));
 sg13g2_dfrbp_1 _15568_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net174),
    .D(_01015_),
    .Q_N(_06296_),
    .Q(\mem.mem[115][0] ));
 sg13g2_dfrbp_1 _15569_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net173),
    .D(_01016_),
    .Q_N(_06295_),
    .Q(\mem.mem[115][1] ));
 sg13g2_dfrbp_1 _15570_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net172),
    .D(_01017_),
    .Q_N(_06294_),
    .Q(\mem.mem[115][2] ));
 sg13g2_dfrbp_1 _15571_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net171),
    .D(_01018_),
    .Q_N(_06293_),
    .Q(\mem.mem[115][3] ));
 sg13g2_dfrbp_1 _15572_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net170),
    .D(_01019_),
    .Q_N(_06292_),
    .Q(\mem.mem[115][4] ));
 sg13g2_dfrbp_1 _15573_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net169),
    .D(_01020_),
    .Q_N(_06291_),
    .Q(\mem.mem[115][5] ));
 sg13g2_dfrbp_1 _15574_ (.CLK(clknet_leaf_27_clk),
    .RESET_B(net168),
    .D(_01021_),
    .Q_N(_06290_),
    .Q(\mem.mem[115][6] ));
 sg13g2_dfrbp_1 _15575_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net167),
    .D(_01022_),
    .Q_N(_06289_),
    .Q(\mem.mem[115][7] ));
 sg13g2_dfrbp_1 _15576_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net166),
    .D(_01023_),
    .Q_N(_06288_),
    .Q(\mem.mem[116][0] ));
 sg13g2_dfrbp_1 _15577_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net165),
    .D(_01024_),
    .Q_N(_06287_),
    .Q(\mem.mem[116][1] ));
 sg13g2_dfrbp_1 _15578_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net164),
    .D(_01025_),
    .Q_N(_06286_),
    .Q(\mem.mem[116][2] ));
 sg13g2_dfrbp_1 _15579_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net163),
    .D(_01026_),
    .Q_N(_06285_),
    .Q(\mem.mem[116][3] ));
 sg13g2_dfrbp_1 _15580_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net162),
    .D(_01027_),
    .Q_N(_06284_),
    .Q(\mem.mem[116][4] ));
 sg13g2_dfrbp_1 _15581_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net161),
    .D(_01028_),
    .Q_N(_06283_),
    .Q(\mem.mem[116][5] ));
 sg13g2_dfrbp_1 _15582_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net160),
    .D(_01029_),
    .Q_N(_06282_),
    .Q(\mem.mem[116][6] ));
 sg13g2_dfrbp_1 _15583_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net159),
    .D(_01030_),
    .Q_N(_06281_),
    .Q(\mem.mem[116][7] ));
 sg13g2_dfrbp_1 _15584_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net158),
    .D(_01031_),
    .Q_N(_06280_),
    .Q(\mem.mem[117][0] ));
 sg13g2_dfrbp_1 _15585_ (.CLK(clknet_leaf_21_clk),
    .RESET_B(net157),
    .D(_01032_),
    .Q_N(_06279_),
    .Q(\mem.mem[117][1] ));
 sg13g2_dfrbp_1 _15586_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net156),
    .D(_01033_),
    .Q_N(_06278_),
    .Q(\mem.mem[117][2] ));
 sg13g2_dfrbp_1 _15587_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net155),
    .D(_01034_),
    .Q_N(_06277_),
    .Q(\mem.mem[117][3] ));
 sg13g2_dfrbp_1 _15588_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net154),
    .D(_01035_),
    .Q_N(_06276_),
    .Q(\mem.mem[117][4] ));
 sg13g2_dfrbp_1 _15589_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net153),
    .D(_01036_),
    .Q_N(_06275_),
    .Q(\mem.mem[117][5] ));
 sg13g2_dfrbp_1 _15590_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net152),
    .D(_01037_),
    .Q_N(_06274_),
    .Q(\mem.mem[117][6] ));
 sg13g2_dfrbp_1 _15591_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net151),
    .D(_01038_),
    .Q_N(_06273_),
    .Q(\mem.mem[117][7] ));
 sg13g2_dfrbp_1 _15592_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net150),
    .D(_01039_),
    .Q_N(_06272_),
    .Q(\mem.mem[118][0] ));
 sg13g2_dfrbp_1 _15593_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net149),
    .D(_01040_),
    .Q_N(_06271_),
    .Q(\mem.mem[118][1] ));
 sg13g2_dfrbp_1 _15594_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net148),
    .D(_01041_),
    .Q_N(_06270_),
    .Q(\mem.mem[118][2] ));
 sg13g2_dfrbp_1 _15595_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net147),
    .D(_01042_),
    .Q_N(_06269_),
    .Q(\mem.mem[118][3] ));
 sg13g2_dfrbp_1 _15596_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net146),
    .D(_01043_),
    .Q_N(_06268_),
    .Q(\mem.mem[118][4] ));
 sg13g2_dfrbp_1 _15597_ (.CLK(clknet_leaf_29_clk),
    .RESET_B(net145),
    .D(_01044_),
    .Q_N(_06267_),
    .Q(\mem.mem[118][5] ));
 sg13g2_dfrbp_1 _15598_ (.CLK(clknet_leaf_31_clk),
    .RESET_B(net144),
    .D(_01045_),
    .Q_N(_06266_),
    .Q(\mem.mem[118][6] ));
 sg13g2_dfrbp_1 _15599_ (.CLK(clknet_leaf_28_clk),
    .RESET_B(net143),
    .D(_01046_),
    .Q_N(_06265_),
    .Q(\mem.mem[118][7] ));
 sg13g2_dfrbp_1 _15600_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net142),
    .D(_01047_),
    .Q_N(_06264_),
    .Q(\mem.mem[11][0] ));
 sg13g2_dfrbp_1 _15601_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net141),
    .D(_01048_),
    .Q_N(_06263_),
    .Q(\mem.mem[11][1] ));
 sg13g2_dfrbp_1 _15602_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net140),
    .D(_01049_),
    .Q_N(_06262_),
    .Q(\mem.mem[11][2] ));
 sg13g2_dfrbp_1 _15603_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net139),
    .D(_01050_),
    .Q_N(_06261_),
    .Q(\mem.mem[11][3] ));
 sg13g2_dfrbp_1 _15604_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net138),
    .D(_01051_),
    .Q_N(_06260_),
    .Q(\mem.mem[11][4] ));
 sg13g2_dfrbp_1 _15605_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net137),
    .D(_01052_),
    .Q_N(_06259_),
    .Q(\mem.mem[11][5] ));
 sg13g2_dfrbp_1 _15606_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net136),
    .D(_01053_),
    .Q_N(_06258_),
    .Q(\mem.mem[11][6] ));
 sg13g2_dfrbp_1 _15607_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net135),
    .D(_01054_),
    .Q_N(_06257_),
    .Q(\mem.mem[11][7] ));
 sg13g2_dfrbp_1 _15608_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net134),
    .D(_01055_),
    .Q_N(_06256_),
    .Q(\mem.mem[120][0] ));
 sg13g2_dfrbp_1 _15609_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net133),
    .D(_01056_),
    .Q_N(_06255_),
    .Q(\mem.mem[120][1] ));
 sg13g2_dfrbp_1 _15610_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net132),
    .D(_01057_),
    .Q_N(_06254_),
    .Q(\mem.mem[120][2] ));
 sg13g2_dfrbp_1 _15611_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net131),
    .D(_01058_),
    .Q_N(_06253_),
    .Q(\mem.mem[120][3] ));
 sg13g2_dfrbp_1 _15612_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net130),
    .D(_01059_),
    .Q_N(_06252_),
    .Q(\mem.mem[120][4] ));
 sg13g2_dfrbp_1 _15613_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net129),
    .D(_01060_),
    .Q_N(_06251_),
    .Q(\mem.mem[120][5] ));
 sg13g2_dfrbp_1 _15614_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net128),
    .D(_01061_),
    .Q_N(_06250_),
    .Q(\mem.mem[120][6] ));
 sg13g2_dfrbp_1 _15615_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net127),
    .D(_01062_),
    .Q_N(_06249_),
    .Q(\mem.mem[120][7] ));
 sg13g2_dfrbp_1 _15616_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net126),
    .D(_01063_),
    .Q_N(_06248_),
    .Q(\mem.mem[121][0] ));
 sg13g2_dfrbp_1 _15617_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net125),
    .D(_01064_),
    .Q_N(_06247_),
    .Q(\mem.mem[121][1] ));
 sg13g2_dfrbp_1 _15618_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net124),
    .D(_01065_),
    .Q_N(_06246_),
    .Q(\mem.mem[121][2] ));
 sg13g2_dfrbp_1 _15619_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net123),
    .D(_01066_),
    .Q_N(_06245_),
    .Q(\mem.mem[121][3] ));
 sg13g2_dfrbp_1 _15620_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net122),
    .D(_01067_),
    .Q_N(_06244_),
    .Q(\mem.mem[121][4] ));
 sg13g2_dfrbp_1 _15621_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net121),
    .D(_01068_),
    .Q_N(_06243_),
    .Q(\mem.mem[121][5] ));
 sg13g2_dfrbp_1 _15622_ (.CLK(clknet_leaf_44_clk),
    .RESET_B(net120),
    .D(_01069_),
    .Q_N(_06242_),
    .Q(\mem.mem[121][6] ));
 sg13g2_dfrbp_1 _15623_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net119),
    .D(_01070_),
    .Q_N(_06241_),
    .Q(\mem.mem[121][7] ));
 sg13g2_dfrbp_1 _15624_ (.CLK(clknet_leaf_42_clk),
    .RESET_B(net118),
    .D(_01071_),
    .Q_N(_06240_),
    .Q(\mem.mem[122][0] ));
 sg13g2_dfrbp_1 _15625_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net117),
    .D(_01072_),
    .Q_N(_06239_),
    .Q(\mem.mem[122][1] ));
 sg13g2_dfrbp_1 _15626_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net116),
    .D(_01073_),
    .Q_N(_06238_),
    .Q(\mem.mem[122][2] ));
 sg13g2_dfrbp_1 _15627_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net115),
    .D(_01074_),
    .Q_N(_06237_),
    .Q(\mem.mem[122][3] ));
 sg13g2_dfrbp_1 _15628_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net114),
    .D(_01075_),
    .Q_N(_06236_),
    .Q(\mem.mem[122][4] ));
 sg13g2_dfrbp_1 _15629_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net113),
    .D(_01076_),
    .Q_N(_06235_),
    .Q(\mem.mem[122][5] ));
 sg13g2_dfrbp_1 _15630_ (.CLK(clknet_leaf_45_clk),
    .RESET_B(net112),
    .D(_01077_),
    .Q_N(_06234_),
    .Q(\mem.mem[122][6] ));
 sg13g2_dfrbp_1 _15631_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net111),
    .D(_01078_),
    .Q_N(_06233_),
    .Q(\mem.mem[122][7] ));
 sg13g2_dfrbp_1 _15632_ (.CLK(clknet_leaf_40_clk),
    .RESET_B(net110),
    .D(_01079_),
    .Q_N(_06232_),
    .Q(\mem.mem[123][0] ));
 sg13g2_dfrbp_1 _15633_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net109),
    .D(_01080_),
    .Q_N(_06231_),
    .Q(\mem.mem[123][1] ));
 sg13g2_dfrbp_1 _15634_ (.CLK(clknet_leaf_37_clk),
    .RESET_B(net108),
    .D(_01081_),
    .Q_N(_06230_),
    .Q(\mem.mem[123][2] ));
 sg13g2_dfrbp_1 _15635_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net107),
    .D(_01082_),
    .Q_N(_06229_),
    .Q(\mem.mem[123][3] ));
 sg13g2_dfrbp_1 _15636_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net106),
    .D(_01083_),
    .Q_N(_06228_),
    .Q(\mem.mem[123][4] ));
 sg13g2_dfrbp_1 _15637_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net105),
    .D(_01084_),
    .Q_N(_06227_),
    .Q(\mem.mem[123][5] ));
 sg13g2_dfrbp_1 _15638_ (.CLK(clknet_leaf_38_clk),
    .RESET_B(net104),
    .D(_01085_),
    .Q_N(_06226_),
    .Q(\mem.mem[123][6] ));
 sg13g2_dfrbp_1 _15639_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net103),
    .D(_01086_),
    .Q_N(_06225_),
    .Q(\mem.mem[123][7] ));
 sg13g2_dfrbp_1 _15640_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net102),
    .D(_01087_),
    .Q_N(_06224_),
    .Q(\mem.mem[124][0] ));
 sg13g2_dfrbp_1 _15641_ (.CLK(clknet_leaf_30_clk),
    .RESET_B(net101),
    .D(_01088_),
    .Q_N(_06223_),
    .Q(\mem.mem[124][1] ));
 sg13g2_dfrbp_1 _15642_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net100),
    .D(_01089_),
    .Q_N(_06222_),
    .Q(\mem.mem[124][2] ));
 sg13g2_dfrbp_1 _15643_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net99),
    .D(_01090_),
    .Q_N(_06221_),
    .Q(\mem.mem[124][3] ));
 sg13g2_dfrbp_1 _15644_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net98),
    .D(_01091_),
    .Q_N(_06220_),
    .Q(\mem.mem[124][4] ));
 sg13g2_dfrbp_1 _15645_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net97),
    .D(_01092_),
    .Q_N(_06219_),
    .Q(\mem.mem[124][5] ));
 sg13g2_dfrbp_1 _15646_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net96),
    .D(_01093_),
    .Q_N(_06218_),
    .Q(\mem.mem[124][6] ));
 sg13g2_dfrbp_1 _15647_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net95),
    .D(_01094_),
    .Q_N(_06217_),
    .Q(\mem.mem[124][7] ));
 sg13g2_dfrbp_1 _15648_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net94),
    .D(_01095_),
    .Q_N(_06216_),
    .Q(\mem.mem[125][0] ));
 sg13g2_dfrbp_1 _15649_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net93),
    .D(_01096_),
    .Q_N(_06215_),
    .Q(\mem.mem[125][1] ));
 sg13g2_dfrbp_1 _15650_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net92),
    .D(_01097_),
    .Q_N(_06214_),
    .Q(\mem.mem[125][2] ));
 sg13g2_dfrbp_1 _15651_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net91),
    .D(_01098_),
    .Q_N(_06213_),
    .Q(\mem.mem[125][3] ));
 sg13g2_dfrbp_1 _15652_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net90),
    .D(_01099_),
    .Q_N(_06212_),
    .Q(\mem.mem[125][4] ));
 sg13g2_dfrbp_1 _15653_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net89),
    .D(_01100_),
    .Q_N(_06211_),
    .Q(\mem.mem[125][5] ));
 sg13g2_dfrbp_1 _15654_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net88),
    .D(_01101_),
    .Q_N(_06210_),
    .Q(\mem.mem[125][6] ));
 sg13g2_dfrbp_1 _15655_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net87),
    .D(_01102_),
    .Q_N(_06209_),
    .Q(\mem.mem[125][7] ));
 sg13g2_dfrbp_1 _15656_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net86),
    .D(_01103_),
    .Q_N(_06208_),
    .Q(\mem.mem[126][0] ));
 sg13g2_dfrbp_1 _15657_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net85),
    .D(_01104_),
    .Q_N(_06207_),
    .Q(\mem.mem[126][1] ));
 sg13g2_dfrbp_1 _15658_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net84),
    .D(_01105_),
    .Q_N(_06206_),
    .Q(\mem.mem[126][2] ));
 sg13g2_dfrbp_1 _15659_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net83),
    .D(_01106_),
    .Q_N(_06205_),
    .Q(\mem.mem[126][3] ));
 sg13g2_dfrbp_1 _15660_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net82),
    .D(_01107_),
    .Q_N(_06204_),
    .Q(\mem.mem[126][4] ));
 sg13g2_dfrbp_1 _15661_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net81),
    .D(_01108_),
    .Q_N(_06203_),
    .Q(\mem.mem[126][5] ));
 sg13g2_dfrbp_1 _15662_ (.CLK(clknet_leaf_35_clk),
    .RESET_B(net80),
    .D(_01109_),
    .Q_N(_06202_),
    .Q(\mem.mem[126][6] ));
 sg13g2_dfrbp_1 _15663_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net79),
    .D(_01110_),
    .Q_N(_06201_),
    .Q(\mem.mem[126][7] ));
 sg13g2_dfrbp_1 _15664_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net78),
    .D(_01111_),
    .Q_N(_06200_),
    .Q(\mem.mem[127][0] ));
 sg13g2_dfrbp_1 _15665_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net77),
    .D(_01112_),
    .Q_N(_06199_),
    .Q(\mem.mem[127][1] ));
 sg13g2_dfrbp_1 _15666_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net76),
    .D(_01113_),
    .Q_N(_06198_),
    .Q(\mem.mem[127][2] ));
 sg13g2_dfrbp_1 _15667_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net75),
    .D(_01114_),
    .Q_N(_06197_),
    .Q(\mem.mem[127][3] ));
 sg13g2_dfrbp_1 _15668_ (.CLK(clknet_leaf_39_clk),
    .RESET_B(net74),
    .D(_01115_),
    .Q_N(_06196_),
    .Q(\mem.mem[127][4] ));
 sg13g2_dfrbp_1 _15669_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net73),
    .D(_01116_),
    .Q_N(_06195_),
    .Q(\mem.mem[127][5] ));
 sg13g2_dfrbp_1 _15670_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net72),
    .D(_01117_),
    .Q_N(_06194_),
    .Q(\mem.mem[127][6] ));
 sg13g2_dfrbp_1 _15671_ (.CLK(clknet_leaf_36_clk),
    .RESET_B(net71),
    .D(_01118_),
    .Q_N(_06193_),
    .Q(\mem.mem[127][7] ));
 sg13g2_dfrbp_1 _15672_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net70),
    .D(_01119_),
    .Q_N(_06192_),
    .Q(\mem.mem[128][0] ));
 sg13g2_dfrbp_1 _15673_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net69),
    .D(_01120_),
    .Q_N(_06191_),
    .Q(\mem.mem[128][1] ));
 sg13g2_dfrbp_1 _15674_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net68),
    .D(_01121_),
    .Q_N(_06190_),
    .Q(\mem.mem[128][2] ));
 sg13g2_dfrbp_1 _15675_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net67),
    .D(_01122_),
    .Q_N(_06189_),
    .Q(\mem.mem[128][3] ));
 sg13g2_dfrbp_1 _15676_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net66),
    .D(_01123_),
    .Q_N(_06188_),
    .Q(\mem.mem[128][4] ));
 sg13g2_dfrbp_1 _15677_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net65),
    .D(_01124_),
    .Q_N(_06187_),
    .Q(\mem.mem[128][5] ));
 sg13g2_dfrbp_1 _15678_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net64),
    .D(_01125_),
    .Q_N(_06186_),
    .Q(\mem.mem[128][6] ));
 sg13g2_dfrbp_1 _15679_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net63),
    .D(_01126_),
    .Q_N(_06185_),
    .Q(\mem.mem[128][7] ));
 sg13g2_dfrbp_1 _15680_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net62),
    .D(_01127_),
    .Q_N(_06184_),
    .Q(\mem.mem[12][0] ));
 sg13g2_dfrbp_1 _15681_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net61),
    .D(_01128_),
    .Q_N(_06183_),
    .Q(\mem.mem[12][1] ));
 sg13g2_dfrbp_1 _15682_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net60),
    .D(_01129_),
    .Q_N(_06182_),
    .Q(\mem.mem[12][2] ));
 sg13g2_dfrbp_1 _15683_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net59),
    .D(_01130_),
    .Q_N(_06181_),
    .Q(\mem.mem[12][3] ));
 sg13g2_dfrbp_1 _15684_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net58),
    .D(_01131_),
    .Q_N(_06180_),
    .Q(\mem.mem[12][4] ));
 sg13g2_dfrbp_1 _15685_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net57),
    .D(_01132_),
    .Q_N(_06179_),
    .Q(\mem.mem[12][5] ));
 sg13g2_dfrbp_1 _15686_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net56),
    .D(_01133_),
    .Q_N(_06178_),
    .Q(\mem.mem[12][6] ));
 sg13g2_dfrbp_1 _15687_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net55),
    .D(_01134_),
    .Q_N(_06177_),
    .Q(\mem.mem[12][7] ));
 sg13g2_dfrbp_1 _15688_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net54),
    .D(_01135_),
    .Q_N(_06176_),
    .Q(\mem.mem[130][0] ));
 sg13g2_dfrbp_1 _15689_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net53),
    .D(_01136_),
    .Q_N(_06175_),
    .Q(\mem.mem[130][1] ));
 sg13g2_dfrbp_1 _15690_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net52),
    .D(_01137_),
    .Q_N(_06174_),
    .Q(\mem.mem[130][2] ));
 sg13g2_dfrbp_1 _15691_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net51),
    .D(_01138_),
    .Q_N(_06173_),
    .Q(\mem.mem[130][3] ));
 sg13g2_dfrbp_1 _15692_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net50),
    .D(_01139_),
    .Q_N(_06172_),
    .Q(\mem.mem[130][4] ));
 sg13g2_dfrbp_1 _15693_ (.CLK(clknet_leaf_167_clk),
    .RESET_B(net49),
    .D(_01140_),
    .Q_N(_06171_),
    .Q(\mem.mem[130][5] ));
 sg13g2_dfrbp_1 _15694_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net48),
    .D(_01141_),
    .Q_N(_06170_),
    .Q(\mem.mem[130][6] ));
 sg13g2_dfrbp_1 _15695_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net47),
    .D(_01142_),
    .Q_N(_06169_),
    .Q(\mem.mem[130][7] ));
 sg13g2_dfrbp_1 _15696_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net46),
    .D(_01143_),
    .Q_N(_06168_),
    .Q(\mem.mem[131][0] ));
 sg13g2_dfrbp_1 _15697_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net45),
    .D(_01144_),
    .Q_N(_06167_),
    .Q(\mem.mem[131][1] ));
 sg13g2_dfrbp_1 _15698_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net44),
    .D(_01145_),
    .Q_N(_06166_),
    .Q(\mem.mem[131][2] ));
 sg13g2_dfrbp_1 _15699_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net43),
    .D(_01146_),
    .Q_N(_06165_),
    .Q(\mem.mem[131][3] ));
 sg13g2_dfrbp_1 _15700_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net42),
    .D(_01147_),
    .Q_N(_06164_),
    .Q(\mem.mem[131][4] ));
 sg13g2_dfrbp_1 _15701_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net41),
    .D(_01148_),
    .Q_N(_06163_),
    .Q(\mem.mem[131][5] ));
 sg13g2_dfrbp_1 _15702_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net40),
    .D(_01149_),
    .Q_N(_06162_),
    .Q(\mem.mem[131][6] ));
 sg13g2_dfrbp_1 _15703_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net39),
    .D(_01150_),
    .Q_N(_06161_),
    .Q(\mem.mem[131][7] ));
 sg13g2_dfrbp_1 _15704_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net38),
    .D(_01151_),
    .Q_N(_06160_),
    .Q(\mem.mem[132][0] ));
 sg13g2_dfrbp_1 _15705_ (.CLK(clknet_leaf_164_clk),
    .RESET_B(net37),
    .D(_01152_),
    .Q_N(_06159_),
    .Q(\mem.mem[132][1] ));
 sg13g2_dfrbp_1 _15706_ (.CLK(clknet_leaf_163_clk),
    .RESET_B(net36),
    .D(_01153_),
    .Q_N(_06158_),
    .Q(\mem.mem[132][2] ));
 sg13g2_dfrbp_1 _15707_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net35),
    .D(_01154_),
    .Q_N(_06157_),
    .Q(\mem.mem[132][3] ));
 sg13g2_dfrbp_1 _15708_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net34),
    .D(_01155_),
    .Q_N(_06156_),
    .Q(\mem.mem[132][4] ));
 sg13g2_dfrbp_1 _15709_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net33),
    .D(_01156_),
    .Q_N(_06155_),
    .Q(\mem.mem[132][5] ));
 sg13g2_dfrbp_1 _15710_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net32),
    .D(_01157_),
    .Q_N(_06154_),
    .Q(\mem.mem[132][6] ));
 sg13g2_dfrbp_1 _15711_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net31),
    .D(_01158_),
    .Q_N(_06153_),
    .Q(\mem.mem[132][7] ));
 sg13g2_dfrbp_1 _15712_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net30),
    .D(_01159_),
    .Q_N(_06152_),
    .Q(\mem.mem[133][0] ));
 sg13g2_dfrbp_1 _15713_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net29),
    .D(_01160_),
    .Q_N(_06151_),
    .Q(\mem.mem[133][1] ));
 sg13g2_dfrbp_1 _15714_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net28),
    .D(_01161_),
    .Q_N(_06150_),
    .Q(\mem.mem[133][2] ));
 sg13g2_dfrbp_1 _15715_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net27),
    .D(_01162_),
    .Q_N(_06149_),
    .Q(\mem.mem[133][3] ));
 sg13g2_dfrbp_1 _15716_ (.CLK(clknet_leaf_149_clk),
    .RESET_B(net26),
    .D(_01163_),
    .Q_N(_06148_),
    .Q(\mem.mem[133][4] ));
 sg13g2_dfrbp_1 _15717_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2127),
    .D(_01164_),
    .Q_N(_06147_),
    .Q(\mem.mem[133][5] ));
 sg13g2_dfrbp_1 _15718_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2126),
    .D(_01165_),
    .Q_N(_06146_),
    .Q(\mem.mem[133][6] ));
 sg13g2_dfrbp_1 _15719_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2125),
    .D(_01166_),
    .Q_N(_06145_),
    .Q(\mem.mem[133][7] ));
 sg13g2_dfrbp_1 _15720_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2124),
    .D(_01167_),
    .Q_N(_06144_),
    .Q(\mem.mem[134][0] ));
 sg13g2_dfrbp_1 _15721_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2123),
    .D(_01168_),
    .Q_N(_06143_),
    .Q(\mem.mem[134][1] ));
 sg13g2_dfrbp_1 _15722_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2122),
    .D(_01169_),
    .Q_N(_06142_),
    .Q(\mem.mem[134][2] ));
 sg13g2_dfrbp_1 _15723_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2121),
    .D(_01170_),
    .Q_N(_06141_),
    .Q(\mem.mem[134][3] ));
 sg13g2_dfrbp_1 _15724_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2120),
    .D(_01171_),
    .Q_N(_06140_),
    .Q(\mem.mem[134][4] ));
 sg13g2_dfrbp_1 _15725_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2119),
    .D(_01172_),
    .Q_N(_06139_),
    .Q(\mem.mem[134][5] ));
 sg13g2_dfrbp_1 _15726_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2118),
    .D(_01173_),
    .Q_N(_06138_),
    .Q(\mem.mem[134][6] ));
 sg13g2_dfrbp_1 _15727_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2117),
    .D(_01174_),
    .Q_N(_06137_),
    .Q(\mem.mem[134][7] ));
 sg13g2_dfrbp_1 _15728_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2116),
    .D(_01175_),
    .Q_N(_06136_),
    .Q(\mem.mem[135][0] ));
 sg13g2_dfrbp_1 _15729_ (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2115),
    .D(_01176_),
    .Q_N(_06135_),
    .Q(\mem.mem[135][1] ));
 sg13g2_dfrbp_1 _15730_ (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2114),
    .D(_01177_),
    .Q_N(_06134_),
    .Q(\mem.mem[135][2] ));
 sg13g2_dfrbp_1 _15731_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2113),
    .D(_01178_),
    .Q_N(_06133_),
    .Q(\mem.mem[135][3] ));
 sg13g2_dfrbp_1 _15732_ (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2112),
    .D(_01179_),
    .Q_N(_06132_),
    .Q(\mem.mem[135][4] ));
 sg13g2_dfrbp_1 _15733_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2111),
    .D(_01180_),
    .Q_N(_06131_),
    .Q(\mem.mem[135][5] ));
 sg13g2_dfrbp_1 _15734_ (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2110),
    .D(_01181_),
    .Q_N(_06130_),
    .Q(\mem.mem[135][6] ));
 sg13g2_dfrbp_1 _15735_ (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2109),
    .D(_01182_),
    .Q_N(_06129_),
    .Q(\mem.mem[135][7] ));
 sg13g2_dfrbp_1 _15736_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2108),
    .D(_01183_),
    .Q_N(_06128_),
    .Q(\mem.mem[136][0] ));
 sg13g2_dfrbp_1 _15737_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2107),
    .D(_01184_),
    .Q_N(_06127_),
    .Q(\mem.mem[136][1] ));
 sg13g2_dfrbp_1 _15738_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2106),
    .D(_01185_),
    .Q_N(_06126_),
    .Q(\mem.mem[136][2] ));
 sg13g2_dfrbp_1 _15739_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2105),
    .D(_01186_),
    .Q_N(_06125_),
    .Q(\mem.mem[136][3] ));
 sg13g2_dfrbp_1 _15740_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2104),
    .D(_01187_),
    .Q_N(_06124_),
    .Q(\mem.mem[136][4] ));
 sg13g2_dfrbp_1 _15741_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2103),
    .D(_01188_),
    .Q_N(_06123_),
    .Q(\mem.mem[136][5] ));
 sg13g2_dfrbp_1 _15742_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2102),
    .D(_01189_),
    .Q_N(_06122_),
    .Q(\mem.mem[136][6] ));
 sg13g2_dfrbp_1 _15743_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2101),
    .D(_01190_),
    .Q_N(_06121_),
    .Q(\mem.mem[136][7] ));
 sg13g2_dfrbp_1 _15744_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2100),
    .D(_01191_),
    .Q_N(_06120_),
    .Q(\mem.mem[137][0] ));
 sg13g2_dfrbp_1 _15745_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2099),
    .D(_01192_),
    .Q_N(_06119_),
    .Q(\mem.mem[137][1] ));
 sg13g2_dfrbp_1 _15746_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2098),
    .D(_01193_),
    .Q_N(_06118_),
    .Q(\mem.mem[137][2] ));
 sg13g2_dfrbp_1 _15747_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2097),
    .D(_01194_),
    .Q_N(_06117_),
    .Q(\mem.mem[137][3] ));
 sg13g2_dfrbp_1 _15748_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2096),
    .D(_01195_),
    .Q_N(_06116_),
    .Q(\mem.mem[137][4] ));
 sg13g2_dfrbp_1 _15749_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2095),
    .D(_01196_),
    .Q_N(_06115_),
    .Q(\mem.mem[137][5] ));
 sg13g2_dfrbp_1 _15750_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2094),
    .D(_01197_),
    .Q_N(_06114_),
    .Q(\mem.mem[137][6] ));
 sg13g2_dfrbp_1 _15751_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2093),
    .D(_01198_),
    .Q_N(_06113_),
    .Q(\mem.mem[137][7] ));
 sg13g2_dfrbp_1 _15752_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2092),
    .D(_01199_),
    .Q_N(_06112_),
    .Q(\mem.mem[138][0] ));
 sg13g2_dfrbp_1 _15753_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2091),
    .D(_01200_),
    .Q_N(_06111_),
    .Q(\mem.mem[138][1] ));
 sg13g2_dfrbp_1 _15754_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2090),
    .D(_01201_),
    .Q_N(_06110_),
    .Q(\mem.mem[138][2] ));
 sg13g2_dfrbp_1 _15755_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2089),
    .D(_01202_),
    .Q_N(_06109_),
    .Q(\mem.mem[138][3] ));
 sg13g2_dfrbp_1 _15756_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2088),
    .D(_01203_),
    .Q_N(_06108_),
    .Q(\mem.mem[138][4] ));
 sg13g2_dfrbp_1 _15757_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2087),
    .D(_01204_),
    .Q_N(_06107_),
    .Q(\mem.mem[138][5] ));
 sg13g2_dfrbp_1 _15758_ (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2086),
    .D(_01205_),
    .Q_N(_06106_),
    .Q(\mem.mem[138][6] ));
 sg13g2_dfrbp_1 _15759_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2085),
    .D(_01206_),
    .Q_N(_06105_),
    .Q(\mem.mem[138][7] ));
 sg13g2_dfrbp_1 _15760_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2084),
    .D(_01207_),
    .Q_N(_06104_),
    .Q(\mem.mem[13][0] ));
 sg13g2_dfrbp_1 _15761_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2083),
    .D(_01208_),
    .Q_N(_06103_),
    .Q(\mem.mem[13][1] ));
 sg13g2_dfrbp_1 _15762_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2082),
    .D(_01209_),
    .Q_N(_06102_),
    .Q(\mem.mem[13][2] ));
 sg13g2_dfrbp_1 _15763_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2081),
    .D(_01210_),
    .Q_N(_06101_),
    .Q(\mem.mem[13][3] ));
 sg13g2_dfrbp_1 _15764_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2080),
    .D(_01211_),
    .Q_N(_06100_),
    .Q(\mem.mem[13][4] ));
 sg13g2_dfrbp_1 _15765_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2079),
    .D(_01212_),
    .Q_N(_06099_),
    .Q(\mem.mem[13][5] ));
 sg13g2_dfrbp_1 _15766_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2078),
    .D(_01213_),
    .Q_N(_06098_),
    .Q(\mem.mem[13][6] ));
 sg13g2_dfrbp_1 _15767_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2077),
    .D(_01214_),
    .Q_N(_06097_),
    .Q(\mem.mem[13][7] ));
 sg13g2_dfrbp_1 _15768_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2076),
    .D(_01215_),
    .Q_N(_06096_),
    .Q(\mem.mem[140][0] ));
 sg13g2_dfrbp_1 _15769_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2075),
    .D(_01216_),
    .Q_N(_06095_),
    .Q(\mem.mem[140][1] ));
 sg13g2_dfrbp_1 _15770_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2074),
    .D(_01217_),
    .Q_N(_06094_),
    .Q(\mem.mem[140][2] ));
 sg13g2_dfrbp_1 _15771_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2073),
    .D(_01218_),
    .Q_N(_06093_),
    .Q(\mem.mem[140][3] ));
 sg13g2_dfrbp_1 _15772_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2072),
    .D(_01219_),
    .Q_N(_06092_),
    .Q(\mem.mem[140][4] ));
 sg13g2_dfrbp_1 _15773_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2071),
    .D(_01220_),
    .Q_N(_06091_),
    .Q(\mem.mem[140][5] ));
 sg13g2_dfrbp_1 _15774_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2070),
    .D(_01221_),
    .Q_N(_06090_),
    .Q(\mem.mem[140][6] ));
 sg13g2_dfrbp_1 _15775_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2069),
    .D(_01222_),
    .Q_N(_06089_),
    .Q(\mem.mem[140][7] ));
 sg13g2_dfrbp_1 _15776_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2068),
    .D(_01223_),
    .Q_N(_06088_),
    .Q(\mem.mem[141][0] ));
 sg13g2_dfrbp_1 _15777_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2067),
    .D(_01224_),
    .Q_N(_06087_),
    .Q(\mem.mem[141][1] ));
 sg13g2_dfrbp_1 _15778_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2066),
    .D(_01225_),
    .Q_N(_06086_),
    .Q(\mem.mem[141][2] ));
 sg13g2_dfrbp_1 _15779_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2065),
    .D(_01226_),
    .Q_N(_06085_),
    .Q(\mem.mem[141][3] ));
 sg13g2_dfrbp_1 _15780_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2064),
    .D(_01227_),
    .Q_N(_06084_),
    .Q(\mem.mem[141][4] ));
 sg13g2_dfrbp_1 _15781_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2063),
    .D(_01228_),
    .Q_N(_06083_),
    .Q(\mem.mem[141][5] ));
 sg13g2_dfrbp_1 _15782_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2062),
    .D(_01229_),
    .Q_N(_06082_),
    .Q(\mem.mem[141][6] ));
 sg13g2_dfrbp_1 _15783_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2061),
    .D(_01230_),
    .Q_N(_06081_),
    .Q(\mem.mem[141][7] ));
 sg13g2_dfrbp_1 _15784_ (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2060),
    .D(_01231_),
    .Q_N(_06080_),
    .Q(\mem.mem[142][0] ));
 sg13g2_dfrbp_1 _15785_ (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2059),
    .D(_01232_),
    .Q_N(_06079_),
    .Q(\mem.mem[142][1] ));
 sg13g2_dfrbp_1 _15786_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2058),
    .D(_01233_),
    .Q_N(_06078_),
    .Q(\mem.mem[142][2] ));
 sg13g2_dfrbp_1 _15787_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2057),
    .D(_01234_),
    .Q_N(_06077_),
    .Q(\mem.mem[142][3] ));
 sg13g2_dfrbp_1 _15788_ (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2056),
    .D(_01235_),
    .Q_N(_06076_),
    .Q(\mem.mem[142][4] ));
 sg13g2_dfrbp_1 _15789_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2055),
    .D(_01236_),
    .Q_N(_06075_),
    .Q(\mem.mem[142][5] ));
 sg13g2_dfrbp_1 _15790_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2054),
    .D(_01237_),
    .Q_N(_06074_),
    .Q(\mem.mem[142][6] ));
 sg13g2_dfrbp_1 _15791_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2053),
    .D(_01238_),
    .Q_N(_06073_),
    .Q(\mem.mem[142][7] ));
 sg13g2_dfrbp_1 _15792_ (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2052),
    .D(_01239_),
    .Q_N(_06072_),
    .Q(\mem.mem[143][0] ));
 sg13g2_dfrbp_1 _15793_ (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2051),
    .D(_01240_),
    .Q_N(_06071_),
    .Q(\mem.mem[143][1] ));
 sg13g2_dfrbp_1 _15794_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2050),
    .D(_01241_),
    .Q_N(_06070_),
    .Q(\mem.mem[143][2] ));
 sg13g2_dfrbp_1 _15795_ (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2049),
    .D(_01242_),
    .Q_N(_06069_),
    .Q(\mem.mem[143][3] ));
 sg13g2_dfrbp_1 _15796_ (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2048),
    .D(_01243_),
    .Q_N(_06068_),
    .Q(\mem.mem[143][4] ));
 sg13g2_dfrbp_1 _15797_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2047),
    .D(_01244_),
    .Q_N(_06067_),
    .Q(\mem.mem[143][5] ));
 sg13g2_dfrbp_1 _15798_ (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2046),
    .D(_01245_),
    .Q_N(_06066_),
    .Q(\mem.mem[143][6] ));
 sg13g2_dfrbp_1 _15799_ (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2045),
    .D(_01246_),
    .Q_N(_06065_),
    .Q(\mem.mem[143][7] ));
 sg13g2_dfrbp_1 _15800_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2044),
    .D(_01247_),
    .Q_N(_06064_),
    .Q(\mem.mem[144][0] ));
 sg13g2_dfrbp_1 _15801_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2043),
    .D(_01248_),
    .Q_N(_06063_),
    .Q(\mem.mem[144][1] ));
 sg13g2_dfrbp_1 _15802_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2042),
    .D(_01249_),
    .Q_N(_06062_),
    .Q(\mem.mem[144][2] ));
 sg13g2_dfrbp_1 _15803_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2041),
    .D(_01250_),
    .Q_N(_06061_),
    .Q(\mem.mem[144][3] ));
 sg13g2_dfrbp_1 _15804_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2040),
    .D(_01251_),
    .Q_N(_06060_),
    .Q(\mem.mem[144][4] ));
 sg13g2_dfrbp_1 _15805_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2039),
    .D(_01252_),
    .Q_N(_06059_),
    .Q(\mem.mem[144][5] ));
 sg13g2_dfrbp_1 _15806_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2038),
    .D(_01253_),
    .Q_N(_06058_),
    .Q(\mem.mem[144][6] ));
 sg13g2_dfrbp_1 _15807_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2037),
    .D(_01254_),
    .Q_N(_06057_),
    .Q(\mem.mem[144][7] ));
 sg13g2_dfrbp_1 _15808_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2036),
    .D(_01255_),
    .Q_N(_06056_),
    .Q(\mem.mem[145][0] ));
 sg13g2_dfrbp_1 _15809_ (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2035),
    .D(_01256_),
    .Q_N(_06055_),
    .Q(\mem.mem[145][1] ));
 sg13g2_dfrbp_1 _15810_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2034),
    .D(_01257_),
    .Q_N(_06054_),
    .Q(\mem.mem[145][2] ));
 sg13g2_dfrbp_1 _15811_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2033),
    .D(_01258_),
    .Q_N(_06053_),
    .Q(\mem.mem[145][3] ));
 sg13g2_dfrbp_1 _15812_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2032),
    .D(_01259_),
    .Q_N(_06052_),
    .Q(\mem.mem[145][4] ));
 sg13g2_dfrbp_1 _15813_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2031),
    .D(_01260_),
    .Q_N(_06051_),
    .Q(\mem.mem[145][5] ));
 sg13g2_dfrbp_1 _15814_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2030),
    .D(_01261_),
    .Q_N(_06050_),
    .Q(\mem.mem[145][6] ));
 sg13g2_dfrbp_1 _15815_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2029),
    .D(_01262_),
    .Q_N(_06049_),
    .Q(\mem.mem[145][7] ));
 sg13g2_dfrbp_1 _15816_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2028),
    .D(_01263_),
    .Q_N(_06048_),
    .Q(\mem.mem[146][0] ));
 sg13g2_dfrbp_1 _15817_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2027),
    .D(_01264_),
    .Q_N(_06047_),
    .Q(\mem.mem[146][1] ));
 sg13g2_dfrbp_1 _15818_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2026),
    .D(_01265_),
    .Q_N(_06046_),
    .Q(\mem.mem[146][2] ));
 sg13g2_dfrbp_1 _15819_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2025),
    .D(_01266_),
    .Q_N(_06045_),
    .Q(\mem.mem[146][3] ));
 sg13g2_dfrbp_1 _15820_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2024),
    .D(_01267_),
    .Q_N(_06044_),
    .Q(\mem.mem[146][4] ));
 sg13g2_dfrbp_1 _15821_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2023),
    .D(_01268_),
    .Q_N(_06043_),
    .Q(\mem.mem[146][5] ));
 sg13g2_dfrbp_1 _15822_ (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2022),
    .D(_01269_),
    .Q_N(_06042_),
    .Q(\mem.mem[146][6] ));
 sg13g2_dfrbp_1 _15823_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2021),
    .D(_01270_),
    .Q_N(_06041_),
    .Q(\mem.mem[146][7] ));
 sg13g2_dfrbp_1 _15824_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2020),
    .D(_01271_),
    .Q_N(_06040_),
    .Q(\mem.mem[147][0] ));
 sg13g2_dfrbp_1 _15825_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2019),
    .D(_01272_),
    .Q_N(_06039_),
    .Q(\mem.mem[147][1] ));
 sg13g2_dfrbp_1 _15826_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2018),
    .D(_01273_),
    .Q_N(_06038_),
    .Q(\mem.mem[147][2] ));
 sg13g2_dfrbp_1 _15827_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2017),
    .D(_01274_),
    .Q_N(_06037_),
    .Q(\mem.mem[147][3] ));
 sg13g2_dfrbp_1 _15828_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2016),
    .D(_01275_),
    .Q_N(_06036_),
    .Q(\mem.mem[147][4] ));
 sg13g2_dfrbp_1 _15829_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2015),
    .D(_01276_),
    .Q_N(_06035_),
    .Q(\mem.mem[147][5] ));
 sg13g2_dfrbp_1 _15830_ (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2014),
    .D(_01277_),
    .Q_N(_06034_),
    .Q(\mem.mem[147][6] ));
 sg13g2_dfrbp_1 _15831_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net2013),
    .D(_01278_),
    .Q_N(_06033_),
    .Q(\mem.mem[147][7] ));
 sg13g2_dfrbp_1 _15832_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2012),
    .D(_01279_),
    .Q_N(_06032_),
    .Q(\mem.mem[148][0] ));
 sg13g2_dfrbp_1 _15833_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2011),
    .D(_01280_),
    .Q_N(_06031_),
    .Q(\mem.mem[148][1] ));
 sg13g2_dfrbp_1 _15834_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2010),
    .D(_01281_),
    .Q_N(_06030_),
    .Q(\mem.mem[148][2] ));
 sg13g2_dfrbp_1 _15835_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2009),
    .D(_01282_),
    .Q_N(_06029_),
    .Q(\mem.mem[148][3] ));
 sg13g2_dfrbp_1 _15836_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2008),
    .D(_01283_),
    .Q_N(_06028_),
    .Q(\mem.mem[148][4] ));
 sg13g2_dfrbp_1 _15837_ (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2007),
    .D(_01284_),
    .Q_N(_06027_),
    .Q(\mem.mem[148][5] ));
 sg13g2_dfrbp_1 _15838_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2006),
    .D(_01285_),
    .Q_N(_06026_),
    .Q(\mem.mem[148][6] ));
 sg13g2_dfrbp_1 _15839_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2005),
    .D(_01286_),
    .Q_N(_06025_),
    .Q(\mem.mem[148][7] ));
 sg13g2_dfrbp_1 _15840_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2004),
    .D(_01287_),
    .Q_N(_06024_),
    .Q(\mem.mem[14][0] ));
 sg13g2_dfrbp_1 _15841_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2003),
    .D(_01288_),
    .Q_N(_06023_),
    .Q(\mem.mem[14][1] ));
 sg13g2_dfrbp_1 _15842_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2002),
    .D(_01289_),
    .Q_N(_06022_),
    .Q(\mem.mem[14][2] ));
 sg13g2_dfrbp_1 _15843_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net2001),
    .D(_01290_),
    .Q_N(_06021_),
    .Q(\mem.mem[14][3] ));
 sg13g2_dfrbp_1 _15844_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2000),
    .D(_01291_),
    .Q_N(_06020_),
    .Q(\mem.mem[14][4] ));
 sg13g2_dfrbp_1 _15845_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1999),
    .D(_01292_),
    .Q_N(_06019_),
    .Q(\mem.mem[14][5] ));
 sg13g2_dfrbp_1 _15846_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1998),
    .D(_01293_),
    .Q_N(_06018_),
    .Q(\mem.mem[14][6] ));
 sg13g2_dfrbp_1 _15847_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1997),
    .D(_01294_),
    .Q_N(_06017_),
    .Q(\mem.mem[14][7] ));
 sg13g2_dfrbp_1 _15848_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1996),
    .D(_01295_),
    .Q_N(_06016_),
    .Q(\mem.mem[150][0] ));
 sg13g2_dfrbp_1 _15849_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1995),
    .D(_01296_),
    .Q_N(_06015_),
    .Q(\mem.mem[150][1] ));
 sg13g2_dfrbp_1 _15850_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1994),
    .D(_01297_),
    .Q_N(_06014_),
    .Q(\mem.mem[150][2] ));
 sg13g2_dfrbp_1 _15851_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1993),
    .D(_01298_),
    .Q_N(_06013_),
    .Q(\mem.mem[150][3] ));
 sg13g2_dfrbp_1 _15852_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1992),
    .D(_01299_),
    .Q_N(_06012_),
    .Q(\mem.mem[150][4] ));
 sg13g2_dfrbp_1 _15853_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1991),
    .D(_01300_),
    .Q_N(_06011_),
    .Q(\mem.mem[150][5] ));
 sg13g2_dfrbp_1 _15854_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1990),
    .D(_01301_),
    .Q_N(_06010_),
    .Q(\mem.mem[150][6] ));
 sg13g2_dfrbp_1 _15855_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1989),
    .D(_01302_),
    .Q_N(_06009_),
    .Q(\mem.mem[150][7] ));
 sg13g2_dfrbp_1 _15856_ (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1988),
    .D(_01303_),
    .Q_N(_06008_),
    .Q(\mem.mem[151][0] ));
 sg13g2_dfrbp_1 _15857_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1987),
    .D(_01304_),
    .Q_N(_06007_),
    .Q(\mem.mem[151][1] ));
 sg13g2_dfrbp_1 _15858_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1986),
    .D(_01305_),
    .Q_N(_06006_),
    .Q(\mem.mem[151][2] ));
 sg13g2_dfrbp_1 _15859_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1985),
    .D(_01306_),
    .Q_N(_06005_),
    .Q(\mem.mem[151][3] ));
 sg13g2_dfrbp_1 _15860_ (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1984),
    .D(_01307_),
    .Q_N(_06004_),
    .Q(\mem.mem[151][4] ));
 sg13g2_dfrbp_1 _15861_ (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1983),
    .D(_01308_),
    .Q_N(_06003_),
    .Q(\mem.mem[151][5] ));
 sg13g2_dfrbp_1 _15862_ (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1982),
    .D(_01309_),
    .Q_N(_06002_),
    .Q(\mem.mem[151][6] ));
 sg13g2_dfrbp_1 _15863_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1981),
    .D(_01310_),
    .Q_N(_06001_),
    .Q(\mem.mem[151][7] ));
 sg13g2_dfrbp_1 _15864_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1980),
    .D(_01311_),
    .Q_N(_06000_),
    .Q(\mem.mem[152][0] ));
 sg13g2_dfrbp_1 _15865_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1979),
    .D(_01312_),
    .Q_N(_05999_),
    .Q(\mem.mem[152][1] ));
 sg13g2_dfrbp_1 _15866_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1978),
    .D(_01313_),
    .Q_N(_05998_),
    .Q(\mem.mem[152][2] ));
 sg13g2_dfrbp_1 _15867_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1977),
    .D(_01314_),
    .Q_N(_05997_),
    .Q(\mem.mem[152][3] ));
 sg13g2_dfrbp_1 _15868_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1976),
    .D(_01315_),
    .Q_N(_05996_),
    .Q(\mem.mem[152][4] ));
 sg13g2_dfrbp_1 _15869_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1975),
    .D(_01316_),
    .Q_N(_05995_),
    .Q(\mem.mem[152][5] ));
 sg13g2_dfrbp_1 _15870_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1974),
    .D(_01317_),
    .Q_N(_05994_),
    .Q(\mem.mem[152][6] ));
 sg13g2_dfrbp_1 _15871_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1973),
    .D(_01318_),
    .Q_N(_05993_),
    .Q(\mem.mem[152][7] ));
 sg13g2_dfrbp_1 _15872_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1972),
    .D(_01319_),
    .Q_N(_05992_),
    .Q(\mem.mem[153][0] ));
 sg13g2_dfrbp_1 _15873_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1971),
    .D(_01320_),
    .Q_N(_05991_),
    .Q(\mem.mem[153][1] ));
 sg13g2_dfrbp_1 _15874_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1970),
    .D(_01321_),
    .Q_N(_05990_),
    .Q(\mem.mem[153][2] ));
 sg13g2_dfrbp_1 _15875_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1969),
    .D(_01322_),
    .Q_N(_05989_),
    .Q(\mem.mem[153][3] ));
 sg13g2_dfrbp_1 _15876_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1968),
    .D(_01323_),
    .Q_N(_05988_),
    .Q(\mem.mem[153][4] ));
 sg13g2_dfrbp_1 _15877_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1967),
    .D(_01324_),
    .Q_N(_05987_),
    .Q(\mem.mem[153][5] ));
 sg13g2_dfrbp_1 _15878_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1966),
    .D(_01325_),
    .Q_N(_05986_),
    .Q(\mem.mem[153][6] ));
 sg13g2_dfrbp_1 _15879_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1965),
    .D(_01326_),
    .Q_N(_05985_),
    .Q(\mem.mem[153][7] ));
 sg13g2_dfrbp_1 _15880_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1964),
    .D(_01327_),
    .Q_N(_05984_),
    .Q(\mem.mem[154][0] ));
 sg13g2_dfrbp_1 _15881_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1963),
    .D(_01328_),
    .Q_N(_05983_),
    .Q(\mem.mem[154][1] ));
 sg13g2_dfrbp_1 _15882_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1962),
    .D(_01329_),
    .Q_N(_05982_),
    .Q(\mem.mem[154][2] ));
 sg13g2_dfrbp_1 _15883_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1961),
    .D(_01330_),
    .Q_N(_05981_),
    .Q(\mem.mem[154][3] ));
 sg13g2_dfrbp_1 _15884_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1960),
    .D(_01331_),
    .Q_N(_05980_),
    .Q(\mem.mem[154][4] ));
 sg13g2_dfrbp_1 _15885_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1959),
    .D(_01332_),
    .Q_N(_05979_),
    .Q(\mem.mem[154][5] ));
 sg13g2_dfrbp_1 _15886_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1958),
    .D(_01333_),
    .Q_N(_05978_),
    .Q(\mem.mem[154][6] ));
 sg13g2_dfrbp_1 _15887_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1957),
    .D(_01334_),
    .Q_N(_05977_),
    .Q(\mem.mem[154][7] ));
 sg13g2_dfrbp_1 _15888_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1956),
    .D(_01335_),
    .Q_N(_05976_),
    .Q(\mem.mem[155][0] ));
 sg13g2_dfrbp_1 _15889_ (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1955),
    .D(_01336_),
    .Q_N(_05975_),
    .Q(\mem.mem[155][1] ));
 sg13g2_dfrbp_1 _15890_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1954),
    .D(_01337_),
    .Q_N(_05974_),
    .Q(\mem.mem[155][2] ));
 sg13g2_dfrbp_1 _15891_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1953),
    .D(_01338_),
    .Q_N(_05973_),
    .Q(\mem.mem[155][3] ));
 sg13g2_dfrbp_1 _15892_ (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1952),
    .D(_01339_),
    .Q_N(_05972_),
    .Q(\mem.mem[155][4] ));
 sg13g2_dfrbp_1 _15893_ (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1951),
    .D(_01340_),
    .Q_N(_05971_),
    .Q(\mem.mem[155][5] ));
 sg13g2_dfrbp_1 _15894_ (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1950),
    .D(_01341_),
    .Q_N(_05970_),
    .Q(\mem.mem[155][6] ));
 sg13g2_dfrbp_1 _15895_ (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1949),
    .D(_01342_),
    .Q_N(_05969_),
    .Q(\mem.mem[155][7] ));
 sg13g2_dfrbp_1 _15896_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1948),
    .D(_01343_),
    .Q_N(_05968_),
    .Q(\mem.mem[156][0] ));
 sg13g2_dfrbp_1 _15897_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1947),
    .D(_01344_),
    .Q_N(_05967_),
    .Q(\mem.mem[156][1] ));
 sg13g2_dfrbp_1 _15898_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1946),
    .D(_01345_),
    .Q_N(_05966_),
    .Q(\mem.mem[156][2] ));
 sg13g2_dfrbp_1 _15899_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1945),
    .D(_01346_),
    .Q_N(_05965_),
    .Q(\mem.mem[156][3] ));
 sg13g2_dfrbp_1 _15900_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1944),
    .D(_01347_),
    .Q_N(_05964_),
    .Q(\mem.mem[156][4] ));
 sg13g2_dfrbp_1 _15901_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1943),
    .D(_01348_),
    .Q_N(_05963_),
    .Q(\mem.mem[156][5] ));
 sg13g2_dfrbp_1 _15902_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1942),
    .D(_01349_),
    .Q_N(_05962_),
    .Q(\mem.mem[156][6] ));
 sg13g2_dfrbp_1 _15903_ (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1941),
    .D(_01350_),
    .Q_N(_05961_),
    .Q(\mem.mem[156][7] ));
 sg13g2_dfrbp_1 _15904_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1940),
    .D(_01351_),
    .Q_N(_05960_),
    .Q(\mem.mem[157][0] ));
 sg13g2_dfrbp_1 _15905_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1939),
    .D(_01352_),
    .Q_N(_05959_),
    .Q(\mem.mem[157][1] ));
 sg13g2_dfrbp_1 _15906_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1938),
    .D(_01353_),
    .Q_N(_05958_),
    .Q(\mem.mem[157][2] ));
 sg13g2_dfrbp_1 _15907_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1937),
    .D(_01354_),
    .Q_N(_05957_),
    .Q(\mem.mem[157][3] ));
 sg13g2_dfrbp_1 _15908_ (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1936),
    .D(_01355_),
    .Q_N(_05956_),
    .Q(\mem.mem[157][4] ));
 sg13g2_dfrbp_1 _15909_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1935),
    .D(_01356_),
    .Q_N(_05955_),
    .Q(\mem.mem[157][5] ));
 sg13g2_dfrbp_1 _15910_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1934),
    .D(_01357_),
    .Q_N(_05954_),
    .Q(\mem.mem[157][6] ));
 sg13g2_dfrbp_1 _15911_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1933),
    .D(_01358_),
    .Q_N(_05953_),
    .Q(\mem.mem[157][7] ));
 sg13g2_dfrbp_1 _15912_ (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1932),
    .D(_01359_),
    .Q_N(_05952_),
    .Q(\mem.mem[158][0] ));
 sg13g2_dfrbp_1 _15913_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1931),
    .D(_01360_),
    .Q_N(_05951_),
    .Q(\mem.mem[158][1] ));
 sg13g2_dfrbp_1 _15914_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1930),
    .D(_01361_),
    .Q_N(_05950_),
    .Q(\mem.mem[158][2] ));
 sg13g2_dfrbp_1 _15915_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1929),
    .D(_01362_),
    .Q_N(_05949_),
    .Q(\mem.mem[158][3] ));
 sg13g2_dfrbp_1 _15916_ (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1928),
    .D(_01363_),
    .Q_N(_05948_),
    .Q(\mem.mem[158][4] ));
 sg13g2_dfrbp_1 _15917_ (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1927),
    .D(_01364_),
    .Q_N(_05947_),
    .Q(\mem.mem[158][5] ));
 sg13g2_dfrbp_1 _15918_ (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1926),
    .D(_01365_),
    .Q_N(_05946_),
    .Q(\mem.mem[158][6] ));
 sg13g2_dfrbp_1 _15919_ (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1925),
    .D(_01366_),
    .Q_N(_05945_),
    .Q(\mem.mem[158][7] ));
 sg13g2_dfrbp_1 _15920_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1924),
    .D(_01367_),
    .Q_N(_05944_),
    .Q(\mem.mem[15][0] ));
 sg13g2_dfrbp_1 _15921_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1923),
    .D(_01368_),
    .Q_N(_05943_),
    .Q(\mem.mem[15][1] ));
 sg13g2_dfrbp_1 _15922_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1922),
    .D(_01369_),
    .Q_N(_05942_),
    .Q(\mem.mem[15][2] ));
 sg13g2_dfrbp_1 _15923_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1921),
    .D(_01370_),
    .Q_N(_05941_),
    .Q(\mem.mem[15][3] ));
 sg13g2_dfrbp_1 _15924_ (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1920),
    .D(_01371_),
    .Q_N(_05940_),
    .Q(\mem.mem[15][4] ));
 sg13g2_dfrbp_1 _15925_ (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1919),
    .D(_01372_),
    .Q_N(_05939_),
    .Q(\mem.mem[15][5] ));
 sg13g2_dfrbp_1 _15926_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1918),
    .D(_01373_),
    .Q_N(_05938_),
    .Q(\mem.mem[15][6] ));
 sg13g2_dfrbp_1 _15927_ (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1917),
    .D(_01374_),
    .Q_N(_05937_),
    .Q(\mem.mem[15][7] ));
 sg13g2_dfrbp_1 _15928_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1916),
    .D(_01375_),
    .Q_N(_05936_),
    .Q(\mem.mem[160][0] ));
 sg13g2_dfrbp_1 _15929_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1915),
    .D(_01376_),
    .Q_N(_05935_),
    .Q(\mem.mem[160][1] ));
 sg13g2_dfrbp_1 _15930_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1914),
    .D(_01377_),
    .Q_N(_05934_),
    .Q(\mem.mem[160][2] ));
 sg13g2_dfrbp_1 _15931_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1913),
    .D(_01378_),
    .Q_N(_05933_),
    .Q(\mem.mem[160][3] ));
 sg13g2_dfrbp_1 _15932_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1912),
    .D(_01379_),
    .Q_N(_05932_),
    .Q(\mem.mem[160][4] ));
 sg13g2_dfrbp_1 _15933_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1911),
    .D(_01380_),
    .Q_N(_05931_),
    .Q(\mem.mem[160][5] ));
 sg13g2_dfrbp_1 _15934_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1910),
    .D(_01381_),
    .Q_N(_05930_),
    .Q(\mem.mem[160][6] ));
 sg13g2_dfrbp_1 _15935_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1909),
    .D(_01382_),
    .Q_N(_05929_),
    .Q(\mem.mem[160][7] ));
 sg13g2_dfrbp_1 _15936_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1908),
    .D(_01383_),
    .Q_N(_05928_),
    .Q(\mem.mem[161][0] ));
 sg13g2_dfrbp_1 _15937_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1907),
    .D(_01384_),
    .Q_N(_05927_),
    .Q(\mem.mem[161][1] ));
 sg13g2_dfrbp_1 _15938_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1906),
    .D(_01385_),
    .Q_N(_05926_),
    .Q(\mem.mem[161][2] ));
 sg13g2_dfrbp_1 _15939_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1905),
    .D(_01386_),
    .Q_N(_05925_),
    .Q(\mem.mem[161][3] ));
 sg13g2_dfrbp_1 _15940_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1904),
    .D(_01387_),
    .Q_N(_05924_),
    .Q(\mem.mem[161][4] ));
 sg13g2_dfrbp_1 _15941_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1903),
    .D(_01388_),
    .Q_N(_05923_),
    .Q(\mem.mem[161][5] ));
 sg13g2_dfrbp_1 _15942_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1902),
    .D(_01389_),
    .Q_N(_05922_),
    .Q(\mem.mem[161][6] ));
 sg13g2_dfrbp_1 _15943_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1901),
    .D(_01390_),
    .Q_N(_05921_),
    .Q(\mem.mem[161][7] ));
 sg13g2_dfrbp_1 _15944_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1900),
    .D(_01391_),
    .Q_N(_05920_),
    .Q(\mem.mem[162][0] ));
 sg13g2_dfrbp_1 _15945_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1899),
    .D(_01392_),
    .Q_N(_05919_),
    .Q(\mem.mem[162][1] ));
 sg13g2_dfrbp_1 _15946_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1898),
    .D(_01393_),
    .Q_N(_05918_),
    .Q(\mem.mem[162][2] ));
 sg13g2_dfrbp_1 _15947_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1897),
    .D(_01394_),
    .Q_N(_05917_),
    .Q(\mem.mem[162][3] ));
 sg13g2_dfrbp_1 _15948_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1896),
    .D(_01395_),
    .Q_N(_05916_),
    .Q(\mem.mem[162][4] ));
 sg13g2_dfrbp_1 _15949_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1895),
    .D(_01396_),
    .Q_N(_05915_),
    .Q(\mem.mem[162][5] ));
 sg13g2_dfrbp_1 _15950_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1894),
    .D(_01397_),
    .Q_N(_05914_),
    .Q(\mem.mem[162][6] ));
 sg13g2_dfrbp_1 _15951_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1893),
    .D(_01398_),
    .Q_N(_05913_),
    .Q(\mem.mem[162][7] ));
 sg13g2_dfrbp_1 _15952_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1892),
    .D(_01399_),
    .Q_N(_05912_),
    .Q(\mem.mem[163][0] ));
 sg13g2_dfrbp_1 _15953_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1891),
    .D(_01400_),
    .Q_N(_05911_),
    .Q(\mem.mem[163][1] ));
 sg13g2_dfrbp_1 _15954_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1890),
    .D(_01401_),
    .Q_N(_05910_),
    .Q(\mem.mem[163][2] ));
 sg13g2_dfrbp_1 _15955_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1889),
    .D(_01402_),
    .Q_N(_05909_),
    .Q(\mem.mem[163][3] ));
 sg13g2_dfrbp_1 _15956_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1888),
    .D(_01403_),
    .Q_N(_05908_),
    .Q(\mem.mem[163][4] ));
 sg13g2_dfrbp_1 _15957_ (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1887),
    .D(_01404_),
    .Q_N(_05907_),
    .Q(\mem.mem[163][5] ));
 sg13g2_dfrbp_1 _15958_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1886),
    .D(_01405_),
    .Q_N(_05906_),
    .Q(\mem.mem[163][6] ));
 sg13g2_dfrbp_1 _15959_ (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1885),
    .D(_01406_),
    .Q_N(_05905_),
    .Q(\mem.mem[163][7] ));
 sg13g2_dfrbp_1 _15960_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1884),
    .D(_01407_),
    .Q_N(_05904_),
    .Q(\mem.mem[164][0] ));
 sg13g2_dfrbp_1 _15961_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1883),
    .D(_01408_),
    .Q_N(_05903_),
    .Q(\mem.mem[164][1] ));
 sg13g2_dfrbp_1 _15962_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1882),
    .D(_01409_),
    .Q_N(_05902_),
    .Q(\mem.mem[164][2] ));
 sg13g2_dfrbp_1 _15963_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1881),
    .D(_01410_),
    .Q_N(_05901_),
    .Q(\mem.mem[164][3] ));
 sg13g2_dfrbp_1 _15964_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1880),
    .D(_01411_),
    .Q_N(_05900_),
    .Q(\mem.mem[164][4] ));
 sg13g2_dfrbp_1 _15965_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1879),
    .D(_01412_),
    .Q_N(_05899_),
    .Q(\mem.mem[164][5] ));
 sg13g2_dfrbp_1 _15966_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1878),
    .D(_01413_),
    .Q_N(_05898_),
    .Q(\mem.mem[164][6] ));
 sg13g2_dfrbp_1 _15967_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1877),
    .D(_01414_),
    .Q_N(_05897_),
    .Q(\mem.mem[164][7] ));
 sg13g2_dfrbp_1 _15968_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1876),
    .D(_01415_),
    .Q_N(_05896_),
    .Q(\mem.mem[165][0] ));
 sg13g2_dfrbp_1 _15969_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1875),
    .D(_01416_),
    .Q_N(_05895_),
    .Q(\mem.mem[165][1] ));
 sg13g2_dfrbp_1 _15970_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1874),
    .D(_01417_),
    .Q_N(_05894_),
    .Q(\mem.mem[165][2] ));
 sg13g2_dfrbp_1 _15971_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1873),
    .D(_01418_),
    .Q_N(_05893_),
    .Q(\mem.mem[165][3] ));
 sg13g2_dfrbp_1 _15972_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1872),
    .D(_01419_),
    .Q_N(_05892_),
    .Q(\mem.mem[165][4] ));
 sg13g2_dfrbp_1 _15973_ (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1871),
    .D(_01420_),
    .Q_N(_05891_),
    .Q(\mem.mem[165][5] ));
 sg13g2_dfrbp_1 _15974_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1870),
    .D(_01421_),
    .Q_N(_05890_),
    .Q(\mem.mem[165][6] ));
 sg13g2_dfrbp_1 _15975_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1869),
    .D(_01422_),
    .Q_N(_05889_),
    .Q(\mem.mem[165][7] ));
 sg13g2_dfrbp_1 _15976_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1868),
    .D(_01423_),
    .Q_N(_05888_),
    .Q(\mem.mem[166][0] ));
 sg13g2_dfrbp_1 _15977_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1867),
    .D(_01424_),
    .Q_N(_05887_),
    .Q(\mem.mem[166][1] ));
 sg13g2_dfrbp_1 _15978_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1866),
    .D(_01425_),
    .Q_N(_05886_),
    .Q(\mem.mem[166][2] ));
 sg13g2_dfrbp_1 _15979_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1865),
    .D(_01426_),
    .Q_N(_05885_),
    .Q(\mem.mem[166][3] ));
 sg13g2_dfrbp_1 _15980_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1864),
    .D(_01427_),
    .Q_N(_05884_),
    .Q(\mem.mem[166][4] ));
 sg13g2_dfrbp_1 _15981_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1863),
    .D(_01428_),
    .Q_N(_05883_),
    .Q(\mem.mem[166][5] ));
 sg13g2_dfrbp_1 _15982_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1862),
    .D(_01429_),
    .Q_N(_05882_),
    .Q(\mem.mem[166][6] ));
 sg13g2_dfrbp_1 _15983_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1861),
    .D(_01430_),
    .Q_N(_05881_),
    .Q(\mem.mem[166][7] ));
 sg13g2_dfrbp_1 _15984_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1860),
    .D(_01431_),
    .Q_N(_05880_),
    .Q(\mem.mem[167][0] ));
 sg13g2_dfrbp_1 _15985_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1859),
    .D(_01432_),
    .Q_N(_05879_),
    .Q(\mem.mem[167][1] ));
 sg13g2_dfrbp_1 _15986_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1858),
    .D(_01433_),
    .Q_N(_05878_),
    .Q(\mem.mem[167][2] ));
 sg13g2_dfrbp_1 _15987_ (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1857),
    .D(_01434_),
    .Q_N(_05877_),
    .Q(\mem.mem[167][3] ));
 sg13g2_dfrbp_1 _15988_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1856),
    .D(_01435_),
    .Q_N(_05876_),
    .Q(\mem.mem[167][4] ));
 sg13g2_dfrbp_1 _15989_ (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1855),
    .D(_01436_),
    .Q_N(_05875_),
    .Q(\mem.mem[167][5] ));
 sg13g2_dfrbp_1 _15990_ (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1854),
    .D(_01437_),
    .Q_N(_05874_),
    .Q(\mem.mem[167][6] ));
 sg13g2_dfrbp_1 _15991_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1853),
    .D(_01438_),
    .Q_N(_05873_),
    .Q(\mem.mem[167][7] ));
 sg13g2_dfrbp_1 _15992_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1852),
    .D(_01439_),
    .Q_N(_05872_),
    .Q(\mem.mem[168][0] ));
 sg13g2_dfrbp_1 _15993_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1851),
    .D(_01440_),
    .Q_N(_05871_),
    .Q(\mem.mem[168][1] ));
 sg13g2_dfrbp_1 _15994_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1850),
    .D(_01441_),
    .Q_N(_05870_),
    .Q(\mem.mem[168][2] ));
 sg13g2_dfrbp_1 _15995_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1849),
    .D(_01442_),
    .Q_N(_05869_),
    .Q(\mem.mem[168][3] ));
 sg13g2_dfrbp_1 _15996_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1848),
    .D(_01443_),
    .Q_N(_05868_),
    .Q(\mem.mem[168][4] ));
 sg13g2_dfrbp_1 _15997_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1847),
    .D(_01444_),
    .Q_N(_05867_),
    .Q(\mem.mem[168][5] ));
 sg13g2_dfrbp_1 _15998_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1846),
    .D(_01445_),
    .Q_N(_05866_),
    .Q(\mem.mem[168][6] ));
 sg13g2_dfrbp_1 _15999_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1845),
    .D(_01446_),
    .Q_N(_05865_),
    .Q(\mem.mem[168][7] ));
 sg13g2_dfrbp_1 _16000_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1844),
    .D(_01447_),
    .Q_N(_05864_),
    .Q(\mem.mem[16][0] ));
 sg13g2_dfrbp_1 _16001_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1843),
    .D(_01448_),
    .Q_N(_05863_),
    .Q(\mem.mem[16][1] ));
 sg13g2_dfrbp_1 _16002_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1842),
    .D(_01449_),
    .Q_N(_05862_),
    .Q(\mem.mem[16][2] ));
 sg13g2_dfrbp_1 _16003_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1841),
    .D(_01450_),
    .Q_N(_05861_),
    .Q(\mem.mem[16][3] ));
 sg13g2_dfrbp_1 _16004_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1840),
    .D(_01451_),
    .Q_N(_05860_),
    .Q(\mem.mem[16][4] ));
 sg13g2_dfrbp_1 _16005_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1839),
    .D(_01452_),
    .Q_N(_05859_),
    .Q(\mem.mem[16][5] ));
 sg13g2_dfrbp_1 _16006_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1838),
    .D(_01453_),
    .Q_N(_05858_),
    .Q(\mem.mem[16][6] ));
 sg13g2_dfrbp_1 _16007_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1837),
    .D(_01454_),
    .Q_N(_05857_),
    .Q(\mem.mem[16][7] ));
 sg13g2_dfrbp_1 _16008_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1836),
    .D(_01455_),
    .Q_N(_05856_),
    .Q(\mem.mem[170][0] ));
 sg13g2_dfrbp_1 _16009_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1835),
    .D(_01456_),
    .Q_N(_05855_),
    .Q(\mem.mem[170][1] ));
 sg13g2_dfrbp_1 _16010_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1834),
    .D(_01457_),
    .Q_N(_05854_),
    .Q(\mem.mem[170][2] ));
 sg13g2_dfrbp_1 _16011_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1833),
    .D(_01458_),
    .Q_N(_05853_),
    .Q(\mem.mem[170][3] ));
 sg13g2_dfrbp_1 _16012_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1832),
    .D(_01459_),
    .Q_N(_05852_),
    .Q(\mem.mem[170][4] ));
 sg13g2_dfrbp_1 _16013_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1831),
    .D(_01460_),
    .Q_N(_05851_),
    .Q(\mem.mem[170][5] ));
 sg13g2_dfrbp_1 _16014_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1830),
    .D(_01461_),
    .Q_N(_05850_),
    .Q(\mem.mem[170][6] ));
 sg13g2_dfrbp_1 _16015_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1829),
    .D(_01462_),
    .Q_N(_05849_),
    .Q(\mem.mem[170][7] ));
 sg13g2_dfrbp_1 _16016_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1828),
    .D(_01463_),
    .Q_N(_05848_),
    .Q(\mem.mem[171][0] ));
 sg13g2_dfrbp_1 _16017_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1827),
    .D(_01464_),
    .Q_N(_05847_),
    .Q(\mem.mem[171][1] ));
 sg13g2_dfrbp_1 _16018_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1826),
    .D(_01465_),
    .Q_N(_05846_),
    .Q(\mem.mem[171][2] ));
 sg13g2_dfrbp_1 _16019_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1825),
    .D(_01466_),
    .Q_N(_05845_),
    .Q(\mem.mem[171][3] ));
 sg13g2_dfrbp_1 _16020_ (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1824),
    .D(_01467_),
    .Q_N(_05844_),
    .Q(\mem.mem[171][4] ));
 sg13g2_dfrbp_1 _16021_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1823),
    .D(_01468_),
    .Q_N(_05843_),
    .Q(\mem.mem[171][5] ));
 sg13g2_dfrbp_1 _16022_ (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1822),
    .D(_01469_),
    .Q_N(_05842_),
    .Q(\mem.mem[171][6] ));
 sg13g2_dfrbp_1 _16023_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1821),
    .D(_01470_),
    .Q_N(_05841_),
    .Q(\mem.mem[171][7] ));
 sg13g2_dfrbp_1 _16024_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1820),
    .D(_01471_),
    .Q_N(_05840_),
    .Q(\mem.mem[172][0] ));
 sg13g2_dfrbp_1 _16025_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1819),
    .D(_01472_),
    .Q_N(_05839_),
    .Q(\mem.mem[172][1] ));
 sg13g2_dfrbp_1 _16026_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1818),
    .D(net2861),
    .Q_N(_05838_),
    .Q(\mem.mem[172][2] ));
 sg13g2_dfrbp_1 _16027_ (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1817),
    .D(_01474_),
    .Q_N(_05837_),
    .Q(\mem.mem[172][3] ));
 sg13g2_dfrbp_1 _16028_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1816),
    .D(_01475_),
    .Q_N(_05836_),
    .Q(\mem.mem[172][4] ));
 sg13g2_dfrbp_1 _16029_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1815),
    .D(_01476_),
    .Q_N(_05835_),
    .Q(\mem.mem[172][5] ));
 sg13g2_dfrbp_1 _16030_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1814),
    .D(_01477_),
    .Q_N(_05834_),
    .Q(\mem.mem[172][6] ));
 sg13g2_dfrbp_1 _16031_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1813),
    .D(_01478_),
    .Q_N(_05833_),
    .Q(\mem.mem[172][7] ));
 sg13g2_dfrbp_1 _16032_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1812),
    .D(_01479_),
    .Q_N(_05832_),
    .Q(\mem.mem[173][0] ));
 sg13g2_dfrbp_1 _16033_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1811),
    .D(_01480_),
    .Q_N(_05831_),
    .Q(\mem.mem[173][1] ));
 sg13g2_dfrbp_1 _16034_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1810),
    .D(_01481_),
    .Q_N(_05830_),
    .Q(\mem.mem[173][2] ));
 sg13g2_dfrbp_1 _16035_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1809),
    .D(_01482_),
    .Q_N(_05829_),
    .Q(\mem.mem[173][3] ));
 sg13g2_dfrbp_1 _16036_ (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1808),
    .D(_01483_),
    .Q_N(_05828_),
    .Q(\mem.mem[173][4] ));
 sg13g2_dfrbp_1 _16037_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1807),
    .D(_01484_),
    .Q_N(_05827_),
    .Q(\mem.mem[173][5] ));
 sg13g2_dfrbp_1 _16038_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1806),
    .D(_01485_),
    .Q_N(_05826_),
    .Q(\mem.mem[173][6] ));
 sg13g2_dfrbp_1 _16039_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1805),
    .D(_01486_),
    .Q_N(_05825_),
    .Q(\mem.mem[173][7] ));
 sg13g2_dfrbp_1 _16040_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1804),
    .D(_01487_),
    .Q_N(_05824_),
    .Q(\mem.mem[174][0] ));
 sg13g2_dfrbp_1 _16041_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1803),
    .D(_01488_),
    .Q_N(_05823_),
    .Q(\mem.mem[174][1] ));
 sg13g2_dfrbp_1 _16042_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1802),
    .D(_01489_),
    .Q_N(_05822_),
    .Q(\mem.mem[174][2] ));
 sg13g2_dfrbp_1 _16043_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1801),
    .D(_01490_),
    .Q_N(_05821_),
    .Q(\mem.mem[174][3] ));
 sg13g2_dfrbp_1 _16044_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1800),
    .D(_01491_),
    .Q_N(_05820_),
    .Q(\mem.mem[174][4] ));
 sg13g2_dfrbp_1 _16045_ (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1799),
    .D(_01492_),
    .Q_N(_05819_),
    .Q(\mem.mem[174][5] ));
 sg13g2_dfrbp_1 _16046_ (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1798),
    .D(_01493_),
    .Q_N(_05818_),
    .Q(\mem.mem[174][6] ));
 sg13g2_dfrbp_1 _16047_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1797),
    .D(_01494_),
    .Q_N(_05817_),
    .Q(\mem.mem[174][7] ));
 sg13g2_dfrbp_1 _16048_ (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1796),
    .D(_01495_),
    .Q_N(_05816_),
    .Q(\mem.mem[175][0] ));
 sg13g2_dfrbp_1 _16049_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1795),
    .D(_01496_),
    .Q_N(_05815_),
    .Q(\mem.mem[175][1] ));
 sg13g2_dfrbp_1 _16050_ (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1794),
    .D(_01497_),
    .Q_N(_05814_),
    .Q(\mem.mem[175][2] ));
 sg13g2_dfrbp_1 _16051_ (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1793),
    .D(_01498_),
    .Q_N(_05813_),
    .Q(\mem.mem[175][3] ));
 sg13g2_dfrbp_1 _16052_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1792),
    .D(_01499_),
    .Q_N(_05812_),
    .Q(\mem.mem[175][4] ));
 sg13g2_dfrbp_1 _16053_ (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1791),
    .D(_01500_),
    .Q_N(_05811_),
    .Q(\mem.mem[175][5] ));
 sg13g2_dfrbp_1 _16054_ (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1790),
    .D(_01501_),
    .Q_N(_05810_),
    .Q(\mem.mem[175][6] ));
 sg13g2_dfrbp_1 _16055_ (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1789),
    .D(_01502_),
    .Q_N(_05809_),
    .Q(\mem.mem[175][7] ));
 sg13g2_dfrbp_1 _16056_ (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1788),
    .D(_01503_),
    .Q_N(_05808_),
    .Q(\mem.mem[176][0] ));
 sg13g2_dfrbp_1 _16057_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1787),
    .D(_01504_),
    .Q_N(_05807_),
    .Q(\mem.mem[176][1] ));
 sg13g2_dfrbp_1 _16058_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1786),
    .D(_01505_),
    .Q_N(_05806_),
    .Q(\mem.mem[176][2] ));
 sg13g2_dfrbp_1 _16059_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1785),
    .D(_01506_),
    .Q_N(_05805_),
    .Q(\mem.mem[176][3] ));
 sg13g2_dfrbp_1 _16060_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1784),
    .D(_01507_),
    .Q_N(_05804_),
    .Q(\mem.mem[176][4] ));
 sg13g2_dfrbp_1 _16061_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1783),
    .D(_01508_),
    .Q_N(_05803_),
    .Q(\mem.mem[176][5] ));
 sg13g2_dfrbp_1 _16062_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1782),
    .D(_01509_),
    .Q_N(_05802_),
    .Q(\mem.mem[176][6] ));
 sg13g2_dfrbp_1 _16063_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1781),
    .D(_01510_),
    .Q_N(_05801_),
    .Q(\mem.mem[176][7] ));
 sg13g2_dfrbp_1 _16064_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1780),
    .D(_01511_),
    .Q_N(_05800_),
    .Q(\mem.mem[177][0] ));
 sg13g2_dfrbp_1 _16065_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1779),
    .D(_01512_),
    .Q_N(_05799_),
    .Q(\mem.mem[177][1] ));
 sg13g2_dfrbp_1 _16066_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1778),
    .D(_01513_),
    .Q_N(_05798_),
    .Q(\mem.mem[177][2] ));
 sg13g2_dfrbp_1 _16067_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1777),
    .D(_01514_),
    .Q_N(_05797_),
    .Q(\mem.mem[177][3] ));
 sg13g2_dfrbp_1 _16068_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1776),
    .D(_01515_),
    .Q_N(_05796_),
    .Q(\mem.mem[177][4] ));
 sg13g2_dfrbp_1 _16069_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1775),
    .D(_01516_),
    .Q_N(_05795_),
    .Q(\mem.mem[177][5] ));
 sg13g2_dfrbp_1 _16070_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1774),
    .D(_01517_),
    .Q_N(_05794_),
    .Q(\mem.mem[177][6] ));
 sg13g2_dfrbp_1 _16071_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1773),
    .D(_01518_),
    .Q_N(_05793_),
    .Q(\mem.mem[177][7] ));
 sg13g2_dfrbp_1 _16072_ (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1772),
    .D(_01519_),
    .Q_N(_05792_),
    .Q(\mem.mem[178][0] ));
 sg13g2_dfrbp_1 _16073_ (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1771),
    .D(_01520_),
    .Q_N(_05791_),
    .Q(\mem.mem[178][1] ));
 sg13g2_dfrbp_1 _16074_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1770),
    .D(_01521_),
    .Q_N(_05790_),
    .Q(\mem.mem[178][2] ));
 sg13g2_dfrbp_1 _16075_ (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1769),
    .D(_01522_),
    .Q_N(_05789_),
    .Q(\mem.mem[178][3] ));
 sg13g2_dfrbp_1 _16076_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1768),
    .D(_01523_),
    .Q_N(_05788_),
    .Q(\mem.mem[178][4] ));
 sg13g2_dfrbp_1 _16077_ (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1767),
    .D(_01524_),
    .Q_N(_05787_),
    .Q(\mem.mem[178][5] ));
 sg13g2_dfrbp_1 _16078_ (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1766),
    .D(_01525_),
    .Q_N(_05786_),
    .Q(\mem.mem[178][6] ));
 sg13g2_dfrbp_1 _16079_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1765),
    .D(_01526_),
    .Q_N(_05785_),
    .Q(\mem.mem[178][7] ));
 sg13g2_dfrbp_1 _16080_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1764),
    .D(_01527_),
    .Q_N(_05784_),
    .Q(\mem.mem[17][0] ));
 sg13g2_dfrbp_1 _16081_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1763),
    .D(_01528_),
    .Q_N(_05783_),
    .Q(\mem.mem[17][1] ));
 sg13g2_dfrbp_1 _16082_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1762),
    .D(_01529_),
    .Q_N(_05782_),
    .Q(\mem.mem[17][2] ));
 sg13g2_dfrbp_1 _16083_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1761),
    .D(_01530_),
    .Q_N(_05781_),
    .Q(\mem.mem[17][3] ));
 sg13g2_dfrbp_1 _16084_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1760),
    .D(_01531_),
    .Q_N(_05780_),
    .Q(\mem.mem[17][4] ));
 sg13g2_dfrbp_1 _16085_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1759),
    .D(_01532_),
    .Q_N(_05779_),
    .Q(\mem.mem[17][5] ));
 sg13g2_dfrbp_1 _16086_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1758),
    .D(_01533_),
    .Q_N(_05778_),
    .Q(\mem.mem[17][6] ));
 sg13g2_dfrbp_1 _16087_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1757),
    .D(_01534_),
    .Q_N(_05777_),
    .Q(\mem.mem[17][7] ));
 sg13g2_dfrbp_1 _16088_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1756),
    .D(_01535_),
    .Q_N(_05776_),
    .Q(\mem.mem[180][0] ));
 sg13g2_dfrbp_1 _16089_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1755),
    .D(_01536_),
    .Q_N(_05775_),
    .Q(\mem.mem[180][1] ));
 sg13g2_dfrbp_1 _16090_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1754),
    .D(_01537_),
    .Q_N(_05774_),
    .Q(\mem.mem[180][2] ));
 sg13g2_dfrbp_1 _16091_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1753),
    .D(_01538_),
    .Q_N(_05773_),
    .Q(\mem.mem[180][3] ));
 sg13g2_dfrbp_1 _16092_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1752),
    .D(_01539_),
    .Q_N(_05772_),
    .Q(\mem.mem[180][4] ));
 sg13g2_dfrbp_1 _16093_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1751),
    .D(_01540_),
    .Q_N(_05771_),
    .Q(\mem.mem[180][5] ));
 sg13g2_dfrbp_1 _16094_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1750),
    .D(_01541_),
    .Q_N(_05770_),
    .Q(\mem.mem[180][6] ));
 sg13g2_dfrbp_1 _16095_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1749),
    .D(_01542_),
    .Q_N(_05769_),
    .Q(\mem.mem[180][7] ));
 sg13g2_dfrbp_1 _16096_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1748),
    .D(_01543_),
    .Q_N(_05768_),
    .Q(\mem.mem[181][0] ));
 sg13g2_dfrbp_1 _16097_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1747),
    .D(_01544_),
    .Q_N(_05767_),
    .Q(\mem.mem[181][1] ));
 sg13g2_dfrbp_1 _16098_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1746),
    .D(_01545_),
    .Q_N(_05766_),
    .Q(\mem.mem[181][2] ));
 sg13g2_dfrbp_1 _16099_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1745),
    .D(_01546_),
    .Q_N(_05765_),
    .Q(\mem.mem[181][3] ));
 sg13g2_dfrbp_1 _16100_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1744),
    .D(_01547_),
    .Q_N(_05764_),
    .Q(\mem.mem[181][4] ));
 sg13g2_dfrbp_1 _16101_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1743),
    .D(_01548_),
    .Q_N(_05763_),
    .Q(\mem.mem[181][5] ));
 sg13g2_dfrbp_1 _16102_ (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1742),
    .D(_01549_),
    .Q_N(_05762_),
    .Q(\mem.mem[181][6] ));
 sg13g2_dfrbp_1 _16103_ (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1741),
    .D(_01550_),
    .Q_N(_05761_),
    .Q(\mem.mem[181][7] ));
 sg13g2_dfrbp_1 _16104_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1740),
    .D(_01551_),
    .Q_N(_05760_),
    .Q(\mem.mem[182][0] ));
 sg13g2_dfrbp_1 _16105_ (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1739),
    .D(_01552_),
    .Q_N(_05759_),
    .Q(\mem.mem[182][1] ));
 sg13g2_dfrbp_1 _16106_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1738),
    .D(_01553_),
    .Q_N(_05758_),
    .Q(\mem.mem[182][2] ));
 sg13g2_dfrbp_1 _16107_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1737),
    .D(_01554_),
    .Q_N(_05757_),
    .Q(\mem.mem[182][3] ));
 sg13g2_dfrbp_1 _16108_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1736),
    .D(_01555_),
    .Q_N(_05756_),
    .Q(\mem.mem[182][4] ));
 sg13g2_dfrbp_1 _16109_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1735),
    .D(_01556_),
    .Q_N(_05755_),
    .Q(\mem.mem[182][5] ));
 sg13g2_dfrbp_1 _16110_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1734),
    .D(_01557_),
    .Q_N(_05754_),
    .Q(\mem.mem[182][6] ));
 sg13g2_dfrbp_1 _16111_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1733),
    .D(_01558_),
    .Q_N(_05753_),
    .Q(\mem.mem[182][7] ));
 sg13g2_dfrbp_1 _16112_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1732),
    .D(_01559_),
    .Q_N(_05752_),
    .Q(\mem.mem[183][0] ));
 sg13g2_dfrbp_1 _16113_ (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1731),
    .D(_01560_),
    .Q_N(_05751_),
    .Q(\mem.mem[183][1] ));
 sg13g2_dfrbp_1 _16114_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1730),
    .D(_01561_),
    .Q_N(_05750_),
    .Q(\mem.mem[183][2] ));
 sg13g2_dfrbp_1 _16115_ (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1729),
    .D(_01562_),
    .Q_N(_05749_),
    .Q(\mem.mem[183][3] ));
 sg13g2_dfrbp_1 _16116_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1728),
    .D(_01563_),
    .Q_N(_05748_),
    .Q(\mem.mem[183][4] ));
 sg13g2_dfrbp_1 _16117_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1727),
    .D(_01564_),
    .Q_N(_05747_),
    .Q(\mem.mem[183][5] ));
 sg13g2_dfrbp_1 _16118_ (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1726),
    .D(_01565_),
    .Q_N(_05746_),
    .Q(\mem.mem[183][6] ));
 sg13g2_dfrbp_1 _16119_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1725),
    .D(_01566_),
    .Q_N(_05745_),
    .Q(\mem.mem[183][7] ));
 sg13g2_dfrbp_1 _16120_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1724),
    .D(_01567_),
    .Q_N(_05744_),
    .Q(\mem.mem[184][0] ));
 sg13g2_dfrbp_1 _16121_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1723),
    .D(_01568_),
    .Q_N(_05743_),
    .Q(\mem.mem[184][1] ));
 sg13g2_dfrbp_1 _16122_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1722),
    .D(_01569_),
    .Q_N(_05742_),
    .Q(\mem.mem[184][2] ));
 sg13g2_dfrbp_1 _16123_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1721),
    .D(_01570_),
    .Q_N(_05741_),
    .Q(\mem.mem[184][3] ));
 sg13g2_dfrbp_1 _16124_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1720),
    .D(_01571_),
    .Q_N(_05740_),
    .Q(\mem.mem[184][4] ));
 sg13g2_dfrbp_1 _16125_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1719),
    .D(_01572_),
    .Q_N(_05739_),
    .Q(\mem.mem[184][5] ));
 sg13g2_dfrbp_1 _16126_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1718),
    .D(_01573_),
    .Q_N(_05738_),
    .Q(\mem.mem[184][6] ));
 sg13g2_dfrbp_1 _16127_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1717),
    .D(_01574_),
    .Q_N(_05737_),
    .Q(\mem.mem[184][7] ));
 sg13g2_dfrbp_1 _16128_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1716),
    .D(_01575_),
    .Q_N(_05736_),
    .Q(\mem.mem[185][0] ));
 sg13g2_dfrbp_1 _16129_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1715),
    .D(_01576_),
    .Q_N(_05735_),
    .Q(\mem.mem[185][1] ));
 sg13g2_dfrbp_1 _16130_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1714),
    .D(_01577_),
    .Q_N(_05734_),
    .Q(\mem.mem[185][2] ));
 sg13g2_dfrbp_1 _16131_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1713),
    .D(_01578_),
    .Q_N(_05733_),
    .Q(\mem.mem[185][3] ));
 sg13g2_dfrbp_1 _16132_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1712),
    .D(_01579_),
    .Q_N(_05732_),
    .Q(\mem.mem[185][4] ));
 sg13g2_dfrbp_1 _16133_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1711),
    .D(_01580_),
    .Q_N(_05731_),
    .Q(\mem.mem[185][5] ));
 sg13g2_dfrbp_1 _16134_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1710),
    .D(_01581_),
    .Q_N(_05730_),
    .Q(\mem.mem[185][6] ));
 sg13g2_dfrbp_1 _16135_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1709),
    .D(_01582_),
    .Q_N(_05729_),
    .Q(\mem.mem[185][7] ));
 sg13g2_dfrbp_1 _16136_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1708),
    .D(_01583_),
    .Q_N(_05728_),
    .Q(\mem.mem[186][0] ));
 sg13g2_dfrbp_1 _16137_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1707),
    .D(_01584_),
    .Q_N(_05727_),
    .Q(\mem.mem[186][1] ));
 sg13g2_dfrbp_1 _16138_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1706),
    .D(_01585_),
    .Q_N(_05726_),
    .Q(\mem.mem[186][2] ));
 sg13g2_dfrbp_1 _16139_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1705),
    .D(_01586_),
    .Q_N(_05725_),
    .Q(\mem.mem[186][3] ));
 sg13g2_dfrbp_1 _16140_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1704),
    .D(_01587_),
    .Q_N(_05724_),
    .Q(\mem.mem[186][4] ));
 sg13g2_dfrbp_1 _16141_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1703),
    .D(_01588_),
    .Q_N(_05723_),
    .Q(\mem.mem[186][5] ));
 sg13g2_dfrbp_1 _16142_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1702),
    .D(_01589_),
    .Q_N(_05722_),
    .Q(\mem.mem[186][6] ));
 sg13g2_dfrbp_1 _16143_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1701),
    .D(_01590_),
    .Q_N(_05721_),
    .Q(\mem.mem[186][7] ));
 sg13g2_dfrbp_1 _16144_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1700),
    .D(_01591_),
    .Q_N(_05720_),
    .Q(\mem.mem[187][0] ));
 sg13g2_dfrbp_1 _16145_ (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1699),
    .D(_01592_),
    .Q_N(_05719_),
    .Q(\mem.mem[187][1] ));
 sg13g2_dfrbp_1 _16146_ (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1698),
    .D(_01593_),
    .Q_N(_05718_),
    .Q(\mem.mem[187][2] ));
 sg13g2_dfrbp_1 _16147_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1697),
    .D(_01594_),
    .Q_N(_05717_),
    .Q(\mem.mem[187][3] ));
 sg13g2_dfrbp_1 _16148_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1696),
    .D(_01595_),
    .Q_N(_05716_),
    .Q(\mem.mem[187][4] ));
 sg13g2_dfrbp_1 _16149_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1695),
    .D(_01596_),
    .Q_N(_05715_),
    .Q(\mem.mem[187][5] ));
 sg13g2_dfrbp_1 _16150_ (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1694),
    .D(_01597_),
    .Q_N(_05714_),
    .Q(\mem.mem[187][6] ));
 sg13g2_dfrbp_1 _16151_ (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1693),
    .D(_01598_),
    .Q_N(_05713_),
    .Q(\mem.mem[187][7] ));
 sg13g2_dfrbp_1 _16152_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1692),
    .D(_01599_),
    .Q_N(_05712_),
    .Q(\mem.mem[188][0] ));
 sg13g2_dfrbp_1 _16153_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1691),
    .D(_01600_),
    .Q_N(_05711_),
    .Q(\mem.mem[188][1] ));
 sg13g2_dfrbp_1 _16154_ (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1690),
    .D(_01601_),
    .Q_N(_05710_),
    .Q(\mem.mem[188][2] ));
 sg13g2_dfrbp_1 _16155_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1689),
    .D(_01602_),
    .Q_N(_05709_),
    .Q(\mem.mem[188][3] ));
 sg13g2_dfrbp_1 _16156_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1688),
    .D(_01603_),
    .Q_N(_05708_),
    .Q(\mem.mem[188][4] ));
 sg13g2_dfrbp_1 _16157_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1687),
    .D(_01604_),
    .Q_N(_05707_),
    .Q(\mem.mem[188][5] ));
 sg13g2_dfrbp_1 _16158_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1686),
    .D(_01605_),
    .Q_N(_05706_),
    .Q(\mem.mem[188][6] ));
 sg13g2_dfrbp_1 _16159_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1685),
    .D(_01606_),
    .Q_N(_05705_),
    .Q(\mem.mem[188][7] ));
 sg13g2_dfrbp_1 _16160_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1684),
    .D(_01607_),
    .Q_N(_05704_),
    .Q(\mem.mem[18][0] ));
 sg13g2_dfrbp_1 _16161_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1683),
    .D(_01608_),
    .Q_N(_05703_),
    .Q(\mem.mem[18][1] ));
 sg13g2_dfrbp_1 _16162_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1682),
    .D(_01609_),
    .Q_N(_05702_),
    .Q(\mem.mem[18][2] ));
 sg13g2_dfrbp_1 _16163_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1681),
    .D(_01610_),
    .Q_N(_05701_),
    .Q(\mem.mem[18][3] ));
 sg13g2_dfrbp_1 _16164_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1680),
    .D(_01611_),
    .Q_N(_05700_),
    .Q(\mem.mem[18][4] ));
 sg13g2_dfrbp_1 _16165_ (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1679),
    .D(_01612_),
    .Q_N(_05699_),
    .Q(\mem.mem[18][5] ));
 sg13g2_dfrbp_1 _16166_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1678),
    .D(_01613_),
    .Q_N(_05698_),
    .Q(\mem.mem[18][6] ));
 sg13g2_dfrbp_1 _16167_ (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1677),
    .D(_01614_),
    .Q_N(_05697_),
    .Q(\mem.mem[18][7] ));
 sg13g2_dfrbp_1 _16168_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1676),
    .D(_01615_),
    .Q_N(_05696_),
    .Q(\mem.mem[190][0] ));
 sg13g2_dfrbp_1 _16169_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1675),
    .D(_01616_),
    .Q_N(_05695_),
    .Q(\mem.mem[190][1] ));
 sg13g2_dfrbp_1 _16170_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1674),
    .D(_01617_),
    .Q_N(_05694_),
    .Q(\mem.mem[190][2] ));
 sg13g2_dfrbp_1 _16171_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1673),
    .D(_01618_),
    .Q_N(_05693_),
    .Q(\mem.mem[190][3] ));
 sg13g2_dfrbp_1 _16172_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1672),
    .D(_01619_),
    .Q_N(_05692_),
    .Q(\mem.mem[190][4] ));
 sg13g2_dfrbp_1 _16173_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1671),
    .D(_01620_),
    .Q_N(_05691_),
    .Q(\mem.mem[190][5] ));
 sg13g2_dfrbp_1 _16174_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1670),
    .D(_01621_),
    .Q_N(_05690_),
    .Q(\mem.mem[190][6] ));
 sg13g2_dfrbp_1 _16175_ (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1669),
    .D(_01622_),
    .Q_N(_05689_),
    .Q(\mem.mem[190][7] ));
 sg13g2_dfrbp_1 _16176_ (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1668),
    .D(_01623_),
    .Q_N(_05688_),
    .Q(\mem.mem[191][0] ));
 sg13g2_dfrbp_1 _16177_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1667),
    .D(_01624_),
    .Q_N(_05687_),
    .Q(\mem.mem[191][1] ));
 sg13g2_dfrbp_1 _16178_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1666),
    .D(_01625_),
    .Q_N(_05686_),
    .Q(\mem.mem[191][2] ));
 sg13g2_dfrbp_1 _16179_ (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1665),
    .D(_01626_),
    .Q_N(_05685_),
    .Q(\mem.mem[191][3] ));
 sg13g2_dfrbp_1 _16180_ (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1664),
    .D(_01627_),
    .Q_N(_05684_),
    .Q(\mem.mem[191][4] ));
 sg13g2_dfrbp_1 _16181_ (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1663),
    .D(_01628_),
    .Q_N(_05683_),
    .Q(\mem.mem[191][5] ));
 sg13g2_dfrbp_1 _16182_ (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1662),
    .D(_01629_),
    .Q_N(_05682_),
    .Q(\mem.mem[191][6] ));
 sg13g2_dfrbp_1 _16183_ (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1661),
    .D(_01630_),
    .Q_N(_05681_),
    .Q(\mem.mem[191][7] ));
 sg13g2_dfrbp_1 _16184_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1660),
    .D(_01631_),
    .Q_N(_05680_),
    .Q(\mem.mem[192][0] ));
 sg13g2_dfrbp_1 _16185_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1659),
    .D(_01632_),
    .Q_N(_05679_),
    .Q(\mem.mem[192][1] ));
 sg13g2_dfrbp_1 _16186_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1658),
    .D(_01633_),
    .Q_N(_05678_),
    .Q(\mem.mem[192][2] ));
 sg13g2_dfrbp_1 _16187_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1657),
    .D(_01634_),
    .Q_N(_05677_),
    .Q(\mem.mem[192][3] ));
 sg13g2_dfrbp_1 _16188_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1656),
    .D(_01635_),
    .Q_N(_05676_),
    .Q(\mem.mem[192][4] ));
 sg13g2_dfrbp_1 _16189_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1655),
    .D(_01636_),
    .Q_N(_05675_),
    .Q(\mem.mem[192][5] ));
 sg13g2_dfrbp_1 _16190_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1654),
    .D(_01637_),
    .Q_N(_05674_),
    .Q(\mem.mem[192][6] ));
 sg13g2_dfrbp_1 _16191_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1653),
    .D(_01638_),
    .Q_N(_05673_),
    .Q(\mem.mem[192][7] ));
 sg13g2_dfrbp_1 _16192_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1652),
    .D(_01639_),
    .Q_N(_05672_),
    .Q(\mem.mem[193][0] ));
 sg13g2_dfrbp_1 _16193_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1651),
    .D(_01640_),
    .Q_N(_05671_),
    .Q(\mem.mem[193][1] ));
 sg13g2_dfrbp_1 _16194_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1650),
    .D(_01641_),
    .Q_N(_05670_),
    .Q(\mem.mem[193][2] ));
 sg13g2_dfrbp_1 _16195_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1649),
    .D(_01642_),
    .Q_N(_05669_),
    .Q(\mem.mem[193][3] ));
 sg13g2_dfrbp_1 _16196_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1648),
    .D(_01643_),
    .Q_N(_05668_),
    .Q(\mem.mem[193][4] ));
 sg13g2_dfrbp_1 _16197_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1647),
    .D(_01644_),
    .Q_N(_05667_),
    .Q(\mem.mem[193][5] ));
 sg13g2_dfrbp_1 _16198_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1646),
    .D(_01645_),
    .Q_N(_05666_),
    .Q(\mem.mem[193][6] ));
 sg13g2_dfrbp_1 _16199_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1645),
    .D(_01646_),
    .Q_N(_05665_),
    .Q(\mem.mem[193][7] ));
 sg13g2_dfrbp_1 _16200_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1644),
    .D(_01647_),
    .Q_N(_05664_),
    .Q(\mem.mem[194][0] ));
 sg13g2_dfrbp_1 _16201_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1643),
    .D(_01648_),
    .Q_N(_05663_),
    .Q(\mem.mem[194][1] ));
 sg13g2_dfrbp_1 _16202_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1642),
    .D(_01649_),
    .Q_N(_05662_),
    .Q(\mem.mem[194][2] ));
 sg13g2_dfrbp_1 _16203_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1641),
    .D(_01650_),
    .Q_N(_05661_),
    .Q(\mem.mem[194][3] ));
 sg13g2_dfrbp_1 _16204_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1640),
    .D(_01651_),
    .Q_N(_05660_),
    .Q(\mem.mem[194][4] ));
 sg13g2_dfrbp_1 _16205_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1639),
    .D(_01652_),
    .Q_N(_05659_),
    .Q(\mem.mem[194][5] ));
 sg13g2_dfrbp_1 _16206_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1638),
    .D(_01653_),
    .Q_N(_05658_),
    .Q(\mem.mem[194][6] ));
 sg13g2_dfrbp_1 _16207_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1637),
    .D(_01654_),
    .Q_N(_05657_),
    .Q(\mem.mem[194][7] ));
 sg13g2_dfrbp_1 _16208_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1636),
    .D(_01655_),
    .Q_N(_05656_),
    .Q(\mem.mem[195][0] ));
 sg13g2_dfrbp_1 _16209_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1635),
    .D(_01656_),
    .Q_N(_05655_),
    .Q(\mem.mem[195][1] ));
 sg13g2_dfrbp_1 _16210_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1634),
    .D(_01657_),
    .Q_N(_05654_),
    .Q(\mem.mem[195][2] ));
 sg13g2_dfrbp_1 _16211_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1633),
    .D(_01658_),
    .Q_N(_05653_),
    .Q(\mem.mem[195][3] ));
 sg13g2_dfrbp_1 _16212_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1632),
    .D(_01659_),
    .Q_N(_05652_),
    .Q(\mem.mem[195][4] ));
 sg13g2_dfrbp_1 _16213_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1631),
    .D(_01660_),
    .Q_N(_05651_),
    .Q(\mem.mem[195][5] ));
 sg13g2_dfrbp_1 _16214_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1630),
    .D(_01661_),
    .Q_N(_05650_),
    .Q(\mem.mem[195][6] ));
 sg13g2_dfrbp_1 _16215_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1629),
    .D(_01662_),
    .Q_N(_05649_),
    .Q(\mem.mem[195][7] ));
 sg13g2_dfrbp_1 _16216_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1628),
    .D(_01663_),
    .Q_N(_05648_),
    .Q(\mem.mem[196][0] ));
 sg13g2_dfrbp_1 _16217_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1627),
    .D(_01664_),
    .Q_N(_05647_),
    .Q(\mem.mem[196][1] ));
 sg13g2_dfrbp_1 _16218_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1626),
    .D(_01665_),
    .Q_N(_05646_),
    .Q(\mem.mem[196][2] ));
 sg13g2_dfrbp_1 _16219_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1625),
    .D(_01666_),
    .Q_N(_05645_),
    .Q(\mem.mem[196][3] ));
 sg13g2_dfrbp_1 _16220_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1624),
    .D(_01667_),
    .Q_N(_05644_),
    .Q(\mem.mem[196][4] ));
 sg13g2_dfrbp_1 _16221_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1623),
    .D(_01668_),
    .Q_N(_05643_),
    .Q(\mem.mem[196][5] ));
 sg13g2_dfrbp_1 _16222_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1622),
    .D(_01669_),
    .Q_N(_05642_),
    .Q(\mem.mem[196][6] ));
 sg13g2_dfrbp_1 _16223_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1621),
    .D(_01670_),
    .Q_N(_05641_),
    .Q(\mem.mem[196][7] ));
 sg13g2_dfrbp_1 _16224_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1620),
    .D(_01671_),
    .Q_N(_05640_),
    .Q(\mem.mem[197][0] ));
 sg13g2_dfrbp_1 _16225_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1619),
    .D(_01672_),
    .Q_N(_05639_),
    .Q(\mem.mem[197][1] ));
 sg13g2_dfrbp_1 _16226_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1618),
    .D(_01673_),
    .Q_N(_05638_),
    .Q(\mem.mem[197][2] ));
 sg13g2_dfrbp_1 _16227_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1617),
    .D(_01674_),
    .Q_N(_05637_),
    .Q(\mem.mem[197][3] ));
 sg13g2_dfrbp_1 _16228_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1616),
    .D(_01675_),
    .Q_N(_05636_),
    .Q(\mem.mem[197][4] ));
 sg13g2_dfrbp_1 _16229_ (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1615),
    .D(_01676_),
    .Q_N(_05635_),
    .Q(\mem.mem[197][5] ));
 sg13g2_dfrbp_1 _16230_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1614),
    .D(_01677_),
    .Q_N(_05634_),
    .Q(\mem.mem[197][6] ));
 sg13g2_dfrbp_1 _16231_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1613),
    .D(_01678_),
    .Q_N(_05633_),
    .Q(\mem.mem[197][7] ));
 sg13g2_dfrbp_1 _16232_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1612),
    .D(_01679_),
    .Q_N(_05632_),
    .Q(\mem.mem[198][0] ));
 sg13g2_dfrbp_1 _16233_ (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1611),
    .D(_01680_),
    .Q_N(_05631_),
    .Q(\mem.mem[198][1] ));
 sg13g2_dfrbp_1 _16234_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1610),
    .D(_01681_),
    .Q_N(_05630_),
    .Q(\mem.mem[198][2] ));
 sg13g2_dfrbp_1 _16235_ (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1609),
    .D(_01682_),
    .Q_N(_05629_),
    .Q(\mem.mem[198][3] ));
 sg13g2_dfrbp_1 _16236_ (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1608),
    .D(_01683_),
    .Q_N(_05628_),
    .Q(\mem.mem[198][4] ));
 sg13g2_dfrbp_1 _16237_ (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1607),
    .D(_01684_),
    .Q_N(_05627_),
    .Q(\mem.mem[198][5] ));
 sg13g2_dfrbp_1 _16238_ (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1606),
    .D(_01685_),
    .Q_N(_05626_),
    .Q(\mem.mem[198][6] ));
 sg13g2_dfrbp_1 _16239_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1605),
    .D(_01686_),
    .Q_N(_05625_),
    .Q(\mem.mem[198][7] ));
 sg13g2_dfrbp_1 _16240_ (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1604),
    .D(_01687_),
    .Q_N(_05624_),
    .Q(\mem.mem[1][0] ));
 sg13g2_dfrbp_1 _16241_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1603),
    .D(_01688_),
    .Q_N(_05623_),
    .Q(\mem.mem[1][1] ));
 sg13g2_dfrbp_1 _16242_ (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1602),
    .D(_01689_),
    .Q_N(_05622_),
    .Q(\mem.mem[1][2] ));
 sg13g2_dfrbp_1 _16243_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1601),
    .D(_01690_),
    .Q_N(_05621_),
    .Q(\mem.mem[1][3] ));
 sg13g2_dfrbp_1 _16244_ (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1600),
    .D(_01691_),
    .Q_N(_05620_),
    .Q(\mem.mem[1][4] ));
 sg13g2_dfrbp_1 _16245_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1599),
    .D(_01692_),
    .Q_N(_05619_),
    .Q(\mem.mem[1][5] ));
 sg13g2_dfrbp_1 _16246_ (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1598),
    .D(_01693_),
    .Q_N(_05618_),
    .Q(\mem.mem[1][6] ));
 sg13g2_dfrbp_1 _16247_ (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1597),
    .D(_01694_),
    .Q_N(_05617_),
    .Q(\mem.mem[1][7] ));
 sg13g2_dfrbp_1 _16248_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1596),
    .D(_01695_),
    .Q_N(_05616_),
    .Q(\mem.mem[200][0] ));
 sg13g2_dfrbp_1 _16249_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1595),
    .D(_01696_),
    .Q_N(_05615_),
    .Q(\mem.mem[200][1] ));
 sg13g2_dfrbp_1 _16250_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1594),
    .D(_01697_),
    .Q_N(_05614_),
    .Q(\mem.mem[200][2] ));
 sg13g2_dfrbp_1 _16251_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1593),
    .D(_01698_),
    .Q_N(_05613_),
    .Q(\mem.mem[200][3] ));
 sg13g2_dfrbp_1 _16252_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1592),
    .D(_01699_),
    .Q_N(_05612_),
    .Q(\mem.mem[200][4] ));
 sg13g2_dfrbp_1 _16253_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1591),
    .D(_01700_),
    .Q_N(_05611_),
    .Q(\mem.mem[200][5] ));
 sg13g2_dfrbp_1 _16254_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1590),
    .D(_01701_),
    .Q_N(_05610_),
    .Q(\mem.mem[200][6] ));
 sg13g2_dfrbp_1 _16255_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1589),
    .D(_01702_),
    .Q_N(_05609_),
    .Q(\mem.mem[200][7] ));
 sg13g2_dfrbp_1 _16256_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1588),
    .D(_01703_),
    .Q_N(_05608_),
    .Q(\mem.mem[201][0] ));
 sg13g2_dfrbp_1 _16257_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1587),
    .D(_01704_),
    .Q_N(_05607_),
    .Q(\mem.mem[201][1] ));
 sg13g2_dfrbp_1 _16258_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1586),
    .D(_01705_),
    .Q_N(_05606_),
    .Q(\mem.mem[201][2] ));
 sg13g2_dfrbp_1 _16259_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1585),
    .D(_01706_),
    .Q_N(_05605_),
    .Q(\mem.mem[201][3] ));
 sg13g2_dfrbp_1 _16260_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1584),
    .D(_01707_),
    .Q_N(_05604_),
    .Q(\mem.mem[201][4] ));
 sg13g2_dfrbp_1 _16261_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1583),
    .D(_01708_),
    .Q_N(_05603_),
    .Q(\mem.mem[201][5] ));
 sg13g2_dfrbp_1 _16262_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1582),
    .D(_01709_),
    .Q_N(_05602_),
    .Q(\mem.mem[201][6] ));
 sg13g2_dfrbp_1 _16263_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1581),
    .D(_01710_),
    .Q_N(_05601_),
    .Q(\mem.mem[201][7] ));
 sg13g2_dfrbp_1 _16264_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1580),
    .D(_01711_),
    .Q_N(_05600_),
    .Q(\mem.mem[202][0] ));
 sg13g2_dfrbp_1 _16265_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1579),
    .D(_01712_),
    .Q_N(_05599_),
    .Q(\mem.mem[202][1] ));
 sg13g2_dfrbp_1 _16266_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1578),
    .D(_01713_),
    .Q_N(_05598_),
    .Q(\mem.mem[202][2] ));
 sg13g2_dfrbp_1 _16267_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1577),
    .D(_01714_),
    .Q_N(_05597_),
    .Q(\mem.mem[202][3] ));
 sg13g2_dfrbp_1 _16268_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1576),
    .D(_01715_),
    .Q_N(_05596_),
    .Q(\mem.mem[202][4] ));
 sg13g2_dfrbp_1 _16269_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1575),
    .D(_01716_),
    .Q_N(_05595_),
    .Q(\mem.mem[202][5] ));
 sg13g2_dfrbp_1 _16270_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1574),
    .D(_01717_),
    .Q_N(_05594_),
    .Q(\mem.mem[202][6] ));
 sg13g2_dfrbp_1 _16271_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1573),
    .D(_01718_),
    .Q_N(_05593_),
    .Q(\mem.mem[202][7] ));
 sg13g2_dfrbp_1 _16272_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1572),
    .D(_01719_),
    .Q_N(_05592_),
    .Q(\mem.mem[203][0] ));
 sg13g2_dfrbp_1 _16273_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1571),
    .D(_01720_),
    .Q_N(_05591_),
    .Q(\mem.mem[203][1] ));
 sg13g2_dfrbp_1 _16274_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1570),
    .D(_01721_),
    .Q_N(_05590_),
    .Q(\mem.mem[203][2] ));
 sg13g2_dfrbp_1 _16275_ (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1569),
    .D(_01722_),
    .Q_N(_05589_),
    .Q(\mem.mem[203][3] ));
 sg13g2_dfrbp_1 _16276_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1568),
    .D(_01723_),
    .Q_N(_05588_),
    .Q(\mem.mem[203][4] ));
 sg13g2_dfrbp_1 _16277_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1567),
    .D(_01724_),
    .Q_N(_05587_),
    .Q(\mem.mem[203][5] ));
 sg13g2_dfrbp_1 _16278_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1566),
    .D(_01725_),
    .Q_N(_05586_),
    .Q(\mem.mem[203][6] ));
 sg13g2_dfrbp_1 _16279_ (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1565),
    .D(_01726_),
    .Q_N(_05585_),
    .Q(\mem.mem[203][7] ));
 sg13g2_dfrbp_1 _16280_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1564),
    .D(_01727_),
    .Q_N(_05584_),
    .Q(\mem.mem[204][0] ));
 sg13g2_dfrbp_1 _16281_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1563),
    .D(_01728_),
    .Q_N(_05583_),
    .Q(\mem.mem[204][1] ));
 sg13g2_dfrbp_1 _16282_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1562),
    .D(_01729_),
    .Q_N(_05582_),
    .Q(\mem.mem[204][2] ));
 sg13g2_dfrbp_1 _16283_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1561),
    .D(_01730_),
    .Q_N(_05581_),
    .Q(\mem.mem[204][3] ));
 sg13g2_dfrbp_1 _16284_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1560),
    .D(_01731_),
    .Q_N(_05580_),
    .Q(\mem.mem[204][4] ));
 sg13g2_dfrbp_1 _16285_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1559),
    .D(_01732_),
    .Q_N(_05579_),
    .Q(\mem.mem[204][5] ));
 sg13g2_dfrbp_1 _16286_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1558),
    .D(_01733_),
    .Q_N(_05578_),
    .Q(\mem.mem[204][6] ));
 sg13g2_dfrbp_1 _16287_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1557),
    .D(_01734_),
    .Q_N(_05577_),
    .Q(\mem.mem[204][7] ));
 sg13g2_dfrbp_1 _16288_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1556),
    .D(_01735_),
    .Q_N(_05576_),
    .Q(\mem.mem[205][0] ));
 sg13g2_dfrbp_1 _16289_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1555),
    .D(_01736_),
    .Q_N(_05575_),
    .Q(\mem.mem[205][1] ));
 sg13g2_dfrbp_1 _16290_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1554),
    .D(_01737_),
    .Q_N(_05574_),
    .Q(\mem.mem[205][2] ));
 sg13g2_dfrbp_1 _16291_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1553),
    .D(_01738_),
    .Q_N(_05573_),
    .Q(\mem.mem[205][3] ));
 sg13g2_dfrbp_1 _16292_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1552),
    .D(_01739_),
    .Q_N(_05572_),
    .Q(\mem.mem[205][4] ));
 sg13g2_dfrbp_1 _16293_ (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1551),
    .D(_01740_),
    .Q_N(_05571_),
    .Q(\mem.mem[205][5] ));
 sg13g2_dfrbp_1 _16294_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1550),
    .D(_01741_),
    .Q_N(_05570_),
    .Q(\mem.mem[205][6] ));
 sg13g2_dfrbp_1 _16295_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1549),
    .D(_01742_),
    .Q_N(_05569_),
    .Q(\mem.mem[205][7] ));
 sg13g2_dfrbp_1 _16296_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1548),
    .D(_01743_),
    .Q_N(_05568_),
    .Q(\mem.mem[206][0] ));
 sg13g2_dfrbp_1 _16297_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1547),
    .D(_01744_),
    .Q_N(_05567_),
    .Q(\mem.mem[206][1] ));
 sg13g2_dfrbp_1 _16298_ (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1546),
    .D(_01745_),
    .Q_N(_05566_),
    .Q(\mem.mem[206][2] ));
 sg13g2_dfrbp_1 _16299_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1545),
    .D(_01746_),
    .Q_N(_05565_),
    .Q(\mem.mem[206][3] ));
 sg13g2_dfrbp_1 _16300_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1544),
    .D(_01747_),
    .Q_N(_05564_),
    .Q(\mem.mem[206][4] ));
 sg13g2_dfrbp_1 _16301_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1543),
    .D(_01748_),
    .Q_N(_05563_),
    .Q(\mem.mem[206][5] ));
 sg13g2_dfrbp_1 _16302_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1542),
    .D(_01749_),
    .Q_N(_05562_),
    .Q(\mem.mem[206][6] ));
 sg13g2_dfrbp_1 _16303_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1541),
    .D(_01750_),
    .Q_N(_05561_),
    .Q(\mem.mem[206][7] ));
 sg13g2_dfrbp_1 _16304_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1540),
    .D(_01751_),
    .Q_N(_05560_),
    .Q(\mem.mem[207][0] ));
 sg13g2_dfrbp_1 _16305_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1539),
    .D(_01752_),
    .Q_N(_05559_),
    .Q(\mem.mem[207][1] ));
 sg13g2_dfrbp_1 _16306_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1538),
    .D(_01753_),
    .Q_N(_05558_),
    .Q(\mem.mem[207][2] ));
 sg13g2_dfrbp_1 _16307_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1537),
    .D(_01754_),
    .Q_N(_05557_),
    .Q(\mem.mem[207][3] ));
 sg13g2_dfrbp_1 _16308_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1536),
    .D(_01755_),
    .Q_N(_05556_),
    .Q(\mem.mem[207][4] ));
 sg13g2_dfrbp_1 _16309_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1535),
    .D(_01756_),
    .Q_N(_05555_),
    .Q(\mem.mem[207][5] ));
 sg13g2_dfrbp_1 _16310_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1534),
    .D(_01757_),
    .Q_N(_05554_),
    .Q(\mem.mem[207][6] ));
 sg13g2_dfrbp_1 _16311_ (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1533),
    .D(_01758_),
    .Q_N(_05553_),
    .Q(\mem.mem[207][7] ));
 sg13g2_dfrbp_1 _16312_ (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1532),
    .D(_01759_),
    .Q_N(_05552_),
    .Q(\mem.mem[208][0] ));
 sg13g2_dfrbp_1 _16313_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1531),
    .D(_01760_),
    .Q_N(_05551_),
    .Q(\mem.mem[208][1] ));
 sg13g2_dfrbp_1 _16314_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1530),
    .D(_01761_),
    .Q_N(_05550_),
    .Q(\mem.mem[208][2] ));
 sg13g2_dfrbp_1 _16315_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1529),
    .D(_01762_),
    .Q_N(_05549_),
    .Q(\mem.mem[208][3] ));
 sg13g2_dfrbp_1 _16316_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1528),
    .D(_01763_),
    .Q_N(_05548_),
    .Q(\mem.mem[208][4] ));
 sg13g2_dfrbp_1 _16317_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1527),
    .D(_01764_),
    .Q_N(_05547_),
    .Q(\mem.mem[208][5] ));
 sg13g2_dfrbp_1 _16318_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1526),
    .D(_01765_),
    .Q_N(_05546_),
    .Q(\mem.mem[208][6] ));
 sg13g2_dfrbp_1 _16319_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1525),
    .D(_01766_),
    .Q_N(_05545_),
    .Q(\mem.mem[208][7] ));
 sg13g2_dfrbp_1 _16320_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1524),
    .D(_01767_),
    .Q_N(_05544_),
    .Q(\mem.mem[20][0] ));
 sg13g2_dfrbp_1 _16321_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1523),
    .D(_01768_),
    .Q_N(_05543_),
    .Q(\mem.mem[20][1] ));
 sg13g2_dfrbp_1 _16322_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1522),
    .D(_01769_),
    .Q_N(_05542_),
    .Q(\mem.mem[20][2] ));
 sg13g2_dfrbp_1 _16323_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1521),
    .D(_01770_),
    .Q_N(_05541_),
    .Q(\mem.mem[20][3] ));
 sg13g2_dfrbp_1 _16324_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1520),
    .D(_01771_),
    .Q_N(_05540_),
    .Q(\mem.mem[20][4] ));
 sg13g2_dfrbp_1 _16325_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1519),
    .D(_01772_),
    .Q_N(_05539_),
    .Q(\mem.mem[20][5] ));
 sg13g2_dfrbp_1 _16326_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1518),
    .D(_01773_),
    .Q_N(_05538_),
    .Q(\mem.mem[20][6] ));
 sg13g2_dfrbp_1 _16327_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1517),
    .D(_01774_),
    .Q_N(_05537_),
    .Q(\mem.mem[20][7] ));
 sg13g2_dfrbp_1 _16328_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1516),
    .D(_01775_),
    .Q_N(_05536_),
    .Q(\mem.mem[210][0] ));
 sg13g2_dfrbp_1 _16329_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1515),
    .D(_01776_),
    .Q_N(_05535_),
    .Q(\mem.mem[210][1] ));
 sg13g2_dfrbp_1 _16330_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1514),
    .D(_01777_),
    .Q_N(_05534_),
    .Q(\mem.mem[210][2] ));
 sg13g2_dfrbp_1 _16331_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1513),
    .D(_01778_),
    .Q_N(_05533_),
    .Q(\mem.mem[210][3] ));
 sg13g2_dfrbp_1 _16332_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1512),
    .D(_01779_),
    .Q_N(_05532_),
    .Q(\mem.mem[210][4] ));
 sg13g2_dfrbp_1 _16333_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1511),
    .D(_01780_),
    .Q_N(_05531_),
    .Q(\mem.mem[210][5] ));
 sg13g2_dfrbp_1 _16334_ (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1510),
    .D(_01781_),
    .Q_N(_05530_),
    .Q(\mem.mem[210][6] ));
 sg13g2_dfrbp_1 _16335_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1509),
    .D(_01782_),
    .Q_N(_05529_),
    .Q(\mem.mem[210][7] ));
 sg13g2_dfrbp_1 _16336_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1508),
    .D(_01783_),
    .Q_N(_05528_),
    .Q(\mem.mem[211][0] ));
 sg13g2_dfrbp_1 _16337_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1507),
    .D(_01784_),
    .Q_N(_05527_),
    .Q(\mem.mem[211][1] ));
 sg13g2_dfrbp_1 _16338_ (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1506),
    .D(_01785_),
    .Q_N(_05526_),
    .Q(\mem.mem[211][2] ));
 sg13g2_dfrbp_1 _16339_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1505),
    .D(_01786_),
    .Q_N(_05525_),
    .Q(\mem.mem[211][3] ));
 sg13g2_dfrbp_1 _16340_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1504),
    .D(_01787_),
    .Q_N(_05524_),
    .Q(\mem.mem[211][4] ));
 sg13g2_dfrbp_1 _16341_ (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1503),
    .D(_01788_),
    .Q_N(_05523_),
    .Q(\mem.mem[211][5] ));
 sg13g2_dfrbp_1 _16342_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1502),
    .D(_01789_),
    .Q_N(_05522_),
    .Q(\mem.mem[211][6] ));
 sg13g2_dfrbp_1 _16343_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1501),
    .D(_01790_),
    .Q_N(_05521_),
    .Q(\mem.mem[211][7] ));
 sg13g2_dfrbp_1 _16344_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1500),
    .D(_01791_),
    .Q_N(_05520_),
    .Q(\mem.mem[212][0] ));
 sg13g2_dfrbp_1 _16345_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1499),
    .D(_01792_),
    .Q_N(_05519_),
    .Q(\mem.mem[212][1] ));
 sg13g2_dfrbp_1 _16346_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1498),
    .D(_01793_),
    .Q_N(_05518_),
    .Q(\mem.mem[212][2] ));
 sg13g2_dfrbp_1 _16347_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1497),
    .D(_01794_),
    .Q_N(_05517_),
    .Q(\mem.mem[212][3] ));
 sg13g2_dfrbp_1 _16348_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1496),
    .D(_01795_),
    .Q_N(_05516_),
    .Q(\mem.mem[212][4] ));
 sg13g2_dfrbp_1 _16349_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1495),
    .D(_01796_),
    .Q_N(_05515_),
    .Q(\mem.mem[212][5] ));
 sg13g2_dfrbp_1 _16350_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1494),
    .D(_01797_),
    .Q_N(_05514_),
    .Q(\mem.mem[212][6] ));
 sg13g2_dfrbp_1 _16351_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1493),
    .D(_01798_),
    .Q_N(_05513_),
    .Q(\mem.mem[212][7] ));
 sg13g2_dfrbp_1 _16352_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1492),
    .D(_01799_),
    .Q_N(_05512_),
    .Q(\mem.mem[213][0] ));
 sg13g2_dfrbp_1 _16353_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1491),
    .D(_01800_),
    .Q_N(_05511_),
    .Q(\mem.mem[213][1] ));
 sg13g2_dfrbp_1 _16354_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1490),
    .D(_01801_),
    .Q_N(_05510_),
    .Q(\mem.mem[213][2] ));
 sg13g2_dfrbp_1 _16355_ (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1489),
    .D(_01802_),
    .Q_N(_05509_),
    .Q(\mem.mem[213][3] ));
 sg13g2_dfrbp_1 _16356_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1488),
    .D(_01803_),
    .Q_N(_05508_),
    .Q(\mem.mem[213][4] ));
 sg13g2_dfrbp_1 _16357_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1487),
    .D(_01804_),
    .Q_N(_05507_),
    .Q(\mem.mem[213][5] ));
 sg13g2_dfrbp_1 _16358_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1486),
    .D(_01805_),
    .Q_N(_05506_),
    .Q(\mem.mem[213][6] ));
 sg13g2_dfrbp_1 _16359_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1485),
    .D(_01806_),
    .Q_N(_05505_),
    .Q(\mem.mem[213][7] ));
 sg13g2_dfrbp_1 _16360_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1484),
    .D(_01807_),
    .Q_N(_05504_),
    .Q(\mem.mem[214][0] ));
 sg13g2_dfrbp_1 _16361_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1483),
    .D(_01808_),
    .Q_N(_05503_),
    .Q(\mem.mem[214][1] ));
 sg13g2_dfrbp_1 _16362_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1482),
    .D(_01809_),
    .Q_N(_05502_),
    .Q(\mem.mem[214][2] ));
 sg13g2_dfrbp_1 _16363_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1481),
    .D(_01810_),
    .Q_N(_05501_),
    .Q(\mem.mem[214][3] ));
 sg13g2_dfrbp_1 _16364_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1480),
    .D(_01811_),
    .Q_N(_05500_),
    .Q(\mem.mem[214][4] ));
 sg13g2_dfrbp_1 _16365_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1479),
    .D(_01812_),
    .Q_N(_05499_),
    .Q(\mem.mem[214][5] ));
 sg13g2_dfrbp_1 _16366_ (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1478),
    .D(_01813_),
    .Q_N(_05498_),
    .Q(\mem.mem[214][6] ));
 sg13g2_dfrbp_1 _16367_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1477),
    .D(_01814_),
    .Q_N(_05497_),
    .Q(\mem.mem[214][7] ));
 sg13g2_dfrbp_1 _16368_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1476),
    .D(_01815_),
    .Q_N(_05496_),
    .Q(\mem.mem[215][0] ));
 sg13g2_dfrbp_1 _16369_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1475),
    .D(_01816_),
    .Q_N(_05495_),
    .Q(\mem.mem[215][1] ));
 sg13g2_dfrbp_1 _16370_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1474),
    .D(_01817_),
    .Q_N(_05494_),
    .Q(\mem.mem[215][2] ));
 sg13g2_dfrbp_1 _16371_ (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1473),
    .D(_01818_),
    .Q_N(_05493_),
    .Q(\mem.mem[215][3] ));
 sg13g2_dfrbp_1 _16372_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1472),
    .D(_01819_),
    .Q_N(_05492_),
    .Q(\mem.mem[215][4] ));
 sg13g2_dfrbp_1 _16373_ (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1471),
    .D(_01820_),
    .Q_N(_05491_),
    .Q(\mem.mem[215][5] ));
 sg13g2_dfrbp_1 _16374_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1470),
    .D(_01821_),
    .Q_N(_05490_),
    .Q(\mem.mem[215][6] ));
 sg13g2_dfrbp_1 _16375_ (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1469),
    .D(_01822_),
    .Q_N(_05489_),
    .Q(\mem.mem[215][7] ));
 sg13g2_dfrbp_1 _16376_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1468),
    .D(_01823_),
    .Q_N(_05488_),
    .Q(\mem.mem[216][0] ));
 sg13g2_dfrbp_1 _16377_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1467),
    .D(_01824_),
    .Q_N(_05487_),
    .Q(\mem.mem[216][1] ));
 sg13g2_dfrbp_1 _16378_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1466),
    .D(_01825_),
    .Q_N(_05486_),
    .Q(\mem.mem[216][2] ));
 sg13g2_dfrbp_1 _16379_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1465),
    .D(_01826_),
    .Q_N(_05485_),
    .Q(\mem.mem[216][3] ));
 sg13g2_dfrbp_1 _16380_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1464),
    .D(_01827_),
    .Q_N(_05484_),
    .Q(\mem.mem[216][4] ));
 sg13g2_dfrbp_1 _16381_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1463),
    .D(_01828_),
    .Q_N(_05483_),
    .Q(\mem.mem[216][5] ));
 sg13g2_dfrbp_1 _16382_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1462),
    .D(_01829_),
    .Q_N(_05482_),
    .Q(\mem.mem[216][6] ));
 sg13g2_dfrbp_1 _16383_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1461),
    .D(_01830_),
    .Q_N(_05481_),
    .Q(\mem.mem[216][7] ));
 sg13g2_dfrbp_1 _16384_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1460),
    .D(_01831_),
    .Q_N(_05480_),
    .Q(\mem.mem[217][0] ));
 sg13g2_dfrbp_1 _16385_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1459),
    .D(_01832_),
    .Q_N(_05479_),
    .Q(\mem.mem[217][1] ));
 sg13g2_dfrbp_1 _16386_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1458),
    .D(_01833_),
    .Q_N(_05478_),
    .Q(\mem.mem[217][2] ));
 sg13g2_dfrbp_1 _16387_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1457),
    .D(_01834_),
    .Q_N(_05477_),
    .Q(\mem.mem[217][3] ));
 sg13g2_dfrbp_1 _16388_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1456),
    .D(_01835_),
    .Q_N(_05476_),
    .Q(\mem.mem[217][4] ));
 sg13g2_dfrbp_1 _16389_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1455),
    .D(_01836_),
    .Q_N(_05475_),
    .Q(\mem.mem[217][5] ));
 sg13g2_dfrbp_1 _16390_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1454),
    .D(_01837_),
    .Q_N(_05474_),
    .Q(\mem.mem[217][6] ));
 sg13g2_dfrbp_1 _16391_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1453),
    .D(_01838_),
    .Q_N(_05473_),
    .Q(\mem.mem[217][7] ));
 sg13g2_dfrbp_1 _16392_ (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1452),
    .D(_01839_),
    .Q_N(_05472_),
    .Q(\mem.mem[218][0] ));
 sg13g2_dfrbp_1 _16393_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1451),
    .D(_01840_),
    .Q_N(_05471_),
    .Q(\mem.mem[218][1] ));
 sg13g2_dfrbp_1 _16394_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1450),
    .D(_01841_),
    .Q_N(_05470_),
    .Q(\mem.mem[218][2] ));
 sg13g2_dfrbp_1 _16395_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1449),
    .D(_01842_),
    .Q_N(_05469_),
    .Q(\mem.mem[218][3] ));
 sg13g2_dfrbp_1 _16396_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1448),
    .D(_01843_),
    .Q_N(_05468_),
    .Q(\mem.mem[218][4] ));
 sg13g2_dfrbp_1 _16397_ (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1447),
    .D(_01844_),
    .Q_N(_05467_),
    .Q(\mem.mem[218][5] ));
 sg13g2_dfrbp_1 _16398_ (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1446),
    .D(_01845_),
    .Q_N(_05466_),
    .Q(\mem.mem[218][6] ));
 sg13g2_dfrbp_1 _16399_ (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1445),
    .D(_01846_),
    .Q_N(_05465_),
    .Q(\mem.mem[218][7] ));
 sg13g2_dfrbp_1 _16400_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1444),
    .D(_01847_),
    .Q_N(_05464_),
    .Q(\mem.mem[21][0] ));
 sg13g2_dfrbp_1 _16401_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1443),
    .D(_01848_),
    .Q_N(_05463_),
    .Q(\mem.mem[21][1] ));
 sg13g2_dfrbp_1 _16402_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1442),
    .D(_01849_),
    .Q_N(_05462_),
    .Q(\mem.mem[21][2] ));
 sg13g2_dfrbp_1 _16403_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1441),
    .D(_01850_),
    .Q_N(_05461_),
    .Q(\mem.mem[21][3] ));
 sg13g2_dfrbp_1 _16404_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1440),
    .D(_01851_),
    .Q_N(_05460_),
    .Q(\mem.mem[21][4] ));
 sg13g2_dfrbp_1 _16405_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1439),
    .D(_01852_),
    .Q_N(_05459_),
    .Q(\mem.mem[21][5] ));
 sg13g2_dfrbp_1 _16406_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1438),
    .D(_01853_),
    .Q_N(_05458_),
    .Q(\mem.mem[21][6] ));
 sg13g2_dfrbp_1 _16407_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1437),
    .D(_01854_),
    .Q_N(_05457_),
    .Q(\mem.mem[21][7] ));
 sg13g2_dfrbp_1 _16408_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1436),
    .D(_01855_),
    .Q_N(_05456_),
    .Q(\mem.mem[220][0] ));
 sg13g2_dfrbp_1 _16409_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1435),
    .D(_01856_),
    .Q_N(_05455_),
    .Q(\mem.mem[220][1] ));
 sg13g2_dfrbp_1 _16410_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1434),
    .D(_01857_),
    .Q_N(_05454_),
    .Q(\mem.mem[220][2] ));
 sg13g2_dfrbp_1 _16411_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1433),
    .D(_01858_),
    .Q_N(_05453_),
    .Q(\mem.mem[220][3] ));
 sg13g2_dfrbp_1 _16412_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1432),
    .D(_01859_),
    .Q_N(_05452_),
    .Q(\mem.mem[220][4] ));
 sg13g2_dfrbp_1 _16413_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1431),
    .D(_01860_),
    .Q_N(_05451_),
    .Q(\mem.mem[220][5] ));
 sg13g2_dfrbp_1 _16414_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1430),
    .D(_01861_),
    .Q_N(_05450_),
    .Q(\mem.mem[220][6] ));
 sg13g2_dfrbp_1 _16415_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1429),
    .D(_01862_),
    .Q_N(_05449_),
    .Q(\mem.mem[220][7] ));
 sg13g2_dfrbp_1 _16416_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1428),
    .D(_01863_),
    .Q_N(_05448_),
    .Q(\mem.mem[221][0] ));
 sg13g2_dfrbp_1 _16417_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1427),
    .D(_01864_),
    .Q_N(_05447_),
    .Q(\mem.mem[221][1] ));
 sg13g2_dfrbp_1 _16418_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1426),
    .D(_01865_),
    .Q_N(_05446_),
    .Q(\mem.mem[221][2] ));
 sg13g2_dfrbp_1 _16419_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1425),
    .D(_01866_),
    .Q_N(_05445_),
    .Q(\mem.mem[221][3] ));
 sg13g2_dfrbp_1 _16420_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1424),
    .D(_01867_),
    .Q_N(_05444_),
    .Q(\mem.mem[221][4] ));
 sg13g2_dfrbp_1 _16421_ (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1423),
    .D(_01868_),
    .Q_N(_05443_),
    .Q(\mem.mem[221][5] ));
 sg13g2_dfrbp_1 _16422_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1422),
    .D(_01869_),
    .Q_N(_05442_),
    .Q(\mem.mem[221][6] ));
 sg13g2_dfrbp_1 _16423_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1421),
    .D(_01870_),
    .Q_N(_05441_),
    .Q(\mem.mem[221][7] ));
 sg13g2_dfrbp_1 _16424_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1420),
    .D(_01871_),
    .Q_N(_05440_),
    .Q(\mem.mem[222][0] ));
 sg13g2_dfrbp_1 _16425_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1419),
    .D(_01872_),
    .Q_N(_05439_),
    .Q(\mem.mem[222][1] ));
 sg13g2_dfrbp_1 _16426_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1418),
    .D(_01873_),
    .Q_N(_05438_),
    .Q(\mem.mem[222][2] ));
 sg13g2_dfrbp_1 _16427_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1417),
    .D(_01874_),
    .Q_N(_05437_),
    .Q(\mem.mem[222][3] ));
 sg13g2_dfrbp_1 _16428_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1416),
    .D(_01875_),
    .Q_N(_05436_),
    .Q(\mem.mem[222][4] ));
 sg13g2_dfrbp_1 _16429_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1415),
    .D(_01876_),
    .Q_N(_05435_),
    .Q(\mem.mem[222][5] ));
 sg13g2_dfrbp_1 _16430_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1414),
    .D(_01877_),
    .Q_N(_05434_),
    .Q(\mem.mem[222][6] ));
 sg13g2_dfrbp_1 _16431_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1413),
    .D(_01878_),
    .Q_N(_05433_),
    .Q(\mem.mem[222][7] ));
 sg13g2_dfrbp_1 _16432_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1412),
    .D(_01879_),
    .Q_N(_05432_),
    .Q(\mem.mem[223][0] ));
 sg13g2_dfrbp_1 _16433_ (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1411),
    .D(_01880_),
    .Q_N(_05431_),
    .Q(\mem.mem[223][1] ));
 sg13g2_dfrbp_1 _16434_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1410),
    .D(_01881_),
    .Q_N(_05430_),
    .Q(\mem.mem[223][2] ));
 sg13g2_dfrbp_1 _16435_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1409),
    .D(_01882_),
    .Q_N(_05429_),
    .Q(\mem.mem[223][3] ));
 sg13g2_dfrbp_1 _16436_ (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1408),
    .D(_01883_),
    .Q_N(_05428_),
    .Q(\mem.mem[223][4] ));
 sg13g2_dfrbp_1 _16437_ (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1407),
    .D(_01884_),
    .Q_N(_05427_),
    .Q(\mem.mem[223][5] ));
 sg13g2_dfrbp_1 _16438_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1406),
    .D(_01885_),
    .Q_N(_05426_),
    .Q(\mem.mem[223][6] ));
 sg13g2_dfrbp_1 _16439_ (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1405),
    .D(_01886_),
    .Q_N(_05425_),
    .Q(\mem.mem[223][7] ));
 sg13g2_dfrbp_1 _16440_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1404),
    .D(_01887_),
    .Q_N(_05424_),
    .Q(\mem.mem[224][0] ));
 sg13g2_dfrbp_1 _16441_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1403),
    .D(_01888_),
    .Q_N(_05423_),
    .Q(\mem.mem[224][1] ));
 sg13g2_dfrbp_1 _16442_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1402),
    .D(_01889_),
    .Q_N(_05422_),
    .Q(\mem.mem[224][2] ));
 sg13g2_dfrbp_1 _16443_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1401),
    .D(_01890_),
    .Q_N(_05421_),
    .Q(\mem.mem[224][3] ));
 sg13g2_dfrbp_1 _16444_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1400),
    .D(_01891_),
    .Q_N(_05420_),
    .Q(\mem.mem[224][4] ));
 sg13g2_dfrbp_1 _16445_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1399),
    .D(_01892_),
    .Q_N(_05419_),
    .Q(\mem.mem[224][5] ));
 sg13g2_dfrbp_1 _16446_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1398),
    .D(_01893_),
    .Q_N(_05418_),
    .Q(\mem.mem[224][6] ));
 sg13g2_dfrbp_1 _16447_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1397),
    .D(_01894_),
    .Q_N(_05417_),
    .Q(\mem.mem[224][7] ));
 sg13g2_dfrbp_1 _16448_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1396),
    .D(_01895_),
    .Q_N(_05416_),
    .Q(\mem.mem[225][0] ));
 sg13g2_dfrbp_1 _16449_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1395),
    .D(_01896_),
    .Q_N(_05415_),
    .Q(\mem.mem[225][1] ));
 sg13g2_dfrbp_1 _16450_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1394),
    .D(_01897_),
    .Q_N(_05414_),
    .Q(\mem.mem[225][2] ));
 sg13g2_dfrbp_1 _16451_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1393),
    .D(_01898_),
    .Q_N(_05413_),
    .Q(\mem.mem[225][3] ));
 sg13g2_dfrbp_1 _16452_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1392),
    .D(_01899_),
    .Q_N(_05412_),
    .Q(\mem.mem[225][4] ));
 sg13g2_dfrbp_1 _16453_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1391),
    .D(_01900_),
    .Q_N(_05411_),
    .Q(\mem.mem[225][5] ));
 sg13g2_dfrbp_1 _16454_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1390),
    .D(_01901_),
    .Q_N(_05410_),
    .Q(\mem.mem[225][6] ));
 sg13g2_dfrbp_1 _16455_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1389),
    .D(_01902_),
    .Q_N(_05409_),
    .Q(\mem.mem[225][7] ));
 sg13g2_dfrbp_1 _16456_ (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1388),
    .D(_01903_),
    .Q_N(_05408_),
    .Q(\mem.mem[226][0] ));
 sg13g2_dfrbp_1 _16457_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1387),
    .D(_01904_),
    .Q_N(_05407_),
    .Q(\mem.mem[226][1] ));
 sg13g2_dfrbp_1 _16458_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1386),
    .D(_01905_),
    .Q_N(_05406_),
    .Q(\mem.mem[226][2] ));
 sg13g2_dfrbp_1 _16459_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1385),
    .D(_01906_),
    .Q_N(_05405_),
    .Q(\mem.mem[226][3] ));
 sg13g2_dfrbp_1 _16460_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1384),
    .D(_01907_),
    .Q_N(_05404_),
    .Q(\mem.mem[226][4] ));
 sg13g2_dfrbp_1 _16461_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1383),
    .D(_01908_),
    .Q_N(_05403_),
    .Q(\mem.mem[226][5] ));
 sg13g2_dfrbp_1 _16462_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1382),
    .D(_01909_),
    .Q_N(_05402_),
    .Q(\mem.mem[226][6] ));
 sg13g2_dfrbp_1 _16463_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1381),
    .D(_01910_),
    .Q_N(_05401_),
    .Q(\mem.mem[226][7] ));
 sg13g2_dfrbp_1 _16464_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1380),
    .D(_01911_),
    .Q_N(_05400_),
    .Q(\mem.mem[227][0] ));
 sg13g2_dfrbp_1 _16465_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1379),
    .D(_01912_),
    .Q_N(_05399_),
    .Q(\mem.mem[227][1] ));
 sg13g2_dfrbp_1 _16466_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1378),
    .D(_01913_),
    .Q_N(_05398_),
    .Q(\mem.mem[227][2] ));
 sg13g2_dfrbp_1 _16467_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1377),
    .D(_01914_),
    .Q_N(_05397_),
    .Q(\mem.mem[227][3] ));
 sg13g2_dfrbp_1 _16468_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1376),
    .D(_01915_),
    .Q_N(_05396_),
    .Q(\mem.mem[227][4] ));
 sg13g2_dfrbp_1 _16469_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1375),
    .D(_01916_),
    .Q_N(_05395_),
    .Q(\mem.mem[227][5] ));
 sg13g2_dfrbp_1 _16470_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1374),
    .D(_01917_),
    .Q_N(_05394_),
    .Q(\mem.mem[227][6] ));
 sg13g2_dfrbp_1 _16471_ (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1373),
    .D(_01918_),
    .Q_N(_05393_),
    .Q(\mem.mem[227][7] ));
 sg13g2_dfrbp_1 _16472_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1372),
    .D(_01919_),
    .Q_N(_05392_),
    .Q(\mem.mem[228][0] ));
 sg13g2_dfrbp_1 _16473_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1371),
    .D(_01920_),
    .Q_N(_05391_),
    .Q(\mem.mem[228][1] ));
 sg13g2_dfrbp_1 _16474_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1370),
    .D(_01921_),
    .Q_N(_05390_),
    .Q(\mem.mem[228][2] ));
 sg13g2_dfrbp_1 _16475_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1369),
    .D(_01922_),
    .Q_N(_05389_),
    .Q(\mem.mem[228][3] ));
 sg13g2_dfrbp_1 _16476_ (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1368),
    .D(_01923_),
    .Q_N(_05388_),
    .Q(\mem.mem[228][4] ));
 sg13g2_dfrbp_1 _16477_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1367),
    .D(_01924_),
    .Q_N(_05387_),
    .Q(\mem.mem[228][5] ));
 sg13g2_dfrbp_1 _16478_ (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1366),
    .D(_01925_),
    .Q_N(_05386_),
    .Q(\mem.mem[228][6] ));
 sg13g2_dfrbp_1 _16479_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1365),
    .D(_01926_),
    .Q_N(_05385_),
    .Q(\mem.mem[228][7] ));
 sg13g2_dfrbp_1 _16480_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1364),
    .D(_01927_),
    .Q_N(_05384_),
    .Q(\mem.mem[22][0] ));
 sg13g2_dfrbp_1 _16481_ (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1363),
    .D(_01928_),
    .Q_N(_05383_),
    .Q(\mem.mem[22][1] ));
 sg13g2_dfrbp_1 _16482_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1362),
    .D(_01929_),
    .Q_N(_05382_),
    .Q(\mem.mem[22][2] ));
 sg13g2_dfrbp_1 _16483_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1361),
    .D(_01930_),
    .Q_N(_05381_),
    .Q(\mem.mem[22][3] ));
 sg13g2_dfrbp_1 _16484_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1360),
    .D(_01931_),
    .Q_N(_05380_),
    .Q(\mem.mem[22][4] ));
 sg13g2_dfrbp_1 _16485_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1359),
    .D(_01932_),
    .Q_N(_05379_),
    .Q(\mem.mem[22][5] ));
 sg13g2_dfrbp_1 _16486_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1358),
    .D(_01933_),
    .Q_N(_05378_),
    .Q(\mem.mem[22][6] ));
 sg13g2_dfrbp_1 _16487_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1357),
    .D(_01934_),
    .Q_N(_05377_),
    .Q(\mem.mem[22][7] ));
 sg13g2_dfrbp_1 _16488_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1356),
    .D(_01935_),
    .Q_N(_05376_),
    .Q(\mem.mem[230][0] ));
 sg13g2_dfrbp_1 _16489_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1355),
    .D(_01936_),
    .Q_N(_05375_),
    .Q(\mem.mem[230][1] ));
 sg13g2_dfrbp_1 _16490_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1354),
    .D(_01937_),
    .Q_N(_05374_),
    .Q(\mem.mem[230][2] ));
 sg13g2_dfrbp_1 _16491_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1353),
    .D(_01938_),
    .Q_N(_05373_),
    .Q(\mem.mem[230][3] ));
 sg13g2_dfrbp_1 _16492_ (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1352),
    .D(_01939_),
    .Q_N(_05372_),
    .Q(\mem.mem[230][4] ));
 sg13g2_dfrbp_1 _16493_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1351),
    .D(_01940_),
    .Q_N(_05371_),
    .Q(\mem.mem[230][5] ));
 sg13g2_dfrbp_1 _16494_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1350),
    .D(_01941_),
    .Q_N(_05370_),
    .Q(\mem.mem[230][6] ));
 sg13g2_dfrbp_1 _16495_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1349),
    .D(_01942_),
    .Q_N(_05369_),
    .Q(\mem.mem[230][7] ));
 sg13g2_dfrbp_1 _16496_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1348),
    .D(_01943_),
    .Q_N(_05368_),
    .Q(\mem.mem[231][0] ));
 sg13g2_dfrbp_1 _16497_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1347),
    .D(_01944_),
    .Q_N(_05367_),
    .Q(\mem.mem[231][1] ));
 sg13g2_dfrbp_1 _16498_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1346),
    .D(_01945_),
    .Q_N(_05366_),
    .Q(\mem.mem[231][2] ));
 sg13g2_dfrbp_1 _16499_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1345),
    .D(_01946_),
    .Q_N(_05365_),
    .Q(\mem.mem[231][3] ));
 sg13g2_dfrbp_1 _16500_ (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1344),
    .D(_01947_),
    .Q_N(_05364_),
    .Q(\mem.mem[231][4] ));
 sg13g2_dfrbp_1 _16501_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1343),
    .D(_01948_),
    .Q_N(_05363_),
    .Q(\mem.mem[231][5] ));
 sg13g2_dfrbp_1 _16502_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1342),
    .D(_01949_),
    .Q_N(_05362_),
    .Q(\mem.mem[231][6] ));
 sg13g2_dfrbp_1 _16503_ (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1341),
    .D(_01950_),
    .Q_N(_05361_),
    .Q(\mem.mem[231][7] ));
 sg13g2_dfrbp_1 _16504_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1340),
    .D(_01951_),
    .Q_N(_05360_),
    .Q(\mem.mem[232][0] ));
 sg13g2_dfrbp_1 _16505_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1339),
    .D(_01952_),
    .Q_N(_05359_),
    .Q(\mem.mem[232][1] ));
 sg13g2_dfrbp_1 _16506_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1338),
    .D(_01953_),
    .Q_N(_05358_),
    .Q(\mem.mem[232][2] ));
 sg13g2_dfrbp_1 _16507_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1337),
    .D(_01954_),
    .Q_N(_05357_),
    .Q(\mem.mem[232][3] ));
 sg13g2_dfrbp_1 _16508_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1336),
    .D(_01955_),
    .Q_N(_05356_),
    .Q(\mem.mem[232][4] ));
 sg13g2_dfrbp_1 _16509_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1335),
    .D(_01956_),
    .Q_N(_05355_),
    .Q(\mem.mem[232][5] ));
 sg13g2_dfrbp_1 _16510_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1334),
    .D(_01957_),
    .Q_N(_05354_),
    .Q(\mem.mem[232][6] ));
 sg13g2_dfrbp_1 _16511_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1333),
    .D(_01958_),
    .Q_N(_05353_),
    .Q(\mem.mem[232][7] ));
 sg13g2_dfrbp_1 _16512_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1332),
    .D(_01959_),
    .Q_N(_05352_),
    .Q(\mem.mem[233][0] ));
 sg13g2_dfrbp_1 _16513_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1331),
    .D(_01960_),
    .Q_N(_05351_),
    .Q(\mem.mem[233][1] ));
 sg13g2_dfrbp_1 _16514_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1330),
    .D(_01961_),
    .Q_N(_05350_),
    .Q(\mem.mem[233][2] ));
 sg13g2_dfrbp_1 _16515_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1329),
    .D(_01962_),
    .Q_N(_05349_),
    .Q(\mem.mem[233][3] ));
 sg13g2_dfrbp_1 _16516_ (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1328),
    .D(_01963_),
    .Q_N(_05348_),
    .Q(\mem.mem[233][4] ));
 sg13g2_dfrbp_1 _16517_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1327),
    .D(_01964_),
    .Q_N(_05347_),
    .Q(\mem.mem[233][5] ));
 sg13g2_dfrbp_1 _16518_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1326),
    .D(_01965_),
    .Q_N(_05346_),
    .Q(\mem.mem[233][6] ));
 sg13g2_dfrbp_1 _16519_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1325),
    .D(_01966_),
    .Q_N(_05345_),
    .Q(\mem.mem[233][7] ));
 sg13g2_dfrbp_1 _16520_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1324),
    .D(_01967_),
    .Q_N(_05344_),
    .Q(\mem.mem[234][0] ));
 sg13g2_dfrbp_1 _16521_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1323),
    .D(_01968_),
    .Q_N(_05343_),
    .Q(\mem.mem[234][1] ));
 sg13g2_dfrbp_1 _16522_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1322),
    .D(_01969_),
    .Q_N(_05342_),
    .Q(\mem.mem[234][2] ));
 sg13g2_dfrbp_1 _16523_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1321),
    .D(_01970_),
    .Q_N(_05341_),
    .Q(\mem.mem[234][3] ));
 sg13g2_dfrbp_1 _16524_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1320),
    .D(_01971_),
    .Q_N(_05340_),
    .Q(\mem.mem[234][4] ));
 sg13g2_dfrbp_1 _16525_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1319),
    .D(_01972_),
    .Q_N(_05339_),
    .Q(\mem.mem[234][5] ));
 sg13g2_dfrbp_1 _16526_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1318),
    .D(_01973_),
    .Q_N(_05338_),
    .Q(\mem.mem[234][6] ));
 sg13g2_dfrbp_1 _16527_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1317),
    .D(_01974_),
    .Q_N(_05337_),
    .Q(\mem.mem[234][7] ));
 sg13g2_dfrbp_1 _16528_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1316),
    .D(_01975_),
    .Q_N(_05336_),
    .Q(\mem.mem[235][0] ));
 sg13g2_dfrbp_1 _16529_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1315),
    .D(_01976_),
    .Q_N(_05335_),
    .Q(\mem.mem[235][1] ));
 sg13g2_dfrbp_1 _16530_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1314),
    .D(_01977_),
    .Q_N(_05334_),
    .Q(\mem.mem[235][2] ));
 sg13g2_dfrbp_1 _16531_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1313),
    .D(_01978_),
    .Q_N(_05333_),
    .Q(\mem.mem[235][3] ));
 sg13g2_dfrbp_1 _16532_ (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1312),
    .D(_01979_),
    .Q_N(_05332_),
    .Q(\mem.mem[235][4] ));
 sg13g2_dfrbp_1 _16533_ (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1311),
    .D(_01980_),
    .Q_N(_05331_),
    .Q(\mem.mem[235][5] ));
 sg13g2_dfrbp_1 _16534_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1310),
    .D(_01981_),
    .Q_N(_05330_),
    .Q(\mem.mem[235][6] ));
 sg13g2_dfrbp_1 _16535_ (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1309),
    .D(_01982_),
    .Q_N(_05329_),
    .Q(\mem.mem[235][7] ));
 sg13g2_dfrbp_1 _16536_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1308),
    .D(_01983_),
    .Q_N(_05328_),
    .Q(\mem.mem[236][0] ));
 sg13g2_dfrbp_1 _16537_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1307),
    .D(_01984_),
    .Q_N(_05327_),
    .Q(\mem.mem[236][1] ));
 sg13g2_dfrbp_1 _16538_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1306),
    .D(_01985_),
    .Q_N(_05326_),
    .Q(\mem.mem[236][2] ));
 sg13g2_dfrbp_1 _16539_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1305),
    .D(_01986_),
    .Q_N(_05325_),
    .Q(\mem.mem[236][3] ));
 sg13g2_dfrbp_1 _16540_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1304),
    .D(_01987_),
    .Q_N(_05324_),
    .Q(\mem.mem[236][4] ));
 sg13g2_dfrbp_1 _16541_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1303),
    .D(_01988_),
    .Q_N(_05323_),
    .Q(\mem.mem[236][5] ));
 sg13g2_dfrbp_1 _16542_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1302),
    .D(_01989_),
    .Q_N(_05322_),
    .Q(\mem.mem[236][6] ));
 sg13g2_dfrbp_1 _16543_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1301),
    .D(_01990_),
    .Q_N(_05321_),
    .Q(\mem.mem[236][7] ));
 sg13g2_dfrbp_1 _16544_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1300),
    .D(_01991_),
    .Q_N(_05320_),
    .Q(\mem.mem[237][0] ));
 sg13g2_dfrbp_1 _16545_ (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1299),
    .D(_01992_),
    .Q_N(_05319_),
    .Q(\mem.mem[237][1] ));
 sg13g2_dfrbp_1 _16546_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1298),
    .D(_01993_),
    .Q_N(_05318_),
    .Q(\mem.mem[237][2] ));
 sg13g2_dfrbp_1 _16547_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1297),
    .D(_01994_),
    .Q_N(_05317_),
    .Q(\mem.mem[237][3] ));
 sg13g2_dfrbp_1 _16548_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1296),
    .D(_01995_),
    .Q_N(_05316_),
    .Q(\mem.mem[237][4] ));
 sg13g2_dfrbp_1 _16549_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1295),
    .D(_01996_),
    .Q_N(_05315_),
    .Q(\mem.mem[237][5] ));
 sg13g2_dfrbp_1 _16550_ (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1294),
    .D(_01997_),
    .Q_N(_05314_),
    .Q(\mem.mem[237][6] ));
 sg13g2_dfrbp_1 _16551_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1293),
    .D(_01998_),
    .Q_N(_05313_),
    .Q(\mem.mem[237][7] ));
 sg13g2_dfrbp_1 _16552_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1292),
    .D(_01999_),
    .Q_N(_05312_),
    .Q(\mem.mem[238][0] ));
 sg13g2_dfrbp_1 _16553_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1291),
    .D(_02000_),
    .Q_N(_05311_),
    .Q(\mem.mem[238][1] ));
 sg13g2_dfrbp_1 _16554_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1290),
    .D(_02001_),
    .Q_N(_05310_),
    .Q(\mem.mem[238][2] ));
 sg13g2_dfrbp_1 _16555_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1289),
    .D(_02002_),
    .Q_N(_05309_),
    .Q(\mem.mem[238][3] ));
 sg13g2_dfrbp_1 _16556_ (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1288),
    .D(_02003_),
    .Q_N(_05308_),
    .Q(\mem.mem[238][4] ));
 sg13g2_dfrbp_1 _16557_ (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1287),
    .D(_02004_),
    .Q_N(_05307_),
    .Q(\mem.mem[238][5] ));
 sg13g2_dfrbp_1 _16558_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1286),
    .D(_02005_),
    .Q_N(_05306_),
    .Q(\mem.mem[238][6] ));
 sg13g2_dfrbp_1 _16559_ (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1285),
    .D(_02006_),
    .Q_N(_05305_),
    .Q(\mem.mem[238][7] ));
 sg13g2_dfrbp_1 _16560_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1284),
    .D(_02007_),
    .Q_N(_05304_),
    .Q(\mem.mem[23][0] ));
 sg13g2_dfrbp_1 _16561_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1283),
    .D(_02008_),
    .Q_N(_05303_),
    .Q(\mem.mem[23][1] ));
 sg13g2_dfrbp_1 _16562_ (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1282),
    .D(_02009_),
    .Q_N(_05302_),
    .Q(\mem.mem[23][2] ));
 sg13g2_dfrbp_1 _16563_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1281),
    .D(_02010_),
    .Q_N(_05301_),
    .Q(\mem.mem[23][3] ));
 sg13g2_dfrbp_1 _16564_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1280),
    .D(_02011_),
    .Q_N(_05300_),
    .Q(\mem.mem[23][4] ));
 sg13g2_dfrbp_1 _16565_ (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1279),
    .D(_02012_),
    .Q_N(_05299_),
    .Q(\mem.mem[23][5] ));
 sg13g2_dfrbp_1 _16566_ (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1278),
    .D(_02013_),
    .Q_N(_05298_),
    .Q(\mem.mem[23][6] ));
 sg13g2_dfrbp_1 _16567_ (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1277),
    .D(_02014_),
    .Q_N(_05297_),
    .Q(\mem.mem[23][7] ));
 sg13g2_dfrbp_1 _16568_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1276),
    .D(_02015_),
    .Q_N(_05296_),
    .Q(\mem.mem[240][0] ));
 sg13g2_dfrbp_1 _16569_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1275),
    .D(_02016_),
    .Q_N(_05295_),
    .Q(\mem.mem[240][1] ));
 sg13g2_dfrbp_1 _16570_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1274),
    .D(_02017_),
    .Q_N(_05294_),
    .Q(\mem.mem[240][2] ));
 sg13g2_dfrbp_1 _16571_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1273),
    .D(_02018_),
    .Q_N(_05293_),
    .Q(\mem.mem[240][3] ));
 sg13g2_dfrbp_1 _16572_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1272),
    .D(_02019_),
    .Q_N(_05292_),
    .Q(\mem.mem[240][4] ));
 sg13g2_dfrbp_1 _16573_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1271),
    .D(_02020_),
    .Q_N(_05291_),
    .Q(\mem.mem[240][5] ));
 sg13g2_dfrbp_1 _16574_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1270),
    .D(_02021_),
    .Q_N(_05290_),
    .Q(\mem.mem[240][6] ));
 sg13g2_dfrbp_1 _16575_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1269),
    .D(_02022_),
    .Q_N(_05289_),
    .Q(\mem.mem[240][7] ));
 sg13g2_dfrbp_1 _16576_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1268),
    .D(_02023_),
    .Q_N(_05288_),
    .Q(\mem.mem[241][0] ));
 sg13g2_dfrbp_1 _16577_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1267),
    .D(_02024_),
    .Q_N(_05287_),
    .Q(\mem.mem[241][1] ));
 sg13g2_dfrbp_1 _16578_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1266),
    .D(_02025_),
    .Q_N(_05286_),
    .Q(\mem.mem[241][2] ));
 sg13g2_dfrbp_1 _16579_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1265),
    .D(_02026_),
    .Q_N(_05285_),
    .Q(\mem.mem[241][3] ));
 sg13g2_dfrbp_1 _16580_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1264),
    .D(_02027_),
    .Q_N(_05284_),
    .Q(\mem.mem[241][4] ));
 sg13g2_dfrbp_1 _16581_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1263),
    .D(_02028_),
    .Q_N(_05283_),
    .Q(\mem.mem[241][5] ));
 sg13g2_dfrbp_1 _16582_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1262),
    .D(_02029_),
    .Q_N(_05282_),
    .Q(\mem.mem[241][6] ));
 sg13g2_dfrbp_1 _16583_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1261),
    .D(_02030_),
    .Q_N(_05281_),
    .Q(\mem.mem[241][7] ));
 sg13g2_dfrbp_1 _16584_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1260),
    .D(_02031_),
    .Q_N(_05280_),
    .Q(\mem.mem[242][0] ));
 sg13g2_dfrbp_1 _16585_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1259),
    .D(_02032_),
    .Q_N(_05279_),
    .Q(\mem.mem[242][1] ));
 sg13g2_dfrbp_1 _16586_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1258),
    .D(_02033_),
    .Q_N(_05278_),
    .Q(\mem.mem[242][2] ));
 sg13g2_dfrbp_1 _16587_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1257),
    .D(_02034_),
    .Q_N(_05277_),
    .Q(\mem.mem[242][3] ));
 sg13g2_dfrbp_1 _16588_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1256),
    .D(_02035_),
    .Q_N(_05276_),
    .Q(\mem.mem[242][4] ));
 sg13g2_dfrbp_1 _16589_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1255),
    .D(_02036_),
    .Q_N(_05275_),
    .Q(\mem.mem[242][5] ));
 sg13g2_dfrbp_1 _16590_ (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1254),
    .D(_02037_),
    .Q_N(_05274_),
    .Q(\mem.mem[242][6] ));
 sg13g2_dfrbp_1 _16591_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1253),
    .D(_02038_),
    .Q_N(_05273_),
    .Q(\mem.mem[242][7] ));
 sg13g2_dfrbp_1 _16592_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1252),
    .D(_02039_),
    .Q_N(_05272_),
    .Q(\mem.mem[243][0] ));
 sg13g2_dfrbp_1 _16593_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1251),
    .D(_02040_),
    .Q_N(_05271_),
    .Q(\mem.mem[243][1] ));
 sg13g2_dfrbp_1 _16594_ (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1250),
    .D(_02041_),
    .Q_N(_05270_),
    .Q(\mem.mem[243][2] ));
 sg13g2_dfrbp_1 _16595_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1249),
    .D(_02042_),
    .Q_N(_05269_),
    .Q(\mem.mem[243][3] ));
 sg13g2_dfrbp_1 _16596_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1248),
    .D(_02043_),
    .Q_N(_05268_),
    .Q(\mem.mem[243][4] ));
 sg13g2_dfrbp_1 _16597_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1247),
    .D(_02044_),
    .Q_N(_05267_),
    .Q(\mem.mem[243][5] ));
 sg13g2_dfrbp_1 _16598_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1246),
    .D(_02045_),
    .Q_N(_05266_),
    .Q(\mem.mem[243][6] ));
 sg13g2_dfrbp_1 _16599_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1245),
    .D(_02046_),
    .Q_N(_05265_),
    .Q(\mem.mem[243][7] ));
 sg13g2_dfrbp_1 _16600_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1244),
    .D(_02047_),
    .Q_N(_05264_),
    .Q(\mem.mem[244][0] ));
 sg13g2_dfrbp_1 _16601_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1243),
    .D(_02048_),
    .Q_N(_05263_),
    .Q(\mem.mem[244][1] ));
 sg13g2_dfrbp_1 _16602_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1242),
    .D(_02049_),
    .Q_N(_05262_),
    .Q(\mem.mem[244][2] ));
 sg13g2_dfrbp_1 _16603_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1241),
    .D(_02050_),
    .Q_N(_05261_),
    .Q(\mem.mem[244][3] ));
 sg13g2_dfrbp_1 _16604_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1240),
    .D(_02051_),
    .Q_N(_05260_),
    .Q(\mem.mem[244][4] ));
 sg13g2_dfrbp_1 _16605_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1239),
    .D(_02052_),
    .Q_N(_05259_),
    .Q(\mem.mem[244][5] ));
 sg13g2_dfrbp_1 _16606_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net661),
    .D(_02053_),
    .Q_N(_05258_),
    .Q(\mem.mem[244][6] ));
 sg13g2_dfrbp_1 _16607_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net659),
    .D(_02054_),
    .Q_N(_05257_),
    .Q(\mem.mem[244][7] ));
 sg13g2_dfrbp_1 _16608_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net657),
    .D(_02055_),
    .Q_N(_05256_),
    .Q(\mem.mem[245][0] ));
 sg13g2_dfrbp_1 _16609_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net655),
    .D(_02056_),
    .Q_N(_05255_),
    .Q(\mem.mem[245][1] ));
 sg13g2_dfrbp_1 _16610_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net653),
    .D(_02057_),
    .Q_N(_05254_),
    .Q(\mem.mem[245][2] ));
 sg13g2_dfrbp_1 _16611_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net651),
    .D(_02058_),
    .Q_N(_05253_),
    .Q(\mem.mem[245][3] ));
 sg13g2_dfrbp_1 _16612_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net649),
    .D(_02059_),
    .Q_N(_05252_),
    .Q(\mem.mem[245][4] ));
 sg13g2_dfrbp_1 _16613_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net647),
    .D(_02060_),
    .Q_N(_05251_),
    .Q(\mem.mem[245][5] ));
 sg13g2_dfrbp_1 _16614_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net645),
    .D(_02061_),
    .Q_N(_05250_),
    .Q(\mem.mem[245][6] ));
 sg13g2_dfrbp_1 _16615_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net643),
    .D(_02062_),
    .Q_N(_05249_),
    .Q(\mem.mem[245][7] ));
 sg13g2_dfrbp_1 _16616_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net641),
    .D(_02063_),
    .Q_N(_05248_),
    .Q(\mem.mem[246][0] ));
 sg13g2_dfrbp_1 _16617_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net639),
    .D(_02064_),
    .Q_N(_05247_),
    .Q(\mem.mem[246][1] ));
 sg13g2_dfrbp_1 _16618_ (.CLK(clknet_leaf_249_clk),
    .RESET_B(net637),
    .D(_02065_),
    .Q_N(_05246_),
    .Q(\mem.mem[246][2] ));
 sg13g2_dfrbp_1 _16619_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net635),
    .D(_02066_),
    .Q_N(_05245_),
    .Q(\mem.mem[246][3] ));
 sg13g2_dfrbp_1 _16620_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net633),
    .D(_02067_),
    .Q_N(_05244_),
    .Q(\mem.mem[246][4] ));
 sg13g2_dfrbp_1 _16621_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net631),
    .D(_02068_),
    .Q_N(_05243_),
    .Q(\mem.mem[246][5] ));
 sg13g2_dfrbp_1 _16622_ (.CLK(clknet_leaf_245_clk),
    .RESET_B(net629),
    .D(_02069_),
    .Q_N(_05242_),
    .Q(\mem.mem[246][6] ));
 sg13g2_dfrbp_1 _16623_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net627),
    .D(_02070_),
    .Q_N(_05241_),
    .Q(\mem.mem[246][7] ));
 sg13g2_dfrbp_1 _16624_ (.CLK(clknet_leaf_247_clk),
    .RESET_B(net625),
    .D(_02071_),
    .Q_N(_05240_),
    .Q(\mem.mem[247][0] ));
 sg13g2_dfrbp_1 _16625_ (.CLK(clknet_leaf_246_clk),
    .RESET_B(net623),
    .D(_02072_),
    .Q_N(_05239_),
    .Q(\mem.mem[247][1] ));
 sg13g2_dfrbp_1 _16626_ (.CLK(clknet_leaf_250_clk),
    .RESET_B(net621),
    .D(_02073_),
    .Q_N(_05238_),
    .Q(\mem.mem[247][2] ));
 sg13g2_dfrbp_1 _16627_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net619),
    .D(_02074_),
    .Q_N(_05237_),
    .Q(\mem.mem[247][3] ));
 sg13g2_dfrbp_1 _16628_ (.CLK(clknet_leaf_251_clk),
    .RESET_B(net617),
    .D(_02075_),
    .Q_N(_05236_),
    .Q(\mem.mem[247][4] ));
 sg13g2_dfrbp_1 _16629_ (.CLK(clknet_leaf_241_clk),
    .RESET_B(net615),
    .D(_02076_),
    .Q_N(_05235_),
    .Q(\mem.mem[247][5] ));
 sg13g2_dfrbp_1 _16630_ (.CLK(clknet_leaf_244_clk),
    .RESET_B(net613),
    .D(_02077_),
    .Q_N(_05234_),
    .Q(\mem.mem[247][6] ));
 sg13g2_dfrbp_1 _16631_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net611),
    .D(_02078_),
    .Q_N(_05233_),
    .Q(\mem.mem[247][7] ));
 sg13g2_dfrbp_1 _16632_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net609),
    .D(_02079_),
    .Q_N(_05232_),
    .Q(\mem.mem[248][0] ));
 sg13g2_dfrbp_1 _16633_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net607),
    .D(_02080_),
    .Q_N(_05231_),
    .Q(\mem.mem[248][1] ));
 sg13g2_dfrbp_1 _16634_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net605),
    .D(_02081_),
    .Q_N(_05230_),
    .Q(\mem.mem[248][2] ));
 sg13g2_dfrbp_1 _16635_ (.CLK(clknet_leaf_252_clk),
    .RESET_B(net603),
    .D(_02082_),
    .Q_N(_05229_),
    .Q(\mem.mem[248][3] ));
 sg13g2_dfrbp_1 _16636_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net601),
    .D(_02083_),
    .Q_N(_05228_),
    .Q(\mem.mem[248][4] ));
 sg13g2_dfrbp_1 _16637_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net599),
    .D(_02084_),
    .Q_N(_05227_),
    .Q(\mem.mem[248][5] ));
 sg13g2_dfrbp_1 _16638_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net597),
    .D(_02085_),
    .Q_N(_05226_),
    .Q(\mem.mem[248][6] ));
 sg13g2_dfrbp_1 _16639_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net595),
    .D(_02086_),
    .Q_N(_05225_),
    .Q(\mem.mem[248][7] ));
 sg13g2_dfrbp_1 _16640_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net593),
    .D(_02087_),
    .Q_N(_05224_),
    .Q(\mem.mem[24][0] ));
 sg13g2_dfrbp_1 _16641_ (.CLK(clknet_leaf_190_clk),
    .RESET_B(net591),
    .D(_02088_),
    .Q_N(_05223_),
    .Q(\mem.mem[24][1] ));
 sg13g2_dfrbp_1 _16642_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net589),
    .D(_02089_),
    .Q_N(_05222_),
    .Q(\mem.mem[24][2] ));
 sg13g2_dfrbp_1 _16643_ (.CLK(clknet_leaf_192_clk),
    .RESET_B(net587),
    .D(_02090_),
    .Q_N(_05221_),
    .Q(\mem.mem[24][3] ));
 sg13g2_dfrbp_1 _16644_ (.CLK(clknet_leaf_189_clk),
    .RESET_B(net585),
    .D(_02091_),
    .Q_N(_05220_),
    .Q(\mem.mem[24][4] ));
 sg13g2_dfrbp_1 _16645_ (.CLK(clknet_leaf_188_clk),
    .RESET_B(net583),
    .D(_02092_),
    .Q_N(_05219_),
    .Q(\mem.mem[24][5] ));
 sg13g2_dfrbp_1 _16646_ (.CLK(clknet_leaf_181_clk),
    .RESET_B(net581),
    .D(_02093_),
    .Q_N(_05218_),
    .Q(\mem.mem[24][6] ));
 sg13g2_dfrbp_1 _16647_ (.CLK(clknet_leaf_182_clk),
    .RESET_B(net579),
    .D(_02094_),
    .Q_N(_05217_),
    .Q(\mem.mem[24][7] ));
 sg13g2_dfrbp_1 _16648_ (.CLK(clknet_leaf_235_clk),
    .RESET_B(net577),
    .D(_02095_),
    .Q_N(_05216_),
    .Q(\mem.mem[250][0] ));
 sg13g2_dfrbp_1 _16649_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net575),
    .D(_02096_),
    .Q_N(_05215_),
    .Q(\mem.mem[250][1] ));
 sg13g2_dfrbp_1 _16650_ (.CLK(clknet_leaf_26_clk),
    .RESET_B(net573),
    .D(_02097_),
    .Q_N(_05214_),
    .Q(\mem.mem[250][2] ));
 sg13g2_dfrbp_1 _16651_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net571),
    .D(_02098_),
    .Q_N(_05213_),
    .Q(\mem.mem[250][3] ));
 sg13g2_dfrbp_1 _16652_ (.CLK(clknet_leaf_236_clk),
    .RESET_B(net569),
    .D(_02099_),
    .Q_N(_05212_),
    .Q(\mem.mem[250][4] ));
 sg13g2_dfrbp_1 _16653_ (.CLK(clknet_leaf_233_clk),
    .RESET_B(net567),
    .D(_02100_),
    .Q_N(_05211_),
    .Q(\mem.mem[250][5] ));
 sg13g2_dfrbp_1 _16654_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net565),
    .D(_02101_),
    .Q_N(_05210_),
    .Q(\mem.mem[250][6] ));
 sg13g2_dfrbp_1 _16655_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net563),
    .D(_02102_),
    .Q_N(_05209_),
    .Q(\mem.mem[250][7] ));
 sg13g2_dfrbp_1 _16656_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net561),
    .D(_02103_),
    .Q_N(_05208_),
    .Q(\mem.mem[251][0] ));
 sg13g2_dfrbp_1 _16657_ (.CLK(clknet_leaf_238_clk),
    .RESET_B(net559),
    .D(_02104_),
    .Q_N(_05207_),
    .Q(\mem.mem[251][1] ));
 sg13g2_dfrbp_1 _16658_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net557),
    .D(_02105_),
    .Q_N(_05206_),
    .Q(\mem.mem[251][2] ));
 sg13g2_dfrbp_1 _16659_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net555),
    .D(_02106_),
    .Q_N(_05205_),
    .Q(\mem.mem[251][3] ));
 sg13g2_dfrbp_1 _16660_ (.CLK(clknet_leaf_237_clk),
    .RESET_B(net553),
    .D(_02107_),
    .Q_N(_05204_),
    .Q(\mem.mem[251][4] ));
 sg13g2_dfrbp_1 _16661_ (.CLK(clknet_leaf_234_clk),
    .RESET_B(net551),
    .D(_02108_),
    .Q_N(_05203_),
    .Q(\mem.mem[251][5] ));
 sg13g2_dfrbp_1 _16662_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net549),
    .D(_02109_),
    .Q_N(_05202_),
    .Q(\mem.mem[251][6] ));
 sg13g2_dfrbp_1 _16663_ (.CLK(clknet_leaf_232_clk),
    .RESET_B(net547),
    .D(_02110_),
    .Q_N(_05201_),
    .Q(\mem.mem[251][7] ));
 sg13g2_dfrbp_1 _16664_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net545),
    .D(_02111_),
    .Q_N(_05200_),
    .Q(\mem.mem[9][0] ));
 sg13g2_dfrbp_1 _16665_ (.CLK(clknet_leaf_218_clk),
    .RESET_B(net359),
    .D(_02112_),
    .Q_N(_05199_),
    .Q(\mem.mem[9][1] ));
 sg13g2_dfrbp_1 _16666_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net357),
    .D(_02113_),
    .Q_N(_05198_),
    .Q(\mem.mem[9][2] ));
 sg13g2_dfrbp_1 _16667_ (.CLK(clknet_leaf_217_clk),
    .RESET_B(net355),
    .D(_02114_),
    .Q_N(_05197_),
    .Q(\mem.mem[9][3] ));
 sg13g2_dfrbp_1 _16668_ (.CLK(clknet_leaf_202_clk),
    .RESET_B(net353),
    .D(_02115_),
    .Q_N(_05196_),
    .Q(\mem.mem[9][4] ));
 sg13g2_dfrbp_1 _16669_ (.CLK(clknet_leaf_168_clk),
    .RESET_B(net351),
    .D(_02116_),
    .Q_N(_05195_),
    .Q(\mem.mem[9][5] ));
 sg13g2_dfrbp_1 _16670_ (.CLK(clknet_leaf_220_clk),
    .RESET_B(net349),
    .D(_02117_),
    .Q_N(_05194_),
    .Q(\mem.mem[9][6] ));
 sg13g2_dfrbp_1 _16671_ (.CLK(clknet_leaf_219_clk),
    .RESET_B(net347),
    .D(_02118_),
    .Q_N(_05193_),
    .Q(\mem.mem[9][7] ));
 sg13g2_dfrbp_1 _16672_ (.CLK(clknet_leaf_89_clk),
    .RESET_B(net345),
    .D(_02119_),
    .Q_N(_00008_),
    .Q(\mem.wr_en ));
 sg13g2_tiehi _15715__27 (.L_HI(net27));
 sg13g2_tiehi _15714__28 (.L_HI(net28));
 sg13g2_tiehi _15713__29 (.L_HI(net29));
 sg13g2_tiehi _15712__30 (.L_HI(net30));
 sg13g2_tiehi _15711__31 (.L_HI(net31));
 sg13g2_tiehi _15710__32 (.L_HI(net32));
 sg13g2_tiehi _15709__33 (.L_HI(net33));
 sg13g2_tiehi _15708__34 (.L_HI(net34));
 sg13g2_tiehi _15707__35 (.L_HI(net35));
 sg13g2_tiehi _15706__36 (.L_HI(net36));
 sg13g2_tiehi _15705__37 (.L_HI(net37));
 sg13g2_tiehi _15704__38 (.L_HI(net38));
 sg13g2_tiehi _15703__39 (.L_HI(net39));
 sg13g2_tiehi _15702__40 (.L_HI(net40));
 sg13g2_tiehi _15701__41 (.L_HI(net41));
 sg13g2_tiehi _15700__42 (.L_HI(net42));
 sg13g2_tiehi _15699__43 (.L_HI(net43));
 sg13g2_tiehi _15698__44 (.L_HI(net44));
 sg13g2_tiehi _15697__45 (.L_HI(net45));
 sg13g2_tiehi _15696__46 (.L_HI(net46));
 sg13g2_tiehi _15695__47 (.L_HI(net47));
 sg13g2_tiehi _15694__48 (.L_HI(net48));
 sg13g2_tiehi _15693__49 (.L_HI(net49));
 sg13g2_tiehi _15692__50 (.L_HI(net50));
 sg13g2_tiehi _15691__51 (.L_HI(net51));
 sg13g2_tiehi _15690__52 (.L_HI(net52));
 sg13g2_tiehi _15689__53 (.L_HI(net53));
 sg13g2_tiehi _15688__54 (.L_HI(net54));
 sg13g2_tiehi _15687__55 (.L_HI(net55));
 sg13g2_tiehi _15686__56 (.L_HI(net56));
 sg13g2_tiehi _15685__57 (.L_HI(net57));
 sg13g2_tiehi _15684__58 (.L_HI(net58));
 sg13g2_tiehi _15683__59 (.L_HI(net59));
 sg13g2_tiehi _15682__60 (.L_HI(net60));
 sg13g2_tiehi _15681__61 (.L_HI(net61));
 sg13g2_tiehi _15680__62 (.L_HI(net62));
 sg13g2_tiehi _15679__63 (.L_HI(net63));
 sg13g2_tiehi _15678__64 (.L_HI(net64));
 sg13g2_tiehi _15677__65 (.L_HI(net65));
 sg13g2_tiehi _15676__66 (.L_HI(net66));
 sg13g2_tiehi _15675__67 (.L_HI(net67));
 sg13g2_tiehi _15674__68 (.L_HI(net68));
 sg13g2_tiehi _15673__69 (.L_HI(net69));
 sg13g2_tiehi _15672__70 (.L_HI(net70));
 sg13g2_tiehi _15671__71 (.L_HI(net71));
 sg13g2_tiehi _15670__72 (.L_HI(net72));
 sg13g2_tiehi _15669__73 (.L_HI(net73));
 sg13g2_tiehi _15668__74 (.L_HI(net74));
 sg13g2_tiehi _15667__75 (.L_HI(net75));
 sg13g2_tiehi _15666__76 (.L_HI(net76));
 sg13g2_tiehi _15665__77 (.L_HI(net77));
 sg13g2_tiehi _15664__78 (.L_HI(net78));
 sg13g2_tiehi _15663__79 (.L_HI(net79));
 sg13g2_tiehi _15662__80 (.L_HI(net80));
 sg13g2_tiehi _15661__81 (.L_HI(net81));
 sg13g2_tiehi _15660__82 (.L_HI(net82));
 sg13g2_tiehi _15659__83 (.L_HI(net83));
 sg13g2_tiehi _15658__84 (.L_HI(net84));
 sg13g2_tiehi _15657__85 (.L_HI(net85));
 sg13g2_tiehi _15656__86 (.L_HI(net86));
 sg13g2_tiehi _15655__87 (.L_HI(net87));
 sg13g2_tiehi _15654__88 (.L_HI(net88));
 sg13g2_tiehi _15653__89 (.L_HI(net89));
 sg13g2_tiehi _15652__90 (.L_HI(net90));
 sg13g2_tiehi _15651__91 (.L_HI(net91));
 sg13g2_tiehi _15650__92 (.L_HI(net92));
 sg13g2_tiehi _15649__93 (.L_HI(net93));
 sg13g2_tiehi _15648__94 (.L_HI(net94));
 sg13g2_tiehi _15647__95 (.L_HI(net95));
 sg13g2_tiehi _15646__96 (.L_HI(net96));
 sg13g2_tiehi _15645__97 (.L_HI(net97));
 sg13g2_tiehi _15644__98 (.L_HI(net98));
 sg13g2_tiehi _15643__99 (.L_HI(net99));
 sg13g2_tiehi _15642__100 (.L_HI(net100));
 sg13g2_tiehi _15641__101 (.L_HI(net101));
 sg13g2_tiehi _15640__102 (.L_HI(net102));
 sg13g2_tiehi _15639__103 (.L_HI(net103));
 sg13g2_tiehi _15638__104 (.L_HI(net104));
 sg13g2_tiehi _15637__105 (.L_HI(net105));
 sg13g2_tiehi _15636__106 (.L_HI(net106));
 sg13g2_tiehi _15635__107 (.L_HI(net107));
 sg13g2_tiehi _15634__108 (.L_HI(net108));
 sg13g2_tiehi _15633__109 (.L_HI(net109));
 sg13g2_tiehi _15632__110 (.L_HI(net110));
 sg13g2_tiehi _15631__111 (.L_HI(net111));
 sg13g2_tiehi _15630__112 (.L_HI(net112));
 sg13g2_tiehi _15629__113 (.L_HI(net113));
 sg13g2_tiehi _15628__114 (.L_HI(net114));
 sg13g2_tiehi _15627__115 (.L_HI(net115));
 sg13g2_tiehi _15626__116 (.L_HI(net116));
 sg13g2_tiehi _15625__117 (.L_HI(net117));
 sg13g2_tiehi _15624__118 (.L_HI(net118));
 sg13g2_tiehi _15623__119 (.L_HI(net119));
 sg13g2_tiehi _15622__120 (.L_HI(net120));
 sg13g2_tiehi _15621__121 (.L_HI(net121));
 sg13g2_tiehi _15620__122 (.L_HI(net122));
 sg13g2_tiehi _15619__123 (.L_HI(net123));
 sg13g2_tiehi _15618__124 (.L_HI(net124));
 sg13g2_tiehi _15617__125 (.L_HI(net125));
 sg13g2_tiehi _15616__126 (.L_HI(net126));
 sg13g2_tiehi _15615__127 (.L_HI(net127));
 sg13g2_tiehi _15614__128 (.L_HI(net128));
 sg13g2_tiehi _15613__129 (.L_HI(net129));
 sg13g2_tiehi _15612__130 (.L_HI(net130));
 sg13g2_tiehi _15611__131 (.L_HI(net131));
 sg13g2_tiehi _15610__132 (.L_HI(net132));
 sg13g2_tiehi _15609__133 (.L_HI(net133));
 sg13g2_tiehi _15608__134 (.L_HI(net134));
 sg13g2_tiehi _15607__135 (.L_HI(net135));
 sg13g2_tiehi _15606__136 (.L_HI(net136));
 sg13g2_tiehi _15605__137 (.L_HI(net137));
 sg13g2_tiehi _15604__138 (.L_HI(net138));
 sg13g2_tiehi _15603__139 (.L_HI(net139));
 sg13g2_tiehi _15602__140 (.L_HI(net140));
 sg13g2_tiehi _15601__141 (.L_HI(net141));
 sg13g2_tiehi _15600__142 (.L_HI(net142));
 sg13g2_tiehi _15599__143 (.L_HI(net143));
 sg13g2_tiehi _15598__144 (.L_HI(net144));
 sg13g2_tiehi _15597__145 (.L_HI(net145));
 sg13g2_tiehi _15596__146 (.L_HI(net146));
 sg13g2_tiehi _15595__147 (.L_HI(net147));
 sg13g2_tiehi _15594__148 (.L_HI(net148));
 sg13g2_tiehi _15593__149 (.L_HI(net149));
 sg13g2_tiehi _15592__150 (.L_HI(net150));
 sg13g2_tiehi _15591__151 (.L_HI(net151));
 sg13g2_tiehi _15590__152 (.L_HI(net152));
 sg13g2_tiehi _15589__153 (.L_HI(net153));
 sg13g2_tiehi _15588__154 (.L_HI(net154));
 sg13g2_tiehi _15587__155 (.L_HI(net155));
 sg13g2_tiehi _15586__156 (.L_HI(net156));
 sg13g2_tiehi _15585__157 (.L_HI(net157));
 sg13g2_tiehi _15584__158 (.L_HI(net158));
 sg13g2_tiehi _15583__159 (.L_HI(net159));
 sg13g2_tiehi _15582__160 (.L_HI(net160));
 sg13g2_tiehi _15581__161 (.L_HI(net161));
 sg13g2_tiehi _15580__162 (.L_HI(net162));
 sg13g2_tiehi _15579__163 (.L_HI(net163));
 sg13g2_tiehi _15578__164 (.L_HI(net164));
 sg13g2_tiehi _15577__165 (.L_HI(net165));
 sg13g2_tiehi _15576__166 (.L_HI(net166));
 sg13g2_tiehi _15575__167 (.L_HI(net167));
 sg13g2_tiehi _15574__168 (.L_HI(net168));
 sg13g2_tiehi _15573__169 (.L_HI(net169));
 sg13g2_tiehi _15572__170 (.L_HI(net170));
 sg13g2_tiehi _15571__171 (.L_HI(net171));
 sg13g2_tiehi _15570__172 (.L_HI(net172));
 sg13g2_tiehi _15569__173 (.L_HI(net173));
 sg13g2_tiehi _15568__174 (.L_HI(net174));
 sg13g2_tiehi _15567__175 (.L_HI(net175));
 sg13g2_tiehi _15566__176 (.L_HI(net176));
 sg13g2_tiehi _15565__177 (.L_HI(net177));
 sg13g2_tiehi _15564__178 (.L_HI(net178));
 sg13g2_tiehi _15563__179 (.L_HI(net179));
 sg13g2_tiehi _15562__180 (.L_HI(net180));
 sg13g2_tiehi _15561__181 (.L_HI(net181));
 sg13g2_tiehi _15560__182 (.L_HI(net182));
 sg13g2_tiehi _15559__183 (.L_HI(net183));
 sg13g2_tiehi _15558__184 (.L_HI(net184));
 sg13g2_tiehi _15557__185 (.L_HI(net185));
 sg13g2_tiehi _15556__186 (.L_HI(net186));
 sg13g2_tiehi _15555__187 (.L_HI(net187));
 sg13g2_tiehi _15554__188 (.L_HI(net188));
 sg13g2_tiehi _15553__189 (.L_HI(net189));
 sg13g2_tiehi _15552__190 (.L_HI(net190));
 sg13g2_tiehi _15551__191 (.L_HI(net191));
 sg13g2_tiehi _15550__192 (.L_HI(net192));
 sg13g2_tiehi _15549__193 (.L_HI(net193));
 sg13g2_tiehi _15548__194 (.L_HI(net194));
 sg13g2_tiehi _15547__195 (.L_HI(net195));
 sg13g2_tiehi _15546__196 (.L_HI(net196));
 sg13g2_tiehi _15545__197 (.L_HI(net197));
 sg13g2_tiehi _15544__198 (.L_HI(net198));
 sg13g2_tiehi _15543__199 (.L_HI(net199));
 sg13g2_tiehi _15542__200 (.L_HI(net200));
 sg13g2_tiehi _15541__201 (.L_HI(net201));
 sg13g2_tiehi _15540__202 (.L_HI(net202));
 sg13g2_tiehi _15539__203 (.L_HI(net203));
 sg13g2_tiehi _15538__204 (.L_HI(net204));
 sg13g2_tiehi _15537__205 (.L_HI(net205));
 sg13g2_tiehi _15536__206 (.L_HI(net206));
 sg13g2_tiehi _15535__207 (.L_HI(net207));
 sg13g2_tiehi _15534__208 (.L_HI(net208));
 sg13g2_tiehi _15533__209 (.L_HI(net209));
 sg13g2_tiehi _15532__210 (.L_HI(net210));
 sg13g2_tiehi _15531__211 (.L_HI(net211));
 sg13g2_tiehi _15530__212 (.L_HI(net212));
 sg13g2_tiehi _15529__213 (.L_HI(net213));
 sg13g2_tiehi _15528__214 (.L_HI(net214));
 sg13g2_tiehi _15527__215 (.L_HI(net215));
 sg13g2_tiehi _15526__216 (.L_HI(net216));
 sg13g2_tiehi _15525__217 (.L_HI(net217));
 sg13g2_tiehi _15524__218 (.L_HI(net218));
 sg13g2_tiehi _15523__219 (.L_HI(net219));
 sg13g2_tiehi _15522__220 (.L_HI(net220));
 sg13g2_tiehi _15521__221 (.L_HI(net221));
 sg13g2_tiehi _15520__222 (.L_HI(net222));
 sg13g2_tiehi _15519__223 (.L_HI(net223));
 sg13g2_tiehi _15518__224 (.L_HI(net224));
 sg13g2_tiehi _15517__225 (.L_HI(net225));
 sg13g2_tiehi _15516__226 (.L_HI(net226));
 sg13g2_tiehi _15515__227 (.L_HI(net227));
 sg13g2_tiehi _15514__228 (.L_HI(net228));
 sg13g2_tiehi _15513__229 (.L_HI(net229));
 sg13g2_tiehi _15512__230 (.L_HI(net230));
 sg13g2_tiehi _15511__231 (.L_HI(net231));
 sg13g2_tiehi _15510__232 (.L_HI(net232));
 sg13g2_tiehi _15509__233 (.L_HI(net233));
 sg13g2_tiehi _15508__234 (.L_HI(net234));
 sg13g2_tiehi _15507__235 (.L_HI(net235));
 sg13g2_tiehi _15506__236 (.L_HI(net236));
 sg13g2_tiehi _15505__237 (.L_HI(net237));
 sg13g2_tiehi _15504__238 (.L_HI(net238));
 sg13g2_tiehi _15503__239 (.L_HI(net239));
 sg13g2_tiehi _15502__240 (.L_HI(net240));
 sg13g2_tiehi _15501__241 (.L_HI(net241));
 sg13g2_tiehi _15500__242 (.L_HI(net242));
 sg13g2_tiehi _15499__243 (.L_HI(net243));
 sg13g2_tiehi _15498__244 (.L_HI(net244));
 sg13g2_tiehi _15497__245 (.L_HI(net245));
 sg13g2_tiehi _15496__246 (.L_HI(net246));
 sg13g2_tiehi _15495__247 (.L_HI(net247));
 sg13g2_tiehi _15494__248 (.L_HI(net248));
 sg13g2_tiehi _15493__249 (.L_HI(net249));
 sg13g2_tiehi _15492__250 (.L_HI(net250));
 sg13g2_tiehi _15491__251 (.L_HI(net251));
 sg13g2_tiehi _15490__252 (.L_HI(net252));
 sg13g2_tiehi _15489__253 (.L_HI(net253));
 sg13g2_tiehi _15488__254 (.L_HI(net254));
 sg13g2_tiehi _15487__255 (.L_HI(net255));
 sg13g2_tiehi _15486__256 (.L_HI(net256));
 sg13g2_tiehi _15485__257 (.L_HI(net257));
 sg13g2_tiehi _15484__258 (.L_HI(net258));
 sg13g2_tiehi _15483__259 (.L_HI(net259));
 sg13g2_tiehi _15482__260 (.L_HI(net260));
 sg13g2_tiehi _15481__261 (.L_HI(net261));
 sg13g2_tiehi _15480__262 (.L_HI(net262));
 sg13g2_tiehi _15479__263 (.L_HI(net263));
 sg13g2_tiehi _15478__264 (.L_HI(net264));
 sg13g2_tiehi _15477__265 (.L_HI(net265));
 sg13g2_tiehi _15476__266 (.L_HI(net266));
 sg13g2_tiehi _15475__267 (.L_HI(net267));
 sg13g2_tiehi _15474__268 (.L_HI(net268));
 sg13g2_tiehi _15473__269 (.L_HI(net269));
 sg13g2_tiehi _15472__270 (.L_HI(net270));
 sg13g2_tiehi _15471__271 (.L_HI(net271));
 sg13g2_tiehi _15470__272 (.L_HI(net272));
 sg13g2_tiehi _15469__273 (.L_HI(net273));
 sg13g2_tiehi _15468__274 (.L_HI(net274));
 sg13g2_tiehi _15467__275 (.L_HI(net275));
 sg13g2_tiehi _15466__276 (.L_HI(net276));
 sg13g2_tiehi _15465__277 (.L_HI(net277));
 sg13g2_tiehi _15464__278 (.L_HI(net278));
 sg13g2_tiehi _15463__279 (.L_HI(net279));
 sg13g2_tiehi _15462__280 (.L_HI(net280));
 sg13g2_tiehi _15461__281 (.L_HI(net281));
 sg13g2_tiehi _15460__282 (.L_HI(net282));
 sg13g2_tiehi _15459__283 (.L_HI(net283));
 sg13g2_tiehi _15458__284 (.L_HI(net284));
 sg13g2_tiehi _15457__285 (.L_HI(net285));
 sg13g2_tiehi _15456__286 (.L_HI(net286));
 sg13g2_tiehi _15455__287 (.L_HI(net287));
 sg13g2_tiehi _15454__288 (.L_HI(net288));
 sg13g2_tiehi _15453__289 (.L_HI(net289));
 sg13g2_tiehi _15452__290 (.L_HI(net290));
 sg13g2_tiehi _15451__291 (.L_HI(net291));
 sg13g2_tiehi _15450__292 (.L_HI(net292));
 sg13g2_tiehi _15449__293 (.L_HI(net293));
 sg13g2_tiehi _15448__294 (.L_HI(net294));
 sg13g2_tiehi _15447__295 (.L_HI(net295));
 sg13g2_tiehi _15446__296 (.L_HI(net296));
 sg13g2_tiehi _15445__297 (.L_HI(net297));
 sg13g2_tiehi _15444__298 (.L_HI(net298));
 sg13g2_tiehi _15443__299 (.L_HI(net299));
 sg13g2_tiehi _15442__300 (.L_HI(net300));
 sg13g2_tiehi _15441__301 (.L_HI(net301));
 sg13g2_tiehi _15440__302 (.L_HI(net302));
 sg13g2_tiehi _15439__303 (.L_HI(net303));
 sg13g2_tiehi _15438__304 (.L_HI(net304));
 sg13g2_tiehi _15437__305 (.L_HI(net305));
 sg13g2_tiehi _15436__306 (.L_HI(net306));
 sg13g2_tiehi _15435__307 (.L_HI(net307));
 sg13g2_tiehi _15434__308 (.L_HI(net308));
 sg13g2_tiehi _15433__309 (.L_HI(net309));
 sg13g2_tiehi _15432__310 (.L_HI(net310));
 sg13g2_tiehi _15431__311 (.L_HI(net311));
 sg13g2_tiehi _15430__312 (.L_HI(net312));
 sg13g2_tiehi _15429__313 (.L_HI(net313));
 sg13g2_tiehi _15428__314 (.L_HI(net314));
 sg13g2_tiehi _15427__315 (.L_HI(net315));
 sg13g2_tiehi _15426__316 (.L_HI(net316));
 sg13g2_tiehi _15425__317 (.L_HI(net317));
 sg13g2_tiehi _15424__318 (.L_HI(net318));
 sg13g2_tiehi _15423__319 (.L_HI(net319));
 sg13g2_tiehi _15422__320 (.L_HI(net320));
 sg13g2_tiehi _15421__321 (.L_HI(net321));
 sg13g2_tiehi _15420__322 (.L_HI(net322));
 sg13g2_tiehi _15419__323 (.L_HI(net323));
 sg13g2_tiehi _15418__324 (.L_HI(net324));
 sg13g2_tiehi _15417__325 (.L_HI(net325));
 sg13g2_tiehi _15416__326 (.L_HI(net326));
 sg13g2_tiehi _15415__327 (.L_HI(net327));
 sg13g2_tiehi _15414__328 (.L_HI(net328));
 sg13g2_tiehi _15413__329 (.L_HI(net329));
 sg13g2_tiehi _15412__330 (.L_HI(net330));
 sg13g2_tiehi _15411__331 (.L_HI(net331));
 sg13g2_tiehi _15410__332 (.L_HI(net332));
 sg13g2_tiehi _15409__333 (.L_HI(net333));
 sg13g2_tiehi _15408__334 (.L_HI(net334));
 sg13g2_tiehi _15407__335 (.L_HI(net335));
 sg13g2_tiehi _15406__336 (.L_HI(net336));
 sg13g2_tiehi _15405__337 (.L_HI(net337));
 sg13g2_tiehi _15404__338 (.L_HI(net338));
 sg13g2_tiehi _15403__339 (.L_HI(net339));
 sg13g2_tiehi _15402__340 (.L_HI(net340));
 sg13g2_tiehi _15401__341 (.L_HI(net341));
 sg13g2_tiehi _15400__342 (.L_HI(net342));
 sg13g2_tiehi _14571__343 (.L_HI(net343));
 sg13g2_tiehi _15399__344 (.L_HI(net344));
 sg13g2_tiehi _16672__345 (.L_HI(net345));
 sg13g2_tiehi _15398__346 (.L_HI(net346));
 sg13g2_tiehi _16671__347 (.L_HI(net347));
 sg13g2_tiehi _15397__348 (.L_HI(net348));
 sg13g2_tiehi _16670__349 (.L_HI(net349));
 sg13g2_tiehi _15396__350 (.L_HI(net350));
 sg13g2_tiehi _16669__351 (.L_HI(net351));
 sg13g2_tiehi _15395__352 (.L_HI(net352));
 sg13g2_tiehi _16668__353 (.L_HI(net353));
 sg13g2_tiehi _15394__354 (.L_HI(net354));
 sg13g2_tiehi _16667__355 (.L_HI(net355));
 sg13g2_tiehi _15393__356 (.L_HI(net356));
 sg13g2_tiehi _16666__357 (.L_HI(net357));
 sg13g2_tiehi _15392__358 (.L_HI(net358));
 sg13g2_tiehi _16665__359 (.L_HI(net359));
 sg13g2_tiehi _15391__360 (.L_HI(net360));
 sg13g2_tiehi _15390__361 (.L_HI(net361));
 sg13g2_tiehi _15389__362 (.L_HI(net362));
 sg13g2_tiehi _15388__363 (.L_HI(net363));
 sg13g2_tiehi _15387__364 (.L_HI(net364));
 sg13g2_tiehi _15386__365 (.L_HI(net365));
 sg13g2_tiehi _15385__366 (.L_HI(net366));
 sg13g2_tiehi _15384__367 (.L_HI(net367));
 sg13g2_tiehi _15383__368 (.L_HI(net368));
 sg13g2_tiehi _15382__369 (.L_HI(net369));
 sg13g2_tiehi _15381__370 (.L_HI(net370));
 sg13g2_tiehi _15380__371 (.L_HI(net371));
 sg13g2_tiehi _15379__372 (.L_HI(net372));
 sg13g2_tiehi _15378__373 (.L_HI(net373));
 sg13g2_tiehi _15377__374 (.L_HI(net374));
 sg13g2_tiehi _15376__375 (.L_HI(net375));
 sg13g2_tiehi _15375__376 (.L_HI(net376));
 sg13g2_tiehi _15374__377 (.L_HI(net377));
 sg13g2_tiehi _15373__378 (.L_HI(net378));
 sg13g2_tiehi _15372__379 (.L_HI(net379));
 sg13g2_tiehi _15371__380 (.L_HI(net380));
 sg13g2_tiehi _15370__381 (.L_HI(net381));
 sg13g2_tiehi _15369__382 (.L_HI(net382));
 sg13g2_tiehi _15368__383 (.L_HI(net383));
 sg13g2_tiehi _15367__384 (.L_HI(net384));
 sg13g2_tiehi _15366__385 (.L_HI(net385));
 sg13g2_tiehi _15365__386 (.L_HI(net386));
 sg13g2_tiehi _15364__387 (.L_HI(net387));
 sg13g2_tiehi _15363__388 (.L_HI(net388));
 sg13g2_tiehi _15362__389 (.L_HI(net389));
 sg13g2_tiehi _15361__390 (.L_HI(net390));
 sg13g2_tiehi _15360__391 (.L_HI(net391));
 sg13g2_tiehi _15359__392 (.L_HI(net392));
 sg13g2_tiehi _15358__393 (.L_HI(net393));
 sg13g2_tiehi _15357__394 (.L_HI(net394));
 sg13g2_tiehi _15356__395 (.L_HI(net395));
 sg13g2_tiehi _15355__396 (.L_HI(net396));
 sg13g2_tiehi _15354__397 (.L_HI(net397));
 sg13g2_tiehi _15353__398 (.L_HI(net398));
 sg13g2_tiehi _15352__399 (.L_HI(net399));
 sg13g2_tiehi _15351__400 (.L_HI(net400));
 sg13g2_tiehi _15350__401 (.L_HI(net401));
 sg13g2_tiehi _15349__402 (.L_HI(net402));
 sg13g2_tiehi _15348__403 (.L_HI(net403));
 sg13g2_tiehi _15347__404 (.L_HI(net404));
 sg13g2_tiehi _15346__405 (.L_HI(net405));
 sg13g2_tiehi _15345__406 (.L_HI(net406));
 sg13g2_tiehi _15344__407 (.L_HI(net407));
 sg13g2_tiehi _15343__408 (.L_HI(net408));
 sg13g2_tiehi _15342__409 (.L_HI(net409));
 sg13g2_tiehi _15341__410 (.L_HI(net410));
 sg13g2_tiehi _15340__411 (.L_HI(net411));
 sg13g2_tiehi _15339__412 (.L_HI(net412));
 sg13g2_tiehi _15338__413 (.L_HI(net413));
 sg13g2_tiehi _15337__414 (.L_HI(net414));
 sg13g2_tiehi _15336__415 (.L_HI(net415));
 sg13g2_tiehi _15335__416 (.L_HI(net416));
 sg13g2_tiehi _15334__417 (.L_HI(net417));
 sg13g2_tiehi _15333__418 (.L_HI(net418));
 sg13g2_tiehi _15332__419 (.L_HI(net419));
 sg13g2_tiehi _15331__420 (.L_HI(net420));
 sg13g2_tiehi _15330__421 (.L_HI(net421));
 sg13g2_tiehi _15329__422 (.L_HI(net422));
 sg13g2_tiehi _15328__423 (.L_HI(net423));
 sg13g2_tiehi _15327__424 (.L_HI(net424));
 sg13g2_tiehi _15326__425 (.L_HI(net425));
 sg13g2_tiehi _15325__426 (.L_HI(net426));
 sg13g2_tiehi _15324__427 (.L_HI(net427));
 sg13g2_tiehi _15323__428 (.L_HI(net428));
 sg13g2_tiehi _15322__429 (.L_HI(net429));
 sg13g2_tiehi _15321__430 (.L_HI(net430));
 sg13g2_tiehi _15320__431 (.L_HI(net431));
 sg13g2_tiehi _15319__432 (.L_HI(net432));
 sg13g2_tiehi _15318__433 (.L_HI(net433));
 sg13g2_tiehi _15317__434 (.L_HI(net434));
 sg13g2_tiehi _15316__435 (.L_HI(net435));
 sg13g2_tiehi _15315__436 (.L_HI(net436));
 sg13g2_tiehi _15314__437 (.L_HI(net437));
 sg13g2_tiehi _15313__438 (.L_HI(net438));
 sg13g2_tiehi _15312__439 (.L_HI(net439));
 sg13g2_tiehi _15311__440 (.L_HI(net440));
 sg13g2_tiehi _15310__441 (.L_HI(net441));
 sg13g2_tiehi _15309__442 (.L_HI(net442));
 sg13g2_tiehi _15308__443 (.L_HI(net443));
 sg13g2_tiehi _15307__444 (.L_HI(net444));
 sg13g2_tiehi _15306__445 (.L_HI(net445));
 sg13g2_tiehi _15305__446 (.L_HI(net446));
 sg13g2_tiehi _15304__447 (.L_HI(net447));
 sg13g2_tiehi _15303__448 (.L_HI(net448));
 sg13g2_tiehi _15302__449 (.L_HI(net449));
 sg13g2_tiehi _15301__450 (.L_HI(net450));
 sg13g2_tiehi _15300__451 (.L_HI(net451));
 sg13g2_tiehi _15299__452 (.L_HI(net452));
 sg13g2_tiehi _15298__453 (.L_HI(net453));
 sg13g2_tiehi _15297__454 (.L_HI(net454));
 sg13g2_tiehi _15296__455 (.L_HI(net455));
 sg13g2_tiehi _15295__456 (.L_HI(net456));
 sg13g2_tiehi _15294__457 (.L_HI(net457));
 sg13g2_tiehi _15293__458 (.L_HI(net458));
 sg13g2_tiehi _15292__459 (.L_HI(net459));
 sg13g2_tiehi _15291__460 (.L_HI(net460));
 sg13g2_tiehi _15290__461 (.L_HI(net461));
 sg13g2_tiehi _15289__462 (.L_HI(net462));
 sg13g2_tiehi _15288__463 (.L_HI(net463));
 sg13g2_tiehi _15287__464 (.L_HI(net464));
 sg13g2_tiehi _15286__465 (.L_HI(net465));
 sg13g2_tiehi _15285__466 (.L_HI(net466));
 sg13g2_tiehi _15284__467 (.L_HI(net467));
 sg13g2_tiehi _15283__468 (.L_HI(net468));
 sg13g2_tiehi _15282__469 (.L_HI(net469));
 sg13g2_tiehi _15281__470 (.L_HI(net470));
 sg13g2_tiehi _15280__471 (.L_HI(net471));
 sg13g2_tiehi _15279__472 (.L_HI(net472));
 sg13g2_tiehi _15278__473 (.L_HI(net473));
 sg13g2_tiehi _15277__474 (.L_HI(net474));
 sg13g2_tiehi _15276__475 (.L_HI(net475));
 sg13g2_tiehi _15275__476 (.L_HI(net476));
 sg13g2_tiehi _15274__477 (.L_HI(net477));
 sg13g2_tiehi _15273__478 (.L_HI(net478));
 sg13g2_tiehi _15272__479 (.L_HI(net479));
 sg13g2_tiehi _15271__480 (.L_HI(net480));
 sg13g2_tiehi _15270__481 (.L_HI(net481));
 sg13g2_tiehi _15269__482 (.L_HI(net482));
 sg13g2_tiehi _15268__483 (.L_HI(net483));
 sg13g2_tiehi _15267__484 (.L_HI(net484));
 sg13g2_tiehi _15266__485 (.L_HI(net485));
 sg13g2_tiehi _15265__486 (.L_HI(net486));
 sg13g2_tiehi _15264__487 (.L_HI(net487));
 sg13g2_tiehi _15263__488 (.L_HI(net488));
 sg13g2_tiehi _15262__489 (.L_HI(net489));
 sg13g2_tiehi _15261__490 (.L_HI(net490));
 sg13g2_tiehi _15260__491 (.L_HI(net491));
 sg13g2_tiehi _15259__492 (.L_HI(net492));
 sg13g2_tiehi _15258__493 (.L_HI(net493));
 sg13g2_tiehi _15257__494 (.L_HI(net494));
 sg13g2_tiehi _15256__495 (.L_HI(net495));
 sg13g2_tiehi _15255__496 (.L_HI(net496));
 sg13g2_tiehi _15254__497 (.L_HI(net497));
 sg13g2_tiehi _15253__498 (.L_HI(net498));
 sg13g2_tiehi _15252__499 (.L_HI(net499));
 sg13g2_tiehi _15251__500 (.L_HI(net500));
 sg13g2_tiehi _15250__501 (.L_HI(net501));
 sg13g2_tiehi _15249__502 (.L_HI(net502));
 sg13g2_tiehi _15248__503 (.L_HI(net503));
 sg13g2_tiehi _15247__504 (.L_HI(net504));
 sg13g2_tiehi _15246__505 (.L_HI(net505));
 sg13g2_tiehi _15245__506 (.L_HI(net506));
 sg13g2_tiehi _15244__507 (.L_HI(net507));
 sg13g2_tiehi _15243__508 (.L_HI(net508));
 sg13g2_tiehi _15242__509 (.L_HI(net509));
 sg13g2_tiehi _15241__510 (.L_HI(net510));
 sg13g2_tiehi _15240__511 (.L_HI(net511));
 sg13g2_tiehi _15239__512 (.L_HI(net512));
 sg13g2_tiehi _15238__513 (.L_HI(net513));
 sg13g2_tiehi _15237__514 (.L_HI(net514));
 sg13g2_tiehi _15236__515 (.L_HI(net515));
 sg13g2_tiehi _15235__516 (.L_HI(net516));
 sg13g2_tiehi _15234__517 (.L_HI(net517));
 sg13g2_tiehi _15233__518 (.L_HI(net518));
 sg13g2_tiehi _15232__519 (.L_HI(net519));
 sg13g2_tiehi _15231__520 (.L_HI(net520));
 sg13g2_tiehi _15230__521 (.L_HI(net521));
 sg13g2_tiehi _15229__522 (.L_HI(net522));
 sg13g2_tiehi _15228__523 (.L_HI(net523));
 sg13g2_tiehi _15227__524 (.L_HI(net524));
 sg13g2_tiehi _15226__525 (.L_HI(net525));
 sg13g2_tiehi _15225__526 (.L_HI(net526));
 sg13g2_tiehi _15224__527 (.L_HI(net527));
 sg13g2_tiehi _15223__528 (.L_HI(net528));
 sg13g2_tiehi _15222__529 (.L_HI(net529));
 sg13g2_tiehi _15221__530 (.L_HI(net530));
 sg13g2_tiehi _15220__531 (.L_HI(net531));
 sg13g2_tiehi _15219__532 (.L_HI(net532));
 sg13g2_tiehi _15218__533 (.L_HI(net533));
 sg13g2_tiehi _15217__534 (.L_HI(net534));
 sg13g2_tiehi _15216__535 (.L_HI(net535));
 sg13g2_tiehi _15215__536 (.L_HI(net536));
 sg13g2_tiehi _15214__537 (.L_HI(net537));
 sg13g2_tiehi _15213__538 (.L_HI(net538));
 sg13g2_tiehi _15212__539 (.L_HI(net539));
 sg13g2_tiehi _15211__540 (.L_HI(net540));
 sg13g2_tiehi _15210__541 (.L_HI(net541));
 sg13g2_tiehi _15209__542 (.L_HI(net542));
 sg13g2_tiehi _15208__543 (.L_HI(net543));
 sg13g2_tiehi _15207__544 (.L_HI(net544));
 sg13g2_tiehi _16664__545 (.L_HI(net545));
 sg13g2_tiehi _15206__546 (.L_HI(net546));
 sg13g2_tiehi _16663__547 (.L_HI(net547));
 sg13g2_tiehi _15205__548 (.L_HI(net548));
 sg13g2_tiehi _16662__549 (.L_HI(net549));
 sg13g2_tiehi _15204__550 (.L_HI(net550));
 sg13g2_tiehi _16661__551 (.L_HI(net551));
 sg13g2_tiehi _15203__552 (.L_HI(net552));
 sg13g2_tiehi _16660__553 (.L_HI(net553));
 sg13g2_tiehi _15202__554 (.L_HI(net554));
 sg13g2_tiehi _16659__555 (.L_HI(net555));
 sg13g2_tiehi _15201__556 (.L_HI(net556));
 sg13g2_tiehi _16658__557 (.L_HI(net557));
 sg13g2_tiehi _15200__558 (.L_HI(net558));
 sg13g2_tiehi _16657__559 (.L_HI(net559));
 sg13g2_tiehi _15199__560 (.L_HI(net560));
 sg13g2_tiehi _16656__561 (.L_HI(net561));
 sg13g2_tiehi _15198__562 (.L_HI(net562));
 sg13g2_tiehi _16655__563 (.L_HI(net563));
 sg13g2_tiehi _15197__564 (.L_HI(net564));
 sg13g2_tiehi _16654__565 (.L_HI(net565));
 sg13g2_tiehi _15196__566 (.L_HI(net566));
 sg13g2_tiehi _16653__567 (.L_HI(net567));
 sg13g2_tiehi _15195__568 (.L_HI(net568));
 sg13g2_tiehi _16652__569 (.L_HI(net569));
 sg13g2_tiehi _15194__570 (.L_HI(net570));
 sg13g2_tiehi _16651__571 (.L_HI(net571));
 sg13g2_tiehi _15193__572 (.L_HI(net572));
 sg13g2_tiehi _16650__573 (.L_HI(net573));
 sg13g2_tiehi _15192__574 (.L_HI(net574));
 sg13g2_tiehi _16649__575 (.L_HI(net575));
 sg13g2_tiehi _15191__576 (.L_HI(net576));
 sg13g2_tiehi _16648__577 (.L_HI(net577));
 sg13g2_tiehi _15190__578 (.L_HI(net578));
 sg13g2_tiehi _16647__579 (.L_HI(net579));
 sg13g2_tiehi _15189__580 (.L_HI(net580));
 sg13g2_tiehi _16646__581 (.L_HI(net581));
 sg13g2_tiehi _15188__582 (.L_HI(net582));
 sg13g2_tiehi _16645__583 (.L_HI(net583));
 sg13g2_tiehi _15187__584 (.L_HI(net584));
 sg13g2_tiehi _16644__585 (.L_HI(net585));
 sg13g2_tiehi _15186__586 (.L_HI(net586));
 sg13g2_tiehi _16643__587 (.L_HI(net587));
 sg13g2_tiehi _15185__588 (.L_HI(net588));
 sg13g2_tiehi _16642__589 (.L_HI(net589));
 sg13g2_tiehi _15184__590 (.L_HI(net590));
 sg13g2_tiehi _16641__591 (.L_HI(net591));
 sg13g2_tiehi _15183__592 (.L_HI(net592));
 sg13g2_tiehi _16640__593 (.L_HI(net593));
 sg13g2_tiehi _15182__594 (.L_HI(net594));
 sg13g2_tiehi _16639__595 (.L_HI(net595));
 sg13g2_tiehi _15181__596 (.L_HI(net596));
 sg13g2_tiehi _16638__597 (.L_HI(net597));
 sg13g2_tiehi _15180__598 (.L_HI(net598));
 sg13g2_tiehi _16637__599 (.L_HI(net599));
 sg13g2_tiehi _15179__600 (.L_HI(net600));
 sg13g2_tiehi _16636__601 (.L_HI(net601));
 sg13g2_tiehi _15178__602 (.L_HI(net602));
 sg13g2_tiehi _16635__603 (.L_HI(net603));
 sg13g2_tiehi _15177__604 (.L_HI(net604));
 sg13g2_tiehi _16634__605 (.L_HI(net605));
 sg13g2_tiehi _15176__606 (.L_HI(net606));
 sg13g2_tiehi _16633__607 (.L_HI(net607));
 sg13g2_tiehi _15175__608 (.L_HI(net608));
 sg13g2_tiehi _16632__609 (.L_HI(net609));
 sg13g2_tiehi _15174__610 (.L_HI(net610));
 sg13g2_tiehi _16631__611 (.L_HI(net611));
 sg13g2_tiehi _15173__612 (.L_HI(net612));
 sg13g2_tiehi _16630__613 (.L_HI(net613));
 sg13g2_tiehi _15172__614 (.L_HI(net614));
 sg13g2_tiehi _16629__615 (.L_HI(net615));
 sg13g2_tiehi _15171__616 (.L_HI(net616));
 sg13g2_tiehi _16628__617 (.L_HI(net617));
 sg13g2_tiehi _15170__618 (.L_HI(net618));
 sg13g2_tiehi _16627__619 (.L_HI(net619));
 sg13g2_tiehi _15169__620 (.L_HI(net620));
 sg13g2_tiehi _16626__621 (.L_HI(net621));
 sg13g2_tiehi _15168__622 (.L_HI(net622));
 sg13g2_tiehi _16625__623 (.L_HI(net623));
 sg13g2_tiehi _15167__624 (.L_HI(net624));
 sg13g2_tiehi _16624__625 (.L_HI(net625));
 sg13g2_tiehi _15166__626 (.L_HI(net626));
 sg13g2_tiehi _16623__627 (.L_HI(net627));
 sg13g2_tiehi _15165__628 (.L_HI(net628));
 sg13g2_tiehi _16622__629 (.L_HI(net629));
 sg13g2_tiehi _15164__630 (.L_HI(net630));
 sg13g2_tiehi _16621__631 (.L_HI(net631));
 sg13g2_tiehi _15163__632 (.L_HI(net632));
 sg13g2_tiehi _16620__633 (.L_HI(net633));
 sg13g2_tiehi _15162__634 (.L_HI(net634));
 sg13g2_tiehi _16619__635 (.L_HI(net635));
 sg13g2_tiehi _15161__636 (.L_HI(net636));
 sg13g2_tiehi _16618__637 (.L_HI(net637));
 sg13g2_tiehi _15160__638 (.L_HI(net638));
 sg13g2_tiehi _16617__639 (.L_HI(net639));
 sg13g2_tiehi _15159__640 (.L_HI(net640));
 sg13g2_tiehi _16616__641 (.L_HI(net641));
 sg13g2_tiehi _15158__642 (.L_HI(net642));
 sg13g2_tiehi _16615__643 (.L_HI(net643));
 sg13g2_tiehi _15157__644 (.L_HI(net644));
 sg13g2_tiehi _16614__645 (.L_HI(net645));
 sg13g2_tiehi _15156__646 (.L_HI(net646));
 sg13g2_tiehi _16613__647 (.L_HI(net647));
 sg13g2_tiehi _15155__648 (.L_HI(net648));
 sg13g2_tiehi _16612__649 (.L_HI(net649));
 sg13g2_tiehi _15154__650 (.L_HI(net650));
 sg13g2_tiehi _16611__651 (.L_HI(net651));
 sg13g2_tiehi _15153__652 (.L_HI(net652));
 sg13g2_tiehi _16610__653 (.L_HI(net653));
 sg13g2_tiehi _15152__654 (.L_HI(net654));
 sg13g2_tiehi _16609__655 (.L_HI(net655));
 sg13g2_tiehi _15151__656 (.L_HI(net656));
 sg13g2_tiehi _16608__657 (.L_HI(net657));
 sg13g2_tiehi _15150__658 (.L_HI(net658));
 sg13g2_tiehi _16607__659 (.L_HI(net659));
 sg13g2_tiehi _15149__660 (.L_HI(net660));
 sg13g2_tiehi _16606__661 (.L_HI(net661));
 sg13g2_tiehi _15148__662 (.L_HI(net662));
 sg13g2_tiehi _15147__663 (.L_HI(net663));
 sg13g2_tiehi _15146__664 (.L_HI(net664));
 sg13g2_tiehi _15145__665 (.L_HI(net665));
 sg13g2_tiehi _15144__666 (.L_HI(net666));
 sg13g2_tiehi _15143__667 (.L_HI(net667));
 sg13g2_tiehi _15142__668 (.L_HI(net668));
 sg13g2_tiehi _15141__669 (.L_HI(net669));
 sg13g2_tiehi _15140__670 (.L_HI(net670));
 sg13g2_tiehi _15139__671 (.L_HI(net671));
 sg13g2_tiehi _15138__672 (.L_HI(net672));
 sg13g2_tiehi _15137__673 (.L_HI(net673));
 sg13g2_tiehi _15136__674 (.L_HI(net674));
 sg13g2_tiehi _15135__675 (.L_HI(net675));
 sg13g2_tiehi _15134__676 (.L_HI(net676));
 sg13g2_tiehi _15133__677 (.L_HI(net677));
 sg13g2_tiehi _15132__678 (.L_HI(net678));
 sg13g2_tiehi _15131__679 (.L_HI(net679));
 sg13g2_tiehi _15130__680 (.L_HI(net680));
 sg13g2_tiehi _15129__681 (.L_HI(net681));
 sg13g2_tiehi _15128__682 (.L_HI(net682));
 sg13g2_tiehi _15127__683 (.L_HI(net683));
 sg13g2_tiehi _15126__684 (.L_HI(net684));
 sg13g2_tiehi _15125__685 (.L_HI(net685));
 sg13g2_tiehi _15124__686 (.L_HI(net686));
 sg13g2_tiehi _15123__687 (.L_HI(net687));
 sg13g2_tiehi _15122__688 (.L_HI(net688));
 sg13g2_tiehi _15121__689 (.L_HI(net689));
 sg13g2_tiehi _15120__690 (.L_HI(net690));
 sg13g2_tiehi _15119__691 (.L_HI(net691));
 sg13g2_tiehi _15118__692 (.L_HI(net692));
 sg13g2_tiehi _15117__693 (.L_HI(net693));
 sg13g2_tiehi _15116__694 (.L_HI(net694));
 sg13g2_tiehi _15115__695 (.L_HI(net695));
 sg13g2_tiehi _15114__696 (.L_HI(net696));
 sg13g2_tiehi _15113__697 (.L_HI(net697));
 sg13g2_tiehi _15112__698 (.L_HI(net698));
 sg13g2_tiehi _15111__699 (.L_HI(net699));
 sg13g2_tiehi _15110__700 (.L_HI(net700));
 sg13g2_tiehi _15109__701 (.L_HI(net701));
 sg13g2_tiehi _15108__702 (.L_HI(net702));
 sg13g2_tiehi _15107__703 (.L_HI(net703));
 sg13g2_tiehi _15106__704 (.L_HI(net704));
 sg13g2_tiehi _15105__705 (.L_HI(net705));
 sg13g2_tiehi _15104__706 (.L_HI(net706));
 sg13g2_tiehi _15103__707 (.L_HI(net707));
 sg13g2_tiehi _15102__708 (.L_HI(net708));
 sg13g2_tiehi _15101__709 (.L_HI(net709));
 sg13g2_tiehi _15100__710 (.L_HI(net710));
 sg13g2_tiehi _15099__711 (.L_HI(net711));
 sg13g2_tiehi _15098__712 (.L_HI(net712));
 sg13g2_tiehi _15097__713 (.L_HI(net713));
 sg13g2_tiehi _15096__714 (.L_HI(net714));
 sg13g2_tiehi _15095__715 (.L_HI(net715));
 sg13g2_tiehi _15094__716 (.L_HI(net716));
 sg13g2_tiehi _15093__717 (.L_HI(net717));
 sg13g2_tiehi _15092__718 (.L_HI(net718));
 sg13g2_tiehi _15091__719 (.L_HI(net719));
 sg13g2_tiehi _15090__720 (.L_HI(net720));
 sg13g2_tiehi _15089__721 (.L_HI(net721));
 sg13g2_tiehi _15088__722 (.L_HI(net722));
 sg13g2_tiehi _15087__723 (.L_HI(net723));
 sg13g2_tiehi _15086__724 (.L_HI(net724));
 sg13g2_tiehi _15085__725 (.L_HI(net725));
 sg13g2_tiehi _15084__726 (.L_HI(net726));
 sg13g2_tiehi _15083__727 (.L_HI(net727));
 sg13g2_tiehi _15082__728 (.L_HI(net728));
 sg13g2_tiehi _15081__729 (.L_HI(net729));
 sg13g2_tiehi _15080__730 (.L_HI(net730));
 sg13g2_tiehi _15079__731 (.L_HI(net731));
 sg13g2_tiehi _15078__732 (.L_HI(net732));
 sg13g2_tiehi _15077__733 (.L_HI(net733));
 sg13g2_tiehi _15076__734 (.L_HI(net734));
 sg13g2_tiehi _15075__735 (.L_HI(net735));
 sg13g2_tiehi _15074__736 (.L_HI(net736));
 sg13g2_tiehi _15073__737 (.L_HI(net737));
 sg13g2_tiehi _15072__738 (.L_HI(net738));
 sg13g2_tiehi _15071__739 (.L_HI(net739));
 sg13g2_tiehi _15070__740 (.L_HI(net740));
 sg13g2_tiehi _15069__741 (.L_HI(net741));
 sg13g2_tiehi _15068__742 (.L_HI(net742));
 sg13g2_tiehi _15067__743 (.L_HI(net743));
 sg13g2_tiehi _15066__744 (.L_HI(net744));
 sg13g2_tiehi _15065__745 (.L_HI(net745));
 sg13g2_tiehi _15064__746 (.L_HI(net746));
 sg13g2_tiehi _15063__747 (.L_HI(net747));
 sg13g2_tiehi _15062__748 (.L_HI(net748));
 sg13g2_tiehi _15061__749 (.L_HI(net749));
 sg13g2_tiehi _15060__750 (.L_HI(net750));
 sg13g2_tiehi _15059__751 (.L_HI(net751));
 sg13g2_tiehi _15058__752 (.L_HI(net752));
 sg13g2_tiehi _15057__753 (.L_HI(net753));
 sg13g2_tiehi _15056__754 (.L_HI(net754));
 sg13g2_tiehi _15055__755 (.L_HI(net755));
 sg13g2_tiehi _15054__756 (.L_HI(net756));
 sg13g2_tiehi _15053__757 (.L_HI(net757));
 sg13g2_tiehi _15052__758 (.L_HI(net758));
 sg13g2_tiehi _15051__759 (.L_HI(net759));
 sg13g2_tiehi _15050__760 (.L_HI(net760));
 sg13g2_tiehi _15049__761 (.L_HI(net761));
 sg13g2_tiehi _15048__762 (.L_HI(net762));
 sg13g2_tiehi _15047__763 (.L_HI(net763));
 sg13g2_tiehi _15046__764 (.L_HI(net764));
 sg13g2_tiehi _15045__765 (.L_HI(net765));
 sg13g2_tiehi _15044__766 (.L_HI(net766));
 sg13g2_tiehi _15043__767 (.L_HI(net767));
 sg13g2_tiehi _15042__768 (.L_HI(net768));
 sg13g2_tiehi _15041__769 (.L_HI(net769));
 sg13g2_tiehi _15040__770 (.L_HI(net770));
 sg13g2_tiehi _15039__771 (.L_HI(net771));
 sg13g2_tiehi _15038__772 (.L_HI(net772));
 sg13g2_tiehi _15037__773 (.L_HI(net773));
 sg13g2_tiehi _15036__774 (.L_HI(net774));
 sg13g2_tiehi _15035__775 (.L_HI(net775));
 sg13g2_tiehi _15034__776 (.L_HI(net776));
 sg13g2_tiehi _15033__777 (.L_HI(net777));
 sg13g2_tiehi _15032__778 (.L_HI(net778));
 sg13g2_tiehi _15031__779 (.L_HI(net779));
 sg13g2_tiehi _15030__780 (.L_HI(net780));
 sg13g2_tiehi _15029__781 (.L_HI(net781));
 sg13g2_tiehi _15028__782 (.L_HI(net782));
 sg13g2_tiehi _15027__783 (.L_HI(net783));
 sg13g2_tiehi _15026__784 (.L_HI(net784));
 sg13g2_tiehi _15025__785 (.L_HI(net785));
 sg13g2_tiehi _15024__786 (.L_HI(net786));
 sg13g2_tiehi _15023__787 (.L_HI(net787));
 sg13g2_tiehi _15022__788 (.L_HI(net788));
 sg13g2_tiehi _15021__789 (.L_HI(net789));
 sg13g2_tiehi _15020__790 (.L_HI(net790));
 sg13g2_tiehi _15019__791 (.L_HI(net791));
 sg13g2_tiehi _15018__792 (.L_HI(net792));
 sg13g2_tiehi _15017__793 (.L_HI(net793));
 sg13g2_tiehi _15016__794 (.L_HI(net794));
 sg13g2_tiehi _15015__795 (.L_HI(net795));
 sg13g2_tiehi _15014__796 (.L_HI(net796));
 sg13g2_tiehi _15013__797 (.L_HI(net797));
 sg13g2_tiehi _15012__798 (.L_HI(net798));
 sg13g2_tiehi _15011__799 (.L_HI(net799));
 sg13g2_tiehi _15010__800 (.L_HI(net800));
 sg13g2_tiehi _15009__801 (.L_HI(net801));
 sg13g2_tiehi _15008__802 (.L_HI(net802));
 sg13g2_tiehi _15007__803 (.L_HI(net803));
 sg13g2_tiehi _15006__804 (.L_HI(net804));
 sg13g2_tiehi _15005__805 (.L_HI(net805));
 sg13g2_tiehi _15004__806 (.L_HI(net806));
 sg13g2_tiehi _15003__807 (.L_HI(net807));
 sg13g2_tiehi _15002__808 (.L_HI(net808));
 sg13g2_tiehi _15001__809 (.L_HI(net809));
 sg13g2_tiehi _15000__810 (.L_HI(net810));
 sg13g2_tiehi _14999__811 (.L_HI(net811));
 sg13g2_tiehi _14998__812 (.L_HI(net812));
 sg13g2_tiehi _14997__813 (.L_HI(net813));
 sg13g2_tiehi _14996__814 (.L_HI(net814));
 sg13g2_tiehi _14995__815 (.L_HI(net815));
 sg13g2_tiehi _14994__816 (.L_HI(net816));
 sg13g2_tiehi _14993__817 (.L_HI(net817));
 sg13g2_tiehi _14992__818 (.L_HI(net818));
 sg13g2_tiehi _14991__819 (.L_HI(net819));
 sg13g2_tiehi _14990__820 (.L_HI(net820));
 sg13g2_tiehi _14989__821 (.L_HI(net821));
 sg13g2_tiehi _14988__822 (.L_HI(net822));
 sg13g2_tiehi _14987__823 (.L_HI(net823));
 sg13g2_tiehi _14986__824 (.L_HI(net824));
 sg13g2_tiehi _14985__825 (.L_HI(net825));
 sg13g2_tiehi _14984__826 (.L_HI(net826));
 sg13g2_tiehi _14983__827 (.L_HI(net827));
 sg13g2_tiehi _14982__828 (.L_HI(net828));
 sg13g2_tiehi _14981__829 (.L_HI(net829));
 sg13g2_tiehi _14980__830 (.L_HI(net830));
 sg13g2_tiehi _14979__831 (.L_HI(net831));
 sg13g2_tiehi _14978__832 (.L_HI(net832));
 sg13g2_tiehi _14977__833 (.L_HI(net833));
 sg13g2_tiehi _14976__834 (.L_HI(net834));
 sg13g2_tiehi _14975__835 (.L_HI(net835));
 sg13g2_tiehi _14974__836 (.L_HI(net836));
 sg13g2_tiehi _14973__837 (.L_HI(net837));
 sg13g2_tiehi _14972__838 (.L_HI(net838));
 sg13g2_tiehi _14971__839 (.L_HI(net839));
 sg13g2_tiehi _14970__840 (.L_HI(net840));
 sg13g2_tiehi _14969__841 (.L_HI(net841));
 sg13g2_tiehi _14968__842 (.L_HI(net842));
 sg13g2_tiehi _14967__843 (.L_HI(net843));
 sg13g2_tiehi _14966__844 (.L_HI(net844));
 sg13g2_tiehi _14965__845 (.L_HI(net845));
 sg13g2_tiehi _14964__846 (.L_HI(net846));
 sg13g2_tiehi _14963__847 (.L_HI(net847));
 sg13g2_tiehi _14962__848 (.L_HI(net848));
 sg13g2_tiehi _14961__849 (.L_HI(net849));
 sg13g2_tiehi _14960__850 (.L_HI(net850));
 sg13g2_tiehi _14959__851 (.L_HI(net851));
 sg13g2_tiehi _14958__852 (.L_HI(net852));
 sg13g2_tiehi _14957__853 (.L_HI(net853));
 sg13g2_tiehi _14956__854 (.L_HI(net854));
 sg13g2_tiehi _14955__855 (.L_HI(net855));
 sg13g2_tiehi _14954__856 (.L_HI(net856));
 sg13g2_tiehi _14953__857 (.L_HI(net857));
 sg13g2_tiehi _14952__858 (.L_HI(net858));
 sg13g2_tiehi _14951__859 (.L_HI(net859));
 sg13g2_tiehi _14950__860 (.L_HI(net860));
 sg13g2_tiehi _14949__861 (.L_HI(net861));
 sg13g2_tiehi _14948__862 (.L_HI(net862));
 sg13g2_tiehi _14947__863 (.L_HI(net863));
 sg13g2_tiehi _14946__864 (.L_HI(net864));
 sg13g2_tiehi _14945__865 (.L_HI(net865));
 sg13g2_tiehi _14944__866 (.L_HI(net866));
 sg13g2_tiehi _14943__867 (.L_HI(net867));
 sg13g2_tiehi _14942__868 (.L_HI(net868));
 sg13g2_tiehi _14941__869 (.L_HI(net869));
 sg13g2_tiehi _14940__870 (.L_HI(net870));
 sg13g2_tiehi _14939__871 (.L_HI(net871));
 sg13g2_tiehi _14938__872 (.L_HI(net872));
 sg13g2_tiehi _14937__873 (.L_HI(net873));
 sg13g2_tiehi _14936__874 (.L_HI(net874));
 sg13g2_tiehi _14935__875 (.L_HI(net875));
 sg13g2_tiehi _14934__876 (.L_HI(net876));
 sg13g2_tiehi _14933__877 (.L_HI(net877));
 sg13g2_tiehi _14932__878 (.L_HI(net878));
 sg13g2_tiehi _14931__879 (.L_HI(net879));
 sg13g2_tiehi _14930__880 (.L_HI(net880));
 sg13g2_tiehi _14929__881 (.L_HI(net881));
 sg13g2_tiehi _14928__882 (.L_HI(net882));
 sg13g2_tiehi _14927__883 (.L_HI(net883));
 sg13g2_tiehi _14926__884 (.L_HI(net884));
 sg13g2_tiehi _14925__885 (.L_HI(net885));
 sg13g2_tiehi _14924__886 (.L_HI(net886));
 sg13g2_tiehi _14923__887 (.L_HI(net887));
 sg13g2_tiehi _14922__888 (.L_HI(net888));
 sg13g2_tiehi _14921__889 (.L_HI(net889));
 sg13g2_tiehi _14920__890 (.L_HI(net890));
 sg13g2_tiehi _14919__891 (.L_HI(net891));
 sg13g2_tiehi _14918__892 (.L_HI(net892));
 sg13g2_tiehi _14917__893 (.L_HI(net893));
 sg13g2_tiehi _14916__894 (.L_HI(net894));
 sg13g2_tiehi _14915__895 (.L_HI(net895));
 sg13g2_tiehi _14914__896 (.L_HI(net896));
 sg13g2_tiehi _14913__897 (.L_HI(net897));
 sg13g2_tiehi _14912__898 (.L_HI(net898));
 sg13g2_tiehi _14911__899 (.L_HI(net899));
 sg13g2_tiehi _14910__900 (.L_HI(net900));
 sg13g2_tiehi _14909__901 (.L_HI(net901));
 sg13g2_tiehi _14908__902 (.L_HI(net902));
 sg13g2_tiehi _14907__903 (.L_HI(net903));
 sg13g2_tiehi _14906__904 (.L_HI(net904));
 sg13g2_tiehi _14905__905 (.L_HI(net905));
 sg13g2_tiehi _14904__906 (.L_HI(net906));
 sg13g2_tiehi _14903__907 (.L_HI(net907));
 sg13g2_tiehi _14902__908 (.L_HI(net908));
 sg13g2_tiehi _14901__909 (.L_HI(net909));
 sg13g2_tiehi _14900__910 (.L_HI(net910));
 sg13g2_tiehi _14899__911 (.L_HI(net911));
 sg13g2_tiehi _14898__912 (.L_HI(net912));
 sg13g2_tiehi _14897__913 (.L_HI(net913));
 sg13g2_tiehi _14896__914 (.L_HI(net914));
 sg13g2_tiehi _14895__915 (.L_HI(net915));
 sg13g2_tiehi _14894__916 (.L_HI(net916));
 sg13g2_tiehi _14893__917 (.L_HI(net917));
 sg13g2_tiehi _14892__918 (.L_HI(net918));
 sg13g2_tiehi _14891__919 (.L_HI(net919));
 sg13g2_tiehi _14890__920 (.L_HI(net920));
 sg13g2_tiehi _14889__921 (.L_HI(net921));
 sg13g2_tiehi _14888__922 (.L_HI(net922));
 sg13g2_tiehi _14887__923 (.L_HI(net923));
 sg13g2_tiehi _14886__924 (.L_HI(net924));
 sg13g2_tiehi _14885__925 (.L_HI(net925));
 sg13g2_tiehi _14884__926 (.L_HI(net926));
 sg13g2_tiehi _14883__927 (.L_HI(net927));
 sg13g2_tiehi _14882__928 (.L_HI(net928));
 sg13g2_tiehi _14881__929 (.L_HI(net929));
 sg13g2_tiehi _14880__930 (.L_HI(net930));
 sg13g2_tiehi _14879__931 (.L_HI(net931));
 sg13g2_tiehi _14878__932 (.L_HI(net932));
 sg13g2_tiehi _14877__933 (.L_HI(net933));
 sg13g2_tiehi _14876__934 (.L_HI(net934));
 sg13g2_tiehi _14875__935 (.L_HI(net935));
 sg13g2_tiehi _14874__936 (.L_HI(net936));
 sg13g2_tiehi _14873__937 (.L_HI(net937));
 sg13g2_tiehi _14872__938 (.L_HI(net938));
 sg13g2_tiehi _14871__939 (.L_HI(net939));
 sg13g2_tiehi _14870__940 (.L_HI(net940));
 sg13g2_tiehi _14869__941 (.L_HI(net941));
 sg13g2_tiehi _14868__942 (.L_HI(net942));
 sg13g2_tiehi _14867__943 (.L_HI(net943));
 sg13g2_tiehi _14866__944 (.L_HI(net944));
 sg13g2_tiehi _14865__945 (.L_HI(net945));
 sg13g2_tiehi _14864__946 (.L_HI(net946));
 sg13g2_tiehi _14863__947 (.L_HI(net947));
 sg13g2_tiehi _14862__948 (.L_HI(net948));
 sg13g2_tiehi _14861__949 (.L_HI(net949));
 sg13g2_tiehi _14860__950 (.L_HI(net950));
 sg13g2_tiehi _14859__951 (.L_HI(net951));
 sg13g2_tiehi _14858__952 (.L_HI(net952));
 sg13g2_tiehi _14857__953 (.L_HI(net953));
 sg13g2_tiehi _14856__954 (.L_HI(net954));
 sg13g2_tiehi _14855__955 (.L_HI(net955));
 sg13g2_tiehi _14854__956 (.L_HI(net956));
 sg13g2_tiehi _14853__957 (.L_HI(net957));
 sg13g2_tiehi _14852__958 (.L_HI(net958));
 sg13g2_tiehi _14851__959 (.L_HI(net959));
 sg13g2_tiehi _14850__960 (.L_HI(net960));
 sg13g2_tiehi _14849__961 (.L_HI(net961));
 sg13g2_tiehi _14848__962 (.L_HI(net962));
 sg13g2_tiehi _14847__963 (.L_HI(net963));
 sg13g2_tiehi _14846__964 (.L_HI(net964));
 sg13g2_tiehi _14845__965 (.L_HI(net965));
 sg13g2_tiehi _14844__966 (.L_HI(net966));
 sg13g2_tiehi _14843__967 (.L_HI(net967));
 sg13g2_tiehi _14842__968 (.L_HI(net968));
 sg13g2_tiehi _14841__969 (.L_HI(net969));
 sg13g2_tiehi _14840__970 (.L_HI(net970));
 sg13g2_tiehi _14839__971 (.L_HI(net971));
 sg13g2_tiehi _14838__972 (.L_HI(net972));
 sg13g2_tiehi _14837__973 (.L_HI(net973));
 sg13g2_tiehi _14836__974 (.L_HI(net974));
 sg13g2_tiehi _14835__975 (.L_HI(net975));
 sg13g2_tiehi _14834__976 (.L_HI(net976));
 sg13g2_tiehi _14833__977 (.L_HI(net977));
 sg13g2_tiehi _14832__978 (.L_HI(net978));
 sg13g2_tiehi _14831__979 (.L_HI(net979));
 sg13g2_tiehi _14830__980 (.L_HI(net980));
 sg13g2_tiehi _14829__981 (.L_HI(net981));
 sg13g2_tiehi _14828__982 (.L_HI(net982));
 sg13g2_tiehi _14827__983 (.L_HI(net983));
 sg13g2_tiehi _14826__984 (.L_HI(net984));
 sg13g2_tiehi _14825__985 (.L_HI(net985));
 sg13g2_tiehi _14824__986 (.L_HI(net986));
 sg13g2_tiehi _14823__987 (.L_HI(net987));
 sg13g2_tiehi _14822__988 (.L_HI(net988));
 sg13g2_tiehi _14821__989 (.L_HI(net989));
 sg13g2_tiehi _14820__990 (.L_HI(net990));
 sg13g2_tiehi _14819__991 (.L_HI(net991));
 sg13g2_tiehi _14818__992 (.L_HI(net992));
 sg13g2_tiehi _14817__993 (.L_HI(net993));
 sg13g2_tiehi _14816__994 (.L_HI(net994));
 sg13g2_tiehi _14815__995 (.L_HI(net995));
 sg13g2_tiehi _14814__996 (.L_HI(net996));
 sg13g2_tiehi _14813__997 (.L_HI(net997));
 sg13g2_tiehi _14812__998 (.L_HI(net998));
 sg13g2_tiehi _14811__999 (.L_HI(net999));
 sg13g2_tiehi _14810__1000 (.L_HI(net1000));
 sg13g2_tiehi _14809__1001 (.L_HI(net1001));
 sg13g2_tiehi _14808__1002 (.L_HI(net1002));
 sg13g2_tiehi _14807__1003 (.L_HI(net1003));
 sg13g2_tiehi _14806__1004 (.L_HI(net1004));
 sg13g2_tiehi _14805__1005 (.L_HI(net1005));
 sg13g2_tiehi _14804__1006 (.L_HI(net1006));
 sg13g2_tiehi _14803__1007 (.L_HI(net1007));
 sg13g2_tiehi _14802__1008 (.L_HI(net1008));
 sg13g2_tiehi _14801__1009 (.L_HI(net1009));
 sg13g2_tiehi _14800__1010 (.L_HI(net1010));
 sg13g2_tiehi _14799__1011 (.L_HI(net1011));
 sg13g2_tiehi _14798__1012 (.L_HI(net1012));
 sg13g2_tiehi _14797__1013 (.L_HI(net1013));
 sg13g2_tiehi _14796__1014 (.L_HI(net1014));
 sg13g2_tiehi _14795__1015 (.L_HI(net1015));
 sg13g2_tiehi _14794__1016 (.L_HI(net1016));
 sg13g2_tiehi _14793__1017 (.L_HI(net1017));
 sg13g2_tiehi _14792__1018 (.L_HI(net1018));
 sg13g2_tiehi _14791__1019 (.L_HI(net1019));
 sg13g2_tiehi _14790__1020 (.L_HI(net1020));
 sg13g2_tiehi _14789__1021 (.L_HI(net1021));
 sg13g2_tiehi _14788__1022 (.L_HI(net1022));
 sg13g2_tiehi _14787__1023 (.L_HI(net1023));
 sg13g2_tiehi _14786__1024 (.L_HI(net1024));
 sg13g2_tiehi _14785__1025 (.L_HI(net1025));
 sg13g2_tiehi _14784__1026 (.L_HI(net1026));
 sg13g2_tiehi _14783__1027 (.L_HI(net1027));
 sg13g2_tiehi _14782__1028 (.L_HI(net1028));
 sg13g2_tiehi _14781__1029 (.L_HI(net1029));
 sg13g2_tiehi _14780__1030 (.L_HI(net1030));
 sg13g2_tiehi _14779__1031 (.L_HI(net1031));
 sg13g2_tiehi _14778__1032 (.L_HI(net1032));
 sg13g2_tiehi _14777__1033 (.L_HI(net1033));
 sg13g2_tiehi _14776__1034 (.L_HI(net1034));
 sg13g2_tiehi _14775__1035 (.L_HI(net1035));
 sg13g2_tiehi _14774__1036 (.L_HI(net1036));
 sg13g2_tiehi _14773__1037 (.L_HI(net1037));
 sg13g2_tiehi _14772__1038 (.L_HI(net1038));
 sg13g2_tiehi _14771__1039 (.L_HI(net1039));
 sg13g2_tiehi _14770__1040 (.L_HI(net1040));
 sg13g2_tiehi _14769__1041 (.L_HI(net1041));
 sg13g2_tiehi _14768__1042 (.L_HI(net1042));
 sg13g2_tiehi _14767__1043 (.L_HI(net1043));
 sg13g2_tiehi _14766__1044 (.L_HI(net1044));
 sg13g2_tiehi _14765__1045 (.L_HI(net1045));
 sg13g2_tiehi _14764__1046 (.L_HI(net1046));
 sg13g2_tiehi _14763__1047 (.L_HI(net1047));
 sg13g2_tiehi _14762__1048 (.L_HI(net1048));
 sg13g2_tiehi _14761__1049 (.L_HI(net1049));
 sg13g2_tiehi _14760__1050 (.L_HI(net1050));
 sg13g2_tiehi _14759__1051 (.L_HI(net1051));
 sg13g2_tiehi _14758__1052 (.L_HI(net1052));
 sg13g2_tiehi _14757__1053 (.L_HI(net1053));
 sg13g2_tiehi _14756__1054 (.L_HI(net1054));
 sg13g2_tiehi _14755__1055 (.L_HI(net1055));
 sg13g2_tiehi _14754__1056 (.L_HI(net1056));
 sg13g2_tiehi _14753__1057 (.L_HI(net1057));
 sg13g2_tiehi _14752__1058 (.L_HI(net1058));
 sg13g2_tiehi _14751__1059 (.L_HI(net1059));
 sg13g2_tiehi _14750__1060 (.L_HI(net1060));
 sg13g2_tiehi _14749__1061 (.L_HI(net1061));
 sg13g2_tiehi _14748__1062 (.L_HI(net1062));
 sg13g2_tiehi _14747__1063 (.L_HI(net1063));
 sg13g2_tiehi _14746__1064 (.L_HI(net1064));
 sg13g2_tiehi _14745__1065 (.L_HI(net1065));
 sg13g2_tiehi _14744__1066 (.L_HI(net1066));
 sg13g2_tiehi _14743__1067 (.L_HI(net1067));
 sg13g2_tiehi _14742__1068 (.L_HI(net1068));
 sg13g2_tiehi _14741__1069 (.L_HI(net1069));
 sg13g2_tiehi _14740__1070 (.L_HI(net1070));
 sg13g2_tiehi _14739__1071 (.L_HI(net1071));
 sg13g2_tiehi _14738__1072 (.L_HI(net1072));
 sg13g2_tiehi _14737__1073 (.L_HI(net1073));
 sg13g2_tiehi _14736__1074 (.L_HI(net1074));
 sg13g2_tiehi _14735__1075 (.L_HI(net1075));
 sg13g2_tiehi _14734__1076 (.L_HI(net1076));
 sg13g2_tiehi _14733__1077 (.L_HI(net1077));
 sg13g2_tiehi _14732__1078 (.L_HI(net1078));
 sg13g2_tiehi _14731__1079 (.L_HI(net1079));
 sg13g2_tiehi _14730__1080 (.L_HI(net1080));
 sg13g2_tiehi _14729__1081 (.L_HI(net1081));
 sg13g2_tiehi _14728__1082 (.L_HI(net1082));
 sg13g2_tiehi _14727__1083 (.L_HI(net1083));
 sg13g2_tiehi _14726__1084 (.L_HI(net1084));
 sg13g2_tiehi _14725__1085 (.L_HI(net1085));
 sg13g2_tiehi _14724__1086 (.L_HI(net1086));
 sg13g2_tiehi _14723__1087 (.L_HI(net1087));
 sg13g2_tiehi _14722__1088 (.L_HI(net1088));
 sg13g2_tiehi _14721__1089 (.L_HI(net1089));
 sg13g2_tiehi _14720__1090 (.L_HI(net1090));
 sg13g2_tiehi _14719__1091 (.L_HI(net1091));
 sg13g2_tiehi _14718__1092 (.L_HI(net1092));
 sg13g2_tiehi _14717__1093 (.L_HI(net1093));
 sg13g2_tiehi _14716__1094 (.L_HI(net1094));
 sg13g2_tiehi _14715__1095 (.L_HI(net1095));
 sg13g2_tiehi _14714__1096 (.L_HI(net1096));
 sg13g2_tiehi _14713__1097 (.L_HI(net1097));
 sg13g2_tiehi _14712__1098 (.L_HI(net1098));
 sg13g2_tiehi _14711__1099 (.L_HI(net1099));
 sg13g2_tiehi _14710__1100 (.L_HI(net1100));
 sg13g2_tiehi _14709__1101 (.L_HI(net1101));
 sg13g2_tiehi _14708__1102 (.L_HI(net1102));
 sg13g2_tiehi _14707__1103 (.L_HI(net1103));
 sg13g2_tiehi _14706__1104 (.L_HI(net1104));
 sg13g2_tiehi _14705__1105 (.L_HI(net1105));
 sg13g2_tiehi _14704__1106 (.L_HI(net1106));
 sg13g2_tiehi _14703__1107 (.L_HI(net1107));
 sg13g2_tiehi _14702__1108 (.L_HI(net1108));
 sg13g2_tiehi _14701__1109 (.L_HI(net1109));
 sg13g2_tiehi _14700__1110 (.L_HI(net1110));
 sg13g2_tiehi _14699__1111 (.L_HI(net1111));
 sg13g2_tiehi _14698__1112 (.L_HI(net1112));
 sg13g2_tiehi _14697__1113 (.L_HI(net1113));
 sg13g2_tiehi _14696__1114 (.L_HI(net1114));
 sg13g2_tiehi _14695__1115 (.L_HI(net1115));
 sg13g2_tiehi _14694__1116 (.L_HI(net1116));
 sg13g2_tiehi _14693__1117 (.L_HI(net1117));
 sg13g2_tiehi _14692__1118 (.L_HI(net1118));
 sg13g2_tiehi _14691__1119 (.L_HI(net1119));
 sg13g2_tiehi _14690__1120 (.L_HI(net1120));
 sg13g2_tiehi _14689__1121 (.L_HI(net1121));
 sg13g2_tiehi _14688__1122 (.L_HI(net1122));
 sg13g2_tiehi _14687__1123 (.L_HI(net1123));
 sg13g2_tiehi _14686__1124 (.L_HI(net1124));
 sg13g2_tiehi _14685__1125 (.L_HI(net1125));
 sg13g2_tiehi _14684__1126 (.L_HI(net1126));
 sg13g2_tiehi _14683__1127 (.L_HI(net1127));
 sg13g2_tiehi _14682__1128 (.L_HI(net1128));
 sg13g2_tiehi _14681__1129 (.L_HI(net1129));
 sg13g2_tiehi _14680__1130 (.L_HI(net1130));
 sg13g2_tiehi _14679__1131 (.L_HI(net1131));
 sg13g2_tiehi _14678__1132 (.L_HI(net1132));
 sg13g2_tiehi _14677__1133 (.L_HI(net1133));
 sg13g2_tiehi _14676__1134 (.L_HI(net1134));
 sg13g2_tiehi _14675__1135 (.L_HI(net1135));
 sg13g2_tiehi _14674__1136 (.L_HI(net1136));
 sg13g2_tiehi _14673__1137 (.L_HI(net1137));
 sg13g2_tiehi _14672__1138 (.L_HI(net1138));
 sg13g2_tiehi _14671__1139 (.L_HI(net1139));
 sg13g2_tiehi _14670__1140 (.L_HI(net1140));
 sg13g2_tiehi _14669__1141 (.L_HI(net1141));
 sg13g2_tiehi _14668__1142 (.L_HI(net1142));
 sg13g2_tiehi _14667__1143 (.L_HI(net1143));
 sg13g2_tiehi _14666__1144 (.L_HI(net1144));
 sg13g2_tiehi _14665__1145 (.L_HI(net1145));
 sg13g2_tiehi _14664__1146 (.L_HI(net1146));
 sg13g2_tiehi _14663__1147 (.L_HI(net1147));
 sg13g2_tiehi _14662__1148 (.L_HI(net1148));
 sg13g2_tiehi _14661__1149 (.L_HI(net1149));
 sg13g2_tiehi _14660__1150 (.L_HI(net1150));
 sg13g2_tiehi _14659__1151 (.L_HI(net1151));
 sg13g2_tiehi _14658__1152 (.L_HI(net1152));
 sg13g2_tiehi _14657__1153 (.L_HI(net1153));
 sg13g2_tiehi _14656__1154 (.L_HI(net1154));
 sg13g2_tiehi _14655__1155 (.L_HI(net1155));
 sg13g2_tiehi _14654__1156 (.L_HI(net1156));
 sg13g2_tiehi _14653__1157 (.L_HI(net1157));
 sg13g2_tiehi _14652__1158 (.L_HI(net1158));
 sg13g2_tiehi _14651__1159 (.L_HI(net1159));
 sg13g2_tiehi _14650__1160 (.L_HI(net1160));
 sg13g2_tiehi _14649__1161 (.L_HI(net1161));
 sg13g2_tiehi _14648__1162 (.L_HI(net1162));
 sg13g2_tiehi _14647__1163 (.L_HI(net1163));
 sg13g2_tiehi _14646__1164 (.L_HI(net1164));
 sg13g2_tiehi _14645__1165 (.L_HI(net1165));
 sg13g2_tiehi _14644__1166 (.L_HI(net1166));
 sg13g2_tiehi _14643__1167 (.L_HI(net1167));
 sg13g2_tiehi _14642__1168 (.L_HI(net1168));
 sg13g2_tiehi _14641__1169 (.L_HI(net1169));
 sg13g2_tiehi _14640__1170 (.L_HI(net1170));
 sg13g2_tiehi _14639__1171 (.L_HI(net1171));
 sg13g2_tiehi _14638__1172 (.L_HI(net1172));
 sg13g2_tiehi _14637__1173 (.L_HI(net1173));
 sg13g2_tiehi _14636__1174 (.L_HI(net1174));
 sg13g2_tiehi _14635__1175 (.L_HI(net1175));
 sg13g2_tiehi _14634__1176 (.L_HI(net1176));
 sg13g2_tiehi _14633__1177 (.L_HI(net1177));
 sg13g2_tiehi _14632__1178 (.L_HI(net1178));
 sg13g2_tiehi _14631__1179 (.L_HI(net1179));
 sg13g2_tiehi _14630__1180 (.L_HI(net1180));
 sg13g2_tiehi _14629__1181 (.L_HI(net1181));
 sg13g2_tiehi _14628__1182 (.L_HI(net1182));
 sg13g2_tiehi _14627__1183 (.L_HI(net1183));
 sg13g2_tiehi _14626__1184 (.L_HI(net1184));
 sg13g2_tiehi _14625__1185 (.L_HI(net1185));
 sg13g2_tiehi _14624__1186 (.L_HI(net1186));
 sg13g2_tiehi _14623__1187 (.L_HI(net1187));
 sg13g2_tiehi _14622__1188 (.L_HI(net1188));
 sg13g2_tiehi _14621__1189 (.L_HI(net1189));
 sg13g2_tiehi _14620__1190 (.L_HI(net1190));
 sg13g2_tiehi _14619__1191 (.L_HI(net1191));
 sg13g2_tiehi _14618__1192 (.L_HI(net1192));
 sg13g2_tiehi _14617__1193 (.L_HI(net1193));
 sg13g2_tiehi _14616__1194 (.L_HI(net1194));
 sg13g2_tiehi _14615__1195 (.L_HI(net1195));
 sg13g2_tiehi _14614__1196 (.L_HI(net1196));
 sg13g2_tiehi _14613__1197 (.L_HI(net1197));
 sg13g2_tiehi _14612__1198 (.L_HI(net1198));
 sg13g2_tiehi _14611__1199 (.L_HI(net1199));
 sg13g2_tiehi _14610__1200 (.L_HI(net1200));
 sg13g2_tiehi _14609__1201 (.L_HI(net1201));
 sg13g2_tiehi _14608__1202 (.L_HI(net1202));
 sg13g2_tiehi _14607__1203 (.L_HI(net1203));
 sg13g2_tiehi _14606__1204 (.L_HI(net1204));
 sg13g2_tiehi _14605__1205 (.L_HI(net1205));
 sg13g2_tiehi _14604__1206 (.L_HI(net1206));
 sg13g2_tiehi _14603__1207 (.L_HI(net1207));
 sg13g2_tiehi _14602__1208 (.L_HI(net1208));
 sg13g2_tiehi _14601__1209 (.L_HI(net1209));
 sg13g2_tiehi _14600__1210 (.L_HI(net1210));
 sg13g2_tiehi _14599__1211 (.L_HI(net1211));
 sg13g2_tiehi _14598__1212 (.L_HI(net1212));
 sg13g2_tiehi _14597__1213 (.L_HI(net1213));
 sg13g2_tiehi _14596__1214 (.L_HI(net1214));
 sg13g2_tiehi _14595__1215 (.L_HI(net1215));
 sg13g2_tiehi _14594__1216 (.L_HI(net1216));
 sg13g2_tiehi _14593__1217 (.L_HI(net1217));
 sg13g2_tiehi _14592__1218 (.L_HI(net1218));
 sg13g2_tiehi _14591__1219 (.L_HI(net1219));
 sg13g2_tiehi _14590__1220 (.L_HI(net1220));
 sg13g2_tiehi _14589__1221 (.L_HI(net1221));
 sg13g2_tiehi _14588__1222 (.L_HI(net1222));
 sg13g2_tiehi _14587__1223 (.L_HI(net1223));
 sg13g2_tiehi _14586__1224 (.L_HI(net1224));
 sg13g2_tiehi _14585__1225 (.L_HI(net1225));
 sg13g2_tiehi _14584__1226 (.L_HI(net1226));
 sg13g2_tiehi _14583__1227 (.L_HI(net1227));
 sg13g2_tiehi _14582__1228 (.L_HI(net1228));
 sg13g2_tiehi _14581__1229 (.L_HI(net1229));
 sg13g2_tiehi _14580__1230 (.L_HI(net1230));
 sg13g2_tiehi _14579__1231 (.L_HI(net1231));
 sg13g2_tiehi _14578__1232 (.L_HI(net1232));
 sg13g2_tiehi _14577__1233 (.L_HI(net1233));
 sg13g2_tiehi _14576__1234 (.L_HI(net1234));
 sg13g2_tiehi _14575__1235 (.L_HI(net1235));
 sg13g2_tiehi _14574__1236 (.L_HI(net1236));
 sg13g2_tiehi _14573__1237 (.L_HI(net1237));
 sg13g2_tiehi _14572__1238 (.L_HI(net1238));
 sg13g2_tiehi _16605__1239 (.L_HI(net1239));
 sg13g2_tiehi _16604__1240 (.L_HI(net1240));
 sg13g2_tiehi _16603__1241 (.L_HI(net1241));
 sg13g2_tiehi _16602__1242 (.L_HI(net1242));
 sg13g2_tiehi _16601__1243 (.L_HI(net1243));
 sg13g2_tiehi _16600__1244 (.L_HI(net1244));
 sg13g2_tiehi _16599__1245 (.L_HI(net1245));
 sg13g2_tiehi _16598__1246 (.L_HI(net1246));
 sg13g2_tiehi _16597__1247 (.L_HI(net1247));
 sg13g2_tiehi _16596__1248 (.L_HI(net1248));
 sg13g2_tiehi _16595__1249 (.L_HI(net1249));
 sg13g2_tiehi _16594__1250 (.L_HI(net1250));
 sg13g2_tiehi _16593__1251 (.L_HI(net1251));
 sg13g2_tiehi _16592__1252 (.L_HI(net1252));
 sg13g2_tiehi _16591__1253 (.L_HI(net1253));
 sg13g2_tiehi _16590__1254 (.L_HI(net1254));
 sg13g2_tiehi _16589__1255 (.L_HI(net1255));
 sg13g2_tiehi _16588__1256 (.L_HI(net1256));
 sg13g2_tiehi _16587__1257 (.L_HI(net1257));
 sg13g2_tiehi _16586__1258 (.L_HI(net1258));
 sg13g2_tiehi _16585__1259 (.L_HI(net1259));
 sg13g2_tiehi _16584__1260 (.L_HI(net1260));
 sg13g2_tiehi _16583__1261 (.L_HI(net1261));
 sg13g2_tiehi _16582__1262 (.L_HI(net1262));
 sg13g2_tiehi _16581__1263 (.L_HI(net1263));
 sg13g2_tiehi _16580__1264 (.L_HI(net1264));
 sg13g2_tiehi _16579__1265 (.L_HI(net1265));
 sg13g2_tiehi _16578__1266 (.L_HI(net1266));
 sg13g2_tiehi _16577__1267 (.L_HI(net1267));
 sg13g2_tiehi _16576__1268 (.L_HI(net1268));
 sg13g2_tiehi _16575__1269 (.L_HI(net1269));
 sg13g2_tiehi _16574__1270 (.L_HI(net1270));
 sg13g2_tiehi _16573__1271 (.L_HI(net1271));
 sg13g2_tiehi _16572__1272 (.L_HI(net1272));
 sg13g2_tiehi _16571__1273 (.L_HI(net1273));
 sg13g2_tiehi _16570__1274 (.L_HI(net1274));
 sg13g2_tiehi _16569__1275 (.L_HI(net1275));
 sg13g2_tiehi _16568__1276 (.L_HI(net1276));
 sg13g2_tiehi _16567__1277 (.L_HI(net1277));
 sg13g2_tiehi _16566__1278 (.L_HI(net1278));
 sg13g2_tiehi _16565__1279 (.L_HI(net1279));
 sg13g2_tiehi _16564__1280 (.L_HI(net1280));
 sg13g2_tiehi _16563__1281 (.L_HI(net1281));
 sg13g2_tiehi _16562__1282 (.L_HI(net1282));
 sg13g2_tiehi _16561__1283 (.L_HI(net1283));
 sg13g2_tiehi _16560__1284 (.L_HI(net1284));
 sg13g2_tiehi _16559__1285 (.L_HI(net1285));
 sg13g2_tiehi _16558__1286 (.L_HI(net1286));
 sg13g2_tiehi _16557__1287 (.L_HI(net1287));
 sg13g2_tiehi _16556__1288 (.L_HI(net1288));
 sg13g2_tiehi _16555__1289 (.L_HI(net1289));
 sg13g2_tiehi _16554__1290 (.L_HI(net1290));
 sg13g2_tiehi _16553__1291 (.L_HI(net1291));
 sg13g2_tiehi _16552__1292 (.L_HI(net1292));
 sg13g2_tiehi _16551__1293 (.L_HI(net1293));
 sg13g2_tiehi _16550__1294 (.L_HI(net1294));
 sg13g2_tiehi _16549__1295 (.L_HI(net1295));
 sg13g2_tiehi _16548__1296 (.L_HI(net1296));
 sg13g2_tiehi _16547__1297 (.L_HI(net1297));
 sg13g2_tiehi _16546__1298 (.L_HI(net1298));
 sg13g2_tiehi _16545__1299 (.L_HI(net1299));
 sg13g2_tiehi _16544__1300 (.L_HI(net1300));
 sg13g2_tiehi _16543__1301 (.L_HI(net1301));
 sg13g2_tiehi _16542__1302 (.L_HI(net1302));
 sg13g2_tiehi _16541__1303 (.L_HI(net1303));
 sg13g2_tiehi _16540__1304 (.L_HI(net1304));
 sg13g2_tiehi _16539__1305 (.L_HI(net1305));
 sg13g2_tiehi _16538__1306 (.L_HI(net1306));
 sg13g2_tiehi _16537__1307 (.L_HI(net1307));
 sg13g2_tiehi _16536__1308 (.L_HI(net1308));
 sg13g2_tiehi _16535__1309 (.L_HI(net1309));
 sg13g2_tiehi _16534__1310 (.L_HI(net1310));
 sg13g2_tiehi _16533__1311 (.L_HI(net1311));
 sg13g2_tiehi _16532__1312 (.L_HI(net1312));
 sg13g2_tiehi _16531__1313 (.L_HI(net1313));
 sg13g2_tiehi _16530__1314 (.L_HI(net1314));
 sg13g2_tiehi _16529__1315 (.L_HI(net1315));
 sg13g2_tiehi _16528__1316 (.L_HI(net1316));
 sg13g2_tiehi _16527__1317 (.L_HI(net1317));
 sg13g2_tiehi _16526__1318 (.L_HI(net1318));
 sg13g2_tiehi _16525__1319 (.L_HI(net1319));
 sg13g2_tiehi _16524__1320 (.L_HI(net1320));
 sg13g2_tiehi _16523__1321 (.L_HI(net1321));
 sg13g2_tiehi _16522__1322 (.L_HI(net1322));
 sg13g2_tiehi _16521__1323 (.L_HI(net1323));
 sg13g2_tiehi _16520__1324 (.L_HI(net1324));
 sg13g2_tiehi _16519__1325 (.L_HI(net1325));
 sg13g2_tiehi _16518__1326 (.L_HI(net1326));
 sg13g2_tiehi _16517__1327 (.L_HI(net1327));
 sg13g2_tiehi _16516__1328 (.L_HI(net1328));
 sg13g2_tiehi _16515__1329 (.L_HI(net1329));
 sg13g2_tiehi _16514__1330 (.L_HI(net1330));
 sg13g2_tiehi _16513__1331 (.L_HI(net1331));
 sg13g2_tiehi _16512__1332 (.L_HI(net1332));
 sg13g2_tiehi _16511__1333 (.L_HI(net1333));
 sg13g2_tiehi _16510__1334 (.L_HI(net1334));
 sg13g2_tiehi _16509__1335 (.L_HI(net1335));
 sg13g2_tiehi _16508__1336 (.L_HI(net1336));
 sg13g2_tiehi _16507__1337 (.L_HI(net1337));
 sg13g2_tiehi _16506__1338 (.L_HI(net1338));
 sg13g2_tiehi _16505__1339 (.L_HI(net1339));
 sg13g2_tiehi _16504__1340 (.L_HI(net1340));
 sg13g2_tiehi _16503__1341 (.L_HI(net1341));
 sg13g2_tiehi _16502__1342 (.L_HI(net1342));
 sg13g2_tiehi _16501__1343 (.L_HI(net1343));
 sg13g2_tiehi _16500__1344 (.L_HI(net1344));
 sg13g2_tiehi _16499__1345 (.L_HI(net1345));
 sg13g2_tiehi _16498__1346 (.L_HI(net1346));
 sg13g2_tiehi _16497__1347 (.L_HI(net1347));
 sg13g2_tiehi _16496__1348 (.L_HI(net1348));
 sg13g2_tiehi _16495__1349 (.L_HI(net1349));
 sg13g2_tiehi _16494__1350 (.L_HI(net1350));
 sg13g2_tiehi _16493__1351 (.L_HI(net1351));
 sg13g2_tiehi _16492__1352 (.L_HI(net1352));
 sg13g2_tiehi _16491__1353 (.L_HI(net1353));
 sg13g2_tiehi _16490__1354 (.L_HI(net1354));
 sg13g2_tiehi _16489__1355 (.L_HI(net1355));
 sg13g2_tiehi _16488__1356 (.L_HI(net1356));
 sg13g2_tiehi _16487__1357 (.L_HI(net1357));
 sg13g2_tiehi _16486__1358 (.L_HI(net1358));
 sg13g2_tiehi _16485__1359 (.L_HI(net1359));
 sg13g2_tiehi _16484__1360 (.L_HI(net1360));
 sg13g2_tiehi _16483__1361 (.L_HI(net1361));
 sg13g2_tiehi _16482__1362 (.L_HI(net1362));
 sg13g2_tiehi _16481__1363 (.L_HI(net1363));
 sg13g2_tiehi _16480__1364 (.L_HI(net1364));
 sg13g2_tiehi _16479__1365 (.L_HI(net1365));
 sg13g2_tiehi _16478__1366 (.L_HI(net1366));
 sg13g2_tiehi _16477__1367 (.L_HI(net1367));
 sg13g2_tiehi _16476__1368 (.L_HI(net1368));
 sg13g2_tiehi _16475__1369 (.L_HI(net1369));
 sg13g2_tiehi _16474__1370 (.L_HI(net1370));
 sg13g2_tiehi _16473__1371 (.L_HI(net1371));
 sg13g2_tiehi _16472__1372 (.L_HI(net1372));
 sg13g2_tiehi _16471__1373 (.L_HI(net1373));
 sg13g2_tiehi _16470__1374 (.L_HI(net1374));
 sg13g2_tiehi _16469__1375 (.L_HI(net1375));
 sg13g2_tiehi _16468__1376 (.L_HI(net1376));
 sg13g2_tiehi _16467__1377 (.L_HI(net1377));
 sg13g2_tiehi _16466__1378 (.L_HI(net1378));
 sg13g2_tiehi _16465__1379 (.L_HI(net1379));
 sg13g2_tiehi _16464__1380 (.L_HI(net1380));
 sg13g2_tiehi _16463__1381 (.L_HI(net1381));
 sg13g2_tiehi _16462__1382 (.L_HI(net1382));
 sg13g2_tiehi _16461__1383 (.L_HI(net1383));
 sg13g2_tiehi _16460__1384 (.L_HI(net1384));
 sg13g2_tiehi _16459__1385 (.L_HI(net1385));
 sg13g2_tiehi _16458__1386 (.L_HI(net1386));
 sg13g2_tiehi _16457__1387 (.L_HI(net1387));
 sg13g2_tiehi _16456__1388 (.L_HI(net1388));
 sg13g2_tiehi _16455__1389 (.L_HI(net1389));
 sg13g2_tiehi _16454__1390 (.L_HI(net1390));
 sg13g2_tiehi _16453__1391 (.L_HI(net1391));
 sg13g2_tiehi _16452__1392 (.L_HI(net1392));
 sg13g2_tiehi _16451__1393 (.L_HI(net1393));
 sg13g2_tiehi _16450__1394 (.L_HI(net1394));
 sg13g2_tiehi _16449__1395 (.L_HI(net1395));
 sg13g2_tiehi _16448__1396 (.L_HI(net1396));
 sg13g2_tiehi _16447__1397 (.L_HI(net1397));
 sg13g2_tiehi _16446__1398 (.L_HI(net1398));
 sg13g2_tiehi _16445__1399 (.L_HI(net1399));
 sg13g2_tiehi _16444__1400 (.L_HI(net1400));
 sg13g2_tiehi _16443__1401 (.L_HI(net1401));
 sg13g2_tiehi _16442__1402 (.L_HI(net1402));
 sg13g2_tiehi _16441__1403 (.L_HI(net1403));
 sg13g2_tiehi _16440__1404 (.L_HI(net1404));
 sg13g2_tiehi _16439__1405 (.L_HI(net1405));
 sg13g2_tiehi _16438__1406 (.L_HI(net1406));
 sg13g2_tiehi _16437__1407 (.L_HI(net1407));
 sg13g2_tiehi _16436__1408 (.L_HI(net1408));
 sg13g2_tiehi _16435__1409 (.L_HI(net1409));
 sg13g2_tiehi _16434__1410 (.L_HI(net1410));
 sg13g2_tiehi _16433__1411 (.L_HI(net1411));
 sg13g2_tiehi _16432__1412 (.L_HI(net1412));
 sg13g2_tiehi _16431__1413 (.L_HI(net1413));
 sg13g2_tiehi _16430__1414 (.L_HI(net1414));
 sg13g2_tiehi _16429__1415 (.L_HI(net1415));
 sg13g2_tiehi _16428__1416 (.L_HI(net1416));
 sg13g2_tiehi _16427__1417 (.L_HI(net1417));
 sg13g2_tiehi _16426__1418 (.L_HI(net1418));
 sg13g2_tiehi _16425__1419 (.L_HI(net1419));
 sg13g2_tiehi _16424__1420 (.L_HI(net1420));
 sg13g2_tiehi _16423__1421 (.L_HI(net1421));
 sg13g2_tiehi _16422__1422 (.L_HI(net1422));
 sg13g2_tiehi _16421__1423 (.L_HI(net1423));
 sg13g2_tiehi _16420__1424 (.L_HI(net1424));
 sg13g2_tiehi _16419__1425 (.L_HI(net1425));
 sg13g2_tiehi _16418__1426 (.L_HI(net1426));
 sg13g2_tiehi _16417__1427 (.L_HI(net1427));
 sg13g2_tiehi _16416__1428 (.L_HI(net1428));
 sg13g2_tiehi _16415__1429 (.L_HI(net1429));
 sg13g2_tiehi _16414__1430 (.L_HI(net1430));
 sg13g2_tiehi _16413__1431 (.L_HI(net1431));
 sg13g2_tiehi _16412__1432 (.L_HI(net1432));
 sg13g2_tiehi _16411__1433 (.L_HI(net1433));
 sg13g2_tiehi _16410__1434 (.L_HI(net1434));
 sg13g2_tiehi _16409__1435 (.L_HI(net1435));
 sg13g2_tiehi _16408__1436 (.L_HI(net1436));
 sg13g2_tiehi _16407__1437 (.L_HI(net1437));
 sg13g2_tiehi _16406__1438 (.L_HI(net1438));
 sg13g2_tiehi _16405__1439 (.L_HI(net1439));
 sg13g2_tiehi _16404__1440 (.L_HI(net1440));
 sg13g2_tiehi _16403__1441 (.L_HI(net1441));
 sg13g2_tiehi _16402__1442 (.L_HI(net1442));
 sg13g2_tiehi _16401__1443 (.L_HI(net1443));
 sg13g2_tiehi _16400__1444 (.L_HI(net1444));
 sg13g2_tiehi _16399__1445 (.L_HI(net1445));
 sg13g2_tiehi _16398__1446 (.L_HI(net1446));
 sg13g2_tiehi _16397__1447 (.L_HI(net1447));
 sg13g2_tiehi _16396__1448 (.L_HI(net1448));
 sg13g2_tiehi _16395__1449 (.L_HI(net1449));
 sg13g2_tiehi _16394__1450 (.L_HI(net1450));
 sg13g2_tiehi _16393__1451 (.L_HI(net1451));
 sg13g2_tiehi _16392__1452 (.L_HI(net1452));
 sg13g2_tiehi _16391__1453 (.L_HI(net1453));
 sg13g2_tiehi _16390__1454 (.L_HI(net1454));
 sg13g2_tiehi _16389__1455 (.L_HI(net1455));
 sg13g2_tiehi _16388__1456 (.L_HI(net1456));
 sg13g2_tiehi _16387__1457 (.L_HI(net1457));
 sg13g2_tiehi _16386__1458 (.L_HI(net1458));
 sg13g2_tiehi _16385__1459 (.L_HI(net1459));
 sg13g2_tiehi _16384__1460 (.L_HI(net1460));
 sg13g2_tiehi _16383__1461 (.L_HI(net1461));
 sg13g2_tiehi _16382__1462 (.L_HI(net1462));
 sg13g2_tiehi _16381__1463 (.L_HI(net1463));
 sg13g2_tiehi _16380__1464 (.L_HI(net1464));
 sg13g2_tiehi _16379__1465 (.L_HI(net1465));
 sg13g2_tiehi _16378__1466 (.L_HI(net1466));
 sg13g2_tiehi _16377__1467 (.L_HI(net1467));
 sg13g2_tiehi _16376__1468 (.L_HI(net1468));
 sg13g2_tiehi _16375__1469 (.L_HI(net1469));
 sg13g2_tiehi _16374__1470 (.L_HI(net1470));
 sg13g2_tiehi _16373__1471 (.L_HI(net1471));
 sg13g2_tiehi _16372__1472 (.L_HI(net1472));
 sg13g2_tiehi _16371__1473 (.L_HI(net1473));
 sg13g2_tiehi _16370__1474 (.L_HI(net1474));
 sg13g2_tiehi _16369__1475 (.L_HI(net1475));
 sg13g2_tiehi _16368__1476 (.L_HI(net1476));
 sg13g2_tiehi _16367__1477 (.L_HI(net1477));
 sg13g2_tiehi _16366__1478 (.L_HI(net1478));
 sg13g2_tiehi _16365__1479 (.L_HI(net1479));
 sg13g2_tiehi _16364__1480 (.L_HI(net1480));
 sg13g2_tiehi _16363__1481 (.L_HI(net1481));
 sg13g2_tiehi _16362__1482 (.L_HI(net1482));
 sg13g2_tiehi _16361__1483 (.L_HI(net1483));
 sg13g2_tiehi _16360__1484 (.L_HI(net1484));
 sg13g2_tiehi _16359__1485 (.L_HI(net1485));
 sg13g2_tiehi _16358__1486 (.L_HI(net1486));
 sg13g2_tiehi _16357__1487 (.L_HI(net1487));
 sg13g2_tiehi _16356__1488 (.L_HI(net1488));
 sg13g2_tiehi _16355__1489 (.L_HI(net1489));
 sg13g2_tiehi _16354__1490 (.L_HI(net1490));
 sg13g2_tiehi _16353__1491 (.L_HI(net1491));
 sg13g2_tiehi _16352__1492 (.L_HI(net1492));
 sg13g2_tiehi _16351__1493 (.L_HI(net1493));
 sg13g2_tiehi _16350__1494 (.L_HI(net1494));
 sg13g2_tiehi _16349__1495 (.L_HI(net1495));
 sg13g2_tiehi _16348__1496 (.L_HI(net1496));
 sg13g2_tiehi _16347__1497 (.L_HI(net1497));
 sg13g2_tiehi _16346__1498 (.L_HI(net1498));
 sg13g2_tiehi _16345__1499 (.L_HI(net1499));
 sg13g2_tiehi _16344__1500 (.L_HI(net1500));
 sg13g2_tiehi _16343__1501 (.L_HI(net1501));
 sg13g2_tiehi _16342__1502 (.L_HI(net1502));
 sg13g2_tiehi _16341__1503 (.L_HI(net1503));
 sg13g2_tiehi _16340__1504 (.L_HI(net1504));
 sg13g2_tiehi _16339__1505 (.L_HI(net1505));
 sg13g2_tiehi _16338__1506 (.L_HI(net1506));
 sg13g2_tiehi _16337__1507 (.L_HI(net1507));
 sg13g2_tiehi _16336__1508 (.L_HI(net1508));
 sg13g2_tiehi _16335__1509 (.L_HI(net1509));
 sg13g2_tiehi _16334__1510 (.L_HI(net1510));
 sg13g2_tiehi _16333__1511 (.L_HI(net1511));
 sg13g2_tiehi _16332__1512 (.L_HI(net1512));
 sg13g2_tiehi _16331__1513 (.L_HI(net1513));
 sg13g2_tiehi _16330__1514 (.L_HI(net1514));
 sg13g2_tiehi _16329__1515 (.L_HI(net1515));
 sg13g2_tiehi _16328__1516 (.L_HI(net1516));
 sg13g2_tiehi _16327__1517 (.L_HI(net1517));
 sg13g2_tiehi _16326__1518 (.L_HI(net1518));
 sg13g2_tiehi _16325__1519 (.L_HI(net1519));
 sg13g2_tiehi _16324__1520 (.L_HI(net1520));
 sg13g2_tiehi _16323__1521 (.L_HI(net1521));
 sg13g2_tiehi _16322__1522 (.L_HI(net1522));
 sg13g2_tiehi _16321__1523 (.L_HI(net1523));
 sg13g2_tiehi _16320__1524 (.L_HI(net1524));
 sg13g2_tiehi _16319__1525 (.L_HI(net1525));
 sg13g2_tiehi _16318__1526 (.L_HI(net1526));
 sg13g2_tiehi _16317__1527 (.L_HI(net1527));
 sg13g2_tiehi _16316__1528 (.L_HI(net1528));
 sg13g2_tiehi _16315__1529 (.L_HI(net1529));
 sg13g2_tiehi _16314__1530 (.L_HI(net1530));
 sg13g2_tiehi _16313__1531 (.L_HI(net1531));
 sg13g2_tiehi _16312__1532 (.L_HI(net1532));
 sg13g2_tiehi _16311__1533 (.L_HI(net1533));
 sg13g2_tiehi _16310__1534 (.L_HI(net1534));
 sg13g2_tiehi _16309__1535 (.L_HI(net1535));
 sg13g2_tiehi _16308__1536 (.L_HI(net1536));
 sg13g2_tiehi _16307__1537 (.L_HI(net1537));
 sg13g2_tiehi _16306__1538 (.L_HI(net1538));
 sg13g2_tiehi _16305__1539 (.L_HI(net1539));
 sg13g2_tiehi _16304__1540 (.L_HI(net1540));
 sg13g2_tiehi _16303__1541 (.L_HI(net1541));
 sg13g2_tiehi _16302__1542 (.L_HI(net1542));
 sg13g2_tiehi _16301__1543 (.L_HI(net1543));
 sg13g2_tiehi _16300__1544 (.L_HI(net1544));
 sg13g2_tiehi _16299__1545 (.L_HI(net1545));
 sg13g2_tiehi _16298__1546 (.L_HI(net1546));
 sg13g2_tiehi _16297__1547 (.L_HI(net1547));
 sg13g2_tiehi _16296__1548 (.L_HI(net1548));
 sg13g2_tiehi _16295__1549 (.L_HI(net1549));
 sg13g2_tiehi _16294__1550 (.L_HI(net1550));
 sg13g2_tiehi _16293__1551 (.L_HI(net1551));
 sg13g2_tiehi _16292__1552 (.L_HI(net1552));
 sg13g2_tiehi _16291__1553 (.L_HI(net1553));
 sg13g2_tiehi _16290__1554 (.L_HI(net1554));
 sg13g2_tiehi _16289__1555 (.L_HI(net1555));
 sg13g2_tiehi _16288__1556 (.L_HI(net1556));
 sg13g2_tiehi _16287__1557 (.L_HI(net1557));
 sg13g2_tiehi _16286__1558 (.L_HI(net1558));
 sg13g2_tiehi _16285__1559 (.L_HI(net1559));
 sg13g2_tiehi _16284__1560 (.L_HI(net1560));
 sg13g2_tiehi _16283__1561 (.L_HI(net1561));
 sg13g2_tiehi _16282__1562 (.L_HI(net1562));
 sg13g2_tiehi _16281__1563 (.L_HI(net1563));
 sg13g2_tiehi _16280__1564 (.L_HI(net1564));
 sg13g2_tiehi _16279__1565 (.L_HI(net1565));
 sg13g2_tiehi _16278__1566 (.L_HI(net1566));
 sg13g2_tiehi _16277__1567 (.L_HI(net1567));
 sg13g2_tiehi _16276__1568 (.L_HI(net1568));
 sg13g2_tiehi _16275__1569 (.L_HI(net1569));
 sg13g2_tiehi _16274__1570 (.L_HI(net1570));
 sg13g2_tiehi _16273__1571 (.L_HI(net1571));
 sg13g2_tiehi _16272__1572 (.L_HI(net1572));
 sg13g2_tiehi _16271__1573 (.L_HI(net1573));
 sg13g2_tiehi _16270__1574 (.L_HI(net1574));
 sg13g2_tiehi _16269__1575 (.L_HI(net1575));
 sg13g2_tiehi _16268__1576 (.L_HI(net1576));
 sg13g2_tiehi _16267__1577 (.L_HI(net1577));
 sg13g2_tiehi _16266__1578 (.L_HI(net1578));
 sg13g2_tiehi _16265__1579 (.L_HI(net1579));
 sg13g2_tiehi _16264__1580 (.L_HI(net1580));
 sg13g2_tiehi _16263__1581 (.L_HI(net1581));
 sg13g2_tiehi _16262__1582 (.L_HI(net1582));
 sg13g2_tiehi _16261__1583 (.L_HI(net1583));
 sg13g2_tiehi _16260__1584 (.L_HI(net1584));
 sg13g2_tiehi _16259__1585 (.L_HI(net1585));
 sg13g2_tiehi _16258__1586 (.L_HI(net1586));
 sg13g2_tiehi _16257__1587 (.L_HI(net1587));
 sg13g2_tiehi _16256__1588 (.L_HI(net1588));
 sg13g2_tiehi _16255__1589 (.L_HI(net1589));
 sg13g2_tiehi _16254__1590 (.L_HI(net1590));
 sg13g2_tiehi _16253__1591 (.L_HI(net1591));
 sg13g2_tiehi _16252__1592 (.L_HI(net1592));
 sg13g2_tiehi _16251__1593 (.L_HI(net1593));
 sg13g2_tiehi _16250__1594 (.L_HI(net1594));
 sg13g2_tiehi _16249__1595 (.L_HI(net1595));
 sg13g2_tiehi _16248__1596 (.L_HI(net1596));
 sg13g2_tiehi _16247__1597 (.L_HI(net1597));
 sg13g2_tiehi _16246__1598 (.L_HI(net1598));
 sg13g2_tiehi _16245__1599 (.L_HI(net1599));
 sg13g2_tiehi _16244__1600 (.L_HI(net1600));
 sg13g2_tiehi _16243__1601 (.L_HI(net1601));
 sg13g2_tiehi _16242__1602 (.L_HI(net1602));
 sg13g2_tiehi _16241__1603 (.L_HI(net1603));
 sg13g2_tiehi _16240__1604 (.L_HI(net1604));
 sg13g2_tiehi _16239__1605 (.L_HI(net1605));
 sg13g2_tiehi _16238__1606 (.L_HI(net1606));
 sg13g2_tiehi _16237__1607 (.L_HI(net1607));
 sg13g2_tiehi _16236__1608 (.L_HI(net1608));
 sg13g2_tiehi _16235__1609 (.L_HI(net1609));
 sg13g2_tiehi _16234__1610 (.L_HI(net1610));
 sg13g2_tiehi _16233__1611 (.L_HI(net1611));
 sg13g2_tiehi _16232__1612 (.L_HI(net1612));
 sg13g2_tiehi _16231__1613 (.L_HI(net1613));
 sg13g2_tiehi _16230__1614 (.L_HI(net1614));
 sg13g2_tiehi _16229__1615 (.L_HI(net1615));
 sg13g2_tiehi _16228__1616 (.L_HI(net1616));
 sg13g2_tiehi _16227__1617 (.L_HI(net1617));
 sg13g2_tiehi _16226__1618 (.L_HI(net1618));
 sg13g2_tiehi _16225__1619 (.L_HI(net1619));
 sg13g2_tiehi _16224__1620 (.L_HI(net1620));
 sg13g2_tiehi _16223__1621 (.L_HI(net1621));
 sg13g2_tiehi _16222__1622 (.L_HI(net1622));
 sg13g2_tiehi _16221__1623 (.L_HI(net1623));
 sg13g2_tiehi _16220__1624 (.L_HI(net1624));
 sg13g2_tiehi _16219__1625 (.L_HI(net1625));
 sg13g2_tiehi _16218__1626 (.L_HI(net1626));
 sg13g2_tiehi _16217__1627 (.L_HI(net1627));
 sg13g2_tiehi _16216__1628 (.L_HI(net1628));
 sg13g2_tiehi _16215__1629 (.L_HI(net1629));
 sg13g2_tiehi _16214__1630 (.L_HI(net1630));
 sg13g2_tiehi _16213__1631 (.L_HI(net1631));
 sg13g2_tiehi _16212__1632 (.L_HI(net1632));
 sg13g2_tiehi _16211__1633 (.L_HI(net1633));
 sg13g2_tiehi _16210__1634 (.L_HI(net1634));
 sg13g2_tiehi _16209__1635 (.L_HI(net1635));
 sg13g2_tiehi _16208__1636 (.L_HI(net1636));
 sg13g2_tiehi _16207__1637 (.L_HI(net1637));
 sg13g2_tiehi _16206__1638 (.L_HI(net1638));
 sg13g2_tiehi _16205__1639 (.L_HI(net1639));
 sg13g2_tiehi _16204__1640 (.L_HI(net1640));
 sg13g2_tiehi _16203__1641 (.L_HI(net1641));
 sg13g2_tiehi _16202__1642 (.L_HI(net1642));
 sg13g2_tiehi _16201__1643 (.L_HI(net1643));
 sg13g2_tiehi _16200__1644 (.L_HI(net1644));
 sg13g2_tiehi _16199__1645 (.L_HI(net1645));
 sg13g2_tiehi _16198__1646 (.L_HI(net1646));
 sg13g2_tiehi _16197__1647 (.L_HI(net1647));
 sg13g2_tiehi _16196__1648 (.L_HI(net1648));
 sg13g2_tiehi _16195__1649 (.L_HI(net1649));
 sg13g2_tiehi _16194__1650 (.L_HI(net1650));
 sg13g2_tiehi _16193__1651 (.L_HI(net1651));
 sg13g2_tiehi _16192__1652 (.L_HI(net1652));
 sg13g2_tiehi _16191__1653 (.L_HI(net1653));
 sg13g2_tiehi _16190__1654 (.L_HI(net1654));
 sg13g2_tiehi _16189__1655 (.L_HI(net1655));
 sg13g2_tiehi _16188__1656 (.L_HI(net1656));
 sg13g2_tiehi _16187__1657 (.L_HI(net1657));
 sg13g2_tiehi _16186__1658 (.L_HI(net1658));
 sg13g2_tiehi _16185__1659 (.L_HI(net1659));
 sg13g2_tiehi _16184__1660 (.L_HI(net1660));
 sg13g2_tiehi _16183__1661 (.L_HI(net1661));
 sg13g2_tiehi _16182__1662 (.L_HI(net1662));
 sg13g2_tiehi _16181__1663 (.L_HI(net1663));
 sg13g2_tiehi _16180__1664 (.L_HI(net1664));
 sg13g2_tiehi _16179__1665 (.L_HI(net1665));
 sg13g2_tiehi _16178__1666 (.L_HI(net1666));
 sg13g2_tiehi _16177__1667 (.L_HI(net1667));
 sg13g2_tiehi _16176__1668 (.L_HI(net1668));
 sg13g2_tiehi _16175__1669 (.L_HI(net1669));
 sg13g2_tiehi _16174__1670 (.L_HI(net1670));
 sg13g2_tiehi _16173__1671 (.L_HI(net1671));
 sg13g2_tiehi _16172__1672 (.L_HI(net1672));
 sg13g2_tiehi _16171__1673 (.L_HI(net1673));
 sg13g2_tiehi _16170__1674 (.L_HI(net1674));
 sg13g2_tiehi _16169__1675 (.L_HI(net1675));
 sg13g2_tiehi _16168__1676 (.L_HI(net1676));
 sg13g2_tiehi _16167__1677 (.L_HI(net1677));
 sg13g2_tiehi _16166__1678 (.L_HI(net1678));
 sg13g2_tiehi _16165__1679 (.L_HI(net1679));
 sg13g2_tiehi _16164__1680 (.L_HI(net1680));
 sg13g2_tiehi _16163__1681 (.L_HI(net1681));
 sg13g2_tiehi _16162__1682 (.L_HI(net1682));
 sg13g2_tiehi _16161__1683 (.L_HI(net1683));
 sg13g2_tiehi _16160__1684 (.L_HI(net1684));
 sg13g2_tiehi _16159__1685 (.L_HI(net1685));
 sg13g2_tiehi _16158__1686 (.L_HI(net1686));
 sg13g2_tiehi _16157__1687 (.L_HI(net1687));
 sg13g2_tiehi _16156__1688 (.L_HI(net1688));
 sg13g2_tiehi _16155__1689 (.L_HI(net1689));
 sg13g2_tiehi _16154__1690 (.L_HI(net1690));
 sg13g2_tiehi _16153__1691 (.L_HI(net1691));
 sg13g2_tiehi _16152__1692 (.L_HI(net1692));
 sg13g2_tiehi _16151__1693 (.L_HI(net1693));
 sg13g2_tiehi _16150__1694 (.L_HI(net1694));
 sg13g2_tiehi _16149__1695 (.L_HI(net1695));
 sg13g2_tiehi _16148__1696 (.L_HI(net1696));
 sg13g2_tiehi _16147__1697 (.L_HI(net1697));
 sg13g2_tiehi _16146__1698 (.L_HI(net1698));
 sg13g2_tiehi _16145__1699 (.L_HI(net1699));
 sg13g2_tiehi _16144__1700 (.L_HI(net1700));
 sg13g2_tiehi _16143__1701 (.L_HI(net1701));
 sg13g2_tiehi _16142__1702 (.L_HI(net1702));
 sg13g2_tiehi _16141__1703 (.L_HI(net1703));
 sg13g2_tiehi _16140__1704 (.L_HI(net1704));
 sg13g2_tiehi _16139__1705 (.L_HI(net1705));
 sg13g2_tiehi _16138__1706 (.L_HI(net1706));
 sg13g2_tiehi _16137__1707 (.L_HI(net1707));
 sg13g2_tiehi _16136__1708 (.L_HI(net1708));
 sg13g2_tiehi _16135__1709 (.L_HI(net1709));
 sg13g2_tiehi _16134__1710 (.L_HI(net1710));
 sg13g2_tiehi _16133__1711 (.L_HI(net1711));
 sg13g2_tiehi _16132__1712 (.L_HI(net1712));
 sg13g2_tiehi _16131__1713 (.L_HI(net1713));
 sg13g2_tiehi _16130__1714 (.L_HI(net1714));
 sg13g2_tiehi _16129__1715 (.L_HI(net1715));
 sg13g2_tiehi _16128__1716 (.L_HI(net1716));
 sg13g2_tiehi _16127__1717 (.L_HI(net1717));
 sg13g2_tiehi _16126__1718 (.L_HI(net1718));
 sg13g2_tiehi _16125__1719 (.L_HI(net1719));
 sg13g2_tiehi _16124__1720 (.L_HI(net1720));
 sg13g2_tiehi _16123__1721 (.L_HI(net1721));
 sg13g2_tiehi _16122__1722 (.L_HI(net1722));
 sg13g2_tiehi _16121__1723 (.L_HI(net1723));
 sg13g2_tiehi _16120__1724 (.L_HI(net1724));
 sg13g2_tiehi _16119__1725 (.L_HI(net1725));
 sg13g2_tiehi _16118__1726 (.L_HI(net1726));
 sg13g2_tiehi _16117__1727 (.L_HI(net1727));
 sg13g2_tiehi _16116__1728 (.L_HI(net1728));
 sg13g2_tiehi _16115__1729 (.L_HI(net1729));
 sg13g2_tiehi _16114__1730 (.L_HI(net1730));
 sg13g2_tiehi _16113__1731 (.L_HI(net1731));
 sg13g2_tiehi _16112__1732 (.L_HI(net1732));
 sg13g2_tiehi _16111__1733 (.L_HI(net1733));
 sg13g2_tiehi _16110__1734 (.L_HI(net1734));
 sg13g2_tiehi _16109__1735 (.L_HI(net1735));
 sg13g2_tiehi _16108__1736 (.L_HI(net1736));
 sg13g2_tiehi _16107__1737 (.L_HI(net1737));
 sg13g2_tiehi _16106__1738 (.L_HI(net1738));
 sg13g2_tiehi _16105__1739 (.L_HI(net1739));
 sg13g2_tiehi _16104__1740 (.L_HI(net1740));
 sg13g2_tiehi _16103__1741 (.L_HI(net1741));
 sg13g2_tiehi _16102__1742 (.L_HI(net1742));
 sg13g2_tiehi _16101__1743 (.L_HI(net1743));
 sg13g2_tiehi _16100__1744 (.L_HI(net1744));
 sg13g2_tiehi _16099__1745 (.L_HI(net1745));
 sg13g2_tiehi _16098__1746 (.L_HI(net1746));
 sg13g2_tiehi _16097__1747 (.L_HI(net1747));
 sg13g2_tiehi _16096__1748 (.L_HI(net1748));
 sg13g2_tiehi _16095__1749 (.L_HI(net1749));
 sg13g2_tiehi _16094__1750 (.L_HI(net1750));
 sg13g2_tiehi _16093__1751 (.L_HI(net1751));
 sg13g2_tiehi _16092__1752 (.L_HI(net1752));
 sg13g2_tiehi _16091__1753 (.L_HI(net1753));
 sg13g2_tiehi _16090__1754 (.L_HI(net1754));
 sg13g2_tiehi _16089__1755 (.L_HI(net1755));
 sg13g2_tiehi _16088__1756 (.L_HI(net1756));
 sg13g2_tiehi _16087__1757 (.L_HI(net1757));
 sg13g2_tiehi _16086__1758 (.L_HI(net1758));
 sg13g2_tiehi _16085__1759 (.L_HI(net1759));
 sg13g2_tiehi _16084__1760 (.L_HI(net1760));
 sg13g2_tiehi _16083__1761 (.L_HI(net1761));
 sg13g2_tiehi _16082__1762 (.L_HI(net1762));
 sg13g2_tiehi _16081__1763 (.L_HI(net1763));
 sg13g2_tiehi _16080__1764 (.L_HI(net1764));
 sg13g2_tiehi _16079__1765 (.L_HI(net1765));
 sg13g2_tiehi _16078__1766 (.L_HI(net1766));
 sg13g2_tiehi _16077__1767 (.L_HI(net1767));
 sg13g2_tiehi _16076__1768 (.L_HI(net1768));
 sg13g2_tiehi _16075__1769 (.L_HI(net1769));
 sg13g2_tiehi _16074__1770 (.L_HI(net1770));
 sg13g2_tiehi _16073__1771 (.L_HI(net1771));
 sg13g2_tiehi _16072__1772 (.L_HI(net1772));
 sg13g2_tiehi _16071__1773 (.L_HI(net1773));
 sg13g2_tiehi _16070__1774 (.L_HI(net1774));
 sg13g2_tiehi _16069__1775 (.L_HI(net1775));
 sg13g2_tiehi _16068__1776 (.L_HI(net1776));
 sg13g2_tiehi _16067__1777 (.L_HI(net1777));
 sg13g2_tiehi _16066__1778 (.L_HI(net1778));
 sg13g2_tiehi _16065__1779 (.L_HI(net1779));
 sg13g2_tiehi _16064__1780 (.L_HI(net1780));
 sg13g2_tiehi _16063__1781 (.L_HI(net1781));
 sg13g2_tiehi _16062__1782 (.L_HI(net1782));
 sg13g2_tiehi _16061__1783 (.L_HI(net1783));
 sg13g2_tiehi _16060__1784 (.L_HI(net1784));
 sg13g2_tiehi _16059__1785 (.L_HI(net1785));
 sg13g2_tiehi _16058__1786 (.L_HI(net1786));
 sg13g2_tiehi _16057__1787 (.L_HI(net1787));
 sg13g2_tiehi _16056__1788 (.L_HI(net1788));
 sg13g2_tiehi _16055__1789 (.L_HI(net1789));
 sg13g2_tiehi _16054__1790 (.L_HI(net1790));
 sg13g2_tiehi _16053__1791 (.L_HI(net1791));
 sg13g2_tiehi _16052__1792 (.L_HI(net1792));
 sg13g2_tiehi _16051__1793 (.L_HI(net1793));
 sg13g2_tiehi _16050__1794 (.L_HI(net1794));
 sg13g2_tiehi _16049__1795 (.L_HI(net1795));
 sg13g2_tiehi _16048__1796 (.L_HI(net1796));
 sg13g2_tiehi _16047__1797 (.L_HI(net1797));
 sg13g2_tiehi _16046__1798 (.L_HI(net1798));
 sg13g2_tiehi _16045__1799 (.L_HI(net1799));
 sg13g2_tiehi _16044__1800 (.L_HI(net1800));
 sg13g2_tiehi _16043__1801 (.L_HI(net1801));
 sg13g2_tiehi _16042__1802 (.L_HI(net1802));
 sg13g2_tiehi _16041__1803 (.L_HI(net1803));
 sg13g2_tiehi _16040__1804 (.L_HI(net1804));
 sg13g2_tiehi _16039__1805 (.L_HI(net1805));
 sg13g2_tiehi _16038__1806 (.L_HI(net1806));
 sg13g2_tiehi _16037__1807 (.L_HI(net1807));
 sg13g2_tiehi _16036__1808 (.L_HI(net1808));
 sg13g2_tiehi _16035__1809 (.L_HI(net1809));
 sg13g2_tiehi _16034__1810 (.L_HI(net1810));
 sg13g2_tiehi _16033__1811 (.L_HI(net1811));
 sg13g2_tiehi _16032__1812 (.L_HI(net1812));
 sg13g2_tiehi _16031__1813 (.L_HI(net1813));
 sg13g2_tiehi _16030__1814 (.L_HI(net1814));
 sg13g2_tiehi _16029__1815 (.L_HI(net1815));
 sg13g2_tiehi _16028__1816 (.L_HI(net1816));
 sg13g2_tiehi _16027__1817 (.L_HI(net1817));
 sg13g2_tiehi _16026__1818 (.L_HI(net1818));
 sg13g2_tiehi _16025__1819 (.L_HI(net1819));
 sg13g2_tiehi _16024__1820 (.L_HI(net1820));
 sg13g2_tiehi _16023__1821 (.L_HI(net1821));
 sg13g2_tiehi _16022__1822 (.L_HI(net1822));
 sg13g2_tiehi _16021__1823 (.L_HI(net1823));
 sg13g2_tiehi _16020__1824 (.L_HI(net1824));
 sg13g2_tiehi _16019__1825 (.L_HI(net1825));
 sg13g2_tiehi _16018__1826 (.L_HI(net1826));
 sg13g2_tiehi _16017__1827 (.L_HI(net1827));
 sg13g2_tiehi _16016__1828 (.L_HI(net1828));
 sg13g2_tiehi _16015__1829 (.L_HI(net1829));
 sg13g2_tiehi _16014__1830 (.L_HI(net1830));
 sg13g2_tiehi _16013__1831 (.L_HI(net1831));
 sg13g2_tiehi _16012__1832 (.L_HI(net1832));
 sg13g2_tiehi _16011__1833 (.L_HI(net1833));
 sg13g2_tiehi _16010__1834 (.L_HI(net1834));
 sg13g2_tiehi _16009__1835 (.L_HI(net1835));
 sg13g2_tiehi _16008__1836 (.L_HI(net1836));
 sg13g2_tiehi _16007__1837 (.L_HI(net1837));
 sg13g2_tiehi _16006__1838 (.L_HI(net1838));
 sg13g2_tiehi _16005__1839 (.L_HI(net1839));
 sg13g2_tiehi _16004__1840 (.L_HI(net1840));
 sg13g2_tiehi _16003__1841 (.L_HI(net1841));
 sg13g2_tiehi _16002__1842 (.L_HI(net1842));
 sg13g2_tiehi _16001__1843 (.L_HI(net1843));
 sg13g2_tiehi _16000__1844 (.L_HI(net1844));
 sg13g2_tiehi _15999__1845 (.L_HI(net1845));
 sg13g2_tiehi _15998__1846 (.L_HI(net1846));
 sg13g2_tiehi _15997__1847 (.L_HI(net1847));
 sg13g2_tiehi _15996__1848 (.L_HI(net1848));
 sg13g2_tiehi _15995__1849 (.L_HI(net1849));
 sg13g2_tiehi _15994__1850 (.L_HI(net1850));
 sg13g2_tiehi _15993__1851 (.L_HI(net1851));
 sg13g2_tiehi _15992__1852 (.L_HI(net1852));
 sg13g2_tiehi _15991__1853 (.L_HI(net1853));
 sg13g2_tiehi _15990__1854 (.L_HI(net1854));
 sg13g2_tiehi _15989__1855 (.L_HI(net1855));
 sg13g2_tiehi _15988__1856 (.L_HI(net1856));
 sg13g2_tiehi _15987__1857 (.L_HI(net1857));
 sg13g2_tiehi _15986__1858 (.L_HI(net1858));
 sg13g2_tiehi _15985__1859 (.L_HI(net1859));
 sg13g2_tiehi _15984__1860 (.L_HI(net1860));
 sg13g2_tiehi _15983__1861 (.L_HI(net1861));
 sg13g2_tiehi _15982__1862 (.L_HI(net1862));
 sg13g2_tiehi _15981__1863 (.L_HI(net1863));
 sg13g2_tiehi _15980__1864 (.L_HI(net1864));
 sg13g2_tiehi _15979__1865 (.L_HI(net1865));
 sg13g2_tiehi _15978__1866 (.L_HI(net1866));
 sg13g2_tiehi _15977__1867 (.L_HI(net1867));
 sg13g2_tiehi _15976__1868 (.L_HI(net1868));
 sg13g2_tiehi _15975__1869 (.L_HI(net1869));
 sg13g2_tiehi _15974__1870 (.L_HI(net1870));
 sg13g2_tiehi _15973__1871 (.L_HI(net1871));
 sg13g2_tiehi _15972__1872 (.L_HI(net1872));
 sg13g2_tiehi _15971__1873 (.L_HI(net1873));
 sg13g2_tiehi _15970__1874 (.L_HI(net1874));
 sg13g2_tiehi _15969__1875 (.L_HI(net1875));
 sg13g2_tiehi _15968__1876 (.L_HI(net1876));
 sg13g2_tiehi _15967__1877 (.L_HI(net1877));
 sg13g2_tiehi _15966__1878 (.L_HI(net1878));
 sg13g2_tiehi _15965__1879 (.L_HI(net1879));
 sg13g2_tiehi _15964__1880 (.L_HI(net1880));
 sg13g2_tiehi _15963__1881 (.L_HI(net1881));
 sg13g2_tiehi _15962__1882 (.L_HI(net1882));
 sg13g2_tiehi _15961__1883 (.L_HI(net1883));
 sg13g2_tiehi _15960__1884 (.L_HI(net1884));
 sg13g2_tiehi _15959__1885 (.L_HI(net1885));
 sg13g2_tiehi _15958__1886 (.L_HI(net1886));
 sg13g2_tiehi _15957__1887 (.L_HI(net1887));
 sg13g2_tiehi _15956__1888 (.L_HI(net1888));
 sg13g2_tiehi _15955__1889 (.L_HI(net1889));
 sg13g2_tiehi _15954__1890 (.L_HI(net1890));
 sg13g2_tiehi _15953__1891 (.L_HI(net1891));
 sg13g2_tiehi _15952__1892 (.L_HI(net1892));
 sg13g2_tiehi _15951__1893 (.L_HI(net1893));
 sg13g2_tiehi _15950__1894 (.L_HI(net1894));
 sg13g2_tiehi _15949__1895 (.L_HI(net1895));
 sg13g2_tiehi _15948__1896 (.L_HI(net1896));
 sg13g2_tiehi _15947__1897 (.L_HI(net1897));
 sg13g2_tiehi _15946__1898 (.L_HI(net1898));
 sg13g2_tiehi _15945__1899 (.L_HI(net1899));
 sg13g2_tiehi _15944__1900 (.L_HI(net1900));
 sg13g2_tiehi _15943__1901 (.L_HI(net1901));
 sg13g2_tiehi _15942__1902 (.L_HI(net1902));
 sg13g2_tiehi _15941__1903 (.L_HI(net1903));
 sg13g2_tiehi _15940__1904 (.L_HI(net1904));
 sg13g2_tiehi _15939__1905 (.L_HI(net1905));
 sg13g2_tiehi _15938__1906 (.L_HI(net1906));
 sg13g2_tiehi _15937__1907 (.L_HI(net1907));
 sg13g2_tiehi _15936__1908 (.L_HI(net1908));
 sg13g2_tiehi _15935__1909 (.L_HI(net1909));
 sg13g2_tiehi _15934__1910 (.L_HI(net1910));
 sg13g2_tiehi _15933__1911 (.L_HI(net1911));
 sg13g2_tiehi _15932__1912 (.L_HI(net1912));
 sg13g2_tiehi _15931__1913 (.L_HI(net1913));
 sg13g2_tiehi _15930__1914 (.L_HI(net1914));
 sg13g2_tiehi _15929__1915 (.L_HI(net1915));
 sg13g2_tiehi _15928__1916 (.L_HI(net1916));
 sg13g2_tiehi _15927__1917 (.L_HI(net1917));
 sg13g2_tiehi _15926__1918 (.L_HI(net1918));
 sg13g2_tiehi _15925__1919 (.L_HI(net1919));
 sg13g2_tiehi _15924__1920 (.L_HI(net1920));
 sg13g2_tiehi _15923__1921 (.L_HI(net1921));
 sg13g2_tiehi _15922__1922 (.L_HI(net1922));
 sg13g2_tiehi _15921__1923 (.L_HI(net1923));
 sg13g2_tiehi _15920__1924 (.L_HI(net1924));
 sg13g2_tiehi _15919__1925 (.L_HI(net1925));
 sg13g2_tiehi _15918__1926 (.L_HI(net1926));
 sg13g2_tiehi _15917__1927 (.L_HI(net1927));
 sg13g2_tiehi _15916__1928 (.L_HI(net1928));
 sg13g2_tiehi _15915__1929 (.L_HI(net1929));
 sg13g2_tiehi _15914__1930 (.L_HI(net1930));
 sg13g2_tiehi _15913__1931 (.L_HI(net1931));
 sg13g2_tiehi _15912__1932 (.L_HI(net1932));
 sg13g2_tiehi _15911__1933 (.L_HI(net1933));
 sg13g2_tiehi _15910__1934 (.L_HI(net1934));
 sg13g2_tiehi _15909__1935 (.L_HI(net1935));
 sg13g2_tiehi _15908__1936 (.L_HI(net1936));
 sg13g2_tiehi _15907__1937 (.L_HI(net1937));
 sg13g2_tiehi _15906__1938 (.L_HI(net1938));
 sg13g2_tiehi _15905__1939 (.L_HI(net1939));
 sg13g2_tiehi _15904__1940 (.L_HI(net1940));
 sg13g2_tiehi _15903__1941 (.L_HI(net1941));
 sg13g2_tiehi _15902__1942 (.L_HI(net1942));
 sg13g2_tiehi _15901__1943 (.L_HI(net1943));
 sg13g2_tiehi _15900__1944 (.L_HI(net1944));
 sg13g2_tiehi _15899__1945 (.L_HI(net1945));
 sg13g2_tiehi _15898__1946 (.L_HI(net1946));
 sg13g2_tiehi _15897__1947 (.L_HI(net1947));
 sg13g2_tiehi _15896__1948 (.L_HI(net1948));
 sg13g2_tiehi _15895__1949 (.L_HI(net1949));
 sg13g2_tiehi _15894__1950 (.L_HI(net1950));
 sg13g2_tiehi _15893__1951 (.L_HI(net1951));
 sg13g2_tiehi _15892__1952 (.L_HI(net1952));
 sg13g2_tiehi _15891__1953 (.L_HI(net1953));
 sg13g2_tiehi _15890__1954 (.L_HI(net1954));
 sg13g2_tiehi _15889__1955 (.L_HI(net1955));
 sg13g2_tiehi _15888__1956 (.L_HI(net1956));
 sg13g2_tiehi _15887__1957 (.L_HI(net1957));
 sg13g2_tiehi _15886__1958 (.L_HI(net1958));
 sg13g2_tiehi _15885__1959 (.L_HI(net1959));
 sg13g2_tiehi _15884__1960 (.L_HI(net1960));
 sg13g2_tiehi _15883__1961 (.L_HI(net1961));
 sg13g2_tiehi _15882__1962 (.L_HI(net1962));
 sg13g2_tiehi _15881__1963 (.L_HI(net1963));
 sg13g2_tiehi _15880__1964 (.L_HI(net1964));
 sg13g2_tiehi _15879__1965 (.L_HI(net1965));
 sg13g2_tiehi _15878__1966 (.L_HI(net1966));
 sg13g2_tiehi _15877__1967 (.L_HI(net1967));
 sg13g2_tiehi _15876__1968 (.L_HI(net1968));
 sg13g2_tiehi _15875__1969 (.L_HI(net1969));
 sg13g2_tiehi _15874__1970 (.L_HI(net1970));
 sg13g2_tiehi _15873__1971 (.L_HI(net1971));
 sg13g2_tiehi _15872__1972 (.L_HI(net1972));
 sg13g2_tiehi _15871__1973 (.L_HI(net1973));
 sg13g2_tiehi _15870__1974 (.L_HI(net1974));
 sg13g2_tiehi _15869__1975 (.L_HI(net1975));
 sg13g2_tiehi _15868__1976 (.L_HI(net1976));
 sg13g2_tiehi _15867__1977 (.L_HI(net1977));
 sg13g2_tiehi _15866__1978 (.L_HI(net1978));
 sg13g2_tiehi _15865__1979 (.L_HI(net1979));
 sg13g2_tiehi _15864__1980 (.L_HI(net1980));
 sg13g2_tiehi _15863__1981 (.L_HI(net1981));
 sg13g2_tiehi _15862__1982 (.L_HI(net1982));
 sg13g2_tiehi _15861__1983 (.L_HI(net1983));
 sg13g2_tiehi _15860__1984 (.L_HI(net1984));
 sg13g2_tiehi _15859__1985 (.L_HI(net1985));
 sg13g2_tiehi _15858__1986 (.L_HI(net1986));
 sg13g2_tiehi _15857__1987 (.L_HI(net1987));
 sg13g2_tiehi _15856__1988 (.L_HI(net1988));
 sg13g2_tiehi _15855__1989 (.L_HI(net1989));
 sg13g2_tiehi _15854__1990 (.L_HI(net1990));
 sg13g2_tiehi _15853__1991 (.L_HI(net1991));
 sg13g2_tiehi _15852__1992 (.L_HI(net1992));
 sg13g2_tiehi _15851__1993 (.L_HI(net1993));
 sg13g2_tiehi _15850__1994 (.L_HI(net1994));
 sg13g2_tiehi _15849__1995 (.L_HI(net1995));
 sg13g2_tiehi _15848__1996 (.L_HI(net1996));
 sg13g2_tiehi _15847__1997 (.L_HI(net1997));
 sg13g2_tiehi _15846__1998 (.L_HI(net1998));
 sg13g2_tiehi _15845__1999 (.L_HI(net1999));
 sg13g2_tiehi _15844__2000 (.L_HI(net2000));
 sg13g2_tiehi _15843__2001 (.L_HI(net2001));
 sg13g2_tiehi _15842__2002 (.L_HI(net2002));
 sg13g2_tiehi _15841__2003 (.L_HI(net2003));
 sg13g2_tiehi _15840__2004 (.L_HI(net2004));
 sg13g2_tiehi _15839__2005 (.L_HI(net2005));
 sg13g2_tiehi _15838__2006 (.L_HI(net2006));
 sg13g2_tiehi _15837__2007 (.L_HI(net2007));
 sg13g2_tiehi _15836__2008 (.L_HI(net2008));
 sg13g2_tiehi _15835__2009 (.L_HI(net2009));
 sg13g2_tiehi _15834__2010 (.L_HI(net2010));
 sg13g2_tiehi _15833__2011 (.L_HI(net2011));
 sg13g2_tiehi _15832__2012 (.L_HI(net2012));
 sg13g2_tiehi _15831__2013 (.L_HI(net2013));
 sg13g2_tiehi _15830__2014 (.L_HI(net2014));
 sg13g2_tiehi _15829__2015 (.L_HI(net2015));
 sg13g2_tiehi _15828__2016 (.L_HI(net2016));
 sg13g2_tiehi _15827__2017 (.L_HI(net2017));
 sg13g2_tiehi _15826__2018 (.L_HI(net2018));
 sg13g2_tiehi _15825__2019 (.L_HI(net2019));
 sg13g2_tiehi _15824__2020 (.L_HI(net2020));
 sg13g2_tiehi _15823__2021 (.L_HI(net2021));
 sg13g2_tiehi _15822__2022 (.L_HI(net2022));
 sg13g2_tiehi _15821__2023 (.L_HI(net2023));
 sg13g2_tiehi _15820__2024 (.L_HI(net2024));
 sg13g2_tiehi _15819__2025 (.L_HI(net2025));
 sg13g2_tiehi _15818__2026 (.L_HI(net2026));
 sg13g2_tiehi _15817__2027 (.L_HI(net2027));
 sg13g2_tiehi _15816__2028 (.L_HI(net2028));
 sg13g2_tiehi _15815__2029 (.L_HI(net2029));
 sg13g2_tiehi _15814__2030 (.L_HI(net2030));
 sg13g2_tiehi _15813__2031 (.L_HI(net2031));
 sg13g2_tiehi _15812__2032 (.L_HI(net2032));
 sg13g2_tiehi _15811__2033 (.L_HI(net2033));
 sg13g2_tiehi _15810__2034 (.L_HI(net2034));
 sg13g2_tiehi _15809__2035 (.L_HI(net2035));
 sg13g2_tiehi _15808__2036 (.L_HI(net2036));
 sg13g2_tiehi _15807__2037 (.L_HI(net2037));
 sg13g2_tiehi _15806__2038 (.L_HI(net2038));
 sg13g2_tiehi _15805__2039 (.L_HI(net2039));
 sg13g2_tiehi _15804__2040 (.L_HI(net2040));
 sg13g2_tiehi _15803__2041 (.L_HI(net2041));
 sg13g2_tiehi _15802__2042 (.L_HI(net2042));
 sg13g2_tiehi _15801__2043 (.L_HI(net2043));
 sg13g2_tiehi _15800__2044 (.L_HI(net2044));
 sg13g2_tiehi _15799__2045 (.L_HI(net2045));
 sg13g2_tiehi _15798__2046 (.L_HI(net2046));
 sg13g2_tiehi _15797__2047 (.L_HI(net2047));
 sg13g2_tiehi _15796__2048 (.L_HI(net2048));
 sg13g2_tiehi _15795__2049 (.L_HI(net2049));
 sg13g2_tiehi _15794__2050 (.L_HI(net2050));
 sg13g2_tiehi _15793__2051 (.L_HI(net2051));
 sg13g2_tiehi _15792__2052 (.L_HI(net2052));
 sg13g2_tiehi _15791__2053 (.L_HI(net2053));
 sg13g2_tiehi _15790__2054 (.L_HI(net2054));
 sg13g2_tiehi _15789__2055 (.L_HI(net2055));
 sg13g2_tiehi _15788__2056 (.L_HI(net2056));
 sg13g2_tiehi _15787__2057 (.L_HI(net2057));
 sg13g2_tiehi _15786__2058 (.L_HI(net2058));
 sg13g2_tiehi _15785__2059 (.L_HI(net2059));
 sg13g2_tiehi _15784__2060 (.L_HI(net2060));
 sg13g2_tiehi _15783__2061 (.L_HI(net2061));
 sg13g2_tiehi _15782__2062 (.L_HI(net2062));
 sg13g2_tiehi _15781__2063 (.L_HI(net2063));
 sg13g2_tiehi _15780__2064 (.L_HI(net2064));
 sg13g2_tiehi _15779__2065 (.L_HI(net2065));
 sg13g2_tiehi _15778__2066 (.L_HI(net2066));
 sg13g2_tiehi _15777__2067 (.L_HI(net2067));
 sg13g2_tiehi _15776__2068 (.L_HI(net2068));
 sg13g2_tiehi _15775__2069 (.L_HI(net2069));
 sg13g2_tiehi _15774__2070 (.L_HI(net2070));
 sg13g2_tiehi _15773__2071 (.L_HI(net2071));
 sg13g2_tiehi _15772__2072 (.L_HI(net2072));
 sg13g2_tiehi _15771__2073 (.L_HI(net2073));
 sg13g2_tiehi _15770__2074 (.L_HI(net2074));
 sg13g2_tiehi _15769__2075 (.L_HI(net2075));
 sg13g2_tiehi _15768__2076 (.L_HI(net2076));
 sg13g2_tiehi _15767__2077 (.L_HI(net2077));
 sg13g2_tiehi _15766__2078 (.L_HI(net2078));
 sg13g2_tiehi _15765__2079 (.L_HI(net2079));
 sg13g2_tiehi _15764__2080 (.L_HI(net2080));
 sg13g2_tiehi _15763__2081 (.L_HI(net2081));
 sg13g2_tiehi _15762__2082 (.L_HI(net2082));
 sg13g2_tiehi _15761__2083 (.L_HI(net2083));
 sg13g2_tiehi _15760__2084 (.L_HI(net2084));
 sg13g2_tiehi _15759__2085 (.L_HI(net2085));
 sg13g2_tiehi _15758__2086 (.L_HI(net2086));
 sg13g2_tiehi _15757__2087 (.L_HI(net2087));
 sg13g2_tiehi _15756__2088 (.L_HI(net2088));
 sg13g2_tiehi _15755__2089 (.L_HI(net2089));
 sg13g2_tiehi _15754__2090 (.L_HI(net2090));
 sg13g2_tiehi _15753__2091 (.L_HI(net2091));
 sg13g2_tiehi _15752__2092 (.L_HI(net2092));
 sg13g2_tiehi _15751__2093 (.L_HI(net2093));
 sg13g2_tiehi _15750__2094 (.L_HI(net2094));
 sg13g2_tiehi _15749__2095 (.L_HI(net2095));
 sg13g2_tiehi _15748__2096 (.L_HI(net2096));
 sg13g2_tiehi _15747__2097 (.L_HI(net2097));
 sg13g2_tiehi _15746__2098 (.L_HI(net2098));
 sg13g2_tiehi _15745__2099 (.L_HI(net2099));
 sg13g2_tiehi _15744__2100 (.L_HI(net2100));
 sg13g2_tiehi _15743__2101 (.L_HI(net2101));
 sg13g2_tiehi _15742__2102 (.L_HI(net2102));
 sg13g2_tiehi _15741__2103 (.L_HI(net2103));
 sg13g2_tiehi _15740__2104 (.L_HI(net2104));
 sg13g2_tiehi _15739__2105 (.L_HI(net2105));
 sg13g2_tiehi _15738__2106 (.L_HI(net2106));
 sg13g2_tiehi _15737__2107 (.L_HI(net2107));
 sg13g2_tiehi _15736__2108 (.L_HI(net2108));
 sg13g2_tiehi _15735__2109 (.L_HI(net2109));
 sg13g2_tiehi _15734__2110 (.L_HI(net2110));
 sg13g2_tiehi _15733__2111 (.L_HI(net2111));
 sg13g2_tiehi _15732__2112 (.L_HI(net2112));
 sg13g2_tiehi _15731__2113 (.L_HI(net2113));
 sg13g2_tiehi _15730__2114 (.L_HI(net2114));
 sg13g2_tiehi _15729__2115 (.L_HI(net2115));
 sg13g2_tiehi _15728__2116 (.L_HI(net2116));
 sg13g2_tiehi _15727__2117 (.L_HI(net2117));
 sg13g2_tiehi _15726__2118 (.L_HI(net2118));
 sg13g2_tiehi _15725__2119 (.L_HI(net2119));
 sg13g2_tiehi _15724__2120 (.L_HI(net2120));
 sg13g2_tiehi _15723__2121 (.L_HI(net2121));
 sg13g2_tiehi _15722__2122 (.L_HI(net2122));
 sg13g2_tiehi _15721__2123 (.L_HI(net2123));
 sg13g2_tiehi _15720__2124 (.L_HI(net2124));
 sg13g2_tiehi _15719__2125 (.L_HI(net2125));
 sg13g2_tiehi _15718__2126 (.L_HI(net2126));
 sg13g2_tiehi _15717__2127 (.L_HI(net2127));
 sg13g2_tiehi tt_um_urish_sic1_2128 (.L_HI(net2128));
 sg13g2_tiehi tt_um_urish_sic1_2129 (.L_HI(net2129));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_urish_sic1_15 (.L_LO(net15));
 sg13g2_tielo tt_um_urish_sic1_16 (.L_LO(net16));
 sg13g2_tielo tt_um_urish_sic1_17 (.L_LO(net17));
 sg13g2_tielo tt_um_urish_sic1_18 (.L_LO(net18));
 sg13g2_tielo tt_um_urish_sic1_19 (.L_LO(net19));
 sg13g2_tielo tt_um_urish_sic1_20 (.L_LO(net20));
 sg13g2_tielo tt_um_urish_sic1_21 (.L_LO(net21));
 sg13g2_tielo tt_um_urish_sic1_22 (.L_LO(net22));
 sg13g2_tielo tt_um_urish_sic1_23 (.L_LO(net23));
 sg13g2_tielo tt_um_urish_sic1_24 (.L_LO(net24));
 sg13g2_tielo tt_um_urish_sic1_25 (.L_LO(net25));
 sg13g2_tiehi _15716__26 (.L_HI(net26));
 sg13g2_buf_2 _18789_ (.A(halted),
    .X(uio_out[1]));
 sg13g2_buf_4 _18790_ (.X(uio_out[4]),
    .A(\mem.out_strobe ));
 sg13g2_buf_4 fanout3010 (.X(net3010),
    .A(_05168_));
 sg13g2_buf_4 fanout3011 (.X(net3011),
    .A(_05160_));
 sg13g2_buf_4 fanout3012 (.X(net3012),
    .A(_05127_));
 sg13g2_buf_4 fanout3013 (.X(net3013),
    .A(_05110_));
 sg13g2_buf_4 fanout3014 (.X(net3014),
    .A(_05045_));
 sg13g2_buf_2 fanout3015 (.A(net3016),
    .X(net3015));
 sg13g2_buf_2 fanout3016 (.A(_02518_),
    .X(net3016));
 sg13g2_buf_2 fanout3017 (.A(net3018),
    .X(net3017));
 sg13g2_buf_2 fanout3018 (.A(net3019),
    .X(net3018));
 sg13g2_buf_2 fanout3019 (.A(_02397_),
    .X(net3019));
 sg13g2_buf_4 fanout3020 (.X(net3020),
    .A(_02384_));
 sg13g2_buf_4 fanout3021 (.X(net3021),
    .A(_02342_));
 sg13g2_buf_4 fanout3022 (.X(net3022),
    .A(_02315_));
 sg13g2_buf_4 fanout3023 (.X(net3023),
    .A(_02269_));
 sg13g2_buf_4 fanout3024 (.X(net3024),
    .A(net3026));
 sg13g2_buf_4 fanout3025 (.X(net3025),
    .A(net3026));
 sg13g2_buf_2 fanout3026 (.A(_05013_),
    .X(net3026));
 sg13g2_buf_4 fanout3027 (.X(net3027),
    .A(_02366_));
 sg13g2_buf_2 fanout3028 (.A(_02366_),
    .X(net3028));
 sg13g2_buf_4 fanout3029 (.X(net3029),
    .A(_02363_));
 sg13g2_buf_2 fanout3030 (.A(_02363_),
    .X(net3030));
 sg13g2_buf_4 fanout3031 (.X(net3031),
    .A(_02355_));
 sg13g2_buf_4 fanout3032 (.X(net3032),
    .A(_02355_));
 sg13g2_buf_16 fanout3033 (.X(net3033),
    .A(_02353_));
 sg13g2_buf_4 fanout3034 (.X(net3034),
    .A(_02351_));
 sg13g2_buf_4 fanout3035 (.X(net3035),
    .A(_02351_));
 sg13g2_buf_16 fanout3036 (.X(net3036),
    .A(_02293_));
 sg13g2_buf_4 fanout3037 (.X(net3037),
    .A(_02292_));
 sg13g2_buf_4 fanout3038 (.X(net3038),
    .A(_02292_));
 sg13g2_buf_8 fanout3039 (.A(_02263_),
    .X(net3039));
 sg13g2_buf_4 fanout3040 (.X(net3040),
    .A(_02263_));
 sg13g2_buf_8 fanout3041 (.A(net3044),
    .X(net3041));
 sg13g2_buf_2 fanout3042 (.A(net3044),
    .X(net3042));
 sg13g2_buf_8 fanout3043 (.A(net3044),
    .X(net3043));
 sg13g2_buf_8 fanout3044 (.A(_02262_),
    .X(net3044));
 sg13g2_buf_2 fanout3045 (.A(net3046),
    .X(net3045));
 sg13g2_buf_2 fanout3046 (.A(_05020_),
    .X(net3046));
 sg13g2_buf_2 fanout3047 (.A(net3048),
    .X(net3047));
 sg13g2_buf_2 fanout3048 (.A(_04920_),
    .X(net3048));
 sg13g2_buf_16 fanout3049 (.X(net3049),
    .A(_02310_));
 sg13g2_buf_4 fanout3050 (.X(net3050),
    .A(_02279_));
 sg13g2_buf_4 fanout3051 (.X(net3051),
    .A(_05006_));
 sg13g2_buf_2 fanout3052 (.A(net3053),
    .X(net3052));
 sg13g2_buf_2 fanout3053 (.A(net3054),
    .X(net3053));
 sg13g2_buf_2 fanout3054 (.A(_04850_),
    .X(net3054));
 sg13g2_buf_2 fanout3055 (.A(_02534_),
    .X(net3055));
 sg13g2_buf_2 fanout3056 (.A(net3057),
    .X(net3056));
 sg13g2_buf_2 fanout3057 (.A(net3058),
    .X(net3057));
 sg13g2_buf_2 fanout3058 (.A(_02413_),
    .X(net3058));
 sg13g2_buf_4 fanout3059 (.X(net3059),
    .A(_02408_));
 sg13g2_buf_2 fanout3060 (.A(_02407_),
    .X(net3060));
 sg13g2_buf_2 fanout3061 (.A(_02403_),
    .X(net3061));
 sg13g2_buf_1 fanout3062 (.A(_02403_),
    .X(net3062));
 sg13g2_buf_2 fanout3063 (.A(net3064),
    .X(net3063));
 sg13g2_buf_4 fanout3064 (.X(net3064),
    .A(_02389_));
 sg13g2_buf_8 fanout3065 (.A(_02383_),
    .X(net3065));
 sg13g2_buf_4 fanout3066 (.X(net3066),
    .A(_02379_));
 sg13g2_buf_4 fanout3067 (.X(net3067),
    .A(net3068));
 sg13g2_buf_4 fanout3068 (.X(net3068),
    .A(_02358_));
 sg13g2_buf_16 fanout3069 (.X(net3069),
    .A(_02345_));
 sg13g2_buf_16 fanout3070 (.X(net3070),
    .A(_02334_));
 sg13g2_buf_8 fanout3071 (.A(_02327_),
    .X(net3071));
 sg13g2_buf_16 fanout3072 (.X(net3072),
    .A(_02321_));
 sg13g2_buf_16 fanout3073 (.X(net3073),
    .A(_02318_));
 sg13g2_buf_8 fanout3074 (.A(_02318_),
    .X(net3074));
 sg13g2_buf_4 fanout3075 (.X(net3075),
    .A(_02313_));
 sg13g2_buf_8 fanout3076 (.A(_02307_),
    .X(net3076));
 sg13g2_buf_8 fanout3077 (.A(_02306_),
    .X(net3077));
 sg13g2_buf_4 fanout3078 (.X(net3078),
    .A(_02299_));
 sg13g2_buf_8 fanout3079 (.A(_02282_),
    .X(net3079));
 sg13g2_buf_4 fanout3080 (.X(net3080),
    .A(_02282_));
 sg13g2_buf_8 fanout3081 (.A(_02278_),
    .X(net3081));
 sg13g2_buf_4 fanout3082 (.X(net3082),
    .A(_02274_));
 sg13g2_buf_4 fanout3083 (.X(net3083),
    .A(_02266_));
 sg13g2_buf_8 fanout3084 (.A(_02248_),
    .X(net3084));
 sg13g2_buf_8 fanout3085 (.A(_02248_),
    .X(net3085));
 sg13g2_buf_2 fanout3086 (.A(_02410_),
    .X(net3086));
 sg13g2_buf_4 fanout3087 (.X(net3087),
    .A(_02256_));
 sg13g2_buf_4 fanout3088 (.X(net3088),
    .A(_02252_));
 sg13g2_buf_8 fanout3089 (.A(_02148_),
    .X(net3089));
 sg13g2_buf_4 fanout3090 (.X(net3090),
    .A(net3091));
 sg13g2_buf_8 fanout3091 (.A(_02147_),
    .X(net3091));
 sg13g2_buf_8 fanout3092 (.A(net3093),
    .X(net3092));
 sg13g2_buf_4 fanout3093 (.X(net3093),
    .A(_02147_));
 sg13g2_buf_8 fanout3094 (.A(net3096),
    .X(net3094));
 sg13g2_buf_4 fanout3095 (.X(net3095),
    .A(net3096));
 sg13g2_buf_8 fanout3096 (.A(_02146_),
    .X(net3096));
 sg13g2_buf_8 fanout3097 (.A(net3100),
    .X(net3097));
 sg13g2_buf_4 fanout3098 (.X(net3098),
    .A(net3100));
 sg13g2_buf_2 fanout3099 (.A(net3100),
    .X(net3099));
 sg13g2_buf_2 fanout3100 (.A(_02146_),
    .X(net3100));
 sg13g2_buf_4 fanout3101 (.X(net3101),
    .A(net3105));
 sg13g2_buf_2 fanout3102 (.A(net3105),
    .X(net3102));
 sg13g2_buf_4 fanout3103 (.X(net3103),
    .A(net3105));
 sg13g2_buf_2 fanout3104 (.A(net3105),
    .X(net3104));
 sg13g2_buf_4 fanout3105 (.X(net3105),
    .A(net3120));
 sg13g2_buf_4 fanout3106 (.X(net3106),
    .A(net3108));
 sg13g2_buf_4 fanout3107 (.X(net3107),
    .A(net3108));
 sg13g2_buf_2 fanout3108 (.A(net3110),
    .X(net3108));
 sg13g2_buf_4 fanout3109 (.X(net3109),
    .A(net3110));
 sg13g2_buf_4 fanout3110 (.X(net3110),
    .A(net3120));
 sg13g2_buf_4 fanout3111 (.X(net3111),
    .A(net3114));
 sg13g2_buf_4 fanout3112 (.X(net3112),
    .A(net3114));
 sg13g2_buf_4 fanout3113 (.X(net3113),
    .A(net3114));
 sg13g2_buf_4 fanout3114 (.X(net3114),
    .A(net3120));
 sg13g2_buf_4 fanout3115 (.X(net3115),
    .A(net3117));
 sg13g2_buf_2 fanout3116 (.A(net3117),
    .X(net3116));
 sg13g2_buf_4 fanout3117 (.X(net3117),
    .A(net3120));
 sg13g2_buf_4 fanout3118 (.X(net3118),
    .A(net3119));
 sg13g2_buf_8 fanout3119 (.A(net3120),
    .X(net3119));
 sg13g2_buf_8 fanout3120 (.A(_02145_),
    .X(net3120));
 sg13g2_buf_2 fanout3121 (.A(net3124),
    .X(net3121));
 sg13g2_buf_2 fanout3122 (.A(net3124),
    .X(net3122));
 sg13g2_buf_4 fanout3123 (.X(net3123),
    .A(net3124));
 sg13g2_buf_2 fanout3124 (.A(net3146),
    .X(net3124));
 sg13g2_buf_4 fanout3125 (.X(net3125),
    .A(net3127));
 sg13g2_buf_2 fanout3126 (.A(net3127),
    .X(net3126));
 sg13g2_buf_4 fanout3127 (.X(net3127),
    .A(net3146));
 sg13g2_buf_4 fanout3128 (.X(net3128),
    .A(net3131));
 sg13g2_buf_4 fanout3129 (.X(net3129),
    .A(net3131));
 sg13g2_buf_2 fanout3130 (.A(net3131),
    .X(net3130));
 sg13g2_buf_2 fanout3131 (.A(net3132),
    .X(net3131));
 sg13g2_buf_2 fanout3132 (.A(net3146),
    .X(net3132));
 sg13g2_buf_4 fanout3133 (.X(net3133),
    .A(net3138));
 sg13g2_buf_4 fanout3134 (.X(net3134),
    .A(net3138));
 sg13g2_buf_2 fanout3135 (.A(net3136),
    .X(net3135));
 sg13g2_buf_2 fanout3136 (.A(net3138),
    .X(net3136));
 sg13g2_buf_2 fanout3137 (.A(net3138),
    .X(net3137));
 sg13g2_buf_4 fanout3138 (.X(net3138),
    .A(net3145));
 sg13g2_buf_4 fanout3139 (.X(net3139),
    .A(net3140));
 sg13g2_buf_4 fanout3140 (.X(net3140),
    .A(net3145));
 sg13g2_buf_2 fanout3141 (.A(net3143),
    .X(net3141));
 sg13g2_buf_2 fanout3142 (.A(net3143),
    .X(net3142));
 sg13g2_buf_2 fanout3143 (.A(net3144),
    .X(net3143));
 sg13g2_buf_4 fanout3144 (.X(net3144),
    .A(net3145));
 sg13g2_buf_2 fanout3145 (.A(net3146),
    .X(net3145));
 sg13g2_buf_4 fanout3146 (.X(net3146),
    .A(_02144_));
 sg13g2_buf_4 fanout3147 (.X(net3147),
    .A(net3148));
 sg13g2_buf_2 fanout3148 (.A(net3149),
    .X(net3148));
 sg13g2_buf_2 fanout3149 (.A(net3174),
    .X(net3149));
 sg13g2_buf_2 fanout3150 (.A(net3153),
    .X(net3150));
 sg13g2_buf_2 fanout3151 (.A(net3153),
    .X(net3151));
 sg13g2_buf_2 fanout3152 (.A(net3153),
    .X(net3152));
 sg13g2_buf_2 fanout3153 (.A(net3174),
    .X(net3153));
 sg13g2_buf_4 fanout3154 (.X(net3154),
    .A(net3159));
 sg13g2_buf_4 fanout3155 (.X(net3155),
    .A(net3157));
 sg13g2_buf_1 fanout3156 (.A(net3157),
    .X(net3156));
 sg13g2_buf_2 fanout3157 (.A(net3159),
    .X(net3157));
 sg13g2_buf_4 fanout3158 (.X(net3158),
    .A(net3159));
 sg13g2_buf_4 fanout3159 (.X(net3159),
    .A(net3174));
 sg13g2_buf_4 fanout3160 (.X(net3160),
    .A(net3165));
 sg13g2_buf_4 fanout3161 (.X(net3161),
    .A(net3164));
 sg13g2_buf_2 fanout3162 (.A(net3163),
    .X(net3162));
 sg13g2_buf_4 fanout3163 (.X(net3163),
    .A(net3164));
 sg13g2_buf_4 fanout3164 (.X(net3164),
    .A(net3165));
 sg13g2_buf_2 fanout3165 (.A(net3174),
    .X(net3165));
 sg13g2_buf_4 fanout3166 (.X(net3166),
    .A(net3169));
 sg13g2_buf_2 fanout3167 (.A(net3168),
    .X(net3167));
 sg13g2_buf_2 fanout3168 (.A(net3169),
    .X(net3168));
 sg13g2_buf_2 fanout3169 (.A(net3173),
    .X(net3169));
 sg13g2_buf_4 fanout3170 (.X(net3170),
    .A(net3172));
 sg13g2_buf_2 fanout3171 (.A(net3172),
    .X(net3171));
 sg13g2_buf_4 fanout3172 (.X(net3172),
    .A(net3173));
 sg13g2_buf_2 fanout3173 (.A(net3174),
    .X(net3173));
 sg13g2_buf_4 fanout3174 (.X(net3174),
    .A(_02144_));
 sg13g2_buf_2 fanout3175 (.A(net3176),
    .X(net3175));
 sg13g2_buf_2 fanout3176 (.A(net3181),
    .X(net3176));
 sg13g2_buf_2 fanout3177 (.A(net3181),
    .X(net3177));
 sg13g2_buf_4 fanout3178 (.X(net3178),
    .A(net3180));
 sg13g2_buf_2 fanout3179 (.A(net3180),
    .X(net3179));
 sg13g2_buf_2 fanout3180 (.A(net3181),
    .X(net3180));
 sg13g2_buf_2 fanout3181 (.A(net3199),
    .X(net3181));
 sg13g2_buf_4 fanout3182 (.X(net3182),
    .A(net3183));
 sg13g2_buf_4 fanout3183 (.X(net3183),
    .A(net3199));
 sg13g2_buf_2 fanout3184 (.A(net3186),
    .X(net3184));
 sg13g2_buf_1 fanout3185 (.A(net3186),
    .X(net3185));
 sg13g2_buf_2 fanout3186 (.A(net3199),
    .X(net3186));
 sg13g2_buf_2 fanout3187 (.A(net3188),
    .X(net3187));
 sg13g2_buf_2 fanout3188 (.A(net3189),
    .X(net3188));
 sg13g2_buf_4 fanout3189 (.X(net3189),
    .A(net3198));
 sg13g2_buf_4 fanout3190 (.X(net3190),
    .A(net3198));
 sg13g2_buf_2 fanout3191 (.A(net3198),
    .X(net3191));
 sg13g2_buf_4 fanout3192 (.X(net3192),
    .A(net3197));
 sg13g2_buf_2 fanout3193 (.A(net3195),
    .X(net3193));
 sg13g2_buf_2 fanout3194 (.A(net3195),
    .X(net3194));
 sg13g2_buf_2 fanout3195 (.A(net3196),
    .X(net3195));
 sg13g2_buf_4 fanout3196 (.X(net3196),
    .A(net3197));
 sg13g2_buf_2 fanout3197 (.A(net3198),
    .X(net3197));
 sg13g2_buf_4 fanout3198 (.X(net3198),
    .A(net3199));
 sg13g2_buf_4 fanout3199 (.X(net3199),
    .A(_02143_));
 sg13g2_buf_2 fanout3200 (.A(net3201),
    .X(net3200));
 sg13g2_buf_2 fanout3201 (.A(net3204),
    .X(net3201));
 sg13g2_buf_2 fanout3202 (.A(net3203),
    .X(net3202));
 sg13g2_buf_2 fanout3203 (.A(net3204),
    .X(net3203));
 sg13g2_buf_2 fanout3204 (.A(net3218),
    .X(net3204));
 sg13g2_buf_2 fanout3205 (.A(net3208),
    .X(net3205));
 sg13g2_buf_2 fanout3206 (.A(net3208),
    .X(net3206));
 sg13g2_buf_2 fanout3207 (.A(net3208),
    .X(net3207));
 sg13g2_buf_2 fanout3208 (.A(net3218),
    .X(net3208));
 sg13g2_buf_4 fanout3209 (.X(net3209),
    .A(net3212));
 sg13g2_buf_4 fanout3210 (.X(net3210),
    .A(net3212));
 sg13g2_buf_2 fanout3211 (.A(net3212),
    .X(net3211));
 sg13g2_buf_2 fanout3212 (.A(net3218),
    .X(net3212));
 sg13g2_buf_2 fanout3213 (.A(net3217),
    .X(net3213));
 sg13g2_buf_2 fanout3214 (.A(net3217),
    .X(net3214));
 sg13g2_buf_2 fanout3215 (.A(net3217),
    .X(net3215));
 sg13g2_buf_1 fanout3216 (.A(net3217),
    .X(net3216));
 sg13g2_buf_2 fanout3217 (.A(net3218),
    .X(net3217));
 sg13g2_buf_4 fanout3218 (.X(net3218),
    .A(_02143_));
 sg13g2_buf_2 fanout3219 (.A(net3221),
    .X(net3219));
 sg13g2_buf_2 fanout3220 (.A(net3221),
    .X(net3220));
 sg13g2_buf_4 fanout3221 (.X(net3221),
    .A(net3237));
 sg13g2_buf_2 fanout3222 (.A(net3223),
    .X(net3222));
 sg13g2_buf_2 fanout3223 (.A(net3227),
    .X(net3223));
 sg13g2_buf_2 fanout3224 (.A(net3226),
    .X(net3224));
 sg13g2_buf_1 fanout3225 (.A(net3226),
    .X(net3225));
 sg13g2_buf_2 fanout3226 (.A(net3227),
    .X(net3226));
 sg13g2_buf_2 fanout3227 (.A(net3237),
    .X(net3227));
 sg13g2_buf_2 fanout3228 (.A(net3231),
    .X(net3228));
 sg13g2_buf_2 fanout3229 (.A(net3231),
    .X(net3229));
 sg13g2_buf_4 fanout3230 (.X(net3230),
    .A(net3231));
 sg13g2_buf_2 fanout3231 (.A(net3237),
    .X(net3231));
 sg13g2_buf_2 fanout3232 (.A(net3233),
    .X(net3232));
 sg13g2_buf_4 fanout3233 (.X(net3233),
    .A(net3237));
 sg13g2_buf_2 fanout3234 (.A(net3236),
    .X(net3234));
 sg13g2_buf_4 fanout3235 (.X(net3235),
    .A(net3236));
 sg13g2_buf_2 fanout3236 (.A(net3237),
    .X(net3236));
 sg13g2_buf_4 fanout3237 (.X(net3237),
    .A(_02143_));
 sg13g2_buf_2 fanout3238 (.A(net3239),
    .X(net3238));
 sg13g2_buf_2 fanout3239 (.A(net3240),
    .X(net3239));
 sg13g2_buf_2 fanout3240 (.A(net3243),
    .X(net3240));
 sg13g2_buf_4 fanout3241 (.X(net3241),
    .A(net3242));
 sg13g2_buf_4 fanout3242 (.X(net3242),
    .A(net3243));
 sg13g2_buf_2 fanout3243 (.A(net3282),
    .X(net3243));
 sg13g2_buf_2 fanout3244 (.A(net3247),
    .X(net3244));
 sg13g2_buf_2 fanout3245 (.A(net3247),
    .X(net3245));
 sg13g2_buf_2 fanout3246 (.A(net3247),
    .X(net3246));
 sg13g2_buf_4 fanout3247 (.X(net3247),
    .A(net3282));
 sg13g2_buf_2 fanout3248 (.A(net3250),
    .X(net3248));
 sg13g2_buf_2 fanout3249 (.A(net3250),
    .X(net3249));
 sg13g2_buf_4 fanout3250 (.X(net3250),
    .A(net3257));
 sg13g2_buf_2 fanout3251 (.A(net3252),
    .X(net3251));
 sg13g2_buf_2 fanout3252 (.A(net3253),
    .X(net3252));
 sg13g2_buf_2 fanout3253 (.A(net3257),
    .X(net3253));
 sg13g2_buf_4 fanout3254 (.X(net3254),
    .A(net3257));
 sg13g2_buf_4 fanout3255 (.X(net3255),
    .A(net3256));
 sg13g2_buf_4 fanout3256 (.X(net3256),
    .A(net3257));
 sg13g2_buf_2 fanout3257 (.A(net3282),
    .X(net3257));
 sg13g2_buf_2 fanout3258 (.A(net3259),
    .X(net3258));
 sg13g2_buf_4 fanout3259 (.X(net3259),
    .A(net3260));
 sg13g2_buf_4 fanout3260 (.X(net3260),
    .A(net3263));
 sg13g2_buf_4 fanout3261 (.X(net3261),
    .A(net3262));
 sg13g2_buf_4 fanout3262 (.X(net3262),
    .A(net3263));
 sg13g2_buf_2 fanout3263 (.A(net3282),
    .X(net3263));
 sg13g2_buf_4 fanout3264 (.X(net3264),
    .A(net3268));
 sg13g2_buf_2 fanout3265 (.A(net3268),
    .X(net3265));
 sg13g2_buf_4 fanout3266 (.X(net3266),
    .A(net3268));
 sg13g2_buf_2 fanout3267 (.A(net3268),
    .X(net3267));
 sg13g2_buf_2 fanout3268 (.A(net3282),
    .X(net3268));
 sg13g2_buf_4 fanout3269 (.X(net3269),
    .A(net3270));
 sg13g2_buf_4 fanout3270 (.X(net3270),
    .A(net3281));
 sg13g2_buf_4 fanout3271 (.X(net3271),
    .A(net3275));
 sg13g2_buf_1 fanout3272 (.A(net3275),
    .X(net3272));
 sg13g2_buf_2 fanout3273 (.A(net3275),
    .X(net3273));
 sg13g2_buf_1 fanout3274 (.A(net3275),
    .X(net3274));
 sg13g2_buf_2 fanout3275 (.A(net3281),
    .X(net3275));
 sg13g2_buf_2 fanout3276 (.A(net3278),
    .X(net3276));
 sg13g2_buf_2 fanout3277 (.A(net3281),
    .X(net3277));
 sg13g2_buf_2 fanout3278 (.A(net3281),
    .X(net3278));
 sg13g2_buf_4 fanout3279 (.X(net3279),
    .A(net3280));
 sg13g2_buf_2 fanout3280 (.A(net3281),
    .X(net3280));
 sg13g2_buf_8 fanout3281 (.A(net3282),
    .X(net3281));
 sg13g2_buf_8 fanout3282 (.A(\mem.data_in[7] ),
    .X(net3282));
 sg13g2_buf_2 fanout3283 (.A(net3287),
    .X(net3283));
 sg13g2_buf_1 fanout3284 (.A(net3287),
    .X(net3284));
 sg13g2_buf_2 fanout3285 (.A(net3287),
    .X(net3285));
 sg13g2_buf_1 fanout3286 (.A(net3287),
    .X(net3286));
 sg13g2_buf_2 fanout3287 (.A(net3289),
    .X(net3287));
 sg13g2_buf_4 fanout3288 (.X(net3288),
    .A(net3289));
 sg13g2_buf_2 fanout3289 (.A(net3308),
    .X(net3289));
 sg13g2_buf_2 fanout3290 (.A(net3293),
    .X(net3290));
 sg13g2_buf_1 fanout3291 (.A(net3293),
    .X(net3291));
 sg13g2_buf_2 fanout3292 (.A(net3293),
    .X(net3292));
 sg13g2_buf_4 fanout3293 (.X(net3293),
    .A(net3308));
 sg13g2_buf_2 fanout3294 (.A(net3296),
    .X(net3294));
 sg13g2_buf_2 fanout3295 (.A(net3296),
    .X(net3295));
 sg13g2_buf_2 fanout3296 (.A(net3308),
    .X(net3296));
 sg13g2_buf_2 fanout3297 (.A(net3302),
    .X(net3297));
 sg13g2_buf_2 fanout3298 (.A(net3299),
    .X(net3298));
 sg13g2_buf_2 fanout3299 (.A(net3301),
    .X(net3299));
 sg13g2_buf_4 fanout3300 (.X(net3300),
    .A(net3301));
 sg13g2_buf_2 fanout3301 (.A(net3302),
    .X(net3301));
 sg13g2_buf_2 fanout3302 (.A(net3308),
    .X(net3302));
 sg13g2_buf_4 fanout3303 (.X(net3303),
    .A(net3307));
 sg13g2_buf_2 fanout3304 (.A(net3307),
    .X(net3304));
 sg13g2_buf_4 fanout3305 (.X(net3305),
    .A(net3307));
 sg13g2_buf_2 fanout3306 (.A(net3307),
    .X(net3306));
 sg13g2_buf_2 fanout3307 (.A(net3308),
    .X(net3307));
 sg13g2_buf_4 fanout3308 (.X(net3308),
    .A(\mem.data_in[6] ));
 sg13g2_buf_4 fanout3309 (.X(net3309),
    .A(net3313));
 sg13g2_buf_4 fanout3310 (.X(net3310),
    .A(net3312));
 sg13g2_buf_2 fanout3311 (.A(net3312),
    .X(net3311));
 sg13g2_buf_2 fanout3312 (.A(net3313),
    .X(net3312));
 sg13g2_buf_2 fanout3313 (.A(net3318),
    .X(net3313));
 sg13g2_buf_2 fanout3314 (.A(net3315),
    .X(net3314));
 sg13g2_buf_2 fanout3315 (.A(net3318),
    .X(net3315));
 sg13g2_buf_2 fanout3316 (.A(net3318),
    .X(net3316));
 sg13g2_buf_4 fanout3317 (.X(net3317),
    .A(net3318));
 sg13g2_buf_4 fanout3318 (.X(net3318),
    .A(\mem.data_in[6] ));
 sg13g2_buf_4 fanout3319 (.X(net3319),
    .A(net3320));
 sg13g2_buf_4 fanout3320 (.X(net3320),
    .A(net3328));
 sg13g2_buf_4 fanout3321 (.X(net3321),
    .A(net3328));
 sg13g2_buf_2 fanout3322 (.A(net3328),
    .X(net3322));
 sg13g2_buf_2 fanout3323 (.A(net3324),
    .X(net3323));
 sg13g2_buf_2 fanout3324 (.A(net3328),
    .X(net3324));
 sg13g2_buf_4 fanout3325 (.X(net3325),
    .A(net3327));
 sg13g2_buf_4 fanout3326 (.X(net3326),
    .A(net3327));
 sg13g2_buf_2 fanout3327 (.A(net3328),
    .X(net3327));
 sg13g2_buf_8 fanout3328 (.A(\mem.data_in[6] ),
    .X(net3328));
 sg13g2_buf_2 fanout3329 (.A(net3335),
    .X(net3329));
 sg13g2_buf_1 fanout3330 (.A(net3335),
    .X(net3330));
 sg13g2_buf_2 fanout3331 (.A(net3335),
    .X(net3331));
 sg13g2_buf_2 fanout3332 (.A(net3334),
    .X(net3332));
 sg13g2_buf_1 fanout3333 (.A(net3334),
    .X(net3333));
 sg13g2_buf_4 fanout3334 (.X(net3334),
    .A(net3335));
 sg13g2_buf_4 fanout3335 (.X(net3335),
    .A(net3341));
 sg13g2_buf_2 fanout3336 (.A(net3338),
    .X(net3336));
 sg13g2_buf_2 fanout3337 (.A(net3338),
    .X(net3337));
 sg13g2_buf_2 fanout3338 (.A(net3341),
    .X(net3338));
 sg13g2_buf_2 fanout3339 (.A(net3341),
    .X(net3339));
 sg13g2_buf_1 fanout3340 (.A(net3341),
    .X(net3340));
 sg13g2_buf_4 fanout3341 (.X(net3341),
    .A(net3352));
 sg13g2_buf_4 fanout3342 (.X(net3342),
    .A(net3343));
 sg13g2_buf_2 fanout3343 (.A(net3352),
    .X(net3343));
 sg13g2_buf_2 fanout3344 (.A(net3346),
    .X(net3344));
 sg13g2_buf_2 fanout3345 (.A(net3346),
    .X(net3345));
 sg13g2_buf_2 fanout3346 (.A(net3352),
    .X(net3346));
 sg13g2_buf_4 fanout3347 (.X(net3347),
    .A(net3348));
 sg13g2_buf_4 fanout3348 (.X(net3348),
    .A(net3351));
 sg13g2_buf_4 fanout3349 (.X(net3349),
    .A(net3351));
 sg13g2_buf_2 fanout3350 (.A(net3351),
    .X(net3350));
 sg13g2_buf_2 fanout3351 (.A(net3352),
    .X(net3351));
 sg13g2_buf_4 fanout3352 (.X(net3352),
    .A(\mem.data_in[5] ));
 sg13g2_buf_4 fanout3353 (.X(net3353),
    .A(net3364));
 sg13g2_buf_2 fanout3354 (.A(net3364),
    .X(net3354));
 sg13g2_buf_2 fanout3355 (.A(net3358),
    .X(net3355));
 sg13g2_buf_2 fanout3356 (.A(net3358),
    .X(net3356));
 sg13g2_buf_2 fanout3357 (.A(net3358),
    .X(net3357));
 sg13g2_buf_2 fanout3358 (.A(net3364),
    .X(net3358));
 sg13g2_buf_4 fanout3359 (.X(net3359),
    .A(net3364));
 sg13g2_buf_2 fanout3360 (.A(net3364),
    .X(net3360));
 sg13g2_buf_4 fanout3361 (.X(net3361),
    .A(net3363));
 sg13g2_buf_1 fanout3362 (.A(net3363),
    .X(net3362));
 sg13g2_buf_2 fanout3363 (.A(net3364),
    .X(net3363));
 sg13g2_buf_8 fanout3364 (.A(\mem.data_in[5] ),
    .X(net3364));
 sg13g2_buf_4 fanout3365 (.X(net3365),
    .A(net3366));
 sg13g2_buf_2 fanout3366 (.A(net3374),
    .X(net3366));
 sg13g2_buf_4 fanout3367 (.X(net3367),
    .A(net3374));
 sg13g2_buf_4 fanout3368 (.X(net3368),
    .A(net3374));
 sg13g2_buf_2 fanout3369 (.A(net3374),
    .X(net3369));
 sg13g2_buf_2 fanout3370 (.A(net3374),
    .X(net3370));
 sg13g2_buf_4 fanout3371 (.X(net3371),
    .A(net3373));
 sg13g2_buf_4 fanout3372 (.X(net3372),
    .A(net3373));
 sg13g2_buf_4 fanout3373 (.X(net3373),
    .A(net3374));
 sg13g2_buf_8 fanout3374 (.A(\mem.data_in[5] ),
    .X(net3374));
 sg13g2_buf_4 fanout3375 (.X(net3375),
    .A(net3386));
 sg13g2_buf_2 fanout3376 (.A(net3386),
    .X(net3376));
 sg13g2_buf_2 fanout3377 (.A(net3379),
    .X(net3377));
 sg13g2_buf_2 fanout3378 (.A(net3379),
    .X(net3378));
 sg13g2_buf_4 fanout3379 (.X(net3379),
    .A(net3386));
 sg13g2_buf_2 fanout3380 (.A(net3383),
    .X(net3380));
 sg13g2_buf_1 fanout3381 (.A(net3383),
    .X(net3381));
 sg13g2_buf_2 fanout3382 (.A(net3383),
    .X(net3382));
 sg13g2_buf_2 fanout3383 (.A(net3385),
    .X(net3383));
 sg13g2_buf_2 fanout3384 (.A(net3385),
    .X(net3384));
 sg13g2_buf_2 fanout3385 (.A(net3386),
    .X(net3385));
 sg13g2_buf_4 fanout3386 (.X(net3386),
    .A(net3421));
 sg13g2_buf_2 fanout3387 (.A(net3388),
    .X(net3387));
 sg13g2_buf_2 fanout3388 (.A(net3389),
    .X(net3388));
 sg13g2_buf_2 fanout3389 (.A(net3390),
    .X(net3389));
 sg13g2_buf_4 fanout3390 (.X(net3390),
    .A(net3396));
 sg13g2_buf_2 fanout3391 (.A(net3396),
    .X(net3391));
 sg13g2_buf_4 fanout3392 (.X(net3392),
    .A(net3394));
 sg13g2_buf_2 fanout3393 (.A(net3394),
    .X(net3393));
 sg13g2_buf_4 fanout3394 (.X(net3394),
    .A(net3395));
 sg13g2_buf_4 fanout3395 (.X(net3395),
    .A(net3396));
 sg13g2_buf_4 fanout3396 (.X(net3396),
    .A(net3421));
 sg13g2_buf_2 fanout3397 (.A(net3399),
    .X(net3397));
 sg13g2_buf_2 fanout3398 (.A(net3399),
    .X(net3398));
 sg13g2_buf_4 fanout3399 (.X(net3399),
    .A(net3402));
 sg13g2_buf_4 fanout3400 (.X(net3400),
    .A(net3401));
 sg13g2_buf_2 fanout3401 (.A(net3402),
    .X(net3401));
 sg13g2_buf_2 fanout3402 (.A(net3421),
    .X(net3402));
 sg13g2_buf_4 fanout3403 (.X(net3403),
    .A(net3407));
 sg13g2_buf_2 fanout3404 (.A(net3407),
    .X(net3404));
 sg13g2_buf_2 fanout3405 (.A(net3407),
    .X(net3405));
 sg13g2_buf_2 fanout3406 (.A(net3407),
    .X(net3406));
 sg13g2_buf_4 fanout3407 (.X(net3407),
    .A(net3421));
 sg13g2_buf_4 fanout3408 (.X(net3408),
    .A(net3420));
 sg13g2_buf_2 fanout3409 (.A(net3420),
    .X(net3409));
 sg13g2_buf_4 fanout3410 (.X(net3410),
    .A(net3412));
 sg13g2_buf_1 fanout3411 (.A(net3412),
    .X(net3411));
 sg13g2_buf_2 fanout3412 (.A(net3420),
    .X(net3412));
 sg13g2_buf_2 fanout3413 (.A(net3415),
    .X(net3413));
 sg13g2_buf_4 fanout3414 (.X(net3414),
    .A(net3415));
 sg13g2_buf_4 fanout3415 (.X(net3415),
    .A(net3420));
 sg13g2_buf_2 fanout3416 (.A(net3419),
    .X(net3416));
 sg13g2_buf_1 fanout3417 (.A(net3419),
    .X(net3417));
 sg13g2_buf_4 fanout3418 (.X(net3418),
    .A(net3419));
 sg13g2_buf_2 fanout3419 (.A(net3420),
    .X(net3419));
 sg13g2_buf_8 fanout3420 (.A(net3421),
    .X(net3420));
 sg13g2_buf_8 fanout3421 (.A(\mem.data_in[4] ),
    .X(net3421));
 sg13g2_buf_2 fanout3422 (.A(net3423),
    .X(net3422));
 sg13g2_buf_2 fanout3423 (.A(net3424),
    .X(net3423));
 sg13g2_buf_2 fanout3424 (.A(net3427),
    .X(net3424));
 sg13g2_buf_4 fanout3425 (.X(net3425),
    .A(net3427));
 sg13g2_buf_2 fanout3426 (.A(net3427),
    .X(net3426));
 sg13g2_buf_2 fanout3427 (.A(net3442),
    .X(net3427));
 sg13g2_buf_2 fanout3428 (.A(net3431),
    .X(net3428));
 sg13g2_buf_2 fanout3429 (.A(net3431),
    .X(net3429));
 sg13g2_buf_2 fanout3430 (.A(net3431),
    .X(net3430));
 sg13g2_buf_4 fanout3431 (.X(net3431),
    .A(net3442));
 sg13g2_buf_2 fanout3432 (.A(net3434),
    .X(net3432));
 sg13g2_buf_1 fanout3433 (.A(net3434),
    .X(net3433));
 sg13g2_buf_2 fanout3434 (.A(net3435),
    .X(net3434));
 sg13g2_buf_4 fanout3435 (.X(net3435),
    .A(net3437));
 sg13g2_buf_4 fanout3436 (.X(net3436),
    .A(net3437));
 sg13g2_buf_2 fanout3437 (.A(net3442),
    .X(net3437));
 sg13g2_buf_4 fanout3438 (.X(net3438),
    .A(net3440));
 sg13g2_buf_2 fanout3439 (.A(net3440),
    .X(net3439));
 sg13g2_buf_4 fanout3440 (.X(net3440),
    .A(net3441));
 sg13g2_buf_2 fanout3441 (.A(net3442),
    .X(net3441));
 sg13g2_buf_4 fanout3442 (.X(net3442),
    .A(net3466));
 sg13g2_buf_4 fanout3443 (.X(net3443),
    .A(net3444));
 sg13g2_buf_4 fanout3444 (.X(net3444),
    .A(net3446));
 sg13g2_buf_4 fanout3445 (.X(net3445),
    .A(net3446));
 sg13g2_buf_2 fanout3446 (.A(net3466),
    .X(net3446));
 sg13g2_buf_2 fanout3447 (.A(net3448),
    .X(net3447));
 sg13g2_buf_2 fanout3448 (.A(net3453),
    .X(net3448));
 sg13g2_buf_4 fanout3449 (.X(net3449),
    .A(net3453));
 sg13g2_buf_2 fanout3450 (.A(net3452),
    .X(net3450));
 sg13g2_buf_4 fanout3451 (.X(net3451),
    .A(net3452));
 sg13g2_buf_2 fanout3452 (.A(net3453),
    .X(net3452));
 sg13g2_buf_2 fanout3453 (.A(net3466),
    .X(net3453));
 sg13g2_buf_4 fanout3454 (.X(net3454),
    .A(net3455));
 sg13g2_buf_4 fanout3455 (.X(net3455),
    .A(net3465));
 sg13g2_buf_4 fanout3456 (.X(net3456),
    .A(net3459));
 sg13g2_buf_1 fanout3457 (.A(net3459),
    .X(net3457));
 sg13g2_buf_4 fanout3458 (.X(net3458),
    .A(net3459));
 sg13g2_buf_2 fanout3459 (.A(net3465),
    .X(net3459));
 sg13g2_buf_2 fanout3460 (.A(net3461),
    .X(net3460));
 sg13g2_buf_4 fanout3461 (.X(net3461),
    .A(net3465));
 sg13g2_buf_4 fanout3462 (.X(net3462),
    .A(net3464));
 sg13g2_buf_4 fanout3463 (.X(net3463),
    .A(net3464));
 sg13g2_buf_2 fanout3464 (.A(net3465),
    .X(net3464));
 sg13g2_buf_4 fanout3465 (.X(net3465),
    .A(net3466));
 sg13g2_buf_8 fanout3466 (.A(\mem.data_in[3] ),
    .X(net3466));
 sg13g2_buf_2 fanout3467 (.A(net3468),
    .X(net3467));
 sg13g2_buf_2 fanout3468 (.A(net3469),
    .X(net3468));
 sg13g2_buf_2 fanout3469 (.A(net3472),
    .X(net3469));
 sg13g2_buf_4 fanout3470 (.X(net3470),
    .A(net3472));
 sg13g2_buf_1 fanout3471 (.A(net3472),
    .X(net3471));
 sg13g2_buf_2 fanout3472 (.A(net3488),
    .X(net3472));
 sg13g2_buf_2 fanout3473 (.A(net3475),
    .X(net3473));
 sg13g2_buf_1 fanout3474 (.A(net3475),
    .X(net3474));
 sg13g2_buf_4 fanout3475 (.X(net3475),
    .A(net3477));
 sg13g2_buf_4 fanout3476 (.X(net3476),
    .A(net3477));
 sg13g2_buf_1 fanout3477 (.A(net3488),
    .X(net3477));
 sg13g2_buf_2 fanout3478 (.A(net3479),
    .X(net3478));
 sg13g2_buf_2 fanout3479 (.A(net3480),
    .X(net3479));
 sg13g2_buf_2 fanout3480 (.A(net3481),
    .X(net3480));
 sg13g2_buf_2 fanout3481 (.A(net3482),
    .X(net3481));
 sg13g2_buf_2 fanout3482 (.A(net3488),
    .X(net3482));
 sg13g2_buf_2 fanout3483 (.A(net3484),
    .X(net3483));
 sg13g2_buf_2 fanout3484 (.A(net3487),
    .X(net3484));
 sg13g2_buf_2 fanout3485 (.A(net3486),
    .X(net3485));
 sg13g2_buf_4 fanout3486 (.X(net3486),
    .A(net3487));
 sg13g2_buf_2 fanout3487 (.A(net3488),
    .X(net3487));
 sg13g2_buf_4 fanout3488 (.X(net3488),
    .A(\mem.data_in[2] ));
 sg13g2_buf_2 fanout3489 (.A(net3491),
    .X(net3489));
 sg13g2_buf_2 fanout3490 (.A(net3491),
    .X(net3490));
 sg13g2_buf_4 fanout3491 (.X(net3491),
    .A(net3494));
 sg13g2_buf_2 fanout3492 (.A(net3493),
    .X(net3492));
 sg13g2_buf_4 fanout3493 (.X(net3493),
    .A(net3494));
 sg13g2_buf_4 fanout3494 (.X(net3494),
    .A(net3512));
 sg13g2_buf_2 fanout3495 (.A(net3496),
    .X(net3495));
 sg13g2_buf_2 fanout3496 (.A(net3497),
    .X(net3496));
 sg13g2_buf_2 fanout3497 (.A(net3512),
    .X(net3497));
 sg13g2_buf_4 fanout3498 (.X(net3498),
    .A(net3512));
 sg13g2_buf_4 fanout3499 (.X(net3499),
    .A(net3501));
 sg13g2_buf_2 fanout3500 (.A(net3501),
    .X(net3500));
 sg13g2_buf_4 fanout3501 (.X(net3501),
    .A(net3511));
 sg13g2_buf_4 fanout3502 (.X(net3502),
    .A(net3503));
 sg13g2_buf_4 fanout3503 (.X(net3503),
    .A(net3511));
 sg13g2_buf_4 fanout3504 (.X(net3504),
    .A(net3505));
 sg13g2_buf_4 fanout3505 (.X(net3505),
    .A(net3511));
 sg13g2_buf_4 fanout3506 (.X(net3506),
    .A(net3510));
 sg13g2_buf_2 fanout3507 (.A(net3510),
    .X(net3507));
 sg13g2_buf_4 fanout3508 (.X(net3508),
    .A(net3510));
 sg13g2_buf_2 fanout3509 (.A(net3510),
    .X(net3509));
 sg13g2_buf_2 fanout3510 (.A(net3511),
    .X(net3510));
 sg13g2_buf_4 fanout3511 (.X(net3511),
    .A(net3512));
 sg13g2_buf_4 fanout3512 (.X(net3512),
    .A(\mem.data_in[2] ));
 sg13g2_buf_4 fanout3513 (.X(net3513),
    .A(net3515));
 sg13g2_buf_2 fanout3514 (.A(net3515),
    .X(net3514));
 sg13g2_buf_2 fanout3515 (.A(net3519),
    .X(net3515));
 sg13g2_buf_2 fanout3516 (.A(net3519),
    .X(net3516));
 sg13g2_buf_2 fanout3517 (.A(net3518),
    .X(net3517));
 sg13g2_buf_2 fanout3518 (.A(net3519),
    .X(net3518));
 sg13g2_buf_2 fanout3519 (.A(net3557),
    .X(net3519));
 sg13g2_buf_2 fanout3520 (.A(net3521),
    .X(net3520));
 sg13g2_buf_1 fanout3521 (.A(net3522),
    .X(net3521));
 sg13g2_buf_4 fanout3522 (.X(net3522),
    .A(net3524));
 sg13g2_buf_4 fanout3523 (.X(net3523),
    .A(net3524));
 sg13g2_buf_2 fanout3524 (.A(net3557),
    .X(net3524));
 sg13g2_buf_4 fanout3525 (.X(net3525),
    .A(net3534));
 sg13g2_buf_4 fanout3526 (.X(net3526),
    .A(net3529));
 sg13g2_buf_2 fanout3527 (.A(net3528),
    .X(net3527));
 sg13g2_buf_4 fanout3528 (.X(net3528),
    .A(net3529));
 sg13g2_buf_2 fanout3529 (.A(net3534),
    .X(net3529));
 sg13g2_buf_2 fanout3530 (.A(net3531),
    .X(net3530));
 sg13g2_buf_4 fanout3531 (.X(net3531),
    .A(net3533));
 sg13g2_buf_4 fanout3532 (.X(net3532),
    .A(net3533));
 sg13g2_buf_4 fanout3533 (.X(net3533),
    .A(net3534));
 sg13g2_buf_2 fanout3534 (.A(net3557),
    .X(net3534));
 sg13g2_buf_4 fanout3535 (.X(net3535),
    .A(net3539));
 sg13g2_buf_4 fanout3536 (.X(net3536),
    .A(net3538));
 sg13g2_buf_2 fanout3537 (.A(net3538),
    .X(net3537));
 sg13g2_buf_4 fanout3538 (.X(net3538),
    .A(net3539));
 sg13g2_buf_2 fanout3539 (.A(net3556),
    .X(net3539));
 sg13g2_buf_4 fanout3540 (.X(net3540),
    .A(net3544));
 sg13g2_buf_2 fanout3541 (.A(net3544),
    .X(net3541));
 sg13g2_buf_4 fanout3542 (.X(net3542),
    .A(net3544));
 sg13g2_buf_2 fanout3543 (.A(net3544),
    .X(net3543));
 sg13g2_buf_2 fanout3544 (.A(net3556),
    .X(net3544));
 sg13g2_buf_4 fanout3545 (.X(net3545),
    .A(net3547));
 sg13g2_buf_1 fanout3546 (.A(net3547),
    .X(net3546));
 sg13g2_buf_4 fanout3547 (.X(net3547),
    .A(net3550));
 sg13g2_buf_4 fanout3548 (.X(net3548),
    .A(net3550));
 sg13g2_buf_4 fanout3549 (.X(net3549),
    .A(net3550));
 sg13g2_buf_4 fanout3550 (.X(net3550),
    .A(net3556));
 sg13g2_buf_2 fanout3551 (.A(net3555),
    .X(net3551));
 sg13g2_buf_4 fanout3552 (.X(net3552),
    .A(net3555));
 sg13g2_buf_2 fanout3553 (.A(net3554),
    .X(net3553));
 sg13g2_buf_2 fanout3554 (.A(net3555),
    .X(net3554));
 sg13g2_buf_4 fanout3555 (.X(net3555),
    .A(net3556));
 sg13g2_buf_8 fanout3556 (.A(net3557),
    .X(net3556));
 sg13g2_buf_4 fanout3557 (.X(net3557),
    .A(\mem.data_in[1] ));
 sg13g2_buf_2 fanout3558 (.A(net3560),
    .X(net3558));
 sg13g2_buf_1 fanout3559 (.A(net3560),
    .X(net3559));
 sg13g2_buf_2 fanout3560 (.A(net3561),
    .X(net3560));
 sg13g2_buf_2 fanout3561 (.A(net3564),
    .X(net3561));
 sg13g2_buf_4 fanout3562 (.X(net3562),
    .A(net3564));
 sg13g2_buf_1 fanout3563 (.A(net3564),
    .X(net3563));
 sg13g2_buf_4 fanout3564 (.X(net3564),
    .A(net3571));
 sg13g2_buf_2 fanout3565 (.A(net3567),
    .X(net3565));
 sg13g2_buf_2 fanout3566 (.A(net3567),
    .X(net3566));
 sg13g2_buf_2 fanout3567 (.A(net3570),
    .X(net3567));
 sg13g2_buf_2 fanout3568 (.A(net3569),
    .X(net3568));
 sg13g2_buf_2 fanout3569 (.A(net3570),
    .X(net3569));
 sg13g2_buf_4 fanout3570 (.X(net3570),
    .A(net3571));
 sg13g2_buf_2 fanout3571 (.A(net3602),
    .X(net3571));
 sg13g2_buf_2 fanout3572 (.A(net3574),
    .X(net3572));
 sg13g2_buf_1 fanout3573 (.A(net3574),
    .X(net3573));
 sg13g2_buf_4 fanout3574 (.X(net3574),
    .A(net3577));
 sg13g2_buf_2 fanout3575 (.A(net3576),
    .X(net3575));
 sg13g2_buf_4 fanout3576 (.X(net3576),
    .A(net3577));
 sg13g2_buf_2 fanout3577 (.A(net3602),
    .X(net3577));
 sg13g2_buf_4 fanout3578 (.X(net3578),
    .A(net3581));
 sg13g2_buf_4 fanout3579 (.X(net3579),
    .A(net3581));
 sg13g2_buf_2 fanout3580 (.A(net3581),
    .X(net3580));
 sg13g2_buf_2 fanout3581 (.A(net3602),
    .X(net3581));
 sg13g2_buf_4 fanout3582 (.X(net3582),
    .A(net3583));
 sg13g2_buf_4 fanout3583 (.X(net3583),
    .A(net3589));
 sg13g2_buf_2 fanout3584 (.A(net3588),
    .X(net3584));
 sg13g2_buf_2 fanout3585 (.A(net3588),
    .X(net3585));
 sg13g2_buf_2 fanout3586 (.A(net3587),
    .X(net3586));
 sg13g2_buf_4 fanout3587 (.X(net3587),
    .A(net3588));
 sg13g2_buf_4 fanout3588 (.X(net3588),
    .A(net3589));
 sg13g2_buf_2 fanout3589 (.A(net3602),
    .X(net3589));
 sg13g2_buf_4 fanout3590 (.X(net3590),
    .A(net3591));
 sg13g2_buf_4 fanout3591 (.X(net3591),
    .A(net3601));
 sg13g2_buf_2 fanout3592 (.A(net3594),
    .X(net3592));
 sg13g2_buf_4 fanout3593 (.X(net3593),
    .A(net3594));
 sg13g2_buf_2 fanout3594 (.A(net3595),
    .X(net3594));
 sg13g2_buf_2 fanout3595 (.A(net3601),
    .X(net3595));
 sg13g2_buf_2 fanout3596 (.A(net3597),
    .X(net3596));
 sg13g2_buf_4 fanout3597 (.X(net3597),
    .A(net3600));
 sg13g2_buf_2 fanout3598 (.A(net3600),
    .X(net3598));
 sg13g2_buf_2 fanout3599 (.A(net3600),
    .X(net3599));
 sg13g2_buf_2 fanout3600 (.A(net3601),
    .X(net3600));
 sg13g2_buf_4 fanout3601 (.X(net3601),
    .A(net3602));
 sg13g2_buf_8 fanout3602 (.A(\mem.data_in[0] ),
    .X(net3602));
 sg13g2_buf_4 fanout3603 (.X(net3603),
    .A(\mem.addr[6] ));
 sg13g2_buf_4 fanout3604 (.X(net3604),
    .A(\mem.addr[4] ));
 sg13g2_buf_4 fanout3605 (.X(net3605),
    .A(\mem.addr[3] ));
 sg13g2_buf_4 fanout3606 (.X(net3606),
    .A(net5222));
 sg13g2_buf_4 fanout3607 (.X(net3607),
    .A(net5218));
 sg13g2_buf_4 fanout3608 (.X(net3608),
    .A(\mem.addr[0] ));
 sg13g2_buf_4 fanout3609 (.X(net3609),
    .A(\state[1] ));
 sg13g2_buf_2 fanout3610 (.A(\state[0] ),
    .X(net3610));
 sg13g2_buf_2 fanout3611 (.A(_00007_),
    .X(net3611));
 sg13g2_buf_4 fanout3612 (.X(net3612),
    .A(net3613));
 sg13g2_buf_2 fanout3613 (.A(net3614),
    .X(net3613));
 sg13g2_buf_8 fanout3614 (.A(_00006_),
    .X(net3614));
 sg13g2_buf_8 fanout3615 (.A(net3619),
    .X(net3615));
 sg13g2_buf_2 fanout3616 (.A(net3617),
    .X(net3616));
 sg13g2_buf_4 fanout3617 (.X(net3617),
    .A(net3619));
 sg13g2_buf_8 fanout3618 (.A(net3619),
    .X(net3618));
 sg13g2_buf_8 fanout3619 (.A(_00005_),
    .X(net3619));
 sg13g2_buf_4 fanout3620 (.X(net3620),
    .A(net3621));
 sg13g2_buf_8 fanout3621 (.A(net3624),
    .X(net3621));
 sg13g2_buf_4 fanout3622 (.X(net3622),
    .A(net3623));
 sg13g2_buf_8 fanout3623 (.A(net3624),
    .X(net3623));
 sg13g2_buf_8 fanout3624 (.A(_00004_),
    .X(net3624));
 sg13g2_buf_8 fanout3625 (.A(net3631),
    .X(net3625));
 sg13g2_buf_8 fanout3626 (.A(net3628),
    .X(net3626));
 sg13g2_buf_2 fanout3627 (.A(net3628),
    .X(net3627));
 sg13g2_buf_4 fanout3628 (.X(net3628),
    .A(net3631));
 sg13g2_buf_4 fanout3629 (.X(net3629),
    .A(net3631));
 sg13g2_buf_4 fanout3630 (.X(net3630),
    .A(net3631));
 sg13g2_buf_8 fanout3631 (.A(_00004_),
    .X(net3631));
 sg13g2_buf_4 fanout3632 (.X(net3632),
    .A(net3633));
 sg13g2_buf_4 fanout3633 (.X(net3633),
    .A(net3637));
 sg13g2_buf_4 fanout3634 (.X(net3634),
    .A(net3635));
 sg13g2_buf_4 fanout3635 (.X(net3635),
    .A(net3637));
 sg13g2_buf_2 fanout3636 (.A(net3637),
    .X(net3636));
 sg13g2_buf_4 fanout3637 (.X(net3637),
    .A(net3642));
 sg13g2_buf_4 fanout3638 (.X(net3638),
    .A(net3642));
 sg13g2_buf_4 fanout3639 (.X(net3639),
    .A(net3642));
 sg13g2_buf_4 fanout3640 (.X(net3640),
    .A(net3641));
 sg13g2_buf_4 fanout3641 (.X(net3641),
    .A(net3642));
 sg13g2_buf_2 fanout3642 (.A(_00003_),
    .X(net3642));
 sg13g2_buf_4 fanout3643 (.X(net3643),
    .A(net3645));
 sg13g2_buf_4 fanout3644 (.X(net3644),
    .A(net3645));
 sg13g2_buf_2 fanout3645 (.A(net3656),
    .X(net3645));
 sg13g2_buf_4 fanout3646 (.X(net3646),
    .A(net3656));
 sg13g2_buf_4 fanout3647 (.X(net3647),
    .A(net3656));
 sg13g2_buf_4 fanout3648 (.X(net3648),
    .A(net3655));
 sg13g2_buf_2 fanout3649 (.A(net3655),
    .X(net3649));
 sg13g2_buf_4 fanout3650 (.X(net3650),
    .A(net3655));
 sg13g2_buf_4 fanout3651 (.X(net3651),
    .A(net3652));
 sg13g2_buf_4 fanout3652 (.X(net3652),
    .A(net3654));
 sg13g2_buf_4 fanout3653 (.X(net3653),
    .A(net3654));
 sg13g2_buf_2 fanout3654 (.A(net3655),
    .X(net3654));
 sg13g2_buf_4 fanout3655 (.X(net3655),
    .A(net3656));
 sg13g2_buf_4 fanout3656 (.X(net3656),
    .A(_00003_));
 sg13g2_buf_4 fanout3657 (.X(net3657),
    .A(net3666));
 sg13g2_buf_2 fanout3658 (.A(net3666),
    .X(net3658));
 sg13g2_buf_2 fanout3659 (.A(net3660),
    .X(net3659));
 sg13g2_buf_4 fanout3660 (.X(net3660),
    .A(net3666));
 sg13g2_buf_2 fanout3661 (.A(net3662),
    .X(net3661));
 sg13g2_buf_2 fanout3662 (.A(net3663),
    .X(net3662));
 sg13g2_buf_4 fanout3663 (.X(net3663),
    .A(net3665));
 sg13g2_buf_4 fanout3664 (.X(net3664),
    .A(net3665));
 sg13g2_buf_2 fanout3665 (.A(net3666),
    .X(net3665));
 sg13g2_buf_4 fanout3666 (.X(net3666),
    .A(net3673));
 sg13g2_buf_4 fanout3667 (.X(net3667),
    .A(net3670));
 sg13g2_buf_4 fanout3668 (.X(net3668),
    .A(net3669));
 sg13g2_buf_4 fanout3669 (.X(net3669),
    .A(net3670));
 sg13g2_buf_4 fanout3670 (.X(net3670),
    .A(net3673));
 sg13g2_buf_4 fanout3671 (.X(net3671),
    .A(net3673));
 sg13g2_buf_2 fanout3672 (.A(net3673),
    .X(net3672));
 sg13g2_buf_4 fanout3673 (.X(net3673),
    .A(_00002_));
 sg13g2_buf_2 fanout3674 (.A(net3675),
    .X(net3674));
 sg13g2_buf_4 fanout3675 (.X(net3675),
    .A(net3676));
 sg13g2_buf_4 fanout3676 (.X(net3676),
    .A(net3681));
 sg13g2_buf_4 fanout3677 (.X(net3677),
    .A(net3680));
 sg13g2_buf_2 fanout3678 (.A(net3680),
    .X(net3678));
 sg13g2_buf_4 fanout3679 (.X(net3679),
    .A(net3680));
 sg13g2_buf_2 fanout3680 (.A(net3681),
    .X(net3680));
 sg13g2_buf_4 fanout3681 (.X(net3681),
    .A(_00002_));
 sg13g2_buf_4 fanout3682 (.X(net3682),
    .A(net3685));
 sg13g2_buf_4 fanout3683 (.X(net3683),
    .A(net3684));
 sg13g2_buf_4 fanout3684 (.X(net3684),
    .A(net3685));
 sg13g2_buf_2 fanout3685 (.A(net3690),
    .X(net3685));
 sg13g2_buf_4 fanout3686 (.X(net3686),
    .A(net3690));
 sg13g2_buf_2 fanout3687 (.A(net3690),
    .X(net3687));
 sg13g2_buf_4 fanout3688 (.X(net3688),
    .A(net3689));
 sg13g2_buf_4 fanout3689 (.X(net3689),
    .A(net3690));
 sg13g2_buf_4 fanout3690 (.X(net3690),
    .A(_00002_));
 sg13g2_buf_4 fanout3691 (.X(net3691),
    .A(net3692));
 sg13g2_buf_4 fanout3692 (.X(net3692),
    .A(net3701));
 sg13g2_buf_4 fanout3693 (.X(net3693),
    .A(net3695));
 sg13g2_buf_2 fanout3694 (.A(net3695),
    .X(net3694));
 sg13g2_buf_4 fanout3695 (.X(net3695),
    .A(net3701));
 sg13g2_buf_4 fanout3696 (.X(net3696),
    .A(net3700));
 sg13g2_buf_4 fanout3697 (.X(net3697),
    .A(net3700));
 sg13g2_buf_4 fanout3698 (.X(net3698),
    .A(net3700));
 sg13g2_buf_2 fanout3699 (.A(net3700),
    .X(net3699));
 sg13g2_buf_2 fanout3700 (.A(net3701),
    .X(net3700));
 sg13g2_buf_2 fanout3701 (.A(net3731),
    .X(net3701));
 sg13g2_buf_4 fanout3702 (.X(net3702),
    .A(net3704));
 sg13g2_buf_1 fanout3703 (.A(net3704),
    .X(net3703));
 sg13g2_buf_4 fanout3704 (.X(net3704),
    .A(net3711));
 sg13g2_buf_4 fanout3705 (.X(net3705),
    .A(net3707));
 sg13g2_buf_2 fanout3706 (.A(net3707),
    .X(net3706));
 sg13g2_buf_4 fanout3707 (.X(net3707),
    .A(net3711));
 sg13g2_buf_4 fanout3708 (.X(net3708),
    .A(net3710));
 sg13g2_buf_2 fanout3709 (.A(net3710),
    .X(net3709));
 sg13g2_buf_2 fanout3710 (.A(net3711),
    .X(net3710));
 sg13g2_buf_2 fanout3711 (.A(net3731),
    .X(net3711));
 sg13g2_buf_4 fanout3712 (.X(net3712),
    .A(net3713));
 sg13g2_buf_4 fanout3713 (.X(net3713),
    .A(net3720));
 sg13g2_buf_4 fanout3714 (.X(net3714),
    .A(net3720));
 sg13g2_buf_4 fanout3715 (.X(net3715),
    .A(net3717));
 sg13g2_buf_4 fanout3716 (.X(net3716),
    .A(net3717));
 sg13g2_buf_2 fanout3717 (.A(net3720),
    .X(net3717));
 sg13g2_buf_4 fanout3718 (.X(net3718),
    .A(net3719));
 sg13g2_buf_4 fanout3719 (.X(net3719),
    .A(net3720));
 sg13g2_buf_2 fanout3720 (.A(net3731),
    .X(net3720));
 sg13g2_buf_4 fanout3721 (.X(net3721),
    .A(net3730));
 sg13g2_buf_2 fanout3722 (.A(net3730),
    .X(net3722));
 sg13g2_buf_2 fanout3723 (.A(net3724),
    .X(net3723));
 sg13g2_buf_2 fanout3724 (.A(net3730),
    .X(net3724));
 sg13g2_buf_4 fanout3725 (.X(net3725),
    .A(net3729));
 sg13g2_buf_4 fanout3726 (.X(net3726),
    .A(net3729));
 sg13g2_buf_2 fanout3727 (.A(net3728),
    .X(net3727));
 sg13g2_buf_4 fanout3728 (.X(net3728),
    .A(net3729));
 sg13g2_buf_2 fanout3729 (.A(net3730),
    .X(net3729));
 sg13g2_buf_2 fanout3730 (.A(net3731),
    .X(net3730));
 sg13g2_buf_4 fanout3731 (.X(net3731),
    .A(_00001_));
 sg13g2_buf_4 fanout3732 (.X(net3732),
    .A(net3733));
 sg13g2_buf_4 fanout3733 (.X(net3733),
    .A(net3736));
 sg13g2_buf_4 fanout3734 (.X(net3734),
    .A(net3736));
 sg13g2_buf_2 fanout3735 (.A(net3736),
    .X(net3735));
 sg13g2_buf_2 fanout3736 (.A(net3741),
    .X(net3736));
 sg13g2_buf_4 fanout3737 (.X(net3737),
    .A(net3738));
 sg13g2_buf_4 fanout3738 (.X(net3738),
    .A(net3741));
 sg13g2_buf_4 fanout3739 (.X(net3739),
    .A(net3740));
 sg13g2_buf_4 fanout3740 (.X(net3740),
    .A(net3741));
 sg13g2_buf_2 fanout3741 (.A(net3770),
    .X(net3741));
 sg13g2_buf_4 fanout3742 (.X(net3742),
    .A(net3745));
 sg13g2_buf_2 fanout3743 (.A(net3744),
    .X(net3743));
 sg13g2_buf_4 fanout3744 (.X(net3744),
    .A(net3745));
 sg13g2_buf_2 fanout3745 (.A(net3770),
    .X(net3745));
 sg13g2_buf_4 fanout3746 (.X(net3746),
    .A(net3747));
 sg13g2_buf_2 fanout3747 (.A(net3750),
    .X(net3747));
 sg13g2_buf_4 fanout3748 (.X(net3748),
    .A(net3749));
 sg13g2_buf_4 fanout3749 (.X(net3749),
    .A(net3750));
 sg13g2_buf_2 fanout3750 (.A(net3770),
    .X(net3750));
 sg13g2_buf_4 fanout3751 (.X(net3751),
    .A(net3752));
 sg13g2_buf_4 fanout3752 (.X(net3752),
    .A(net3754));
 sg13g2_buf_4 fanout3753 (.X(net3753),
    .A(net3754));
 sg13g2_buf_2 fanout3754 (.A(net3770),
    .X(net3754));
 sg13g2_buf_4 fanout3755 (.X(net3755),
    .A(net3759));
 sg13g2_buf_4 fanout3756 (.X(net3756),
    .A(net3759));
 sg13g2_buf_4 fanout3757 (.X(net3757),
    .A(net3759));
 sg13g2_buf_4 fanout3758 (.X(net3758),
    .A(net3759));
 sg13g2_buf_2 fanout3759 (.A(net3770),
    .X(net3759));
 sg13g2_buf_4 fanout3760 (.X(net3760),
    .A(net3764));
 sg13g2_buf_2 fanout3761 (.A(net3764),
    .X(net3761));
 sg13g2_buf_4 fanout3762 (.X(net3762),
    .A(net3763));
 sg13g2_buf_4 fanout3763 (.X(net3763),
    .A(net3764));
 sg13g2_buf_2 fanout3764 (.A(net3769),
    .X(net3764));
 sg13g2_buf_4 fanout3765 (.X(net3765),
    .A(net3766));
 sg13g2_buf_4 fanout3766 (.X(net3766),
    .A(net3769));
 sg13g2_buf_4 fanout3767 (.X(net3767),
    .A(net3768));
 sg13g2_buf_4 fanout3768 (.X(net3768),
    .A(net3769));
 sg13g2_buf_2 fanout3769 (.A(net3770),
    .X(net3769));
 sg13g2_buf_8 fanout3770 (.A(_00001_),
    .X(net3770));
 sg13g2_buf_4 fanout3771 (.X(net3771),
    .A(net3773));
 sg13g2_buf_4 fanout3772 (.X(net3772),
    .A(net3773));
 sg13g2_buf_2 fanout3773 (.A(net3782),
    .X(net3773));
 sg13g2_buf_4 fanout3774 (.X(net3774),
    .A(net3776));
 sg13g2_buf_2 fanout3775 (.A(net3776),
    .X(net3775));
 sg13g2_buf_2 fanout3776 (.A(net3782),
    .X(net3776));
 sg13g2_buf_4 fanout3777 (.X(net3777),
    .A(net3778));
 sg13g2_buf_4 fanout3778 (.X(net3778),
    .A(net3781));
 sg13g2_buf_2 fanout3779 (.A(net3780),
    .X(net3779));
 sg13g2_buf_4 fanout3780 (.X(net3780),
    .A(net3781));
 sg13g2_buf_4 fanout3781 (.X(net3781),
    .A(net3782));
 sg13g2_buf_2 fanout3782 (.A(net3796),
    .X(net3782));
 sg13g2_buf_2 fanout3783 (.A(net3786),
    .X(net3783));
 sg13g2_buf_2 fanout3784 (.A(net3786),
    .X(net3784));
 sg13g2_buf_2 fanout3785 (.A(net3786),
    .X(net3785));
 sg13g2_buf_2 fanout3786 (.A(net3789),
    .X(net3786));
 sg13g2_buf_2 fanout3787 (.A(net3788),
    .X(net3787));
 sg13g2_buf_8 fanout3788 (.A(net3789),
    .X(net3788));
 sg13g2_buf_2 fanout3789 (.A(net3796),
    .X(net3789));
 sg13g2_buf_4 fanout3790 (.X(net3790),
    .A(net3792));
 sg13g2_buf_4 fanout3791 (.X(net3791),
    .A(net3792));
 sg13g2_buf_2 fanout3792 (.A(net3796),
    .X(net3792));
 sg13g2_buf_4 fanout3793 (.X(net3793),
    .A(net3794));
 sg13g2_buf_2 fanout3794 (.A(net3795),
    .X(net3794));
 sg13g2_buf_2 fanout3795 (.A(net3796),
    .X(net3795));
 sg13g2_buf_4 fanout3796 (.X(net3796),
    .A(net3815));
 sg13g2_buf_4 fanout3797 (.X(net3797),
    .A(net3799));
 sg13g2_buf_4 fanout3798 (.X(net3798),
    .A(net3799));
 sg13g2_buf_2 fanout3799 (.A(net3807),
    .X(net3799));
 sg13g2_buf_4 fanout3800 (.X(net3800),
    .A(net3807));
 sg13g2_buf_1 fanout3801 (.A(net3807),
    .X(net3801));
 sg13g2_buf_4 fanout3802 (.X(net3802),
    .A(net3803));
 sg13g2_buf_8 fanout3803 (.A(net3806),
    .X(net3803));
 sg13g2_buf_4 fanout3804 (.X(net3804),
    .A(net3806));
 sg13g2_buf_2 fanout3805 (.A(net3806),
    .X(net3805));
 sg13g2_buf_2 fanout3806 (.A(net3807),
    .X(net3806));
 sg13g2_buf_2 fanout3807 (.A(net3815),
    .X(net3807));
 sg13g2_buf_4 fanout3808 (.X(net3808),
    .A(net3811));
 sg13g2_buf_2 fanout3809 (.A(net3811),
    .X(net3809));
 sg13g2_buf_1 fanout3810 (.A(net3811),
    .X(net3810));
 sg13g2_buf_2 fanout3811 (.A(net3814),
    .X(net3811));
 sg13g2_buf_4 fanout3812 (.X(net3812),
    .A(net3814));
 sg13g2_buf_2 fanout3813 (.A(net3814),
    .X(net3813));
 sg13g2_buf_4 fanout3814 (.X(net3814),
    .A(net3815));
 sg13g2_buf_4 fanout3815 (.X(net3815),
    .A(net3992));
 sg13g2_buf_2 fanout3816 (.A(net3818),
    .X(net3816));
 sg13g2_buf_2 fanout3817 (.A(net3818),
    .X(net3817));
 sg13g2_buf_4 fanout3818 (.X(net3818),
    .A(net3819));
 sg13g2_buf_8 fanout3819 (.A(net3840),
    .X(net3819));
 sg13g2_buf_4 fanout3820 (.X(net3820),
    .A(net3823));
 sg13g2_buf_2 fanout3821 (.A(net3822),
    .X(net3821));
 sg13g2_buf_2 fanout3822 (.A(net3823),
    .X(net3822));
 sg13g2_buf_2 fanout3823 (.A(net3826),
    .X(net3823));
 sg13g2_buf_2 fanout3824 (.A(net3825),
    .X(net3824));
 sg13g2_buf_4 fanout3825 (.X(net3825),
    .A(net3826));
 sg13g2_buf_1 fanout3826 (.A(net3840),
    .X(net3826));
 sg13g2_buf_2 fanout3827 (.A(net3828),
    .X(net3827));
 sg13g2_buf_4 fanout3828 (.X(net3828),
    .A(net3829));
 sg13g2_buf_2 fanout3829 (.A(net3839),
    .X(net3829));
 sg13g2_buf_2 fanout3830 (.A(net3832),
    .X(net3830));
 sg13g2_buf_2 fanout3831 (.A(net3832),
    .X(net3831));
 sg13g2_buf_4 fanout3832 (.X(net3832),
    .A(net3839));
 sg13g2_buf_4 fanout3833 (.X(net3833),
    .A(net3834));
 sg13g2_buf_4 fanout3834 (.X(net3834),
    .A(net3839));
 sg13g2_buf_2 fanout3835 (.A(net3837),
    .X(net3835));
 sg13g2_buf_2 fanout3836 (.A(net3837),
    .X(net3836));
 sg13g2_buf_2 fanout3837 (.A(net3838),
    .X(net3837));
 sg13g2_buf_2 fanout3838 (.A(net3839),
    .X(net3838));
 sg13g2_buf_2 fanout3839 (.A(net3840),
    .X(net3839));
 sg13g2_buf_4 fanout3840 (.X(net3840),
    .A(net3992));
 sg13g2_buf_4 fanout3841 (.X(net3841),
    .A(net3845));
 sg13g2_buf_4 fanout3842 (.X(net3842),
    .A(net3844));
 sg13g2_buf_1 fanout3843 (.A(net3844),
    .X(net3843));
 sg13g2_buf_2 fanout3844 (.A(net3845),
    .X(net3844));
 sg13g2_buf_2 fanout3845 (.A(net3863),
    .X(net3845));
 sg13g2_buf_2 fanout3846 (.A(net3847),
    .X(net3846));
 sg13g2_buf_2 fanout3847 (.A(net3848),
    .X(net3847));
 sg13g2_buf_4 fanout3848 (.X(net3848),
    .A(net3863));
 sg13g2_buf_4 fanout3849 (.X(net3849),
    .A(net3853));
 sg13g2_buf_2 fanout3850 (.A(net3853),
    .X(net3850));
 sg13g2_buf_4 fanout3851 (.X(net3851),
    .A(net3852));
 sg13g2_buf_4 fanout3852 (.X(net3852),
    .A(net3853));
 sg13g2_buf_2 fanout3853 (.A(net3863),
    .X(net3853));
 sg13g2_buf_2 fanout3854 (.A(net3857),
    .X(net3854));
 sg13g2_buf_1 fanout3855 (.A(net3856),
    .X(net3855));
 sg13g2_buf_2 fanout3856 (.A(net3857),
    .X(net3856));
 sg13g2_buf_4 fanout3857 (.X(net3857),
    .A(net3862));
 sg13g2_buf_2 fanout3858 (.A(net3859),
    .X(net3858));
 sg13g2_buf_2 fanout3859 (.A(net3862),
    .X(net3859));
 sg13g2_buf_4 fanout3860 (.X(net3860),
    .A(net3862));
 sg13g2_buf_2 fanout3861 (.A(net3862),
    .X(net3861));
 sg13g2_buf_2 fanout3862 (.A(net3863),
    .X(net3862));
 sg13g2_buf_2 fanout3863 (.A(net3992),
    .X(net3863));
 sg13g2_buf_2 fanout3864 (.A(net3866),
    .X(net3864));
 sg13g2_buf_2 fanout3865 (.A(net3866),
    .X(net3865));
 sg13g2_buf_4 fanout3866 (.X(net3866),
    .A(net3871));
 sg13g2_buf_4 fanout3867 (.X(net3867),
    .A(net3870));
 sg13g2_buf_2 fanout3868 (.A(net3870),
    .X(net3868));
 sg13g2_buf_2 fanout3869 (.A(net3870),
    .X(net3869));
 sg13g2_buf_2 fanout3870 (.A(net3871),
    .X(net3870));
 sg13g2_buf_2 fanout3871 (.A(net3893),
    .X(net3871));
 sg13g2_buf_2 fanout3872 (.A(net3874),
    .X(net3872));
 sg13g2_buf_2 fanout3873 (.A(net3874),
    .X(net3873));
 sg13g2_buf_4 fanout3874 (.X(net3874),
    .A(net3878));
 sg13g2_buf_2 fanout3875 (.A(net3878),
    .X(net3875));
 sg13g2_buf_2 fanout3876 (.A(net3878),
    .X(net3876));
 sg13g2_buf_4 fanout3877 (.X(net3877),
    .A(net3878));
 sg13g2_buf_2 fanout3878 (.A(net3893),
    .X(net3878));
 sg13g2_buf_4 fanout3879 (.X(net3879),
    .A(net3882));
 sg13g2_buf_4 fanout3880 (.X(net3880),
    .A(net3882));
 sg13g2_buf_1 fanout3881 (.A(net3882),
    .X(net3881));
 sg13g2_buf_2 fanout3882 (.A(net3885),
    .X(net3882));
 sg13g2_buf_4 fanout3883 (.X(net3883),
    .A(net3885));
 sg13g2_buf_4 fanout3884 (.X(net3884),
    .A(net3885));
 sg13g2_buf_2 fanout3885 (.A(net3893),
    .X(net3885));
 sg13g2_buf_4 fanout3886 (.X(net3886),
    .A(net3887));
 sg13g2_buf_4 fanout3887 (.X(net3887),
    .A(net3892));
 sg13g2_buf_2 fanout3888 (.A(net3892),
    .X(net3888));
 sg13g2_buf_1 fanout3889 (.A(net3892),
    .X(net3889));
 sg13g2_buf_2 fanout3890 (.A(net3891),
    .X(net3890));
 sg13g2_buf_2 fanout3891 (.A(net3892),
    .X(net3891));
 sg13g2_buf_2 fanout3892 (.A(net3893),
    .X(net3892));
 sg13g2_buf_4 fanout3893 (.X(net3893),
    .A(net3992));
 sg13g2_buf_2 fanout3894 (.A(net3896),
    .X(net3894));
 sg13g2_buf_2 fanout3895 (.A(net3896),
    .X(net3895));
 sg13g2_buf_4 fanout3896 (.X(net3896),
    .A(net3899));
 sg13g2_buf_2 fanout3897 (.A(net3898),
    .X(net3897));
 sg13g2_buf_4 fanout3898 (.X(net3898),
    .A(net3899));
 sg13g2_buf_2 fanout3899 (.A(net3924),
    .X(net3899));
 sg13g2_buf_4 fanout3900 (.X(net3900),
    .A(net3902));
 sg13g2_buf_2 fanout3901 (.A(net3902),
    .X(net3901));
 sg13g2_buf_4 fanout3902 (.X(net3902),
    .A(net3924));
 sg13g2_buf_2 fanout3903 (.A(net3906),
    .X(net3903));
 sg13g2_buf_2 fanout3904 (.A(net3906),
    .X(net3904));
 sg13g2_buf_2 fanout3905 (.A(net3906),
    .X(net3905));
 sg13g2_buf_2 fanout3906 (.A(net3924),
    .X(net3906));
 sg13g2_buf_2 fanout3907 (.A(net3908),
    .X(net3907));
 sg13g2_buf_1 fanout3908 (.A(net3909),
    .X(net3908));
 sg13g2_buf_2 fanout3909 (.A(net3910),
    .X(net3909));
 sg13g2_buf_4 fanout3910 (.X(net3910),
    .A(net3923));
 sg13g2_buf_2 fanout3911 (.A(net3912),
    .X(net3911));
 sg13g2_buf_2 fanout3912 (.A(net3923),
    .X(net3912));
 sg13g2_buf_2 fanout3913 (.A(net3914),
    .X(net3913));
 sg13g2_buf_2 fanout3914 (.A(net3923),
    .X(net3914));
 sg13g2_buf_4 fanout3915 (.X(net3915),
    .A(net3922));
 sg13g2_buf_1 fanout3916 (.A(net3922),
    .X(net3916));
 sg13g2_buf_2 fanout3917 (.A(net3918),
    .X(net3917));
 sg13g2_buf_2 fanout3918 (.A(net3922),
    .X(net3918));
 sg13g2_buf_4 fanout3919 (.X(net3919),
    .A(net3921));
 sg13g2_buf_1 fanout3920 (.A(net3921),
    .X(net3920));
 sg13g2_buf_4 fanout3921 (.X(net3921),
    .A(net3922));
 sg13g2_buf_2 fanout3922 (.A(net3923),
    .X(net3922));
 sg13g2_buf_2 fanout3923 (.A(net3924),
    .X(net3923));
 sg13g2_buf_2 fanout3924 (.A(net3992),
    .X(net3924));
 sg13g2_buf_4 fanout3925 (.X(net3925),
    .A(net3938));
 sg13g2_buf_4 fanout3926 (.X(net3926),
    .A(net3938));
 sg13g2_buf_4 fanout3927 (.X(net3927),
    .A(net3930));
 sg13g2_buf_2 fanout3928 (.A(net3930),
    .X(net3928));
 sg13g2_buf_4 fanout3929 (.X(net3929),
    .A(net3930));
 sg13g2_buf_2 fanout3930 (.A(net3938),
    .X(net3930));
 sg13g2_buf_2 fanout3931 (.A(net3932),
    .X(net3931));
 sg13g2_buf_4 fanout3932 (.X(net3932),
    .A(net3937));
 sg13g2_buf_2 fanout3933 (.A(net3934),
    .X(net3933));
 sg13g2_buf_2 fanout3934 (.A(net3937),
    .X(net3934));
 sg13g2_buf_2 fanout3935 (.A(net3937),
    .X(net3935));
 sg13g2_buf_2 fanout3936 (.A(net3937),
    .X(net3936));
 sg13g2_buf_1 fanout3937 (.A(net3938),
    .X(net3937));
 sg13g2_buf_2 fanout3938 (.A(net3991),
    .X(net3938));
 sg13g2_buf_4 fanout3939 (.X(net3939),
    .A(net3942));
 sg13g2_buf_2 fanout3940 (.A(net3941),
    .X(net3940));
 sg13g2_buf_2 fanout3941 (.A(net3942),
    .X(net3941));
 sg13g2_buf_2 fanout3942 (.A(net3954),
    .X(net3942));
 sg13g2_buf_4 fanout3943 (.X(net3943),
    .A(net3954));
 sg13g2_buf_4 fanout3944 (.X(net3944),
    .A(net3954));
 sg13g2_buf_4 fanout3945 (.X(net3945),
    .A(net3953));
 sg13g2_buf_1 fanout3946 (.A(net3953),
    .X(net3946));
 sg13g2_buf_4 fanout3947 (.X(net3947),
    .A(net3953));
 sg13g2_buf_2 fanout3948 (.A(net3952),
    .X(net3948));
 sg13g2_buf_2 fanout3949 (.A(net3952),
    .X(net3949));
 sg13g2_buf_4 fanout3950 (.X(net3950),
    .A(net3952));
 sg13g2_buf_2 fanout3951 (.A(net3952),
    .X(net3951));
 sg13g2_buf_1 fanout3952 (.A(net3953),
    .X(net3952));
 sg13g2_buf_2 fanout3953 (.A(net3954),
    .X(net3953));
 sg13g2_buf_2 fanout3954 (.A(net3991),
    .X(net3954));
 sg13g2_buf_2 fanout3955 (.A(net3958),
    .X(net3955));
 sg13g2_buf_1 fanout3956 (.A(net3958),
    .X(net3956));
 sg13g2_buf_4 fanout3957 (.X(net3957),
    .A(net3958));
 sg13g2_buf_2 fanout3958 (.A(net3973),
    .X(net3958));
 sg13g2_buf_2 fanout3959 (.A(net3960),
    .X(net3959));
 sg13g2_buf_2 fanout3960 (.A(net3963),
    .X(net3960));
 sg13g2_buf_2 fanout3961 (.A(net3962),
    .X(net3961));
 sg13g2_buf_2 fanout3962 (.A(net3963),
    .X(net3962));
 sg13g2_buf_1 fanout3963 (.A(net3973),
    .X(net3963));
 sg13g2_buf_2 fanout3964 (.A(net3966),
    .X(net3964));
 sg13g2_buf_2 fanout3965 (.A(net3966),
    .X(net3965));
 sg13g2_buf_2 fanout3966 (.A(net3967),
    .X(net3966));
 sg13g2_buf_4 fanout3967 (.X(net3967),
    .A(net3973));
 sg13g2_buf_2 fanout3968 (.A(net3972),
    .X(net3968));
 sg13g2_buf_2 fanout3969 (.A(net3971),
    .X(net3969));
 sg13g2_buf_1 fanout3970 (.A(net3971),
    .X(net3970));
 sg13g2_buf_2 fanout3971 (.A(net3972),
    .X(net3971));
 sg13g2_buf_2 fanout3972 (.A(net3973),
    .X(net3972));
 sg13g2_buf_2 fanout3973 (.A(net3991),
    .X(net3973));
 sg13g2_buf_2 fanout3974 (.A(net3977),
    .X(net3974));
 sg13g2_buf_2 fanout3975 (.A(net3977),
    .X(net3975));
 sg13g2_buf_2 fanout3976 (.A(net3977),
    .X(net3976));
 sg13g2_buf_2 fanout3977 (.A(net3990),
    .X(net3977));
 sg13g2_buf_4 fanout3978 (.X(net3978),
    .A(net3980));
 sg13g2_buf_4 fanout3979 (.X(net3979),
    .A(net3990));
 sg13g2_buf_2 fanout3980 (.A(net3990),
    .X(net3980));
 sg13g2_buf_2 fanout3981 (.A(net3989),
    .X(net3981));
 sg13g2_buf_2 fanout3982 (.A(net3989),
    .X(net3982));
 sg13g2_buf_4 fanout3983 (.X(net3983),
    .A(net3989));
 sg13g2_buf_4 fanout3984 (.X(net3984),
    .A(net3988));
 sg13g2_buf_1 fanout3985 (.A(net3988),
    .X(net3985));
 sg13g2_buf_4 fanout3986 (.X(net3986),
    .A(net3988));
 sg13g2_buf_2 fanout3987 (.A(net3988),
    .X(net3987));
 sg13g2_buf_2 fanout3988 (.A(net3989),
    .X(net3988));
 sg13g2_buf_2 fanout3989 (.A(net3990),
    .X(net3989));
 sg13g2_buf_2 fanout3990 (.A(net3991),
    .X(net3990));
 sg13g2_buf_4 fanout3991 (.X(net3991),
    .A(net3992));
 sg13g2_buf_8 fanout3992 (.A(_00000_),
    .X(net3992));
 sg13g2_buf_4 fanout3993 (.X(net3993),
    .A(_02198_));
 sg13g2_buf_2 fanout3994 (.A(net3995),
    .X(net3994));
 sg13g2_buf_2 fanout3995 (.A(_02184_),
    .X(net3995));
 sg13g2_buf_4 fanout3996 (.X(net3996),
    .A(net3998));
 sg13g2_buf_2 fanout3997 (.A(net3998),
    .X(net3997));
 sg13g2_buf_1 fanout3998 (.A(_02184_),
    .X(net3998));
 sg13g2_buf_2 fanout3999 (.A(net13),
    .X(net3999));
 sg13g2_buf_2 fanout4000 (.A(net4001),
    .X(net4000));
 sg13g2_buf_2 fanout4001 (.A(uio_in[2]),
    .X(net4001));
 sg13g2_buf_2 fanout4002 (.A(net4005),
    .X(net4002));
 sg13g2_buf_2 fanout4003 (.A(net4005),
    .X(net4003));
 sg13g2_buf_2 fanout4004 (.A(net4005),
    .X(net4004));
 sg13g2_buf_2 fanout4005 (.A(rst_n),
    .X(net4005));
 sg13g2_buf_2 fanout4006 (.A(net4010),
    .X(net4006));
 sg13g2_buf_2 fanout4007 (.A(net4010),
    .X(net4007));
 sg13g2_buf_4 fanout4008 (.X(net4008),
    .A(net4010));
 sg13g2_buf_2 fanout4009 (.A(net4010),
    .X(net4009));
 sg13g2_buf_2 fanout4010 (.A(rst_n),
    .X(net4010));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[3]),
    .X(net10));
 sg13g2_buf_4 input11 (.X(net11),
    .A(uio_in[5]));
 sg13g2_buf_4 input12 (.X(net12),
    .A(uio_in[6]));
 sg13g2_buf_2 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tielo tt_um_urish_sic1_14 (.L_LO(net14));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_2 clkbuf_leaf_42_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_2 clkbuf_leaf_43_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_2 clkbuf_leaf_44_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_2 clkbuf_leaf_45_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_2 clkbuf_leaf_46_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_2 clkbuf_leaf_47_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_2 clkbuf_leaf_48_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_2 clkbuf_leaf_49_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_2 clkbuf_leaf_50_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_2 clkbuf_leaf_51_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_2 clkbuf_leaf_52_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_2 clkbuf_leaf_53_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_2 clkbuf_leaf_54_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_2 clkbuf_leaf_55_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_2 clkbuf_leaf_56_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_2 clkbuf_leaf_57_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_2 clkbuf_leaf_58_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_2 clkbuf_leaf_59_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_2 clkbuf_leaf_60_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_2 clkbuf_leaf_61_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_2 clkbuf_leaf_62_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_2 clkbuf_leaf_63_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_2 clkbuf_leaf_64_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_2 clkbuf_leaf_65_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_2 clkbuf_leaf_66_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_2 clkbuf_leaf_67_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_2 clkbuf_leaf_68_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_2 clkbuf_leaf_69_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_2 clkbuf_leaf_70_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_2 clkbuf_leaf_71_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_2 clkbuf_leaf_72_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_2 clkbuf_leaf_73_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_2 clkbuf_leaf_74_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_2 clkbuf_leaf_75_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_2 clkbuf_leaf_76_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_2 clkbuf_leaf_77_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_2 clkbuf_leaf_78_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_2 clkbuf_leaf_79_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_2 clkbuf_leaf_80_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_2 clkbuf_leaf_81_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_2 clkbuf_leaf_82_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_2 clkbuf_leaf_83_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_2 clkbuf_leaf_84_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_2 clkbuf_leaf_85_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_2 clkbuf_leaf_86_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_2 clkbuf_leaf_87_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_2 clkbuf_leaf_88_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_2 clkbuf_leaf_89_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_2 clkbuf_leaf_90_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_2 clkbuf_leaf_91_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_2 clkbuf_leaf_92_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_2 clkbuf_leaf_93_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_2 clkbuf_leaf_94_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_2 clkbuf_leaf_95_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_2 clkbuf_leaf_96_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_2 clkbuf_leaf_97_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_2 clkbuf_leaf_98_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_2 clkbuf_leaf_99_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_2 clkbuf_leaf_100_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_2 clkbuf_leaf_101_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_2 clkbuf_leaf_102_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_2 clkbuf_leaf_103_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_2 clkbuf_leaf_104_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_2 clkbuf_leaf_105_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_2 clkbuf_leaf_106_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_2 clkbuf_leaf_107_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_2 clkbuf_leaf_108_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_2 clkbuf_leaf_109_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_2 clkbuf_leaf_110_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_2 clkbuf_leaf_111_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_2 clkbuf_leaf_112_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_2 clkbuf_leaf_113_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_2 clkbuf_leaf_114_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_2 clkbuf_leaf_115_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_2 clkbuf_leaf_116_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_2 clkbuf_leaf_117_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_2 clkbuf_leaf_118_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_2 clkbuf_leaf_119_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_2 clkbuf_leaf_120_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_2 clkbuf_leaf_121_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_2 clkbuf_leaf_122_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_2 clkbuf_leaf_123_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_2 clkbuf_leaf_124_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_2 clkbuf_leaf_125_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_2 clkbuf_leaf_126_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_2 clkbuf_leaf_127_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_2 clkbuf_leaf_128_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_2 clkbuf_leaf_129_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_2 clkbuf_leaf_130_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_2 clkbuf_leaf_131_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_2 clkbuf_leaf_132_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_2 clkbuf_leaf_133_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_2 clkbuf_leaf_134_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_2 clkbuf_leaf_135_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_2 clkbuf_leaf_136_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_2 clkbuf_leaf_137_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_2 clkbuf_leaf_138_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_2 clkbuf_leaf_139_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_2 clkbuf_leaf_140_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_2 clkbuf_leaf_141_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_2 clkbuf_leaf_142_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_2 clkbuf_leaf_143_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_2 clkbuf_leaf_144_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_2 clkbuf_leaf_145_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_2 clkbuf_leaf_146_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_2 clkbuf_leaf_147_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_2 clkbuf_leaf_148_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_2 clkbuf_leaf_149_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_2 clkbuf_leaf_150_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_2 clkbuf_leaf_151_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_2 clkbuf_leaf_152_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_2 clkbuf_leaf_153_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_2 clkbuf_leaf_154_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_2 clkbuf_leaf_155_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_2 clkbuf_leaf_156_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_2 clkbuf_leaf_157_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_2 clkbuf_leaf_158_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_2 clkbuf_leaf_159_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_2 clkbuf_leaf_160_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_2 clkbuf_leaf_161_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_2 clkbuf_leaf_162_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_2 clkbuf_leaf_163_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_2 clkbuf_leaf_164_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_2 clkbuf_leaf_165_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_2 clkbuf_leaf_166_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_2 clkbuf_leaf_167_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_2 clkbuf_leaf_168_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_2 clkbuf_leaf_169_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_2 clkbuf_leaf_170_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_2 clkbuf_leaf_171_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_2 clkbuf_leaf_172_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_2 clkbuf_leaf_173_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_2 clkbuf_leaf_174_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_2 clkbuf_leaf_175_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_2 clkbuf_leaf_176_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_2 clkbuf_leaf_177_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_2 clkbuf_leaf_178_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_2 clkbuf_leaf_179_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_2 clkbuf_leaf_180_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_2 clkbuf_leaf_181_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_2 clkbuf_leaf_182_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_2 clkbuf_leaf_183_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_2 clkbuf_leaf_184_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_2 clkbuf_leaf_185_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_2 clkbuf_leaf_186_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_2 clkbuf_leaf_187_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_2 clkbuf_leaf_188_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_2 clkbuf_leaf_189_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_2 clkbuf_leaf_190_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_2 clkbuf_leaf_191_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_2 clkbuf_leaf_192_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_2 clkbuf_leaf_193_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_2 clkbuf_leaf_194_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_2 clkbuf_leaf_195_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_2 clkbuf_leaf_196_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_2 clkbuf_leaf_197_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_2 clkbuf_leaf_198_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_2 clkbuf_leaf_199_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_2 clkbuf_leaf_200_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_2 clkbuf_leaf_201_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_2 clkbuf_leaf_202_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_2 clkbuf_leaf_203_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_2 clkbuf_leaf_204_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_2 clkbuf_leaf_205_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_2 clkbuf_leaf_206_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_2 clkbuf_leaf_207_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_2 clkbuf_leaf_208_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_2 clkbuf_leaf_209_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_2 clkbuf_leaf_210_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_2 clkbuf_leaf_211_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_2 clkbuf_leaf_212_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_2 clkbuf_leaf_213_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_2 clkbuf_leaf_214_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_2 clkbuf_leaf_215_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_2 clkbuf_leaf_216_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_2 clkbuf_leaf_217_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_2 clkbuf_leaf_218_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_2 clkbuf_leaf_219_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_2 clkbuf_leaf_220_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_2 clkbuf_leaf_221_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_2 clkbuf_leaf_222_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_2 clkbuf_leaf_223_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_2 clkbuf_leaf_224_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_2 clkbuf_leaf_225_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_2 clkbuf_leaf_226_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_2 clkbuf_leaf_227_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_2 clkbuf_leaf_228_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_2 clkbuf_leaf_229_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_2 clkbuf_leaf_230_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_2 clkbuf_leaf_231_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_2 clkbuf_leaf_232_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_2 clkbuf_leaf_233_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_2 clkbuf_leaf_234_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_2 clkbuf_leaf_235_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_2 clkbuf_leaf_236_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_2 clkbuf_leaf_237_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_2 clkbuf_leaf_238_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_2 clkbuf_leaf_239_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_2 clkbuf_leaf_240_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_2 clkbuf_leaf_241_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_2 clkbuf_leaf_242_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_2 clkbuf_leaf_243_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_2 clkbuf_leaf_244_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_2 clkbuf_leaf_245_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_2 clkbuf_leaf_246_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_2 clkbuf_leaf_247_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_2 clkbuf_leaf_248_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_2 clkbuf_leaf_249_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_2 clkbuf_leaf_250_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_2 clkbuf_leaf_251_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_2 clkbuf_leaf_252_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_2 clkbuf_leaf_253_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_2 clkbuf_leaf_254_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_2 clkbuf_leaf_255_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_2 clkbuf_leaf_256_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_2 clkbuf_leaf_257_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_2 clkbuf_leaf_258_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_2 clkbuf_leaf_259_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_2 clkbuf_leaf_260_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_2 clkbuf_leaf_261_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_2 clkbuf_leaf_262_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_2 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_2 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_2 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_2 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_2 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_2 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_2 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_2 clkbuf_6_0__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_0__leaf_clk));
 sg13g2_buf_2 clkbuf_6_1__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_1__leaf_clk));
 sg13g2_buf_2 clkbuf_6_2__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_2__leaf_clk));
 sg13g2_buf_2 clkbuf_6_3__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_3__leaf_clk));
 sg13g2_buf_2 clkbuf_6_4__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_4__leaf_clk));
 sg13g2_buf_2 clkbuf_6_5__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_5__leaf_clk));
 sg13g2_buf_2 clkbuf_6_6__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_6__leaf_clk));
 sg13g2_buf_2 clkbuf_6_7__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_6_7__leaf_clk));
 sg13g2_buf_2 clkbuf_6_8__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_8__leaf_clk));
 sg13g2_buf_2 clkbuf_6_9__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_9__leaf_clk));
 sg13g2_buf_2 clkbuf_6_10__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_10__leaf_clk));
 sg13g2_buf_2 clkbuf_6_11__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_11__leaf_clk));
 sg13g2_buf_2 clkbuf_6_12__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_12__leaf_clk));
 sg13g2_buf_2 clkbuf_6_13__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_13__leaf_clk));
 sg13g2_buf_2 clkbuf_6_14__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_14__leaf_clk));
 sg13g2_buf_2 clkbuf_6_15__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_6_15__leaf_clk));
 sg13g2_buf_2 clkbuf_6_16__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_16__leaf_clk));
 sg13g2_buf_2 clkbuf_6_17__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_17__leaf_clk));
 sg13g2_buf_2 clkbuf_6_18__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_18__leaf_clk));
 sg13g2_buf_2 clkbuf_6_19__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_19__leaf_clk));
 sg13g2_buf_2 clkbuf_6_20__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_20__leaf_clk));
 sg13g2_buf_2 clkbuf_6_21__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_21__leaf_clk));
 sg13g2_buf_2 clkbuf_6_22__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_22__leaf_clk));
 sg13g2_buf_2 clkbuf_6_23__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_6_23__leaf_clk));
 sg13g2_buf_2 clkbuf_6_24__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_24__leaf_clk));
 sg13g2_buf_2 clkbuf_6_25__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_25__leaf_clk));
 sg13g2_buf_2 clkbuf_6_26__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_26__leaf_clk));
 sg13g2_buf_2 clkbuf_6_27__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_27__leaf_clk));
 sg13g2_buf_2 clkbuf_6_28__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_28__leaf_clk));
 sg13g2_buf_2 clkbuf_6_29__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_29__leaf_clk));
 sg13g2_buf_2 clkbuf_6_30__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_30__leaf_clk));
 sg13g2_buf_2 clkbuf_6_31__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_6_31__leaf_clk));
 sg13g2_buf_2 clkbuf_6_32__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_32__leaf_clk));
 sg13g2_buf_2 clkbuf_6_33__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_33__leaf_clk));
 sg13g2_buf_2 clkbuf_6_34__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_34__leaf_clk));
 sg13g2_buf_2 clkbuf_6_35__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_35__leaf_clk));
 sg13g2_buf_2 clkbuf_6_36__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_36__leaf_clk));
 sg13g2_buf_2 clkbuf_6_37__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_37__leaf_clk));
 sg13g2_buf_2 clkbuf_6_38__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_38__leaf_clk));
 sg13g2_buf_2 clkbuf_6_39__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_6_39__leaf_clk));
 sg13g2_buf_2 clkbuf_6_40__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_40__leaf_clk));
 sg13g2_buf_2 clkbuf_6_41__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_41__leaf_clk));
 sg13g2_buf_2 clkbuf_6_42__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_42__leaf_clk));
 sg13g2_buf_2 clkbuf_6_43__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_43__leaf_clk));
 sg13g2_buf_2 clkbuf_6_44__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_44__leaf_clk));
 sg13g2_buf_2 clkbuf_6_45__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_45__leaf_clk));
 sg13g2_buf_2 clkbuf_6_46__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_46__leaf_clk));
 sg13g2_buf_2 clkbuf_6_47__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_6_47__leaf_clk));
 sg13g2_buf_2 clkbuf_6_48__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_48__leaf_clk));
 sg13g2_buf_2 clkbuf_6_49__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_49__leaf_clk));
 sg13g2_buf_2 clkbuf_6_50__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_50__leaf_clk));
 sg13g2_buf_2 clkbuf_6_51__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_51__leaf_clk));
 sg13g2_buf_2 clkbuf_6_52__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_52__leaf_clk));
 sg13g2_buf_2 clkbuf_6_53__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_53__leaf_clk));
 sg13g2_buf_2 clkbuf_6_54__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_54__leaf_clk));
 sg13g2_buf_2 clkbuf_6_55__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_6_55__leaf_clk));
 sg13g2_buf_2 clkbuf_6_56__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_56__leaf_clk));
 sg13g2_buf_2 clkbuf_6_57__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_57__leaf_clk));
 sg13g2_buf_2 clkbuf_6_58__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_58__leaf_clk));
 sg13g2_buf_2 clkbuf_6_59__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_59__leaf_clk));
 sg13g2_buf_2 clkbuf_6_60__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_60__leaf_clk));
 sg13g2_buf_2 clkbuf_6_61__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_61__leaf_clk));
 sg13g2_buf_2 clkbuf_6_62__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_62__leaf_clk));
 sg13g2_buf_2 clkbuf_6_63__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_6_63__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_6_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_6_2__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_6_3__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_6_4__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_6_5__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_6_6__leaf_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_2 clkload7 (.A(clknet_6_9__leaf_clk));
 sg13g2_buf_2 clkload8 (.A(clknet_6_10__leaf_clk));
 sg13g2_buf_2 clkload9 (.A(clknet_6_11__leaf_clk));
 sg13g2_buf_2 clkload10 (.A(clknet_6_12__leaf_clk));
 sg13g2_buf_2 clkload11 (.A(clknet_6_13__leaf_clk));
 sg13g2_buf_2 clkload12 (.A(clknet_6_14__leaf_clk));
 sg13g2_buf_2 clkload13 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_2 clkload14 (.A(clknet_6_17__leaf_clk));
 sg13g2_buf_2 clkload15 (.A(clknet_6_18__leaf_clk));
 sg13g2_buf_2 clkload16 (.A(clknet_6_19__leaf_clk));
 sg13g2_buf_2 clkload17 (.A(clknet_6_20__leaf_clk));
 sg13g2_buf_2 clkload18 (.A(clknet_6_21__leaf_clk));
 sg13g2_buf_2 clkload19 (.A(clknet_6_22__leaf_clk));
 sg13g2_buf_2 clkload20 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_2 clkload21 (.A(clknet_6_25__leaf_clk));
 sg13g2_buf_2 clkload22 (.A(clknet_6_26__leaf_clk));
 sg13g2_buf_2 clkload23 (.A(clknet_6_27__leaf_clk));
 sg13g2_buf_2 clkload24 (.A(clknet_6_28__leaf_clk));
 sg13g2_buf_2 clkload25 (.A(clknet_6_29__leaf_clk));
 sg13g2_buf_2 clkload26 (.A(clknet_6_30__leaf_clk));
 sg13g2_buf_2 clkload27 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_2 clkload28 (.A(clknet_6_33__leaf_clk));
 sg13g2_buf_2 clkload29 (.A(clknet_6_34__leaf_clk));
 sg13g2_buf_2 clkload30 (.A(clknet_6_35__leaf_clk));
 sg13g2_buf_2 clkload31 (.A(clknet_6_36__leaf_clk));
 sg13g2_buf_2 clkload32 (.A(clknet_6_37__leaf_clk));
 sg13g2_buf_2 clkload33 (.A(clknet_6_38__leaf_clk));
 sg13g2_buf_2 clkload34 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_2 clkload35 (.A(clknet_6_41__leaf_clk));
 sg13g2_buf_2 clkload36 (.A(clknet_6_42__leaf_clk));
 sg13g2_buf_2 clkload37 (.A(clknet_6_43__leaf_clk));
 sg13g2_buf_2 clkload38 (.A(clknet_6_44__leaf_clk));
 sg13g2_buf_2 clkload39 (.A(clknet_6_45__leaf_clk));
 sg13g2_buf_2 clkload40 (.A(clknet_6_46__leaf_clk));
 sg13g2_buf_2 clkload41 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_2 clkload42 (.A(clknet_6_49__leaf_clk));
 sg13g2_buf_2 clkload43 (.A(clknet_6_50__leaf_clk));
 sg13g2_buf_2 clkload44 (.A(clknet_6_51__leaf_clk));
 sg13g2_buf_2 clkload45 (.A(clknet_6_52__leaf_clk));
 sg13g2_buf_2 clkload46 (.A(clknet_6_53__leaf_clk));
 sg13g2_buf_2 clkload47 (.A(clknet_6_54__leaf_clk));
 sg13g2_buf_2 clkload48 (.A(clknet_6_55__leaf_clk));
 sg13g2_inv_2 clkload49 (.A(clknet_leaf_262_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\mem.wr_en ),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold2 (.A(_00838_),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold3 (.A(\mem.mem[196][4] ),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold4 (.A(\C[7] ),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold5 (.A(\mem.mem[140][5] ),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold6 (.A(\mem.mem[68][5] ),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold7 (.A(\mem.mem[78][6] ),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold8 (.A(\mem.mem[70][6] ),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold9 (.A(\mem.mem[98][5] ),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold10 (.A(\mem.mem[134][5] ),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold11 (.A(\mem.mem[44][6] ),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold12 (.A(\C[2] ),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold13 (.A(\mem.mem[228][4] ),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold14 (.A(\mem.mem[212][4] ),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold15 (.A(\mem.mem[76][6] ),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold16 (.A(\mem.mem[206][6] ),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold17 (.A(\mem.mem[132][5] ),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold18 (.A(\mem.mem[68][6] ),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold19 (.A(\mem.uo_out[2] ),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold20 (.A(\mem.mem[212][5] ),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold21 (.A(\mem.mem[206][5] ),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold22 (.A(\mem.mem[228][5] ),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold23 (.A(\mem.mem[84][4] ),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold24 (.A(\mem.mem[72][1] ),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold25 (.A(\mem.mem[176][2] ),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold26 (.A(\mem.mem[94][5] ),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold27 (.A(\mem.mem[76][2] ),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold28 (.A(\mem.mem[130][5] ),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold29 (.A(\mem.mem[44][5] ),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold30 (.A(\mem.mem[196][5] ),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold31 (.A(\mem.mem[70][4] ),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold32 (.A(\mem.mem[70][5] ),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold33 (.A(\mem.mem[88][6] ),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold34 (.A(\mem.mem[116][5] ),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold35 (.A(\mem.mem[38][2] ),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold36 (.A(\mem.mem[228][3] ),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold37 (.A(\mem.mem[62][6] ),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold38 (.A(\mem.uo_out[5] ),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold39 (.A(\mem.mem[244][1] ),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold40 (.A(\mem.mem[132][7] ),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold41 (.A(\mem.mem[144][2] ),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold42 (.A(\mem.mem[62][5] ),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold43 (.A(\mem.mem[116][6] ),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold44 (.A(\mem.mem[46][7] ),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold45 (.A(\mem.mem[56][3] ),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold46 (.A(\mem.mem[84][6] ),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold47 (.A(\mem.mem[116][1] ),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold48 (.A(\mem.uo_out[6] ),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold49 (.A(\mem.mem[140][0] ),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold50 (.A(\mem.mem[52][0] ),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold51 (.A(\mem.mem[62][7] ),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold52 (.A(\mem.mem[116][2] ),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold53 (.A(\mem.mem[52][6] ),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold54 (.A(\mem.mem[46][6] ),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold55 (.A(\mem.mem[52][5] ),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold56 (.A(\mem.mem[94][6] ),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold57 (.A(\mem.mem[140][4] ),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold58 (.A(\mem.mem[40][2] ),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold59 (.A(\mem.mem[228][0] ),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold60 (.A(\mem.mem[98][1] ),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold61 (.A(\mem.mem[136][2] ),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold62 (.A(\mem.mem[222][7] ),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold63 (.A(\mem.mem[244][5] ),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold64 (.A(\mem.mem[116][4] ),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold65 (.A(\mem.mem[69][4] ),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold66 (.A(\mem.mem[136][3] ),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold67 (.A(\mem.mem[104][5] ),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold68 (.A(\mem.mem[249][2] ),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold69 (.A(\mem.mem[191][6] ),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold70 (.A(\mem.mem[160][5] ),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold71 (.A(\mem.mem[206][2] ),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold72 (.A(\mem.mem[56][0] ),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold73 (.A(\mem.mem[228][6] ),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold74 (.A(\mem.uo_out[0] ),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold75 (.A(_00839_),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold76 (.A(\mem.mem[176][1] ),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold77 (.A(\mem.mem[246][6] ),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold78 (.A(\mem.mem[160][3] ),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold79 (.A(\mem.mem[176][5] ),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold80 (.A(\mem.mem[98][7] ),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold81 (.A(\mem.mem[212][7] ),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold82 (.A(\mem.mem[63][4] ),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold83 (.A(\mem.mem[136][1] ),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold84 (.A(\mem.mem[88][3] ),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold85 (.A(\mem.mem[133][1] ),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold86 (.A(\mem.mem[250][5] ),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold87 (.A(\mem.mem[144][3] ),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold88 (.A(\mem.mem[95][0] ),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold89 (.A(\mem.mem[132][0] ),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold90 (.A(\mem.mem[159][0] ),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold91 (.A(\mem.mem[239][0] ),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold92 (.A(\mem.mem[174][5] ),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold93 (.A(\mem.mem[4][2] ),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold94 (.A(\mem.mem[241][2] ),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold95 (.A(\mem.mem[223][5] ),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold96 (.A(\mem.mem[245][2] ),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold97 (.A(\mem.mem[110][6] ),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold98 (.A(\mem.mem[129][1] ),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold99 (.A(\mem.mem[116][0] ),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold100 (.A(\mem.mem[212][6] ),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold101 (.A(\mem.mem[196][7] ),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold102 (.A(\mem.mem[252][7] ),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold103 (.A(\mem.mem[245][1] ),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold104 (.A(\mem.mem[241][6] ),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold105 (.A(\mem.mem[116][7] ),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold106 (.A(\mem.mem[120][4] ),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold107 (.A(\mem.mem[232][7] ),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold108 (.A(\mem.mem[193][3] ),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold109 (.A(\mem.mem[245][5] ),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold110 (.A(\mem.mem[113][1] ),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold111 (.A(\mem.mem[251][6] ),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold112 (.A(\mem.mem[249][5] ),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold113 (.A(\mem.mem[52][2] ),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold114 (.A(\mem.mem[246][0] ),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold115 (.A(\mem.mem[81][7] ),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold116 (.A(\mem.mem[28][6] ),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold117 (.A(\mem.mem[196][2] ),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold118 (.A(\mem.mem[132][4] ),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold119 (.A(\mem.mem[209][3] ),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold120 (.A(\mem.mem[143][2] ),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold121 (.A(\mem.mem[228][1] ),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold122 (.A(\mem.mem[63][1] ),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold123 (.A(\mem.mem[70][7] ),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold124 (.A(\mem.mem[252][1] ),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold125 (.A(\mem.mem[138][0] ),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold126 (.A(\mem.mem[251][4] ),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold127 (.A(\mem.mem[249][0] ),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold128 (.A(\mem.mem[63][7] ),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold129 (.A(\mem.mem[131][6] ),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold130 (.A(\mem.mem[175][6] ),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold131 (.A(\mem.mem[232][0] ),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold132 (.A(\mem.mem[223][7] ),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold133 (.A(\mem.mem[93][1] ),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold134 (.A(\mem.mem[193][6] ),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold135 (.A(\mem.mem[28][7] ),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold136 (.A(\mem.mem[207][7] ),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold137 (.A(\mem.mem[104][1] ),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold138 (.A(\mem.mem[88][1] ),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold139 (.A(\mem.mem[196][1] ),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold140 (.A(\mem.mem[252][4] ),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold141 (.A(\mem.mem[175][4] ),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold142 (.A(\mem.mem[94][1] ),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold143 (.A(\mem.mem[248][4] ),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold144 (.A(\mem.mem[241][3] ),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold145 (.A(\mem.mem[136][0] ),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold146 (.A(\mem.mem[239][6] ),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold147 (.A(\mem.mem[251][0] ),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold148 (.A(\mem.mem[15][5] ),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold149 (.A(\mem.mem[131][3] ),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold150 (.A(\mem.mem[121][5] ),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold151 (.A(\mem.mem[191][4] ),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold152 (.A(\mem.mem[138][1] ),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold153 (.A(\mem.mem[56][6] ),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold154 (.A(\mem.mem[63][6] ),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold155 (.A(\mem.mem[136][4] ),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold156 (.A(\mem.mem[205][1] ),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold157 (.A(\mem.mem[244][0] ),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold158 (.A(\mem.mem[140][6] ),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold159 (.A(\mem.mem[84][7] ),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold160 (.A(\mem.mem[68][7] ),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold161 (.A(\mem.mem[94][4] ),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold162 (.A(\mem.mem[73][6] ),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold163 (.A(\mem.mem[88][2] ),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold164 (.A(\mem.mem[76][0] ),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold165 (.A(\mem.mem[175][7] ),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold166 (.A(\mem.mem[79][5] ),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold167 (.A(\mem.mem[65][0] ),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold168 (.A(\mem.mem[129][7] ),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold169 (.A(\mem.mem[111][7] ),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold170 (.A(\mem.mem[63][5] ),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold171 (.A(\mem.mem[245][3] ),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold172 (.A(\mem.mem[113][3] ),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold173 (.A(\mem.mem[127][1] ),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold174 (.A(\mem.mem[79][0] ),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold175 (.A(\mem.mem[223][3] ),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold176 (.A(\mem.mem[98][4] ),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold177 (.A(\mem.mem[97][7] ),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold178 (.A(\mem.mem[175][0] ),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold179 (.A(\mem.mem[212][1] ),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold180 (.A(\mem.mem[104][2] ),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold181 (.A(\mem.mem[137][2] ),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold182 (.A(\mem.mem[131][7] ),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold183 (.A(\mem.mem[134][0] ),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold184 (.A(\mem.mem[133][6] ),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold185 (.A(\mem.mem[93][2] ),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold186 (.A(\mem.mem[209][6] ),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold187 (.A(\mem.mem[89][7] ),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold188 (.A(\mem.mem[95][4] ),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold189 (.A(\mem.mem[206][1] ),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold190 (.A(\mem.mem[160][2] ),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold191 (.A(\mem.mem[200][2] ),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold192 (.A(\mem.mem[200][1] ),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold193 (.A(\mem.mem[252][2] ),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold194 (.A(\mem.mem[72][7] ),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold195 (.A(\mem.mem[209][7] ),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold196 (.A(\mem.mem[207][1] ),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold197 (.A(\mem.mem[225][1] ),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold198 (.A(\mem.mem[56][1] ),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold199 (.A(\mem.mem[28][5] ),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold200 (.A(\mem.mem[228][7] ),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold201 (.A(\mem.mem[130][7] ),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold202 (.A(\mem.mem[250][0] ),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold203 (.A(\mem.mem[252][0] ),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold204 (.A(\mem.mem[52][4] ),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold205 (.A(\mem.mem[201][1] ),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold206 (.A(\mem.mem[133][7] ),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold207 (.A(\mem.mem[127][2] ),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold208 (.A(\mem.mem[93][0] ),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold209 (.A(\mem.mem[121][1] ),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold210 (.A(\mem.mem[73][5] ),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold211 (.A(\mem.mem[44][4] ),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold212 (.A(\mem.mem[138][5] ),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold213 (.A(\mem.mem[223][6] ),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold214 (.A(\mem.mem[137][6] ),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold215 (.A(\mem.mem[78][5] ),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold216 (.A(\mem.mem[246][1] ),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold217 (.A(\mem.mem[111][6] ),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold218 (.A(\mem.mem[111][2] ),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold219 (.A(\mem.mem[244][6] ),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold220 (.A(\mem.mem[65][5] ),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold221 (.A(\mem.mem[251][3] ),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold222 (.A(\mem.mem[72][0] ),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold223 (.A(\mem.mem[134][6] ),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold224 (.A(\mem.mem[212][0] ),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold225 (.A(\mem.mem[120][2] ),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold226 (.A(\mem.mem[132][3] ),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold227 (.A(\mem.mem[121][2] ),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold228 (.A(\mem.mem[134][3] ),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold229 (.A(\mem.mem[95][3] ),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold230 (.A(\mem.mem[69][0] ),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold231 (.A(\mem.mem[143][4] ),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold232 (.A(\mem.uo_out[4] ),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold233 (.A(\mem.mem[131][2] ),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold234 (.A(\mem.mem[97][4] ),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold235 (.A(\mem.mem[232][1] ),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold236 (.A(\mem.mem[127][6] ),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold237 (.A(\mem.mem[76][4] ),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold238 (.A(\mem.mem[129][3] ),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold239 (.A(\mem.mem[200][0] ),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold240 (.A(\mem.mem[196][3] ),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold241 (.A(\mem.mem[232][3] ),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold242 (.A(\mem.mem[176][4] ),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold243 (.A(\mem.mem[143][7] ),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold244 (.A(\mem.mem[76][1] ),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold245 (.A(\mem.mem[95][1] ),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold246 (.A(\mem.mem[78][2] ),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold247 (.A(\mem.mem[143][1] ),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold248 (.A(\mem.mem[206][4] ),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold249 (.A(\mem.mem[98][3] ),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold250 (.A(\mem.mem[176][6] ),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold251 (.A(\mem.mem[201][6] ),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold252 (.A(\mem.mem[121][3] ),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold253 (.A(\mem.mem[134][2] ),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold254 (.A(\mem.mem[113][4] ),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold255 (.A(\mem.mem[113][5] ),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold256 (.A(\mem.mem[73][4] ),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold257 (.A(\mem.mem[68][1] ),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold258 (.A(\mem.mem[98][2] ),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold259 (.A(\mem.mem[137][1] ),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold260 (.A(\mem.mem[159][5] ),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold261 (.A(\mem.mem[239][7] ),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold262 (.A(\mem.mem[241][5] ),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold263 (.A(\mem.mem[245][7] ),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold264 (.A(\mem.mem[40][4] ),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold265 (.A(\mem.mem[176][7] ),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold266 (.A(\mem.mem[65][3] ),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold267 (.A(\mem.mem[193][0] ),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold268 (.A(\mem.mem[251][2] ),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold269 (.A(\mem.mem[249][4] ),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold270 (.A(\mem.mem[70][0] ),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold271 (.A(\mem.mem[132][1] ),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold272 (.A(\mem.mem[134][4] ),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold273 (.A(\mem.mem[250][7] ),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold274 (.A(\mem.mem[120][5] ),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold275 (.A(\mem.mem[251][5] ),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold276 (.A(\mem.mem[143][0] ),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold277 (.A(\mem.mem[28][2] ),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold278 (.A(\mem.mem[244][4] ),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold279 (.A(\mem.mem[44][0] ),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold280 (.A(\mem.mem[15][7] ),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold281 (.A(\mem.mem[52][7] ),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold282 (.A(\mem.mem[200][6] ),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold283 (.A(\mem.mem[97][5] ),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold284 (.A(\mem.mem[84][0] ),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold285 (.A(\mem.mem[79][3] ),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold286 (.A(\mem.mem[239][1] ),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold287 (.A(\mem.mem[133][3] ),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold288 (.A(\mem.mem[127][4] ),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold289 (.A(\mem.mem[40][6] ),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold290 (.A(\mem.mem[249][3] ),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold291 (.A(\mem.mem[251][1] ),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold292 (.A(\mem.mem[246][2] ),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold293 (.A(\mem.mem[28][4] ),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold294 (.A(\mem.mem[193][7] ),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold295 (.A(\mem.mem[137][0] ),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold296 (.A(\mem.mem[223][2] ),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold297 (.A(\mem.mem[63][3] ),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold298 (.A(\mem.mem[132][2] ),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold299 (.A(\mem.mem[249][7] ),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold300 (.A(\mem.mem[127][7] ),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold301 (.A(\mem.mem[131][4] ),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold302 (.A(\mem.mem[193][2] ),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold303 (.A(\mem.mem[138][4] ),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold304 (.A(\mem.mem[84][3] ),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold305 (.A(\mem.mem[79][6] ),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold306 (.A(\mem.mem[76][3] ),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold307 (.A(\mem.mem[72][6] ),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold308 (.A(\mem.mem[52][3] ),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold309 (.A(\mem.mem[138][7] ),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold310 (.A(\mem.mem[94][3] ),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold311 (.A(\mem.mem[44][7] ),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold312 (.A(\mem.mem[246][4] ),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold313 (.A(\mem.mem[56][4] ),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold314 (.A(\mem.mem[249][6] ),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold315 (.A(\mem.mem[81][4] ),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold316 (.A(\mem.mem[132][6] ),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold317 (.A(\mem.mem[65][7] ),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold318 (.A(\mem.mem[207][0] ),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold319 (.A(\mem.mem[223][1] ),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold320 (.A(\mem.mem[130][6] ),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold321 (.A(\mem.mem[249][1] ),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold322 (.A(\mem.mem[225][2] ),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold323 (.A(\mem.mem[246][3] ),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold324 (.A(\mem.mem[40][3] ),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold325 (.A(\mem.mem[65][2] ),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold326 (.A(\mem.mem[68][2] ),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold327 (.A(\mem.mem[104][0] ),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold328 (.A(\mem.mem[160][4] ),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold329 (.A(\mem.mem[190][7] ),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold330 (.A(\mem.mem[120][1] ),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold331 (.A(\mem.mem[191][0] ),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold332 (.A(\mem.mem[28][3] ),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold333 (.A(\mem.mem[201][4] ),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold334 (.A(\mem.mem[111][1] ),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold335 (.A(\mem.mem[250][2] ),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold336 (.A(\mem.mem[28][0] ),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold337 (.A(\mem.mem[225][6] ),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold338 (.A(\mem.mem[250][6] ),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold339 (.A(\mem.mem[89][0] ),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold340 (.A(\mem.mem[73][7] ),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold341 (.A(\mem.mem[40][5] ),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold342 (.A(\mem.mem[206][7] ),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold343 (.A(\mem.mem[191][1] ),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold344 (.A(\mem.mem[138][2] ),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold345 (.A(\mem.mem[239][4] ),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold346 (.A(\mem.mem[78][3] ),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold347 (.A(\mem.mem[245][6] ),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold348 (.A(\mem.mem[73][0] ),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold349 (.A(\mem.mem[70][1] ),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold350 (.A(\mem.mem[130][1] ),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold351 (.A(\mem.mem[95][7] ),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold352 (.A(\mem.mem[93][4] ),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold353 (.A(\mem.mem[250][1] ),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold354 (.A(\mem.mem[28][1] ),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold355 (.A(\mem.mem[160][1] ),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold356 (.A(\mem.mem[104][3] ),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold357 (.A(\mem.mem[89][6] ),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold358 (.A(\mem.mem[130][3] ),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold359 (.A(\mem.mem[248][3] ),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold360 (.A(\mem.mem[129][2] ),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold361 (.A(\mem.mem[121][6] ),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold362 (.A(\mem.mem[176][0] ),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold363 (.A(\mem.mem[196][6] ),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold364 (.A(\mem.mem[144][5] ),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold365 (.A(\mem.mem[79][7] ),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold366 (.A(\mem.mem[78][4] ),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold367 (.A(\mem.mem[73][2] ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold368 (.A(\mem.mem[245][4] ),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold369 (.A(\mem.mem[79][1] ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold370 (.A(\mem.mem[127][5] ),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold371 (.A(\mem.mem[68][0] ),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold372 (.A(\mem.mem[73][1] ),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold373 (.A(\mem.mem[144][0] ),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold374 (.A(\mem.mem[81][0] ),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold375 (.A(\mem.mem[212][3] ),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold376 (.A(\mem.mem[207][6] ),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold377 (.A(\mem.mem[140][2] ),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold378 (.A(\mem.mem[207][2] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold379 (.A(\mem.mem[40][1] ),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold380 (.A(\mem.mem[206][0] ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold381 (.A(\mem.mem[201][2] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold382 (.A(\mem.mem[73][3] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold383 (.A(\mem.mem[113][7] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold384 (.A(\mem.mem[134][1] ),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold385 (.A(\mem.mem[95][5] ),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold386 (.A(\mem.mem[143][3] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold387 (.A(\mem.mem[133][4] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold388 (.A(\mem.mem[248][7] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold389 (.A(\mem.mem[205][4] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold390 (.A(\mem.mem[159][6] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold391 (.A(\mem.mem[69][2] ),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold392 (.A(\mem.mem[93][7] ),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold393 (.A(\mem.mem[131][1] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold394 (.A(\mem.mem[113][2] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold395 (.A(\mem.mem[209][2] ),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold396 (.A(\mem.mem[97][6] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold397 (.A(\mem.mem[137][4] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold398 (.A(\mem.mem[97][0] ),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold399 (.A(\mem.mem[209][1] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold400 (.A(\mem.mem[130][0] ),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold401 (.A(\mem.mem[140][3] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold402 (.A(\mem.mem[97][3] ),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold403 (.A(\mem.mem[225][7] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold404 (.A(\mem.mem[200][7] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold405 (.A(\mem.mem[129][6] ),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold406 (.A(\mem.mem[84][1] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold407 (.A(\mem.mem[72][4] ),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold408 (.A(\mem.mem[104][6] ),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold409 (.A(\mem.mem[201][0] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold410 (.A(\mem.mem[44][2] ),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold411 (.A(\mem.mem[252][3] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold412 (.A(\mem.mem[205][7] ),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold413 (.A(\mem.mem[160][7] ),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold414 (.A(\mem.mem[79][4] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold415 (.A(\mem.mem[205][2] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold416 (.A(\mem.mem[137][5] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold417 (.A(\mem.mem[40][0] ),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold418 (.A(\mem.mem[68][3] ),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold419 (.A(\mem.mem[138][6] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold420 (.A(\mem.mem[136][5] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold421 (.A(\mem.mem[143][5] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold422 (.A(\mem.mem[72][3] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold423 (.A(\mem.mem[246][5] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold424 (.A(\mem.mem[160][0] ),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold425 (.A(\mem.mem[121][0] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold426 (.A(\mem.mem[176][3] ),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold427 (.A(\mem.mem[69][1] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold428 (.A(\mem.mem[248][2] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold429 (.A(\mem.mem[252][5] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold430 (.A(\mem.mem[89][3] ),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold431 (.A(\mem.mem[159][7] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold432 (.A(\mem.mem[191][5] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold433 (.A(\mem.mem[250][3] ),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold434 (.A(\mem.mem[245][0] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold435 (.A(\mem.mem[140][7] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold436 (.A(\mem.mem[250][4] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold437 (.A(\mem.mem[225][0] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold438 (.A(\mem.mem[223][0] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold439 (.A(\mem.mem[120][3] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold440 (.A(\mem.mem[232][5] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold441 (.A(\mem.mem[248][1] ),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold442 (.A(\mem.mem[120][0] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold443 (.A(\mem.mem[15][1] ),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold444 (.A(\mem.mem[200][4] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold445 (.A(\mem.mem[241][7] ),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold446 (.A(\mem.mem[97][2] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold447 (.A(\mem.mem[81][3] ),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold448 (.A(\mem.mem[138][3] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold449 (.A(\mem.mem[72][5] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold450 (.A(\mem.mem[68][4] ),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold451 (.A(\mem.mem[244][3] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold452 (.A(\mem.mem[69][3] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold453 (.A(\mem.mem[16][1] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold454 (.A(\mem.mem[111][5] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold455 (.A(\mem.mem[40][7] ),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold456 (.A(\mem.mem[69][7] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold457 (.A(\mem.mem[248][0] ),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold458 (.A(\mem.mem[134][7] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold459 (.A(\mem.mem[209][0] ),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold460 (.A(\mem.mem[239][5] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold461 (.A(\mem.mem[56][5] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold462 (.A(\mem.mem[191][3] ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold463 (.A(\mem.mem[95][2] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold464 (.A(\mem.mem[225][3] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold465 (.A(\mem.mem[78][1] ),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold466 (.A(\mem.mem[56][2] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold467 (.A(\mem.mem[88][0] ),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold468 (.A(\mem.mem[204][5] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold469 (.A(\mem.mem[252][6] ),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold470 (.A(\mem.mem[241][1] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold471 (.A(\mem.mem[159][2] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold472 (.A(\mem.mem[63][0] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold473 (.A(\mem.mem[201][5] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold474 (.A(\mem.mem[120][6] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold475 (.A(\mem.mem[20][4] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold476 (.A(\mem.mem[130][4] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold477 (.A(\mem.mem[121][4] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold478 (.A(\mem.mem[127][3] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold479 (.A(\mem.mem[186][1] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold480 (.A(\mem.mem[244][7] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold481 (.A(\mem.mem[175][2] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold482 (.A(\mem.mem[79][2] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold483 (.A(\mem.mem[140][1] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold484 (.A(\mem.mem[223][4] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold485 (.A(\mem.mem[212][2] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold486 (.A(\mem.mem[89][4] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold487 (.A(\C[6] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold488 (.A(\mem.mem[78][0] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold489 (.A(\mem.mem[193][5] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold490 (.A(\mem.mem[201][3] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold491 (.A(\mem.mem[72][2] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold492 (.A(\mem.mem[159][1] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold493 (.A(\mem.mem[201][7] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold494 (.A(\mem.mem[228][2] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold495 (.A(\mem.mem[70][3] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold496 (.A(\mem.mem[6][5] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold497 (.A(\mem.mem[180][6] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold498 (.A(\mem.mem[225][5] ),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold499 (.A(\mem.mem[88][7] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold500 (.A(\mem.mem[232][2] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold501 (.A(\mem.mem[111][4] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold502 (.A(\mem.uo_out[7] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold503 (.A(\mem.mem[22][3] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold504 (.A(\mem.mem[108][6] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold505 (.A(\mem.mem[246][7] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold506 (.A(\mem.mem[65][1] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold507 (.A(\mem.mem[76][5] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold508 (.A(\mem.mem[20][6] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold509 (.A(\mem.mem[131][5] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold510 (.A(\mem.mem[236][4] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold511 (.A(\mem.mem[207][3] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold512 (.A(\mem.mem[48][3] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold513 (.A(\mem.mem[121][7] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold514 (.A(\mem.mem[191][7] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold515 (.A(\mem.mem[230][2] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold516 (.A(\mem.mem[44][3] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold517 (.A(\mem.mem[136][6] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold518 (.A(\mem.mem[112][0] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold519 (.A(\mem.mem[251][7] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold520 (.A(\mem.mem[196][0] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold521 (.A(\mem.mem[63][2] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold522 (.A(\mem.mem[81][6] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold523 (.A(\mem.mem[225][4] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold524 (.A(\mem.mem[193][4] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold525 (.A(\mem.mem[137][3] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold526 (.A(\A[7] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold527 (.A(_00602_),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold528 (.A(\mem.mem[104][4] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold529 (.A(\mem.mem[93][3] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold530 (.A(\mem.mem[18][1] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold531 (.A(\mem.mem[76][7] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold532 (.A(\mem.mem[113][6] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold533 (.A(\mem.mem[81][5] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold534 (.A(\mem.mem[131][0] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold535 (.A(\mem.mem[193][1] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold536 (.A(\mem.mem[104][7] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold537 (.A(\mem.mem[164][2] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold538 (.A(\mem.mem[159][3] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold539 (.A(\mem.mem[241][4] ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold540 (.A(\mem.mem[133][5] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold541 (.A(\mem.mem[133][2] ),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold542 (.A(\mem.mem[81][1] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold543 (.A(\mem.mem[162][2] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold544 (.A(\A[2] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold545 (.A(_00597_),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold546 (.A(\mem.mem[69][5] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold547 (.A(\mem.mem[144][6] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold548 (.A(\mem.mem[207][5] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold549 (.A(\mem.mem[65][4] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold550 (.A(\mem.mem[206][3] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold551 (.A(\mem.mem[56][7] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold552 (.A(\mem.mem[89][2] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold553 (.A(\mem.mem[93][5] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold554 (.A(\mem.mem[64][5] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold555 (.A(\mem.mem[148][6] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold556 (.A(\mem.mem[144][1] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold557 (.A(\mem.mem[239][2] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold558 (.A(\mem.mem[248][5] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold559 (.A(\mem.mem[89][5] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold560 (.A(\mem.mem[144][4] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold561 (.A(\mem.mem[200][3] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold562 (.A(\mem.mem[144][7] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold563 (.A(\mem.mem[192][5] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold564 (.A(\mem.mem[96][1] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold565 (.A(\mem.mem[175][5] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold566 (.A(\mem.mem[15][3] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold567 (.A(\mem.mem[209][5] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold568 (.A(\mem.mem[111][0] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold569 (.A(\mem.mem[174][3] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold570 (.A(\mem.mem[22][4] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold571 (.A(\mem.mem[97][1] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold572 (.A(\mem.mem[2][5] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold573 (.A(\mem.mem[168][4] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold574 (.A(\mem.mem[182][2] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold575 (.A(\mem.mem[92][5] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold576 (.A(\mem.mem[16][6] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold577 (.A(\mem.mem[95][6] ),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold578 (.A(\mem.mem[62][2] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold579 (.A(\mem.mem[172][5] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold580 (.A(\mem.mem[114][0] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold581 (.A(\mem.mem[6][4] ),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold582 (.A(\mem.mem[15][0] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold583 (.A(\mem.mem[244][2] ),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold584 (.A(\mem.mem[16][4] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold585 (.A(\mem.mem[94][0] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold586 (.A(\mem.mem[98][0] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold587 (.A(\mem.mem[230][5] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold588 (.A(\mem.mem[46][5] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold589 (.A(\mem.mem[84][2] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold590 (.A(\mem.mem[207][4] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold591 (.A(\mem.mem[70][2] ),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold592 (.A(\mem.mem[0][6] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold593 (.A(\mem.mem[232][4] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold594 (.A(\mem.mem[205][6] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold595 (.A(\mem.mem[98][6] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold596 (.A(\mem.mem[208][4] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold597 (.A(\mem.mem[150][5] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold598 (.A(\mem.mem[84][5] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold599 (.A(\mem.mem[216][1] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold600 (.A(\mem.mem[86][1] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold601 (.A(\mem.mem[12][5] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold602 (.A(\mem.mem[48][2] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold603 (.A(\mem.mem[22][7] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold604 (.A(\mem.mem[60][7] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold605 (.A(\mem.mem[111][3] ),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold606 (.A(\mem.mem[4][6] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold607 (.A(\mem.mem[88][4] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold608 (.A(\mem.mem[137][7] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold609 (.A(\mem.mem[222][4] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold610 (.A(\mem.mem[92][4] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold611 (.A(\mem.mem[15][4] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold612 (.A(\mem.mem[93][6] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold613 (.A(\mem.mem[15][6] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold614 (.A(\mem.mem[178][2] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold615 (.A(\mem.mem[129][0] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold616 (.A(\mem.mem[218][1] ),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold617 (.A(\mem.mem[214][5] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold618 (.A(\mem.mem[116][3] ),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold619 (.A(\mem.mem[166][6] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold620 (.A(\mem.mem[133][0] ),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold621 (.A(\mem.mem[126][0] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold622 (.A(\mem.mem[136][7] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold623 (.A(\mem.mem[89][1] ),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold624 (.A(\mem.mem[130][2] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold625 (.A(\mem.mem[69][6] ),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold626 (.A(\mem.mem[241][0] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold627 (.A(\mem.mem[154][4] ),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold628 (.A(\mem.mem[175][1] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold629 (.A(\mem.mem[65][6] ),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold630 (.A(\mem.mem[18][4] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold631 (.A(\mem.mem[20][7] ),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold632 (.A(\mem.mem[188][6] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold633 (.A(\mem.mem[14][0] ),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold634 (.A(\mem.mem[198][4] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold635 (.A(\mem.mem[175][3] ),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold636 (.A(\mem.mem[129][4] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold637 (.A(\mem.mem[172][6] ),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold638 (.A(\mem.mem[191][2] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold639 (.A(\mem.mem[194][4] ),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold640 (.A(\mem.mem[143][6] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold641 (.A(\mem.mem[81][2] ),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold642 (.A(\mem.mem[174][1] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold643 (.A(\mem.mem[238][1] ),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold644 (.A(\mem.mem[216][2] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold645 (.A(\mem.mem[204][2] ),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold646 (.A(\mem.mem[186][4] ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold647 (.A(\mem.mem[78][7] ),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold648 (.A(\mem.mem[38][1] ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold649 (.A(\mem.mem[248][6] ),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold650 (.A(\mem.mem[6][6] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold651 (.A(\mem.mem[159][4] ),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold652 (.A(\mem.mem[92][6] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold653 (.A(\A[6] ),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold654 (.A(_00601_),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold655 (.A(\mem.mem[184][0] ),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold656 (.A(\mem.mem[224][0] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold657 (.A(\mem.mem[110][0] ),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold658 (.A(\mem.mem[74][1] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold659 (.A(\mem.mem[0][4] ),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold660 (.A(\mem.mem[194][5] ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold661 (.A(\mem.mem[14][4] ),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold662 (.A(\mem.mem[62][0] ),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold663 (.A(\mem.mem[129][5] ),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold664 (.A(\mem.mem[152][1] ),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold665 (.A(\mem.mem[12][4] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold666 (.A(\mem.mem[170][4] ),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold667 (.A(\mem.mem[232][6] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold668 (.A(\mem.mem[194][1] ),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold669 (.A(\mem.mem[198][6] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold670 (.A(\mem.mem[220][7] ),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold671 (.A(\mem.mem[2][6] ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold672 (.A(\mem.mem[205][3] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold673 (.A(\mem.mem[205][0] ),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold674 (.A(\mem.mem[184][1] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold675 (.A(\mem.mem[180][0] ),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold676 (.A(\mem.mem[236][0] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold677 (.A(\mem.mem[160][6] ),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold678 (.A(\mem.mem[100][5] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold679 (.A(\mem.mem[127][0] ),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold680 (.A(\mem.mem[52][1] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold681 (.A(\mem.mem[44][1] ),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold682 (.A(\mem.mem[96][5] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold683 (.A(\mem.mem[106][5] ),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold684 (.A(\mem.mem[66][6] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold685 (.A(\mem.mem[58][3] ),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold686 (.A(\mem.mem[239][3] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold687 (.A(\mem.mem[50][3] ),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold688 (.A(\mem.mem[210][5] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold689 (.A(\mem.mem[86][4] ),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold690 (.A(\mem.mem[113][0] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold691 (.A(\mem.mem[208][2] ),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold692 (.A(\mem.mem[230][4] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold693 (.A(\mem.mem[226][4] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold694 (.A(\mem.mem[204][6] ),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold695 (.A(\mem.mem[124][5] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold696 (.A(\mem.mem[0][5] ),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold697 (.A(\mem.mem[46][0] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold698 (.A(\mem.mem[124][0] ),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold699 (.A(\mem.mem[4][5] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold700 (.A(\mem.mem[192][4] ),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold701 (.A(\mem.mem[208][5] ),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold702 (.A(\mem.mem[128][5] ),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold703 (.A(\mem.mem[238][3] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold704 (.A(\mem.mem[180][2] ),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold705 (.A(\mem.mem[2][4] ),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold706 (.A(\mem.mem[209][4] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold707 (.A(\mem.mem[188][2] ),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold708 (.A(\mem.mem[15][2] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold709 (.A(\mem.mem[224][4] ),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold710 (.A(\mem.mem[20][3] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold711 (.A(\mem.mem[205][5] ),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold712 (.A(\mem.mem[236][5] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold713 (.A(\mem.mem[14][6] ),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold714 (.A(\mem.mem[88][5] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold715 (.A(\mem.mem[12][6] ),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold716 (.A(\mem.mem[172][0] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold717 (.A(\mem.mem[50][2] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold718 (.A(\mem.mem[200][5] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold719 (.A(\mem.mem[22][6] ),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold720 (.A(\mem.mem[142][6] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold721 (.A(\mem.mem[142][5] ),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold722 (.A(\mem.mem[80][3] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold723 (.A(\mem.mem[54][1] ),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold724 (.A(\mem.mem[226][5] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold725 (.A(\mem.mem[18][6] ),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold726 (.A(\mem.mem[152][3] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold727 (.A(\mem.mem[110][2] ),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold728 (.A(\mem.mem[192][7] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold729 (.A(\mem.mem[226][0] ),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold730 (.A(\mem.mem[214][4] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold731 (.A(\mem.mem[172][2] ),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold732 (.A(_01473_),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold733 (.A(\mem.mem[90][6] ),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold734 (.A(\mem.mem[198][5] ),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold735 (.A(\mem.mem[186][0] ),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold736 (.A(\mem.mem[220][4] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold737 (.A(\mem.mem[174][2] ),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold738 (.A(\mem.mem[36][6] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold739 (.A(\mem.mem[92][7] ),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold740 (.A(\mem.mem[120][7] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold741 (.A(\mem.mem[110][5] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold742 (.A(\mem.mem[154][1] ),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold743 (.A(\mem.mem[110][4] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold744 (.A(\mem.mem[184][4] ),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold745 (.A(\mem.mem[4][0] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold746 (.A(\mem.mem[182][6] ),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold747 (.A(\mem.mem[60][2] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold748 (.A(\mem.mem[166][0] ),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold749 (.A(\mem.mem[192][1] ),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold750 (.A(\mem.mem[238][5] ),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold751 (.A(\mem.mem[142][3] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold752 (.A(\mem.mem[157][2] ),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold753 (.A(\mem.mem[158][3] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold754 (.A(\mem.mem[164][3] ),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold755 (.A(\mem.mem[36][5] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold756 (.A(\mem.mem[82][3] ),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold757 (.A(\mem.mem[54][7] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold758 (.A(\mem.mem[20][2] ),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold759 (.A(\mem.mem[210][4] ),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold760 (.A(\mem.mem[102][3] ),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold761 (.A(\mem.mem[208][7] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold762 (.A(\mem.mem[36][7] ),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold763 (.A(\mem.mem[149][5] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold764 (.A(\mem.mem[213][2] ),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold765 (.A(\mem.mem[238][4] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold766 (.A(\mem.mem[53][3] ),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold767 (.A(\mem.mem[156][4] ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold768 (.A(\mem.mem[0][0] ),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold769 (.A(\mem.mem[172][4] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold770 (.A(\mem.mem[122][2] ),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold771 (.A(\mem.mem[184][7] ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold772 (.A(\mem.mem[222][1] ),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold773 (.A(\mem.mem[157][5] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold774 (.A(\mem.mem[164][5] ),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold775 (.A(\mem.mem[50][7] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold776 (.A(\mem.mem[94][2] ),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold777 (.A(\mem.mem[135][0] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold778 (.A(\mem.mem[166][4] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold779 (.A(\mem.mem[150][4] ),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold780 (.A(\mem.mem[103][0] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold781 (.A(\mem.mem[30][2] ),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold782 (.A(\mem.mem[48][4] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold783 (.A(\mem.mem[151][1] ),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold784 (.A(\mem.mem[33][4] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold785 (.A(\mem.mem[109][0] ),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold786 (.A(\mem.mem[92][3] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold787 (.A(\mem.mem[163][0] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold788 (.A(\mem.mem[167][4] ),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold789 (.A(\mem.mem[25][4] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold790 (.A(\mem.mem[158][1] ),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold791 (.A(\mem.mem[96][7] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold792 (.A(\mem.mem[64][6] ),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold793 (.A(\mem.mem[170][3] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold794 (.A(\mem.mem[36][4] ),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold795 (.A(\mem.mem[170][1] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold796 (.A(\mem.mem[110][7] ),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold797 (.A(\mem.mem[48][6] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold798 (.A(\mem.mem[5][0] ),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold799 (.A(\mem.mem[118][1] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold800 (.A(\mem.mem[148][7] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold801 (.A(\mem.mem[59][6] ),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold802 (.A(\mem.mem[106][0] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold803 (.A(\mem.mem[242][3] ),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold804 (.A(\mem.mem[183][1] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold805 (.A(\mem.mem[25][7] ),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold806 (.A(\mem.mem[192][6] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold807 (.A(\mem.mem[218][5] ),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold808 (.A(\mem.mem[231][0] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold809 (.A(\mem.mem[156][2] ),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold810 (.A(\mem.mem[74][3] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold811 (.A(\mem.mem[186][3] ),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold812 (.A(\mem.mem[100][4] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold813 (.A(\mem.mem[161][7] ),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold814 (.A(\mem.mem[27][6] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold815 (.A(\mem.mem[106][3] ),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold816 (.A(\mem.mem[153][2] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold817 (.A(\mem.mem[103][5] ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold818 (.A(\mem.mem[14][1] ),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold819 (.A(\mem.mem[230][1] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold820 (.A(\mem.mem[197][6] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold821 (.A(\mem.mem[222][0] ),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold822 (.A(\mem.mem[218][0] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold823 (.A(\mem.mem[182][4] ),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold824 (.A(\mem.mem[37][1] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold825 (.A(\mem.mem[180][7] ),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold826 (.A(\mem.mem[148][2] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold827 (.A(\mem.mem[74][5] ),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold828 (.A(\mem.mem[59][0] ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold829 (.A(\mem.mem[105][1] ),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold830 (.A(\mem.mem[57][0] ),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold831 (.A(\mem.mem[33][2] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold832 (.A(\mem.mem[39][6] ),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold833 (.A(\mem.mem[96][3] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold834 (.A(\mem.mem[216][5] ),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold835 (.A(\mem.mem[237][3] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold836 (.A(\mem.mem[16][7] ),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold837 (.A(\mem.mem[234][2] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold838 (.A(\mem.mem[16][5] ),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold839 (.A(\mem.mem[210][2] ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold840 (.A(\mem.mem[100][6] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold841 (.A(\mem.mem[96][4] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold842 (.A(\mem.mem[96][6] ),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold843 (.A(\mem.mem[38][7] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold844 (.A(\mem.mem[20][5] ),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold845 (.A(\mem.mem[25][6] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold846 (.A(\mem.mem[150][0] ),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold847 (.A(\mem.mem[16][0] ),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold848 (.A(\mem.mem[187][7] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold849 (.A(\mem.mem[107][0] ),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold850 (.A(\mem.mem[224][6] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold851 (.A(\mem.mem[220][5] ),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold852 (.A(\mem.mem[165][4] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold853 (.A(\mem.mem[157][0] ),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold854 (.A(\mem.mem[199][1] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold855 (.A(\mem.mem[149][7] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold856 (.A(\mem.mem[60][0] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold857 (.A(\mem.mem[151][6] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold858 (.A(\mem.mem[42][6] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold859 (.A(\mem.mem[177][6] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold860 (.A(\mem.mem[231][1] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold861 (.A(\mem.mem[100][0] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold862 (.A(\mem.mem[215][0] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold863 (.A(\mem.mem[27][5] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold864 (.A(\mem.mem[187][3] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold865 (.A(\mem.mem[107][1] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold866 (.A(\mem.mem[43][4] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold867 (.A(\mem.mem[155][2] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold868 (.A(\mem.mem[112][6] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold869 (.A(\mem.mem[123][2] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold870 (.A(\mem.mem[112][4] ),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold871 (.A(\mem.mem[142][4] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold872 (.A(\mem.mem[210][3] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold873 (.A(\mem.mem[234][4] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold874 (.A(\mem.mem[181][1] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold875 (.A(\mem.mem[142][1] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold876 (.A(\mem.mem[161][2] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold877 (.A(\mem.mem[163][5] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold878 (.A(\mem.mem[126][6] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold879 (.A(\mem.mem[203][1] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold880 (.A(\mem.mem[32][5] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold881 (.A(\mem.mem[171][7] ),
    .X(net4011));
 sg13g2_dlygate4sd3_1 hold882 (.A(\mem.mem[157][6] ),
    .X(net4012));
 sg13g2_dlygate4sd3_1 hold883 (.A(\mem.mem[224][3] ),
    .X(net4013));
 sg13g2_dlygate4sd3_1 hold884 (.A(\mem.mem[21][1] ),
    .X(net4014));
 sg13g2_dlygate4sd3_1 hold885 (.A(\mem.mem[202][7] ),
    .X(net4015));
 sg13g2_dlygate4sd3_1 hold886 (.A(\mem.mem[148][3] ),
    .X(net4016));
 sg13g2_dlygate4sd3_1 hold887 (.A(\mem.mem[185][5] ),
    .X(net4017));
 sg13g2_dlygate4sd3_1 hold888 (.A(\mem.mem[43][6] ),
    .X(net4018));
 sg13g2_dlygate4sd3_1 hold889 (.A(\mem.mem[66][5] ),
    .X(net4019));
 sg13g2_dlygate4sd3_1 hold890 (.A(\mem.mem[23][0] ),
    .X(net4020));
 sg13g2_dlygate4sd3_1 hold891 (.A(\mem.mem[142][0] ),
    .X(net4021));
 sg13g2_dlygate4sd3_1 hold892 (.A(\mem.mem[18][3] ),
    .X(net4022));
 sg13g2_dlygate4sd3_1 hold893 (.A(\mem.mem[60][6] ),
    .X(net4023));
 sg13g2_dlygate4sd3_1 hold894 (.A(\mem.mem[211][1] ),
    .X(net4024));
 sg13g2_dlygate4sd3_1 hold895 (.A(\mem.mem[238][7] ),
    .X(net4025));
 sg13g2_dlygate4sd3_1 hold896 (.A(\mem.mem[247][7] ),
    .X(net4026));
 sg13g2_dlygate4sd3_1 hold897 (.A(\mem.mem[31][6] ),
    .X(net4027));
 sg13g2_dlygate4sd3_1 hold898 (.A(\mem.mem[153][0] ),
    .X(net4028));
 sg13g2_dlygate4sd3_1 hold899 (.A(\mem.mem[48][5] ),
    .X(net4029));
 sg13g2_dlygate4sd3_1 hold900 (.A(\mem.mem[188][7] ),
    .X(net4030));
 sg13g2_dlygate4sd3_1 hold901 (.A(\mem.mem[231][7] ),
    .X(net4031));
 sg13g2_dlygate4sd3_1 hold902 (.A(\mem.mem[224][5] ),
    .X(net4032));
 sg13g2_dlygate4sd3_1 hold903 (.A(\mem.mem[21][0] ),
    .X(net4033));
 sg13g2_dlygate4sd3_1 hold904 (.A(\mem.mem[151][4] ),
    .X(net4034));
 sg13g2_dlygate4sd3_1 hold905 (.A(\mem.mem[94][7] ),
    .X(net4035));
 sg13g2_dlygate4sd3_1 hold906 (.A(\mem.mem[198][7] ),
    .X(net4036));
 sg13g2_dlygate4sd3_1 hold907 (.A(\mem.mem[128][6] ),
    .X(net4037));
 sg13g2_dlygate4sd3_1 hold908 (.A(\mem.mem[122][1] ),
    .X(net4038));
 sg13g2_dlygate4sd3_1 hold909 (.A(\mem.mem[170][5] ),
    .X(net4039));
 sg13g2_dlygate4sd3_1 hold910 (.A(\mem.mem[218][7] ),
    .X(net4040));
 sg13g2_dlygate4sd3_1 hold911 (.A(\mem.mem[38][5] ),
    .X(net4041));
 sg13g2_dlygate4sd3_1 hold912 (.A(\mem.mem[102][0] ),
    .X(net4042));
 sg13g2_dlygate4sd3_1 hold913 (.A(\mem.mem[202][3] ),
    .X(net4043));
 sg13g2_dlygate4sd3_1 hold914 (.A(\mem.mem[55][7] ),
    .X(net4044));
 sg13g2_dlygate4sd3_1 hold915 (.A(\mem.mem[32][6] ),
    .X(net4045));
 sg13g2_dlygate4sd3_1 hold916 (.A(\mem.mem[155][7] ),
    .X(net4046));
 sg13g2_dlygate4sd3_1 hold917 (.A(\mem.mem[163][1] ),
    .X(net4047));
 sg13g2_dlygate4sd3_1 hold918 (.A(\mem.mem[190][5] ),
    .X(net4048));
 sg13g2_dlygate4sd3_1 hold919 (.A(\mem.mem[123][5] ),
    .X(net4049));
 sg13g2_dlygate4sd3_1 hold920 (.A(\mem.mem[123][6] ),
    .X(net4050));
 sg13g2_dlygate4sd3_1 hold921 (.A(\mem.mem[158][0] ),
    .X(net4051));
 sg13g2_dlygate4sd3_1 hold922 (.A(\mem.mem[221][0] ),
    .X(net4052));
 sg13g2_dlygate4sd3_1 hold923 (.A(\mem.mem[240][0] ),
    .X(net4053));
 sg13g2_dlygate4sd3_1 hold924 (.A(\mem.mem[4][1] ),
    .X(net4054));
 sg13g2_dlygate4sd3_1 hold925 (.A(\mem.mem[59][2] ),
    .X(net4055));
 sg13g2_dlygate4sd3_1 hold926 (.A(\mem.mem[114][5] ),
    .X(net4056));
 sg13g2_dlygate4sd3_1 hold927 (.A(\mem.mem[101][7] ),
    .X(net4057));
 sg13g2_dlygate4sd3_1 hold928 (.A(\mem.mem[235][0] ),
    .X(net4058));
 sg13g2_dlygate4sd3_1 hold929 (.A(\mem.mem[204][0] ),
    .X(net4059));
 sg13g2_dlygate4sd3_1 hold930 (.A(\mem.mem[230][7] ),
    .X(net4060));
 sg13g2_dlygate4sd3_1 hold931 (.A(\mem.mem[152][4] ),
    .X(net4061));
 sg13g2_dlygate4sd3_1 hold932 (.A(\mem.mem[199][2] ),
    .X(net4062));
 sg13g2_dlygate4sd3_1 hold933 (.A(\mem.mem[199][3] ),
    .X(net4063));
 sg13g2_dlygate4sd3_1 hold934 (.A(\mem.mem[99][3] ),
    .X(net4064));
 sg13g2_dlygate4sd3_1 hold935 (.A(\mem.mem[100][3] ),
    .X(net4065));
 sg13g2_dlygate4sd3_1 hold936 (.A(\mem.mem[33][0] ),
    .X(net4066));
 sg13g2_dlygate4sd3_1 hold937 (.A(\mem.mem[184][2] ),
    .X(net4067));
 sg13g2_dlygate4sd3_1 hold938 (.A(\mem.mem[221][2] ),
    .X(net4068));
 sg13g2_dlygate4sd3_1 hold939 (.A(\mem.mem[197][2] ),
    .X(net4069));
 sg13g2_dlygate4sd3_1 hold940 (.A(\mem.mem[165][5] ),
    .X(net4070));
 sg13g2_dlygate4sd3_1 hold941 (.A(\mem.mem[82][7] ),
    .X(net4071));
 sg13g2_dlygate4sd3_1 hold942 (.A(\mem.mem[150][7] ),
    .X(net4072));
 sg13g2_dlygate4sd3_1 hold943 (.A(\mem.mem[219][2] ),
    .X(net4073));
 sg13g2_dlygate4sd3_1 hold944 (.A(\mem.mem[90][0] ),
    .X(net4074));
 sg13g2_dlygate4sd3_1 hold945 (.A(\mem.mem[156][5] ),
    .X(net4075));
 sg13g2_dlygate4sd3_1 hold946 (.A(\mem.mem[31][4] ),
    .X(net4076));
 sg13g2_dlygate4sd3_1 hold947 (.A(\mem.mem[210][7] ),
    .X(net4077));
 sg13g2_dlygate4sd3_1 hold948 (.A(\mem.mem[43][0] ),
    .X(net4078));
 sg13g2_dlygate4sd3_1 hold949 (.A(\mem.mem[146][7] ),
    .X(net4079));
 sg13g2_dlygate4sd3_1 hold950 (.A(\mem.mem[218][3] ),
    .X(net4080));
 sg13g2_dlygate4sd3_1 hold951 (.A(\mem.mem[7][0] ),
    .X(net4081));
 sg13g2_dlygate4sd3_1 hold952 (.A(\mem.mem[105][0] ),
    .X(net4082));
 sg13g2_dlygate4sd3_1 hold953 (.A(\mem.mem[148][1] ),
    .X(net4083));
 sg13g2_dlygate4sd3_1 hold954 (.A(\mem.mem[229][7] ),
    .X(net4084));
 sg13g2_dlygate4sd3_1 hold955 (.A(\mem.mem[99][6] ),
    .X(net4085));
 sg13g2_dlygate4sd3_1 hold956 (.A(\mem.mem[203][5] ),
    .X(net4086));
 sg13g2_dlygate4sd3_1 hold957 (.A(\mem.mem[155][3] ),
    .X(net4087));
 sg13g2_dlygate4sd3_1 hold958 (.A(\mem.mem[179][5] ),
    .X(net4088));
 sg13g2_dlygate4sd3_1 hold959 (.A(\mem.mem[24][6] ),
    .X(net4089));
 sg13g2_dlygate4sd3_1 hold960 (.A(\mem.mem[57][4] ),
    .X(net4090));
 sg13g2_dlygate4sd3_1 hold961 (.A(\mem.mem[61][4] ),
    .X(net4091));
 sg13g2_dlygate4sd3_1 hold962 (.A(\mem.mem[86][6] ),
    .X(net4092));
 sg13g2_dlygate4sd3_1 hold963 (.A(\mem.mem[83][5] ),
    .X(net4093));
 sg13g2_dlygate4sd3_1 hold964 (.A(\mem.mem[47][1] ),
    .X(net4094));
 sg13g2_dlygate4sd3_1 hold965 (.A(\mem.mem[101][6] ),
    .X(net4095));
 sg13g2_dlygate4sd3_1 hold966 (.A(\mem.mem[82][0] ),
    .X(net4096));
 sg13g2_dlygate4sd3_1 hold967 (.A(\mem.mem[216][6] ),
    .X(net4097));
 sg13g2_dlygate4sd3_1 hold968 (.A(\mem.mem[215][6] ),
    .X(net4098));
 sg13g2_dlygate4sd3_1 hold969 (.A(\mem.mem[166][1] ),
    .X(net4099));
 sg13g2_dlygate4sd3_1 hold970 (.A(\mem.mem[32][4] ),
    .X(net4100));
 sg13g2_dlygate4sd3_1 hold971 (.A(\mem.mem[198][0] ),
    .X(net4101));
 sg13g2_dlygate4sd3_1 hold972 (.A(\mem.mem[183][4] ),
    .X(net4102));
 sg13g2_dlygate4sd3_1 hold973 (.A(\mem.mem[177][0] ),
    .X(net4103));
 sg13g2_dlygate4sd3_1 hold974 (.A(\mem.mem[177][7] ),
    .X(net4104));
 sg13g2_dlygate4sd3_1 hold975 (.A(\mem.mem[67][1] ),
    .X(net4105));
 sg13g2_dlygate4sd3_1 hold976 (.A(\mem.mem[82][1] ),
    .X(net4106));
 sg13g2_dlygate4sd3_1 hold977 (.A(\mem.mem[21][5] ),
    .X(net4107));
 sg13g2_dlygate4sd3_1 hold978 (.A(\mem.mem[109][4] ),
    .X(net4108));
 sg13g2_dlygate4sd3_1 hold979 (.A(\mem.mem[181][7] ),
    .X(net4109));
 sg13g2_dlygate4sd3_1 hold980 (.A(\mem.mem[39][0] ),
    .X(net4110));
 sg13g2_dlygate4sd3_1 hold981 (.A(\mem.mem[39][2] ),
    .X(net4111));
 sg13g2_dlygate4sd3_1 hold982 (.A(\mem.mem[235][4] ),
    .X(net4112));
 sg13g2_dlygate4sd3_1 hold983 (.A(\mem.mem[31][0] ),
    .X(net4113));
 sg13g2_dlygate4sd3_1 hold984 (.A(\mem.mem[146][6] ),
    .X(net4114));
 sg13g2_dlygate4sd3_1 hold985 (.A(\mem.mem[151][7] ),
    .X(net4115));
 sg13g2_dlygate4sd3_1 hold986 (.A(\mem.mem[11][3] ),
    .X(net4116));
 sg13g2_dlygate4sd3_1 hold987 (.A(\mem.mem[222][3] ),
    .X(net4117));
 sg13g2_dlygate4sd3_1 hold988 (.A(\mem.mem[107][3] ),
    .X(net4118));
 sg13g2_dlygate4sd3_1 hold989 (.A(\mem.mem[135][2] ),
    .X(net4119));
 sg13g2_dlygate4sd3_1 hold990 (.A(\mem.mem[171][6] ),
    .X(net4120));
 sg13g2_dlygate4sd3_1 hold991 (.A(\mem.mem[29][1] ),
    .X(net4121));
 sg13g2_dlygate4sd3_1 hold992 (.A(\mem.mem[139][2] ),
    .X(net4122));
 sg13g2_dlygate4sd3_1 hold993 (.A(\mem.mem[47][3] ),
    .X(net4123));
 sg13g2_dlygate4sd3_1 hold994 (.A(\mem.mem[172][7] ),
    .X(net4124));
 sg13g2_dlygate4sd3_1 hold995 (.A(\mem.mem[187][6] ),
    .X(net4125));
 sg13g2_dlygate4sd3_1 hold996 (.A(\mem.mem[204][1] ),
    .X(net4126));
 sg13g2_dlygate4sd3_1 hold997 (.A(\mem.mem[80][0] ),
    .X(net4127));
 sg13g2_dlygate4sd3_1 hold998 (.A(\mem.mem[13][1] ),
    .X(net4128));
 sg13g2_dlygate4sd3_1 hold999 (.A(\mem.mem[243][3] ),
    .X(net4129));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\mem.mem[162][6] ),
    .X(net4130));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\mem.mem[4][3] ),
    .X(net4131));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\mem.mem[10][6] ),
    .X(net4132));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\mem.mem[158][4] ),
    .X(net4133));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\mem.mem[162][7] ),
    .X(net4134));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\mem.mem[150][6] ),
    .X(net4135));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\mem.mem[149][1] ),
    .X(net4136));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\mem.mem[22][5] ),
    .X(net4137));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\mem.mem[35][6] ),
    .X(net4138));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\mem.mem[185][2] ),
    .X(net4139));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\mem.mem[57][1] ),
    .X(net4140));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\mem.mem[49][4] ),
    .X(net4141));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\mem.mem[7][7] ),
    .X(net4142));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\mem.mem[233][0] ),
    .X(net4143));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\mem.mem[216][3] ),
    .X(net4144));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\mem.mem[90][5] ),
    .X(net4145));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\mem.mem[181][5] ),
    .X(net4146));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\mem.mem[219][6] ),
    .X(net4147));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\mem.mem[219][4] ),
    .X(net4148));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\mem.mem[145][1] ),
    .X(net4149));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\mem.mem[38][0] ),
    .X(net4150));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\mem.mem[236][6] ),
    .X(net4151));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\mem.mem[227][6] ),
    .X(net4152));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\mem.mem[188][3] ),
    .X(net4153));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\mem.mem[220][2] ),
    .X(net4154));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\mem.mem[211][0] ),
    .X(net4155));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\mem.mem[29][6] ),
    .X(net4156));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\mem.mem[167][7] ),
    .X(net4157));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\mem.mem[36][1] ),
    .X(net4158));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\mem.mem[19][7] ),
    .X(net4159));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\mem.mem[53][0] ),
    .X(net4160));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\mem.mem[24][2] ),
    .X(net4161));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\mem.mem[4][7] ),
    .X(net4162));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\mem.mem[184][6] ),
    .X(net4163));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\mem.mem[243][2] ),
    .X(net4164));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\mem.mem[135][7] ),
    .X(net4165));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\mem.mem[30][7] ),
    .X(net4166));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\mem.mem[117][6] ),
    .X(net4167));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\mem.mem[31][3] ),
    .X(net4168));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\mem.mem[77][1] ),
    .X(net4169));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\mem.mem[192][2] ),
    .X(net4170));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\mem.mem[55][6] ),
    .X(net4171));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\mem.mem[8][6] ),
    .X(net4172));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\mem.mem[86][7] ),
    .X(net4173));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\mem.mem[106][7] ),
    .X(net4174));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\mem.mem[83][4] ),
    .X(net4175));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\mem.mem[49][1] ),
    .X(net4176));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\mem.mem[170][7] ),
    .X(net4177));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\mem.mem[12][7] ),
    .X(net4178));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\mem.mem[103][1] ),
    .X(net4179));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\mem.mem[161][5] ),
    .X(net4180));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\mem.mem[9][6] ),
    .X(net4181));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\mem.mem[102][4] ),
    .X(net4182));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\mem.mem[235][3] ),
    .X(net4183));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\mem.mem[64][0] ),
    .X(net4184));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\mem.mem[62][4] ),
    .X(net4185));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\mem.mem[197][0] ),
    .X(net4186));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\mem.mem[114][3] ),
    .X(net4187));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\mem.mem[114][7] ),
    .X(net4188));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\mem.mem[103][3] ),
    .X(net4189));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\mem.mem[26][2] ),
    .X(net4190));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\mem.mem[158][7] ),
    .X(net4191));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\mem.mem[115][7] ),
    .X(net4192));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\mem.mem[213][6] ),
    .X(net4193));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\mem.mem[0][7] ),
    .X(net4194));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\mem.mem[18][5] ),
    .X(net4195));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\mem.mem[162][5] ),
    .X(net4196));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\mem.mem[147][5] ),
    .X(net4197));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\mem.mem[125][6] ),
    .X(net4198));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\mem.mem[182][3] ),
    .X(net4199));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\mem.mem[119][2] ),
    .X(net4200));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\mem.mem[55][5] ),
    .X(net4201));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\mem.mem[38][4] ),
    .X(net4202));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\mem.mem[102][1] ),
    .X(net4203));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\mem.mem[141][4] ),
    .X(net4204));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\mem.mem[49][5] ),
    .X(net4205));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\mem.mem[195][3] ),
    .X(net4206));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\mem.mem[46][4] ),
    .X(net4207));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\mem.mem[179][0] ),
    .X(net4208));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\mem.mem[142][7] ),
    .X(net4209));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\mem.mem[240][5] ),
    .X(net4210));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\mem.mem[8][2] ),
    .X(net4211));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\mem.mem[168][3] ),
    .X(net4212));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\mem.mem[247][6] ),
    .X(net4213));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\mem.mem[114][6] ),
    .X(net4214));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\mem.mem[22][1] ),
    .X(net4215));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\mem.mem[224][2] ),
    .X(net4216));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\mem.mem[64][1] ),
    .X(net4217));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\mem.mem[114][4] ),
    .X(net4218));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\mem.mem[155][5] ),
    .X(net4219));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\mem.mem[114][2] ),
    .X(net4220));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\mem.mem[87][0] ),
    .X(net4221));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\mem.mem[26][1] ),
    .X(net4222));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\mem.mem[217][0] ),
    .X(net4223));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\mem.mem[67][3] ),
    .X(net4224));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\mem.mem[112][2] ),
    .X(net4225));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\mem.mem[54][4] ),
    .X(net4226));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\mem.mem[123][7] ),
    .X(net4227));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\mem.mem[189][4] ),
    .X(net4228));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\mem.mem[173][0] ),
    .X(net4229));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\mem.mem[167][2] ),
    .X(net4230));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\mem.mem[60][1] ),
    .X(net4231));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\mem.mem[14][7] ),
    .X(net4232));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\mem.mem[43][7] ),
    .X(net4233));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\mem.mem[31][2] ),
    .X(net4234));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\mem.mem[218][2] ),
    .X(net4235));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\mem.mem[71][0] ),
    .X(net4236));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\mem.mem[233][1] ),
    .X(net4237));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\mem.mem[11][5] ),
    .X(net4238));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\mem.mem[226][3] ),
    .X(net4239));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\mem.mem[60][3] ),
    .X(net4240));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\mem.mem[30][6] ),
    .X(net4241));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\mem.mem[85][1] ),
    .X(net4242));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\mem.mem[118][4] ),
    .X(net4243));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\mem.mem[58][5] ),
    .X(net4244));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\mem.mem[2][3] ),
    .X(net4245));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\mem.mem[49][7] ),
    .X(net4246));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\mem.mem[145][5] ),
    .X(net4247));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\mem.mem[118][2] ),
    .X(net4248));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\mem.mem[42][7] ),
    .X(net4249));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\mem.mem[112][7] ),
    .X(net4250));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\mem.mem[37][5] ),
    .X(net4251));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\mem.mem[139][5] ),
    .X(net4252));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\mem.mem[168][0] ),
    .X(net4253));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\mem.mem[118][6] ),
    .X(net4254));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\mem.mem[190][1] ),
    .X(net4255));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\mem.mem[124][6] ),
    .X(net4256));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\mem.mem[99][0] ),
    .X(net4257));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\mem.mem[7][5] ),
    .X(net4258));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\mem.mem[145][2] ),
    .X(net4259));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\mem.mem[51][6] ),
    .X(net4260));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\mem.mem[42][2] ),
    .X(net4261));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\mem.mem[231][6] ),
    .X(net4262));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\mem.mem[141][6] ),
    .X(net4263));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\mem.mem[145][3] ),
    .X(net4264));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\mem.mem[23][7] ),
    .X(net4265));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\mem.mem[45][0] ),
    .X(net4266));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\mem.mem[183][6] ),
    .X(net4267));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\mem.mem[247][2] ),
    .X(net4268));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\mem.mem[34][5] ),
    .X(net4269));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\mem.mem[173][1] ),
    .X(net4270));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\mem.mem[64][3] ),
    .X(net4271));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\mem.mem[107][4] ),
    .X(net4272));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\mem.mem[122][6] ),
    .X(net4273));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\mem.mem[29][7] ),
    .X(net4274));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\mem.mem[141][1] ),
    .X(net4275));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\mem.mem[173][6] ),
    .X(net4276));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\mem.mem[211][7] ),
    .X(net4277));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\mem.mem[29][4] ),
    .X(net4278));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\mem.mem[122][4] ),
    .X(net4279));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\mem.mem[67][7] ),
    .X(net4280));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\mem.mem[240][4] ),
    .X(net4281));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\mem.mem[9][3] ),
    .X(net4282));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\mem.mem[109][6] ),
    .X(net4283));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\mem.mem[182][0] ),
    .X(net4284));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\mem.mem[23][1] ),
    .X(net4285));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\mem.mem[231][5] ),
    .X(net4286));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\mem.mem[240][2] ),
    .X(net4287));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\mem.mem[167][0] ),
    .X(net4288));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\mem.mem[8][5] ),
    .X(net4289));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\mem.mem[154][2] ),
    .X(net4290));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\mem.mem[149][6] ),
    .X(net4291));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\mem.mem[109][2] ),
    .X(net4292));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\mem.mem[188][4] ),
    .X(net4293));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\mem.mem[17][7] ),
    .X(net4294));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\mem.mem[217][3] ),
    .X(net4295));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\mem.mem[8][0] ),
    .X(net4296));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\mem.mem[192][0] ),
    .X(net4297));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\mem.mem[148][0] ),
    .X(net4298));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\mem.mem[61][0] ),
    .X(net4299));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\mem.mem[156][3] ),
    .X(net4300));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\mem.mem[114][1] ),
    .X(net4301));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\mem.mem[135][6] ),
    .X(net4302));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\mem.mem[80][2] ),
    .X(net4303));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\mem.mem[135][1] ),
    .X(net4304));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\mem.mem[174][7] ),
    .X(net4305));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\mem.mem[158][5] ),
    .X(net4306));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\mem.mem[38][3] ),
    .X(net4307));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\mem.mem[74][7] ),
    .X(net4308));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\mem.mem[30][4] ),
    .X(net4309));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\mem.mem[247][1] ),
    .X(net4310));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\mem.mem[195][1] ),
    .X(net4311));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\mem.mem[13][0] ),
    .X(net4312));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\mem.mem[51][4] ),
    .X(net4313));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\mem.mem[180][5] ),
    .X(net4314));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\mem.mem[33][5] ),
    .X(net4315));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\mem.mem[178][4] ),
    .X(net4316));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\mem.mem[139][7] ),
    .X(net4317));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\mem.mem[203][0] ),
    .X(net4318));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\mem.mem[11][4] ),
    .X(net4319));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\mem.mem[155][4] ),
    .X(net4320));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\mem.mem[54][3] ),
    .X(net4321));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\mem.mem[172][3] ),
    .X(net4322));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\mem.mem[45][7] ),
    .X(net4323));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\mem.mem[169][7] ),
    .X(net4324));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\mem.mem[101][0] ),
    .X(net4325));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\mem.mem[247][3] ),
    .X(net4326));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\mem.mem[152][7] ),
    .X(net4327));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\mem.mem[107][6] ),
    .X(net4328));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\mem.mem[92][0] ),
    .X(net4329));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\mem.mem[83][1] ),
    .X(net4330));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\mem.mem[37][4] ),
    .X(net4331));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\mem.mem[108][7] ),
    .X(net4332));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\mem.mem[39][7] ),
    .X(net4333));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\mem.mem[192][3] ),
    .X(net4334));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\mem.mem[6][3] ),
    .X(net4335));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\mem.mem[42][4] ),
    .X(net4336));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\mem.mem[233][7] ),
    .X(net4337));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\mem.mem[194][3] ),
    .X(net4338));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\mem.mem[10][0] ),
    .X(net4339));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\mem.mem[208][6] ),
    .X(net4340));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\mem.mem[235][2] ),
    .X(net4341));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\mem.mem[188][0] ),
    .X(net4342));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\mem.mem[230][3] ),
    .X(net4343));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\mem.mem[211][2] ),
    .X(net4344));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\mem.mem[57][3] ),
    .X(net4345));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\mem.mem[12][1] ),
    .X(net4346));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\mem.mem[91][2] ),
    .X(net4347));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\mem.mem[0][3] ),
    .X(net4348));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\mem.mem[77][0] ),
    .X(net4349));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\mem.mem[7][2] ),
    .X(net4350));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\mem.mem[164][7] ),
    .X(net4351));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\mem.mem[64][4] ),
    .X(net4352));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\mem.mem[6][2] ),
    .X(net4353));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\mem.mem[75][2] ),
    .X(net4354));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\mem.mem[45][2] ),
    .X(net4355));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\mem.mem[108][2] ),
    .X(net4356));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\mem.mem[77][4] ),
    .X(net4357));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\mem.mem[32][1] ),
    .X(net4358));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\mem.mem[165][0] ),
    .X(net4359));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\mem.mem[61][6] ),
    .X(net4360));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\mem.mem[240][6] ),
    .X(net4361));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\mem.mem[124][2] ),
    .X(net4362));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\mem.mem[179][2] ),
    .X(net4363));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\mem.mem[0][1] ),
    .X(net4364));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\mem.mem[53][6] ),
    .X(net4365));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\mem.mem[54][5] ),
    .X(net4366));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\mem.mem[27][0] ),
    .X(net4367));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\mem.mem[234][1] ),
    .X(net4368));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\mem.mem[174][6] ),
    .X(net4369));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\mem.mem[117][7] ),
    .X(net4370));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\mem.mem[190][2] ),
    .X(net4371));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\mem.mem[210][0] ),
    .X(net4372));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\mem.mem[3][3] ),
    .X(net4373));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\mem.mem[115][0] ),
    .X(net4374));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\mem.mem[55][3] ),
    .X(net4375));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\mem.mem[59][1] ),
    .X(net4376));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\mem.mem[202][2] ),
    .X(net4377));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\mem.mem[247][5] ),
    .X(net4378));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\mem.mem[151][3] ),
    .X(net4379));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\mem.mem[233][2] ),
    .X(net4380));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\mem.mem[195][5] ),
    .X(net4381));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\mem.mem[141][5] ),
    .X(net4382));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\mem.mem[173][2] ),
    .X(net4383));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\mem.mem[46][2] ),
    .X(net4384));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\mem.mem[139][1] ),
    .X(net4385));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\mem.mem[1][3] ),
    .X(net4386));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\mem.mem[9][2] ),
    .X(net4387));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\mem.mem[33][6] ),
    .X(net4388));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\mem.mem[60][4] ),
    .X(net4389));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\mem.mem[213][5] ),
    .X(net4390));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\mem.mem[16][3] ),
    .X(net4391));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\mem.mem[80][7] ),
    .X(net4392));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\mem.mem[57][6] ),
    .X(net4393));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\mem.mem[42][5] ),
    .X(net4394));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\mem.mem[231][3] ),
    .X(net4395));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\mem.mem[57][7] ),
    .X(net4396));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\mem.mem[85][6] ),
    .X(net4397));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\mem.mem[42][0] ),
    .X(net4398));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\mem.mem[169][0] ),
    .X(net4399));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\mem.mem[166][5] ),
    .X(net4400));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\mem.mem[106][1] ),
    .X(net4401));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\mem.mem[125][2] ),
    .X(net4402));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\mem.mem[90][4] ),
    .X(net4403));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\mem.mem[199][5] ),
    .X(net4404));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\mem.mem[32][0] ),
    .X(net4405));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\mem.mem[229][2] ),
    .X(net4406));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\mem.mem[178][0] ),
    .X(net4407));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\mem.mem[42][3] ),
    .X(net4408));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\mem.mem[171][3] ),
    .X(net4409));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\mem.mem[152][2] ),
    .X(net4410));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\mem.mem[152][6] ),
    .X(net4411));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\mem.mem[181][3] ),
    .X(net4412));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\mem.mem[18][7] ),
    .X(net4413));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\mem.mem[224][1] ),
    .X(net4414));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\mem.mem[86][0] ),
    .X(net4415));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\mem.mem[182][5] ),
    .X(net4416));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\mem.mem[105][7] ),
    .X(net4417));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\mem.mem[190][0] ),
    .X(net4418));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\mem.mem[83][6] ),
    .X(net4419));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\mem.mem[91][3] ),
    .X(net4420));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\mem.mem[183][2] ),
    .X(net4421));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\mem.mem[115][4] ),
    .X(net4422));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\mem.mem[220][0] ),
    .X(net4423));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\mem.mem[237][2] ),
    .X(net4424));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\mem.mem[217][7] ),
    .X(net4425));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\mem.mem[211][5] ),
    .X(net4426));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\mem.mem[243][7] ),
    .X(net4427));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\mem.mem[217][5] ),
    .X(net4428));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\mem.mem[41][4] ),
    .X(net4429));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\mem.mem[18][2] ),
    .X(net4430));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\mem.mem[11][2] ),
    .X(net4431));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\mem.mem[91][1] ),
    .X(net4432));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\mem.mem[53][1] ),
    .X(net4433));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\mem.mem[213][3] ),
    .X(net4434));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\mem.mem[22][2] ),
    .X(net4435));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\mem.mem[167][6] ),
    .X(net4436));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\mem.mem[122][5] ),
    .X(net4437));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\mem.mem[158][6] ),
    .X(net4438));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\mem.mem[92][1] ),
    .X(net4439));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\mem.mem[58][0] ),
    .X(net4440));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\mem.mem[177][3] ),
    .X(net4441));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\mem.mem[29][3] ),
    .X(net4442));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\mem.mem[9][1] ),
    .X(net4443));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\mem.mem[119][1] ),
    .X(net4444));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\mem.mem[161][1] ),
    .X(net4445));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\mem.mem[169][6] ),
    .X(net4446));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\mem.mem[151][2] ),
    .X(net4447));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\mem.mem[187][5] ),
    .X(net4448));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\mem.mem[54][6] ),
    .X(net4449));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\mem.mem[19][0] ),
    .X(net4450));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\mem.mem[234][5] ),
    .X(net4451));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\mem.mem[67][4] ),
    .X(net4452));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\mem.mem[24][3] ),
    .X(net4453));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\mem.mem[39][3] ),
    .X(net4454));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\mem.mem[119][5] ),
    .X(net4455));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\mem.mem[75][5] ),
    .X(net4456));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\mem.mem[221][3] ),
    .X(net4457));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\mem.mem[162][4] ),
    .X(net4458));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\mem.mem[2][0] ),
    .X(net4459));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\mem.mem[226][1] ),
    .X(net4460));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\mem.mem[27][2] ),
    .X(net4461));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\mem.mem[198][2] ),
    .X(net4462));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\mem.mem[163][4] ),
    .X(net4463));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\mem.mem[237][5] ),
    .X(net4464));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\mem.mem[194][7] ),
    .X(net4465));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\mem.mem[77][3] ),
    .X(net4466));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\mem.mem[35][4] ),
    .X(net4467));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\mem.mem[199][7] ),
    .X(net4468));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\mem.mem[208][0] ),
    .X(net4469));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\mem.mem[237][1] ),
    .X(net4470));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\mem.mem[149][0] ),
    .X(net4471));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\mem.mem[64][7] ),
    .X(net4472));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\mem.mem[24][4] ),
    .X(net4473));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\mem.mem[183][0] ),
    .X(net4474));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\mem.mem[202][0] ),
    .X(net4475));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\mem.mem[57][2] ),
    .X(net4476));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\mem.mem[128][0] ),
    .X(net4477));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\mem.mem[8][1] ),
    .X(net4478));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\mem.mem[167][5] ),
    .X(net4479));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\mem.mem[219][7] ),
    .X(net4480));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\mem.mem[181][6] ),
    .X(net4481));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\mem.mem[61][2] ),
    .X(net4482));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\mem.mem[161][4] ),
    .X(net4483));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\mem.mem[177][5] ),
    .X(net4484));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\mem.mem[154][3] ),
    .X(net4485));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\mem.mem[172][1] ),
    .X(net4486));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\mem.mem[115][3] ),
    .X(net4487));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\mem.mem[219][3] ),
    .X(net4488));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\mem.mem[117][3] ),
    .X(net4489));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\mem.mem[2][1] ),
    .X(net4490));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\mem.mem[197][4] ),
    .X(net4491));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\mem.mem[145][7] ),
    .X(net4492));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\mem.mem[139][0] ),
    .X(net4493));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\mem.mem[1][5] ),
    .X(net4494));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\mem.mem[54][0] ),
    .X(net4495));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\mem.mem[22][0] ),
    .X(net4496));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\mem.mem[216][0] ),
    .X(net4497));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\mem.mem[103][2] ),
    .X(net4498));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\mem.mem[222][2] ),
    .X(net4499));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\mem.mem[60][5] ),
    .X(net4500));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\mem.mem[215][2] ),
    .X(net4501));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\mem.mem[237][0] ),
    .X(net4502));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\mem.mem[119][7] ),
    .X(net4503));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\mem.mem[141][7] ),
    .X(net4504));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\mem.mem[66][4] ),
    .X(net4505));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\mem.mem[145][6] ),
    .X(net4506));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\mem.mem[234][6] ),
    .X(net4507));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\mem.mem[141][2] ),
    .X(net4508));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\mem.mem[48][1] ),
    .X(net4509));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\mem.mem[1][2] ),
    .X(net4510));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\mem.mem[75][7] ),
    .X(net4511));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\mem.mem[19][5] ),
    .X(net4512));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\mem.mem[237][7] ),
    .X(net4513));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\mem.mem[149][3] ),
    .X(net4514));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\mem.mem[213][0] ),
    .X(net4515));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\mem.mem[51][1] ),
    .X(net4516));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\mem.mem[145][0] ),
    .X(net4517));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\mem.mem[2][2] ),
    .X(net4518));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\mem.mem[217][6] ),
    .X(net4519));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\mem.mem[14][5] ),
    .X(net4520));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\mem.mem[234][3] ),
    .X(net4521));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\mem.mem[233][6] ),
    .X(net4522));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\mem.mem[208][1] ),
    .X(net4523));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\mem.mem[85][4] ),
    .X(net4524));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\mem.mem[16][2] ),
    .X(net4525));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\mem.mem[58][7] ),
    .X(net4526));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\mem.mem[58][1] ),
    .X(net4527));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\mem.mem[215][1] ),
    .X(net4528));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\mem.mem[75][6] ),
    .X(net4529));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\mem.mem[112][5] ),
    .X(net4530));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\mem.mem[37][2] ),
    .X(net4531));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\mem.mem[101][5] ),
    .X(net4532));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\mem.mem[49][0] ),
    .X(net4533));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\mem.mem[235][5] ),
    .X(net4534));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\mem.mem[66][3] ),
    .X(net4535));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\mem.mem[119][0] ),
    .X(net4536));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\mem.mem[9][7] ),
    .X(net4537));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\mem.mem[150][3] ),
    .X(net4538));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\mem.mem[115][1] ),
    .X(net4539));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\mem.mem[229][6] ),
    .X(net4540));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\mem.mem[147][3] ),
    .X(net4541));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\mem.mem[103][6] ),
    .X(net4542));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\mem.mem[164][6] ),
    .X(net4543));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\mem.mem[12][0] ),
    .X(net4544));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\mem.mem[99][4] ),
    .X(net4545));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\mem.mem[36][3] ),
    .X(net4546));
 sg13g2_dlygate4sd3_1 hold1417 (.A(\mem.mem[85][7] ),
    .X(net4547));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\mem.mem[230][0] ),
    .X(net4548));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\mem.mem[108][0] ),
    .X(net4549));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\mem.mem[125][4] ),
    .X(net4550));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\mem.mem[33][3] ),
    .X(net4551));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\mem.mem[32][7] ),
    .X(net4552));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\mem.mem[173][7] ),
    .X(net4553));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\mem.mem[183][3] ),
    .X(net4554));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\mem.mem[55][0] ),
    .X(net4555));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\mem.mem[35][3] ),
    .X(net4556));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\mem.mem[165][6] ),
    .X(net4557));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\mem.mem[61][1] ),
    .X(net4558));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\mem.mem[157][7] ),
    .X(net4559));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\mem.mem[158][2] ),
    .X(net4560));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\mem.mem[55][4] ),
    .X(net4561));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\mem.mem[125][1] ),
    .X(net4562));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\mem.mem[77][2] ),
    .X(net4563));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\mem.mem[181][0] ),
    .X(net4564));
 sg13g2_dlygate4sd3_1 hold1435 (.A(\mem.mem[153][7] ),
    .X(net4565));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\mem.mem[34][4] ),
    .X(net4566));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\mem.mem[242][7] ),
    .X(net4567));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\mem.mem[74][0] ),
    .X(net4568));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\mem.mem[87][4] ),
    .X(net4569));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\mem.mem[156][0] ),
    .X(net4570));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\mem.mem[80][5] ),
    .X(net4571));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\mem.mem[45][4] ),
    .X(net4572));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\mem.mem[210][6] ),
    .X(net4573));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\mem.mem[234][0] ),
    .X(net4574));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\mem.mem[186][7] ),
    .X(net4575));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\mem.mem[247][4] ),
    .X(net4576));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\mem.mem[169][1] ),
    .X(net4577));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\mem.mem[19][3] ),
    .X(net4578));
 sg13g2_dlygate4sd3_1 hold1449 (.A(\mem.mem[189][6] ),
    .X(net4579));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\mem.mem[128][2] ),
    .X(net4580));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\mem.uo_out[3] ),
    .X(net4581));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\mem.mem[217][2] ),
    .X(net4582));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\mem.mem[112][3] ),
    .X(net4583));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\mem.mem[83][2] ),
    .X(net4584));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\mem.mem[35][1] ),
    .X(net4585));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\mem.mem[30][5] ),
    .X(net4586));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\mem.mem[87][6] ),
    .X(net4587));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\mem.mem[34][2] ),
    .X(net4588));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\mem.mem[149][4] ),
    .X(net4589));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\mem.mem[55][2] ),
    .X(net4590));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\mem.mem[211][4] ),
    .X(net4591));
 sg13g2_dlygate4sd3_1 hold1462 (.A(\mem.mem[198][3] ),
    .X(net4592));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\mem.mem[99][2] ),
    .X(net4593));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\mem.mem[145][4] ),
    .X(net4594));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\mem.mem[35][7] ),
    .X(net4595));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\mem.mem[174][0] ),
    .X(net4596));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\mem.mem[229][0] ),
    .X(net4597));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\mem.mem[36][0] ),
    .X(net4598));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\mem.mem[3][1] ),
    .X(net4599));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\mem.mem[157][3] ),
    .X(net4600));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\mem.mem[170][6] ),
    .X(net4601));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\mem.mem[96][0] ),
    .X(net4602));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\mem.mem[164][4] ),
    .X(net4603));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\mem.mem[190][3] ),
    .X(net4604));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\mem.mem[29][0] ),
    .X(net4605));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\mem.mem[10][7] ),
    .X(net4606));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\mem.mem[243][6] ),
    .X(net4607));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\mem.mem[231][2] ),
    .X(net4608));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\mem.mem[195][2] ),
    .X(net4609));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\mem.mem[146][0] ),
    .X(net4610));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\mem.mem[50][0] ),
    .X(net4611));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\mem.mem[23][4] ),
    .X(net4612));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\mem.mem[100][7] ),
    .X(net4613));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\mem.mem[202][4] ),
    .X(net4614));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\mem.mem[161][0] ),
    .X(net4615));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\mem.mem[147][2] ),
    .X(net4616));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\mem.mem[109][5] ),
    .X(net4617));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\mem.mem[77][5] ),
    .X(net4618));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\mem.mem[106][4] ),
    .X(net4619));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\mem.mem[227][1] ),
    .X(net4620));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\mem.mem[230][6] ),
    .X(net4621));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\mem.mem[49][2] ),
    .X(net4622));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\mem.mem[43][2] ),
    .X(net4623));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\mem.mem[39][5] ),
    .X(net4624));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\mem.mem[168][7] ),
    .X(net4625));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\mem.mem[26][4] ),
    .X(net4626));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\mem.mem[53][7] ),
    .X(net4627));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\mem.mem[126][2] ),
    .X(net4628));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\mem.mem[10][2] ),
    .X(net4629));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\mem.mem[142][2] ),
    .X(net4630));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\mem.mem[186][2] ),
    .X(net4631));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\mem.mem[103][7] ),
    .X(net4632));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\mem.mem[102][2] ),
    .X(net4633));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\mem.mem[119][4] ),
    .X(net4634));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\mem.mem[126][1] ),
    .X(net4635));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\mem.mem[87][3] ),
    .X(net4636));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\mem.mem[226][6] ),
    .X(net4637));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\mem.mem[96][2] ),
    .X(net4638));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\mem.mem[174][4] ),
    .X(net4639));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\mem.mem[238][6] ),
    .X(net4640));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\mem.mem[109][3] ),
    .X(net4641));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\mem.mem[141][0] ),
    .X(net4642));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\mem.mem[153][4] ),
    .X(net4643));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\mem.mem[202][5] ),
    .X(net4644));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\mem.mem[115][5] ),
    .X(net4645));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\mem.mem[75][3] ),
    .X(net4646));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\mem.mem[151][5] ),
    .X(net4647));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\mem.mem[62][3] ),
    .X(net4648));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\mem.mem[141][3] ),
    .X(net4649));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\mem.mem[71][2] ),
    .X(net4650));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\mem.mem[183][5] ),
    .X(net4651));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\mem.mem[53][4] ),
    .X(net4652));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\mem.mem[233][3] ),
    .X(net4653));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\mem.mem[26][0] ),
    .X(net4654));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\mem.mem[168][2] ),
    .X(net4655));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\mem.mem[92][2] ),
    .X(net4656));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\mem.mem[218][6] ),
    .X(net4657));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\mem.mem[221][4] ),
    .X(net4658));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\mem.mem[199][6] ),
    .X(net4659));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\mem.mem[180][1] ),
    .X(net4660));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\mem.mem[82][5] ),
    .X(net4661));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\mem.mem[117][4] ),
    .X(net4662));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\mem.mem[178][1] ),
    .X(net4663));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\mem.mem[117][1] ),
    .X(net4664));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\mem.mem[48][0] ),
    .X(net4665));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\mem.mem[165][3] ),
    .X(net4666));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\mem.mem[197][3] ),
    .X(net4667));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\mem.mem[66][7] ),
    .X(net4668));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\mem.mem[107][7] ),
    .X(net4669));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\mem.mem[146][2] ),
    .X(net4670));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\mem.mem[102][5] ),
    .X(net4671));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\mem.mem[128][4] ),
    .X(net4672));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\mem.mem[197][1] ),
    .X(net4673));
 sg13g2_dlygate4sd3_1 hold1544 (.A(\mem.mem[126][7] ),
    .X(net4674));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\mem.mem[1][1] ),
    .X(net4675));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\mem.mem[179][3] ),
    .X(net4676));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\mem.mem[162][1] ),
    .X(net4677));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\mem.mem[109][1] ),
    .X(net4678));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\mem.mem[41][0] ),
    .X(net4679));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\mem.mem[35][0] ),
    .X(net4680));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\mem.mem[58][2] ),
    .X(net4681));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\mem.mem[214][7] ),
    .X(net4682));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\mem.mem[14][3] ),
    .X(net4683));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\mem.mem[19][2] ),
    .X(net4684));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\mem.mem[26][3] ),
    .X(net4685));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\mem.mem[162][0] ),
    .X(net4686));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\mem.mem[43][1] ),
    .X(net4687));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\mem.mem[153][5] ),
    .X(net4688));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\mem.mem[224][7] ),
    .X(net4689));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\mem.mem[185][7] ),
    .X(net4690));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\mem.mem[13][3] ),
    .X(net4691));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\mem.mem[117][2] ),
    .X(net4692));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\mem.mem[148][5] ),
    .X(net4693));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\mem.mem[202][6] ),
    .X(net4694));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\mem.mem[197][7] ),
    .X(net4695));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\mem.mem[146][4] ),
    .X(net4696));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\mem.mem[71][1] ),
    .X(net4697));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\mem.mem[118][7] ),
    .X(net4698));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\mem.mem[9][4] ),
    .X(net4699));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\mem.mem[171][1] ),
    .X(net4700));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\mem.mem[108][5] ),
    .X(net4701));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\mem.mem[153][6] ),
    .X(net4702));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\mem.mem[171][0] ),
    .X(net4703));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\mem.mem[128][7] ),
    .X(net4704));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\mem.mem[105][4] ),
    .X(net4705));
 sg13g2_dlygate4sd3_1 hold1576 (.A(\mem.mem[85][2] ),
    .X(net4706));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\mem.mem[166][7] ),
    .X(net4707));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\mem.mem[119][6] ),
    .X(net4708));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\mem.mem[29][5] ),
    .X(net4709));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\mem.mem[242][5] ),
    .X(net4710));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\mem.mem[117][0] ),
    .X(net4711));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\mem.mem[240][1] ),
    .X(net4712));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\mem.mem[124][4] ),
    .X(net4713));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\mem.mem[8][7] ),
    .X(net4714));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\mem.mem[236][2] ),
    .X(net4715));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\mem.mem[179][1] ),
    .X(net4716));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\mem.mem[236][1] ),
    .X(net4717));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\mem.mem[118][0] ),
    .X(net4718));
 sg13g2_dlygate4sd3_1 hold1589 (.A(\mem.mem[165][1] ),
    .X(net4719));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\mem.mem[170][0] ),
    .X(net4720));
 sg13g2_dlygate4sd3_1 hold1591 (.A(\mem.mem[126][3] ),
    .X(net4721));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\mem.mem[171][5] ),
    .X(net4722));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\mem.mem[50][4] ),
    .X(net4723));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\mem.mem[214][6] ),
    .X(net4724));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\mem.mem[154][5] ),
    .X(net4725));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\mem.mem[26][7] ),
    .X(net4726));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\mem.mem[236][3] ),
    .X(net4727));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\mem.mem[118][3] ),
    .X(net4728));
 sg13g2_dlygate4sd3_1 hold1599 (.A(\mem.mem[25][1] ),
    .X(net4729));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\mem.mem[27][3] ),
    .X(net4730));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\mem.mem[23][3] ),
    .X(net4731));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\mem.mem[227][3] ),
    .X(net4732));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\mem.mem[55][1] ),
    .X(net4733));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\mem.mem[13][7] ),
    .X(net4734));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\mem.mem[31][1] ),
    .X(net4735));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\mem.mem[214][1] ),
    .X(net4736));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\mem.mem[87][7] ),
    .X(net4737));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\mem.mem[204][7] ),
    .X(net4738));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\mem.mem[32][2] ),
    .X(net4739));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\mem.mem[242][6] ),
    .X(net4740));
 sg13g2_dlygate4sd3_1 hold1611 (.A(\mem.mem[41][2] ),
    .X(net4741));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\mem.mem[189][0] ),
    .X(net4742));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\mem.mem[233][4] ),
    .X(net4743));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\mem.mem[211][6] ),
    .X(net4744));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\mem.mem[87][2] ),
    .X(net4745));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\mem.mem[156][6] ),
    .X(net4746));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\mem.mem[146][1] ),
    .X(net4747));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\mem.mem[105][3] ),
    .X(net4748));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\mem.mem[115][2] ),
    .X(net4749));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\mem.mem[243][1] ),
    .X(net4750));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\mem.mem[199][4] ),
    .X(net4751));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\mem.mem[53][5] ),
    .X(net4752));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\mem.mem[32][3] ),
    .X(net4753));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\mem.mem[34][1] ),
    .X(net4754));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\mem.mem[5][1] ),
    .X(net4755));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\mem.mem[126][4] ),
    .X(net4756));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\mem.mem[222][5] ),
    .X(net4757));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\mem.mem[169][3] ),
    .X(net4758));
 sg13g2_dlygate4sd3_1 hold1629 (.A(\mem.mem[195][6] ),
    .X(net4759));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\mem.mem[50][1] ),
    .X(net4760));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\mem.mem[57][5] ),
    .X(net4761));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\mem.mem[105][5] ),
    .X(net4762));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\mem.mem[147][1] ),
    .X(net4763));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\mem.mem[100][2] ),
    .X(net4764));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\mem.mem[10][1] ),
    .X(net4765));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\mem.mem[18][0] ),
    .X(net4766));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\mem.mem[86][3] ),
    .X(net4767));
 sg13g2_dlygate4sd3_1 hold1638 (.A(\mem.mem[186][5] ),
    .X(net4768));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\mem.mem[77][7] ),
    .X(net4769));
 sg13g2_dlygate4sd3_1 hold1640 (.A(\mem.mem[19][1] ),
    .X(net4770));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\mem.mem[167][1] ),
    .X(net4771));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\mem.mem[135][4] ),
    .X(net4772));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\mem.mem[185][6] ),
    .X(net4773));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\mem.mem[173][3] ),
    .X(net4774));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\mem.mem[50][5] ),
    .X(net4775));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\mem.mem[178][5] ),
    .X(net4776));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\mem.mem[219][1] ),
    .X(net4777));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\mem.mem[155][0] ),
    .X(net4778));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\mem.mem[59][4] ),
    .X(net4779));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\mem.mem[49][6] ),
    .X(net4780));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\mem.mem[11][6] ),
    .X(net4781));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\mem.mem[203][6] ),
    .X(net4782));
 sg13g2_dlygate4sd3_1 hold1653 (.A(\mem.mem[37][3] ),
    .X(net4783));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\mem.mem[85][0] ),
    .X(net4784));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\mem.mem[5][2] ),
    .X(net4785));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\mem.mem[126][5] ),
    .X(net4786));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\mem.mem[215][7] ),
    .X(net4787));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\mem.mem[154][6] ),
    .X(net4788));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\mem.mem[101][3] ),
    .X(net4789));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\mem.mem[75][1] ),
    .X(net4790));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\mem.mem[105][6] ),
    .X(net4791));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\mem.mem[34][7] ),
    .X(net4792));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\mem.mem[10][5] ),
    .X(net4793));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\mem.mem[210][1] ),
    .X(net4794));
 sg13g2_dlygate4sd3_1 hold1665 (.A(\mem.mem[189][1] ),
    .X(net4795));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\mem.mem[148][4] ),
    .X(net4796));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\mem.mem[165][7] ),
    .X(net4797));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\mem.mem[214][3] ),
    .X(net4798));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\mem.mem[125][3] ),
    .X(net4799));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\mem.mem[17][0] ),
    .X(net4800));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\mem.mem[153][1] ),
    .X(net4801));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\mem.mem[20][0] ),
    .X(net4802));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\mem.mem[161][3] ),
    .X(net4803));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\mem.mem[100][1] ),
    .X(net4804));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\mem.mem[154][0] ),
    .X(net4805));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\mem.mem[180][3] ),
    .X(net4806));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\mem.mem[123][3] ),
    .X(net4807));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\mem.mem[208][3] ),
    .X(net4808));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\mem.mem[1][0] ),
    .X(net4809));
 sg13g2_dlygate4sd3_1 hold1680 (.A(\mem.mem[33][1] ),
    .X(net4810));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\mem.mem[101][1] ),
    .X(net4811));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\mem.mem[10][3] ),
    .X(net4812));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\mem.mem[67][6] ),
    .X(net4813));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\mem.mem[87][1] ),
    .X(net4814));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\mem.mem[14][2] ),
    .X(net4815));
 sg13g2_dlygate4sd3_1 hold1686 (.A(\mem.mem[203][7] ),
    .X(net4816));
 sg13g2_dlygate4sd3_1 hold1687 (.A(\mem.mem[169][5] ),
    .X(net4817));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\mem.mem[198][1] ),
    .X(net4818));
 sg13g2_dlygate4sd3_1 hold1689 (.A(\mem.mem[38][6] ),
    .X(net4819));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\mem.mem[12][3] ),
    .X(net4820));
 sg13g2_dlygate4sd3_1 hold1691 (.A(\mem.mem[109][7] ),
    .X(net4821));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\mem.mem[128][1] ),
    .X(net4822));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\mem.mem[5][6] ),
    .X(net4823));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\mem.mem[185][1] ),
    .X(net4824));
 sg13g2_dlygate4sd3_1 hold1695 (.A(\mem.mem[157][1] ),
    .X(net4825));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\mem.mem[51][7] ),
    .X(net4826));
 sg13g2_dlygate4sd3_1 hold1697 (.A(\mem.mem[166][3] ),
    .X(net4827));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\mem.mem[146][3] ),
    .X(net4828));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\mem.mem[128][3] ),
    .X(net4829));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\mem.mem[227][4] ),
    .X(net4830));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\mem.mem[47][4] ),
    .X(net4831));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\mem.mem[47][7] ),
    .X(net4832));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\mem.mem[29][2] ),
    .X(net4833));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\mem.mem[197][5] ),
    .X(net4834));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\mem.mem[151][0] ),
    .X(net4835));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\mem.mem[75][0] ),
    .X(net4836));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\mem.mem[182][7] ),
    .X(net4837));
 sg13g2_dlygate4sd3_1 hold1708 (.A(\mem.mem[46][3] ),
    .X(net4838));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\mem.mem[35][5] ),
    .X(net4839));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\mem.mem[91][6] ),
    .X(net4840));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\mem.mem[166][2] ),
    .X(net4841));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\mem.mem[71][6] ),
    .X(net4842));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\mem.mem[64][2] ),
    .X(net4843));
 sg13g2_dlygate4sd3_1 hold1714 (.A(\mem.mem[31][5] ),
    .X(net4844));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\mem.mem[168][1] ),
    .X(net4845));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\mem.mem[177][1] ),
    .X(net4846));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\mem.mem[42][1] ),
    .X(net4847));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\mem.mem[156][1] ),
    .X(net4848));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\mem.mem[235][6] ),
    .X(net4849));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\mem_A[2] ),
    .X(net4850));
 sg13g2_dlygate4sd3_1 hold1721 (.A(_00648_),
    .X(net4851));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\mem.mem[169][4] ),
    .X(net4852));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\mem.mem[25][2] ),
    .X(net4853));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\mem.mem[2][7] ),
    .X(net4854));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\mem.mem[50][6] ),
    .X(net4855));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\mem.mem[204][3] ),
    .X(net4856));
 sg13g2_dlygate4sd3_1 hold1727 (.A(\mem.mem[90][2] ),
    .X(net4857));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\mem.mem[45][1] ),
    .X(net4858));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\mem.mem[20][1] ),
    .X(net4859));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\mem.mem[75][4] ),
    .X(net4860));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\mem.mem[83][3] ),
    .X(net4861));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\mem.mem[162][3] ),
    .X(net4862));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\mem.mem[164][0] ),
    .X(net4863));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\mem.mem[213][4] ),
    .X(net4864));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\mem.mem[8][3] ),
    .X(net4865));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\mem.mem[215][5] ),
    .X(net4866));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\mem.mem[66][0] ),
    .X(net4867));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\mem.mem[152][5] ),
    .X(net4868));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\mem.mem[219][0] ),
    .X(net4869));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\mem.mem[34][6] ),
    .X(net4870));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\mem.mem[211][3] ),
    .X(net4871));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\mem.mem[51][0] ),
    .X(net4872));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\mem.mem[139][4] ),
    .X(net4873));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\mem.mem[51][3] ),
    .X(net4874));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\mem.mem[195][0] ),
    .X(net4875));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\mem.mem[203][3] ),
    .X(net4876));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\mem.mem[45][3] ),
    .X(net4877));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\mem.mem[23][5] ),
    .X(net4878));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\mem.mem[99][7] ),
    .X(net4879));
 sg13g2_dlygate4sd3_1 hold1750 (.A(\mem.mem[0][2] ),
    .X(net4880));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\mem.mem[3][4] ),
    .X(net4881));
 sg13g2_dlygate4sd3_1 hold1752 (.A(\mem.mem[187][1] ),
    .X(net4882));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\mem.mem[231][4] ),
    .X(net4883));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\mem.mem[106][2] ),
    .X(net4884));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\mem.mem[13][4] ),
    .X(net4885));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\mem.mem[9][5] ),
    .X(net4886));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\mem.mem[83][7] ),
    .X(net4887));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\mem.mem[247][0] ),
    .X(net4888));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\mem.mem[21][4] ),
    .X(net4889));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\mem.mem[82][6] ),
    .X(net4890));
 sg13g2_dlygate4sd3_1 hold1761 (.A(\mem.mem[26][5] ),
    .X(net4891));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\mem.mem[87][5] ),
    .X(net4892));
 sg13g2_dlygate4sd3_1 hold1763 (.A(\mem.mem[67][5] ),
    .X(net4893));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\mem.mem[67][2] ),
    .X(net4894));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\mem.mem[122][3] ),
    .X(net4895));
 sg13g2_dlygate4sd3_1 hold1766 (.A(\mem.mem[17][5] ),
    .X(net4896));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\mem.mem[152][0] ),
    .X(net4897));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\mem.mem[41][3] ),
    .X(net4898));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\mem.mem[226][2] ),
    .X(net4899));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\mem.mem[6][1] ),
    .X(net4900));
 sg13g2_dlygate4sd3_1 hold1771 (.A(\mem.mem[24][5] ),
    .X(net4901));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\mem.mem[6][7] ),
    .X(net4902));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\mem.mem[163][6] ),
    .X(net4903));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\mem.mem[203][2] ),
    .X(net4904));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\mem.mem[118][5] ),
    .X(net4905));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\mem.mem[41][6] ),
    .X(net4906));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\mem.mem[163][3] ),
    .X(net4907));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\mem.mem[74][2] ),
    .X(net4908));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\mem.mem[85][3] ),
    .X(net4909));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\mem.mem[123][1] ),
    .X(net4910));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\mem.mem[6][0] ),
    .X(net4911));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\mem.mem[61][3] ),
    .X(net4912));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\mem.mem[199][0] ),
    .X(net4913));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\mem.mem[242][2] ),
    .X(net4914));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\mem.mem[115][6] ),
    .X(net4915));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\mem.mem[12][2] ),
    .X(net4916));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\mem.mem[58][4] ),
    .X(net4917));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\mem.mem[21][2] ),
    .X(net4918));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\mem.mem[47][2] ),
    .X(net4919));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\mem.mem[238][2] ),
    .X(net4920));
 sg13g2_dlygate4sd3_1 hold1791 (.A(\mem.mem[188][1] ),
    .X(net4921));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\mem.mem[217][1] ),
    .X(net4922));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\mem.mem[10][4] ),
    .X(net4923));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\mem.mem[171][4] ),
    .X(net4924));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\mem.mem[185][3] ),
    .X(net4925));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\mem.mem[243][5] ),
    .X(net4926));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\mem.mem[123][0] ),
    .X(net4927));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\mem.mem[242][1] ),
    .X(net4928));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\mem.mem[17][2] ),
    .X(net4929));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\mem.mem[58][6] ),
    .X(net4930));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\mem.mem[220][1] ),
    .X(net4931));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\mem.mem[240][7] ),
    .X(net4932));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\mem.mem[24][0] ),
    .X(net4933));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\mem.mem[91][7] ),
    .X(net4934));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\mem.mem[27][7] ),
    .X(net4935));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\mem.mem[220][6] ),
    .X(net4936));
 sg13g2_dlygate4sd3_1 hold1807 (.A(\mem.mem[5][3] ),
    .X(net4937));
 sg13g2_dlygate4sd3_1 hold1808 (.A(\mem.mem[4][4] ),
    .X(net4938));
 sg13g2_dlygate4sd3_1 hold1809 (.A(\mem.mem[47][5] ),
    .X(net4939));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\mem.mem[203][4] ),
    .X(net4940));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\mem.mem[243][0] ),
    .X(net4941));
 sg13g2_dlygate4sd3_1 hold1812 (.A(\mem.mem[171][2] ),
    .X(net4942));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\mem.mem[23][2] ),
    .X(net4943));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\mem.mem[74][4] ),
    .X(net4944));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\mem.mem[178][7] ),
    .X(net4945));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\mem.mem[119][3] ),
    .X(net4946));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\mem.mem[221][6] ),
    .X(net4947));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\mem.mem[71][5] ),
    .X(net4948));
 sg13g2_dlygate4sd3_1 hold1819 (.A(\mem.mem[46][1] ),
    .X(net4949));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\mem.mem[86][2] ),
    .X(net4950));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\mem.mem[5][5] ),
    .X(net4951));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\mem.mem[170][2] ),
    .X(net4952));
 sg13g2_dlygate4sd3_1 hold1823 (.A(\mem.mem[167][3] ),
    .X(net4953));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\mem.mem[1][4] ),
    .X(net4954));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\mem.mem[185][4] ),
    .X(net4955));
 sg13g2_dlygate4sd3_1 hold1826 (.A(\mem.mem[213][7] ),
    .X(net4956));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\mem.mem[147][6] ),
    .X(net4957));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\mem.mem[19][4] ),
    .X(net4958));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\mem.mem[26][6] ),
    .X(net4959));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\mem.mem[80][1] ),
    .X(net4960));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\mem.mem[195][7] ),
    .X(net4961));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\mem.mem[155][1] ),
    .X(net4962));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\mem.mem[135][5] ),
    .X(net4963));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\mem.mem[27][1] ),
    .X(net4964));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\mem.mem[101][2] ),
    .X(net4965));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\mem.mem[106][6] ),
    .X(net4966));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\mem.mem[125][7] ),
    .X(net4967));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\mem.mem[41][7] ),
    .X(net4968));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\mem.mem[36][2] ),
    .X(net4969));
 sg13g2_dlygate4sd3_1 hold1840 (.A(\mem.mem[99][1] ),
    .X(net4970));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\mem.mem[123][4] ),
    .X(net4971));
 sg13g2_dlygate4sd3_1 hold1842 (.A(\mem.mem[218][4] ),
    .X(net4972));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\mem.mem[213][1] ),
    .X(net4973));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\mem.mem[235][1] ),
    .X(net4974));
 sg13g2_dlygate4sd3_1 hold1845 (.A(\mem.mem[242][4] ),
    .X(net4975));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\mem.mem[216][4] ),
    .X(net4976));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\mem.mem[43][3] ),
    .X(net4977));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\mem.mem[39][4] ),
    .X(net4978));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\mem.mem[169][2] ),
    .X(net4979));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\mem.mem[91][0] ),
    .X(net4980));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\mem.mem[233][5] ),
    .X(net4981));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\mem.mem[33][7] ),
    .X(net4982));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\mem.mem[117][5] ),
    .X(net4983));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\mem.mem[189][5] ),
    .X(net4984));
 sg13g2_dlygate4sd3_1 hold1855 (.A(\mem.mem[157][4] ),
    .X(net4985));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\mem.mem[31][7] ),
    .X(net4986));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\mem.mem[154][7] ),
    .X(net4987));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\mem.mem[74][6] ),
    .X(net4988));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\mem.mem[110][1] ),
    .X(net4989));
 sg13g2_dlygate4sd3_1 hold1860 (.A(\mem.mem[101][4] ),
    .X(net4990));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\mem.mem[189][7] ),
    .X(net4991));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\mem.mem[112][1] ),
    .X(net4992));
 sg13g2_dlygate4sd3_1 hold1863 (.A(\mem.mem[11][7] ),
    .X(net4993));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\mem.mem[13][6] ),
    .X(net4994));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\mem.mem[24][1] ),
    .X(net4995));
 sg13g2_dlygate4sd3_1 hold1866 (.A(\mem.mem[45][5] ),
    .X(net4996));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\mem.mem[156][7] ),
    .X(net4997));
 sg13g2_dlygate4sd3_1 hold1868 (.A(\mem.mem[229][5] ),
    .X(net4998));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\mem.mem[61][5] ),
    .X(net4999));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\mem.mem[188][5] ),
    .X(net5000));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\mem.mem[229][1] ),
    .X(net5001));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\mem.mem[11][1] ),
    .X(net5002));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\mem.mem[71][4] ),
    .X(net5003));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\mem.mem[66][2] ),
    .X(net5004));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\mem.mem[3][6] ),
    .X(net5005));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\mem.mem[173][5] ),
    .X(net5006));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\mem.mem[5][7] ),
    .X(net5007));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\mem.mem[24][7] ),
    .X(net5008));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\mem.mem[51][2] ),
    .X(net5009));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\mem.mem[102][6] ),
    .X(net5010));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\mem.mem[177][2] ),
    .X(net5011));
 sg13g2_dlygate4sd3_1 hold1882 (.A(\mem.mem[221][5] ),
    .X(net5012));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\mem.mem[34][3] ),
    .X(net5013));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\mem.mem[90][1] ),
    .X(net5014));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\mem.mem[178][6] ),
    .X(net5015));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\mem.mem[3][7] ),
    .X(net5016));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\mem.mem[37][0] ),
    .X(net5017));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\mem.mem[226][7] ),
    .X(net5018));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\mem.mem[187][4] ),
    .X(net5019));
 sg13g2_dlygate4sd3_1 hold1890 (.A(\mem.mem[82][2] ),
    .X(net5020));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\mem.mem[150][2] ),
    .X(net5021));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\mem.mem[7][3] ),
    .X(net5022));
 sg13g2_dlygate4sd3_1 hold1893 (.A(\mem.mem[103][4] ),
    .X(net5023));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\mem.mem[11][0] ),
    .X(net5024));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\mem.mem[47][0] ),
    .X(net5025));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\mem.mem[240][3] ),
    .X(net5026));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\mem.mem[21][6] ),
    .X(net5027));
 sg13g2_dlygate4sd3_1 hold1898 (.A(\mem.mem[163][2] ),
    .X(net5028));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\mem.mem[227][0] ),
    .X(net5029));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\mem.mem[91][5] ),
    .X(net5030));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\mem.mem[147][4] ),
    .X(net5031));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\mem.mem[222][6] ),
    .X(net5032));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\mem.mem[173][4] ),
    .X(net5033));
 sg13g2_dlygate4sd3_1 hold1904 (.A(\mem.mem[214][2] ),
    .X(net5034));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\mem.mem[165][2] ),
    .X(net5035));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\mem.mem[59][5] ),
    .X(net5036));
 sg13g2_dlygate4sd3_1 hold1907 (.A(\mem.mem[71][3] ),
    .X(net5037));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\mem.mem[49][3] ),
    .X(net5038));
 sg13g2_dlygate4sd3_1 hold1909 (.A(\mem.mem[59][7] ),
    .X(net5039));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\mem.uo_out[1] ),
    .X(net5040));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\mem.mem[227][5] ),
    .X(net5041));
 sg13g2_dlygate4sd3_1 hold1912 (.A(\mem.mem[37][7] ),
    .X(net5042));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\mem.mem[186][6] ),
    .X(net5043));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\mem.mem[19][6] ),
    .X(net5044));
 sg13g2_dlygate4sd3_1 hold1915 (.A(\mem.mem[82][4] ),
    .X(net5045));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\mem.mem[107][5] ),
    .X(net5046));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\mem.mem[215][3] ),
    .X(net5047));
 sg13g2_dlygate4sd3_1 hold1918 (.A(\mem.mem[236][7] ),
    .X(net5048));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\mem.mem[30][1] ),
    .X(net5049));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\mem.mem[181][4] ),
    .X(net5050));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\mem.mem[184][3] ),
    .X(net5051));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\mem.mem[91][4] ),
    .X(net5052));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\mem.mem[66][1] ),
    .X(net5053));
 sg13g2_dlygate4sd3_1 hold1924 (.A(\mem.mem[215][4] ),
    .X(net5054));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\mem.mem[194][6] ),
    .X(net5055));
 sg13g2_dlygate4sd3_1 hold1926 (.A(\mem.mem[190][4] ),
    .X(net5056));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\mem.mem[48][7] ),
    .X(net5057));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\mem.mem[124][7] ),
    .X(net5058));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\mem.mem[30][0] ),
    .X(net5059));
 sg13g2_dlygate4sd3_1 hold1930 (.A(\mem.mem[214][0] ),
    .X(net5060));
 sg13g2_dlygate4sd3_1 hold1931 (.A(\mem.mem[147][7] ),
    .X(net5061));
 sg13g2_dlygate4sd3_1 hold1932 (.A(\mem.mem[39][1] ),
    .X(net5062));
 sg13g2_dlygate4sd3_1 hold1933 (.A(\mem.mem[17][3] ),
    .X(net5063));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\mem.mem[229][3] ),
    .X(net5064));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\mem.mem[179][6] ),
    .X(net5065));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\mem.mem[83][0] ),
    .X(net5066));
 sg13g2_dlygate4sd3_1 hold1937 (.A(\mem.mem[179][4] ),
    .X(net5067));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\mem.mem[45][6] ),
    .X(net5068));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\mem.mem[146][5] ),
    .X(net5069));
 sg13g2_dlygate4sd3_1 hold1940 (.A(\mem.mem[237][6] ),
    .X(net5070));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\mem.mem[62][1] ),
    .X(net5071));
 sg13g2_dlygate4sd3_1 hold1942 (.A(\mem.mem[153][3] ),
    .X(net5072));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\mem.mem[189][2] ),
    .X(net5073));
 sg13g2_dlygate4sd3_1 hold1944 (.A(\mem.mem[217][4] ),
    .X(net5074));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\mem.mem[3][0] ),
    .X(net5075));
 sg13g2_dlygate4sd3_1 hold1946 (.A(\mem.mem[107][2] ),
    .X(net5076));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\mem.mem[227][7] ),
    .X(net5077));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\mem.mem[124][3] ),
    .X(net5078));
 sg13g2_dlygate4sd3_1 hold1949 (.A(\mem.mem[187][2] ),
    .X(net5079));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\mem.mem[3][2] ),
    .X(net5080));
 sg13g2_dlygate4sd3_1 hold1951 (.A(\mem.mem[122][0] ),
    .X(net5081));
 sg13g2_dlygate4sd3_1 hold1952 (.A(\mem.mem[30][3] ),
    .X(net5082));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\mem.mem[168][5] ),
    .X(net5083));
 sg13g2_dlygate4sd3_1 hold1954 (.A(\mem.mem[181][2] ),
    .X(net5084));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\mem.mem[80][4] ),
    .X(net5085));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\mem.mem[139][3] ),
    .X(net5086));
 sg13g2_dlygate4sd3_1 hold1957 (.A(\mem.mem[51][5] ),
    .X(net5087));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\mem.mem[168][6] ),
    .X(net5088));
 sg13g2_dlygate4sd3_1 hold1959 (.A(\mem.mem[161][6] ),
    .X(net5089));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\mem.mem[59][3] ),
    .X(net5090));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\mem.mem[9][0] ),
    .X(net5091));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\mem.mem[43][5] ),
    .X(net5092));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\mem.mem[90][3] ),
    .X(net5093));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\mem.mem[139][6] ),
    .X(net5094));
 sg13g2_dlygate4sd3_1 hold1965 (.A(\mem.mem[5][4] ),
    .X(net5095));
 sg13g2_dlygate4sd3_1 hold1966 (.A(\mem.mem[25][0] ),
    .X(net5096));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\mem.mem[189][3] ),
    .X(net5097));
 sg13g2_dlygate4sd3_1 hold1968 (.A(\mem_A[7] ),
    .X(net5098));
 sg13g2_dlygate4sd3_1 hold1969 (.A(_00653_),
    .X(net5099));
 sg13g2_dlygate4sd3_1 hold1970 (.A(\mem.mem[86][5] ),
    .X(net5100));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\mem.mem[147][0] ),
    .X(net5101));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\mem.mem[194][2] ),
    .X(net5102));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\mem.mem[135][3] ),
    .X(net5103));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\mem.mem[221][7] ),
    .X(net5104));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\mem.mem[216][7] ),
    .X(net5105));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\mem.mem[178][3] ),
    .X(net5106));
 sg13g2_dlygate4sd3_1 hold1977 (.A(\mem.mem[27][4] ),
    .X(net5107));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\mem.mem[41][1] ),
    .X(net5108));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\mem.mem[13][5] ),
    .X(net5109));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\mem.mem[185][0] ),
    .X(net5110));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\mem.mem[204][4] ),
    .X(net5111));
 sg13g2_dlygate4sd3_1 hold1982 (.A(\mem.mem[155][6] ),
    .X(net5112));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\mem.mem[37][6] ),
    .X(net5113));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\mem.mem[34][0] ),
    .X(net5114));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\mem.mem[190][6] ),
    .X(net5115));
 sg13g2_dlygate4sd3_1 hold1986 (.A(\mem.mem[187][0] ),
    .X(net5116));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\mem.mem[124][1] ),
    .X(net5117));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\mem.mem[229][4] ),
    .X(net5118));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\mem.mem[194][0] ),
    .X(net5119));
 sg13g2_dlygate4sd3_1 hold1990 (.A(\mem.mem[71][7] ),
    .X(net5120));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\mem.mem[105][2] ),
    .X(net5121));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\mem.mem[35][2] ),
    .X(net5122));
 sg13g2_dlygate4sd3_1 hold1993 (.A(\mem.mem[163][7] ),
    .X(net5123));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\mem.mem[149][2] ),
    .X(net5124));
 sg13g2_dlygate4sd3_1 hold1995 (.A(\mem.mem[90][7] ),
    .X(net5125));
 sg13g2_dlygate4sd3_1 hold1996 (.A(\mem.mem[108][1] ),
    .X(net5126));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\mem.mem[99][5] ),
    .X(net5127));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\mem.mem[164][1] ),
    .X(net5128));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\mem.mem[195][4] ),
    .X(net5129));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\mem.mem[25][3] ),
    .X(net5130));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\mem.mem[3][5] ),
    .X(net5131));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\mem.mem[220][3] ),
    .X(net5132));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\mem.mem[182][1] ),
    .X(net5133));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\mem.mem[7][4] ),
    .X(net5134));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\mem.mem[110][3] ),
    .X(net5135));
 sg13g2_dlygate4sd3_1 hold2006 (.A(\mem.mem[219][5] ),
    .X(net5136));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\mem.mem[177][4] ),
    .X(net5137));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\mem.mem[85][5] ),
    .X(net5138));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\mem.mem[242][0] ),
    .X(net5139));
 sg13g2_dlygate4sd3_1 hold2010 (.A(\mem.mem[77][6] ),
    .X(net5140));
 sg13g2_dlygate4sd3_1 hold2011 (.A(\mem.mem[237][4] ),
    .X(net5141));
 sg13g2_dlygate4sd3_1 hold2012 (.A(\mem.mem[150][1] ),
    .X(net5142));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\mem.mem[17][6] ),
    .X(net5143));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\mem.mem[183][7] ),
    .X(net5144));
 sg13g2_dlygate4sd3_1 hold2015 (.A(\mem.mem[227][2] ),
    .X(net5145));
 sg13g2_dlygate4sd3_1 hold2016 (.A(\mem.mem[234][7] ),
    .X(net5146));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\mem.mem[1][7] ),
    .X(net5147));
 sg13g2_dlygate4sd3_1 hold2018 (.A(\mem.mem[125][0] ),
    .X(net5148));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\mem.mem[221][1] ),
    .X(net5149));
 sg13g2_dlygate4sd3_1 hold2020 (.A(\mem.mem[80][6] ),
    .X(net5150));
 sg13g2_dlygate4sd3_1 hold2021 (.A(\mem.mem[25][5] ),
    .X(net5151));
 sg13g2_dlygate4sd3_1 hold2022 (.A(\mem.mem[17][1] ),
    .X(net5152));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\mem.mem[8][4] ),
    .X(net5153));
 sg13g2_dlygate4sd3_1 hold2024 (.A(\mem.mem[202][1] ),
    .X(net5154));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\mem.mem[235][7] ),
    .X(net5155));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\mem.mem[21][7] ),
    .X(net5156));
 sg13g2_dlygate4sd3_1 hold2027 (.A(\mem.mem[7][1] ),
    .X(net5157));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\mem.mem[238][0] ),
    .X(net5158));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\mem.mem[61][7] ),
    .X(net5159));
 sg13g2_dlygate4sd3_1 hold2030 (.A(\mem.mem[122][7] ),
    .X(net5160));
 sg13g2_dlygate4sd3_1 hold2031 (.A(\mem.mem[243][4] ),
    .X(net5161));
 sg13g2_dlygate4sd3_1 hold2032 (.A(\mem.mem[23][6] ),
    .X(net5162));
 sg13g2_dlygate4sd3_1 hold2033 (.A(\mem.mem[108][4] ),
    .X(net5163));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\mem.mem[47][6] ),
    .X(net5164));
 sg13g2_dlygate4sd3_1 hold2035 (.A(\mem.mem[7][6] ),
    .X(net5165));
 sg13g2_dlygate4sd3_1 hold2036 (.A(\mem.mem[184][5] ),
    .X(net5166));
 sg13g2_dlygate4sd3_1 hold2037 (.A(\mem_A[1] ),
    .X(net5167));
 sg13g2_dlygate4sd3_1 hold2038 (.A(\mem.mem[108][3] ),
    .X(net5168));
 sg13g2_dlygate4sd3_1 hold2039 (.A(\mem.mem[67][0] ),
    .X(net5169));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\mem.mem[1][6] ),
    .X(net5170));
 sg13g2_dlygate4sd3_1 hold2041 (.A(\mem.mem[21][3] ),
    .X(net5171));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\C[4] ),
    .X(net5172));
 sg13g2_dlygate4sd3_1 hold2043 (.A(\mem.mem[53][2] ),
    .X(net5173));
 sg13g2_dlygate4sd3_1 hold2044 (.A(\mem.mem[17][4] ),
    .X(net5174));
 sg13g2_dlygate4sd3_1 hold2045 (.A(\mem.mem[54][2] ),
    .X(net5175));
 sg13g2_dlygate4sd3_1 hold2046 (.A(\mem.mem[41][5] ),
    .X(net5176));
 sg13g2_dlygate4sd3_1 hold2047 (.A(\mem.mem[102][7] ),
    .X(net5177));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\mem.mem[180][4] ),
    .X(net5178));
 sg13g2_dlygate4sd3_1 hold2049 (.A(\mem.mem[125][5] ),
    .X(net5179));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\mem.mem[179][7] ),
    .X(net5180));
 sg13g2_dlygate4sd3_1 hold2051 (.A(\C[3] ),
    .X(net5181));
 sg13g2_dlygate4sd3_1 hold2052 (.A(\A[0] ),
    .X(net5182));
 sg13g2_dlygate4sd3_1 hold2053 (.A(\mem.mem[13][2] ),
    .X(net5183));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\B[4] ),
    .X(net5184));
 sg13g2_dlygate4sd3_1 hold2055 (.A(\B[5] ),
    .X(net5185));
 sg13g2_dlygate4sd3_1 hold2056 (.A(\B[3] ),
    .X(net5186));
 sg13g2_dlygate4sd3_1 hold2057 (.A(\state[0] ),
    .X(net5187));
 sg13g2_dlygate4sd3_1 hold2058 (.A(_02388_),
    .X(net5188));
 sg13g2_dlygate4sd3_1 hold2059 (.A(_00621_),
    .X(net5189));
 sg13g2_dlygate4sd3_1 hold2060 (.A(\C[5] ),
    .X(net5190));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\A[3] ),
    .X(net5191));
 sg13g2_dlygate4sd3_1 hold2062 (.A(\B[7] ),
    .X(net5192));
 sg13g2_dlygate4sd3_1 hold2063 (.A(\A[4] ),
    .X(net5193));
 sg13g2_dlygate4sd3_1 hold2064 (.A(\A[1] ),
    .X(net5194));
 sg13g2_dlygate4sd3_1 hold2065 (.A(_00596_),
    .X(net5195));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\B[0] ),
    .X(net5196));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\A[5] ),
    .X(net5197));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\C[1] ),
    .X(net5198));
 sg13g2_dlygate4sd3_1 hold2069 (.A(\B[1] ),
    .X(net5199));
 sg13g2_dlygate4sd3_1 hold2070 (.A(\C[0] ),
    .X(net5200));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\mem_A[6] ),
    .X(net5201));
 sg13g2_dlygate4sd3_1 hold2072 (.A(_00652_),
    .X(net5202));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\mem_A[0] ),
    .X(net5203));
 sg13g2_dlygate4sd3_1 hold2074 (.A(\B[6] ),
    .X(net5204));
 sg13g2_dlygate4sd3_1 hold2075 (.A(\B[2] ),
    .X(net5205));
 sg13g2_dlygate4sd3_1 hold2076 (.A(\mem.addr[4] ),
    .X(net5206));
 sg13g2_dlygate4sd3_1 hold2077 (.A(\mem_A[4] ),
    .X(net5207));
 sg13g2_dlygate4sd3_1 hold2078 (.A(\mem_A[3] ),
    .X(net5208));
 sg13g2_dlygate4sd3_1 hold2079 (.A(\mem_A[5] ),
    .X(net5209));
 sg13g2_dlygate4sd3_1 hold2080 (.A(prev_run),
    .X(net5210));
 sg13g2_dlygate4sd3_1 hold2081 (.A(_02396_),
    .X(net5211));
 sg13g2_dlygate4sd3_1 hold2082 (.A(\PC[0] ),
    .X(net5212));
 sg13g2_dlygate4sd3_1 hold2083 (.A(_04883_),
    .X(net5213));
 sg13g2_dlygate4sd3_1 hold2084 (.A(_00622_),
    .X(net5214));
 sg13g2_dlygate4sd3_1 hold2085 (.A(\mem.addr[0] ),
    .X(net5215));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\PC[1] ),
    .X(net5216));
 sg13g2_dlygate4sd3_1 hold2087 (.A(\PC[6] ),
    .X(net5217));
 sg13g2_dlygate4sd3_1 hold2088 (.A(\mem.addr[1] ),
    .X(net5218));
 sg13g2_dlygate4sd3_1 hold2089 (.A(_00012_),
    .X(net5219));
 sg13g2_dlygate4sd3_1 hold2090 (.A(_00017_),
    .X(net5220));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\PC[4] ),
    .X(net5221));
 sg13g2_dlygate4sd3_1 hold2092 (.A(\mem.addr[2] ),
    .X(net5222));
 sg13g2_dlygate4sd3_1 hold2093 (.A(\PC[5] ),
    .X(net5223));
 sg13g2_dlygate4sd3_1 hold2094 (.A(\mem.addr[5] ),
    .X(net5224));
 sg13g2_dlygate4sd3_1 hold2095 (.A(_00016_),
    .X(net5225));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\mem.addr[7] ),
    .X(net5226));
 sg13g2_antennanp ANTENNA_1 (.A(_03950_));
 sg13g2_antennanp ANTENNA_2 (.A(_04528_));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(net3049));
 sg13g2_antennanp ANTENNA_6 (.A(net3049));
 sg13g2_antennanp ANTENNA_7 (.A(net3049));
 sg13g2_antennanp ANTENNA_8 (.A(net3049));
 sg13g2_antennanp ANTENNA_9 (.A(net3049));
 sg13g2_antennanp ANTENNA_10 (.A(net3049));
 sg13g2_antennanp ANTENNA_11 (.A(net3049));
 sg13g2_antennanp ANTENNA_12 (.A(net3049));
 sg13g2_antennanp ANTENNA_13 (.A(net3065));
 sg13g2_antennanp ANTENNA_14 (.A(net3065));
 sg13g2_antennanp ANTENNA_15 (.A(net3065));
 sg13g2_antennanp ANTENNA_16 (.A(net3065));
 sg13g2_antennanp ANTENNA_17 (.A(net3065));
 sg13g2_antennanp ANTENNA_18 (.A(net3065));
 sg13g2_antennanp ANTENNA_19 (.A(net3065));
 sg13g2_antennanp ANTENNA_20 (.A(net3065));
 sg13g2_antennanp ANTENNA_21 (.A(net3065));
 sg13g2_antennanp ANTENNA_22 (.A(net3065));
 sg13g2_antennanp ANTENNA_23 (.A(net3065));
 sg13g2_antennanp ANTENNA_24 (.A(net3065));
 sg13g2_antennanp ANTENNA_25 (.A(net3065));
 sg13g2_antennanp ANTENNA_26 (.A(net3065));
 sg13g2_antennanp ANTENNA_27 (.A(net3065));
 sg13g2_antennanp ANTENNA_28 (.A(net3065));
 sg13g2_antennanp ANTENNA_29 (.A(net3065));
 sg13g2_antennanp ANTENNA_30 (.A(net3065));
 sg13g2_antennanp ANTENNA_31 (.A(net3065));
 sg13g2_antennanp ANTENNA_32 (.A(net3065));
 sg13g2_antennanp ANTENNA_33 (.A(net3077));
 sg13g2_antennanp ANTENNA_34 (.A(net3077));
 sg13g2_antennanp ANTENNA_35 (.A(net3077));
 sg13g2_antennanp ANTENNA_36 (.A(net3077));
 sg13g2_antennanp ANTENNA_37 (.A(net3077));
 sg13g2_antennanp ANTENNA_38 (.A(net3077));
 sg13g2_antennanp ANTENNA_39 (.A(net3077));
 sg13g2_antennanp ANTENNA_40 (.A(net3077));
 sg13g2_antennanp ANTENNA_41 (.A(net3077));
 sg13g2_antennanp ANTENNA_42 (.A(net3077));
 sg13g2_antennanp ANTENNA_43 (.A(net3077));
 sg13g2_antennanp ANTENNA_44 (.A(net3077));
 sg13g2_antennanp ANTENNA_45 (.A(net3077));
 sg13g2_antennanp ANTENNA_46 (.A(net3077));
 sg13g2_antennanp ANTENNA_47 (.A(net3077));
 sg13g2_antennanp ANTENNA_48 (.A(net3077));
 sg13g2_antennanp ANTENNA_49 (.A(net3077));
 sg13g2_antennanp ANTENNA_50 (.A(net3077));
 sg13g2_antennanp ANTENNA_51 (.A(net3077));
 sg13g2_antennanp ANTENNA_52 (.A(net3077));
 sg13g2_antennanp ANTENNA_53 (.A(net3077));
 sg13g2_antennanp ANTENNA_54 (.A(net3077));
 sg13g2_antennanp ANTENNA_55 (.A(net3077));
 sg13g2_antennanp ANTENNA_56 (.A(net3077));
 sg13g2_antennanp ANTENNA_57 (.A(net3077));
 sg13g2_antennanp ANTENNA_58 (.A(net3077));
 sg13g2_antennanp ANTENNA_59 (.A(net3077));
 sg13g2_antennanp ANTENNA_60 (.A(net3077));
 sg13g2_antennanp ANTENNA_61 (.A(net3731));
 sg13g2_antennanp ANTENNA_62 (.A(net3731));
 sg13g2_antennanp ANTENNA_63 (.A(net3731));
 sg13g2_antennanp ANTENNA_64 (.A(net3731));
 sg13g2_antennanp ANTENNA_65 (.A(net3731));
 sg13g2_antennanp ANTENNA_66 (.A(net3731));
 sg13g2_antennanp ANTENNA_67 (.A(net3731));
 sg13g2_antennanp ANTENNA_68 (.A(net3731));
 sg13g2_antennanp ANTENNA_69 (.A(net3731));
 sg13g2_antennanp ANTENNA_70 (.A(net3731));
 sg13g2_antennanp ANTENNA_71 (.A(_02973_));
 sg13g2_antennanp ANTENNA_72 (.A(_03211_));
 sg13g2_antennanp ANTENNA_73 (.A(_03950_));
 sg13g2_antennanp ANTENNA_74 (.A(_04528_));
 sg13g2_antennanp ANTENNA_75 (.A(clk));
 sg13g2_antennanp ANTENNA_76 (.A(clk));
 sg13g2_antennanp ANTENNA_77 (.A(net3049));
 sg13g2_antennanp ANTENNA_78 (.A(net3049));
 sg13g2_antennanp ANTENNA_79 (.A(net3049));
 sg13g2_antennanp ANTENNA_80 (.A(net3049));
 sg13g2_antennanp ANTENNA_81 (.A(net3049));
 sg13g2_antennanp ANTENNA_82 (.A(net3049));
 sg13g2_antennanp ANTENNA_83 (.A(net3049));
 sg13g2_antennanp ANTENNA_84 (.A(net3049));
 sg13g2_antennanp ANTENNA_85 (.A(net3073));
 sg13g2_antennanp ANTENNA_86 (.A(net3073));
 sg13g2_antennanp ANTENNA_87 (.A(net3073));
 sg13g2_antennanp ANTENNA_88 (.A(net3073));
 sg13g2_antennanp ANTENNA_89 (.A(net3073));
 sg13g2_antennanp ANTENNA_90 (.A(net3073));
 sg13g2_antennanp ANTENNA_91 (.A(net3073));
 sg13g2_antennanp ANTENNA_92 (.A(net3073));
 sg13g2_antennanp ANTENNA_93 (.A(net3073));
 sg13g2_antennanp ANTENNA_94 (.A(net3073));
 sg13g2_antennanp ANTENNA_95 (.A(net3073));
 sg13g2_antennanp ANTENNA_96 (.A(net3073));
 sg13g2_antennanp ANTENNA_97 (.A(net3073));
 sg13g2_antennanp ANTENNA_98 (.A(net3073));
 sg13g2_antennanp ANTENNA_99 (.A(net3073));
 sg13g2_antennanp ANTENNA_100 (.A(net3073));
 sg13g2_antennanp ANTENNA_101 (.A(net3077));
 sg13g2_antennanp ANTENNA_102 (.A(net3077));
 sg13g2_antennanp ANTENNA_103 (.A(net3077));
 sg13g2_antennanp ANTENNA_104 (.A(net3077));
 sg13g2_antennanp ANTENNA_105 (.A(net3077));
 sg13g2_antennanp ANTENNA_106 (.A(net3077));
 sg13g2_antennanp ANTENNA_107 (.A(net3077));
 sg13g2_antennanp ANTENNA_108 (.A(net3077));
 sg13g2_antennanp ANTENNA_109 (.A(net3077));
 sg13g2_antennanp ANTENNA_110 (.A(net3077));
 sg13g2_antennanp ANTENNA_111 (.A(net3077));
 sg13g2_antennanp ANTENNA_112 (.A(net3077));
 sg13g2_antennanp ANTENNA_113 (.A(net3077));
 sg13g2_antennanp ANTENNA_114 (.A(net3077));
 sg13g2_antennanp ANTENNA_115 (.A(net3077));
 sg13g2_antennanp ANTENNA_116 (.A(net3077));
 sg13g2_antennanp ANTENNA_117 (.A(net3077));
 sg13g2_antennanp ANTENNA_118 (.A(net3077));
 sg13g2_antennanp ANTENNA_119 (.A(net3731));
 sg13g2_antennanp ANTENNA_120 (.A(net3731));
 sg13g2_antennanp ANTENNA_121 (.A(net3731));
 sg13g2_antennanp ANTENNA_122 (.A(net3731));
 sg13g2_antennanp ANTENNA_123 (.A(net3731));
 sg13g2_antennanp ANTENNA_124 (.A(net3731));
 sg13g2_antennanp ANTENNA_125 (.A(net3731));
 sg13g2_antennanp ANTENNA_126 (.A(net3731));
 sg13g2_antennanp ANTENNA_127 (.A(net3731));
 sg13g2_antennanp ANTENNA_128 (.A(net3731));
 sg13g2_antennanp ANTENNA_129 (.A(_02973_));
 sg13g2_antennanp ANTENNA_130 (.A(_03211_));
 sg13g2_antennanp ANTENNA_131 (.A(_03233_));
 sg13g2_antennanp ANTENNA_132 (.A(_03950_));
 sg13g2_antennanp ANTENNA_133 (.A(_04528_));
 sg13g2_antennanp ANTENNA_134 (.A(clk));
 sg13g2_antennanp ANTENNA_135 (.A(clk));
 sg13g2_antennanp ANTENNA_136 (.A(net3077));
 sg13g2_antennanp ANTENNA_137 (.A(net3077));
 sg13g2_antennanp ANTENNA_138 (.A(net3077));
 sg13g2_antennanp ANTENNA_139 (.A(net3077));
 sg13g2_antennanp ANTENNA_140 (.A(net3077));
 sg13g2_antennanp ANTENNA_141 (.A(net3077));
 sg13g2_antennanp ANTENNA_142 (.A(net3077));
 sg13g2_antennanp ANTENNA_143 (.A(net3077));
 sg13g2_antennanp ANTENNA_144 (.A(net3077));
 sg13g2_antennanp ANTENNA_145 (.A(net3077));
 sg13g2_antennanp ANTENNA_146 (.A(net3077));
 sg13g2_antennanp ANTENNA_147 (.A(net3077));
 sg13g2_antennanp ANTENNA_148 (.A(net3077));
 sg13g2_antennanp ANTENNA_149 (.A(net3077));
 sg13g2_antennanp ANTENNA_150 (.A(net3077));
 sg13g2_antennanp ANTENNA_151 (.A(net3077));
 sg13g2_antennanp ANTENNA_152 (.A(net3077));
 sg13g2_antennanp ANTENNA_153 (.A(net3731));
 sg13g2_antennanp ANTENNA_154 (.A(net3731));
 sg13g2_antennanp ANTENNA_155 (.A(net3731));
 sg13g2_antennanp ANTENNA_156 (.A(net3731));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_4 FILLER_0_14 ();
 sg13g2_fill_2 FILLER_0_48 ();
 sg13g2_fill_1 FILLER_0_50 ();
 sg13g2_fill_2 FILLER_0_91 ();
 sg13g2_fill_1 FILLER_0_111 ();
 sg13g2_fill_2 FILLER_0_193 ();
 sg13g2_fill_1 FILLER_0_195 ();
 sg13g2_fill_1 FILLER_0_209 ();
 sg13g2_fill_2 FILLER_0_240 ();
 sg13g2_fill_1 FILLER_0_255 ();
 sg13g2_fill_2 FILLER_0_319 ();
 sg13g2_fill_1 FILLER_0_321 ();
 sg13g2_fill_1 FILLER_0_343 ();
 sg13g2_fill_2 FILLER_0_387 ();
 sg13g2_fill_1 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_448 ();
 sg13g2_fill_2 FILLER_0_515 ();
 sg13g2_fill_2 FILLER_0_535 ();
 sg13g2_fill_2 FILLER_0_613 ();
 sg13g2_fill_2 FILLER_0_654 ();
 sg13g2_fill_1 FILLER_0_656 ();
 sg13g2_fill_1 FILLER_0_676 ();
 sg13g2_fill_1 FILLER_0_761 ();
 sg13g2_fill_2 FILLER_0_811 ();
 sg13g2_fill_1 FILLER_0_813 ();
 sg13g2_decap_8 FILLER_0_859 ();
 sg13g2_fill_1 FILLER_0_901 ();
 sg13g2_decap_8 FILLER_0_929 ();
 sg13g2_fill_1 FILLER_0_936 ();
 sg13g2_fill_1 FILLER_0_941 ();
 sg13g2_fill_2 FILLER_0_970 ();
 sg13g2_fill_2 FILLER_0_1012 ();
 sg13g2_fill_1 FILLER_0_1014 ();
 sg13g2_fill_2 FILLER_0_1043 ();
 sg13g2_fill_1 FILLER_0_1045 ();
 sg13g2_fill_1 FILLER_0_1050 ();
 sg13g2_fill_2 FILLER_0_1099 ();
 sg13g2_decap_8 FILLER_0_1128 ();
 sg13g2_decap_8 FILLER_0_1135 ();
 sg13g2_fill_2 FILLER_0_1142 ();
 sg13g2_decap_8 FILLER_0_1148 ();
 sg13g2_fill_2 FILLER_0_1155 ();
 sg13g2_fill_1 FILLER_0_1157 ();
 sg13g2_fill_2 FILLER_0_1204 ();
 sg13g2_fill_2 FILLER_0_1253 ();
 sg13g2_decap_8 FILLER_0_1323 ();
 sg13g2_fill_2 FILLER_0_1330 ();
 sg13g2_fill_2 FILLER_0_1340 ();
 sg13g2_fill_2 FILLER_0_1371 ();
 sg13g2_fill_1 FILLER_0_1373 ();
 sg13g2_fill_2 FILLER_0_1436 ();
 sg13g2_fill_1 FILLER_0_1438 ();
 sg13g2_fill_2 FILLER_0_1598 ();
 sg13g2_fill_1 FILLER_0_1600 ();
 sg13g2_decap_8 FILLER_0_1614 ();
 sg13g2_decap_8 FILLER_0_1621 ();
 sg13g2_decap_8 FILLER_0_1628 ();
 sg13g2_decap_8 FILLER_0_1635 ();
 sg13g2_decap_8 FILLER_0_1642 ();
 sg13g2_decap_8 FILLER_0_1649 ();
 sg13g2_decap_8 FILLER_0_1656 ();
 sg13g2_decap_8 FILLER_0_1663 ();
 sg13g2_decap_8 FILLER_0_1670 ();
 sg13g2_decap_8 FILLER_0_1677 ();
 sg13g2_decap_8 FILLER_0_1684 ();
 sg13g2_decap_8 FILLER_0_1691 ();
 sg13g2_decap_8 FILLER_0_1698 ();
 sg13g2_decap_8 FILLER_0_1705 ();
 sg13g2_decap_8 FILLER_0_1712 ();
 sg13g2_decap_8 FILLER_0_1719 ();
 sg13g2_decap_8 FILLER_0_1726 ();
 sg13g2_decap_8 FILLER_0_1733 ();
 sg13g2_decap_8 FILLER_0_1740 ();
 sg13g2_decap_8 FILLER_0_1747 ();
 sg13g2_decap_8 FILLER_0_1754 ();
 sg13g2_decap_8 FILLER_0_1761 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_1_7 ();
 sg13g2_fill_2 FILLER_1_70 ();
 sg13g2_fill_1 FILLER_1_72 ();
 sg13g2_fill_2 FILLER_1_213 ();
 sg13g2_fill_2 FILLER_1_326 ();
 sg13g2_fill_1 FILLER_1_328 ();
 sg13g2_fill_2 FILLER_1_365 ();
 sg13g2_fill_1 FILLER_1_367 ();
 sg13g2_fill_2 FILLER_1_466 ();
 sg13g2_fill_2 FILLER_1_583 ();
 sg13g2_fill_2 FILLER_1_634 ();
 sg13g2_fill_1 FILLER_1_636 ();
 sg13g2_fill_2 FILLER_1_719 ();
 sg13g2_fill_1 FILLER_1_721 ();
 sg13g2_fill_2 FILLER_1_790 ();
 sg13g2_fill_1 FILLER_1_792 ();
 sg13g2_decap_4 FILLER_1_864 ();
 sg13g2_fill_2 FILLER_1_990 ();
 sg13g2_fill_1 FILLER_1_1080 ();
 sg13g2_decap_4 FILLER_1_1133 ();
 sg13g2_fill_1 FILLER_1_1137 ();
 sg13g2_fill_1 FILLER_1_1450 ();
 sg13g2_fill_1 FILLER_1_1477 ();
 sg13g2_fill_1 FILLER_1_1554 ();
 sg13g2_fill_2 FILLER_1_1585 ();
 sg13g2_fill_1 FILLER_1_1587 ();
 sg13g2_fill_1 FILLER_1_1618 ();
 sg13g2_decap_8 FILLER_1_1628 ();
 sg13g2_fill_2 FILLER_1_1635 ();
 sg13g2_decap_8 FILLER_1_1641 ();
 sg13g2_decap_8 FILLER_1_1648 ();
 sg13g2_decap_8 FILLER_1_1655 ();
 sg13g2_decap_8 FILLER_1_1662 ();
 sg13g2_decap_4 FILLER_1_1669 ();
 sg13g2_fill_2 FILLER_1_1673 ();
 sg13g2_decap_8 FILLER_1_1679 ();
 sg13g2_decap_8 FILLER_1_1686 ();
 sg13g2_decap_8 FILLER_1_1693 ();
 sg13g2_decap_8 FILLER_1_1700 ();
 sg13g2_decap_8 FILLER_1_1707 ();
 sg13g2_decap_8 FILLER_1_1714 ();
 sg13g2_decap_8 FILLER_1_1721 ();
 sg13g2_decap_8 FILLER_1_1728 ();
 sg13g2_decap_8 FILLER_1_1735 ();
 sg13g2_decap_8 FILLER_1_1742 ();
 sg13g2_decap_8 FILLER_1_1749 ();
 sg13g2_decap_8 FILLER_1_1756 ();
 sg13g2_decap_4 FILLER_1_1763 ();
 sg13g2_fill_1 FILLER_1_1767 ();
 sg13g2_decap_4 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_29 ();
 sg13g2_fill_2 FILLER_2_40 ();
 sg13g2_fill_1 FILLER_2_42 ();
 sg13g2_fill_2 FILLER_2_72 ();
 sg13g2_fill_1 FILLER_2_84 ();
 sg13g2_fill_1 FILLER_2_95 ();
 sg13g2_fill_2 FILLER_2_131 ();
 sg13g2_fill_1 FILLER_2_143 ();
 sg13g2_fill_2 FILLER_2_168 ();
 sg13g2_fill_2 FILLER_2_254 ();
 sg13g2_fill_2 FILLER_2_291 ();
 sg13g2_fill_1 FILLER_2_293 ();
 sg13g2_fill_2 FILLER_2_318 ();
 sg13g2_fill_2 FILLER_2_339 ();
 sg13g2_fill_2 FILLER_2_373 ();
 sg13g2_fill_2 FILLER_2_424 ();
 sg13g2_fill_2 FILLER_2_490 ();
 sg13g2_fill_1 FILLER_2_492 ();
 sg13g2_fill_1 FILLER_2_537 ();
 sg13g2_fill_2 FILLER_2_599 ();
 sg13g2_fill_2 FILLER_2_611 ();
 sg13g2_fill_2 FILLER_2_632 ();
 sg13g2_fill_1 FILLER_2_663 ();
 sg13g2_fill_1 FILLER_2_685 ();
 sg13g2_fill_1 FILLER_2_700 ();
 sg13g2_fill_1 FILLER_2_797 ();
 sg13g2_decap_4 FILLER_2_842 ();
 sg13g2_fill_2 FILLER_2_846 ();
 sg13g2_decap_8 FILLER_2_920 ();
 sg13g2_decap_8 FILLER_2_927 ();
 sg13g2_fill_2 FILLER_2_987 ();
 sg13g2_fill_1 FILLER_2_989 ();
 sg13g2_fill_2 FILLER_2_1000 ();
 sg13g2_fill_1 FILLER_2_1002 ();
 sg13g2_decap_4 FILLER_2_1046 ();
 sg13g2_fill_1 FILLER_2_1050 ();
 sg13g2_fill_1 FILLER_2_1121 ();
 sg13g2_fill_1 FILLER_2_1183 ();
 sg13g2_decap_8 FILLER_2_1194 ();
 sg13g2_fill_2 FILLER_2_1210 ();
 sg13g2_fill_1 FILLER_2_1227 ();
 sg13g2_fill_1 FILLER_2_1271 ();
 sg13g2_fill_1 FILLER_2_1295 ();
 sg13g2_fill_2 FILLER_2_1340 ();
 sg13g2_fill_1 FILLER_2_1342 ();
 sg13g2_fill_2 FILLER_2_1377 ();
 sg13g2_fill_1 FILLER_2_1379 ();
 sg13g2_fill_2 FILLER_2_1395 ();
 sg13g2_fill_2 FILLER_2_1476 ();
 sg13g2_fill_1 FILLER_2_1478 ();
 sg13g2_fill_1 FILLER_2_1505 ();
 sg13g2_fill_2 FILLER_2_1542 ();
 sg13g2_fill_1 FILLER_2_1544 ();
 sg13g2_fill_1 FILLER_2_1578 ();
 sg13g2_decap_8 FILLER_2_1647 ();
 sg13g2_decap_4 FILLER_2_1654 ();
 sg13g2_fill_1 FILLER_2_1658 ();
 sg13g2_fill_2 FILLER_2_1672 ();
 sg13g2_decap_4 FILLER_2_1689 ();
 sg13g2_decap_8 FILLER_2_1702 ();
 sg13g2_decap_8 FILLER_2_1709 ();
 sg13g2_decap_8 FILLER_2_1716 ();
 sg13g2_decap_8 FILLER_2_1723 ();
 sg13g2_decap_8 FILLER_2_1730 ();
 sg13g2_decap_8 FILLER_2_1737 ();
 sg13g2_decap_8 FILLER_2_1744 ();
 sg13g2_decap_8 FILLER_2_1751 ();
 sg13g2_decap_8 FILLER_2_1758 ();
 sg13g2_fill_2 FILLER_2_1765 ();
 sg13g2_fill_1 FILLER_2_1767 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_27 ();
 sg13g2_fill_1 FILLER_3_29 ();
 sg13g2_fill_2 FILLER_3_70 ();
 sg13g2_fill_2 FILLER_3_121 ();
 sg13g2_fill_1 FILLER_3_123 ();
 sg13g2_fill_1 FILLER_3_133 ();
 sg13g2_fill_2 FILLER_3_196 ();
 sg13g2_fill_2 FILLER_3_252 ();
 sg13g2_fill_1 FILLER_3_254 ();
 sg13g2_fill_2 FILLER_3_277 ();
 sg13g2_fill_2 FILLER_3_340 ();
 sg13g2_fill_1 FILLER_3_342 ();
 sg13g2_fill_1 FILLER_3_417 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_fill_2 FILLER_3_562 ();
 sg13g2_fill_1 FILLER_3_564 ();
 sg13g2_fill_2 FILLER_3_686 ();
 sg13g2_fill_1 FILLER_3_688 ();
 sg13g2_fill_1 FILLER_3_750 ();
 sg13g2_fill_2 FILLER_3_756 ();
 sg13g2_fill_1 FILLER_3_758 ();
 sg13g2_fill_1 FILLER_3_966 ();
 sg13g2_fill_2 FILLER_3_986 ();
 sg13g2_fill_2 FILLER_3_1024 ();
 sg13g2_fill_1 FILLER_3_1026 ();
 sg13g2_fill_2 FILLER_3_1053 ();
 sg13g2_fill_2 FILLER_3_1117 ();
 sg13g2_fill_1 FILLER_3_1147 ();
 sg13g2_fill_2 FILLER_3_1184 ();
 sg13g2_fill_1 FILLER_3_1186 ();
 sg13g2_fill_1 FILLER_3_1213 ();
 sg13g2_fill_1 FILLER_3_1301 ();
 sg13g2_fill_2 FILLER_3_1354 ();
 sg13g2_fill_1 FILLER_3_1356 ();
 sg13g2_fill_2 FILLER_3_1492 ();
 sg13g2_fill_1 FILLER_3_1494 ();
 sg13g2_fill_2 FILLER_3_1515 ();
 sg13g2_fill_2 FILLER_3_1542 ();
 sg13g2_fill_2 FILLER_3_1615 ();
 sg13g2_fill_1 FILLER_3_1617 ();
 sg13g2_fill_2 FILLER_3_1641 ();
 sg13g2_fill_2 FILLER_3_1679 ();
 sg13g2_fill_1 FILLER_3_1681 ();
 sg13g2_decap_8 FILLER_3_1717 ();
 sg13g2_decap_8 FILLER_3_1724 ();
 sg13g2_decap_8 FILLER_3_1731 ();
 sg13g2_decap_8 FILLER_3_1738 ();
 sg13g2_decap_8 FILLER_3_1745 ();
 sg13g2_decap_8 FILLER_3_1752 ();
 sg13g2_decap_8 FILLER_3_1759 ();
 sg13g2_fill_2 FILLER_3_1766 ();
 sg13g2_fill_1 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_153 ();
 sg13g2_fill_1 FILLER_4_155 ();
 sg13g2_fill_2 FILLER_4_177 ();
 sg13g2_fill_2 FILLER_4_231 ();
 sg13g2_fill_2 FILLER_4_259 ();
 sg13g2_fill_1 FILLER_4_261 ();
 sg13g2_fill_2 FILLER_4_298 ();
 sg13g2_fill_2 FILLER_4_322 ();
 sg13g2_fill_2 FILLER_4_345 ();
 sg13g2_fill_2 FILLER_4_479 ();
 sg13g2_fill_1 FILLER_4_524 ();
 sg13g2_fill_2 FILLER_4_570 ();
 sg13g2_fill_1 FILLER_4_572 ();
 sg13g2_fill_2 FILLER_4_587 ();
 sg13g2_fill_2 FILLER_4_628 ();
 sg13g2_fill_1 FILLER_4_630 ();
 sg13g2_fill_2 FILLER_4_653 ();
 sg13g2_fill_1 FILLER_4_665 ();
 sg13g2_fill_1 FILLER_4_670 ();
 sg13g2_fill_2 FILLER_4_704 ();
 sg13g2_fill_1 FILLER_4_770 ();
 sg13g2_fill_2 FILLER_4_799 ();
 sg13g2_fill_1 FILLER_4_801 ();
 sg13g2_fill_2 FILLER_4_823 ();
 sg13g2_fill_1 FILLER_4_825 ();
 sg13g2_fill_1 FILLER_4_849 ();
 sg13g2_fill_1 FILLER_4_863 ();
 sg13g2_fill_2 FILLER_4_919 ();
 sg13g2_fill_1 FILLER_4_926 ();
 sg13g2_fill_2 FILLER_4_935 ();
 sg13g2_fill_2 FILLER_4_963 ();
 sg13g2_fill_1 FILLER_4_965 ();
 sg13g2_fill_2 FILLER_4_1002 ();
 sg13g2_fill_2 FILLER_4_1013 ();
 sg13g2_fill_1 FILLER_4_1015 ();
 sg13g2_fill_2 FILLER_4_1126 ();
 sg13g2_fill_1 FILLER_4_1128 ();
 sg13g2_fill_2 FILLER_4_1137 ();
 sg13g2_fill_2 FILLER_4_1149 ();
 sg13g2_fill_1 FILLER_4_1151 ();
 sg13g2_fill_2 FILLER_4_1206 ();
 sg13g2_fill_2 FILLER_4_1235 ();
 sg13g2_fill_1 FILLER_4_1246 ();
 sg13g2_fill_2 FILLER_4_1260 ();
 sg13g2_fill_2 FILLER_4_1276 ();
 sg13g2_fill_1 FILLER_4_1278 ();
 sg13g2_fill_1 FILLER_4_1329 ();
 sg13g2_fill_2 FILLER_4_1395 ();
 sg13g2_fill_1 FILLER_4_1397 ();
 sg13g2_fill_2 FILLER_4_1460 ();
 sg13g2_fill_1 FILLER_4_1462 ();
 sg13g2_fill_2 FILLER_4_1499 ();
 sg13g2_fill_1 FILLER_4_1501 ();
 sg13g2_fill_2 FILLER_4_1528 ();
 sg13g2_fill_1 FILLER_4_1530 ();
 sg13g2_fill_2 FILLER_4_1539 ();
 sg13g2_fill_2 FILLER_4_1577 ();
 sg13g2_fill_1 FILLER_4_1579 ();
 sg13g2_fill_2 FILLER_4_1609 ();
 sg13g2_fill_1 FILLER_4_1611 ();
 sg13g2_fill_2 FILLER_4_1683 ();
 sg13g2_decap_8 FILLER_4_1721 ();
 sg13g2_decap_8 FILLER_4_1728 ();
 sg13g2_decap_8 FILLER_4_1735 ();
 sg13g2_decap_8 FILLER_4_1742 ();
 sg13g2_decap_8 FILLER_4_1749 ();
 sg13g2_decap_8 FILLER_4_1756 ();
 sg13g2_decap_4 FILLER_4_1763 ();
 sg13g2_fill_1 FILLER_4_1767 ();
 sg13g2_fill_1 FILLER_5_40 ();
 sg13g2_fill_1 FILLER_5_67 ();
 sg13g2_fill_1 FILLER_5_98 ();
 sg13g2_fill_1 FILLER_5_109 ();
 sg13g2_fill_1 FILLER_5_119 ();
 sg13g2_fill_2 FILLER_5_204 ();
 sg13g2_fill_2 FILLER_5_233 ();
 sg13g2_fill_1 FILLER_5_235 ();
 sg13g2_fill_2 FILLER_5_250 ();
 sg13g2_fill_1 FILLER_5_252 ();
 sg13g2_fill_2 FILLER_5_273 ();
 sg13g2_fill_2 FILLER_5_299 ();
 sg13g2_fill_1 FILLER_5_337 ();
 sg13g2_fill_2 FILLER_5_353 ();
 sg13g2_fill_2 FILLER_5_364 ();
 sg13g2_fill_1 FILLER_5_366 ();
 sg13g2_fill_2 FILLER_5_397 ();
 sg13g2_fill_1 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_449 ();
 sg13g2_fill_1 FILLER_5_461 ();
 sg13g2_fill_1 FILLER_5_488 ();
 sg13g2_fill_2 FILLER_5_498 ();
 sg13g2_fill_2 FILLER_5_526 ();
 sg13g2_fill_2 FILLER_5_538 ();
 sg13g2_fill_2 FILLER_5_601 ();
 sg13g2_fill_1 FILLER_5_603 ();
 sg13g2_fill_2 FILLER_5_623 ();
 sg13g2_fill_1 FILLER_5_634 ();
 sg13g2_fill_2 FILLER_5_684 ();
 sg13g2_fill_2 FILLER_5_738 ();
 sg13g2_fill_1 FILLER_5_740 ();
 sg13g2_fill_1 FILLER_5_764 ();
 sg13g2_fill_1 FILLER_5_837 ();
 sg13g2_fill_2 FILLER_5_942 ();
 sg13g2_fill_1 FILLER_5_944 ();
 sg13g2_fill_2 FILLER_5_983 ();
 sg13g2_fill_1 FILLER_5_985 ();
 sg13g2_fill_2 FILLER_5_1008 ();
 sg13g2_fill_1 FILLER_5_1033 ();
 sg13g2_fill_2 FILLER_5_1065 ();
 sg13g2_fill_2 FILLER_5_1077 ();
 sg13g2_fill_1 FILLER_5_1079 ();
 sg13g2_fill_2 FILLER_5_1110 ();
 sg13g2_fill_1 FILLER_5_1112 ();
 sg13g2_fill_2 FILLER_5_1174 ();
 sg13g2_fill_2 FILLER_5_1221 ();
 sg13g2_fill_1 FILLER_5_1223 ();
 sg13g2_fill_2 FILLER_5_1260 ();
 sg13g2_fill_1 FILLER_5_1262 ();
 sg13g2_fill_2 FILLER_5_1282 ();
 sg13g2_fill_1 FILLER_5_1284 ();
 sg13g2_fill_2 FILLER_5_1322 ();
 sg13g2_fill_1 FILLER_5_1324 ();
 sg13g2_fill_1 FILLER_5_1345 ();
 sg13g2_fill_1 FILLER_5_1377 ();
 sg13g2_fill_2 FILLER_5_1470 ();
 sg13g2_fill_1 FILLER_5_1482 ();
 sg13g2_fill_2 FILLER_5_1529 ();
 sg13g2_fill_2 FILLER_5_1535 ();
 sg13g2_fill_1 FILLER_5_1547 ();
 sg13g2_fill_1 FILLER_5_1572 ();
 sg13g2_fill_2 FILLER_5_1588 ();
 sg13g2_fill_1 FILLER_5_1590 ();
 sg13g2_fill_1 FILLER_5_1622 ();
 sg13g2_decap_4 FILLER_5_1633 ();
 sg13g2_fill_1 FILLER_5_1637 ();
 sg13g2_fill_1 FILLER_5_1668 ();
 sg13g2_fill_2 FILLER_5_1700 ();
 sg13g2_decap_8 FILLER_5_1728 ();
 sg13g2_decap_8 FILLER_5_1735 ();
 sg13g2_decap_8 FILLER_5_1742 ();
 sg13g2_decap_8 FILLER_5_1749 ();
 sg13g2_decap_8 FILLER_5_1756 ();
 sg13g2_decap_4 FILLER_5_1763 ();
 sg13g2_fill_1 FILLER_5_1767 ();
 sg13g2_fill_2 FILLER_6_26 ();
 sg13g2_fill_2 FILLER_6_74 ();
 sg13g2_fill_2 FILLER_6_95 ();
 sg13g2_fill_2 FILLER_6_138 ();
 sg13g2_fill_2 FILLER_6_150 ();
 sg13g2_fill_2 FILLER_6_166 ();
 sg13g2_fill_1 FILLER_6_168 ();
 sg13g2_fill_2 FILLER_6_184 ();
 sg13g2_fill_1 FILLER_6_186 ();
 sg13g2_fill_1 FILLER_6_263 ();
 sg13g2_fill_1 FILLER_6_295 ();
 sg13g2_fill_1 FILLER_6_368 ();
 sg13g2_fill_2 FILLER_6_424 ();
 sg13g2_fill_1 FILLER_6_426 ();
 sg13g2_fill_2 FILLER_6_467 ();
 sg13g2_fill_2 FILLER_6_527 ();
 sg13g2_fill_2 FILLER_6_565 ();
 sg13g2_fill_2 FILLER_6_650 ();
 sg13g2_fill_1 FILLER_6_652 ();
 sg13g2_fill_2 FILLER_6_661 ();
 sg13g2_fill_1 FILLER_6_663 ();
 sg13g2_fill_2 FILLER_6_683 ();
 sg13g2_fill_2 FILLER_6_690 ();
 sg13g2_fill_1 FILLER_6_702 ();
 sg13g2_fill_1 FILLER_6_769 ();
 sg13g2_fill_2 FILLER_6_775 ();
 sg13g2_decap_4 FILLER_6_807 ();
 sg13g2_decap_8 FILLER_6_852 ();
 sg13g2_decap_4 FILLER_6_901 ();
 sg13g2_fill_2 FILLER_6_905 ();
 sg13g2_fill_1 FILLER_6_935 ();
 sg13g2_fill_2 FILLER_6_972 ();
 sg13g2_fill_1 FILLER_6_974 ();
 sg13g2_decap_8 FILLER_6_1134 ();
 sg13g2_decap_4 FILLER_6_1141 ();
 sg13g2_fill_1 FILLER_6_1145 ();
 sg13g2_fill_2 FILLER_6_1164 ();
 sg13g2_fill_1 FILLER_6_1166 ();
 sg13g2_fill_2 FILLER_6_1226 ();
 sg13g2_fill_2 FILLER_6_1258 ();
 sg13g2_fill_2 FILLER_6_1305 ();
 sg13g2_fill_2 FILLER_6_1413 ();
 sg13g2_fill_2 FILLER_6_1446 ();
 sg13g2_fill_1 FILLER_6_1474 ();
 sg13g2_fill_1 FILLER_6_1531 ();
 sg13g2_fill_2 FILLER_6_1549 ();
 sg13g2_fill_1 FILLER_6_1551 ();
 sg13g2_fill_2 FILLER_6_1569 ();
 sg13g2_fill_1 FILLER_6_1571 ();
 sg13g2_decap_8 FILLER_6_1727 ();
 sg13g2_decap_8 FILLER_6_1734 ();
 sg13g2_decap_8 FILLER_6_1741 ();
 sg13g2_decap_8 FILLER_6_1748 ();
 sg13g2_decap_8 FILLER_6_1755 ();
 sg13g2_decap_4 FILLER_6_1762 ();
 sg13g2_fill_2 FILLER_6_1766 ();
 sg13g2_fill_1 FILLER_7_43 ();
 sg13g2_fill_1 FILLER_7_70 ();
 sg13g2_fill_2 FILLER_7_140 ();
 sg13g2_fill_1 FILLER_7_142 ();
 sg13g2_fill_2 FILLER_7_205 ();
 sg13g2_fill_2 FILLER_7_246 ();
 sg13g2_fill_1 FILLER_7_248 ();
 sg13g2_fill_2 FILLER_7_263 ();
 sg13g2_fill_1 FILLER_7_265 ();
 sg13g2_fill_1 FILLER_7_294 ();
 sg13g2_fill_1 FILLER_7_351 ();
 sg13g2_fill_1 FILLER_7_379 ();
 sg13g2_fill_2 FILLER_7_399 ();
 sg13g2_fill_1 FILLER_7_459 ();
 sg13g2_fill_2 FILLER_7_469 ();
 sg13g2_fill_2 FILLER_7_499 ();
 sg13g2_fill_2 FILLER_7_516 ();
 sg13g2_fill_1 FILLER_7_526 ();
 sg13g2_fill_2 FILLER_7_546 ();
 sg13g2_fill_2 FILLER_7_584 ();
 sg13g2_fill_1 FILLER_7_586 ();
 sg13g2_fill_2 FILLER_7_613 ();
 sg13g2_fill_1 FILLER_7_615 ();
 sg13g2_fill_2 FILLER_7_671 ();
 sg13g2_fill_1 FILLER_7_673 ();
 sg13g2_fill_2 FILLER_7_714 ();
 sg13g2_fill_2 FILLER_7_751 ();
 sg13g2_fill_1 FILLER_7_753 ();
 sg13g2_fill_2 FILLER_7_790 ();
 sg13g2_fill_1 FILLER_7_822 ();
 sg13g2_decap_4 FILLER_7_836 ();
 sg13g2_fill_2 FILLER_7_840 ();
 sg13g2_decap_4 FILLER_7_913 ();
 sg13g2_fill_2 FILLER_7_917 ();
 sg13g2_fill_2 FILLER_7_924 ();
 sg13g2_fill_1 FILLER_7_931 ();
 sg13g2_fill_2 FILLER_7_987 ();
 sg13g2_fill_1 FILLER_7_998 ();
 sg13g2_fill_2 FILLER_7_1012 ();
 sg13g2_fill_2 FILLER_7_1083 ();
 sg13g2_fill_1 FILLER_7_1121 ();
 sg13g2_fill_2 FILLER_7_1153 ();
 sg13g2_fill_1 FILLER_7_1155 ();
 sg13g2_fill_1 FILLER_7_1196 ();
 sg13g2_fill_2 FILLER_7_1251 ();
 sg13g2_fill_2 FILLER_7_1263 ();
 sg13g2_fill_2 FILLER_7_1291 ();
 sg13g2_fill_1 FILLER_7_1293 ();
 sg13g2_fill_2 FILLER_7_1349 ();
 sg13g2_fill_1 FILLER_7_1390 ();
 sg13g2_fill_2 FILLER_7_1421 ();
 sg13g2_fill_1 FILLER_7_1423 ();
 sg13g2_fill_2 FILLER_7_1434 ();
 sg13g2_fill_1 FILLER_7_1436 ();
 sg13g2_fill_2 FILLER_7_1457 ();
 sg13g2_fill_1 FILLER_7_1459 ();
 sg13g2_fill_2 FILLER_7_1474 ();
 sg13g2_fill_1 FILLER_7_1476 ();
 sg13g2_fill_1 FILLER_7_1487 ();
 sg13g2_fill_2 FILLER_7_1512 ();
 sg13g2_fill_2 FILLER_7_1552 ();
 sg13g2_fill_1 FILLER_7_1554 ();
 sg13g2_fill_1 FILLER_7_1624 ();
 sg13g2_fill_1 FILLER_7_1682 ();
 sg13g2_decap_4 FILLER_7_1697 ();
 sg13g2_fill_1 FILLER_7_1701 ();
 sg13g2_decap_8 FILLER_7_1723 ();
 sg13g2_decap_8 FILLER_7_1730 ();
 sg13g2_decap_8 FILLER_7_1737 ();
 sg13g2_decap_8 FILLER_7_1744 ();
 sg13g2_decap_8 FILLER_7_1751 ();
 sg13g2_decap_8 FILLER_7_1758 ();
 sg13g2_fill_2 FILLER_7_1765 ();
 sg13g2_fill_1 FILLER_7_1767 ();
 sg13g2_fill_2 FILLER_8_55 ();
 sg13g2_fill_2 FILLER_8_124 ();
 sg13g2_fill_2 FILLER_8_149 ();
 sg13g2_fill_1 FILLER_8_151 ();
 sg13g2_fill_2 FILLER_8_188 ();
 sg13g2_fill_1 FILLER_8_190 ();
 sg13g2_fill_2 FILLER_8_300 ();
 sg13g2_fill_1 FILLER_8_302 ();
 sg13g2_fill_1 FILLER_8_363 ();
 sg13g2_fill_1 FILLER_8_486 ();
 sg13g2_fill_2 FILLER_8_527 ();
 sg13g2_fill_2 FILLER_8_565 ();
 sg13g2_fill_1 FILLER_8_567 ();
 sg13g2_fill_2 FILLER_8_597 ();
 sg13g2_fill_1 FILLER_8_664 ();
 sg13g2_fill_2 FILLER_8_717 ();
 sg13g2_fill_1 FILLER_8_719 ();
 sg13g2_fill_2 FILLER_8_786 ();
 sg13g2_fill_1 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_839 ();
 sg13g2_decap_8 FILLER_8_846 ();
 sg13g2_fill_2 FILLER_8_857 ();
 sg13g2_fill_2 FILLER_8_883 ();
 sg13g2_fill_2 FILLER_8_903 ();
 sg13g2_decap_4 FILLER_8_914 ();
 sg13g2_decap_4 FILLER_8_944 ();
 sg13g2_fill_1 FILLER_8_1020 ();
 sg13g2_fill_1 FILLER_8_1087 ();
 sg13g2_fill_1 FILLER_8_1154 ();
 sg13g2_fill_2 FILLER_8_1163 ();
 sg13g2_fill_1 FILLER_8_1165 ();
 sg13g2_fill_2 FILLER_8_1180 ();
 sg13g2_fill_1 FILLER_8_1182 ();
 sg13g2_fill_2 FILLER_8_1197 ();
 sg13g2_fill_1 FILLER_8_1199 ();
 sg13g2_fill_1 FILLER_8_1261 ();
 sg13g2_decap_4 FILLER_8_1298 ();
 sg13g2_fill_2 FILLER_8_1331 ();
 sg13g2_fill_1 FILLER_8_1333 ();
 sg13g2_fill_2 FILLER_8_1386 ();
 sg13g2_fill_1 FILLER_8_1388 ();
 sg13g2_fill_2 FILLER_8_1408 ();
 sg13g2_fill_2 FILLER_8_1446 ();
 sg13g2_fill_2 FILLER_8_1474 ();
 sg13g2_fill_2 FILLER_8_1536 ();
 sg13g2_fill_2 FILLER_8_1564 ();
 sg13g2_fill_1 FILLER_8_1594 ();
 sg13g2_fill_2 FILLER_8_1619 ();
 sg13g2_fill_1 FILLER_8_1621 ();
 sg13g2_fill_2 FILLER_8_1683 ();
 sg13g2_fill_1 FILLER_8_1685 ();
 sg13g2_decap_8 FILLER_8_1731 ();
 sg13g2_decap_8 FILLER_8_1738 ();
 sg13g2_decap_4 FILLER_8_1745 ();
 sg13g2_fill_2 FILLER_8_1749 ();
 sg13g2_decap_8 FILLER_8_1755 ();
 sg13g2_decap_4 FILLER_8_1762 ();
 sg13g2_fill_2 FILLER_8_1766 ();
 sg13g2_fill_1 FILLER_9_26 ();
 sg13g2_fill_1 FILLER_9_67 ();
 sg13g2_fill_2 FILLER_9_113 ();
 sg13g2_fill_1 FILLER_9_115 ();
 sg13g2_fill_2 FILLER_9_159 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_fill_2 FILLER_9_172 ();
 sg13g2_fill_1 FILLER_9_174 ();
 sg13g2_fill_2 FILLER_9_211 ();
 sg13g2_fill_2 FILLER_9_256 ();
 sg13g2_fill_2 FILLER_9_267 ();
 sg13g2_fill_2 FILLER_9_343 ();
 sg13g2_fill_1 FILLER_9_345 ();
 sg13g2_fill_1 FILLER_9_404 ();
 sg13g2_decap_8 FILLER_9_409 ();
 sg13g2_fill_1 FILLER_9_416 ();
 sg13g2_fill_2 FILLER_9_493 ();
 sg13g2_fill_2 FILLER_9_565 ();
 sg13g2_fill_1 FILLER_9_621 ();
 sg13g2_fill_2 FILLER_9_632 ();
 sg13g2_fill_2 FILLER_9_672 ();
 sg13g2_fill_2 FILLER_9_687 ();
 sg13g2_fill_2 FILLER_9_725 ();
 sg13g2_fill_2 FILLER_9_814 ();
 sg13g2_fill_1 FILLER_9_816 ();
 sg13g2_fill_2 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_838 ();
 sg13g2_fill_2 FILLER_9_845 ();
 sg13g2_fill_1 FILLER_9_847 ();
 sg13g2_fill_2 FILLER_9_883 ();
 sg13g2_fill_1 FILLER_9_885 ();
 sg13g2_fill_1 FILLER_9_931 ();
 sg13g2_fill_1 FILLER_9_995 ();
 sg13g2_fill_2 FILLER_9_1010 ();
 sg13g2_fill_2 FILLER_9_1051 ();
 sg13g2_fill_1 FILLER_9_1085 ();
 sg13g2_fill_2 FILLER_9_1109 ();
 sg13g2_fill_1 FILLER_9_1172 ();
 sg13g2_fill_1 FILLER_9_1213 ();
 sg13g2_fill_2 FILLER_9_1236 ();
 sg13g2_fill_2 FILLER_9_1251 ();
 sg13g2_fill_1 FILLER_9_1253 ();
 sg13g2_fill_1 FILLER_9_1264 ();
 sg13g2_decap_8 FILLER_9_1291 ();
 sg13g2_decap_8 FILLER_9_1298 ();
 sg13g2_fill_1 FILLER_9_1305 ();
 sg13g2_fill_2 FILLER_9_1342 ();
 sg13g2_fill_1 FILLER_9_1344 ();
 sg13g2_fill_2 FILLER_9_1349 ();
 sg13g2_fill_1 FILLER_9_1370 ();
 sg13g2_fill_2 FILLER_9_1420 ();
 sg13g2_fill_2 FILLER_9_1437 ();
 sg13g2_fill_1 FILLER_9_1439 ();
 sg13g2_fill_2 FILLER_9_1457 ();
 sg13g2_fill_1 FILLER_9_1467 ();
 sg13g2_fill_1 FILLER_9_1513 ();
 sg13g2_fill_1 FILLER_9_1523 ();
 sg13g2_fill_2 FILLER_9_1542 ();
 sg13g2_fill_2 FILLER_9_1567 ();
 sg13g2_fill_1 FILLER_9_1569 ();
 sg13g2_fill_2 FILLER_9_1633 ();
 sg13g2_fill_1 FILLER_9_1684 ();
 sg13g2_fill_1 FILLER_9_1695 ();
 sg13g2_decap_4 FILLER_9_1740 ();
 sg13g2_fill_2 FILLER_9_1744 ();
 sg13g2_decap_4 FILLER_9_1764 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_38 ();
 sg13g2_fill_2 FILLER_10_48 ();
 sg13g2_fill_1 FILLER_10_50 ();
 sg13g2_fill_2 FILLER_10_204 ();
 sg13g2_fill_1 FILLER_10_206 ();
 sg13g2_fill_2 FILLER_10_309 ();
 sg13g2_fill_1 FILLER_10_311 ();
 sg13g2_fill_2 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_419 ();
 sg13g2_decap_4 FILLER_10_426 ();
 sg13g2_fill_1 FILLER_10_436 ();
 sg13g2_fill_2 FILLER_10_482 ();
 sg13g2_fill_1 FILLER_10_520 ();
 sg13g2_fill_1 FILLER_10_544 ();
 sg13g2_fill_2 FILLER_10_676 ();
 sg13g2_fill_1 FILLER_10_678 ();
 sg13g2_fill_2 FILLER_10_741 ();
 sg13g2_fill_1 FILLER_10_758 ();
 sg13g2_decap_4 FILLER_10_817 ();
 sg13g2_fill_2 FILLER_10_857 ();
 sg13g2_fill_2 FILLER_10_967 ();
 sg13g2_fill_2 FILLER_10_1095 ();
 sg13g2_fill_1 FILLER_10_1132 ();
 sg13g2_fill_1 FILLER_10_1250 ();
 sg13g2_fill_2 FILLER_10_1278 ();
 sg13g2_fill_1 FILLER_10_1280 ();
 sg13g2_fill_2 FILLER_10_1338 ();
 sg13g2_fill_2 FILLER_10_1344 ();
 sg13g2_fill_1 FILLER_10_1356 ();
 sg13g2_fill_2 FILLER_10_1366 ();
 sg13g2_fill_1 FILLER_10_1368 ();
 sg13g2_fill_2 FILLER_10_1382 ();
 sg13g2_fill_1 FILLER_10_1384 ();
 sg13g2_fill_2 FILLER_10_1434 ();
 sg13g2_fill_1 FILLER_10_1436 ();
 sg13g2_fill_2 FILLER_10_1451 ();
 sg13g2_fill_1 FILLER_10_1453 ();
 sg13g2_fill_2 FILLER_10_1458 ();
 sg13g2_fill_2 FILLER_10_1496 ();
 sg13g2_fill_1 FILLER_10_1498 ();
 sg13g2_fill_2 FILLER_10_1534 ();
 sg13g2_fill_2 FILLER_10_1553 ();
 sg13g2_fill_2 FILLER_10_1583 ();
 sg13g2_fill_1 FILLER_10_1585 ();
 sg13g2_fill_1 FILLER_10_1619 ();
 sg13g2_fill_1 FILLER_10_1661 ();
 sg13g2_fill_2 FILLER_10_1686 ();
 sg13g2_fill_1 FILLER_10_1688 ();
 sg13g2_fill_1 FILLER_10_1725 ();
 sg13g2_fill_1 FILLER_10_1736 ();
 sg13g2_fill_1 FILLER_10_1767 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_36 ();
 sg13g2_fill_1 FILLER_11_50 ();
 sg13g2_fill_2 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_79 ();
 sg13g2_fill_1 FILLER_11_99 ();
 sg13g2_fill_2 FILLER_11_118 ();
 sg13g2_fill_2 FILLER_11_181 ();
 sg13g2_fill_1 FILLER_11_183 ();
 sg13g2_fill_2 FILLER_11_263 ();
 sg13g2_fill_1 FILLER_11_265 ();
 sg13g2_fill_2 FILLER_11_271 ();
 sg13g2_fill_1 FILLER_11_273 ();
 sg13g2_fill_1 FILLER_11_279 ();
 sg13g2_fill_1 FILLER_11_310 ();
 sg13g2_fill_2 FILLER_11_354 ();
 sg13g2_fill_2 FILLER_11_392 ();
 sg13g2_fill_1 FILLER_11_436 ();
 sg13g2_fill_2 FILLER_11_447 ();
 sg13g2_fill_1 FILLER_11_449 ();
 sg13g2_fill_2 FILLER_11_478 ();
 sg13g2_fill_1 FILLER_11_480 ();
 sg13g2_fill_1 FILLER_11_491 ();
 sg13g2_fill_2 FILLER_11_527 ();
 sg13g2_fill_1 FILLER_11_529 ();
 sg13g2_fill_1 FILLER_11_596 ();
 sg13g2_fill_1 FILLER_11_602 ();
 sg13g2_fill_2 FILLER_11_629 ();
 sg13g2_fill_2 FILLER_11_685 ();
 sg13g2_fill_1 FILLER_11_687 ();
 sg13g2_fill_2 FILLER_11_720 ();
 sg13g2_decap_4 FILLER_11_832 ();
 sg13g2_fill_1 FILLER_11_836 ();
 sg13g2_fill_2 FILLER_11_850 ();
 sg13g2_fill_2 FILLER_11_927 ();
 sg13g2_fill_1 FILLER_11_929 ();
 sg13g2_decap_8 FILLER_11_938 ();
 sg13g2_fill_1 FILLER_11_1039 ();
 sg13g2_fill_2 FILLER_11_1075 ();
 sg13g2_fill_1 FILLER_11_1086 ();
 sg13g2_fill_2 FILLER_11_1092 ();
 sg13g2_fill_1 FILLER_11_1231 ();
 sg13g2_fill_2 FILLER_11_1283 ();
 sg13g2_fill_1 FILLER_11_1285 ();
 sg13g2_fill_2 FILLER_11_1300 ();
 sg13g2_fill_1 FILLER_11_1302 ();
 sg13g2_fill_2 FILLER_11_1308 ();
 sg13g2_fill_1 FILLER_11_1310 ();
 sg13g2_fill_2 FILLER_11_1415 ();
 sg13g2_fill_2 FILLER_11_1522 ();
 sg13g2_fill_1 FILLER_11_1524 ();
 sg13g2_fill_2 FILLER_11_1551 ();
 sg13g2_fill_1 FILLER_11_1553 ();
 sg13g2_fill_1 FILLER_11_1585 ();
 sg13g2_fill_1 FILLER_11_1590 ();
 sg13g2_fill_2 FILLER_11_1629 ();
 sg13g2_fill_1 FILLER_11_1631 ();
 sg13g2_fill_2 FILLER_11_1657 ();
 sg13g2_fill_1 FILLER_11_1695 ();
 sg13g2_fill_2 FILLER_11_1766 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_fill_1 FILLER_12_79 ();
 sg13g2_fill_2 FILLER_12_106 ();
 sg13g2_fill_1 FILLER_12_108 ();
 sg13g2_fill_1 FILLER_12_207 ();
 sg13g2_fill_2 FILLER_12_230 ();
 sg13g2_fill_1 FILLER_12_327 ();
 sg13g2_fill_1 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_429 ();
 sg13g2_fill_2 FILLER_12_462 ();
 sg13g2_fill_1 FILLER_12_464 ();
 sg13g2_fill_2 FILLER_12_574 ();
 sg13g2_fill_2 FILLER_12_648 ();
 sg13g2_fill_1 FILLER_12_685 ();
 sg13g2_fill_2 FILLER_12_704 ();
 sg13g2_fill_2 FILLER_12_745 ();
 sg13g2_fill_1 FILLER_12_747 ();
 sg13g2_fill_1 FILLER_12_776 ();
 sg13g2_fill_1 FILLER_12_803 ();
 sg13g2_decap_4 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_918 ();
 sg13g2_fill_2 FILLER_12_932 ();
 sg13g2_fill_1 FILLER_12_934 ();
 sg13g2_fill_2 FILLER_12_993 ();
 sg13g2_fill_2 FILLER_12_1049 ();
 sg13g2_fill_1 FILLER_12_1051 ();
 sg13g2_fill_2 FILLER_12_1103 ();
 sg13g2_fill_1 FILLER_12_1105 ();
 sg13g2_fill_2 FILLER_12_1111 ();
 sg13g2_fill_2 FILLER_12_1153 ();
 sg13g2_fill_1 FILLER_12_1155 ();
 sg13g2_fill_2 FILLER_12_1192 ();
 sg13g2_decap_8 FILLER_12_1264 ();
 sg13g2_decap_8 FILLER_12_1271 ();
 sg13g2_fill_2 FILLER_12_1278 ();
 sg13g2_fill_2 FILLER_12_1288 ();
 sg13g2_fill_1 FILLER_12_1290 ();
 sg13g2_fill_2 FILLER_12_1336 ();
 sg13g2_fill_1 FILLER_12_1338 ();
 sg13g2_fill_1 FILLER_12_1353 ();
 sg13g2_decap_4 FILLER_12_1364 ();
 sg13g2_fill_1 FILLER_12_1447 ();
 sg13g2_fill_2 FILLER_12_1475 ();
 sg13g2_fill_1 FILLER_12_1477 ();
 sg13g2_fill_2 FILLER_12_1528 ();
 sg13g2_fill_1 FILLER_12_1530 ();
 sg13g2_fill_2 FILLER_12_1564 ();
 sg13g2_fill_2 FILLER_12_1602 ();
 sg13g2_fill_1 FILLER_12_1604 ();
 sg13g2_fill_1 FILLER_12_1663 ();
 sg13g2_fill_2 FILLER_12_1747 ();
 sg13g2_fill_1 FILLER_12_1767 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_33 ();
 sg13g2_fill_1 FILLER_13_35 ();
 sg13g2_fill_2 FILLER_13_81 ();
 sg13g2_fill_1 FILLER_13_83 ();
 sg13g2_fill_2 FILLER_13_122 ();
 sg13g2_fill_1 FILLER_13_124 ();
 sg13g2_fill_2 FILLER_13_135 ();
 sg13g2_fill_1 FILLER_13_137 ();
 sg13g2_decap_4 FILLER_13_175 ();
 sg13g2_fill_1 FILLER_13_189 ();
 sg13g2_fill_2 FILLER_13_199 ();
 sg13g2_fill_1 FILLER_13_201 ();
 sg13g2_fill_2 FILLER_13_254 ();
 sg13g2_fill_1 FILLER_13_256 ();
 sg13g2_fill_2 FILLER_13_316 ();
 sg13g2_fill_1 FILLER_13_318 ();
 sg13g2_fill_2 FILLER_13_362 ();
 sg13g2_fill_1 FILLER_13_364 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_fill_1 FILLER_13_441 ();
 sg13g2_fill_2 FILLER_13_461 ();
 sg13g2_fill_2 FILLER_13_482 ();
 sg13g2_decap_4 FILLER_13_497 ();
 sg13g2_fill_2 FILLER_13_501 ();
 sg13g2_fill_2 FILLER_13_529 ();
 sg13g2_fill_2 FILLER_13_622 ();
 sg13g2_fill_2 FILLER_13_637 ();
 sg13g2_fill_1 FILLER_13_639 ();
 sg13g2_fill_2 FILLER_13_650 ();
 sg13g2_fill_1 FILLER_13_671 ();
 sg13g2_fill_1 FILLER_13_730 ();
 sg13g2_fill_1 FILLER_13_783 ();
 sg13g2_fill_1 FILLER_13_807 ();
 sg13g2_fill_2 FILLER_13_828 ();
 sg13g2_decap_4 FILLER_13_853 ();
 sg13g2_fill_2 FILLER_13_857 ();
 sg13g2_decap_4 FILLER_13_869 ();
 sg13g2_fill_1 FILLER_13_873 ();
 sg13g2_fill_1 FILLER_13_884 ();
 sg13g2_fill_2 FILLER_13_919 ();
 sg13g2_fill_2 FILLER_13_930 ();
 sg13g2_fill_2 FILLER_13_942 ();
 sg13g2_fill_2 FILLER_13_964 ();
 sg13g2_fill_1 FILLER_13_1002 ();
 sg13g2_fill_2 FILLER_13_1027 ();
 sg13g2_fill_1 FILLER_13_1029 ();
 sg13g2_decap_8 FILLER_13_1071 ();
 sg13g2_decap_4 FILLER_13_1108 ();
 sg13g2_fill_2 FILLER_13_1151 ();
 sg13g2_fill_1 FILLER_13_1153 ();
 sg13g2_fill_2 FILLER_13_1186 ();
 sg13g2_fill_1 FILLER_13_1277 ();
 sg13g2_fill_2 FILLER_13_1288 ();
 sg13g2_fill_2 FILLER_13_1366 ();
 sg13g2_fill_1 FILLER_13_1402 ();
 sg13g2_fill_2 FILLER_13_1407 ();
 sg13g2_fill_2 FILLER_13_1428 ();
 sg13g2_fill_1 FILLER_13_1430 ();
 sg13g2_fill_2 FILLER_13_1511 ();
 sg13g2_fill_1 FILLER_13_1513 ();
 sg13g2_fill_1 FILLER_13_1536 ();
 sg13g2_fill_1 FILLER_13_1560 ();
 sg13g2_fill_2 FILLER_13_1598 ();
 sg13g2_fill_1 FILLER_13_1614 ();
 sg13g2_fill_1 FILLER_13_1720 ();
 sg13g2_fill_1 FILLER_13_1741 ();
 sg13g2_fill_2 FILLER_14_46 ();
 sg13g2_fill_1 FILLER_14_48 ();
 sg13g2_fill_1 FILLER_14_64 ();
 sg13g2_fill_2 FILLER_14_100 ();
 sg13g2_fill_1 FILLER_14_102 ();
 sg13g2_fill_2 FILLER_14_168 ();
 sg13g2_fill_2 FILLER_14_218 ();
 sg13g2_fill_1 FILLER_14_259 ();
 sg13g2_fill_1 FILLER_14_278 ();
 sg13g2_fill_1 FILLER_14_305 ();
 sg13g2_fill_1 FILLER_14_356 ();
 sg13g2_fill_1 FILLER_14_407 ();
 sg13g2_fill_1 FILLER_14_434 ();
 sg13g2_fill_2 FILLER_14_466 ();
 sg13g2_fill_2 FILLER_14_494 ();
 sg13g2_fill_2 FILLER_14_504 ();
 sg13g2_fill_2 FILLER_14_510 ();
 sg13g2_fill_1 FILLER_14_512 ();
 sg13g2_fill_2 FILLER_14_527 ();
 sg13g2_fill_1 FILLER_14_596 ();
 sg13g2_fill_2 FILLER_14_614 ();
 sg13g2_fill_1 FILLER_14_723 ();
 sg13g2_fill_2 FILLER_14_906 ();
 sg13g2_fill_1 FILLER_14_953 ();
 sg13g2_fill_2 FILLER_14_1018 ();
 sg13g2_fill_2 FILLER_14_1043 ();
 sg13g2_fill_1 FILLER_14_1072 ();
 sg13g2_fill_2 FILLER_14_1077 ();
 sg13g2_fill_1 FILLER_14_1121 ();
 sg13g2_fill_1 FILLER_14_1148 ();
 sg13g2_fill_1 FILLER_14_1159 ();
 sg13g2_fill_2 FILLER_14_1191 ();
 sg13g2_fill_1 FILLER_14_1212 ();
 sg13g2_fill_2 FILLER_14_1240 ();
 sg13g2_fill_1 FILLER_14_1303 ();
 sg13g2_fill_2 FILLER_14_1329 ();
 sg13g2_fill_1 FILLER_14_1349 ();
 sg13g2_fill_1 FILLER_14_1360 ();
 sg13g2_fill_1 FILLER_14_1376 ();
 sg13g2_fill_1 FILLER_14_1406 ();
 sg13g2_fill_2 FILLER_14_1412 ();
 sg13g2_fill_2 FILLER_14_1426 ();
 sg13g2_fill_1 FILLER_14_1464 ();
 sg13g2_fill_2 FILLER_14_1505 ();
 sg13g2_fill_1 FILLER_14_1507 ();
 sg13g2_fill_2 FILLER_14_1512 ();
 sg13g2_fill_1 FILLER_14_1514 ();
 sg13g2_fill_1 FILLER_14_1520 ();
 sg13g2_fill_1 FILLER_14_1530 ();
 sg13g2_fill_1 FILLER_14_1560 ();
 sg13g2_decap_4 FILLER_14_1571 ();
 sg13g2_fill_1 FILLER_14_1575 ();
 sg13g2_fill_2 FILLER_14_1647 ();
 sg13g2_fill_1 FILLER_14_1649 ();
 sg13g2_fill_1 FILLER_14_1660 ();
 sg13g2_fill_2 FILLER_14_1666 ();
 sg13g2_fill_1 FILLER_14_1704 ();
 sg13g2_fill_2 FILLER_14_1736 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_15 ();
 sg13g2_fill_1 FILLER_15_40 ();
 sg13g2_fill_1 FILLER_15_87 ();
 sg13g2_fill_2 FILLER_15_184 ();
 sg13g2_fill_1 FILLER_15_186 ();
 sg13g2_fill_1 FILLER_15_196 ();
 sg13g2_fill_2 FILLER_15_217 ();
 sg13g2_fill_1 FILLER_15_219 ();
 sg13g2_fill_2 FILLER_15_226 ();
 sg13g2_fill_2 FILLER_15_289 ();
 sg13g2_fill_1 FILLER_15_305 ();
 sg13g2_fill_2 FILLER_15_332 ();
 sg13g2_fill_1 FILLER_15_334 ();
 sg13g2_fill_1 FILLER_15_367 ();
 sg13g2_fill_2 FILLER_15_377 ();
 sg13g2_fill_1 FILLER_15_379 ();
 sg13g2_fill_2 FILLER_15_433 ();
 sg13g2_fill_2 FILLER_15_452 ();
 sg13g2_fill_2 FILLER_15_467 ();
 sg13g2_fill_2 FILLER_15_521 ();
 sg13g2_fill_1 FILLER_15_523 ();
 sg13g2_decap_8 FILLER_15_528 ();
 sg13g2_fill_2 FILLER_15_535 ();
 sg13g2_decap_4 FILLER_15_584 ();
 sg13g2_fill_1 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_634 ();
 sg13g2_decap_8 FILLER_15_641 ();
 sg13g2_fill_2 FILLER_15_648 ();
 sg13g2_fill_2 FILLER_15_664 ();
 sg13g2_fill_1 FILLER_15_666 ();
 sg13g2_fill_1 FILLER_15_684 ();
 sg13g2_fill_1 FILLER_15_727 ();
 sg13g2_decap_4 FILLER_15_745 ();
 sg13g2_fill_1 FILLER_15_749 ();
 sg13g2_fill_2 FILLER_15_776 ();
 sg13g2_fill_1 FILLER_15_778 ();
 sg13g2_fill_2 FILLER_15_808 ();
 sg13g2_fill_2 FILLER_15_825 ();
 sg13g2_fill_2 FILLER_15_841 ();
 sg13g2_fill_1 FILLER_15_843 ();
 sg13g2_fill_1 FILLER_15_866 ();
 sg13g2_fill_2 FILLER_15_886 ();
 sg13g2_fill_1 FILLER_15_888 ();
 sg13g2_fill_1 FILLER_15_902 ();
 sg13g2_fill_2 FILLER_15_927 ();
 sg13g2_decap_4 FILLER_15_943 ();
 sg13g2_fill_2 FILLER_15_1009 ();
 sg13g2_decap_8 FILLER_15_1088 ();
 sg13g2_decap_4 FILLER_15_1095 ();
 sg13g2_fill_2 FILLER_15_1183 ();
 sg13g2_fill_1 FILLER_15_1185 ();
 sg13g2_decap_4 FILLER_15_1195 ();
 sg13g2_fill_1 FILLER_15_1251 ();
 sg13g2_decap_4 FILLER_15_1257 ();
 sg13g2_fill_1 FILLER_15_1292 ();
 sg13g2_fill_1 FILLER_15_1319 ();
 sg13g2_fill_2 FILLER_15_1339 ();
 sg13g2_fill_2 FILLER_15_1360 ();
 sg13g2_fill_1 FILLER_15_1362 ();
 sg13g2_decap_4 FILLER_15_1382 ();
 sg13g2_fill_1 FILLER_15_1386 ();
 sg13g2_fill_2 FILLER_15_1429 ();
 sg13g2_fill_1 FILLER_15_1431 ();
 sg13g2_fill_2 FILLER_15_1442 ();
 sg13g2_fill_2 FILLER_15_1485 ();
 sg13g2_fill_2 FILLER_15_1528 ();
 sg13g2_fill_1 FILLER_15_1540 ();
 sg13g2_fill_1 FILLER_15_1547 ();
 sg13g2_fill_1 FILLER_15_1566 ();
 sg13g2_decap_8 FILLER_15_1575 ();
 sg13g2_decap_4 FILLER_15_1582 ();
 sg13g2_fill_1 FILLER_15_1586 ();
 sg13g2_fill_1 FILLER_15_1591 ();
 sg13g2_fill_2 FILLER_15_1610 ();
 sg13g2_fill_2 FILLER_15_1622 ();
 sg13g2_fill_1 FILLER_15_1624 ();
 sg13g2_fill_1 FILLER_15_1661 ();
 sg13g2_fill_2 FILLER_15_1694 ();
 sg13g2_fill_1 FILLER_15_1696 ();
 sg13g2_fill_1 FILLER_15_1730 ();
 sg13g2_fill_1 FILLER_15_1750 ();
 sg13g2_fill_1 FILLER_16_26 ();
 sg13g2_fill_1 FILLER_16_53 ();
 sg13g2_fill_2 FILLER_16_141 ();
 sg13g2_fill_1 FILLER_16_151 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_2 FILLER_16_168 ();
 sg13g2_fill_2 FILLER_16_204 ();
 sg13g2_fill_2 FILLER_16_247 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_fill_2 FILLER_16_323 ();
 sg13g2_fill_2 FILLER_16_396 ();
 sg13g2_fill_1 FILLER_16_398 ();
 sg13g2_fill_1 FILLER_16_446 ();
 sg13g2_decap_4 FILLER_16_539 ();
 sg13g2_fill_2 FILLER_16_574 ();
 sg13g2_fill_1 FILLER_16_598 ();
 sg13g2_decap_8 FILLER_16_650 ();
 sg13g2_fill_2 FILLER_16_688 ();
 sg13g2_fill_1 FILLER_16_690 ();
 sg13g2_fill_2 FILLER_16_722 ();
 sg13g2_fill_1 FILLER_16_734 ();
 sg13g2_decap_4 FILLER_16_752 ();
 sg13g2_fill_1 FILLER_16_756 ();
 sg13g2_fill_1 FILLER_16_767 ();
 sg13g2_fill_2 FILLER_16_829 ();
 sg13g2_fill_2 FILLER_16_876 ();
 sg13g2_fill_1 FILLER_16_878 ();
 sg13g2_fill_2 FILLER_16_905 ();
 sg13g2_fill_1 FILLER_16_938 ();
 sg13g2_fill_2 FILLER_16_965 ();
 sg13g2_fill_2 FILLER_16_1141 ();
 sg13g2_fill_1 FILLER_16_1182 ();
 sg13g2_fill_2 FILLER_16_1192 ();
 sg13g2_fill_2 FILLER_16_1238 ();
 sg13g2_fill_1 FILLER_16_1240 ();
 sg13g2_fill_1 FILLER_16_1267 ();
 sg13g2_fill_1 FILLER_16_1318 ();
 sg13g2_fill_1 FILLER_16_1375 ();
 sg13g2_fill_1 FILLER_16_1402 ();
 sg13g2_decap_4 FILLER_16_1422 ();
 sg13g2_fill_2 FILLER_16_1434 ();
 sg13g2_decap_8 FILLER_16_1558 ();
 sg13g2_fill_2 FILLER_16_1565 ();
 sg13g2_fill_1 FILLER_16_1585 ();
 sg13g2_fill_1 FILLER_16_1616 ();
 sg13g2_fill_2 FILLER_16_1653 ();
 sg13g2_fill_1 FILLER_16_1655 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_47 ();
 sg13g2_fill_2 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_86 ();
 sg13g2_fill_2 FILLER_17_93 ();
 sg13g2_fill_2 FILLER_17_100 ();
 sg13g2_fill_1 FILLER_17_102 ();
 sg13g2_fill_2 FILLER_17_121 ();
 sg13g2_fill_2 FILLER_17_137 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_212 ();
 sg13g2_fill_1 FILLER_17_222 ();
 sg13g2_fill_2 FILLER_17_227 ();
 sg13g2_fill_2 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_288 ();
 sg13g2_fill_2 FILLER_17_391 ();
 sg13g2_fill_2 FILLER_17_410 ();
 sg13g2_decap_8 FILLER_17_429 ();
 sg13g2_fill_1 FILLER_17_477 ();
 sg13g2_fill_1 FILLER_17_514 ();
 sg13g2_decap_4 FILLER_17_574 ();
 sg13g2_fill_1 FILLER_17_578 ();
 sg13g2_decap_8 FILLER_17_645 ();
 sg13g2_fill_1 FILLER_17_652 ();
 sg13g2_decap_4 FILLER_17_657 ();
 sg13g2_fill_2 FILLER_17_661 ();
 sg13g2_fill_2 FILLER_17_676 ();
 sg13g2_fill_1 FILLER_17_678 ();
 sg13g2_fill_2 FILLER_17_824 ();
 sg13g2_fill_1 FILLER_17_826 ();
 sg13g2_fill_2 FILLER_17_842 ();
 sg13g2_decap_4 FILLER_17_884 ();
 sg13g2_fill_2 FILLER_17_888 ();
 sg13g2_fill_2 FILLER_17_894 ();
 sg13g2_fill_2 FILLER_17_900 ();
 sg13g2_fill_2 FILLER_17_916 ();
 sg13g2_fill_1 FILLER_17_918 ();
 sg13g2_fill_1 FILLER_17_938 ();
 sg13g2_fill_2 FILLER_17_963 ();
 sg13g2_fill_1 FILLER_17_965 ();
 sg13g2_fill_1 FILLER_17_982 ();
 sg13g2_fill_1 FILLER_17_1001 ();
 sg13g2_fill_2 FILLER_17_1022 ();
 sg13g2_fill_1 FILLER_17_1024 ();
 sg13g2_fill_1 FILLER_17_1033 ();
 sg13g2_fill_2 FILLER_17_1047 ();
 sg13g2_fill_2 FILLER_17_1098 ();
 sg13g2_fill_2 FILLER_17_1105 ();
 sg13g2_fill_1 FILLER_17_1107 ();
 sg13g2_fill_1 FILLER_17_1117 ();
 sg13g2_fill_1 FILLER_17_1128 ();
 sg13g2_decap_8 FILLER_17_1201 ();
 sg13g2_fill_1 FILLER_17_1234 ();
 sg13g2_fill_1 FILLER_17_1259 ();
 sg13g2_fill_1 FILLER_17_1265 ();
 sg13g2_fill_2 FILLER_17_1295 ();
 sg13g2_fill_2 FILLER_17_1333 ();
 sg13g2_fill_2 FILLER_17_1398 ();
 sg13g2_fill_1 FILLER_17_1418 ();
 sg13g2_fill_1 FILLER_17_1428 ();
 sg13g2_fill_2 FILLER_17_1433 ();
 sg13g2_fill_1 FILLER_17_1448 ();
 sg13g2_fill_2 FILLER_17_1463 ();
 sg13g2_fill_1 FILLER_17_1465 ();
 sg13g2_fill_1 FILLER_17_1533 ();
 sg13g2_decap_4 FILLER_17_1548 ();
 sg13g2_fill_2 FILLER_17_1572 ();
 sg13g2_fill_1 FILLER_17_1574 ();
 sg13g2_fill_2 FILLER_17_1648 ();
 sg13g2_fill_1 FILLER_17_1650 ();
 sg13g2_fill_2 FILLER_17_1665 ();
 sg13g2_fill_1 FILLER_17_1688 ();
 sg13g2_fill_2 FILLER_17_1710 ();
 sg13g2_fill_1 FILLER_17_1712 ();
 sg13g2_fill_2 FILLER_18_26 ();
 sg13g2_fill_1 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_59 ();
 sg13g2_fill_2 FILLER_18_89 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_fill_2 FILLER_18_210 ();
 sg13g2_fill_1 FILLER_18_237 ();
 sg13g2_decap_4 FILLER_18_256 ();
 sg13g2_fill_2 FILLER_18_260 ();
 sg13g2_fill_2 FILLER_18_270 ();
 sg13g2_fill_1 FILLER_18_293 ();
 sg13g2_fill_1 FILLER_18_313 ();
 sg13g2_fill_2 FILLER_18_344 ();
 sg13g2_fill_1 FILLER_18_346 ();
 sg13g2_fill_2 FILLER_18_372 ();
 sg13g2_fill_2 FILLER_18_382 ();
 sg13g2_fill_1 FILLER_18_384 ();
 sg13g2_fill_1 FILLER_18_390 ();
 sg13g2_decap_4 FILLER_18_440 ();
 sg13g2_fill_1 FILLER_18_514 ();
 sg13g2_fill_2 FILLER_18_536 ();
 sg13g2_fill_1 FILLER_18_559 ();
 sg13g2_fill_2 FILLER_18_578 ();
 sg13g2_fill_1 FILLER_18_580 ();
 sg13g2_fill_2 FILLER_18_645 ();
 sg13g2_fill_2 FILLER_18_688 ();
 sg13g2_fill_1 FILLER_18_690 ();
 sg13g2_fill_2 FILLER_18_717 ();
 sg13g2_fill_1 FILLER_18_760 ();
 sg13g2_fill_2 FILLER_18_776 ();
 sg13g2_fill_2 FILLER_18_882 ();
 sg13g2_fill_1 FILLER_18_884 ();
 sg13g2_fill_1 FILLER_18_911 ();
 sg13g2_fill_2 FILLER_18_938 ();
 sg13g2_fill_1 FILLER_18_981 ();
 sg13g2_fill_2 FILLER_18_1018 ();
 sg13g2_fill_1 FILLER_18_1020 ();
 sg13g2_fill_2 FILLER_18_1070 ();
 sg13g2_fill_1 FILLER_18_1072 ();
 sg13g2_decap_4 FILLER_18_1099 ();
 sg13g2_fill_2 FILLER_18_1138 ();
 sg13g2_fill_1 FILLER_18_1140 ();
 sg13g2_fill_1 FILLER_18_1190 ();
 sg13g2_fill_2 FILLER_18_1235 ();
 sg13g2_fill_1 FILLER_18_1237 ();
 sg13g2_fill_2 FILLER_18_1246 ();
 sg13g2_fill_2 FILLER_18_1271 ();
 sg13g2_fill_1 FILLER_18_1273 ();
 sg13g2_fill_2 FILLER_18_1279 ();
 sg13g2_fill_1 FILLER_18_1429 ();
 sg13g2_fill_2 FILLER_18_1479 ();
 sg13g2_fill_1 FILLER_18_1481 ();
 sg13g2_fill_1 FILLER_18_1523 ();
 sg13g2_fill_2 FILLER_18_1529 ();
 sg13g2_fill_2 FILLER_18_1579 ();
 sg13g2_fill_2 FILLER_18_1609 ();
 sg13g2_fill_1 FILLER_18_1721 ();
 sg13g2_fill_2 FILLER_18_1766 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_4 ();
 sg13g2_fill_2 FILLER_19_89 ();
 sg13g2_decap_4 FILLER_19_147 ();
 sg13g2_fill_2 FILLER_19_191 ();
 sg13g2_fill_1 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_243 ();
 sg13g2_decap_8 FILLER_19_250 ();
 sg13g2_fill_2 FILLER_19_257 ();
 sg13g2_fill_2 FILLER_19_277 ();
 sg13g2_fill_2 FILLER_19_322 ();
 sg13g2_fill_1 FILLER_19_324 ();
 sg13g2_fill_2 FILLER_19_335 ();
 sg13g2_fill_1 FILLER_19_337 ();
 sg13g2_fill_2 FILLER_19_388 ();
 sg13g2_fill_2 FILLER_19_420 ();
 sg13g2_fill_1 FILLER_19_448 ();
 sg13g2_fill_2 FILLER_19_472 ();
 sg13g2_fill_1 FILLER_19_474 ();
 sg13g2_fill_2 FILLER_19_506 ();
 sg13g2_fill_1 FILLER_19_513 ();
 sg13g2_fill_1 FILLER_19_519 ();
 sg13g2_fill_1 FILLER_19_541 ();
 sg13g2_fill_2 FILLER_19_639 ();
 sg13g2_fill_1 FILLER_19_641 ();
 sg13g2_fill_2 FILLER_19_658 ();
 sg13g2_decap_4 FILLER_19_726 ();
 sg13g2_fill_1 FILLER_19_753 ();
 sg13g2_fill_2 FILLER_19_780 ();
 sg13g2_fill_1 FILLER_19_782 ();
 sg13g2_fill_2 FILLER_19_837 ();
 sg13g2_fill_1 FILLER_19_839 ();
 sg13g2_fill_2 FILLER_19_868 ();
 sg13g2_fill_1 FILLER_19_870 ();
 sg13g2_fill_2 FILLER_19_877 ();
 sg13g2_fill_1 FILLER_19_889 ();
 sg13g2_decap_4 FILLER_19_948 ();
 sg13g2_fill_2 FILLER_19_952 ();
 sg13g2_decap_8 FILLER_19_972 ();
 sg13g2_fill_1 FILLER_19_979 ();
 sg13g2_fill_2 FILLER_19_984 ();
 sg13g2_fill_2 FILLER_19_1007 ();
 sg13g2_fill_1 FILLER_19_1009 ();
 sg13g2_fill_2 FILLER_19_1031 ();
 sg13g2_fill_1 FILLER_19_1041 ();
 sg13g2_fill_2 FILLER_19_1051 ();
 sg13g2_fill_1 FILLER_19_1066 ();
 sg13g2_decap_8 FILLER_19_1100 ();
 sg13g2_fill_1 FILLER_19_1107 ();
 sg13g2_fill_2 FILLER_19_1138 ();
 sg13g2_fill_1 FILLER_19_1150 ();
 sg13g2_fill_2 FILLER_19_1196 ();
 sg13g2_fill_1 FILLER_19_1198 ();
 sg13g2_fill_2 FILLER_19_1209 ();
 sg13g2_fill_2 FILLER_19_1237 ();
 sg13g2_fill_1 FILLER_19_1239 ();
 sg13g2_fill_1 FILLER_19_1279 ();
 sg13g2_fill_2 FILLER_19_1306 ();
 sg13g2_fill_1 FILLER_19_1308 ();
 sg13g2_fill_2 FILLER_19_1313 ();
 sg13g2_fill_1 FILLER_19_1315 ();
 sg13g2_fill_2 FILLER_19_1320 ();
 sg13g2_fill_1 FILLER_19_1322 ();
 sg13g2_decap_4 FILLER_19_1364 ();
 sg13g2_fill_1 FILLER_19_1368 ();
 sg13g2_fill_2 FILLER_19_1379 ();
 sg13g2_fill_1 FILLER_19_1459 ();
 sg13g2_fill_1 FILLER_19_1561 ();
 sg13g2_fill_2 FILLER_19_1567 ();
 sg13g2_fill_1 FILLER_19_1569 ();
 sg13g2_fill_2 FILLER_19_1616 ();
 sg13g2_fill_2 FILLER_19_1640 ();
 sg13g2_fill_1 FILLER_19_1642 ();
 sg13g2_decap_8 FILLER_19_1666 ();
 sg13g2_decap_4 FILLER_19_1673 ();
 sg13g2_fill_1 FILLER_19_1677 ();
 sg13g2_fill_1 FILLER_19_1696 ();
 sg13g2_fill_2 FILLER_19_1723 ();
 sg13g2_fill_1 FILLER_19_1725 ();
 sg13g2_fill_2 FILLER_20_61 ();
 sg13g2_fill_1 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_128 ();
 sg13g2_fill_1 FILLER_20_142 ();
 sg13g2_fill_2 FILLER_20_158 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_2 FILLER_20_208 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_decap_8 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_230 ();
 sg13g2_fill_2 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_238 ();
 sg13g2_fill_2 FILLER_20_298 ();
 sg13g2_fill_1 FILLER_20_318 ();
 sg13g2_fill_1 FILLER_20_325 ();
 sg13g2_fill_2 FILLER_20_332 ();
 sg13g2_fill_1 FILLER_20_334 ();
 sg13g2_fill_2 FILLER_20_352 ();
 sg13g2_fill_1 FILLER_20_354 ();
 sg13g2_fill_1 FILLER_20_364 ();
 sg13g2_fill_2 FILLER_20_506 ();
 sg13g2_fill_1 FILLER_20_534 ();
 sg13g2_fill_2 FILLER_20_631 ();
 sg13g2_fill_1 FILLER_20_633 ();
 sg13g2_fill_1 FILLER_20_677 ();
 sg13g2_decap_4 FILLER_20_723 ();
 sg13g2_fill_2 FILLER_20_813 ();
 sg13g2_fill_1 FILLER_20_815 ();
 sg13g2_fill_2 FILLER_20_826 ();
 sg13g2_fill_2 FILLER_20_867 ();
 sg13g2_fill_1 FILLER_20_869 ();
 sg13g2_decap_4 FILLER_20_916 ();
 sg13g2_fill_2 FILLER_20_920 ();
 sg13g2_decap_4 FILLER_20_944 ();
 sg13g2_fill_2 FILLER_20_958 ();
 sg13g2_fill_2 FILLER_20_995 ();
 sg13g2_fill_1 FILLER_20_1023 ();
 sg13g2_fill_1 FILLER_20_1047 ();
 sg13g2_fill_1 FILLER_20_1057 ();
 sg13g2_fill_2 FILLER_20_1068 ();
 sg13g2_fill_2 FILLER_20_1111 ();
 sg13g2_fill_1 FILLER_20_1123 ();
 sg13g2_fill_2 FILLER_20_1147 ();
 sg13g2_fill_2 FILLER_20_1202 ();
 sg13g2_decap_4 FILLER_20_1231 ();
 sg13g2_fill_2 FILLER_20_1270 ();
 sg13g2_fill_1 FILLER_20_1331 ();
 sg13g2_fill_1 FILLER_20_1474 ();
 sg13g2_fill_2 FILLER_20_1540 ();
 sg13g2_fill_1 FILLER_20_1617 ();
 sg13g2_fill_2 FILLER_20_1658 ();
 sg13g2_fill_1 FILLER_20_1660 ();
 sg13g2_fill_1 FILLER_20_1671 ();
 sg13g2_fill_1 FILLER_20_1720 ();
 sg13g2_fill_2 FILLER_20_1765 ();
 sg13g2_fill_1 FILLER_20_1767 ();
 sg13g2_fill_2 FILLER_21_61 ();
 sg13g2_fill_2 FILLER_21_78 ();
 sg13g2_fill_2 FILLER_21_89 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_fill_2 FILLER_21_144 ();
 sg13g2_fill_1 FILLER_21_146 ();
 sg13g2_fill_2 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_231 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_fill_2 FILLER_21_344 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_421 ();
 sg13g2_fill_1 FILLER_21_446 ();
 sg13g2_fill_2 FILLER_21_454 ();
 sg13g2_fill_1 FILLER_21_456 ();
 sg13g2_decap_8 FILLER_21_467 ();
 sg13g2_fill_1 FILLER_21_474 ();
 sg13g2_decap_4 FILLER_21_515 ();
 sg13g2_decap_8 FILLER_21_523 ();
 sg13g2_fill_2 FILLER_21_530 ();
 sg13g2_fill_2 FILLER_21_545 ();
 sg13g2_fill_2 FILLER_21_561 ();
 sg13g2_fill_1 FILLER_21_604 ();
 sg13g2_fill_2 FILLER_21_614 ();
 sg13g2_fill_1 FILLER_21_652 ();
 sg13g2_fill_1 FILLER_21_686 ();
 sg13g2_decap_4 FILLER_21_743 ();
 sg13g2_fill_2 FILLER_21_747 ();
 sg13g2_fill_2 FILLER_21_877 ();
 sg13g2_fill_2 FILLER_21_891 ();
 sg13g2_fill_2 FILLER_21_923 ();
 sg13g2_fill_1 FILLER_21_925 ();
 sg13g2_fill_2 FILLER_21_1063 ();
 sg13g2_fill_2 FILLER_21_1095 ();
 sg13g2_fill_1 FILLER_21_1132 ();
 sg13g2_fill_1 FILLER_21_1154 ();
 sg13g2_fill_1 FILLER_21_1182 ();
 sg13g2_fill_1 FILLER_21_1209 ();
 sg13g2_fill_2 FILLER_21_1236 ();
 sg13g2_fill_1 FILLER_21_1312 ();
 sg13g2_fill_1 FILLER_21_1337 ();
 sg13g2_fill_2 FILLER_21_1409 ();
 sg13g2_fill_1 FILLER_21_1411 ();
 sg13g2_decap_4 FILLER_21_1537 ();
 sg13g2_fill_2 FILLER_21_1541 ();
 sg13g2_fill_1 FILLER_21_1569 ();
 sg13g2_fill_2 FILLER_21_1654 ();
 sg13g2_fill_2 FILLER_21_1690 ();
 sg13g2_fill_1 FILLER_21_1692 ();
 sg13g2_fill_2 FILLER_21_1740 ();
 sg13g2_fill_2 FILLER_22_34 ();
 sg13g2_fill_1 FILLER_22_66 ();
 sg13g2_decap_4 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_97 ();
 sg13g2_fill_1 FILLER_22_129 ();
 sg13g2_fill_1 FILLER_22_153 ();
 sg13g2_decap_4 FILLER_22_183 ();
 sg13g2_fill_2 FILLER_22_187 ();
 sg13g2_fill_1 FILLER_22_202 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_225 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_fill_2 FILLER_22_270 ();
 sg13g2_fill_1 FILLER_22_295 ();
 sg13g2_fill_2 FILLER_22_358 ();
 sg13g2_fill_2 FILLER_22_411 ();
 sg13g2_fill_2 FILLER_22_422 ();
 sg13g2_fill_1 FILLER_22_424 ();
 sg13g2_fill_2 FILLER_22_433 ();
 sg13g2_fill_1 FILLER_22_435 ();
 sg13g2_fill_2 FILLER_22_513 ();
 sg13g2_fill_1 FILLER_22_515 ();
 sg13g2_fill_1 FILLER_22_524 ();
 sg13g2_fill_1 FILLER_22_573 ();
 sg13g2_decap_4 FILLER_22_677 ();
 sg13g2_fill_2 FILLER_22_681 ();
 sg13g2_fill_1 FILLER_22_718 ();
 sg13g2_fill_1 FILLER_22_755 ();
 sg13g2_fill_2 FILLER_22_797 ();
 sg13g2_fill_1 FILLER_22_799 ();
 sg13g2_fill_2 FILLER_22_833 ();
 sg13g2_fill_2 FILLER_22_880 ();
 sg13g2_fill_2 FILLER_22_888 ();
 sg13g2_fill_1 FILLER_22_890 ();
 sg13g2_fill_2 FILLER_22_910 ();
 sg13g2_fill_1 FILLER_22_912 ();
 sg13g2_fill_1 FILLER_22_960 ();
 sg13g2_fill_1 FILLER_22_1003 ();
 sg13g2_fill_2 FILLER_22_1044 ();
 sg13g2_fill_1 FILLER_22_1046 ();
 sg13g2_fill_2 FILLER_22_1080 ();
 sg13g2_fill_1 FILLER_22_1082 ();
 sg13g2_decap_4 FILLER_22_1109 ();
 sg13g2_fill_1 FILLER_22_1153 ();
 sg13g2_fill_1 FILLER_22_1184 ();
 sg13g2_fill_1 FILLER_22_1198 ();
 sg13g2_fill_2 FILLER_22_1212 ();
 sg13g2_fill_2 FILLER_22_1224 ();
 sg13g2_fill_1 FILLER_22_1286 ();
 sg13g2_decap_8 FILLER_22_1323 ();
 sg13g2_fill_1 FILLER_22_1330 ();
 sg13g2_fill_2 FILLER_22_1360 ();
 sg13g2_fill_1 FILLER_22_1371 ();
 sg13g2_fill_2 FILLER_22_1387 ();
 sg13g2_fill_1 FILLER_22_1399 ();
 sg13g2_fill_2 FILLER_22_1433 ();
 sg13g2_decap_4 FILLER_22_1555 ();
 sg13g2_fill_1 FILLER_22_1578 ();
 sg13g2_decap_4 FILLER_22_1615 ();
 sg13g2_fill_2 FILLER_22_1619 ();
 sg13g2_fill_1 FILLER_22_1640 ();
 sg13g2_fill_2 FILLER_22_1651 ();
 sg13g2_fill_1 FILLER_22_1658 ();
 sg13g2_fill_1 FILLER_22_1664 ();
 sg13g2_fill_2 FILLER_22_1698 ();
 sg13g2_fill_1 FILLER_22_1700 ();
 sg13g2_fill_2 FILLER_22_1710 ();
 sg13g2_fill_2 FILLER_22_1725 ();
 sg13g2_fill_1 FILLER_22_1727 ();
 sg13g2_fill_2 FILLER_22_1766 ();
 sg13g2_fill_1 FILLER_23_26 ();
 sg13g2_fill_1 FILLER_23_37 ();
 sg13g2_fill_2 FILLER_23_66 ();
 sg13g2_fill_1 FILLER_23_68 ();
 sg13g2_fill_1 FILLER_23_108 ();
 sg13g2_decap_8 FILLER_23_113 ();
 sg13g2_fill_2 FILLER_23_120 ();
 sg13g2_fill_1 FILLER_23_122 ();
 sg13g2_decap_4 FILLER_23_154 ();
 sg13g2_fill_1 FILLER_23_158 ();
 sg13g2_decap_4 FILLER_23_208 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_342 ();
 sg13g2_fill_1 FILLER_23_378 ();
 sg13g2_fill_2 FILLER_23_397 ();
 sg13g2_fill_1 FILLER_23_404 ();
 sg13g2_fill_2 FILLER_23_449 ();
 sg13g2_fill_1 FILLER_23_460 ();
 sg13g2_fill_2 FILLER_23_503 ();
 sg13g2_fill_2 FILLER_23_541 ();
 sg13g2_fill_2 FILLER_23_579 ();
 sg13g2_fill_1 FILLER_23_581 ();
 sg13g2_fill_2 FILLER_23_592 ();
 sg13g2_fill_1 FILLER_23_594 ();
 sg13g2_fill_2 FILLER_23_671 ();
 sg13g2_fill_1 FILLER_23_673 ();
 sg13g2_fill_2 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_755 ();
 sg13g2_fill_2 FILLER_23_762 ();
 sg13g2_fill_1 FILLER_23_798 ();
 sg13g2_fill_2 FILLER_23_846 ();
 sg13g2_fill_2 FILLER_23_882 ();
 sg13g2_fill_2 FILLER_23_950 ();
 sg13g2_fill_1 FILLER_23_952 ();
 sg13g2_fill_1 FILLER_23_1095 ();
 sg13g2_fill_1 FILLER_23_1155 ();
 sg13g2_fill_2 FILLER_23_1166 ();
 sg13g2_fill_1 FILLER_23_1217 ();
 sg13g2_fill_1 FILLER_23_1273 ();
 sg13g2_fill_2 FILLER_23_1318 ();
 sg13g2_fill_2 FILLER_23_1389 ();
 sg13g2_fill_2 FILLER_23_1482 ();
 sg13g2_fill_1 FILLER_23_1484 ();
 sg13g2_decap_8 FILLER_23_1531 ();
 sg13g2_fill_1 FILLER_23_1538 ();
 sg13g2_fill_2 FILLER_23_1552 ();
 sg13g2_fill_1 FILLER_23_1558 ();
 sg13g2_fill_1 FILLER_23_1580 ();
 sg13g2_fill_1 FILLER_23_1615 ();
 sg13g2_fill_2 FILLER_23_1650 ();
 sg13g2_fill_2 FILLER_23_1679 ();
 sg13g2_fill_1 FILLER_23_1738 ();
 sg13g2_fill_2 FILLER_23_1765 ();
 sg13g2_fill_1 FILLER_23_1767 ();
 sg13g2_fill_2 FILLER_24_26 ();
 sg13g2_fill_2 FILLER_24_82 ();
 sg13g2_fill_1 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_142 ();
 sg13g2_decap_4 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_184 ();
 sg13g2_fill_2 FILLER_24_242 ();
 sg13g2_fill_1 FILLER_24_244 ();
 sg13g2_fill_1 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_311 ();
 sg13g2_fill_2 FILLER_24_338 ();
 sg13g2_fill_1 FILLER_24_380 ();
 sg13g2_fill_2 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_403 ();
 sg13g2_decap_4 FILLER_24_446 ();
 sg13g2_fill_2 FILLER_24_510 ();
 sg13g2_fill_1 FILLER_24_512 ();
 sg13g2_fill_2 FILLER_24_573 ();
 sg13g2_fill_2 FILLER_24_600 ();
 sg13g2_fill_2 FILLER_24_641 ();
 sg13g2_fill_2 FILLER_24_650 ();
 sg13g2_fill_2 FILLER_24_665 ();
 sg13g2_fill_2 FILLER_24_693 ();
 sg13g2_fill_1 FILLER_24_695 ();
 sg13g2_fill_2 FILLER_24_731 ();
 sg13g2_fill_1 FILLER_24_759 ();
 sg13g2_fill_2 FILLER_24_817 ();
 sg13g2_fill_2 FILLER_24_866 ();
 sg13g2_fill_1 FILLER_24_868 ();
 sg13g2_decap_4 FILLER_24_888 ();
 sg13g2_decap_4 FILLER_24_917 ();
 sg13g2_fill_1 FILLER_24_921 ();
 sg13g2_fill_2 FILLER_24_931 ();
 sg13g2_fill_2 FILLER_24_947 ();
 sg13g2_fill_1 FILLER_24_949 ();
 sg13g2_fill_2 FILLER_24_976 ();
 sg13g2_fill_2 FILLER_24_993 ();
 sg13g2_fill_2 FILLER_24_1028 ();
 sg13g2_fill_1 FILLER_24_1030 ();
 sg13g2_fill_2 FILLER_24_1045 ();
 sg13g2_fill_1 FILLER_24_1117 ();
 sg13g2_fill_1 FILLER_24_1200 ();
 sg13g2_fill_2 FILLER_24_1229 ();
 sg13g2_fill_1 FILLER_24_1257 ();
 sg13g2_decap_4 FILLER_24_1283 ();
 sg13g2_fill_2 FILLER_24_1287 ();
 sg13g2_fill_2 FILLER_24_1335 ();
 sg13g2_fill_1 FILLER_24_1337 ();
 sg13g2_fill_1 FILLER_24_1363 ();
 sg13g2_fill_2 FILLER_24_1434 ();
 sg13g2_fill_2 FILLER_24_1445 ();
 sg13g2_fill_1 FILLER_24_1447 ();
 sg13g2_fill_2 FILLER_24_1454 ();
 sg13g2_fill_2 FILLER_24_1482 ();
 sg13g2_fill_1 FILLER_24_1508 ();
 sg13g2_decap_4 FILLER_24_1535 ();
 sg13g2_decap_4 FILLER_24_1554 ();
 sg13g2_fill_1 FILLER_24_1558 ();
 sg13g2_fill_1 FILLER_24_1575 ();
 sg13g2_fill_2 FILLER_24_1586 ();
 sg13g2_fill_1 FILLER_24_1588 ();
 sg13g2_fill_2 FILLER_24_1633 ();
 sg13g2_fill_1 FILLER_24_1635 ();
 sg13g2_fill_1 FILLER_24_1660 ();
 sg13g2_fill_1 FILLER_24_1691 ();
 sg13g2_fill_2 FILLER_24_1728 ();
 sg13g2_fill_1 FILLER_24_1730 ();
 sg13g2_fill_1 FILLER_24_1741 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_2 FILLER_25_41 ();
 sg13g2_decap_4 FILLER_25_146 ();
 sg13g2_fill_2 FILLER_25_150 ();
 sg13g2_fill_2 FILLER_25_178 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_fill_2 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_317 ();
 sg13g2_fill_2 FILLER_25_345 ();
 sg13g2_fill_1 FILLER_25_347 ();
 sg13g2_decap_4 FILLER_25_465 ();
 sg13g2_fill_2 FILLER_25_657 ();
 sg13g2_decap_4 FILLER_25_669 ();
 sg13g2_fill_2 FILLER_25_686 ();
 sg13g2_fill_1 FILLER_25_717 ();
 sg13g2_fill_1 FILLER_25_758 ();
 sg13g2_fill_2 FILLER_25_764 ();
 sg13g2_fill_1 FILLER_25_788 ();
 sg13g2_fill_2 FILLER_25_821 ();
 sg13g2_fill_1 FILLER_25_823 ();
 sg13g2_decap_4 FILLER_25_910 ();
 sg13g2_fill_1 FILLER_25_914 ();
 sg13g2_fill_1 FILLER_25_1079 ();
 sg13g2_fill_1 FILLER_25_1125 ();
 sg13g2_fill_2 FILLER_25_1139 ();
 sg13g2_fill_1 FILLER_25_1141 ();
 sg13g2_fill_2 FILLER_25_1167 ();
 sg13g2_fill_1 FILLER_25_1169 ();
 sg13g2_decap_4 FILLER_25_1183 ();
 sg13g2_fill_2 FILLER_25_1266 ();
 sg13g2_fill_1 FILLER_25_1268 ();
 sg13g2_fill_1 FILLER_25_1364 ();
 sg13g2_fill_2 FILLER_25_1453 ();
 sg13g2_fill_1 FILLER_25_1455 ();
 sg13g2_fill_1 FILLER_25_1534 ();
 sg13g2_decap_4 FILLER_25_1540 ();
 sg13g2_fill_1 FILLER_25_1544 ();
 sg13g2_fill_2 FILLER_25_1576 ();
 sg13g2_fill_1 FILLER_25_1604 ();
 sg13g2_fill_2 FILLER_25_1610 ();
 sg13g2_fill_1 FILLER_25_1653 ();
 sg13g2_fill_1 FILLER_25_1694 ();
 sg13g2_fill_1 FILLER_25_1767 ();
 sg13g2_fill_2 FILLER_26_31 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_fill_2 FILLER_26_60 ();
 sg13g2_fill_1 FILLER_26_88 ();
 sg13g2_fill_2 FILLER_26_143 ();
 sg13g2_fill_1 FILLER_26_145 ();
 sg13g2_fill_2 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_192 ();
 sg13g2_fill_1 FILLER_26_194 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_fill_2 FILLER_26_289 ();
 sg13g2_fill_1 FILLER_26_328 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_fill_2 FILLER_26_342 ();
 sg13g2_fill_2 FILLER_26_349 ();
 sg13g2_fill_1 FILLER_26_351 ();
 sg13g2_fill_1 FILLER_26_405 ();
 sg13g2_fill_2 FILLER_26_432 ();
 sg13g2_fill_2 FILLER_26_443 ();
 sg13g2_fill_1 FILLER_26_445 ();
 sg13g2_decap_8 FILLER_26_450 ();
 sg13g2_fill_2 FILLER_26_526 ();
 sg13g2_fill_1 FILLER_26_528 ();
 sg13g2_fill_1 FILLER_26_659 ();
 sg13g2_fill_2 FILLER_26_691 ();
 sg13g2_fill_2 FILLER_26_728 ();
 sg13g2_fill_2 FILLER_26_744 ();
 sg13g2_fill_2 FILLER_26_770 ();
 sg13g2_fill_1 FILLER_26_772 ();
 sg13g2_fill_2 FILLER_26_830 ();
 sg13g2_fill_1 FILLER_26_832 ();
 sg13g2_decap_4 FILLER_26_869 ();
 sg13g2_fill_2 FILLER_26_887 ();
 sg13g2_fill_1 FILLER_26_889 ();
 sg13g2_fill_2 FILLER_26_903 ();
 sg13g2_decap_8 FILLER_26_911 ();
 sg13g2_decap_8 FILLER_26_918 ();
 sg13g2_fill_1 FILLER_26_925 ();
 sg13g2_fill_1 FILLER_26_930 ();
 sg13g2_decap_4 FILLER_26_940 ();
 sg13g2_fill_1 FILLER_26_944 ();
 sg13g2_fill_1 FILLER_26_986 ();
 sg13g2_fill_2 FILLER_26_1004 ();
 sg13g2_fill_1 FILLER_26_1026 ();
 sg13g2_fill_2 FILLER_26_1084 ();
 sg13g2_fill_1 FILLER_26_1086 ();
 sg13g2_fill_1 FILLER_26_1122 ();
 sg13g2_fill_1 FILLER_26_1153 ();
 sg13g2_decap_8 FILLER_26_1250 ();
 sg13g2_fill_1 FILLER_26_1257 ();
 sg13g2_fill_2 FILLER_26_1267 ();
 sg13g2_fill_2 FILLER_26_1284 ();
 sg13g2_fill_1 FILLER_26_1286 ();
 sg13g2_fill_2 FILLER_26_1296 ();
 sg13g2_fill_2 FILLER_26_1346 ();
 sg13g2_fill_2 FILLER_26_1371 ();
 sg13g2_fill_2 FILLER_26_1405 ();
 sg13g2_fill_1 FILLER_26_1407 ();
 sg13g2_fill_2 FILLER_26_1429 ();
 sg13g2_fill_2 FILLER_26_1441 ();
 sg13g2_fill_1 FILLER_26_1534 ();
 sg13g2_fill_2 FILLER_26_1560 ();
 sg13g2_fill_1 FILLER_26_1624 ();
 sg13g2_fill_2 FILLER_26_1652 ();
 sg13g2_fill_1 FILLER_26_1654 ();
 sg13g2_fill_1 FILLER_26_1668 ();
 sg13g2_fill_2 FILLER_26_1720 ();
 sg13g2_fill_1 FILLER_26_1722 ();
 sg13g2_fill_1 FILLER_26_1728 ();
 sg13g2_fill_1 FILLER_26_1767 ();
 sg13g2_fill_2 FILLER_27_50 ();
 sg13g2_fill_1 FILLER_27_159 ();
 sg13g2_fill_2 FILLER_27_170 ();
 sg13g2_fill_1 FILLER_27_172 ();
 sg13g2_fill_2 FILLER_27_206 ();
 sg13g2_fill_1 FILLER_27_276 ();
 sg13g2_fill_1 FILLER_27_291 ();
 sg13g2_fill_2 FILLER_27_307 ();
 sg13g2_fill_2 FILLER_27_371 ();
 sg13g2_fill_2 FILLER_27_411 ();
 sg13g2_decap_4 FILLER_27_439 ();
 sg13g2_fill_1 FILLER_27_443 ();
 sg13g2_fill_2 FILLER_27_480 ();
 sg13g2_fill_1 FILLER_27_482 ();
 sg13g2_fill_2 FILLER_27_596 ();
 sg13g2_fill_1 FILLER_27_598 ();
 sg13g2_fill_2 FILLER_27_630 ();
 sg13g2_fill_1 FILLER_27_632 ();
 sg13g2_fill_2 FILLER_27_664 ();
 sg13g2_fill_1 FILLER_27_680 ();
 sg13g2_fill_2 FILLER_27_695 ();
 sg13g2_fill_1 FILLER_27_697 ();
 sg13g2_fill_2 FILLER_27_717 ();
 sg13g2_fill_1 FILLER_27_779 ();
 sg13g2_fill_2 FILLER_27_789 ();
 sg13g2_fill_1 FILLER_27_791 ();
 sg13g2_fill_1 FILLER_27_817 ();
 sg13g2_fill_2 FILLER_27_842 ();
 sg13g2_fill_1 FILLER_27_880 ();
 sg13g2_fill_2 FILLER_27_933 ();
 sg13g2_fill_1 FILLER_27_935 ();
 sg13g2_fill_1 FILLER_27_951 ();
 sg13g2_fill_2 FILLER_27_1039 ();
 sg13g2_fill_1 FILLER_27_1046 ();
 sg13g2_fill_1 FILLER_27_1066 ();
 sg13g2_fill_1 FILLER_27_1090 ();
 sg13g2_fill_2 FILLER_27_1127 ();
 sg13g2_fill_1 FILLER_27_1129 ();
 sg13g2_decap_8 FILLER_27_1179 ();
 sg13g2_fill_1 FILLER_27_1186 ();
 sg13g2_fill_2 FILLER_27_1300 ();
 sg13g2_fill_1 FILLER_27_1302 ();
 sg13g2_fill_1 FILLER_27_1381 ();
 sg13g2_fill_2 FILLER_27_1469 ();
 sg13g2_fill_1 FILLER_27_1471 ();
 sg13g2_fill_1 FILLER_27_1490 ();
 sg13g2_fill_2 FILLER_27_1525 ();
 sg13g2_fill_1 FILLER_27_1527 ();
 sg13g2_fill_1 FILLER_27_1554 ();
 sg13g2_fill_1 FILLER_27_1608 ();
 sg13g2_fill_2 FILLER_27_1619 ();
 sg13g2_fill_2 FILLER_27_1631 ();
 sg13g2_fill_1 FILLER_27_1633 ();
 sg13g2_fill_1 FILLER_27_1656 ();
 sg13g2_fill_2 FILLER_27_1687 ();
 sg13g2_fill_1 FILLER_27_1689 ();
 sg13g2_fill_2 FILLER_27_1720 ();
 sg13g2_fill_1 FILLER_27_1722 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_15 ();
 sg13g2_fill_2 FILLER_28_51 ();
 sg13g2_fill_1 FILLER_28_53 ();
 sg13g2_fill_1 FILLER_28_64 ();
 sg13g2_decap_8 FILLER_28_86 ();
 sg13g2_fill_1 FILLER_28_93 ();
 sg13g2_fill_2 FILLER_28_123 ();
 sg13g2_fill_1 FILLER_28_196 ();
 sg13g2_fill_2 FILLER_28_255 ();
 sg13g2_fill_1 FILLER_28_352 ();
 sg13g2_fill_2 FILLER_28_422 ();
 sg13g2_decap_8 FILLER_28_432 ();
 sg13g2_fill_1 FILLER_28_470 ();
 sg13g2_fill_1 FILLER_28_543 ();
 sg13g2_fill_2 FILLER_28_641 ();
 sg13g2_fill_1 FILLER_28_643 ();
 sg13g2_fill_2 FILLER_28_670 ();
 sg13g2_fill_1 FILLER_28_703 ();
 sg13g2_fill_1 FILLER_28_730 ();
 sg13g2_fill_2 FILLER_28_796 ();
 sg13g2_fill_2 FILLER_28_824 ();
 sg13g2_fill_2 FILLER_28_861 ();
 sg13g2_fill_1 FILLER_28_863 ();
 sg13g2_fill_2 FILLER_28_873 ();
 sg13g2_fill_1 FILLER_28_875 ();
 sg13g2_decap_8 FILLER_28_933 ();
 sg13g2_fill_1 FILLER_28_982 ();
 sg13g2_fill_2 FILLER_28_1155 ();
 sg13g2_fill_1 FILLER_28_1157 ();
 sg13g2_fill_2 FILLER_28_1189 ();
 sg13g2_fill_2 FILLER_28_1217 ();
 sg13g2_fill_1 FILLER_28_1219 ();
 sg13g2_fill_1 FILLER_28_1246 ();
 sg13g2_decap_4 FILLER_28_1273 ();
 sg13g2_fill_1 FILLER_28_1306 ();
 sg13g2_decap_4 FILLER_28_1326 ();
 sg13g2_fill_1 FILLER_28_1330 ();
 sg13g2_decap_4 FILLER_28_1339 ();
 sg13g2_fill_1 FILLER_28_1343 ();
 sg13g2_fill_1 FILLER_28_1397 ();
 sg13g2_fill_2 FILLER_28_1411 ();
 sg13g2_fill_1 FILLER_28_1413 ();
 sg13g2_fill_2 FILLER_28_1441 ();
 sg13g2_fill_1 FILLER_28_1443 ();
 sg13g2_fill_2 FILLER_28_1472 ();
 sg13g2_fill_1 FILLER_28_1474 ();
 sg13g2_fill_2 FILLER_28_1485 ();
 sg13g2_fill_2 FILLER_28_1521 ();
 sg13g2_fill_1 FILLER_28_1523 ();
 sg13g2_fill_2 FILLER_28_1584 ();
 sg13g2_fill_1 FILLER_28_1586 ();
 sg13g2_fill_1 FILLER_28_1613 ();
 sg13g2_fill_1 FILLER_28_1650 ();
 sg13g2_decap_4 FILLER_28_1708 ();
 sg13g2_fill_1 FILLER_28_1712 ();
 sg13g2_fill_2 FILLER_28_1723 ();
 sg13g2_fill_2 FILLER_28_1766 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_decap_4 FILLER_29_50 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_fill_1 FILLER_29_71 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_fill_1 FILLER_29_154 ();
 sg13g2_fill_2 FILLER_29_165 ();
 sg13g2_fill_2 FILLER_29_186 ();
 sg13g2_fill_2 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_fill_2 FILLER_29_237 ();
 sg13g2_fill_1 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_fill_1 FILLER_29_286 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_fill_2 FILLER_29_378 ();
 sg13g2_fill_2 FILLER_29_388 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_fill_2 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_430 ();
 sg13g2_fill_1 FILLER_29_432 ();
 sg13g2_fill_1 FILLER_29_469 ();
 sg13g2_fill_1 FILLER_29_494 ();
 sg13g2_fill_2 FILLER_29_581 ();
 sg13g2_fill_1 FILLER_29_583 ();
 sg13g2_fill_2 FILLER_29_615 ();
 sg13g2_fill_1 FILLER_29_617 ();
 sg13g2_fill_2 FILLER_29_662 ();
 sg13g2_decap_4 FILLER_29_672 ();
 sg13g2_fill_1 FILLER_29_676 ();
 sg13g2_fill_1 FILLER_29_682 ();
 sg13g2_fill_1 FILLER_29_687 ();
 sg13g2_fill_2 FILLER_29_693 ();
 sg13g2_fill_2 FILLER_29_703 ();
 sg13g2_fill_1 FILLER_29_705 ();
 sg13g2_fill_2 FILLER_29_720 ();
 sg13g2_fill_1 FILLER_29_735 ();
 sg13g2_decap_4 FILLER_29_812 ();
 sg13g2_fill_1 FILLER_29_895 ();
 sg13g2_fill_1 FILLER_29_968 ();
 sg13g2_fill_2 FILLER_29_979 ();
 sg13g2_fill_2 FILLER_29_1019 ();
 sg13g2_fill_1 FILLER_29_1021 ();
 sg13g2_fill_2 FILLER_29_1037 ();
 sg13g2_fill_1 FILLER_29_1039 ();
 sg13g2_fill_2 FILLER_29_1055 ();
 sg13g2_fill_1 FILLER_29_1057 ();
 sg13g2_decap_8 FILLER_29_1104 ();
 sg13g2_fill_2 FILLER_29_1141 ();
 sg13g2_fill_1 FILLER_29_1230 ();
 sg13g2_fill_2 FILLER_29_1240 ();
 sg13g2_fill_1 FILLER_29_1242 ();
 sg13g2_fill_1 FILLER_29_1256 ();
 sg13g2_decap_8 FILLER_29_1274 ();
 sg13g2_decap_4 FILLER_29_1281 ();
 sg13g2_fill_2 FILLER_29_1285 ();
 sg13g2_fill_2 FILLER_29_1323 ();
 sg13g2_fill_1 FILLER_29_1325 ();
 sg13g2_decap_4 FILLER_29_1344 ();
 sg13g2_fill_2 FILLER_29_1417 ();
 sg13g2_fill_1 FILLER_29_1428 ();
 sg13g2_fill_2 FILLER_29_1439 ();
 sg13g2_fill_1 FILLER_29_1441 ();
 sg13g2_fill_2 FILLER_29_1456 ();
 sg13g2_fill_2 FILLER_29_1493 ();
 sg13g2_fill_2 FILLER_29_1526 ();
 sg13g2_fill_2 FILLER_29_1557 ();
 sg13g2_fill_1 FILLER_29_1559 ();
 sg13g2_fill_2 FILLER_29_1584 ();
 sg13g2_fill_2 FILLER_29_1658 ();
 sg13g2_fill_1 FILLER_29_1670 ();
 sg13g2_fill_2 FILLER_29_1680 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_103 ();
 sg13g2_fill_1 FILLER_30_105 ();
 sg13g2_fill_2 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_131 ();
 sg13g2_fill_2 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_212 ();
 sg13g2_fill_2 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_311 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_fill_2 FILLER_30_345 ();
 sg13g2_decap_4 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_428 ();
 sg13g2_fill_1 FILLER_30_435 ();
 sg13g2_fill_1 FILLER_30_468 ();
 sg13g2_fill_1 FILLER_30_567 ();
 sg13g2_fill_1 FILLER_30_582 ();
 sg13g2_fill_1 FILLER_30_606 ();
 sg13g2_fill_1 FILLER_30_653 ();
 sg13g2_decap_4 FILLER_30_664 ();
 sg13g2_fill_1 FILLER_30_668 ();
 sg13g2_fill_2 FILLER_30_686 ();
 sg13g2_fill_1 FILLER_30_688 ();
 sg13g2_fill_2 FILLER_30_734 ();
 sg13g2_fill_1 FILLER_30_736 ();
 sg13g2_fill_1 FILLER_30_824 ();
 sg13g2_fill_2 FILLER_30_856 ();
 sg13g2_fill_1 FILLER_30_858 ();
 sg13g2_decap_4 FILLER_30_869 ();
 sg13g2_fill_1 FILLER_30_873 ();
 sg13g2_fill_2 FILLER_30_883 ();
 sg13g2_fill_1 FILLER_30_943 ();
 sg13g2_fill_2 FILLER_30_977 ();
 sg13g2_fill_2 FILLER_30_1010 ();
 sg13g2_fill_1 FILLER_30_1012 ();
 sg13g2_fill_2 FILLER_30_1044 ();
 sg13g2_fill_1 FILLER_30_1103 ();
 sg13g2_decap_8 FILLER_30_1112 ();
 sg13g2_fill_1 FILLER_30_1119 ();
 sg13g2_fill_2 FILLER_30_1215 ();
 sg13g2_fill_1 FILLER_30_1217 ();
 sg13g2_fill_1 FILLER_30_1244 ();
 sg13g2_decap_4 FILLER_30_1285 ();
 sg13g2_fill_2 FILLER_30_1289 ();
 sg13g2_fill_2 FILLER_30_1301 ();
 sg13g2_fill_1 FILLER_30_1393 ();
 sg13g2_fill_1 FILLER_30_1398 ();
 sg13g2_fill_1 FILLER_30_1471 ();
 sg13g2_decap_4 FILLER_30_1512 ();
 sg13g2_fill_1 FILLER_30_1516 ();
 sg13g2_fill_1 FILLER_30_1633 ();
 sg13g2_fill_2 FILLER_30_1648 ();
 sg13g2_fill_1 FILLER_30_1650 ();
 sg13g2_fill_2 FILLER_30_1687 ();
 sg13g2_fill_1 FILLER_31_35 ();
 sg13g2_decap_4 FILLER_31_80 ();
 sg13g2_fill_2 FILLER_31_129 ();
 sg13g2_fill_1 FILLER_31_131 ();
 sg13g2_fill_1 FILLER_31_137 ();
 sg13g2_fill_2 FILLER_31_157 ();
 sg13g2_fill_1 FILLER_31_159 ();
 sg13g2_fill_1 FILLER_31_197 ();
 sg13g2_fill_2 FILLER_31_208 ();
 sg13g2_fill_1 FILLER_31_210 ();
 sg13g2_fill_2 FILLER_31_230 ();
 sg13g2_fill_1 FILLER_31_232 ();
 sg13g2_fill_2 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_356 ();
 sg13g2_fill_2 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_408 ();
 sg13g2_fill_1 FILLER_31_412 ();
 sg13g2_decap_4 FILLER_31_421 ();
 sg13g2_fill_2 FILLER_31_425 ();
 sg13g2_fill_2 FILLER_31_473 ();
 sg13g2_fill_2 FILLER_31_549 ();
 sg13g2_fill_2 FILLER_31_575 ();
 sg13g2_fill_1 FILLER_31_577 ();
 sg13g2_fill_1 FILLER_31_614 ();
 sg13g2_decap_4 FILLER_31_649 ();
 sg13g2_fill_1 FILLER_31_653 ();
 sg13g2_fill_2 FILLER_31_706 ();
 sg13g2_fill_1 FILLER_31_712 ();
 sg13g2_fill_2 FILLER_31_759 ();
 sg13g2_fill_2 FILLER_31_776 ();
 sg13g2_fill_1 FILLER_31_792 ();
 sg13g2_fill_2 FILLER_31_807 ();
 sg13g2_fill_1 FILLER_31_809 ();
 sg13g2_fill_2 FILLER_31_815 ();
 sg13g2_fill_2 FILLER_31_881 ();
 sg13g2_fill_2 FILLER_31_896 ();
 sg13g2_fill_1 FILLER_31_898 ();
 sg13g2_decap_4 FILLER_31_906 ();
 sg13g2_fill_1 FILLER_31_910 ();
 sg13g2_fill_1 FILLER_31_941 ();
 sg13g2_decap_8 FILLER_31_961 ();
 sg13g2_fill_2 FILLER_31_973 ();
 sg13g2_fill_1 FILLER_31_1039 ();
 sg13g2_fill_2 FILLER_31_1055 ();
 sg13g2_fill_1 FILLER_31_1057 ();
 sg13g2_fill_2 FILLER_31_1077 ();
 sg13g2_fill_2 FILLER_31_1136 ();
 sg13g2_fill_1 FILLER_31_1138 ();
 sg13g2_fill_1 FILLER_31_1192 ();
 sg13g2_fill_2 FILLER_31_1260 ();
 sg13g2_fill_1 FILLER_31_1280 ();
 sg13g2_decap_8 FILLER_31_1321 ();
 sg13g2_decap_8 FILLER_31_1328 ();
 sg13g2_decap_8 FILLER_31_1335 ();
 sg13g2_fill_2 FILLER_31_1342 ();
 sg13g2_fill_1 FILLER_31_1344 ();
 sg13g2_fill_2 FILLER_31_1359 ();
 sg13g2_decap_4 FILLER_31_1397 ();
 sg13g2_fill_2 FILLER_31_1401 ();
 sg13g2_fill_2 FILLER_31_1412 ();
 sg13g2_fill_2 FILLER_31_1423 ();
 sg13g2_fill_2 FILLER_31_1435 ();
 sg13g2_fill_1 FILLER_31_1437 ();
 sg13g2_fill_2 FILLER_31_1451 ();
 sg13g2_fill_1 FILLER_31_1458 ();
 sg13g2_decap_4 FILLER_31_1477 ();
 sg13g2_fill_2 FILLER_31_1513 ();
 sg13g2_fill_2 FILLER_31_1560 ();
 sg13g2_fill_1 FILLER_31_1575 ();
 sg13g2_fill_2 FILLER_31_1595 ();
 sg13g2_fill_2 FILLER_31_1623 ();
 sg13g2_fill_1 FILLER_31_1625 ();
 sg13g2_fill_1 FILLER_31_1686 ();
 sg13g2_fill_1 FILLER_31_1711 ();
 sg13g2_fill_2 FILLER_31_1717 ();
 sg13g2_fill_1 FILLER_31_1719 ();
 sg13g2_fill_1 FILLER_31_1739 ();
 sg13g2_fill_1 FILLER_31_1767 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_11 ();
 sg13g2_fill_2 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_111 ();
 sg13g2_fill_1 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_279 ();
 sg13g2_fill_1 FILLER_32_288 ();
 sg13g2_fill_2 FILLER_32_353 ();
 sg13g2_fill_2 FILLER_32_375 ();
 sg13g2_fill_2 FILLER_32_403 ();
 sg13g2_fill_1 FILLER_32_405 ();
 sg13g2_fill_2 FILLER_32_414 ();
 sg13g2_decap_4 FILLER_32_432 ();
 sg13g2_fill_1 FILLER_32_436 ();
 sg13g2_decap_4 FILLER_32_441 ();
 sg13g2_fill_2 FILLER_32_475 ();
 sg13g2_fill_2 FILLER_32_504 ();
 sg13g2_fill_2 FILLER_32_530 ();
 sg13g2_fill_2 FILLER_32_542 ();
 sg13g2_fill_1 FILLER_32_544 ();
 sg13g2_fill_1 FILLER_32_550 ();
 sg13g2_fill_2 FILLER_32_577 ();
 sg13g2_decap_4 FILLER_32_615 ();
 sg13g2_decap_8 FILLER_32_660 ();
 sg13g2_fill_2 FILLER_32_667 ();
 sg13g2_fill_1 FILLER_32_805 ();
 sg13g2_fill_1 FILLER_32_873 ();
 sg13g2_fill_2 FILLER_32_892 ();
 sg13g2_fill_2 FILLER_32_905 ();
 sg13g2_fill_1 FILLER_32_907 ();
 sg13g2_fill_2 FILLER_32_944 ();
 sg13g2_fill_1 FILLER_32_946 ();
 sg13g2_fill_2 FILLER_32_977 ();
 sg13g2_fill_2 FILLER_32_988 ();
 sg13g2_fill_1 FILLER_32_990 ();
 sg13g2_fill_1 FILLER_32_1013 ();
 sg13g2_fill_1 FILLER_32_1049 ();
 sg13g2_fill_2 FILLER_32_1098 ();
 sg13g2_fill_1 FILLER_32_1100 ();
 sg13g2_fill_2 FILLER_32_1111 ();
 sg13g2_fill_2 FILLER_32_1177 ();
 sg13g2_fill_1 FILLER_32_1179 ();
 sg13g2_fill_1 FILLER_32_1268 ();
 sg13g2_fill_2 FILLER_32_1384 ();
 sg13g2_fill_2 FILLER_32_1506 ();
 sg13g2_fill_2 FILLER_32_1548 ();
 sg13g2_fill_1 FILLER_32_1580 ();
 sg13g2_decap_4 FILLER_32_1603 ();
 sg13g2_fill_1 FILLER_32_1607 ();
 sg13g2_fill_1 FILLER_32_1665 ();
 sg13g2_fill_2 FILLER_32_1701 ();
 sg13g2_fill_2 FILLER_32_1707 ();
 sg13g2_fill_1 FILLER_32_1709 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_33 ();
 sg13g2_fill_1 FILLER_33_35 ();
 sg13g2_fill_1 FILLER_33_60 ();
 sg13g2_fill_1 FILLER_33_85 ();
 sg13g2_fill_2 FILLER_33_110 ();
 sg13g2_fill_1 FILLER_33_170 ();
 sg13g2_fill_1 FILLER_33_196 ();
 sg13g2_decap_4 FILLER_33_233 ();
 sg13g2_fill_2 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_268 ();
 sg13g2_decap_4 FILLER_33_295 ();
 sg13g2_fill_2 FILLER_33_308 ();
 sg13g2_fill_2 FILLER_33_327 ();
 sg13g2_fill_1 FILLER_33_445 ();
 sg13g2_fill_1 FILLER_33_455 ();
 sg13g2_fill_2 FILLER_33_480 ();
 sg13g2_fill_1 FILLER_33_482 ();
 sg13g2_fill_2 FILLER_33_523 ();
 sg13g2_fill_2 FILLER_33_556 ();
 sg13g2_decap_4 FILLER_33_598 ();
 sg13g2_fill_1 FILLER_33_602 ();
 sg13g2_fill_1 FILLER_33_612 ();
 sg13g2_fill_2 FILLER_33_621 ();
 sg13g2_fill_1 FILLER_33_623 ();
 sg13g2_fill_1 FILLER_33_643 ();
 sg13g2_decap_8 FILLER_33_661 ();
 sg13g2_fill_2 FILLER_33_673 ();
 sg13g2_decap_4 FILLER_33_724 ();
 sg13g2_fill_1 FILLER_33_728 ();
 sg13g2_fill_2 FILLER_33_753 ();
 sg13g2_fill_1 FILLER_33_755 ();
 sg13g2_fill_1 FILLER_33_774 ();
 sg13g2_fill_2 FILLER_33_811 ();
 sg13g2_fill_1 FILLER_33_852 ();
 sg13g2_fill_1 FILLER_33_873 ();
 sg13g2_decap_4 FILLER_33_900 ();
 sg13g2_fill_1 FILLER_33_904 ();
 sg13g2_fill_1 FILLER_33_923 ();
 sg13g2_fill_2 FILLER_33_963 ();
 sg13g2_fill_1 FILLER_33_995 ();
 sg13g2_fill_2 FILLER_33_1010 ();
 sg13g2_fill_1 FILLER_33_1012 ();
 sg13g2_fill_2 FILLER_33_1032 ();
 sg13g2_fill_1 FILLER_33_1070 ();
 sg13g2_fill_2 FILLER_33_1097 ();
 sg13g2_fill_1 FILLER_33_1149 ();
 sg13g2_fill_2 FILLER_33_1206 ();
 sg13g2_fill_1 FILLER_33_1244 ();
 sg13g2_fill_2 FILLER_33_1274 ();
 sg13g2_fill_2 FILLER_33_1304 ();
 sg13g2_fill_1 FILLER_33_1306 ();
 sg13g2_decap_8 FILLER_33_1338 ();
 sg13g2_fill_1 FILLER_33_1345 ();
 sg13g2_decap_8 FILLER_33_1350 ();
 sg13g2_fill_1 FILLER_33_1385 ();
 sg13g2_decap_8 FILLER_33_1426 ();
 sg13g2_fill_2 FILLER_33_1433 ();
 sg13g2_fill_1 FILLER_33_1435 ();
 sg13g2_decap_8 FILLER_33_1454 ();
 sg13g2_fill_2 FILLER_33_1461 ();
 sg13g2_decap_4 FILLER_33_1487 ();
 sg13g2_fill_2 FILLER_33_1491 ();
 sg13g2_fill_1 FILLER_33_1537 ();
 sg13g2_fill_2 FILLER_33_1550 ();
 sg13g2_decap_8 FILLER_33_1597 ();
 sg13g2_fill_2 FILLER_33_1614 ();
 sg13g2_fill_1 FILLER_33_1635 ();
 sg13g2_fill_1 FILLER_33_1672 ();
 sg13g2_fill_1 FILLER_33_1767 ();
 sg13g2_fill_2 FILLER_34_84 ();
 sg13g2_fill_1 FILLER_34_86 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_fill_1 FILLER_34_150 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_fill_1 FILLER_34_283 ();
 sg13g2_fill_2 FILLER_34_392 ();
 sg13g2_fill_2 FILLER_34_478 ();
 sg13g2_fill_1 FILLER_34_480 ();
 sg13g2_fill_2 FILLER_34_491 ();
 sg13g2_fill_1 FILLER_34_493 ();
 sg13g2_fill_1 FILLER_34_571 ();
 sg13g2_fill_1 FILLER_34_581 ();
 sg13g2_fill_2 FILLER_34_595 ();
 sg13g2_fill_2 FILLER_34_623 ();
 sg13g2_fill_1 FILLER_34_625 ();
 sg13g2_fill_2 FILLER_34_657 ();
 sg13g2_fill_2 FILLER_34_701 ();
 sg13g2_decap_8 FILLER_34_725 ();
 sg13g2_fill_2 FILLER_34_732 ();
 sg13g2_fill_1 FILLER_34_734 ();
 sg13g2_fill_2 FILLER_34_776 ();
 sg13g2_fill_2 FILLER_34_788 ();
 sg13g2_fill_1 FILLER_34_790 ();
 sg13g2_fill_2 FILLER_34_823 ();
 sg13g2_fill_2 FILLER_34_959 ();
 sg13g2_fill_1 FILLER_34_961 ();
 sg13g2_fill_1 FILLER_34_1026 ();
 sg13g2_fill_2 FILLER_34_1103 ();
 sg13g2_decap_8 FILLER_34_1178 ();
 sg13g2_fill_1 FILLER_34_1185 ();
 sg13g2_fill_2 FILLER_34_1226 ();
 sg13g2_fill_2 FILLER_34_1245 ();
 sg13g2_fill_1 FILLER_34_1252 ();
 sg13g2_fill_2 FILLER_34_1297 ();
 sg13g2_decap_8 FILLER_34_1343 ();
 sg13g2_fill_1 FILLER_34_1397 ();
 sg13g2_fill_2 FILLER_34_1417 ();
 sg13g2_fill_1 FILLER_34_1419 ();
 sg13g2_fill_1 FILLER_34_1461 ();
 sg13g2_decap_4 FILLER_34_1484 ();
 sg13g2_fill_2 FILLER_34_1488 ();
 sg13g2_fill_1 FILLER_34_1498 ();
 sg13g2_fill_1 FILLER_34_1533 ();
 sg13g2_fill_1 FILLER_34_1562 ();
 sg13g2_fill_2 FILLER_34_1638 ();
 sg13g2_fill_1 FILLER_34_1640 ();
 sg13g2_fill_2 FILLER_34_1663 ();
 sg13g2_fill_1 FILLER_34_1665 ();
 sg13g2_fill_2 FILLER_34_1702 ();
 sg13g2_fill_2 FILLER_34_1719 ();
 sg13g2_fill_1 FILLER_34_1721 ();
 sg13g2_fill_1 FILLER_34_1732 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_1 FILLER_35_37 ();
 sg13g2_fill_2 FILLER_35_64 ();
 sg13g2_fill_1 FILLER_35_66 ();
 sg13g2_fill_2 FILLER_35_93 ();
 sg13g2_fill_1 FILLER_35_95 ();
 sg13g2_fill_1 FILLER_35_111 ();
 sg13g2_fill_2 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_195 ();
 sg13g2_decap_4 FILLER_35_215 ();
 sg13g2_fill_1 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_262 ();
 sg13g2_decap_8 FILLER_35_290 ();
 sg13g2_fill_2 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_451 ();
 sg13g2_fill_2 FILLER_35_457 ();
 sg13g2_fill_1 FILLER_35_459 ();
 sg13g2_fill_2 FILLER_35_490 ();
 sg13g2_fill_1 FILLER_35_492 ();
 sg13g2_fill_1 FILLER_35_512 ();
 sg13g2_decap_4 FILLER_35_545 ();
 sg13g2_fill_1 FILLER_35_549 ();
 sg13g2_decap_8 FILLER_35_591 ();
 sg13g2_fill_2 FILLER_35_598 ();
 sg13g2_fill_2 FILLER_35_604 ();
 sg13g2_fill_1 FILLER_35_606 ();
 sg13g2_fill_1 FILLER_35_639 ();
 sg13g2_decap_8 FILLER_35_649 ();
 sg13g2_fill_2 FILLER_35_666 ();
 sg13g2_fill_1 FILLER_35_731 ();
 sg13g2_fill_1 FILLER_35_782 ();
 sg13g2_fill_1 FILLER_35_809 ();
 sg13g2_fill_2 FILLER_35_868 ();
 sg13g2_fill_1 FILLER_35_880 ();
 sg13g2_fill_2 FILLER_35_909 ();
 sg13g2_fill_1 FILLER_35_921 ();
 sg13g2_fill_2 FILLER_35_965 ();
 sg13g2_fill_2 FILLER_35_977 ();
 sg13g2_fill_1 FILLER_35_979 ();
 sg13g2_fill_2 FILLER_35_999 ();
 sg13g2_fill_1 FILLER_35_1001 ();
 sg13g2_fill_2 FILLER_35_1033 ();
 sg13g2_fill_1 FILLER_35_1035 ();
 sg13g2_fill_1 FILLER_35_1088 ();
 sg13g2_decap_4 FILLER_35_1156 ();
 sg13g2_fill_2 FILLER_35_1160 ();
 sg13g2_decap_4 FILLER_35_1175 ();
 sg13g2_fill_1 FILLER_35_1179 ();
 sg13g2_fill_2 FILLER_35_1233 ();
 sg13g2_fill_2 FILLER_35_1285 ();
 sg13g2_fill_1 FILLER_35_1287 ();
 sg13g2_fill_1 FILLER_35_1324 ();
 sg13g2_decap_4 FILLER_35_1359 ();
 sg13g2_fill_1 FILLER_35_1363 ();
 sg13g2_decap_4 FILLER_35_1385 ();
 sg13g2_fill_1 FILLER_35_1397 ();
 sg13g2_decap_4 FILLER_35_1424 ();
 sg13g2_fill_1 FILLER_35_1467 ();
 sg13g2_decap_4 FILLER_35_1494 ();
 sg13g2_fill_1 FILLER_35_1529 ();
 sg13g2_fill_2 FILLER_35_1540 ();
 sg13g2_fill_2 FILLER_35_1590 ();
 sg13g2_fill_1 FILLER_35_1610 ();
 sg13g2_fill_1 FILLER_35_1621 ();
 sg13g2_fill_1 FILLER_35_1627 ();
 sg13g2_fill_1 FILLER_35_1661 ();
 sg13g2_fill_2 FILLER_35_1699 ();
 sg13g2_fill_1 FILLER_35_1727 ();
 sg13g2_fill_1 FILLER_35_1767 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_30 ();
 sg13g2_fill_1 FILLER_36_32 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_fill_2 FILLER_36_139 ();
 sg13g2_fill_1 FILLER_36_151 ();
 sg13g2_fill_2 FILLER_36_190 ();
 sg13g2_fill_1 FILLER_36_192 ();
 sg13g2_decap_4 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_36_214 ();
 sg13g2_decap_4 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_277 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_354 ();
 sg13g2_fill_1 FILLER_36_364 ();
 sg13g2_fill_2 FILLER_36_373 ();
 sg13g2_fill_2 FILLER_36_411 ();
 sg13g2_fill_2 FILLER_36_489 ();
 sg13g2_fill_2 FILLER_36_501 ();
 sg13g2_fill_1 FILLER_36_546 ();
 sg13g2_fill_1 FILLER_36_583 ();
 sg13g2_fill_2 FILLER_36_615 ();
 sg13g2_fill_2 FILLER_36_631 ();
 sg13g2_fill_1 FILLER_36_633 ();
 sg13g2_fill_1 FILLER_36_647 ();
 sg13g2_decap_8 FILLER_36_665 ();
 sg13g2_fill_1 FILLER_36_672 ();
 sg13g2_decap_4 FILLER_36_719 ();
 sg13g2_fill_2 FILLER_36_723 ();
 sg13g2_fill_1 FILLER_36_792 ();
 sg13g2_fill_2 FILLER_36_854 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_fill_1 FILLER_36_949 ();
 sg13g2_fill_1 FILLER_36_986 ();
 sg13g2_decap_8 FILLER_36_1026 ();
 sg13g2_fill_2 FILLER_36_1059 ();
 sg13g2_decap_8 FILLER_36_1091 ();
 sg13g2_fill_2 FILLER_36_1098 ();
 sg13g2_fill_2 FILLER_36_1104 ();
 sg13g2_fill_1 FILLER_36_1106 ();
 sg13g2_fill_1 FILLER_36_1129 ();
 sg13g2_fill_2 FILLER_36_1144 ();
 sg13g2_fill_2 FILLER_36_1252 ();
 sg13g2_fill_1 FILLER_36_1307 ();
 sg13g2_fill_2 FILLER_36_1321 ();
 sg13g2_fill_1 FILLER_36_1323 ();
 sg13g2_fill_2 FILLER_36_1334 ();
 sg13g2_fill_2 FILLER_36_1359 ();
 sg13g2_fill_1 FILLER_36_1361 ();
 sg13g2_fill_2 FILLER_36_1372 ();
 sg13g2_fill_1 FILLER_36_1374 ();
 sg13g2_fill_1 FILLER_36_1401 ();
 sg13g2_fill_1 FILLER_36_1467 ();
 sg13g2_fill_1 FILLER_36_1481 ();
 sg13g2_fill_2 FILLER_36_1492 ();
 sg13g2_fill_1 FILLER_36_1494 ();
 sg13g2_fill_2 FILLER_36_1511 ();
 sg13g2_fill_2 FILLER_36_1518 ();
 sg13g2_fill_1 FILLER_36_1550 ();
 sg13g2_fill_1 FILLER_36_1641 ();
 sg13g2_fill_1 FILLER_36_1678 ();
 sg13g2_fill_2 FILLER_36_1766 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_decap_4 FILLER_37_31 ();
 sg13g2_fill_2 FILLER_37_35 ();
 sg13g2_decap_4 FILLER_37_80 ();
 sg13g2_fill_1 FILLER_37_84 ();
 sg13g2_fill_1 FILLER_37_112 ();
 sg13g2_fill_1 FILLER_37_174 ();
 sg13g2_decap_8 FILLER_37_219 ();
 sg13g2_fill_2 FILLER_37_230 ();
 sg13g2_fill_1 FILLER_37_232 ();
 sg13g2_fill_2 FILLER_37_259 ();
 sg13g2_fill_1 FILLER_37_261 ();
 sg13g2_fill_2 FILLER_37_284 ();
 sg13g2_fill_1 FILLER_37_286 ();
 sg13g2_fill_1 FILLER_37_297 ();
 sg13g2_fill_2 FILLER_37_348 ();
 sg13g2_fill_1 FILLER_37_350 ();
 sg13g2_decap_4 FILLER_37_361 ();
 sg13g2_fill_2 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_419 ();
 sg13g2_fill_1 FILLER_37_421 ();
 sg13g2_fill_1 FILLER_37_467 ();
 sg13g2_fill_1 FILLER_37_512 ();
 sg13g2_fill_1 FILLER_37_576 ();
 sg13g2_fill_2 FILLER_37_594 ();
 sg13g2_fill_2 FILLER_37_700 ();
 sg13g2_fill_1 FILLER_37_702 ();
 sg13g2_fill_2 FILLER_37_721 ();
 sg13g2_fill_1 FILLER_37_723 ();
 sg13g2_decap_8 FILLER_37_732 ();
 sg13g2_fill_1 FILLER_37_739 ();
 sg13g2_decap_4 FILLER_37_748 ();
 sg13g2_fill_2 FILLER_37_761 ();
 sg13g2_fill_1 FILLER_37_772 ();
 sg13g2_decap_4 FILLER_37_777 ();
 sg13g2_fill_2 FILLER_37_781 ();
 sg13g2_fill_2 FILLER_37_813 ();
 sg13g2_fill_2 FILLER_37_897 ();
 sg13g2_fill_2 FILLER_37_995 ();
 sg13g2_fill_1 FILLER_37_997 ();
 sg13g2_fill_1 FILLER_37_1011 ();
 sg13g2_decap_4 FILLER_37_1026 ();
 sg13g2_fill_1 FILLER_37_1030 ();
 sg13g2_fill_1 FILLER_37_1054 ();
 sg13g2_fill_1 FILLER_37_1078 ();
 sg13g2_fill_2 FILLER_37_1089 ();
 sg13g2_fill_2 FILLER_37_1095 ();
 sg13g2_fill_2 FILLER_37_1107 ();
 sg13g2_decap_4 FILLER_37_1153 ();
 sg13g2_fill_1 FILLER_37_1157 ();
 sg13g2_fill_2 FILLER_37_1185 ();
 sg13g2_fill_1 FILLER_37_1187 ();
 sg13g2_fill_2 FILLER_37_1291 ();
 sg13g2_fill_1 FILLER_37_1293 ();
 sg13g2_fill_2 FILLER_37_1308 ();
 sg13g2_fill_2 FILLER_37_1345 ();
 sg13g2_fill_1 FILLER_37_1347 ();
 sg13g2_decap_4 FILLER_37_1434 ();
 sg13g2_fill_2 FILLER_37_1438 ();
 sg13g2_fill_1 FILLER_37_1466 ();
 sg13g2_fill_1 FILLER_37_1472 ();
 sg13g2_fill_1 FILLER_37_1494 ();
 sg13g2_fill_1 FILLER_37_1610 ();
 sg13g2_fill_2 FILLER_37_1657 ();
 sg13g2_fill_1 FILLER_37_1659 ();
 sg13g2_decap_4 FILLER_37_1685 ();
 sg13g2_fill_1 FILLER_37_1689 ();
 sg13g2_fill_2 FILLER_37_1709 ();
 sg13g2_fill_1 FILLER_37_1711 ();
 sg13g2_fill_2 FILLER_37_1726 ();
 sg13g2_fill_1 FILLER_37_1728 ();
 sg13g2_fill_2 FILLER_37_1739 ();
 sg13g2_fill_1 FILLER_37_1767 ();
 sg13g2_fill_2 FILLER_38_36 ();
 sg13g2_fill_2 FILLER_38_85 ();
 sg13g2_fill_1 FILLER_38_97 ();
 sg13g2_decap_4 FILLER_38_102 ();
 sg13g2_fill_1 FILLER_38_111 ();
 sg13g2_fill_2 FILLER_38_121 ();
 sg13g2_fill_2 FILLER_38_138 ();
 sg13g2_fill_2 FILLER_38_150 ();
 sg13g2_fill_1 FILLER_38_152 ();
 sg13g2_decap_4 FILLER_38_175 ();
 sg13g2_fill_1 FILLER_38_179 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_fill_1 FILLER_38_296 ();
 sg13g2_fill_1 FILLER_38_323 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_412 ();
 sg13g2_decap_4 FILLER_38_419 ();
 sg13g2_fill_2 FILLER_38_427 ();
 sg13g2_fill_2 FILLER_38_571 ();
 sg13g2_fill_2 FILLER_38_614 ();
 sg13g2_fill_1 FILLER_38_616 ();
 sg13g2_fill_2 FILLER_38_668 ();
 sg13g2_fill_1 FILLER_38_670 ();
 sg13g2_fill_1 FILLER_38_684 ();
 sg13g2_fill_1 FILLER_38_695 ();
 sg13g2_fill_2 FILLER_38_717 ();
 sg13g2_fill_1 FILLER_38_771 ();
 sg13g2_fill_1 FILLER_38_777 ();
 sg13g2_fill_2 FILLER_38_832 ();
 sg13g2_fill_1 FILLER_38_862 ();
 sg13g2_fill_1 FILLER_38_881 ();
 sg13g2_fill_2 FILLER_38_891 ();
 sg13g2_fill_1 FILLER_38_926 ();
 sg13g2_fill_2 FILLER_38_937 ();
 sg13g2_fill_2 FILLER_38_975 ();
 sg13g2_fill_1 FILLER_38_977 ();
 sg13g2_fill_2 FILLER_38_1014 ();
 sg13g2_fill_2 FILLER_38_1047 ();
 sg13g2_fill_1 FILLER_38_1049 ();
 sg13g2_fill_2 FILLER_38_1205 ();
 sg13g2_fill_1 FILLER_38_1207 ();
 sg13g2_fill_1 FILLER_38_1234 ();
 sg13g2_fill_1 FILLER_38_1250 ();
 sg13g2_fill_2 FILLER_38_1285 ();
 sg13g2_fill_1 FILLER_38_1287 ();
 sg13g2_decap_8 FILLER_38_1314 ();
 sg13g2_fill_2 FILLER_38_1325 ();
 sg13g2_decap_4 FILLER_38_1348 ();
 sg13g2_fill_1 FILLER_38_1352 ();
 sg13g2_fill_2 FILLER_38_1361 ();
 sg13g2_fill_2 FILLER_38_1396 ();
 sg13g2_fill_1 FILLER_38_1398 ();
 sg13g2_fill_2 FILLER_38_1414 ();
 sg13g2_fill_1 FILLER_38_1416 ();
 sg13g2_fill_1 FILLER_38_1443 ();
 sg13g2_fill_2 FILLER_38_1448 ();
 sg13g2_fill_1 FILLER_38_1450 ();
 sg13g2_decap_8 FILLER_38_1491 ();
 sg13g2_decap_4 FILLER_38_1498 ();
 sg13g2_decap_4 FILLER_38_1507 ();
 sg13g2_decap_8 FILLER_38_1515 ();
 sg13g2_fill_2 FILLER_38_1522 ();
 sg13g2_fill_1 FILLER_38_1534 ();
 sg13g2_fill_1 FILLER_38_1545 ();
 sg13g2_fill_2 FILLER_38_1560 ();
 sg13g2_fill_2 FILLER_38_1570 ();
 sg13g2_fill_2 FILLER_38_1585 ();
 sg13g2_fill_2 FILLER_38_1645 ();
 sg13g2_fill_1 FILLER_38_1647 ();
 sg13g2_fill_1 FILLER_38_1688 ();
 sg13g2_fill_2 FILLER_38_1707 ();
 sg13g2_fill_2 FILLER_38_1766 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_34 ();
 sg13g2_fill_2 FILLER_39_73 ();
 sg13g2_fill_1 FILLER_39_114 ();
 sg13g2_fill_2 FILLER_39_141 ();
 sg13g2_decap_8 FILLER_39_169 ();
 sg13g2_decap_8 FILLER_39_180 ();
 sg13g2_decap_4 FILLER_39_187 ();
 sg13g2_fill_2 FILLER_39_217 ();
 sg13g2_fill_1 FILLER_39_219 ();
 sg13g2_decap_4 FILLER_39_294 ();
 sg13g2_fill_2 FILLER_39_298 ();
 sg13g2_fill_1 FILLER_39_309 ();
 sg13g2_fill_2 FILLER_39_344 ();
 sg13g2_fill_1 FILLER_39_346 ();
 sg13g2_fill_1 FILLER_39_360 ();
 sg13g2_fill_2 FILLER_39_397 ();
 sg13g2_fill_1 FILLER_39_399 ();
 sg13g2_fill_2 FILLER_39_550 ();
 sg13g2_fill_1 FILLER_39_552 ();
 sg13g2_fill_2 FILLER_39_573 ();
 sg13g2_fill_2 FILLER_39_581 ();
 sg13g2_fill_2 FILLER_39_596 ();
 sg13g2_fill_2 FILLER_39_656 ();
 sg13g2_fill_1 FILLER_39_658 ();
 sg13g2_fill_2 FILLER_39_682 ();
 sg13g2_fill_2 FILLER_39_714 ();
 sg13g2_fill_2 FILLER_39_790 ();
 sg13g2_decap_8 FILLER_39_850 ();
 sg13g2_fill_1 FILLER_39_934 ();
 sg13g2_fill_1 FILLER_39_966 ();
 sg13g2_fill_1 FILLER_39_976 ();
 sg13g2_fill_2 FILLER_39_994 ();
 sg13g2_fill_1 FILLER_39_996 ();
 sg13g2_fill_2 FILLER_39_1011 ();
 sg13g2_decap_8 FILLER_39_1031 ();
 sg13g2_fill_1 FILLER_39_1038 ();
 sg13g2_fill_1 FILLER_39_1054 ();
 sg13g2_fill_1 FILLER_39_1069 ();
 sg13g2_fill_1 FILLER_39_1144 ();
 sg13g2_fill_1 FILLER_39_1225 ();
 sg13g2_fill_1 FILLER_39_1240 ();
 sg13g2_fill_1 FILLER_39_1257 ();
 sg13g2_fill_2 FILLER_39_1269 ();
 sg13g2_decap_4 FILLER_39_1275 ();
 sg13g2_fill_1 FILLER_39_1335 ();
 sg13g2_fill_2 FILLER_39_1378 ();
 sg13g2_fill_1 FILLER_39_1380 ();
 sg13g2_fill_1 FILLER_39_1427 ();
 sg13g2_fill_2 FILLER_39_1468 ();
 sg13g2_fill_1 FILLER_39_1470 ();
 sg13g2_fill_1 FILLER_39_1480 ();
 sg13g2_fill_1 FILLER_39_1516 ();
 sg13g2_fill_2 FILLER_39_1521 ();
 sg13g2_fill_1 FILLER_39_1523 ();
 sg13g2_fill_2 FILLER_39_1534 ();
 sg13g2_fill_1 FILLER_39_1536 ();
 sg13g2_fill_1 FILLER_39_1603 ();
 sg13g2_fill_2 FILLER_39_1634 ();
 sg13g2_fill_1 FILLER_39_1636 ();
 sg13g2_fill_1 FILLER_39_1671 ();
 sg13g2_fill_2 FILLER_39_1744 ();
 sg13g2_fill_2 FILLER_40_26 ();
 sg13g2_decap_4 FILLER_40_68 ();
 sg13g2_fill_2 FILLER_40_151 ();
 sg13g2_fill_1 FILLER_40_153 ();
 sg13g2_fill_2 FILLER_40_162 ();
 sg13g2_fill_1 FILLER_40_164 ();
 sg13g2_decap_8 FILLER_40_211 ();
 sg13g2_fill_2 FILLER_40_218 ();
 sg13g2_fill_1 FILLER_40_220 ();
 sg13g2_decap_4 FILLER_40_256 ();
 sg13g2_fill_1 FILLER_40_260 ();
 sg13g2_fill_2 FILLER_40_285 ();
 sg13g2_fill_1 FILLER_40_292 ();
 sg13g2_fill_2 FILLER_40_316 ();
 sg13g2_decap_4 FILLER_40_323 ();
 sg13g2_fill_2 FILLER_40_382 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_2 FILLER_40_421 ();
 sg13g2_fill_1 FILLER_40_423 ();
 sg13g2_fill_2 FILLER_40_437 ();
 sg13g2_fill_1 FILLER_40_439 ();
 sg13g2_fill_2 FILLER_40_463 ();
 sg13g2_fill_1 FILLER_40_465 ();
 sg13g2_decap_4 FILLER_40_484 ();
 sg13g2_decap_4 FILLER_40_515 ();
 sg13g2_fill_2 FILLER_40_546 ();
 sg13g2_fill_1 FILLER_40_548 ();
 sg13g2_fill_2 FILLER_40_561 ();
 sg13g2_fill_2 FILLER_40_587 ();
 sg13g2_fill_2 FILLER_40_617 ();
 sg13g2_fill_1 FILLER_40_619 ();
 sg13g2_decap_4 FILLER_40_639 ();
 sg13g2_fill_2 FILLER_40_643 ();
 sg13g2_decap_4 FILLER_40_671 ();
 sg13g2_fill_2 FILLER_40_722 ();
 sg13g2_fill_1 FILLER_40_724 ();
 sg13g2_fill_2 FILLER_40_754 ();
 sg13g2_fill_1 FILLER_40_756 ();
 sg13g2_fill_1 FILLER_40_786 ();
 sg13g2_fill_1 FILLER_40_813 ();
 sg13g2_fill_2 FILLER_40_843 ();
 sg13g2_fill_1 FILLER_40_894 ();
 sg13g2_fill_2 FILLER_40_926 ();
 sg13g2_fill_2 FILLER_40_957 ();
 sg13g2_fill_2 FILLER_40_995 ();
 sg13g2_fill_1 FILLER_40_997 ();
 sg13g2_fill_1 FILLER_40_1024 ();
 sg13g2_decap_8 FILLER_40_1030 ();
 sg13g2_fill_2 FILLER_40_1037 ();
 sg13g2_fill_1 FILLER_40_1039 ();
 sg13g2_fill_1 FILLER_40_1076 ();
 sg13g2_fill_2 FILLER_40_1147 ();
 sg13g2_fill_2 FILLER_40_1167 ();
 sg13g2_fill_1 FILLER_40_1169 ();
 sg13g2_fill_2 FILLER_40_1180 ();
 sg13g2_fill_1 FILLER_40_1182 ();
 sg13g2_fill_1 FILLER_40_1214 ();
 sg13g2_decap_4 FILLER_40_1241 ();
 sg13g2_fill_1 FILLER_40_1245 ();
 sg13g2_fill_2 FILLER_40_1269 ();
 sg13g2_fill_2 FILLER_40_1281 ();
 sg13g2_fill_1 FILLER_40_1283 ();
 sg13g2_decap_4 FILLER_40_1316 ();
 sg13g2_fill_1 FILLER_40_1343 ();
 sg13g2_fill_2 FILLER_40_1390 ();
 sg13g2_fill_1 FILLER_40_1396 ();
 sg13g2_decap_8 FILLER_40_1406 ();
 sg13g2_fill_2 FILLER_40_1426 ();
 sg13g2_fill_1 FILLER_40_1428 ();
 sg13g2_decap_8 FILLER_40_1551 ();
 sg13g2_decap_8 FILLER_40_1558 ();
 sg13g2_decap_4 FILLER_40_1565 ();
 sg13g2_fill_2 FILLER_40_1569 ();
 sg13g2_fill_2 FILLER_40_1575 ();
 sg13g2_fill_2 FILLER_40_1591 ();
 sg13g2_fill_2 FILLER_40_1619 ();
 sg13g2_fill_1 FILLER_40_1650 ();
 sg13g2_fill_2 FILLER_40_1660 ();
 sg13g2_decap_8 FILLER_40_1702 ();
 sg13g2_decap_8 FILLER_40_1709 ();
 sg13g2_fill_1 FILLER_40_1716 ();
 sg13g2_fill_2 FILLER_40_1738 ();
 sg13g2_fill_1 FILLER_40_1740 ();
 sg13g2_fill_1 FILLER_40_1767 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_fill_1 FILLER_41_9 ();
 sg13g2_fill_2 FILLER_41_84 ();
 sg13g2_fill_1 FILLER_41_86 ();
 sg13g2_decap_4 FILLER_41_101 ();
 sg13g2_fill_1 FILLER_41_115 ();
 sg13g2_fill_2 FILLER_41_142 ();
 sg13g2_fill_1 FILLER_41_144 ();
 sg13g2_decap_4 FILLER_41_155 ();
 sg13g2_fill_1 FILLER_41_163 ();
 sg13g2_decap_4 FILLER_41_174 ();
 sg13g2_fill_2 FILLER_41_178 ();
 sg13g2_fill_2 FILLER_41_236 ();
 sg13g2_decap_8 FILLER_41_269 ();
 sg13g2_fill_1 FILLER_41_310 ();
 sg13g2_fill_2 FILLER_41_321 ();
 sg13g2_fill_2 FILLER_41_367 ();
 sg13g2_fill_1 FILLER_41_369 ();
 sg13g2_decap_8 FILLER_41_396 ();
 sg13g2_decap_4 FILLER_41_403 ();
 sg13g2_fill_1 FILLER_41_407 ();
 sg13g2_fill_1 FILLER_41_444 ();
 sg13g2_fill_2 FILLER_41_471 ();
 sg13g2_decap_8 FILLER_41_551 ();
 sg13g2_fill_1 FILLER_41_558 ();
 sg13g2_fill_1 FILLER_41_574 ();
 sg13g2_decap_4 FILLER_41_635 ();
 sg13g2_fill_2 FILLER_41_639 ();
 sg13g2_decap_8 FILLER_41_651 ();
 sg13g2_fill_2 FILLER_41_667 ();
 sg13g2_fill_1 FILLER_41_669 ();
 sg13g2_fill_2 FILLER_41_680 ();
 sg13g2_fill_1 FILLER_41_682 ();
 sg13g2_decap_4 FILLER_41_696 ();
 sg13g2_fill_2 FILLER_41_740 ();
 sg13g2_fill_1 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_806 ();
 sg13g2_decap_4 FILLER_41_875 ();
 sg13g2_fill_1 FILLER_41_879 ();
 sg13g2_fill_2 FILLER_41_942 ();
 sg13g2_fill_1 FILLER_41_944 ();
 sg13g2_decap_8 FILLER_41_993 ();
 sg13g2_decap_8 FILLER_41_1000 ();
 sg13g2_fill_1 FILLER_41_1007 ();
 sg13g2_decap_8 FILLER_41_1043 ();
 sg13g2_fill_1 FILLER_41_1050 ();
 sg13g2_fill_2 FILLER_41_1055 ();
 sg13g2_fill_2 FILLER_41_1078 ();
 sg13g2_fill_2 FILLER_41_1131 ();
 sg13g2_fill_2 FILLER_41_1152 ();
 sg13g2_decap_4 FILLER_41_1220 ();
 sg13g2_fill_2 FILLER_41_1224 ();
 sg13g2_decap_8 FILLER_41_1230 ();
 sg13g2_decap_4 FILLER_41_1237 ();
 sg13g2_fill_1 FILLER_41_1241 ();
 sg13g2_decap_4 FILLER_41_1287 ();
 sg13g2_fill_1 FILLER_41_1321 ();
 sg13g2_fill_2 FILLER_41_1374 ();
 sg13g2_decap_8 FILLER_41_1380 ();
 sg13g2_fill_2 FILLER_41_1387 ();
 sg13g2_fill_2 FILLER_41_1413 ();
 sg13g2_fill_1 FILLER_41_1437 ();
 sg13g2_fill_2 FILLER_41_1492 ();
 sg13g2_fill_2 FILLER_41_1504 ();
 sg13g2_fill_2 FILLER_41_1520 ();
 sg13g2_fill_1 FILLER_41_1522 ();
 sg13g2_decap_8 FILLER_41_1540 ();
 sg13g2_fill_2 FILLER_41_1547 ();
 sg13g2_fill_1 FILLER_41_1549 ();
 sg13g2_fill_2 FILLER_41_1634 ();
 sg13g2_fill_2 FILLER_41_1668 ();
 sg13g2_fill_1 FILLER_41_1679 ();
 sg13g2_fill_1 FILLER_41_1693 ();
 sg13g2_decap_8 FILLER_41_1699 ();
 sg13g2_fill_1 FILLER_41_1706 ();
 sg13g2_fill_2 FILLER_41_1733 ();
 sg13g2_fill_1 FILLER_41_1735 ();
 sg13g2_fill_2 FILLER_41_1766 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_4 FILLER_42_7 ();
 sg13g2_fill_2 FILLER_42_37 ();
 sg13g2_fill_1 FILLER_42_39 ();
 sg13g2_decap_4 FILLER_42_77 ();
 sg13g2_fill_2 FILLER_42_104 ();
 sg13g2_fill_2 FILLER_42_145 ();
 sg13g2_fill_1 FILLER_42_147 ();
 sg13g2_fill_2 FILLER_42_174 ();
 sg13g2_decap_4 FILLER_42_190 ();
 sg13g2_fill_1 FILLER_42_247 ();
 sg13g2_decap_8 FILLER_42_288 ();
 sg13g2_fill_2 FILLER_42_338 ();
 sg13g2_fill_1 FILLER_42_340 ();
 sg13g2_fill_2 FILLER_42_360 ();
 sg13g2_decap_4 FILLER_42_435 ();
 sg13g2_fill_1 FILLER_42_439 ();
 sg13g2_fill_2 FILLER_42_461 ();
 sg13g2_fill_2 FILLER_42_481 ();
 sg13g2_fill_2 FILLER_42_509 ();
 sg13g2_fill_1 FILLER_42_511 ();
 sg13g2_fill_1 FILLER_42_592 ();
 sg13g2_fill_2 FILLER_42_602 ();
 sg13g2_fill_2 FILLER_42_613 ();
 sg13g2_fill_1 FILLER_42_615 ();
 sg13g2_fill_2 FILLER_42_652 ();
 sg13g2_decap_4 FILLER_42_692 ();
 sg13g2_fill_2 FILLER_42_696 ();
 sg13g2_fill_2 FILLER_42_724 ();
 sg13g2_fill_1 FILLER_42_726 ();
 sg13g2_fill_1 FILLER_42_753 ();
 sg13g2_fill_2 FILLER_42_758 ();
 sg13g2_decap_4 FILLER_42_812 ();
 sg13g2_fill_1 FILLER_42_816 ();
 sg13g2_fill_1 FILLER_42_846 ();
 sg13g2_decap_4 FILLER_42_876 ();
 sg13g2_decap_4 FILLER_42_956 ();
 sg13g2_fill_1 FILLER_42_960 ();
 sg13g2_decap_4 FILLER_42_989 ();
 sg13g2_fill_1 FILLER_42_1019 ();
 sg13g2_fill_2 FILLER_42_1069 ();
 sg13g2_fill_2 FILLER_42_1112 ();
 sg13g2_fill_1 FILLER_42_1114 ();
 sg13g2_fill_2 FILLER_42_1170 ();
 sg13g2_fill_1 FILLER_42_1172 ();
 sg13g2_fill_1 FILLER_42_1203 ();
 sg13g2_fill_2 FILLER_42_1240 ();
 sg13g2_fill_1 FILLER_42_1242 ();
 sg13g2_fill_2 FILLER_42_1263 ();
 sg13g2_fill_1 FILLER_42_1265 ();
 sg13g2_fill_1 FILLER_42_1324 ();
 sg13g2_fill_1 FILLER_42_1339 ();
 sg13g2_fill_1 FILLER_42_1368 ();
 sg13g2_fill_1 FILLER_42_1413 ();
 sg13g2_decap_8 FILLER_42_1552 ();
 sg13g2_fill_1 FILLER_42_1559 ();
 sg13g2_fill_2 FILLER_42_1602 ();
 sg13g2_fill_1 FILLER_42_1604 ();
 sg13g2_fill_2 FILLER_42_1665 ();
 sg13g2_decap_4 FILLER_42_1702 ();
 sg13g2_fill_2 FILLER_42_1706 ();
 sg13g2_fill_2 FILLER_42_1728 ();
 sg13g2_fill_2 FILLER_42_1740 ();
 sg13g2_fill_2 FILLER_43_30 ();
 sg13g2_fill_1 FILLER_43_32 ();
 sg13g2_fill_1 FILLER_43_120 ();
 sg13g2_fill_1 FILLER_43_144 ();
 sg13g2_fill_1 FILLER_43_175 ();
 sg13g2_fill_2 FILLER_43_214 ();
 sg13g2_fill_1 FILLER_43_216 ();
 sg13g2_fill_1 FILLER_43_267 ();
 sg13g2_fill_1 FILLER_43_310 ();
 sg13g2_fill_2 FILLER_43_329 ();
 sg13g2_fill_2 FILLER_43_355 ();
 sg13g2_decap_4 FILLER_43_410 ();
 sg13g2_decap_4 FILLER_43_437 ();
 sg13g2_fill_1 FILLER_43_441 ();
 sg13g2_decap_4 FILLER_43_478 ();
 sg13g2_fill_2 FILLER_43_482 ();
 sg13g2_fill_2 FILLER_43_504 ();
 sg13g2_fill_1 FILLER_43_506 ();
 sg13g2_fill_2 FILLER_43_516 ();
 sg13g2_fill_1 FILLER_43_528 ();
 sg13g2_fill_1 FILLER_43_542 ();
 sg13g2_decap_8 FILLER_43_564 ();
 sg13g2_fill_2 FILLER_43_610 ();
 sg13g2_fill_1 FILLER_43_612 ();
 sg13g2_fill_1 FILLER_43_623 ();
 sg13g2_fill_1 FILLER_43_650 ();
 sg13g2_decap_8 FILLER_43_659 ();
 sg13g2_fill_2 FILLER_43_726 ();
 sg13g2_fill_1 FILLER_43_728 ();
 sg13g2_decap_4 FILLER_43_779 ();
 sg13g2_fill_1 FILLER_43_793 ();
 sg13g2_decap_4 FILLER_43_820 ();
 sg13g2_fill_1 FILLER_43_824 ();
 sg13g2_fill_2 FILLER_43_861 ();
 sg13g2_decap_4 FILLER_43_880 ();
 sg13g2_fill_2 FILLER_43_884 ();
 sg13g2_fill_2 FILLER_43_912 ();
 sg13g2_fill_2 FILLER_43_952 ();
 sg13g2_fill_1 FILLER_43_954 ();
 sg13g2_fill_2 FILLER_43_986 ();
 sg13g2_fill_2 FILLER_43_998 ();
 sg13g2_fill_1 FILLER_43_1000 ();
 sg13g2_fill_2 FILLER_43_1014 ();
 sg13g2_fill_2 FILLER_43_1035 ();
 sg13g2_fill_1 FILLER_43_1081 ();
 sg13g2_decap_4 FILLER_43_1086 ();
 sg13g2_fill_1 FILLER_43_1090 ();
 sg13g2_fill_1 FILLER_43_1101 ();
 sg13g2_decap_8 FILLER_43_1106 ();
 sg13g2_decap_8 FILLER_43_1123 ();
 sg13g2_decap_4 FILLER_43_1130 ();
 sg13g2_fill_1 FILLER_43_1134 ();
 sg13g2_fill_2 FILLER_43_1148 ();
 sg13g2_fill_2 FILLER_43_1164 ();
 sg13g2_fill_1 FILLER_43_1166 ();
 sg13g2_fill_2 FILLER_43_1176 ();
 sg13g2_fill_2 FILLER_43_1210 ();
 sg13g2_decap_4 FILLER_43_1229 ();
 sg13g2_fill_1 FILLER_43_1233 ();
 sg13g2_decap_4 FILLER_43_1242 ();
 sg13g2_fill_1 FILLER_43_1246 ();
 sg13g2_fill_2 FILLER_43_1306 ();
 sg13g2_fill_2 FILLER_43_1336 ();
 sg13g2_fill_2 FILLER_43_1342 ();
 sg13g2_fill_1 FILLER_43_1344 ();
 sg13g2_decap_8 FILLER_43_1396 ();
 sg13g2_decap_8 FILLER_43_1403 ();
 sg13g2_fill_1 FILLER_43_1410 ();
 sg13g2_fill_1 FILLER_43_1421 ();
 sg13g2_fill_2 FILLER_43_1437 ();
 sg13g2_fill_1 FILLER_43_1439 ();
 sg13g2_fill_2 FILLER_43_1454 ();
 sg13g2_fill_2 FILLER_43_1470 ();
 sg13g2_fill_1 FILLER_43_1472 ();
 sg13g2_fill_2 FILLER_43_1497 ();
 sg13g2_fill_1 FILLER_43_1509 ();
 sg13g2_decap_4 FILLER_43_1524 ();
 sg13g2_decap_4 FILLER_43_1532 ();
 sg13g2_fill_1 FILLER_43_1536 ();
 sg13g2_fill_1 FILLER_43_1593 ();
 sg13g2_fill_2 FILLER_43_1656 ();
 sg13g2_fill_1 FILLER_43_1658 ();
 sg13g2_fill_1 FILLER_43_1688 ();
 sg13g2_fill_2 FILLER_43_1715 ();
 sg13g2_fill_2 FILLER_43_1765 ();
 sg13g2_fill_1 FILLER_43_1767 ();
 sg13g2_fill_1 FILLER_44_46 ();
 sg13g2_fill_1 FILLER_44_61 ();
 sg13g2_decap_8 FILLER_44_89 ();
 sg13g2_fill_2 FILLER_44_96 ();
 sg13g2_fill_2 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_fill_2 FILLER_44_189 ();
 sg13g2_fill_1 FILLER_44_191 ();
 sg13g2_decap_4 FILLER_44_241 ();
 sg13g2_fill_1 FILLER_44_254 ();
 sg13g2_fill_2 FILLER_44_323 ();
 sg13g2_fill_1 FILLER_44_360 ();
 sg13g2_decap_4 FILLER_44_552 ();
 sg13g2_fill_1 FILLER_44_560 ();
 sg13g2_fill_2 FILLER_44_596 ();
 sg13g2_fill_1 FILLER_44_616 ();
 sg13g2_fill_2 FILLER_44_653 ();
 sg13g2_decap_8 FILLER_44_747 ();
 sg13g2_fill_2 FILLER_44_758 ();
 sg13g2_fill_1 FILLER_44_790 ();
 sg13g2_fill_1 FILLER_44_813 ();
 sg13g2_fill_2 FILLER_44_824 ();
 sg13g2_fill_1 FILLER_44_826 ();
 sg13g2_fill_1 FILLER_44_854 ();
 sg13g2_decap_4 FILLER_44_891 ();
 sg13g2_fill_2 FILLER_44_895 ();
 sg13g2_decap_8 FILLER_44_901 ();
 sg13g2_decap_4 FILLER_44_908 ();
 sg13g2_fill_2 FILLER_44_912 ();
 sg13g2_fill_2 FILLER_44_922 ();
 sg13g2_fill_1 FILLER_44_924 ();
 sg13g2_fill_1 FILLER_44_943 ();
 sg13g2_fill_1 FILLER_44_969 ();
 sg13g2_fill_2 FILLER_44_1054 ();
 sg13g2_fill_1 FILLER_44_1056 ();
 sg13g2_fill_1 FILLER_44_1083 ();
 sg13g2_fill_2 FILLER_44_1118 ();
 sg13g2_fill_1 FILLER_44_1120 ();
 sg13g2_fill_2 FILLER_44_1151 ();
 sg13g2_fill_1 FILLER_44_1153 ();
 sg13g2_fill_1 FILLER_44_1216 ();
 sg13g2_fill_2 FILLER_44_1279 ();
 sg13g2_fill_1 FILLER_44_1326 ();
 sg13g2_fill_2 FILLER_44_1363 ();
 sg13g2_fill_1 FILLER_44_1365 ();
 sg13g2_fill_1 FILLER_44_1379 ();
 sg13g2_fill_2 FILLER_44_1390 ();
 sg13g2_fill_1 FILLER_44_1392 ();
 sg13g2_fill_1 FILLER_44_1429 ();
 sg13g2_fill_1 FILLER_44_1466 ();
 sg13g2_fill_2 FILLER_44_1487 ();
 sg13g2_fill_2 FILLER_44_1525 ();
 sg13g2_decap_4 FILLER_44_1532 ();
 sg13g2_fill_2 FILLER_44_1546 ();
 sg13g2_fill_2 FILLER_44_1573 ();
 sg13g2_fill_1 FILLER_44_1575 ();
 sg13g2_fill_2 FILLER_44_1605 ();
 sg13g2_fill_2 FILLER_44_1617 ();
 sg13g2_fill_1 FILLER_44_1619 ();
 sg13g2_decap_4 FILLER_44_1715 ();
 sg13g2_fill_2 FILLER_44_1740 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_fill_2 FILLER_45_58 ();
 sg13g2_fill_2 FILLER_45_121 ();
 sg13g2_fill_1 FILLER_45_123 ();
 sg13g2_fill_2 FILLER_45_143 ();
 sg13g2_fill_1 FILLER_45_169 ();
 sg13g2_fill_1 FILLER_45_176 ();
 sg13g2_fill_1 FILLER_45_208 ();
 sg13g2_fill_2 FILLER_45_252 ();
 sg13g2_fill_1 FILLER_45_254 ();
 sg13g2_fill_2 FILLER_45_263 ();
 sg13g2_decap_4 FILLER_45_288 ();
 sg13g2_fill_1 FILLER_45_339 ();
 sg13g2_fill_2 FILLER_45_350 ();
 sg13g2_fill_1 FILLER_45_352 ();
 sg13g2_fill_1 FILLER_45_373 ();
 sg13g2_fill_1 FILLER_45_404 ();
 sg13g2_decap_4 FILLER_45_476 ();
 sg13g2_fill_2 FILLER_45_484 ();
 sg13g2_decap_4 FILLER_45_513 ();
 sg13g2_fill_1 FILLER_45_517 ();
 sg13g2_fill_1 FILLER_45_535 ();
 sg13g2_fill_1 FILLER_45_544 ();
 sg13g2_fill_1 FILLER_45_646 ();
 sg13g2_fill_2 FILLER_45_666 ();
 sg13g2_fill_1 FILLER_45_681 ();
 sg13g2_decap_4 FILLER_45_695 ();
 sg13g2_fill_1 FILLER_45_743 ();
 sg13g2_decap_8 FILLER_45_770 ();
 sg13g2_fill_1 FILLER_45_777 ();
 sg13g2_fill_2 FILLER_45_856 ();
 sg13g2_decap_4 FILLER_45_883 ();
 sg13g2_fill_2 FILLER_45_923 ();
 sg13g2_fill_1 FILLER_45_925 ();
 sg13g2_fill_1 FILLER_45_931 ();
 sg13g2_decap_4 FILLER_45_954 ();
 sg13g2_fill_1 FILLER_45_994 ();
 sg13g2_fill_2 FILLER_45_1030 ();
 sg13g2_fill_1 FILLER_45_1036 ();
 sg13g2_fill_2 FILLER_45_1076 ();
 sg13g2_fill_2 FILLER_45_1088 ();
 sg13g2_fill_2 FILLER_45_1104 ();
 sg13g2_fill_1 FILLER_45_1130 ();
 sg13g2_fill_2 FILLER_45_1145 ();
 sg13g2_fill_1 FILLER_45_1147 ();
 sg13g2_fill_2 FILLER_45_1166 ();
 sg13g2_fill_1 FILLER_45_1168 ();
 sg13g2_fill_2 FILLER_45_1192 ();
 sg13g2_decap_8 FILLER_45_1198 ();
 sg13g2_fill_1 FILLER_45_1205 ();
 sg13g2_fill_2 FILLER_45_1227 ();
 sg13g2_fill_2 FILLER_45_1271 ();
 sg13g2_fill_2 FILLER_45_1287 ();
 sg13g2_fill_2 FILLER_45_1294 ();
 sg13g2_fill_1 FILLER_45_1296 ();
 sg13g2_fill_1 FILLER_45_1336 ();
 sg13g2_fill_2 FILLER_45_1351 ();
 sg13g2_fill_2 FILLER_45_1423 ();
 sg13g2_fill_1 FILLER_45_1437 ();
 sg13g2_decap_8 FILLER_45_1442 ();
 sg13g2_fill_2 FILLER_45_1449 ();
 sg13g2_fill_2 FILLER_45_1464 ();
 sg13g2_fill_1 FILLER_45_1480 ();
 sg13g2_decap_4 FILLER_45_1486 ();
 sg13g2_fill_2 FILLER_45_1490 ();
 sg13g2_fill_2 FILLER_45_1600 ();
 sg13g2_fill_2 FILLER_45_1610 ();
 sg13g2_fill_1 FILLER_45_1612 ();
 sg13g2_fill_1 FILLER_45_1632 ();
 sg13g2_fill_1 FILLER_45_1639 ();
 sg13g2_fill_2 FILLER_45_1650 ();
 sg13g2_fill_1 FILLER_45_1652 ();
 sg13g2_fill_1 FILLER_45_1715 ();
 sg13g2_fill_2 FILLER_45_1766 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_95 ();
 sg13g2_fill_2 FILLER_46_102 ();
 sg13g2_fill_1 FILLER_46_104 ();
 sg13g2_fill_1 FILLER_46_140 ();
 sg13g2_fill_2 FILLER_46_187 ();
 sg13g2_fill_1 FILLER_46_189 ();
 sg13g2_fill_1 FILLER_46_214 ();
 sg13g2_fill_1 FILLER_46_261 ();
 sg13g2_fill_1 FILLER_46_279 ();
 sg13g2_fill_2 FILLER_46_306 ();
 sg13g2_fill_2 FILLER_46_350 ();
 sg13g2_fill_2 FILLER_46_368 ();
 sg13g2_fill_1 FILLER_46_370 ();
 sg13g2_fill_2 FILLER_46_406 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_fill_2 FILLER_46_435 ();
 sg13g2_fill_1 FILLER_46_437 ();
 sg13g2_fill_2 FILLER_46_474 ();
 sg13g2_decap_4 FILLER_46_489 ();
 sg13g2_fill_2 FILLER_46_566 ();
 sg13g2_fill_1 FILLER_46_618 ();
 sg13g2_fill_1 FILLER_46_689 ();
 sg13g2_fill_1 FILLER_46_736 ();
 sg13g2_fill_1 FILLER_46_750 ();
 sg13g2_fill_1 FILLER_46_774 ();
 sg13g2_decap_4 FILLER_46_811 ();
 sg13g2_decap_4 FILLER_46_823 ();
 sg13g2_fill_1 FILLER_46_827 ();
 sg13g2_fill_2 FILLER_46_845 ();
 sg13g2_fill_1 FILLER_46_847 ();
 sg13g2_decap_8 FILLER_46_892 ();
 sg13g2_fill_1 FILLER_46_899 ();
 sg13g2_fill_2 FILLER_46_926 ();
 sg13g2_fill_2 FILLER_46_954 ();
 sg13g2_fill_1 FILLER_46_993 ();
 sg13g2_decap_4 FILLER_46_1007 ();
 sg13g2_fill_1 FILLER_46_1051 ();
 sg13g2_fill_1 FILLER_46_1075 ();
 sg13g2_fill_2 FILLER_46_1086 ();
 sg13g2_fill_1 FILLER_46_1088 ();
 sg13g2_fill_2 FILLER_46_1181 ();
 sg13g2_fill_2 FILLER_46_1225 ();
 sg13g2_fill_1 FILLER_46_1227 ();
 sg13g2_fill_2 FILLER_46_1232 ();
 sg13g2_fill_1 FILLER_46_1238 ();
 sg13g2_fill_1 FILLER_46_1243 ();
 sg13g2_decap_4 FILLER_46_1257 ();
 sg13g2_fill_1 FILLER_46_1269 ();
 sg13g2_decap_4 FILLER_46_1274 ();
 sg13g2_fill_2 FILLER_46_1283 ();
 sg13g2_fill_1 FILLER_46_1285 ();
 sg13g2_fill_1 FILLER_46_1330 ();
 sg13g2_fill_2 FILLER_46_1354 ();
 sg13g2_fill_1 FILLER_46_1356 ();
 sg13g2_fill_2 FILLER_46_1366 ();
 sg13g2_fill_1 FILLER_46_1382 ();
 sg13g2_fill_2 FILLER_46_1436 ();
 sg13g2_fill_1 FILLER_46_1438 ();
 sg13g2_fill_1 FILLER_46_1453 ();
 sg13g2_fill_1 FILLER_46_1480 ();
 sg13g2_decap_4 FILLER_46_1489 ();
 sg13g2_fill_2 FILLER_46_1501 ();
 sg13g2_decap_4 FILLER_46_1516 ();
 sg13g2_fill_2 FILLER_46_1520 ();
 sg13g2_fill_1 FILLER_46_1536 ();
 sg13g2_fill_1 FILLER_46_1569 ();
 sg13g2_fill_2 FILLER_46_1579 ();
 sg13g2_fill_2 FILLER_46_1591 ();
 sg13g2_fill_2 FILLER_46_1619 ();
 sg13g2_fill_1 FILLER_46_1682 ();
 sg13g2_fill_1 FILLER_46_1692 ();
 sg13g2_fill_1 FILLER_46_1702 ();
 sg13g2_fill_1 FILLER_46_1729 ();
 sg13g2_fill_1 FILLER_46_1767 ();
 sg13g2_fill_2 FILLER_47_26 ();
 sg13g2_fill_2 FILLER_47_54 ();
 sg13g2_fill_1 FILLER_47_56 ();
 sg13g2_fill_2 FILLER_47_192 ();
 sg13g2_fill_1 FILLER_47_194 ();
 sg13g2_fill_1 FILLER_47_204 ();
 sg13g2_fill_1 FILLER_47_244 ();
 sg13g2_fill_2 FILLER_47_276 ();
 sg13g2_fill_1 FILLER_47_278 ();
 sg13g2_fill_2 FILLER_47_330 ();
 sg13g2_fill_2 FILLER_47_394 ();
 sg13g2_fill_1 FILLER_47_396 ();
 sg13g2_fill_1 FILLER_47_415 ();
 sg13g2_fill_2 FILLER_47_471 ();
 sg13g2_fill_2 FILLER_47_514 ();
 sg13g2_fill_1 FILLER_47_516 ();
 sg13g2_fill_1 FILLER_47_531 ();
 sg13g2_fill_2 FILLER_47_568 ();
 sg13g2_fill_1 FILLER_47_570 ();
 sg13g2_fill_2 FILLER_47_607 ();
 sg13g2_fill_1 FILLER_47_609 ();
 sg13g2_fill_1 FILLER_47_623 ();
 sg13g2_fill_2 FILLER_47_643 ();
 sg13g2_fill_2 FILLER_47_649 ();
 sg13g2_fill_1 FILLER_47_651 ();
 sg13g2_fill_1 FILLER_47_662 ();
 sg13g2_fill_1 FILLER_47_676 ();
 sg13g2_fill_2 FILLER_47_687 ();
 sg13g2_fill_1 FILLER_47_689 ();
 sg13g2_fill_2 FILLER_47_726 ();
 sg13g2_fill_2 FILLER_47_743 ();
 sg13g2_fill_2 FILLER_47_775 ();
 sg13g2_fill_1 FILLER_47_795 ();
 sg13g2_decap_4 FILLER_47_800 ();
 sg13g2_fill_1 FILLER_47_804 ();
 sg13g2_fill_1 FILLER_47_859 ();
 sg13g2_fill_1 FILLER_47_891 ();
 sg13g2_fill_1 FILLER_47_906 ();
 sg13g2_fill_1 FILLER_47_921 ();
 sg13g2_fill_2 FILLER_47_955 ();
 sg13g2_fill_2 FILLER_47_1029 ();
 sg13g2_fill_1 FILLER_47_1031 ();
 sg13g2_fill_2 FILLER_47_1056 ();
 sg13g2_fill_1 FILLER_47_1058 ();
 sg13g2_decap_4 FILLER_47_1089 ();
 sg13g2_fill_2 FILLER_47_1093 ();
 sg13g2_fill_1 FILLER_47_1104 ();
 sg13g2_fill_2 FILLER_47_1114 ();
 sg13g2_fill_2 FILLER_47_1154 ();
 sg13g2_fill_2 FILLER_47_1161 ();
 sg13g2_fill_1 FILLER_47_1163 ();
 sg13g2_fill_2 FILLER_47_1173 ();
 sg13g2_fill_1 FILLER_47_1175 ();
 sg13g2_fill_2 FILLER_47_1210 ();
 sg13g2_fill_1 FILLER_47_1212 ();
 sg13g2_decap_4 FILLER_47_1285 ();
 sg13g2_fill_2 FILLER_47_1289 ();
 sg13g2_decap_4 FILLER_47_1300 ();
 sg13g2_fill_2 FILLER_47_1304 ();
 sg13g2_decap_4 FILLER_47_1319 ();
 sg13g2_fill_1 FILLER_47_1405 ();
 sg13g2_fill_2 FILLER_47_1412 ();
 sg13g2_fill_1 FILLER_47_1414 ();
 sg13g2_fill_2 FILLER_47_1475 ();
 sg13g2_fill_1 FILLER_47_1477 ();
 sg13g2_fill_2 FILLER_47_1525 ();
 sg13g2_fill_1 FILLER_47_1527 ();
 sg13g2_fill_2 FILLER_47_1603 ();
 sg13g2_fill_1 FILLER_47_1605 ();
 sg13g2_fill_2 FILLER_47_1630 ();
 sg13g2_fill_1 FILLER_47_1632 ();
 sg13g2_fill_2 FILLER_47_1647 ();
 sg13g2_fill_1 FILLER_47_1649 ();
 sg13g2_fill_2 FILLER_47_1699 ();
 sg13g2_fill_1 FILLER_47_1701 ();
 sg13g2_fill_2 FILLER_47_1716 ();
 sg13g2_fill_2 FILLER_47_1727 ();
 sg13g2_fill_2 FILLER_47_1765 ();
 sg13g2_fill_1 FILLER_47_1767 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_34 ();
 sg13g2_fill_1 FILLER_48_36 ();
 sg13g2_fill_1 FILLER_48_58 ();
 sg13g2_decap_8 FILLER_48_82 ();
 sg13g2_fill_2 FILLER_48_89 ();
 sg13g2_fill_2 FILLER_48_113 ();
 sg13g2_fill_2 FILLER_48_150 ();
 sg13g2_fill_1 FILLER_48_152 ();
 sg13g2_fill_2 FILLER_48_205 ();
 sg13g2_fill_1 FILLER_48_207 ();
 sg13g2_fill_2 FILLER_48_235 ();
 sg13g2_fill_1 FILLER_48_237 ();
 sg13g2_fill_1 FILLER_48_268 ();
 sg13g2_fill_2 FILLER_48_306 ();
 sg13g2_fill_1 FILLER_48_308 ();
 sg13g2_fill_1 FILLER_48_318 ();
 sg13g2_fill_2 FILLER_48_329 ();
 sg13g2_fill_1 FILLER_48_331 ();
 sg13g2_fill_2 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_fill_1 FILLER_48_409 ();
 sg13g2_fill_2 FILLER_48_445 ();
 sg13g2_fill_1 FILLER_48_447 ();
 sg13g2_fill_1 FILLER_48_478 ();
 sg13g2_fill_2 FILLER_48_489 ();
 sg13g2_fill_2 FILLER_48_531 ();
 sg13g2_fill_1 FILLER_48_533 ();
 sg13g2_fill_1 FILLER_48_552 ();
 sg13g2_fill_2 FILLER_48_571 ();
 sg13g2_fill_2 FILLER_48_624 ();
 sg13g2_fill_1 FILLER_48_655 ();
 sg13g2_fill_2 FILLER_48_708 ();
 sg13g2_fill_2 FILLER_48_719 ();
 sg13g2_fill_2 FILLER_48_780 ();
 sg13g2_fill_1 FILLER_48_782 ();
 sg13g2_fill_2 FILLER_48_798 ();
 sg13g2_fill_2 FILLER_48_826 ();
 sg13g2_fill_2 FILLER_48_841 ();
 sg13g2_fill_1 FILLER_48_859 ();
 sg13g2_decap_4 FILLER_48_896 ();
 sg13g2_fill_2 FILLER_48_900 ();
 sg13g2_fill_2 FILLER_48_946 ();
 sg13g2_fill_2 FILLER_48_958 ();
 sg13g2_fill_1 FILLER_48_960 ();
 sg13g2_fill_2 FILLER_48_971 ();
 sg13g2_fill_1 FILLER_48_1003 ();
 sg13g2_fill_1 FILLER_48_1013 ();
 sg13g2_fill_2 FILLER_48_1066 ();
 sg13g2_fill_1 FILLER_48_1076 ();
 sg13g2_fill_1 FILLER_48_1117 ();
 sg13g2_decap_4 FILLER_48_1133 ();
 sg13g2_fill_1 FILLER_48_1213 ();
 sg13g2_fill_1 FILLER_48_1227 ();
 sg13g2_fill_2 FILLER_48_1266 ();
 sg13g2_decap_8 FILLER_48_1304 ();
 sg13g2_fill_1 FILLER_48_1333 ();
 sg13g2_fill_1 FILLER_48_1387 ();
 sg13g2_fill_1 FILLER_48_1414 ();
 sg13g2_fill_2 FILLER_48_1423 ();
 sg13g2_fill_1 FILLER_48_1497 ();
 sg13g2_fill_2 FILLER_48_1528 ();
 sg13g2_fill_1 FILLER_48_1548 ();
 sg13g2_fill_1 FILLER_48_1588 ();
 sg13g2_fill_1 FILLER_48_1644 ();
 sg13g2_fill_1 FILLER_48_1659 ();
 sg13g2_fill_2 FILLER_48_1701 ();
 sg13g2_fill_2 FILLER_48_1738 ();
 sg13g2_fill_2 FILLER_48_1766 ();
 sg13g2_fill_2 FILLER_49_50 ();
 sg13g2_fill_1 FILLER_49_52 ();
 sg13g2_fill_2 FILLER_49_150 ();
 sg13g2_fill_1 FILLER_49_152 ();
 sg13g2_fill_2 FILLER_49_180 ();
 sg13g2_fill_2 FILLER_49_212 ();
 sg13g2_fill_1 FILLER_49_214 ();
 sg13g2_fill_2 FILLER_49_325 ();
 sg13g2_fill_2 FILLER_49_334 ();
 sg13g2_fill_1 FILLER_49_336 ();
 sg13g2_fill_2 FILLER_49_347 ();
 sg13g2_fill_1 FILLER_49_374 ();
 sg13g2_fill_2 FILLER_49_400 ();
 sg13g2_fill_1 FILLER_49_428 ();
 sg13g2_fill_1 FILLER_49_525 ();
 sg13g2_fill_1 FILLER_49_576 ();
 sg13g2_fill_2 FILLER_49_602 ();
 sg13g2_fill_1 FILLER_49_624 ();
 sg13g2_fill_2 FILLER_49_636 ();
 sg13g2_decap_8 FILLER_49_675 ();
 sg13g2_decap_8 FILLER_49_682 ();
 sg13g2_fill_2 FILLER_49_708 ();
 sg13g2_fill_2 FILLER_49_769 ();
 sg13g2_fill_2 FILLER_49_785 ();
 sg13g2_fill_2 FILLER_49_848 ();
 sg13g2_fill_2 FILLER_49_888 ();
 sg13g2_fill_2 FILLER_49_922 ();
 sg13g2_fill_1 FILLER_49_983 ();
 sg13g2_fill_2 FILLER_49_1064 ();
 sg13g2_fill_1 FILLER_49_1066 ();
 sg13g2_fill_2 FILLER_49_1085 ();
 sg13g2_fill_1 FILLER_49_1087 ();
 sg13g2_fill_1 FILLER_49_1128 ();
 sg13g2_fill_2 FILLER_49_1200 ();
 sg13g2_fill_1 FILLER_49_1202 ();
 sg13g2_fill_2 FILLER_49_1208 ();
 sg13g2_fill_1 FILLER_49_1269 ();
 sg13g2_fill_2 FILLER_49_1298 ();
 sg13g2_decap_4 FILLER_49_1329 ();
 sg13g2_decap_4 FILLER_49_1364 ();
 sg13g2_fill_2 FILLER_49_1368 ();
 sg13g2_fill_2 FILLER_49_1379 ();
 sg13g2_fill_1 FILLER_49_1381 ();
 sg13g2_fill_1 FILLER_49_1445 ();
 sg13g2_fill_1 FILLER_49_1459 ();
 sg13g2_fill_2 FILLER_49_1479 ();
 sg13g2_fill_2 FILLER_49_1501 ();
 sg13g2_fill_1 FILLER_49_1503 ();
 sg13g2_fill_2 FILLER_49_1538 ();
 sg13g2_fill_1 FILLER_49_1540 ();
 sg13g2_fill_2 FILLER_49_1560 ();
 sg13g2_fill_1 FILLER_49_1598 ();
 sg13g2_fill_2 FILLER_49_1624 ();
 sg13g2_fill_1 FILLER_49_1626 ();
 sg13g2_fill_1 FILLER_49_1661 ();
 sg13g2_fill_1 FILLER_49_1667 ();
 sg13g2_decap_4 FILLER_49_1700 ();
 sg13g2_fill_1 FILLER_49_1704 ();
 sg13g2_fill_2 FILLER_49_1746 ();
 sg13g2_fill_1 FILLER_49_1748 ();
 sg13g2_fill_1 FILLER_49_1767 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_29 ();
 sg13g2_fill_2 FILLER_50_70 ();
 sg13g2_fill_1 FILLER_50_72 ();
 sg13g2_fill_2 FILLER_50_78 ();
 sg13g2_fill_1 FILLER_50_80 ();
 sg13g2_fill_1 FILLER_50_117 ();
 sg13g2_fill_1 FILLER_50_173 ();
 sg13g2_fill_2 FILLER_50_209 ();
 sg13g2_fill_1 FILLER_50_211 ();
 sg13g2_fill_1 FILLER_50_258 ();
 sg13g2_fill_2 FILLER_50_264 ();
 sg13g2_fill_1 FILLER_50_266 ();
 sg13g2_fill_2 FILLER_50_281 ();
 sg13g2_fill_1 FILLER_50_283 ();
 sg13g2_fill_2 FILLER_50_292 ();
 sg13g2_fill_1 FILLER_50_294 ();
 sg13g2_fill_2 FILLER_50_322 ();
 sg13g2_fill_2 FILLER_50_332 ();
 sg13g2_fill_2 FILLER_50_343 ();
 sg13g2_fill_1 FILLER_50_345 ();
 sg13g2_fill_2 FILLER_50_500 ();
 sg13g2_decap_4 FILLER_50_545 ();
 sg13g2_fill_1 FILLER_50_549 ();
 sg13g2_decap_4 FILLER_50_574 ();
 sg13g2_fill_1 FILLER_50_578 ();
 sg13g2_decap_8 FILLER_50_666 ();
 sg13g2_fill_2 FILLER_50_673 ();
 sg13g2_fill_2 FILLER_50_685 ();
 sg13g2_fill_1 FILLER_50_687 ();
 sg13g2_fill_1 FILLER_50_692 ();
 sg13g2_fill_1 FILLER_50_777 ();
 sg13g2_fill_2 FILLER_50_787 ();
 sg13g2_fill_2 FILLER_50_804 ();
 sg13g2_fill_2 FILLER_50_820 ();
 sg13g2_fill_2 FILLER_50_832 ();
 sg13g2_fill_2 FILLER_50_843 ();
 sg13g2_fill_2 FILLER_50_850 ();
 sg13g2_fill_2 FILLER_50_888 ();
 sg13g2_fill_1 FILLER_50_890 ();
 sg13g2_fill_1 FILLER_50_936 ();
 sg13g2_fill_2 FILLER_50_958 ();
 sg13g2_fill_1 FILLER_50_960 ();
 sg13g2_fill_2 FILLER_50_1016 ();
 sg13g2_fill_1 FILLER_50_1028 ();
 sg13g2_fill_2 FILLER_50_1127 ();
 sg13g2_fill_2 FILLER_50_1161 ();
 sg13g2_fill_2 FILLER_50_1227 ();
 sg13g2_fill_1 FILLER_50_1229 ();
 sg13g2_fill_2 FILLER_50_1269 ();
 sg13g2_fill_1 FILLER_50_1271 ();
 sg13g2_decap_4 FILLER_50_1308 ();
 sg13g2_fill_2 FILLER_50_1409 ();
 sg13g2_fill_1 FILLER_50_1411 ();
 sg13g2_decap_4 FILLER_50_1540 ();
 sg13g2_fill_1 FILLER_50_1593 ();
 sg13g2_fill_2 FILLER_50_1602 ();
 sg13g2_decap_4 FILLER_50_1619 ();
 sg13g2_fill_2 FILLER_50_1654 ();
 sg13g2_fill_1 FILLER_50_1656 ();
 sg13g2_fill_2 FILLER_50_1688 ();
 sg13g2_fill_2 FILLER_50_1716 ();
 sg13g2_fill_1 FILLER_50_1718 ();
 sg13g2_fill_1 FILLER_50_1728 ();
 sg13g2_fill_2 FILLER_50_1759 ();
 sg13g2_fill_1 FILLER_50_1761 ();
 sg13g2_fill_2 FILLER_50_1766 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_6 ();
 sg13g2_fill_1 FILLER_51_78 ();
 sg13g2_fill_2 FILLER_51_92 ();
 sg13g2_fill_1 FILLER_51_94 ();
 sg13g2_fill_2 FILLER_51_157 ();
 sg13g2_fill_2 FILLER_51_178 ();
 sg13g2_fill_2 FILLER_51_184 ();
 sg13g2_fill_1 FILLER_51_186 ();
 sg13g2_fill_2 FILLER_51_217 ();
 sg13g2_fill_1 FILLER_51_219 ();
 sg13g2_fill_1 FILLER_51_246 ();
 sg13g2_fill_1 FILLER_51_302 ();
 sg13g2_fill_1 FILLER_51_331 ();
 sg13g2_decap_4 FILLER_51_342 ();
 sg13g2_fill_2 FILLER_51_356 ();
 sg13g2_fill_1 FILLER_51_358 ();
 sg13g2_fill_1 FILLER_51_395 ();
 sg13g2_decap_8 FILLER_51_521 ();
 sg13g2_fill_1 FILLER_51_528 ();
 sg13g2_fill_2 FILLER_51_555 ();
 sg13g2_fill_1 FILLER_51_557 ();
 sg13g2_fill_1 FILLER_51_580 ();
 sg13g2_fill_1 FILLER_51_614 ();
 sg13g2_decap_8 FILLER_51_703 ();
 sg13g2_fill_1 FILLER_51_757 ();
 sg13g2_fill_2 FILLER_51_762 ();
 sg13g2_fill_2 FILLER_51_795 ();
 sg13g2_fill_1 FILLER_51_797 ();
 sg13g2_fill_2 FILLER_51_824 ();
 sg13g2_fill_1 FILLER_51_826 ();
 sg13g2_fill_1 FILLER_51_853 ();
 sg13g2_fill_2 FILLER_51_906 ();
 sg13g2_fill_1 FILLER_51_908 ();
 sg13g2_fill_1 FILLER_51_917 ();
 sg13g2_fill_2 FILLER_51_944 ();
 sg13g2_fill_1 FILLER_51_946 ();
 sg13g2_fill_2 FILLER_51_987 ();
 sg13g2_fill_1 FILLER_51_989 ();
 sg13g2_decap_4 FILLER_51_1016 ();
 sg13g2_fill_2 FILLER_51_1050 ();
 sg13g2_fill_2 FILLER_51_1082 ();
 sg13g2_fill_1 FILLER_51_1084 ();
 sg13g2_fill_2 FILLER_51_1095 ();
 sg13g2_fill_1 FILLER_51_1101 ();
 sg13g2_fill_2 FILLER_51_1137 ();
 sg13g2_fill_1 FILLER_51_1139 ();
 sg13g2_fill_2 FILLER_51_1166 ();
 sg13g2_fill_1 FILLER_51_1208 ();
 sg13g2_fill_2 FILLER_51_1255 ();
 sg13g2_fill_1 FILLER_51_1257 ();
 sg13g2_fill_1 FILLER_51_1312 ();
 sg13g2_fill_2 FILLER_51_1355 ();
 sg13g2_fill_1 FILLER_51_1392 ();
 sg13g2_fill_1 FILLER_51_1475 ();
 sg13g2_fill_1 FILLER_51_1508 ();
 sg13g2_fill_1 FILLER_51_1524 ();
 sg13g2_fill_2 FILLER_51_1530 ();
 sg13g2_fill_1 FILLER_51_1532 ();
 sg13g2_fill_2 FILLER_51_1543 ();
 sg13g2_fill_2 FILLER_51_1566 ();
 sg13g2_fill_1 FILLER_51_1582 ();
 sg13g2_fill_2 FILLER_51_1652 ();
 sg13g2_fill_1 FILLER_51_1654 ();
 sg13g2_fill_1 FILLER_51_1665 ();
 sg13g2_fill_2 FILLER_51_1680 ();
 sg13g2_fill_2 FILLER_51_1705 ();
 sg13g2_fill_2 FILLER_51_1739 ();
 sg13g2_fill_1 FILLER_51_1741 ();
 sg13g2_fill_2 FILLER_52_97 ();
 sg13g2_fill_1 FILLER_52_99 ();
 sg13g2_fill_2 FILLER_52_126 ();
 sg13g2_fill_1 FILLER_52_214 ();
 sg13g2_fill_2 FILLER_52_237 ();
 sg13g2_fill_2 FILLER_52_302 ();
 sg13g2_fill_1 FILLER_52_304 ();
 sg13g2_fill_2 FILLER_52_336 ();
 sg13g2_fill_2 FILLER_52_364 ();
 sg13g2_fill_2 FILLER_52_402 ();
 sg13g2_fill_1 FILLER_52_404 ();
 sg13g2_fill_2 FILLER_52_479 ();
 sg13g2_fill_1 FILLER_52_481 ();
 sg13g2_fill_2 FILLER_52_505 ();
 sg13g2_fill_1 FILLER_52_543 ();
 sg13g2_fill_1 FILLER_52_570 ();
 sg13g2_fill_1 FILLER_52_597 ();
 sg13g2_fill_2 FILLER_52_629 ();
 sg13g2_fill_2 FILLER_52_641 ();
 sg13g2_fill_2 FILLER_52_662 ();
 sg13g2_fill_1 FILLER_52_664 ();
 sg13g2_decap_8 FILLER_52_673 ();
 sg13g2_fill_2 FILLER_52_680 ();
 sg13g2_fill_1 FILLER_52_690 ();
 sg13g2_decap_4 FILLER_52_700 ();
 sg13g2_fill_1 FILLER_52_723 ();
 sg13g2_fill_2 FILLER_52_760 ();
 sg13g2_fill_1 FILLER_52_762 ();
 sg13g2_fill_2 FILLER_52_771 ();
 sg13g2_fill_1 FILLER_52_773 ();
 sg13g2_fill_1 FILLER_52_783 ();
 sg13g2_decap_4 FILLER_52_859 ();
 sg13g2_decap_8 FILLER_52_897 ();
 sg13g2_decap_4 FILLER_52_904 ();
 sg13g2_decap_8 FILLER_52_912 ();
 sg13g2_fill_2 FILLER_52_943 ();
 sg13g2_fill_1 FILLER_52_945 ();
 sg13g2_fill_1 FILLER_52_1012 ();
 sg13g2_fill_2 FILLER_52_1023 ();
 sg13g2_fill_1 FILLER_52_1025 ();
 sg13g2_decap_4 FILLER_52_1081 ();
 sg13g2_fill_2 FILLER_52_1085 ();
 sg13g2_fill_1 FILLER_52_1113 ();
 sg13g2_fill_2 FILLER_52_1128 ();
 sg13g2_fill_1 FILLER_52_1135 ();
 sg13g2_decap_4 FILLER_52_1164 ();
 sg13g2_fill_1 FILLER_52_1168 ();
 sg13g2_fill_2 FILLER_52_1197 ();
 sg13g2_fill_1 FILLER_52_1199 ();
 sg13g2_fill_2 FILLER_52_1259 ();
 sg13g2_fill_2 FILLER_52_1276 ();
 sg13g2_fill_1 FILLER_52_1278 ();
 sg13g2_fill_2 FILLER_52_1297 ();
 sg13g2_fill_1 FILLER_52_1299 ();
 sg13g2_decap_8 FILLER_52_1326 ();
 sg13g2_fill_1 FILLER_52_1333 ();
 sg13g2_fill_2 FILLER_52_1355 ();
 sg13g2_fill_1 FILLER_52_1357 ();
 sg13g2_fill_1 FILLER_52_1559 ();
 sg13g2_fill_2 FILLER_52_1596 ();
 sg13g2_fill_1 FILLER_52_1598 ();
 sg13g2_fill_1 FILLER_52_1692 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_2 ();
 sg13g2_fill_2 FILLER_53_64 ();
 sg13g2_fill_2 FILLER_53_79 ();
 sg13g2_fill_1 FILLER_53_94 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_fill_2 FILLER_53_166 ();
 sg13g2_fill_2 FILLER_53_207 ();
 sg13g2_fill_1 FILLER_53_209 ();
 sg13g2_fill_1 FILLER_53_271 ();
 sg13g2_decap_8 FILLER_53_308 ();
 sg13g2_fill_1 FILLER_53_315 ();
 sg13g2_fill_1 FILLER_53_424 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_decap_4 FILLER_53_440 ();
 sg13g2_fill_1 FILLER_53_444 ();
 sg13g2_fill_1 FILLER_53_476 ();
 sg13g2_fill_1 FILLER_53_480 ();
 sg13g2_decap_8 FILLER_53_486 ();
 sg13g2_fill_2 FILLER_53_493 ();
 sg13g2_fill_1 FILLER_53_495 ();
 sg13g2_fill_1 FILLER_53_580 ();
 sg13g2_decap_4 FILLER_53_594 ();
 sg13g2_fill_2 FILLER_53_611 ();
 sg13g2_fill_1 FILLER_53_613 ();
 sg13g2_fill_2 FILLER_53_618 ();
 sg13g2_fill_1 FILLER_53_634 ();
 sg13g2_decap_4 FILLER_53_670 ();
 sg13g2_fill_2 FILLER_53_674 ();
 sg13g2_fill_1 FILLER_53_681 ();
 sg13g2_fill_2 FILLER_53_716 ();
 sg13g2_decap_8 FILLER_53_737 ();
 sg13g2_fill_2 FILLER_53_744 ();
 sg13g2_fill_2 FILLER_53_765 ();
 sg13g2_fill_1 FILLER_53_767 ();
 sg13g2_fill_2 FILLER_53_773 ();
 sg13g2_fill_2 FILLER_53_789 ();
 sg13g2_fill_1 FILLER_53_791 ();
 sg13g2_fill_2 FILLER_53_815 ();
 sg13g2_fill_1 FILLER_53_817 ();
 sg13g2_fill_2 FILLER_53_836 ();
 sg13g2_decap_4 FILLER_53_868 ();
 sg13g2_fill_1 FILLER_53_872 ();
 sg13g2_fill_1 FILLER_53_923 ();
 sg13g2_fill_2 FILLER_53_959 ();
 sg13g2_fill_2 FILLER_53_975 ();
 sg13g2_fill_1 FILLER_53_977 ();
 sg13g2_fill_1 FILLER_53_1018 ();
 sg13g2_fill_1 FILLER_53_1054 ();
 sg13g2_fill_2 FILLER_53_1079 ();
 sg13g2_fill_1 FILLER_53_1081 ();
 sg13g2_decap_4 FILLER_53_1092 ();
 sg13g2_fill_1 FILLER_53_1096 ();
 sg13g2_fill_1 FILLER_53_1115 ();
 sg13g2_fill_2 FILLER_53_1130 ();
 sg13g2_fill_1 FILLER_53_1132 ();
 sg13g2_fill_2 FILLER_53_1169 ();
 sg13g2_fill_2 FILLER_53_1175 ();
 sg13g2_fill_1 FILLER_53_1177 ();
 sg13g2_fill_2 FILLER_53_1260 ();
 sg13g2_fill_1 FILLER_53_1272 ();
 sg13g2_fill_2 FILLER_53_1308 ();
 sg13g2_decap_4 FILLER_53_1340 ();
 sg13g2_fill_2 FILLER_53_1348 ();
 sg13g2_fill_2 FILLER_53_1410 ();
 sg13g2_fill_1 FILLER_53_1412 ();
 sg13g2_decap_4 FILLER_53_1449 ();
 sg13g2_fill_2 FILLER_53_1453 ();
 sg13g2_fill_1 FILLER_53_1465 ();
 sg13g2_fill_1 FILLER_53_1549 ();
 sg13g2_fill_1 FILLER_53_1608 ();
 sg13g2_fill_2 FILLER_53_1727 ();
 sg13g2_fill_2 FILLER_53_1739 ();
 sg13g2_fill_1 FILLER_53_1741 ();
 sg13g2_fill_1 FILLER_54_30 ();
 sg13g2_fill_1 FILLER_54_71 ();
 sg13g2_fill_1 FILLER_54_98 ();
 sg13g2_fill_1 FILLER_54_140 ();
 sg13g2_fill_2 FILLER_54_176 ();
 sg13g2_fill_1 FILLER_54_178 ();
 sg13g2_fill_1 FILLER_54_268 ();
 sg13g2_fill_2 FILLER_54_278 ();
 sg13g2_fill_2 FILLER_54_289 ();
 sg13g2_fill_1 FILLER_54_291 ();
 sg13g2_fill_1 FILLER_54_301 ();
 sg13g2_fill_2 FILLER_54_353 ();
 sg13g2_fill_1 FILLER_54_355 ();
 sg13g2_fill_2 FILLER_54_360 ();
 sg13g2_fill_1 FILLER_54_362 ();
 sg13g2_fill_2 FILLER_54_388 ();
 sg13g2_fill_1 FILLER_54_450 ();
 sg13g2_fill_1 FILLER_54_480 ();
 sg13g2_fill_2 FILLER_54_560 ();
 sg13g2_fill_1 FILLER_54_562 ();
 sg13g2_fill_1 FILLER_54_579 ();
 sg13g2_fill_1 FILLER_54_608 ();
 sg13g2_fill_1 FILLER_54_620 ();
 sg13g2_decap_4 FILLER_54_661 ();
 sg13g2_decap_4 FILLER_54_681 ();
 sg13g2_fill_1 FILLER_54_691 ();
 sg13g2_decap_4 FILLER_54_696 ();
 sg13g2_fill_1 FILLER_54_700 ();
 sg13g2_fill_1 FILLER_54_720 ();
 sg13g2_fill_2 FILLER_54_737 ();
 sg13g2_fill_2 FILLER_54_765 ();
 sg13g2_decap_4 FILLER_54_803 ();
 sg13g2_fill_2 FILLER_54_807 ();
 sg13g2_fill_1 FILLER_54_835 ();
 sg13g2_decap_4 FILLER_54_913 ();
 sg13g2_fill_2 FILLER_54_944 ();
 sg13g2_fill_1 FILLER_54_946 ();
 sg13g2_fill_1 FILLER_54_1006 ();
 sg13g2_fill_2 FILLER_54_1048 ();
 sg13g2_fill_1 FILLER_54_1050 ();
 sg13g2_decap_4 FILLER_54_1095 ();
 sg13g2_fill_1 FILLER_54_1099 ();
 sg13g2_fill_2 FILLER_54_1160 ();
 sg13g2_fill_2 FILLER_54_1171 ();
 sg13g2_fill_2 FILLER_54_1216 ();
 sg13g2_fill_2 FILLER_54_1294 ();
 sg13g2_fill_1 FILLER_54_1296 ();
 sg13g2_decap_8 FILLER_54_1307 ();
 sg13g2_fill_1 FILLER_54_1314 ();
 sg13g2_decap_4 FILLER_54_1319 ();
 sg13g2_fill_2 FILLER_54_1323 ();
 sg13g2_fill_1 FILLER_54_1329 ();
 sg13g2_fill_2 FILLER_54_1349 ();
 sg13g2_fill_1 FILLER_54_1351 ();
 sg13g2_fill_2 FILLER_54_1366 ();
 sg13g2_decap_8 FILLER_54_1425 ();
 sg13g2_fill_2 FILLER_54_1432 ();
 sg13g2_fill_1 FILLER_54_1434 ();
 sg13g2_fill_2 FILLER_54_1440 ();
 sg13g2_fill_1 FILLER_54_1483 ();
 sg13g2_fill_1 FILLER_54_1489 ();
 sg13g2_fill_2 FILLER_54_1542 ();
 sg13g2_fill_1 FILLER_54_1580 ();
 sg13g2_decap_4 FILLER_54_1589 ();
 sg13g2_fill_2 FILLER_54_1593 ();
 sg13g2_fill_1 FILLER_54_1696 ();
 sg13g2_fill_2 FILLER_54_1721 ();
 sg13g2_fill_2 FILLER_54_1766 ();
 sg13g2_fill_2 FILLER_55_60 ();
 sg13g2_fill_2 FILLER_55_80 ();
 sg13g2_fill_1 FILLER_55_95 ();
 sg13g2_fill_2 FILLER_55_139 ();
 sg13g2_fill_1 FILLER_55_159 ();
 sg13g2_fill_2 FILLER_55_205 ();
 sg13g2_fill_2 FILLER_55_217 ();
 sg13g2_fill_1 FILLER_55_219 ();
 sg13g2_fill_1 FILLER_55_260 ();
 sg13g2_fill_2 FILLER_55_297 ();
 sg13g2_fill_1 FILLER_55_299 ();
 sg13g2_fill_2 FILLER_55_316 ();
 sg13g2_fill_1 FILLER_55_334 ();
 sg13g2_fill_2 FILLER_55_390 ();
 sg13g2_decap_8 FILLER_55_418 ();
 sg13g2_decap_8 FILLER_55_425 ();
 sg13g2_fill_2 FILLER_55_432 ();
 sg13g2_fill_1 FILLER_55_462 ();
 sg13g2_decap_4 FILLER_55_467 ();
 sg13g2_fill_2 FILLER_55_495 ();
 sg13g2_fill_1 FILLER_55_497 ();
 sg13g2_decap_4 FILLER_55_537 ();
 sg13g2_fill_1 FILLER_55_541 ();
 sg13g2_fill_1 FILLER_55_554 ();
 sg13g2_decap_4 FILLER_55_560 ();
 sg13g2_decap_4 FILLER_55_572 ();
 sg13g2_fill_1 FILLER_55_576 ();
 sg13g2_fill_2 FILLER_55_614 ();
 sg13g2_decap_4 FILLER_55_650 ();
 sg13g2_fill_2 FILLER_55_654 ();
 sg13g2_fill_1 FILLER_55_664 ();
 sg13g2_fill_2 FILLER_55_742 ();
 sg13g2_fill_1 FILLER_55_744 ();
 sg13g2_fill_1 FILLER_55_771 ();
 sg13g2_fill_1 FILLER_55_787 ();
 sg13g2_fill_2 FILLER_55_798 ();
 sg13g2_fill_1 FILLER_55_800 ();
 sg13g2_fill_1 FILLER_55_807 ();
 sg13g2_decap_4 FILLER_55_885 ();
 sg13g2_fill_2 FILLER_55_915 ();
 sg13g2_fill_2 FILLER_55_936 ();
 sg13g2_fill_1 FILLER_55_938 ();
 sg13g2_fill_1 FILLER_55_943 ();
 sg13g2_fill_1 FILLER_55_953 ();
 sg13g2_decap_4 FILLER_55_984 ();
 sg13g2_fill_1 FILLER_55_988 ();
 sg13g2_fill_2 FILLER_55_1019 ();
 sg13g2_fill_1 FILLER_55_1026 ();
 sg13g2_fill_2 FILLER_55_1057 ();
 sg13g2_decap_4 FILLER_55_1101 ();
 sg13g2_fill_2 FILLER_55_1110 ();
 sg13g2_fill_1 FILLER_55_1112 ();
 sg13g2_fill_1 FILLER_55_1121 ();
 sg13g2_fill_1 FILLER_55_1160 ();
 sg13g2_fill_1 FILLER_55_1197 ();
 sg13g2_fill_1 FILLER_55_1224 ();
 sg13g2_fill_2 FILLER_55_1235 ();
 sg13g2_fill_1 FILLER_55_1237 ();
 sg13g2_fill_2 FILLER_55_1272 ();
 sg13g2_fill_1 FILLER_55_1274 ();
 sg13g2_fill_2 FILLER_55_1284 ();
 sg13g2_fill_1 FILLER_55_1308 ();
 sg13g2_decap_4 FILLER_55_1335 ();
 sg13g2_fill_2 FILLER_55_1339 ();
 sg13g2_fill_1 FILLER_55_1409 ();
 sg13g2_fill_1 FILLER_55_1451 ();
 sg13g2_fill_1 FILLER_55_1466 ();
 sg13g2_fill_2 FILLER_55_1489 ();
 sg13g2_fill_1 FILLER_55_1491 ();
 sg13g2_fill_2 FILLER_55_1515 ();
 sg13g2_fill_1 FILLER_55_1553 ();
 sg13g2_fill_2 FILLER_55_1564 ();
 sg13g2_fill_1 FILLER_55_1566 ();
 sg13g2_fill_2 FILLER_55_1641 ();
 sg13g2_fill_2 FILLER_55_1693 ();
 sg13g2_fill_1 FILLER_55_1695 ();
 sg13g2_fill_1 FILLER_55_1710 ();
 sg13g2_fill_1 FILLER_55_1737 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_167 ();
 sg13g2_fill_1 FILLER_56_195 ();
 sg13g2_fill_1 FILLER_56_243 ();
 sg13g2_fill_2 FILLER_56_363 ();
 sg13g2_fill_2 FILLER_56_405 ();
 sg13g2_fill_2 FILLER_56_423 ();
 sg13g2_fill_1 FILLER_56_425 ();
 sg13g2_decap_8 FILLER_56_434 ();
 sg13g2_decap_4 FILLER_56_441 ();
 sg13g2_fill_1 FILLER_56_445 ();
 sg13g2_fill_2 FILLER_56_507 ();
 sg13g2_fill_1 FILLER_56_514 ();
 sg13g2_fill_2 FILLER_56_541 ();
 sg13g2_fill_1 FILLER_56_543 ();
 sg13g2_decap_4 FILLER_56_579 ();
 sg13g2_fill_1 FILLER_56_604 ();
 sg13g2_fill_2 FILLER_56_620 ();
 sg13g2_decap_4 FILLER_56_628 ();
 sg13g2_decap_8 FILLER_56_672 ();
 sg13g2_decap_4 FILLER_56_679 ();
 sg13g2_fill_1 FILLER_56_683 ();
 sg13g2_fill_2 FILLER_56_688 ();
 sg13g2_fill_1 FILLER_56_690 ();
 sg13g2_fill_2 FILLER_56_704 ();
 sg13g2_decap_4 FILLER_56_733 ();
 sg13g2_decap_4 FILLER_56_742 ();
 sg13g2_fill_2 FILLER_56_753 ();
 sg13g2_fill_2 FILLER_56_761 ();
 sg13g2_fill_2 FILLER_56_769 ();
 sg13g2_fill_2 FILLER_56_779 ();
 sg13g2_fill_1 FILLER_56_836 ();
 sg13g2_fill_1 FILLER_56_847 ();
 sg13g2_fill_1 FILLER_56_910 ();
 sg13g2_fill_1 FILLER_56_974 ();
 sg13g2_fill_1 FILLER_56_1002 ();
 sg13g2_fill_2 FILLER_56_1023 ();
 sg13g2_fill_1 FILLER_56_1025 ();
 sg13g2_decap_8 FILLER_56_1062 ();
 sg13g2_fill_1 FILLER_56_1069 ();
 sg13g2_fill_2 FILLER_56_1078 ();
 sg13g2_fill_2 FILLER_56_1086 ();
 sg13g2_fill_1 FILLER_56_1088 ();
 sg13g2_fill_1 FILLER_56_1144 ();
 sg13g2_fill_2 FILLER_56_1164 ();
 sg13g2_fill_1 FILLER_56_1166 ();
 sg13g2_fill_1 FILLER_56_1188 ();
 sg13g2_fill_2 FILLER_56_1212 ();
 sg13g2_fill_1 FILLER_56_1222 ();
 sg13g2_fill_2 FILLER_56_1227 ();
 sg13g2_fill_2 FILLER_56_1265 ();
 sg13g2_fill_1 FILLER_56_1267 ();
 sg13g2_fill_2 FILLER_56_1334 ();
 sg13g2_fill_1 FILLER_56_1336 ();
 sg13g2_fill_1 FILLER_56_1370 ();
 sg13g2_fill_1 FILLER_56_1425 ();
 sg13g2_fill_1 FILLER_56_1439 ();
 sg13g2_fill_2 FILLER_56_1485 ();
 sg13g2_fill_2 FILLER_56_1563 ();
 sg13g2_fill_2 FILLER_56_1575 ();
 sg13g2_fill_1 FILLER_56_1590 ();
 sg13g2_fill_2 FILLER_56_1605 ();
 sg13g2_fill_1 FILLER_56_1648 ();
 sg13g2_fill_1 FILLER_56_1731 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_52 ();
 sg13g2_fill_2 FILLER_57_99 ();
 sg13g2_fill_1 FILLER_57_101 ();
 sg13g2_fill_2 FILLER_57_116 ();
 sg13g2_fill_1 FILLER_57_118 ();
 sg13g2_fill_2 FILLER_57_124 ();
 sg13g2_fill_2 FILLER_57_131 ();
 sg13g2_fill_1 FILLER_57_138 ();
 sg13g2_fill_2 FILLER_57_220 ();
 sg13g2_fill_1 FILLER_57_222 ();
 sg13g2_fill_2 FILLER_57_232 ();
 sg13g2_fill_1 FILLER_57_234 ();
 sg13g2_fill_2 FILLER_57_288 ();
 sg13g2_fill_2 FILLER_57_375 ();
 sg13g2_fill_1 FILLER_57_377 ();
 sg13g2_fill_1 FILLER_57_470 ();
 sg13g2_fill_1 FILLER_57_493 ();
 sg13g2_fill_1 FILLER_57_509 ();
 sg13g2_fill_2 FILLER_57_520 ();
 sg13g2_fill_2 FILLER_57_549 ();
 sg13g2_fill_2 FILLER_57_582 ();
 sg13g2_fill_1 FILLER_57_584 ();
 sg13g2_fill_2 FILLER_57_627 ();
 sg13g2_fill_1 FILLER_57_662 ();
 sg13g2_decap_4 FILLER_57_667 ();
 sg13g2_fill_1 FILLER_57_671 ();
 sg13g2_fill_2 FILLER_57_680 ();
 sg13g2_fill_2 FILLER_57_704 ();
 sg13g2_fill_2 FILLER_57_719 ();
 sg13g2_decap_4 FILLER_57_738 ();
 sg13g2_decap_4 FILLER_57_754 ();
 sg13g2_fill_1 FILLER_57_758 ();
 sg13g2_decap_4 FILLER_57_770 ();
 sg13g2_fill_2 FILLER_57_774 ();
 sg13g2_fill_1 FILLER_57_788 ();
 sg13g2_decap_4 FILLER_57_795 ();
 sg13g2_fill_2 FILLER_57_799 ();
 sg13g2_fill_1 FILLER_57_821 ();
 sg13g2_fill_2 FILLER_57_828 ();
 sg13g2_fill_1 FILLER_57_830 ();
 sg13g2_decap_4 FILLER_57_841 ();
 sg13g2_decap_4 FILLER_57_867 ();
 sg13g2_fill_2 FILLER_57_871 ();
 sg13g2_fill_1 FILLER_57_883 ();
 sg13g2_fill_1 FILLER_57_920 ();
 sg13g2_fill_2 FILLER_57_939 ();
 sg13g2_fill_2 FILLER_57_950 ();
 sg13g2_fill_1 FILLER_57_952 ();
 sg13g2_fill_2 FILLER_57_967 ();
 sg13g2_fill_2 FILLER_57_999 ();
 sg13g2_fill_1 FILLER_57_1028 ();
 sg13g2_fill_2 FILLER_57_1047 ();
 sg13g2_fill_1 FILLER_57_1049 ();
 sg13g2_fill_2 FILLER_57_1067 ();
 sg13g2_fill_2 FILLER_57_1140 ();
 sg13g2_decap_4 FILLER_57_1184 ();
 sg13g2_fill_1 FILLER_57_1329 ();
 sg13g2_fill_1 FILLER_57_1340 ();
 sg13g2_fill_1 FILLER_57_1389 ();
 sg13g2_fill_2 FILLER_57_1414 ();
 sg13g2_fill_2 FILLER_57_1447 ();
 sg13g2_decap_4 FILLER_57_1511 ();
 sg13g2_fill_2 FILLER_57_1515 ();
 sg13g2_decap_4 FILLER_57_1525 ();
 sg13g2_fill_1 FILLER_57_1529 ();
 sg13g2_fill_1 FILLER_57_1540 ();
 sg13g2_fill_1 FILLER_57_1581 ();
 sg13g2_fill_2 FILLER_57_1630 ();
 sg13g2_fill_1 FILLER_57_1632 ();
 sg13g2_fill_1 FILLER_57_1665 ();
 sg13g2_fill_1 FILLER_57_1687 ();
 sg13g2_fill_2 FILLER_57_1710 ();
 sg13g2_fill_1 FILLER_57_1712 ();
 sg13g2_fill_1 FILLER_57_1722 ();
 sg13g2_fill_2 FILLER_57_1765 ();
 sg13g2_fill_1 FILLER_57_1767 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_86 ();
 sg13g2_fill_1 FILLER_58_96 ();
 sg13g2_fill_2 FILLER_58_146 ();
 sg13g2_fill_1 FILLER_58_148 ();
 sg13g2_fill_2 FILLER_58_162 ();
 sg13g2_fill_2 FILLER_58_172 ();
 sg13g2_fill_1 FILLER_58_178 ();
 sg13g2_fill_2 FILLER_58_237 ();
 sg13g2_fill_1 FILLER_58_336 ();
 sg13g2_fill_2 FILLER_58_356 ();
 sg13g2_decap_8 FILLER_58_413 ();
 sg13g2_decap_8 FILLER_58_429 ();
 sg13g2_fill_2 FILLER_58_436 ();
 sg13g2_fill_1 FILLER_58_438 ();
 sg13g2_fill_2 FILLER_58_443 ();
 sg13g2_fill_1 FILLER_58_455 ();
 sg13g2_fill_1 FILLER_58_497 ();
 sg13g2_fill_1 FILLER_58_506 ();
 sg13g2_fill_2 FILLER_58_533 ();
 sg13g2_fill_2 FILLER_58_595 ();
 sg13g2_fill_1 FILLER_58_597 ();
 sg13g2_fill_1 FILLER_58_633 ();
 sg13g2_fill_1 FILLER_58_705 ();
 sg13g2_decap_8 FILLER_58_741 ();
 sg13g2_fill_2 FILLER_58_748 ();
 sg13g2_fill_1 FILLER_58_768 ();
 sg13g2_decap_4 FILLER_58_788 ();
 sg13g2_fill_2 FILLER_58_802 ();
 sg13g2_decap_8 FILLER_58_830 ();
 sg13g2_fill_1 FILLER_58_837 ();
 sg13g2_fill_2 FILLER_58_872 ();
 sg13g2_fill_1 FILLER_58_874 ();
 sg13g2_fill_1 FILLER_58_906 ();
 sg13g2_fill_2 FILLER_58_919 ();
 sg13g2_fill_2 FILLER_58_934 ();
 sg13g2_fill_1 FILLER_58_936 ();
 sg13g2_fill_2 FILLER_58_1018 ();
 sg13g2_fill_1 FILLER_58_1080 ();
 sg13g2_fill_2 FILLER_58_1094 ();
 sg13g2_decap_4 FILLER_58_1121 ();
 sg13g2_fill_2 FILLER_58_1138 ();
 sg13g2_fill_2 FILLER_58_1145 ();
 sg13g2_fill_2 FILLER_58_1157 ();
 sg13g2_fill_1 FILLER_58_1163 ();
 sg13g2_decap_4 FILLER_58_1177 ();
 sg13g2_fill_1 FILLER_58_1181 ();
 sg13g2_decap_4 FILLER_58_1297 ();
 sg13g2_fill_1 FILLER_58_1301 ();
 sg13g2_fill_1 FILLER_58_1456 ();
 sg13g2_fill_2 FILLER_58_1466 ();
 sg13g2_fill_1 FILLER_58_1468 ();
 sg13g2_fill_1 FILLER_58_1483 ();
 sg13g2_fill_2 FILLER_58_1500 ();
 sg13g2_fill_1 FILLER_58_1502 ();
 sg13g2_decap_8 FILLER_58_1509 ();
 sg13g2_fill_1 FILLER_58_1591 ();
 sg13g2_fill_2 FILLER_58_1611 ();
 sg13g2_fill_1 FILLER_58_1649 ();
 sg13g2_fill_2 FILLER_58_1702 ();
 sg13g2_fill_2 FILLER_58_1735 ();
 sg13g2_fill_1 FILLER_58_1767 ();
 sg13g2_fill_1 FILLER_59_26 ();
 sg13g2_fill_2 FILLER_59_126 ();
 sg13g2_fill_1 FILLER_59_174 ();
 sg13g2_fill_2 FILLER_59_211 ();
 sg13g2_fill_2 FILLER_59_239 ();
 sg13g2_fill_1 FILLER_59_241 ();
 sg13g2_fill_1 FILLER_59_269 ();
 sg13g2_fill_1 FILLER_59_279 ();
 sg13g2_fill_1 FILLER_59_301 ();
 sg13g2_fill_1 FILLER_59_352 ();
 sg13g2_fill_2 FILLER_59_387 ();
 sg13g2_decap_4 FILLER_59_460 ();
 sg13g2_fill_1 FILLER_59_503 ();
 sg13g2_fill_2 FILLER_59_552 ();
 sg13g2_fill_1 FILLER_59_554 ();
 sg13g2_decap_8 FILLER_59_559 ();
 sg13g2_fill_1 FILLER_59_566 ();
 sg13g2_fill_1 FILLER_59_593 ();
 sg13g2_fill_1 FILLER_59_603 ();
 sg13g2_fill_1 FILLER_59_612 ();
 sg13g2_fill_2 FILLER_59_632 ();
 sg13g2_decap_4 FILLER_59_642 ();
 sg13g2_fill_1 FILLER_59_646 ();
 sg13g2_decap_4 FILLER_59_651 ();
 sg13g2_fill_2 FILLER_59_655 ();
 sg13g2_decap_8 FILLER_59_665 ();
 sg13g2_fill_2 FILLER_59_672 ();
 sg13g2_fill_1 FILLER_59_674 ();
 sg13g2_decap_8 FILLER_59_695 ();
 sg13g2_fill_2 FILLER_59_702 ();
 sg13g2_decap_4 FILLER_59_738 ();
 sg13g2_fill_1 FILLER_59_777 ();
 sg13g2_decap_8 FILLER_59_823 ();
 sg13g2_fill_2 FILLER_59_858 ();
 sg13g2_fill_1 FILLER_59_860 ();
 sg13g2_decap_4 FILLER_59_880 ();
 sg13g2_fill_1 FILLER_59_892 ();
 sg13g2_decap_4 FILLER_59_921 ();
 sg13g2_fill_1 FILLER_59_925 ();
 sg13g2_fill_2 FILLER_59_962 ();
 sg13g2_fill_1 FILLER_59_964 ();
 sg13g2_fill_1 FILLER_59_969 ();
 sg13g2_fill_2 FILLER_59_988 ();
 sg13g2_fill_2 FILLER_59_1038 ();
 sg13g2_fill_1 FILLER_59_1049 ();
 sg13g2_decap_4 FILLER_59_1125 ();
 sg13g2_fill_1 FILLER_59_1129 ();
 sg13g2_decap_4 FILLER_59_1138 ();
 sg13g2_fill_1 FILLER_59_1196 ();
 sg13g2_fill_2 FILLER_59_1263 ();
 sg13g2_fill_1 FILLER_59_1293 ();
 sg13g2_fill_2 FILLER_59_1347 ();
 sg13g2_fill_1 FILLER_59_1349 ();
 sg13g2_fill_2 FILLER_59_1396 ();
 sg13g2_decap_8 FILLER_59_1480 ();
 sg13g2_fill_1 FILLER_59_1487 ();
 sg13g2_fill_2 FILLER_59_1514 ();
 sg13g2_fill_2 FILLER_59_1524 ();
 sg13g2_fill_2 FILLER_59_1536 ();
 sg13g2_fill_1 FILLER_59_1538 ();
 sg13g2_fill_2 FILLER_59_1543 ();
 sg13g2_fill_1 FILLER_59_1570 ();
 sg13g2_fill_2 FILLER_59_1589 ();
 sg13g2_fill_1 FILLER_59_1591 ();
 sg13g2_fill_2 FILLER_59_1633 ();
 sg13g2_fill_1 FILLER_59_1635 ();
 sg13g2_decap_8 FILLER_59_1648 ();
 sg13g2_fill_1 FILLER_59_1655 ();
 sg13g2_fill_2 FILLER_59_1696 ();
 sg13g2_fill_1 FILLER_59_1698 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_2 ();
 sg13g2_fill_2 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_9 ();
 sg13g2_fill_2 FILLER_60_46 ();
 sg13g2_fill_1 FILLER_60_48 ();
 sg13g2_fill_1 FILLER_60_68 ();
 sg13g2_fill_2 FILLER_60_87 ();
 sg13g2_fill_1 FILLER_60_108 ();
 sg13g2_fill_2 FILLER_60_138 ();
 sg13g2_fill_1 FILLER_60_140 ();
 sg13g2_fill_2 FILLER_60_256 ();
 sg13g2_fill_1 FILLER_60_335 ();
 sg13g2_fill_1 FILLER_60_346 ();
 sg13g2_fill_2 FILLER_60_368 ();
 sg13g2_fill_1 FILLER_60_386 ();
 sg13g2_fill_2 FILLER_60_430 ();
 sg13g2_fill_1 FILLER_60_432 ();
 sg13g2_fill_2 FILLER_60_443 ();
 sg13g2_fill_2 FILLER_60_488 ();
 sg13g2_fill_1 FILLER_60_524 ();
 sg13g2_decap_8 FILLER_60_555 ();
 sg13g2_fill_2 FILLER_60_570 ();
 sg13g2_fill_1 FILLER_60_576 ();
 sg13g2_fill_2 FILLER_60_581 ();
 sg13g2_fill_1 FILLER_60_583 ();
 sg13g2_fill_2 FILLER_60_610 ();
 sg13g2_fill_1 FILLER_60_612 ();
 sg13g2_fill_2 FILLER_60_628 ();
 sg13g2_fill_1 FILLER_60_635 ();
 sg13g2_decap_4 FILLER_60_647 ();
 sg13g2_fill_1 FILLER_60_651 ();
 sg13g2_fill_1 FILLER_60_656 ();
 sg13g2_fill_2 FILLER_60_673 ();
 sg13g2_fill_1 FILLER_60_701 ();
 sg13g2_fill_2 FILLER_60_756 ();
 sg13g2_fill_1 FILLER_60_758 ();
 sg13g2_fill_2 FILLER_60_805 ();
 sg13g2_decap_4 FILLER_60_812 ();
 sg13g2_decap_4 FILLER_60_822 ();
 sg13g2_fill_1 FILLER_60_826 ();
 sg13g2_fill_2 FILLER_60_863 ();
 sg13g2_fill_1 FILLER_60_865 ();
 sg13g2_decap_8 FILLER_60_892 ();
 sg13g2_fill_2 FILLER_60_977 ();
 sg13g2_fill_1 FILLER_60_979 ();
 sg13g2_fill_2 FILLER_60_1020 ();
 sg13g2_decap_8 FILLER_60_1071 ();
 sg13g2_fill_1 FILLER_60_1078 ();
 sg13g2_fill_1 FILLER_60_1092 ();
 sg13g2_fill_2 FILLER_60_1120 ();
 sg13g2_fill_2 FILLER_60_1153 ();
 sg13g2_decap_4 FILLER_60_1207 ();
 sg13g2_fill_2 FILLER_60_1211 ();
 sg13g2_fill_2 FILLER_60_1223 ();
 sg13g2_decap_8 FILLER_60_1244 ();
 sg13g2_fill_2 FILLER_60_1251 ();
 sg13g2_fill_1 FILLER_60_1292 ();
 sg13g2_fill_2 FILLER_60_1299 ();
 sg13g2_fill_1 FILLER_60_1301 ();
 sg13g2_decap_4 FILLER_60_1312 ();
 sg13g2_fill_1 FILLER_60_1316 ();
 sg13g2_decap_4 FILLER_60_1408 ();
 sg13g2_fill_2 FILLER_60_1421 ();
 sg13g2_fill_1 FILLER_60_1423 ();
 sg13g2_fill_2 FILLER_60_1450 ();
 sg13g2_fill_2 FILLER_60_1469 ();
 sg13g2_decap_4 FILLER_60_1484 ();
 sg13g2_fill_1 FILLER_60_1488 ();
 sg13g2_fill_1 FILLER_60_1498 ();
 sg13g2_fill_2 FILLER_60_1503 ();
 sg13g2_decap_4 FILLER_60_1509 ();
 sg13g2_fill_1 FILLER_60_1513 ();
 sg13g2_fill_1 FILLER_60_1573 ();
 sg13g2_fill_1 FILLER_60_1600 ();
 sg13g2_decap_4 FILLER_60_1637 ();
 sg13g2_fill_2 FILLER_60_1654 ();
 sg13g2_fill_1 FILLER_60_1656 ();
 sg13g2_decap_8 FILLER_60_1666 ();
 sg13g2_decap_8 FILLER_60_1673 ();
 sg13g2_decap_4 FILLER_60_1685 ();
 sg13g2_fill_1 FILLER_60_1720 ();
 sg13g2_fill_1 FILLER_60_1767 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_87 ();
 sg13g2_fill_1 FILLER_61_89 ();
 sg13g2_fill_2 FILLER_61_116 ();
 sg13g2_fill_1 FILLER_61_118 ();
 sg13g2_fill_2 FILLER_61_145 ();
 sg13g2_fill_1 FILLER_61_147 ();
 sg13g2_fill_1 FILLER_61_175 ();
 sg13g2_fill_1 FILLER_61_198 ();
 sg13g2_fill_1 FILLER_61_209 ();
 sg13g2_fill_2 FILLER_61_248 ();
 sg13g2_fill_1 FILLER_61_266 ();
 sg13g2_fill_1 FILLER_61_286 ();
 sg13g2_fill_2 FILLER_61_308 ();
 sg13g2_fill_2 FILLER_61_336 ();
 sg13g2_fill_1 FILLER_61_338 ();
 sg13g2_decap_4 FILLER_61_378 ();
 sg13g2_fill_1 FILLER_61_382 ();
 sg13g2_fill_2 FILLER_61_397 ();
 sg13g2_fill_1 FILLER_61_399 ();
 sg13g2_fill_1 FILLER_61_433 ();
 sg13g2_fill_2 FILLER_61_439 ();
 sg13g2_fill_1 FILLER_61_441 ();
 sg13g2_fill_2 FILLER_61_486 ();
 sg13g2_fill_1 FILLER_61_493 ();
 sg13g2_fill_2 FILLER_61_499 ();
 sg13g2_fill_2 FILLER_61_539 ();
 sg13g2_fill_2 FILLER_61_567 ();
 sg13g2_fill_1 FILLER_61_569 ();
 sg13g2_fill_1 FILLER_61_589 ();
 sg13g2_fill_1 FILLER_61_609 ();
 sg13g2_decap_8 FILLER_61_672 ();
 sg13g2_fill_2 FILLER_61_705 ();
 sg13g2_fill_2 FILLER_61_715 ();
 sg13g2_fill_2 FILLER_61_720 ();
 sg13g2_fill_2 FILLER_61_730 ();
 sg13g2_fill_1 FILLER_61_736 ();
 sg13g2_fill_2 FILLER_61_804 ();
 sg13g2_fill_1 FILLER_61_806 ();
 sg13g2_fill_2 FILLER_61_811 ();
 sg13g2_fill_1 FILLER_61_835 ();
 sg13g2_fill_2 FILLER_61_885 ();
 sg13g2_fill_2 FILLER_61_897 ();
 sg13g2_fill_1 FILLER_61_908 ();
 sg13g2_decap_4 FILLER_61_919 ();
 sg13g2_fill_1 FILLER_61_923 ();
 sg13g2_fill_2 FILLER_61_989 ();
 sg13g2_fill_1 FILLER_61_991 ();
 sg13g2_fill_1 FILLER_61_1028 ();
 sg13g2_fill_2 FILLER_61_1037 ();
 sg13g2_decap_4 FILLER_61_1072 ();
 sg13g2_decap_8 FILLER_61_1125 ();
 sg13g2_fill_1 FILLER_61_1132 ();
 sg13g2_decap_8 FILLER_61_1137 ();
 sg13g2_fill_1 FILLER_61_1178 ();
 sg13g2_fill_2 FILLER_61_1188 ();
 sg13g2_fill_1 FILLER_61_1190 ();
 sg13g2_fill_1 FILLER_61_1241 ();
 sg13g2_fill_2 FILLER_61_1268 ();
 sg13g2_decap_8 FILLER_61_1322 ();
 sg13g2_decap_4 FILLER_61_1329 ();
 sg13g2_fill_1 FILLER_61_1364 ();
 sg13g2_fill_2 FILLER_61_1378 ();
 sg13g2_fill_1 FILLER_61_1380 ();
 sg13g2_fill_2 FILLER_61_1394 ();
 sg13g2_decap_8 FILLER_61_1425 ();
 sg13g2_fill_2 FILLER_61_1432 ();
 sg13g2_fill_2 FILLER_61_1448 ();
 sg13g2_decap_8 FILLER_61_1486 ();
 sg13g2_fill_2 FILLER_61_1493 ();
 sg13g2_fill_2 FILLER_61_1521 ();
 sg13g2_fill_1 FILLER_61_1523 ();
 sg13g2_fill_1 FILLER_61_1550 ();
 sg13g2_fill_2 FILLER_61_1561 ();
 sg13g2_fill_1 FILLER_61_1563 ();
 sg13g2_fill_1 FILLER_61_1569 ();
 sg13g2_fill_2 FILLER_61_1583 ();
 sg13g2_fill_2 FILLER_61_1597 ();
 sg13g2_fill_1 FILLER_61_1599 ();
 sg13g2_decap_4 FILLER_61_1612 ();
 sg13g2_fill_1 FILLER_61_1616 ();
 sg13g2_fill_1 FILLER_61_1634 ();
 sg13g2_fill_2 FILLER_61_1680 ();
 sg13g2_fill_2 FILLER_61_1696 ();
 sg13g2_fill_1 FILLER_61_1734 ();
 sg13g2_fill_2 FILLER_61_1765 ();
 sg13g2_fill_1 FILLER_61_1767 ();
 sg13g2_fill_2 FILLER_62_40 ();
 sg13g2_fill_1 FILLER_62_42 ();
 sg13g2_fill_2 FILLER_62_132 ();
 sg13g2_fill_1 FILLER_62_134 ();
 sg13g2_fill_2 FILLER_62_145 ();
 sg13g2_fill_2 FILLER_62_155 ();
 sg13g2_fill_1 FILLER_62_157 ();
 sg13g2_fill_1 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_214 ();
 sg13g2_fill_1 FILLER_62_255 ();
 sg13g2_fill_1 FILLER_62_309 ();
 sg13g2_decap_8 FILLER_62_336 ();
 sg13g2_decap_4 FILLER_62_343 ();
 sg13g2_fill_2 FILLER_62_347 ();
 sg13g2_fill_2 FILLER_62_358 ();
 sg13g2_fill_2 FILLER_62_457 ();
 sg13g2_fill_1 FILLER_62_459 ();
 sg13g2_fill_1 FILLER_62_480 ();
 sg13g2_fill_2 FILLER_62_515 ();
 sg13g2_fill_2 FILLER_62_549 ();
 sg13g2_fill_1 FILLER_62_551 ();
 sg13g2_fill_2 FILLER_62_560 ();
 sg13g2_decap_4 FILLER_62_571 ();
 sg13g2_decap_4 FILLER_62_584 ();
 sg13g2_fill_2 FILLER_62_588 ();
 sg13g2_fill_2 FILLER_62_594 ();
 sg13g2_fill_2 FILLER_62_611 ();
 sg13g2_decap_4 FILLER_62_630 ();
 sg13g2_decap_4 FILLER_62_650 ();
 sg13g2_fill_2 FILLER_62_654 ();
 sg13g2_fill_2 FILLER_62_666 ();
 sg13g2_fill_2 FILLER_62_704 ();
 sg13g2_fill_1 FILLER_62_716 ();
 sg13g2_fill_2 FILLER_62_723 ();
 sg13g2_fill_2 FILLER_62_744 ();
 sg13g2_fill_1 FILLER_62_746 ();
 sg13g2_fill_1 FILLER_62_765 ();
 sg13g2_fill_1 FILLER_62_849 ();
 sg13g2_fill_2 FILLER_62_921 ();
 sg13g2_fill_1 FILLER_62_923 ();
 sg13g2_fill_1 FILLER_62_1005 ();
 sg13g2_fill_1 FILLER_62_1011 ();
 sg13g2_fill_1 FILLER_62_1021 ();
 sg13g2_fill_2 FILLER_62_1042 ();
 sg13g2_fill_1 FILLER_62_1044 ();
 sg13g2_decap_4 FILLER_62_1126 ();
 sg13g2_fill_1 FILLER_62_1155 ();
 sg13g2_fill_2 FILLER_62_1211 ();
 sg13g2_fill_2 FILLER_62_1251 ();
 sg13g2_fill_2 FILLER_62_1257 ();
 sg13g2_fill_1 FILLER_62_1259 ();
 sg13g2_decap_8 FILLER_62_1266 ();
 sg13g2_decap_8 FILLER_62_1273 ();
 sg13g2_fill_1 FILLER_62_1299 ();
 sg13g2_fill_2 FILLER_62_1314 ();
 sg13g2_fill_1 FILLER_62_1360 ();
 sg13g2_decap_4 FILLER_62_1379 ();
 sg13g2_fill_1 FILLER_62_1387 ();
 sg13g2_fill_2 FILLER_62_1410 ();
 sg13g2_fill_1 FILLER_62_1461 ();
 sg13g2_decap_4 FILLER_62_1488 ();
 sg13g2_fill_2 FILLER_62_1496 ();
 sg13g2_fill_1 FILLER_62_1498 ();
 sg13g2_fill_1 FILLER_62_1525 ();
 sg13g2_fill_2 FILLER_62_1603 ();
 sg13g2_fill_1 FILLER_62_1605 ();
 sg13g2_fill_1 FILLER_62_1614 ();
 sg13g2_fill_2 FILLER_62_1673 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_59 ();
 sg13g2_fill_2 FILLER_63_78 ();
 sg13g2_fill_1 FILLER_63_116 ();
 sg13g2_fill_2 FILLER_63_194 ();
 sg13g2_fill_2 FILLER_63_209 ();
 sg13g2_fill_2 FILLER_63_296 ();
 sg13g2_fill_1 FILLER_63_298 ();
 sg13g2_fill_2 FILLER_63_323 ();
 sg13g2_decap_4 FILLER_63_333 ();
 sg13g2_decap_4 FILLER_63_345 ();
 sg13g2_fill_2 FILLER_63_349 ();
 sg13g2_fill_2 FILLER_63_400 ();
 sg13g2_fill_1 FILLER_63_402 ();
 sg13g2_fill_2 FILLER_63_432 ();
 sg13g2_fill_1 FILLER_63_434 ();
 sg13g2_fill_1 FILLER_63_525 ();
 sg13g2_fill_1 FILLER_63_552 ();
 sg13g2_decap_4 FILLER_63_569 ();
 sg13g2_fill_1 FILLER_63_634 ();
 sg13g2_decap_8 FILLER_63_639 ();
 sg13g2_decap_8 FILLER_63_646 ();
 sg13g2_decap_4 FILLER_63_653 ();
 sg13g2_fill_1 FILLER_63_657 ();
 sg13g2_fill_2 FILLER_63_684 ();
 sg13g2_fill_2 FILLER_63_699 ();
 sg13g2_fill_1 FILLER_63_764 ();
 sg13g2_fill_2 FILLER_63_791 ();
 sg13g2_fill_2 FILLER_63_807 ();
 sg13g2_fill_1 FILLER_63_809 ();
 sg13g2_fill_2 FILLER_63_828 ();
 sg13g2_fill_1 FILLER_63_830 ();
 sg13g2_fill_1 FILLER_63_886 ();
 sg13g2_fill_2 FILLER_63_891 ();
 sg13g2_fill_1 FILLER_63_893 ();
 sg13g2_fill_2 FILLER_63_903 ();
 sg13g2_fill_1 FILLER_63_905 ();
 sg13g2_decap_8 FILLER_63_910 ();
 sg13g2_decap_4 FILLER_63_917 ();
 sg13g2_fill_1 FILLER_63_921 ();
 sg13g2_fill_2 FILLER_63_1129 ();
 sg13g2_fill_2 FILLER_63_1170 ();
 sg13g2_decap_4 FILLER_63_1267 ();
 sg13g2_fill_2 FILLER_63_1271 ();
 sg13g2_fill_1 FILLER_63_1277 ();
 sg13g2_fill_1 FILLER_63_1344 ();
 sg13g2_fill_2 FILLER_63_1430 ();
 sg13g2_fill_2 FILLER_63_1451 ();
 sg13g2_fill_2 FILLER_63_1482 ();
 sg13g2_fill_1 FILLER_63_1484 ();
 sg13g2_fill_2 FILLER_63_1494 ();
 sg13g2_fill_1 FILLER_63_1496 ();
 sg13g2_fill_2 FILLER_63_1507 ();
 sg13g2_fill_1 FILLER_63_1622 ();
 sg13g2_fill_1 FILLER_63_1647 ();
 sg13g2_fill_1 FILLER_63_1701 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_61 ();
 sg13g2_fill_2 FILLER_64_88 ();
 sg13g2_fill_2 FILLER_64_109 ();
 sg13g2_fill_1 FILLER_64_111 ();
 sg13g2_fill_2 FILLER_64_135 ();
 sg13g2_fill_2 FILLER_64_158 ();
 sg13g2_fill_1 FILLER_64_160 ();
 sg13g2_fill_2 FILLER_64_189 ();
 sg13g2_fill_1 FILLER_64_191 ();
 sg13g2_fill_1 FILLER_64_218 ();
 sg13g2_decap_4 FILLER_64_253 ();
 sg13g2_fill_1 FILLER_64_257 ();
 sg13g2_decap_4 FILLER_64_297 ();
 sg13g2_fill_1 FILLER_64_301 ();
 sg13g2_fill_2 FILLER_64_316 ();
 sg13g2_fill_1 FILLER_64_318 ();
 sg13g2_fill_1 FILLER_64_327 ();
 sg13g2_fill_2 FILLER_64_340 ();
 sg13g2_fill_2 FILLER_64_354 ();
 sg13g2_fill_2 FILLER_64_405 ();
 sg13g2_fill_2 FILLER_64_468 ();
 sg13g2_fill_1 FILLER_64_470 ();
 sg13g2_fill_2 FILLER_64_481 ();
 sg13g2_decap_8 FILLER_64_526 ();
 sg13g2_fill_2 FILLER_64_538 ();
 sg13g2_decap_8 FILLER_64_563 ();
 sg13g2_decap_4 FILLER_64_570 ();
 sg13g2_fill_1 FILLER_64_574 ();
 sg13g2_fill_1 FILLER_64_590 ();
 sg13g2_fill_2 FILLER_64_654 ();
 sg13g2_fill_1 FILLER_64_656 ();
 sg13g2_fill_1 FILLER_64_667 ();
 sg13g2_fill_2 FILLER_64_735 ();
 sg13g2_fill_1 FILLER_64_737 ();
 sg13g2_fill_2 FILLER_64_757 ();
 sg13g2_fill_2 FILLER_64_801 ();
 sg13g2_fill_1 FILLER_64_803 ();
 sg13g2_fill_1 FILLER_64_835 ();
 sg13g2_fill_1 FILLER_64_872 ();
 sg13g2_decap_8 FILLER_64_899 ();
 sg13g2_decap_8 FILLER_64_906 ();
 sg13g2_fill_1 FILLER_64_913 ();
 sg13g2_fill_2 FILLER_64_997 ();
 sg13g2_fill_2 FILLER_64_1054 ();
 sg13g2_fill_2 FILLER_64_1075 ();
 sg13g2_decap_4 FILLER_64_1122 ();
 sg13g2_fill_1 FILLER_64_1141 ();
 sg13g2_fill_2 FILLER_64_1151 ();
 sg13g2_fill_1 FILLER_64_1153 ();
 sg13g2_fill_2 FILLER_64_1229 ();
 sg13g2_fill_2 FILLER_64_1250 ();
 sg13g2_fill_2 FILLER_64_1275 ();
 sg13g2_fill_1 FILLER_64_1300 ();
 sg13g2_fill_1 FILLER_64_1320 ();
 sg13g2_fill_1 FILLER_64_1384 ();
 sg13g2_fill_2 FILLER_64_1466 ();
 sg13g2_fill_1 FILLER_64_1526 ();
 sg13g2_fill_2 FILLER_64_1537 ();
 sg13g2_fill_1 FILLER_64_1539 ();
 sg13g2_fill_2 FILLER_64_1576 ();
 sg13g2_fill_1 FILLER_64_1578 ();
 sg13g2_fill_2 FILLER_64_1584 ();
 sg13g2_fill_1 FILLER_64_1629 ();
 sg13g2_fill_2 FILLER_64_1743 ();
 sg13g2_fill_1 FILLER_64_1767 ();
 sg13g2_fill_2 FILLER_65_70 ();
 sg13g2_fill_1 FILLER_65_92 ();
 sg13g2_fill_2 FILLER_65_142 ();
 sg13g2_fill_1 FILLER_65_170 ();
 sg13g2_fill_2 FILLER_65_211 ();
 sg13g2_fill_1 FILLER_65_246 ();
 sg13g2_fill_1 FILLER_65_303 ();
 sg13g2_fill_2 FILLER_65_423 ();
 sg13g2_fill_2 FILLER_65_448 ();
 sg13g2_decap_4 FILLER_65_486 ();
 sg13g2_fill_1 FILLER_65_526 ();
 sg13g2_fill_2 FILLER_65_540 ();
 sg13g2_fill_1 FILLER_65_550 ();
 sg13g2_fill_2 FILLER_65_567 ();
 sg13g2_fill_1 FILLER_65_569 ();
 sg13g2_fill_2 FILLER_65_662 ();
 sg13g2_decap_4 FILLER_65_690 ();
 sg13g2_fill_1 FILLER_65_694 ();
 sg13g2_fill_1 FILLER_65_714 ();
 sg13g2_fill_1 FILLER_65_761 ();
 sg13g2_fill_1 FILLER_65_785 ();
 sg13g2_fill_2 FILLER_65_817 ();
 sg13g2_fill_2 FILLER_65_824 ();
 sg13g2_decap_4 FILLER_65_894 ();
 sg13g2_fill_2 FILLER_65_956 ();
 sg13g2_fill_2 FILLER_65_1016 ();
 sg13g2_fill_2 FILLER_65_1119 ();
 sg13g2_fill_1 FILLER_65_1121 ();
 sg13g2_fill_1 FILLER_65_1173 ();
 sg13g2_fill_1 FILLER_65_1191 ();
 sg13g2_fill_1 FILLER_65_1201 ();
 sg13g2_fill_1 FILLER_65_1408 ();
 sg13g2_fill_2 FILLER_65_1445 ();
 sg13g2_fill_1 FILLER_65_1447 ();
 sg13g2_fill_2 FILLER_65_1515 ();
 sg13g2_fill_1 FILLER_65_1517 ();
 sg13g2_fill_2 FILLER_65_1566 ();
 sg13g2_fill_2 FILLER_65_1589 ();
 sg13g2_fill_1 FILLER_65_1591 ();
 sg13g2_fill_2 FILLER_65_1602 ();
 sg13g2_fill_1 FILLER_65_1604 ();
 sg13g2_fill_1 FILLER_65_1638 ();
 sg13g2_fill_2 FILLER_65_1653 ();
 sg13g2_fill_1 FILLER_65_1683 ();
 sg13g2_fill_1 FILLER_65_1698 ();
 sg13g2_fill_1 FILLER_65_1716 ();
 sg13g2_fill_1 FILLER_65_1736 ();
 sg13g2_fill_1 FILLER_65_1767 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_28 ();
 sg13g2_fill_2 FILLER_66_60 ();
 sg13g2_fill_1 FILLER_66_62 ();
 sg13g2_fill_2 FILLER_66_89 ();
 sg13g2_fill_1 FILLER_66_91 ();
 sg13g2_fill_2 FILLER_66_153 ();
 sg13g2_fill_2 FILLER_66_200 ();
 sg13g2_fill_1 FILLER_66_202 ();
 sg13g2_fill_1 FILLER_66_235 ();
 sg13g2_fill_2 FILLER_66_244 ();
 sg13g2_fill_1 FILLER_66_261 ();
 sg13g2_fill_2 FILLER_66_324 ();
 sg13g2_fill_1 FILLER_66_326 ();
 sg13g2_decap_4 FILLER_66_365 ();
 sg13g2_fill_1 FILLER_66_377 ();
 sg13g2_fill_2 FILLER_66_410 ();
 sg13g2_fill_1 FILLER_66_412 ();
 sg13g2_fill_1 FILLER_66_441 ();
 sg13g2_fill_1 FILLER_66_454 ();
 sg13g2_fill_2 FILLER_66_470 ();
 sg13g2_fill_2 FILLER_66_486 ();
 sg13g2_fill_1 FILLER_66_488 ();
 sg13g2_fill_2 FILLER_66_518 ();
 sg13g2_fill_2 FILLER_66_525 ();
 sg13g2_fill_2 FILLER_66_550 ();
 sg13g2_decap_8 FILLER_66_561 ();
 sg13g2_decap_8 FILLER_66_568 ();
 sg13g2_fill_1 FILLER_66_575 ();
 sg13g2_fill_1 FILLER_66_600 ();
 sg13g2_fill_2 FILLER_66_643 ();
 sg13g2_fill_1 FILLER_66_645 ();
 sg13g2_fill_2 FILLER_66_682 ();
 sg13g2_fill_1 FILLER_66_684 ();
 sg13g2_fill_1 FILLER_66_749 ();
 sg13g2_fill_2 FILLER_66_772 ();
 sg13g2_fill_1 FILLER_66_774 ();
 sg13g2_fill_1 FILLER_66_783 ();
 sg13g2_fill_2 FILLER_66_809 ();
 sg13g2_fill_1 FILLER_66_811 ();
 sg13g2_fill_2 FILLER_66_842 ();
 sg13g2_fill_2 FILLER_66_875 ();
 sg13g2_fill_1 FILLER_66_877 ();
 sg13g2_decap_8 FILLER_66_890 ();
 sg13g2_decap_8 FILLER_66_897 ();
 sg13g2_fill_2 FILLER_66_904 ();
 sg13g2_fill_1 FILLER_66_906 ();
 sg13g2_fill_1 FILLER_66_1009 ();
 sg13g2_fill_1 FILLER_66_1030 ();
 sg13g2_fill_2 FILLER_66_1208 ();
 sg13g2_fill_2 FILLER_66_1219 ();
 sg13g2_fill_2 FILLER_66_1241 ();
 sg13g2_fill_1 FILLER_66_1246 ();
 sg13g2_fill_2 FILLER_66_1256 ();
 sg13g2_fill_1 FILLER_66_1303 ();
 sg13g2_fill_2 FILLER_66_1338 ();
 sg13g2_fill_1 FILLER_66_1340 ();
 sg13g2_fill_2 FILLER_66_1360 ();
 sg13g2_fill_2 FILLER_66_1377 ();
 sg13g2_fill_2 FILLER_66_1408 ();
 sg13g2_fill_2 FILLER_66_1419 ();
 sg13g2_fill_1 FILLER_66_1443 ();
 sg13g2_fill_2 FILLER_66_1471 ();
 sg13g2_decap_8 FILLER_66_1478 ();
 sg13g2_fill_2 FILLER_66_1485 ();
 sg13g2_fill_1 FILLER_66_1487 ();
 sg13g2_decap_4 FILLER_66_1492 ();
 sg13g2_fill_2 FILLER_66_1496 ();
 sg13g2_decap_4 FILLER_66_1503 ();
 sg13g2_fill_2 FILLER_66_1516 ();
 sg13g2_decap_4 FILLER_66_1534 ();
 sg13g2_fill_2 FILLER_66_1538 ();
 sg13g2_decap_4 FILLER_66_1555 ();
 sg13g2_fill_1 FILLER_66_1559 ();
 sg13g2_fill_2 FILLER_66_1596 ();
 sg13g2_fill_2 FILLER_66_1737 ();
 sg13g2_fill_2 FILLER_66_1765 ();
 sg13g2_fill_1 FILLER_66_1767 ();
 sg13g2_fill_2 FILLER_67_4 ();
 sg13g2_fill_1 FILLER_67_6 ();
 sg13g2_fill_1 FILLER_67_56 ();
 sg13g2_fill_1 FILLER_67_67 ();
 sg13g2_fill_2 FILLER_67_129 ();
 sg13g2_fill_1 FILLER_67_201 ();
 sg13g2_fill_2 FILLER_67_210 ();
 sg13g2_fill_1 FILLER_67_212 ();
 sg13g2_fill_2 FILLER_67_222 ();
 sg13g2_fill_1 FILLER_67_224 ();
 sg13g2_fill_1 FILLER_67_287 ();
 sg13g2_fill_1 FILLER_67_297 ();
 sg13g2_fill_1 FILLER_67_318 ();
 sg13g2_fill_2 FILLER_67_352 ();
 sg13g2_fill_1 FILLER_67_354 ();
 sg13g2_fill_1 FILLER_67_400 ();
 sg13g2_fill_2 FILLER_67_433 ();
 sg13g2_fill_1 FILLER_67_435 ();
 sg13g2_fill_2 FILLER_67_485 ();
 sg13g2_fill_2 FILLER_67_527 ();
 sg13g2_fill_1 FILLER_67_529 ();
 sg13g2_fill_2 FILLER_67_557 ();
 sg13g2_fill_1 FILLER_67_565 ();
 sg13g2_fill_2 FILLER_67_605 ();
 sg13g2_fill_1 FILLER_67_607 ();
 sg13g2_fill_1 FILLER_67_616 ();
 sg13g2_fill_1 FILLER_67_743 ();
 sg13g2_fill_1 FILLER_67_784 ();
 sg13g2_fill_2 FILLER_67_826 ();
 sg13g2_fill_1 FILLER_67_828 ();
 sg13g2_fill_1 FILLER_67_883 ();
 sg13g2_fill_1 FILLER_67_924 ();
 sg13g2_fill_2 FILLER_67_934 ();
 sg13g2_fill_2 FILLER_67_1011 ();
 sg13g2_fill_2 FILLER_67_1029 ();
 sg13g2_fill_1 FILLER_67_1046 ();
 sg13g2_fill_1 FILLER_67_1059 ();
 sg13g2_fill_2 FILLER_67_1094 ();
 sg13g2_fill_1 FILLER_67_1118 ();
 sg13g2_fill_1 FILLER_67_1213 ();
 sg13g2_fill_2 FILLER_67_1233 ();
 sg13g2_fill_2 FILLER_67_1249 ();
 sg13g2_fill_1 FILLER_67_1251 ();
 sg13g2_fill_1 FILLER_67_1260 ();
 sg13g2_decap_4 FILLER_67_1295 ();
 sg13g2_fill_1 FILLER_67_1299 ();
 sg13g2_fill_1 FILLER_67_1357 ();
 sg13g2_fill_2 FILLER_67_1394 ();
 sg13g2_fill_1 FILLER_67_1396 ();
 sg13g2_fill_2 FILLER_67_1428 ();
 sg13g2_fill_1 FILLER_67_1430 ();
 sg13g2_fill_2 FILLER_67_1440 ();
 sg13g2_fill_1 FILLER_67_1442 ();
 sg13g2_fill_1 FILLER_67_1453 ();
 sg13g2_fill_1 FILLER_67_1490 ();
 sg13g2_fill_1 FILLER_67_1536 ();
 sg13g2_fill_2 FILLER_67_1573 ();
 sg13g2_fill_1 FILLER_67_1575 ();
 sg13g2_fill_2 FILLER_67_1602 ();
 sg13g2_fill_1 FILLER_67_1627 ();
 sg13g2_fill_2 FILLER_67_1704 ();
 sg13g2_fill_1 FILLER_67_1706 ();
 sg13g2_fill_2 FILLER_67_1740 ();
 sg13g2_fill_1 FILLER_68_76 ();
 sg13g2_fill_1 FILLER_68_147 ();
 sg13g2_fill_1 FILLER_68_184 ();
 sg13g2_fill_1 FILLER_68_203 ();
 sg13g2_fill_1 FILLER_68_212 ();
 sg13g2_fill_1 FILLER_68_249 ();
 sg13g2_fill_1 FILLER_68_258 ();
 sg13g2_fill_1 FILLER_68_268 ();
 sg13g2_fill_1 FILLER_68_279 ();
 sg13g2_fill_1 FILLER_68_329 ();
 sg13g2_fill_1 FILLER_68_389 ();
 sg13g2_fill_2 FILLER_68_405 ();
 sg13g2_fill_1 FILLER_68_407 ();
 sg13g2_fill_1 FILLER_68_500 ();
 sg13g2_fill_1 FILLER_68_527 ();
 sg13g2_decap_8 FILLER_68_565 ();
 sg13g2_fill_1 FILLER_68_572 ();
 sg13g2_fill_2 FILLER_68_587 ();
 sg13g2_fill_2 FILLER_68_604 ();
 sg13g2_fill_1 FILLER_68_615 ();
 sg13g2_fill_2 FILLER_68_657 ();
 sg13g2_fill_1 FILLER_68_659 ();
 sg13g2_fill_2 FILLER_68_669 ();
 sg13g2_fill_2 FILLER_68_675 ();
 sg13g2_fill_1 FILLER_68_749 ();
 sg13g2_fill_2 FILLER_68_795 ();
 sg13g2_fill_1 FILLER_68_797 ();
 sg13g2_fill_2 FILLER_68_812 ();
 sg13g2_fill_2 FILLER_68_832 ();
 sg13g2_fill_1 FILLER_68_834 ();
 sg13g2_fill_2 FILLER_68_864 ();
 sg13g2_fill_1 FILLER_68_866 ();
 sg13g2_decap_8 FILLER_68_909 ();
 sg13g2_fill_1 FILLER_68_916 ();
 sg13g2_fill_2 FILLER_68_969 ();
 sg13g2_fill_1 FILLER_68_1048 ();
 sg13g2_fill_1 FILLER_68_1065 ();
 sg13g2_fill_2 FILLER_68_1075 ();
 sg13g2_fill_2 FILLER_68_1103 ();
 sg13g2_fill_1 FILLER_68_1105 ();
 sg13g2_decap_4 FILLER_68_1114 ();
 sg13g2_fill_2 FILLER_68_1127 ();
 sg13g2_fill_1 FILLER_68_1129 ();
 sg13g2_fill_1 FILLER_68_1134 ();
 sg13g2_fill_2 FILLER_68_1145 ();
 sg13g2_fill_1 FILLER_68_1147 ();
 sg13g2_fill_2 FILLER_68_1163 ();
 sg13g2_fill_1 FILLER_68_1165 ();
 sg13g2_fill_1 FILLER_68_1180 ();
 sg13g2_fill_1 FILLER_68_1221 ();
 sg13g2_fill_1 FILLER_68_1278 ();
 sg13g2_fill_1 FILLER_68_1305 ();
 sg13g2_fill_1 FILLER_68_1310 ();
 sg13g2_fill_1 FILLER_68_1323 ();
 sg13g2_fill_1 FILLER_68_1333 ();
 sg13g2_fill_1 FILLER_68_1399 ();
 sg13g2_fill_2 FILLER_68_1409 ();
 sg13g2_fill_1 FILLER_68_1447 ();
 sg13g2_fill_1 FILLER_68_1461 ();
 sg13g2_fill_2 FILLER_68_1490 ();
 sg13g2_fill_2 FILLER_68_1518 ();
 sg13g2_fill_2 FILLER_68_1527 ();
 sg13g2_fill_1 FILLER_68_1529 ();
 sg13g2_fill_1 FILLER_68_1556 ();
 sg13g2_fill_2 FILLER_68_1581 ();
 sg13g2_fill_1 FILLER_68_1583 ();
 sg13g2_fill_1 FILLER_68_1693 ();
 sg13g2_fill_2 FILLER_68_1729 ();
 sg13g2_fill_1 FILLER_68_1741 ();
 sg13g2_fill_2 FILLER_69_36 ();
 sg13g2_fill_1 FILLER_69_38 ();
 sg13g2_fill_2 FILLER_69_74 ();
 sg13g2_fill_2 FILLER_69_157 ();
 sg13g2_fill_1 FILLER_69_159 ();
 sg13g2_fill_2 FILLER_69_188 ();
 sg13g2_fill_1 FILLER_69_190 ();
 sg13g2_fill_1 FILLER_69_211 ();
 sg13g2_fill_2 FILLER_69_221 ();
 sg13g2_fill_2 FILLER_69_251 ();
 sg13g2_fill_2 FILLER_69_309 ();
 sg13g2_fill_1 FILLER_69_386 ();
 sg13g2_fill_2 FILLER_69_419 ();
 sg13g2_fill_2 FILLER_69_438 ();
 sg13g2_fill_1 FILLER_69_440 ();
 sg13g2_fill_1 FILLER_69_446 ();
 sg13g2_fill_2 FILLER_69_476 ();
 sg13g2_fill_1 FILLER_69_478 ();
 sg13g2_fill_1 FILLER_69_494 ();
 sg13g2_decap_8 FILLER_69_500 ();
 sg13g2_fill_2 FILLER_69_547 ();
 sg13g2_fill_2 FILLER_69_644 ();
 sg13g2_fill_1 FILLER_69_690 ();
 sg13g2_fill_1 FILLER_69_704 ();
 sg13g2_fill_1 FILLER_69_723 ();
 sg13g2_fill_2 FILLER_69_829 ();
 sg13g2_fill_1 FILLER_69_831 ();
 sg13g2_fill_1 FILLER_69_867 ();
 sg13g2_fill_2 FILLER_69_916 ();
 sg13g2_fill_2 FILLER_69_940 ();
 sg13g2_fill_2 FILLER_69_956 ();
 sg13g2_fill_1 FILLER_69_983 ();
 sg13g2_fill_1 FILLER_69_1007 ();
 sg13g2_fill_1 FILLER_69_1135 ();
 sg13g2_fill_2 FILLER_69_1157 ();
 sg13g2_fill_1 FILLER_69_1159 ();
 sg13g2_fill_1 FILLER_69_1186 ();
 sg13g2_fill_2 FILLER_69_1288 ();
 sg13g2_fill_1 FILLER_69_1318 ();
 sg13g2_fill_2 FILLER_69_1423 ();
 sg13g2_fill_1 FILLER_69_1425 ();
 sg13g2_fill_2 FILLER_69_1439 ();
 sg13g2_fill_1 FILLER_69_1441 ();
 sg13g2_fill_1 FILLER_69_1447 ();
 sg13g2_fill_2 FILLER_69_1488 ();
 sg13g2_fill_2 FILLER_69_1591 ();
 sg13g2_fill_1 FILLER_69_1593 ();
 sg13g2_fill_1 FILLER_69_1604 ();
 sg13g2_fill_2 FILLER_69_1631 ();
 sg13g2_fill_1 FILLER_69_1633 ();
 sg13g2_fill_1 FILLER_69_1647 ();
 sg13g2_fill_1 FILLER_69_1657 ();
 sg13g2_fill_2 FILLER_69_1662 ();
 sg13g2_fill_1 FILLER_69_1676 ();
 sg13g2_fill_1 FILLER_69_1687 ();
 sg13g2_fill_2 FILLER_69_1706 ();
 sg13g2_fill_2 FILLER_69_1744 ();
 sg13g2_fill_2 FILLER_70_4 ();
 sg13g2_fill_1 FILLER_70_55 ();
 sg13g2_fill_1 FILLER_70_105 ();
 sg13g2_fill_2 FILLER_70_110 ();
 sg13g2_fill_1 FILLER_70_112 ();
 sg13g2_fill_2 FILLER_70_164 ();
 sg13g2_fill_2 FILLER_70_247 ();
 sg13g2_fill_2 FILLER_70_254 ();
 sg13g2_fill_1 FILLER_70_290 ();
 sg13g2_fill_1 FILLER_70_308 ();
 sg13g2_fill_1 FILLER_70_328 ();
 sg13g2_fill_1 FILLER_70_362 ();
 sg13g2_fill_2 FILLER_70_429 ();
 sg13g2_fill_1 FILLER_70_457 ();
 sg13g2_fill_1 FILLER_70_467 ();
 sg13g2_fill_1 FILLER_70_507 ();
 sg13g2_fill_2 FILLER_70_514 ();
 sg13g2_fill_1 FILLER_70_521 ();
 sg13g2_fill_1 FILLER_70_558 ();
 sg13g2_decap_4 FILLER_70_563 ();
 sg13g2_fill_1 FILLER_70_567 ();
 sg13g2_fill_2 FILLER_70_611 ();
 sg13g2_fill_1 FILLER_70_613 ();
 sg13g2_fill_1 FILLER_70_619 ();
 sg13g2_fill_1 FILLER_70_652 ();
 sg13g2_fill_2 FILLER_70_663 ();
 sg13g2_fill_1 FILLER_70_670 ();
 sg13g2_fill_1 FILLER_70_681 ();
 sg13g2_fill_1 FILLER_70_716 ();
 sg13g2_fill_2 FILLER_70_786 ();
 sg13g2_fill_1 FILLER_70_828 ();
 sg13g2_decap_4 FILLER_70_900 ();
 sg13g2_decap_8 FILLER_70_908 ();
 sg13g2_fill_1 FILLER_70_956 ();
 sg13g2_fill_1 FILLER_70_1017 ();
 sg13g2_fill_2 FILLER_70_1069 ();
 sg13g2_fill_2 FILLER_70_1104 ();
 sg13g2_fill_2 FILLER_70_1161 ();
 sg13g2_fill_2 FILLER_70_1231 ();
 sg13g2_fill_1 FILLER_70_1233 ();
 sg13g2_fill_2 FILLER_70_1260 ();
 sg13g2_fill_1 FILLER_70_1283 ();
 sg13g2_fill_2 FILLER_70_1322 ();
 sg13g2_fill_2 FILLER_70_1328 ();
 sg13g2_fill_2 FILLER_70_1334 ();
 sg13g2_fill_2 FILLER_70_1359 ();
 sg13g2_fill_1 FILLER_70_1361 ();
 sg13g2_fill_1 FILLER_70_1372 ();
 sg13g2_fill_1 FILLER_70_1396 ();
 sg13g2_fill_2 FILLER_70_1446 ();
 sg13g2_fill_2 FILLER_70_1467 ();
 sg13g2_fill_1 FILLER_70_1510 ();
 sg13g2_fill_2 FILLER_70_1537 ();
 sg13g2_fill_1 FILLER_70_1570 ();
 sg13g2_fill_1 FILLER_70_1634 ();
 sg13g2_fill_2 FILLER_70_1652 ();
 sg13g2_fill_1 FILLER_70_1664 ();
 sg13g2_fill_1 FILLER_70_1669 ();
 sg13g2_decap_4 FILLER_70_1679 ();
 sg13g2_fill_2 FILLER_70_1683 ();
 sg13g2_fill_2 FILLER_70_1729 ();
 sg13g2_fill_1 FILLER_70_1750 ();
 sg13g2_fill_2 FILLER_70_1765 ();
 sg13g2_fill_1 FILLER_70_1767 ();
 sg13g2_fill_1 FILLER_71_63 ();
 sg13g2_fill_2 FILLER_71_89 ();
 sg13g2_fill_2 FILLER_71_131 ();
 sg13g2_fill_1 FILLER_71_133 ();
 sg13g2_fill_2 FILLER_71_152 ();
 sg13g2_fill_1 FILLER_71_154 ();
 sg13g2_fill_1 FILLER_71_212 ();
 sg13g2_fill_2 FILLER_71_217 ();
 sg13g2_fill_1 FILLER_71_219 ();
 sg13g2_fill_2 FILLER_71_269 ();
 sg13g2_fill_2 FILLER_71_289 ();
 sg13g2_fill_2 FILLER_71_296 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_fill_2 FILLER_71_472 ();
 sg13g2_fill_2 FILLER_71_494 ();
 sg13g2_fill_2 FILLER_71_522 ();
 sg13g2_decap_8 FILLER_71_557 ();
 sg13g2_fill_1 FILLER_71_564 ();
 sg13g2_fill_2 FILLER_71_622 ();
 sg13g2_fill_1 FILLER_71_624 ();
 sg13g2_fill_1 FILLER_71_651 ();
 sg13g2_fill_2 FILLER_71_804 ();
 sg13g2_fill_1 FILLER_71_806 ();
 sg13g2_fill_2 FILLER_71_853 ();
 sg13g2_fill_2 FILLER_71_873 ();
 sg13g2_decap_8 FILLER_71_919 ();
 sg13g2_decap_8 FILLER_71_930 ();
 sg13g2_fill_2 FILLER_71_937 ();
 sg13g2_fill_1 FILLER_71_939 ();
 sg13g2_fill_1 FILLER_71_963 ();
 sg13g2_fill_2 FILLER_71_983 ();
 sg13g2_fill_1 FILLER_71_1026 ();
 sg13g2_fill_2 FILLER_71_1086 ();
 sg13g2_fill_1 FILLER_71_1119 ();
 sg13g2_fill_2 FILLER_71_1134 ();
 sg13g2_fill_1 FILLER_71_1136 ();
 sg13g2_fill_2 FILLER_71_1155 ();
 sg13g2_fill_1 FILLER_71_1215 ();
 sg13g2_fill_1 FILLER_71_1234 ();
 sg13g2_fill_1 FILLER_71_1275 ();
 sg13g2_fill_1 FILLER_71_1338 ();
 sg13g2_fill_1 FILLER_71_1343 ();
 sg13g2_fill_1 FILLER_71_1367 ();
 sg13g2_fill_2 FILLER_71_1424 ();
 sg13g2_fill_1 FILLER_71_1448 ();
 sg13g2_fill_2 FILLER_71_1486 ();
 sg13g2_fill_1 FILLER_71_1503 ();
 sg13g2_fill_1 FILLER_71_1567 ();
 sg13g2_fill_2 FILLER_71_1598 ();
 sg13g2_fill_2 FILLER_71_1705 ();
 sg13g2_fill_2 FILLER_71_1765 ();
 sg13g2_fill_1 FILLER_71_1767 ();
 sg13g2_fill_2 FILLER_72_26 ();
 sg13g2_fill_2 FILLER_72_80 ();
 sg13g2_fill_2 FILLER_72_147 ();
 sg13g2_fill_1 FILLER_72_149 ();
 sg13g2_fill_2 FILLER_72_155 ();
 sg13g2_fill_1 FILLER_72_351 ();
 sg13g2_fill_2 FILLER_72_372 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_fill_1 FILLER_72_413 ();
 sg13g2_fill_2 FILLER_72_419 ();
 sg13g2_fill_1 FILLER_72_421 ();
 sg13g2_decap_4 FILLER_72_426 ();
 sg13g2_fill_2 FILLER_72_441 ();
 sg13g2_fill_1 FILLER_72_443 ();
 sg13g2_fill_1 FILLER_72_459 ();
 sg13g2_fill_1 FILLER_72_473 ();
 sg13g2_fill_1 FILLER_72_507 ();
 sg13g2_fill_2 FILLER_72_542 ();
 sg13g2_fill_1 FILLER_72_570 ();
 sg13g2_fill_2 FILLER_72_584 ();
 sg13g2_fill_1 FILLER_72_586 ();
 sg13g2_fill_2 FILLER_72_602 ();
 sg13g2_fill_2 FILLER_72_618 ();
 sg13g2_fill_1 FILLER_72_620 ();
 sg13g2_fill_1 FILLER_72_702 ();
 sg13g2_fill_2 FILLER_72_739 ();
 sg13g2_fill_1 FILLER_72_803 ();
 sg13g2_fill_2 FILLER_72_812 ();
 sg13g2_fill_2 FILLER_72_840 ();
 sg13g2_fill_1 FILLER_72_842 ();
 sg13g2_decap_4 FILLER_72_879 ();
 sg13g2_decap_4 FILLER_72_919 ();
 sg13g2_fill_2 FILLER_72_923 ();
 sg13g2_fill_2 FILLER_72_1019 ();
 sg13g2_fill_2 FILLER_72_1026 ();
 sg13g2_fill_1 FILLER_72_1046 ();
 sg13g2_fill_2 FILLER_72_1119 ();
 sg13g2_fill_1 FILLER_72_1155 ();
 sg13g2_fill_2 FILLER_72_1180 ();
 sg13g2_fill_1 FILLER_72_1244 ();
 sg13g2_fill_1 FILLER_72_1249 ();
 sg13g2_fill_1 FILLER_72_1254 ();
 sg13g2_fill_1 FILLER_72_1295 ();
 sg13g2_fill_2 FILLER_72_1306 ();
 sg13g2_fill_1 FILLER_72_1348 ();
 sg13g2_fill_2 FILLER_72_1456 ();
 sg13g2_fill_2 FILLER_72_1494 ();
 sg13g2_fill_1 FILLER_72_1572 ();
 sg13g2_fill_2 FILLER_72_1583 ();
 sg13g2_fill_2 FILLER_72_1591 ();
 sg13g2_fill_2 FILLER_72_1612 ();
 sg13g2_fill_1 FILLER_72_1614 ();
 sg13g2_decap_8 FILLER_72_1663 ();
 sg13g2_fill_2 FILLER_72_1670 ();
 sg13g2_fill_2 FILLER_72_1708 ();
 sg13g2_fill_2 FILLER_72_1758 ();
 sg13g2_fill_2 FILLER_73_55 ();
 sg13g2_fill_1 FILLER_73_78 ();
 sg13g2_fill_2 FILLER_73_103 ();
 sg13g2_fill_1 FILLER_73_105 ();
 sg13g2_fill_2 FILLER_73_153 ();
 sg13g2_fill_2 FILLER_73_165 ();
 sg13g2_fill_1 FILLER_73_167 ();
 sg13g2_fill_2 FILLER_73_289 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_fill_1 FILLER_73_310 ();
 sg13g2_fill_1 FILLER_73_343 ();
 sg13g2_fill_1 FILLER_73_363 ();
 sg13g2_fill_1 FILLER_73_384 ();
 sg13g2_fill_2 FILLER_73_399 ();
 sg13g2_fill_2 FILLER_73_411 ();
 sg13g2_fill_1 FILLER_73_428 ();
 sg13g2_fill_1 FILLER_73_447 ();
 sg13g2_fill_2 FILLER_73_458 ();
 sg13g2_fill_1 FILLER_73_460 ();
 sg13g2_fill_1 FILLER_73_467 ();
 sg13g2_fill_2 FILLER_73_473 ();
 sg13g2_fill_1 FILLER_73_475 ();
 sg13g2_fill_1 FILLER_73_546 ();
 sg13g2_fill_2 FILLER_73_574 ();
 sg13g2_fill_1 FILLER_73_576 ();
 sg13g2_fill_2 FILLER_73_601 ();
 sg13g2_fill_2 FILLER_73_696 ();
 sg13g2_fill_1 FILLER_73_718 ();
 sg13g2_fill_2 FILLER_73_739 ();
 sg13g2_fill_1 FILLER_73_782 ();
 sg13g2_fill_1 FILLER_73_823 ();
 sg13g2_fill_1 FILLER_73_834 ();
 sg13g2_decap_4 FILLER_73_844 ();
 sg13g2_fill_1 FILLER_73_848 ();
 sg13g2_fill_2 FILLER_73_885 ();
 sg13g2_fill_1 FILLER_73_913 ();
 sg13g2_fill_2 FILLER_73_1083 ();
 sg13g2_fill_2 FILLER_73_1094 ();
 sg13g2_fill_1 FILLER_73_1096 ();
 sg13g2_fill_2 FILLER_73_1144 ();
 sg13g2_fill_2 FILLER_73_1160 ();
 sg13g2_decap_4 FILLER_73_1216 ();
 sg13g2_fill_2 FILLER_73_1220 ();
 sg13g2_fill_2 FILLER_73_1231 ();
 sg13g2_fill_1 FILLER_73_1233 ();
 sg13g2_fill_2 FILLER_73_1243 ();
 sg13g2_fill_2 FILLER_73_1258 ();
 sg13g2_fill_2 FILLER_73_1331 ();
 sg13g2_fill_2 FILLER_73_1365 ();
 sg13g2_fill_1 FILLER_73_1367 ();
 sg13g2_fill_2 FILLER_73_1376 ();
 sg13g2_fill_1 FILLER_73_1378 ();
 sg13g2_fill_2 FILLER_73_1402 ();
 sg13g2_fill_1 FILLER_73_1404 ();
 sg13g2_fill_1 FILLER_73_1458 ();
 sg13g2_fill_1 FILLER_73_1667 ();
 sg13g2_fill_2 FILLER_73_1694 ();
 sg13g2_fill_2 FILLER_73_1716 ();
 sg13g2_fill_1 FILLER_73_1748 ();
 sg13g2_decap_8 FILLER_73_1757 ();
 sg13g2_decap_4 FILLER_73_1764 ();
 sg13g2_fill_1 FILLER_74_4 ();
 sg13g2_fill_1 FILLER_74_50 ();
 sg13g2_fill_2 FILLER_74_77 ();
 sg13g2_fill_1 FILLER_74_79 ();
 sg13g2_fill_2 FILLER_74_110 ();
 sg13g2_fill_2 FILLER_74_142 ();
 sg13g2_fill_2 FILLER_74_152 ();
 sg13g2_fill_1 FILLER_74_154 ();
 sg13g2_fill_1 FILLER_74_248 ();
 sg13g2_fill_1 FILLER_74_368 ();
 sg13g2_fill_1 FILLER_74_378 ();
 sg13g2_fill_1 FILLER_74_416 ();
 sg13g2_fill_2 FILLER_74_423 ();
 sg13g2_fill_1 FILLER_74_425 ();
 sg13g2_fill_1 FILLER_74_434 ();
 sg13g2_fill_2 FILLER_74_489 ();
 sg13g2_fill_1 FILLER_74_495 ();
 sg13g2_decap_8 FILLER_74_533 ();
 sg13g2_decap_4 FILLER_74_540 ();
 sg13g2_fill_1 FILLER_74_570 ();
 sg13g2_fill_1 FILLER_74_625 ();
 sg13g2_fill_2 FILLER_74_639 ();
 sg13g2_fill_2 FILLER_74_759 ();
 sg13g2_fill_2 FILLER_74_769 ();
 sg13g2_fill_1 FILLER_74_771 ();
 sg13g2_decap_4 FILLER_74_780 ();
 sg13g2_fill_1 FILLER_74_794 ();
 sg13g2_fill_2 FILLER_74_812 ();
 sg13g2_fill_1 FILLER_74_814 ();
 sg13g2_fill_2 FILLER_74_851 ();
 sg13g2_fill_1 FILLER_74_874 ();
 sg13g2_decap_4 FILLER_74_911 ();
 sg13g2_fill_1 FILLER_74_915 ();
 sg13g2_decap_4 FILLER_74_921 ();
 sg13g2_fill_1 FILLER_74_925 ();
 sg13g2_fill_1 FILLER_74_962 ();
 sg13g2_fill_1 FILLER_74_1007 ();
 sg13g2_fill_1 FILLER_74_1017 ();
 sg13g2_fill_1 FILLER_74_1072 ();
 sg13g2_fill_2 FILLER_74_1099 ();
 sg13g2_fill_1 FILLER_74_1101 ();
 sg13g2_fill_1 FILLER_74_1128 ();
 sg13g2_fill_2 FILLER_74_1134 ();
 sg13g2_fill_1 FILLER_74_1136 ();
 sg13g2_decap_8 FILLER_74_1201 ();
 sg13g2_decap_4 FILLER_74_1208 ();
 sg13g2_fill_1 FILLER_74_1212 ();
 sg13g2_fill_2 FILLER_74_1217 ();
 sg13g2_fill_2 FILLER_74_1265 ();
 sg13g2_fill_2 FILLER_74_1326 ();
 sg13g2_fill_1 FILLER_74_1328 ();
 sg13g2_fill_1 FILLER_74_1347 ();
 sg13g2_fill_2 FILLER_74_1416 ();
 sg13g2_fill_1 FILLER_74_1418 ();
 sg13g2_fill_2 FILLER_74_1432 ();
 sg13g2_fill_1 FILLER_74_1528 ();
 sg13g2_fill_2 FILLER_74_1551 ();
 sg13g2_fill_1 FILLER_74_1553 ();
 sg13g2_fill_2 FILLER_74_1567 ();
 sg13g2_fill_1 FILLER_74_1569 ();
 sg13g2_fill_2 FILLER_74_1583 ();
 sg13g2_fill_1 FILLER_74_1585 ();
 sg13g2_fill_2 FILLER_74_1605 ();
 sg13g2_fill_1 FILLER_74_1607 ();
 sg13g2_fill_2 FILLER_74_1629 ();
 sg13g2_fill_1 FILLER_74_1631 ();
 sg13g2_fill_2 FILLER_74_1650 ();
 sg13g2_fill_2 FILLER_74_1656 ();
 sg13g2_fill_2 FILLER_74_1672 ();
 sg13g2_fill_1 FILLER_74_1674 ();
 sg13g2_fill_2 FILLER_74_1706 ();
 sg13g2_decap_8 FILLER_74_1744 ();
 sg13g2_decap_8 FILLER_74_1751 ();
 sg13g2_decap_8 FILLER_74_1758 ();
 sg13g2_fill_2 FILLER_74_1765 ();
 sg13g2_fill_1 FILLER_74_1767 ();
 sg13g2_fill_1 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_71 ();
 sg13g2_fill_1 FILLER_75_149 ();
 sg13g2_fill_1 FILLER_75_204 ();
 sg13g2_fill_1 FILLER_75_410 ();
 sg13g2_fill_1 FILLER_75_416 ();
 sg13g2_fill_2 FILLER_75_425 ();
 sg13g2_fill_1 FILLER_75_427 ();
 sg13g2_fill_1 FILLER_75_434 ();
 sg13g2_fill_1 FILLER_75_464 ();
 sg13g2_fill_1 FILLER_75_473 ();
 sg13g2_fill_1 FILLER_75_486 ();
 sg13g2_fill_1 FILLER_75_495 ();
 sg13g2_fill_1 FILLER_75_517 ();
 sg13g2_decap_8 FILLER_75_522 ();
 sg13g2_decap_8 FILLER_75_529 ();
 sg13g2_fill_1 FILLER_75_536 ();
 sg13g2_fill_2 FILLER_75_564 ();
 sg13g2_fill_1 FILLER_75_566 ();
 sg13g2_fill_1 FILLER_75_585 ();
 sg13g2_fill_2 FILLER_75_596 ();
 sg13g2_fill_1 FILLER_75_598 ();
 sg13g2_fill_2 FILLER_75_612 ();
 sg13g2_fill_2 FILLER_75_624 ();
 sg13g2_fill_1 FILLER_75_691 ();
 sg13g2_fill_2 FILLER_75_711 ();
 sg13g2_fill_2 FILLER_75_759 ();
 sg13g2_fill_2 FILLER_75_817 ();
 sg13g2_fill_1 FILLER_75_828 ();
 sg13g2_fill_2 FILLER_75_834 ();
 sg13g2_fill_2 FILLER_75_903 ();
 sg13g2_fill_2 FILLER_75_945 ();
 sg13g2_fill_1 FILLER_75_978 ();
 sg13g2_fill_2 FILLER_75_1085 ();
 sg13g2_fill_2 FILLER_75_1125 ();
 sg13g2_fill_1 FILLER_75_1127 ();
 sg13g2_fill_1 FILLER_75_1163 ();
 sg13g2_fill_2 FILLER_75_1200 ();
 sg13g2_fill_2 FILLER_75_1242 ();
 sg13g2_fill_1 FILLER_75_1266 ();
 sg13g2_fill_1 FILLER_75_1318 ();
 sg13g2_fill_2 FILLER_75_1397 ();
 sg13g2_fill_2 FILLER_75_1435 ();
 sg13g2_fill_2 FILLER_75_1451 ();
 sg13g2_fill_2 FILLER_75_1468 ();
 sg13g2_fill_1 FILLER_75_1470 ();
 sg13g2_fill_2 FILLER_75_1500 ();
 sg13g2_fill_1 FILLER_75_1502 ();
 sg13g2_fill_2 FILLER_75_1512 ();
 sg13g2_fill_2 FILLER_75_1545 ();
 sg13g2_fill_2 FILLER_75_1570 ();
 sg13g2_fill_1 FILLER_75_1582 ();
 sg13g2_fill_1 FILLER_75_1619 ();
 sg13g2_fill_1 FILLER_75_1661 ();
 sg13g2_decap_4 FILLER_75_1719 ();
 sg13g2_fill_1 FILLER_75_1723 ();
 sg13g2_decap_8 FILLER_75_1750 ();
 sg13g2_decap_8 FILLER_75_1757 ();
 sg13g2_decap_4 FILLER_75_1764 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_5 ();
 sg13g2_fill_2 FILLER_76_47 ();
 sg13g2_fill_1 FILLER_76_49 ();
 sg13g2_fill_2 FILLER_76_60 ();
 sg13g2_fill_1 FILLER_76_114 ();
 sg13g2_fill_2 FILLER_76_139 ();
 sg13g2_fill_1 FILLER_76_141 ();
 sg13g2_fill_1 FILLER_76_168 ();
 sg13g2_fill_2 FILLER_76_202 ();
 sg13g2_fill_1 FILLER_76_217 ();
 sg13g2_fill_2 FILLER_76_246 ();
 sg13g2_fill_1 FILLER_76_248 ();
 sg13g2_fill_1 FILLER_76_259 ();
 sg13g2_fill_1 FILLER_76_312 ();
 sg13g2_fill_2 FILLER_76_391 ();
 sg13g2_fill_1 FILLER_76_428 ();
 sg13g2_fill_1 FILLER_76_465 ();
 sg13g2_fill_2 FILLER_76_532 ();
 sg13g2_fill_1 FILLER_76_534 ();
 sg13g2_fill_1 FILLER_76_561 ();
 sg13g2_fill_2 FILLER_76_583 ();
 sg13g2_fill_2 FILLER_76_660 ();
 sg13g2_fill_1 FILLER_76_662 ();
 sg13g2_fill_2 FILLER_76_689 ();
 sg13g2_fill_2 FILLER_76_814 ();
 sg13g2_fill_1 FILLER_76_831 ();
 sg13g2_fill_2 FILLER_76_841 ();
 sg13g2_fill_2 FILLER_76_857 ();
 sg13g2_fill_1 FILLER_76_873 ();
 sg13g2_decap_4 FILLER_76_910 ();
 sg13g2_fill_1 FILLER_76_914 ();
 sg13g2_fill_2 FILLER_76_944 ();
 sg13g2_fill_1 FILLER_76_956 ();
 sg13g2_fill_2 FILLER_76_1009 ();
 sg13g2_fill_1 FILLER_76_1011 ();
 sg13g2_fill_1 FILLER_76_1033 ();
 sg13g2_fill_1 FILLER_76_1042 ();
 sg13g2_fill_2 FILLER_76_1115 ();
 sg13g2_fill_2 FILLER_76_1172 ();
 sg13g2_fill_1 FILLER_76_1227 ();
 sg13g2_fill_1 FILLER_76_1300 ();
 sg13g2_fill_2 FILLER_76_1310 ();
 sg13g2_fill_1 FILLER_76_1312 ();
 sg13g2_fill_2 FILLER_76_1328 ();
 sg13g2_fill_2 FILLER_76_1361 ();
 sg13g2_fill_1 FILLER_76_1363 ();
 sg13g2_fill_2 FILLER_76_1373 ();
 sg13g2_fill_1 FILLER_76_1375 ();
 sg13g2_fill_1 FILLER_76_1404 ();
 sg13g2_fill_2 FILLER_76_1460 ();
 sg13g2_fill_1 FILLER_76_1462 ();
 sg13g2_fill_1 FILLER_76_1585 ();
 sg13g2_fill_2 FILLER_76_1617 ();
 sg13g2_fill_1 FILLER_76_1619 ();
 sg13g2_fill_1 FILLER_76_1691 ();
 sg13g2_decap_8 FILLER_76_1713 ();
 sg13g2_decap_8 FILLER_76_1746 ();
 sg13g2_decap_8 FILLER_76_1753 ();
 sg13g2_decap_8 FILLER_76_1760 ();
 sg13g2_fill_1 FILLER_76_1767 ();
 sg13g2_fill_2 FILLER_77_35 ();
 sg13g2_fill_2 FILLER_77_63 ();
 sg13g2_fill_1 FILLER_77_65 ();
 sg13g2_fill_1 FILLER_77_142 ();
 sg13g2_fill_1 FILLER_77_148 ();
 sg13g2_fill_1 FILLER_77_190 ();
 sg13g2_fill_1 FILLER_77_217 ();
 sg13g2_fill_2 FILLER_77_309 ();
 sg13g2_fill_2 FILLER_77_337 ();
 sg13g2_fill_1 FILLER_77_402 ();
 sg13g2_fill_2 FILLER_77_416 ();
 sg13g2_fill_2 FILLER_77_445 ();
 sg13g2_fill_2 FILLER_77_475 ();
 sg13g2_fill_1 FILLER_77_492 ();
 sg13g2_fill_2 FILLER_77_612 ();
 sg13g2_fill_2 FILLER_77_654 ();
 sg13g2_fill_1 FILLER_77_656 ();
 sg13g2_fill_2 FILLER_77_661 ();
 sg13g2_fill_2 FILLER_77_701 ();
 sg13g2_fill_1 FILLER_77_791 ();
 sg13g2_fill_1 FILLER_77_884 ();
 sg13g2_fill_2 FILLER_77_899 ();
 sg13g2_fill_2 FILLER_77_922 ();
 sg13g2_fill_2 FILLER_77_1021 ();
 sg13g2_fill_1 FILLER_77_1079 ();
 sg13g2_fill_2 FILLER_77_1089 ();
 sg13g2_decap_4 FILLER_77_1117 ();
 sg13g2_fill_1 FILLER_77_1121 ();
 sg13g2_fill_2 FILLER_77_1172 ();
 sg13g2_fill_1 FILLER_77_1174 ();
 sg13g2_fill_2 FILLER_77_1198 ();
 sg13g2_fill_1 FILLER_77_1200 ();
 sg13g2_fill_1 FILLER_77_1255 ();
 sg13g2_fill_2 FILLER_77_1342 ();
 sg13g2_fill_1 FILLER_77_1375 ();
 sg13g2_fill_1 FILLER_77_1381 ();
 sg13g2_fill_2 FILLER_77_1412 ();
 sg13g2_fill_2 FILLER_77_1440 ();
 sg13g2_fill_2 FILLER_77_1492 ();
 sg13g2_fill_2 FILLER_77_1525 ();
 sg13g2_fill_1 FILLER_77_1527 ();
 sg13g2_fill_2 FILLER_77_1554 ();
 sg13g2_fill_2 FILLER_77_1592 ();
 sg13g2_fill_2 FILLER_77_1660 ();
 sg13g2_fill_2 FILLER_77_1672 ();
 sg13g2_fill_1 FILLER_77_1674 ();
 sg13g2_fill_1 FILLER_77_1711 ();
 sg13g2_decap_4 FILLER_77_1722 ();
 sg13g2_fill_1 FILLER_77_1726 ();
 sg13g2_decap_8 FILLER_77_1740 ();
 sg13g2_decap_8 FILLER_77_1747 ();
 sg13g2_decap_8 FILLER_77_1754 ();
 sg13g2_decap_8 FILLER_77_1761 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_6 ();
 sg13g2_fill_1 FILLER_78_8 ();
 sg13g2_fill_1 FILLER_78_51 ();
 sg13g2_fill_1 FILLER_78_82 ();
 sg13g2_fill_2 FILLER_78_97 ();
 sg13g2_fill_1 FILLER_78_99 ();
 sg13g2_fill_2 FILLER_78_126 ();
 sg13g2_fill_1 FILLER_78_128 ();
 sg13g2_fill_2 FILLER_78_155 ();
 sg13g2_fill_1 FILLER_78_157 ();
 sg13g2_fill_1 FILLER_78_207 ();
 sg13g2_fill_2 FILLER_78_273 ();
 sg13g2_fill_1 FILLER_78_275 ();
 sg13g2_fill_2 FILLER_78_300 ();
 sg13g2_fill_1 FILLER_78_464 ();
 sg13g2_fill_2 FILLER_78_490 ();
 sg13g2_fill_1 FILLER_78_497 ();
 sg13g2_fill_1 FILLER_78_508 ();
 sg13g2_fill_2 FILLER_78_557 ();
 sg13g2_fill_2 FILLER_78_574 ();
 sg13g2_fill_2 FILLER_78_590 ();
 sg13g2_fill_2 FILLER_78_601 ();
 sg13g2_fill_1 FILLER_78_727 ();
 sg13g2_fill_2 FILLER_78_754 ();
 sg13g2_fill_1 FILLER_78_756 ();
 sg13g2_fill_2 FILLER_78_767 ();
 sg13g2_fill_1 FILLER_78_769 ();
 sg13g2_fill_2 FILLER_78_820 ();
 sg13g2_fill_1 FILLER_78_854 ();
 sg13g2_decap_4 FILLER_78_881 ();
 sg13g2_fill_2 FILLER_78_965 ();
 sg13g2_fill_2 FILLER_78_976 ();
 sg13g2_fill_2 FILLER_78_1012 ();
 sg13g2_fill_1 FILLER_78_1014 ();
 sg13g2_fill_1 FILLER_78_1039 ();
 sg13g2_fill_2 FILLER_78_1157 ();
 sg13g2_fill_1 FILLER_78_1199 ();
 sg13g2_fill_2 FILLER_78_1226 ();
 sg13g2_fill_2 FILLER_78_1253 ();
 sg13g2_fill_1 FILLER_78_1255 ();
 sg13g2_fill_1 FILLER_78_1290 ();
 sg13g2_fill_2 FILLER_78_1306 ();
 sg13g2_fill_1 FILLER_78_1308 ();
 sg13g2_fill_2 FILLER_78_1329 ();
 sg13g2_fill_1 FILLER_78_1336 ();
 sg13g2_fill_1 FILLER_78_1368 ();
 sg13g2_fill_2 FILLER_78_1403 ();
 sg13g2_fill_1 FILLER_78_1405 ();
 sg13g2_fill_2 FILLER_78_1420 ();
 sg13g2_fill_2 FILLER_78_1453 ();
 sg13g2_fill_1 FILLER_78_1455 ();
 sg13g2_fill_1 FILLER_78_1495 ();
 sg13g2_fill_2 FILLER_78_1554 ();
 sg13g2_fill_2 FILLER_78_1608 ();
 sg13g2_fill_2 FILLER_78_1636 ();
 sg13g2_fill_2 FILLER_78_1664 ();
 sg13g2_fill_2 FILLER_78_1692 ();
 sg13g2_fill_1 FILLER_78_1694 ();
 sg13g2_decap_8 FILLER_78_1736 ();
 sg13g2_decap_8 FILLER_78_1743 ();
 sg13g2_decap_8 FILLER_78_1750 ();
 sg13g2_decap_8 FILLER_78_1757 ();
 sg13g2_decap_4 FILLER_78_1764 ();
 sg13g2_fill_1 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_9 ();
 sg13g2_fill_1 FILLER_79_104 ();
 sg13g2_fill_2 FILLER_79_119 ();
 sg13g2_fill_1 FILLER_79_121 ();
 sg13g2_fill_1 FILLER_79_173 ();
 sg13g2_fill_1 FILLER_79_214 ();
 sg13g2_fill_2 FILLER_79_229 ();
 sg13g2_fill_2 FILLER_79_364 ();
 sg13g2_fill_1 FILLER_79_423 ();
 sg13g2_fill_2 FILLER_79_502 ();
 sg13g2_fill_2 FILLER_79_512 ();
 sg13g2_fill_1 FILLER_79_514 ();
 sg13g2_fill_2 FILLER_79_611 ();
 sg13g2_fill_1 FILLER_79_613 ();
 sg13g2_fill_2 FILLER_79_633 ();
 sg13g2_fill_2 FILLER_79_667 ();
 sg13g2_fill_1 FILLER_79_669 ();
 sg13g2_fill_1 FILLER_79_689 ();
 sg13g2_fill_2 FILLER_79_747 ();
 sg13g2_fill_1 FILLER_79_749 ();
 sg13g2_fill_2 FILLER_79_805 ();
 sg13g2_fill_1 FILLER_79_859 ();
 sg13g2_fill_1 FILLER_79_911 ();
 sg13g2_fill_2 FILLER_79_921 ();
 sg13g2_fill_1 FILLER_79_923 ();
 sg13g2_fill_2 FILLER_79_934 ();
 sg13g2_fill_1 FILLER_79_958 ();
 sg13g2_fill_1 FILLER_79_1133 ();
 sg13g2_fill_2 FILLER_79_1188 ();
 sg13g2_fill_1 FILLER_79_1190 ();
 sg13g2_fill_2 FILLER_79_1217 ();
 sg13g2_fill_1 FILLER_79_1219 ();
 sg13g2_fill_1 FILLER_79_1362 ();
 sg13g2_fill_1 FILLER_79_1508 ();
 sg13g2_fill_2 FILLER_79_1580 ();
 sg13g2_fill_1 FILLER_79_1592 ();
 sg13g2_fill_2 FILLER_79_1630 ();
 sg13g2_fill_1 FILLER_79_1632 ();
 sg13g2_decap_8 FILLER_79_1668 ();
 sg13g2_fill_2 FILLER_79_1692 ();
 sg13g2_fill_1 FILLER_79_1694 ();
 sg13g2_decap_8 FILLER_79_1708 ();
 sg13g2_decap_4 FILLER_79_1715 ();
 sg13g2_fill_1 FILLER_79_1719 ();
 sg13g2_decap_8 FILLER_79_1733 ();
 sg13g2_decap_8 FILLER_79_1740 ();
 sg13g2_decap_8 FILLER_79_1747 ();
 sg13g2_decap_8 FILLER_79_1754 ();
 sg13g2_decap_8 FILLER_79_1761 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_14 ();
 sg13g2_fill_2 FILLER_80_45 ();
 sg13g2_fill_1 FILLER_80_74 ();
 sg13g2_fill_2 FILLER_80_134 ();
 sg13g2_fill_2 FILLER_80_149 ();
 sg13g2_fill_1 FILLER_80_151 ();
 sg13g2_fill_2 FILLER_80_161 ();
 sg13g2_fill_2 FILLER_80_280 ();
 sg13g2_fill_2 FILLER_80_299 ();
 sg13g2_fill_1 FILLER_80_301 ();
 sg13g2_fill_2 FILLER_80_342 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_fill_2 FILLER_80_357 ();
 sg13g2_fill_2 FILLER_80_395 ();
 sg13g2_fill_1 FILLER_80_397 ();
 sg13g2_decap_8 FILLER_80_439 ();
 sg13g2_decap_4 FILLER_80_446 ();
 sg13g2_fill_1 FILLER_80_450 ();
 sg13g2_decap_4 FILLER_80_459 ();
 sg13g2_fill_1 FILLER_80_496 ();
 sg13g2_fill_2 FILLER_80_597 ();
 sg13g2_fill_1 FILLER_80_599 ();
 sg13g2_fill_2 FILLER_80_640 ();
 sg13g2_fill_1 FILLER_80_642 ();
 sg13g2_fill_2 FILLER_80_786 ();
 sg13g2_fill_1 FILLER_80_788 ();
 sg13g2_fill_2 FILLER_80_815 ();
 sg13g2_fill_2 FILLER_80_837 ();
 sg13g2_fill_2 FILLER_80_862 ();
 sg13g2_fill_1 FILLER_80_864 ();
 sg13g2_fill_2 FILLER_80_878 ();
 sg13g2_fill_1 FILLER_80_928 ();
 sg13g2_fill_2 FILLER_80_959 ();
 sg13g2_decap_4 FILLER_80_984 ();
 sg13g2_fill_2 FILLER_80_988 ();
 sg13g2_fill_2 FILLER_80_1051 ();
 sg13g2_fill_1 FILLER_80_1053 ();
 sg13g2_fill_1 FILLER_80_1093 ();
 sg13g2_fill_1 FILLER_80_1111 ();
 sg13g2_fill_2 FILLER_80_1150 ();
 sg13g2_fill_1 FILLER_80_1152 ();
 sg13g2_fill_2 FILLER_80_1162 ();
 sg13g2_fill_2 FILLER_80_1199 ();
 sg13g2_fill_1 FILLER_80_1254 ();
 sg13g2_fill_1 FILLER_80_1307 ();
 sg13g2_fill_2 FILLER_80_1333 ();
 sg13g2_fill_1 FILLER_80_1350 ();
 sg13g2_fill_1 FILLER_80_1360 ();
 sg13g2_fill_2 FILLER_80_1404 ();
 sg13g2_fill_1 FILLER_80_1406 ();
 sg13g2_fill_2 FILLER_80_1459 ();
 sg13g2_fill_2 FILLER_80_1484 ();
 sg13g2_fill_2 FILLER_80_1515 ();
 sg13g2_fill_1 FILLER_80_1517 ();
 sg13g2_fill_1 FILLER_80_1553 ();
 sg13g2_fill_1 FILLER_80_1585 ();
 sg13g2_fill_1 FILLER_80_1638 ();
 sg13g2_decap_8 FILLER_80_1664 ();
 sg13g2_decap_8 FILLER_80_1671 ();
 sg13g2_decap_8 FILLER_80_1678 ();
 sg13g2_decap_8 FILLER_80_1685 ();
 sg13g2_decap_8 FILLER_80_1692 ();
 sg13g2_decap_8 FILLER_80_1699 ();
 sg13g2_decap_8 FILLER_80_1706 ();
 sg13g2_decap_8 FILLER_80_1713 ();
 sg13g2_decap_8 FILLER_80_1720 ();
 sg13g2_decap_8 FILLER_80_1727 ();
 sg13g2_decap_8 FILLER_80_1734 ();
 sg13g2_decap_8 FILLER_80_1741 ();
 sg13g2_decap_8 FILLER_80_1748 ();
 sg13g2_decap_8 FILLER_80_1755 ();
 sg13g2_decap_4 FILLER_80_1762 ();
 sg13g2_fill_2 FILLER_80_1766 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net2128;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net16;
 assign uio_oe[4] = net2129;
 assign uio_oe[5] = net17;
 assign uio_oe[6] = net18;
 assign uio_oe[7] = net19;
 assign uio_out[0] = net20;
 assign uio_out[2] = net21;
 assign uio_out[3] = net22;
 assign uio_out[5] = net23;
 assign uio_out[6] = net24;
 assign uio_out[7] = net25;
endmodule
