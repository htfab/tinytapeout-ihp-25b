module tt_um_alif_single_dualleak (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire params_ready;
 wire spike_out;
 wire \system_inst.leak_cycles_1[0] ;
 wire \system_inst.leak_cycles_1[1] ;
 wire \system_inst.leak_cycles_1[2] ;
 wire \system_inst.leak_cycles_1[3] ;
 wire \system_inst.leak_cycles_2[0] ;
 wire \system_inst.leak_cycles_2[1] ;
 wire \system_inst.leak_cycles_2[2] ;
 wire \system_inst.leak_cycles_2[3] ;
 wire \system_inst.leak_rate_1[0] ;
 wire \system_inst.leak_rate_1[1] ;
 wire \system_inst.leak_rate_1[2] ;
 wire \system_inst.leak_rate_1[3] ;
 wire \system_inst.leak_rate_1[4] ;
 wire \system_inst.leak_rate_1[5] ;
 wire \system_inst.leak_rate_1[6] ;
 wire \system_inst.leak_rate_1[7] ;
 wire \system_inst.leak_rate_2[0] ;
 wire \system_inst.leak_rate_2[1] ;
 wire \system_inst.leak_rate_2[2] ;
 wire \system_inst.leak_rate_2[3] ;
 wire \system_inst.leak_rate_2[4] ;
 wire \system_inst.leak_rate_2[5] ;
 wire \system_inst.leak_rate_2[6] ;
 wire \system_inst.leak_rate_2[7] ;
 wire \system_inst.loader.bit_count[0] ;
 wire \system_inst.loader.bit_count[1] ;
 wire \system_inst.loader.bit_count[2] ;
 wire \system_inst.loader.current_state[0] ;
 wire \system_inst.loader.current_state[1] ;
 wire \system_inst.loader.current_state[2] ;
 wire \system_inst.loader.current_state[3] ;
 wire \system_inst.loader.current_state[4] ;
 wire \system_inst.loader.current_state[5] ;
 wire \system_inst.loader.current_state[6] ;
 wire \system_inst.loader.shift_reg[0] ;
 wire \system_inst.loader.shift_reg[1] ;
 wire \system_inst.loader.shift_reg[2] ;
 wire \system_inst.loader.shift_reg[3] ;
 wire \system_inst.loader.shift_reg[4] ;
 wire \system_inst.loader.shift_reg[5] ;
 wire \system_inst.loader.shift_reg[6] ;
 wire \system_inst.loader.threshold_min[0] ;
 wire \system_inst.loader.threshold_min[1] ;
 wire \system_inst.loader.threshold_min[2] ;
 wire \system_inst.loader.threshold_min[3] ;
 wire \system_inst.loader.threshold_min[4] ;
 wire \system_inst.loader.threshold_min[5] ;
 wire \system_inst.loader.threshold_min[6] ;
 wire \system_inst.loader.threshold_min[7] ;
 wire \system_inst.loader.weight_a[0] ;
 wire \system_inst.loader.weight_a[1] ;
 wire \system_inst.loader.weight_a[2] ;
 wire \system_inst.neuron.leak_counter_1[0] ;
 wire \system_inst.neuron.leak_counter_1[1] ;
 wire \system_inst.neuron.leak_counter_1[2] ;
 wire \system_inst.neuron.leak_counter_1[3] ;
 wire \system_inst.neuron.leak_counter_2[0] ;
 wire \system_inst.neuron.leak_counter_2[1] ;
 wire \system_inst.neuron.leak_counter_2[2] ;
 wire \system_inst.neuron.leak_counter_2[3] ;
 wire \system_inst.neuron.refr_cnt[0] ;
 wire \system_inst.neuron.refr_cnt[1] ;
 wire \system_inst.neuron.refr_cnt[2] ;
 wire \system_inst.neuron.refr_cnt[3] ;
 wire \system_inst.neuron.threshold[0] ;
 wire \system_inst.neuron.threshold[1] ;
 wire \system_inst.neuron.threshold[2] ;
 wire \system_inst.neuron.threshold[3] ;
 wire \system_inst.neuron.threshold[4] ;
 wire \system_inst.neuron.threshold[5] ;
 wire \system_inst.neuron.threshold[6] ;
 wire \system_inst.neuron.threshold[7] ;
 wire \system_inst.neuron.v_mem[0] ;
 wire \system_inst.neuron.v_mem[1] ;
 wire \system_inst.neuron.v_mem[2] ;
 wire \system_inst.neuron.v_mem[3] ;
 wire \system_inst.neuron.v_mem[4] ;
 wire \system_inst.neuron.v_mem[5] ;
 wire \system_inst.neuron.v_mem[6] ;
 wire \system_inst.neuron.v_mem[7] ;
 wire \system_inst.neuron.v_mem[8] ;
 wire clknet_0_clk;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;

 sg13g2_inv_1 _0979_ (.Y(_0139_),
    .A(\system_inst.neuron.leak_counter_1[2] ));
 sg13g2_inv_1 _0980_ (.Y(_0140_),
    .A(net254));
 sg13g2_inv_2 _0981_ (.Y(_0141_),
    .A(net139));
 sg13g2_inv_2 _0982_ (.Y(_0142_),
    .A(net204));
 sg13g2_inv_1 _0983_ (.Y(_0143_),
    .A(net226));
 sg13g2_inv_2 _0984_ (.Y(_0144_),
    .A(\system_inst.loader.shift_reg[2] ));
 sg13g2_inv_4 _0985_ (.A(net239),
    .Y(_0145_));
 sg13g2_inv_4 _0986_ (.A(net250),
    .Y(_0146_));
 sg13g2_inv_1 _0987_ (.Y(_0147_),
    .A(\system_inst.leak_cycles_2[3] ));
 sg13g2_inv_1 _0988_ (.Y(_0148_),
    .A(net135));
 sg13g2_inv_4 _0989_ (.A(net4),
    .Y(_0149_));
 sg13g2_inv_1 _0990_ (.Y(_0150_),
    .A(net128));
 sg13g2_inv_1 _0991_ (.Y(_0151_),
    .A(\system_inst.loader.threshold_min[5] ));
 sg13g2_inv_1 _0992_ (.Y(_0152_),
    .A(net230));
 sg13g2_inv_1 _0993_ (.Y(_0153_),
    .A(net246));
 sg13g2_inv_1 _0994_ (.Y(_0154_),
    .A(net264));
 sg13g2_inv_1 _0995_ (.Y(_0155_),
    .A(net194));
 sg13g2_inv_1 _0996_ (.Y(_0156_),
    .A(net261));
 sg13g2_inv_1 _0997_ (.Y(_0157_),
    .A(\system_inst.neuron.leak_counter_2[2] ));
 sg13g2_inv_1 _0998_ (.Y(_0158_),
    .A(\system_inst.neuron.leak_counter_2[1] ));
 sg13g2_inv_1 _0999_ (.Y(_0159_),
    .A(\system_inst.neuron.threshold[7] ));
 sg13g2_inv_2 _1000_ (.Y(_0160_),
    .A(net244));
 sg13g2_inv_2 _1001_ (.Y(_0161_),
    .A(_0010_));
 sg13g2_inv_1 _1002_ (.Y(_0162_),
    .A(net253));
 sg13g2_inv_2 _1003_ (.Y(_0163_),
    .A(_0011_));
 sg13g2_inv_2 _1004_ (.Y(_0164_),
    .A(net252));
 sg13g2_inv_1 _1005_ (.Y(_0165_),
    .A(\system_inst.neuron.threshold[3] ));
 sg13g2_inv_1 _1006_ (.Y(_0166_),
    .A(_0012_));
 sg13g2_inv_2 _1007_ (.Y(_0167_),
    .A(net176));
 sg13g2_inv_1 _1008_ (.Y(_0168_),
    .A(_0013_));
 sg13g2_inv_2 _1009_ (.Y(_0169_),
    .A(\system_inst.neuron.threshold[1] ));
 sg13g2_inv_1 _1010_ (.Y(_0170_),
    .A(_0026_));
 sg13g2_inv_1 _1011_ (.Y(_0171_),
    .A(\system_inst.neuron.threshold[0] ));
 sg13g2_inv_1 _1012_ (.Y(_0172_),
    .A(net192));
 sg13g2_inv_1 _1013_ (.Y(_0173_),
    .A(\system_inst.loader.current_state[0] ));
 sg13g2_inv_1 _1014_ (.Y(_0174_),
    .A(net133));
 sg13g2_inv_1 _1015_ (.Y(_0175_),
    .A(_0033_));
 sg13g2_and2_1 _1016_ (.A(net1),
    .B(net3),
    .X(_0176_));
 sg13g2_nand2_1 _1017_ (.Y(_0177_),
    .A(net191),
    .B(_0176_));
 sg13g2_nand2b_1 _1018_ (.Y(_0178_),
    .B(net191),
    .A_N(net1));
 sg13g2_nor2_1 _1019_ (.A(net132),
    .B(_0178_),
    .Y(_0179_));
 sg13g2_a21oi_1 _1020_ (.A1(net191),
    .A2(net178),
    .Y(_0000_),
    .B1(_0179_));
 sg13g2_nand2_1 _1021_ (.Y(_0180_),
    .A(net124),
    .B(net120));
 sg13g2_nor2_2 _1022_ (.A(_0030_),
    .B(_0180_),
    .Y(_0181_));
 sg13g2_o21ai_1 _1023_ (.B1(_0178_),
    .Y(_0182_),
    .A1(_0177_),
    .A2(_0181_));
 sg13g2_nand3_1 _1024_ (.B(net178),
    .C(net172),
    .A(net118),
    .Y(_0183_));
 sg13g2_inv_1 _1025_ (.Y(_0184_),
    .A(_0183_));
 sg13g2_a22oi_1 _1026_ (.Y(_0185_),
    .B1(_0184_),
    .B2(net192),
    .A2(_0182_),
    .A1(net127));
 sg13g2_inv_1 _1027_ (.Y(_0002_),
    .A(_0185_));
 sg13g2_and3_1 _1028_ (.X(_0186_),
    .A(\system_inst.loader.current_state[5] ),
    .B(net178),
    .C(net172));
 sg13g2_a22oi_1 _1029_ (.Y(_0187_),
    .B1(_0186_),
    .B2(net191),
    .A2(_0182_),
    .A1(net133));
 sg13g2_inv_1 _1030_ (.Y(_0003_),
    .A(net134));
 sg13g2_nand2_1 _1031_ (.Y(_0188_),
    .A(net118),
    .B(_0182_));
 sg13g2_o21ai_1 _1032_ (.B1(_0188_),
    .Y(_0004_),
    .A1(_0173_),
    .A2(_0177_));
 sg13g2_and3_2 _1033_ (.X(_0189_),
    .A(\system_inst.loader.current_state[1] ),
    .B(net178),
    .C(net172));
 sg13g2_nand3_1 _1034_ (.B(net178),
    .C(net172),
    .A(net202),
    .Y(_0190_));
 sg13g2_a22oi_1 _1035_ (.Y(_0191_),
    .B1(_0189_),
    .B2(net191),
    .A2(_0182_),
    .A1(net137));
 sg13g2_inv_1 _1036_ (.Y(_0005_),
    .A(net138));
 sg13g2_and3_1 _1037_ (.X(_0192_),
    .A(net127),
    .B(net178),
    .C(net172));
 sg13g2_a22oi_1 _1038_ (.Y(_0193_),
    .B1(net168),
    .B2(net191),
    .A2(_0182_),
    .A1(net130));
 sg13g2_inv_1 _1039_ (.Y(_0006_),
    .A(_0193_));
 sg13g2_and3_1 _1040_ (.X(_0194_),
    .A(\system_inst.loader.current_state[6] ),
    .B(net178),
    .C(net172));
 sg13g2_a22oi_1 _1041_ (.Y(_0195_),
    .B1(net166),
    .B2(net191),
    .A2(_0182_),
    .A1(net202));
 sg13g2_inv_1 _1042_ (.Y(_0001_),
    .A(_0195_));
 sg13g2_nor2b_1 _1043_ (.A(net177),
    .B_N(\system_inst.neuron.v_mem[0] ),
    .Y(uo_out[1]));
 sg13g2_nor2b_1 _1044_ (.A(net177),
    .B_N(\system_inst.neuron.v_mem[1] ),
    .Y(uo_out[2]));
 sg13g2_nor2b_1 _1045_ (.A(net177),
    .B_N(\system_inst.neuron.v_mem[2] ),
    .Y(uo_out[3]));
 sg13g2_nor2b_1 _1046_ (.A(net177),
    .B_N(\system_inst.neuron.v_mem[3] ),
    .Y(uo_out[4]));
 sg13g2_nor2b_1 _1047_ (.A(net177),
    .B_N(\system_inst.neuron.v_mem[4] ),
    .Y(uo_out[5]));
 sg13g2_nor2b_1 _1048_ (.A(net177),
    .B_N(\system_inst.neuron.v_mem[5] ),
    .Y(uo_out[6]));
 sg13g2_nor2b_1 _1049_ (.A(net177),
    .B_N(\system_inst.neuron.v_mem[6] ),
    .Y(uo_out[7]));
 sg13g2_and2_2 _1050_ (.A(net270),
    .B(net1),
    .X(_0196_));
 sg13g2_nand2_2 _1051_ (.Y(_0197_),
    .A(net271),
    .B(net1));
 sg13g2_nor2_1 _1052_ (.A(\system_inst.leak_cycles_2[1] ),
    .B(_0158_),
    .Y(_0198_));
 sg13g2_nand2b_1 _1053_ (.Y(_0199_),
    .B(\system_inst.leak_cycles_2[0] ),
    .A_N(\system_inst.neuron.leak_counter_2[0] ));
 sg13g2_a22oi_1 _1054_ (.Y(_0200_),
    .B1(_0158_),
    .B2(\system_inst.leak_cycles_2[1] ),
    .A2(_0157_),
    .A1(\system_inst.leak_cycles_2[2] ));
 sg13g2_o21ai_1 _1055_ (.B1(_0200_),
    .Y(_0201_),
    .A1(_0198_),
    .A2(_0199_));
 sg13g2_a22oi_1 _1056_ (.Y(_0202_),
    .B1(\system_inst.neuron.leak_counter_2[2] ),
    .B2(_0148_),
    .A2(\system_inst.neuron.leak_counter_2[3] ),
    .A1(_0147_));
 sg13g2_nand2_1 _1057_ (.Y(_0203_),
    .A(_0201_),
    .B(_0202_));
 sg13g2_o21ai_1 _1058_ (.B1(_0203_),
    .Y(_0204_),
    .A1(_0147_),
    .A2(\system_inst.neuron.leak_counter_2[3] ));
 sg13g2_inv_2 _1059_ (.Y(_0205_),
    .A(net159));
 sg13g2_o21ai_1 _1060_ (.B1(net188),
    .Y(_0206_),
    .A1(_0197_),
    .A2(net160));
 sg13g2_xnor2_1 _1061_ (.Y(_0207_),
    .A(net203),
    .B(_0196_));
 sg13g2_nor2_1 _1062_ (.A(_0206_),
    .B(_0207_),
    .Y(_0039_));
 sg13g2_and3_1 _1063_ (.X(_0208_),
    .A(net115),
    .B(net203),
    .C(_0196_));
 sg13g2_a21oi_1 _1064_ (.A1(\system_inst.neuron.leak_counter_2[0] ),
    .A2(_0196_),
    .Y(_0209_),
    .B1(net115));
 sg13g2_nor3_1 _1065_ (.A(_0206_),
    .B(_0208_),
    .C(net116),
    .Y(_0040_));
 sg13g2_nand2_1 _1066_ (.Y(_0210_),
    .A(\system_inst.neuron.leak_counter_2[2] ),
    .B(_0208_));
 sg13g2_xnor2_1 _1067_ (.Y(_0211_),
    .A(net216),
    .B(_0208_));
 sg13g2_nor2_1 _1068_ (.A(_0206_),
    .B(_0211_),
    .Y(_0041_));
 sg13g2_xor2_1 _1069_ (.B(_0210_),
    .A(net213),
    .X(_0212_));
 sg13g2_nor2_1 _1070_ (.A(_0206_),
    .B(net214),
    .Y(_0042_));
 sg13g2_or2_1 _1071_ (.X(_0213_),
    .B(\system_inst.neuron.refr_cnt[0] ),
    .A(\system_inst.neuron.refr_cnt[1] ));
 sg13g2_nor2_1 _1072_ (.A(\system_inst.neuron.refr_cnt[2] ),
    .B(_0213_),
    .Y(_0214_));
 sg13g2_nor3_2 _1073_ (.A(\system_inst.neuron.refr_cnt[3] ),
    .B(\system_inst.neuron.refr_cnt[2] ),
    .C(_0213_),
    .Y(_0215_));
 sg13g2_and2_2 _1074_ (.A(net2),
    .B(_0196_),
    .X(_0216_));
 sg13g2_nand2_1 _1075_ (.Y(_0217_),
    .A(_0215_),
    .B(_0216_));
 sg13g2_a21oi_1 _1076_ (.A1(_0215_),
    .A2(_0216_),
    .Y(_0218_),
    .B1(net181));
 sg13g2_inv_1 _1077_ (.Y(_0219_),
    .A(net163));
 sg13g2_nand2_1 _1078_ (.Y(_0220_),
    .A(net114),
    .B(_0218_));
 sg13g2_nand2b_1 _1079_ (.Y(_0221_),
    .B(\system_inst.leak_cycles_1[3] ),
    .A_N(\system_inst.neuron.leak_counter_1[3] ));
 sg13g2_nand2_1 _1080_ (.Y(_0222_),
    .A(\system_inst.neuron.leak_counter_1[1] ),
    .B(_0150_));
 sg13g2_nor2b_1 _1081_ (.A(\system_inst.neuron.leak_counter_1[0] ),
    .B_N(\system_inst.leak_cycles_1[0] ),
    .Y(_0223_));
 sg13g2_nor2_1 _1082_ (.A(\system_inst.neuron.leak_counter_1[1] ),
    .B(_0150_),
    .Y(_0224_));
 sg13g2_a221oi_1 _1083_ (.B2(_0223_),
    .C1(_0224_),
    .B1(_0222_),
    .A1(_0139_),
    .Y(_0225_),
    .A2(\system_inst.leak_cycles_1[2] ));
 sg13g2_nand2b_1 _1084_ (.Y(_0226_),
    .B(\system_inst.neuron.leak_counter_1[3] ),
    .A_N(\system_inst.leak_cycles_1[3] ));
 sg13g2_o21ai_1 _1085_ (.B1(_0226_),
    .Y(_0227_),
    .A1(_0139_),
    .A2(\system_inst.leak_cycles_1[2] ));
 sg13g2_o21ai_1 _1086_ (.B1(_0221_),
    .Y(_0228_),
    .A1(_0225_),
    .A2(_0227_));
 sg13g2_inv_4 _1087_ (.A(net162),
    .Y(_0229_));
 sg13g2_and3_1 _1088_ (.X(_0230_),
    .A(net174),
    .B(\system_inst.neuron.v_mem[4] ),
    .C(net7));
 sg13g2_nand3_1 _1089_ (.B(\system_inst.neuron.v_mem[4] ),
    .C(net7),
    .A(net174),
    .Y(_0231_));
 sg13g2_nand2_1 _1090_ (.Y(_0232_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net8));
 sg13g2_a21oi_1 _1091_ (.A1(net174),
    .A2(net7),
    .Y(_0233_),
    .B1(\system_inst.neuron.v_mem[4] ));
 sg13g2_nor2_1 _1092_ (.A(_0230_),
    .B(_0233_),
    .Y(_0234_));
 sg13g2_o21ai_1 _1093_ (.B1(_0231_),
    .Y(_0235_),
    .A1(_0232_),
    .A2(_0233_));
 sg13g2_nand2_1 _1094_ (.Y(_0236_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net9));
 sg13g2_nand3_1 _1095_ (.B(\system_inst.neuron.v_mem[5] ),
    .C(net8),
    .A(net174),
    .Y(_0237_));
 sg13g2_a21o_1 _1096_ (.A2(net8),
    .A1(net174),
    .B1(\system_inst.neuron.v_mem[5] ),
    .X(_0238_));
 sg13g2_nand2_1 _1097_ (.Y(_0239_),
    .A(_0237_),
    .B(_0238_));
 sg13g2_xor2_1 _1098_ (.B(_0239_),
    .A(_0236_),
    .X(_0240_));
 sg13g2_nand2_1 _1099_ (.Y(_0241_),
    .A(_0235_),
    .B(_0240_));
 sg13g2_nand2_1 _1100_ (.Y(_0242_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net10));
 sg13g2_xnor2_1 _1101_ (.Y(_0243_),
    .A(_0235_),
    .B(_0240_));
 sg13g2_or2_1 _1102_ (.X(_0244_),
    .B(_0243_),
    .A(_0242_));
 sg13g2_o21ai_1 _1103_ (.B1(_0237_),
    .Y(_0245_),
    .A1(_0236_),
    .A2(_0239_));
 sg13g2_nand2_1 _1104_ (.Y(_0246_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net10));
 sg13g2_nand3_1 _1105_ (.B(\system_inst.neuron.v_mem[6] ),
    .C(net9),
    .A(net174),
    .Y(_0247_));
 sg13g2_a21o_1 _1106_ (.A2(net9),
    .A1(net174),
    .B1(\system_inst.neuron.v_mem[6] ),
    .X(_0248_));
 sg13g2_nand2_1 _1107_ (.Y(_0249_),
    .A(_0247_),
    .B(_0248_));
 sg13g2_xor2_1 _1108_ (.B(_0249_),
    .A(_0246_),
    .X(_0250_));
 sg13g2_nand2_1 _1109_ (.Y(_0251_),
    .A(_0245_),
    .B(_0250_));
 sg13g2_xnor2_1 _1110_ (.Y(_0252_),
    .A(_0245_),
    .B(_0250_));
 sg13g2_a21oi_1 _1111_ (.A1(_0241_),
    .A2(_0244_),
    .Y(_0253_),
    .B1(_0252_));
 sg13g2_nand3_1 _1112_ (.B(_0244_),
    .C(_0252_),
    .A(_0241_),
    .Y(_0254_));
 sg13g2_nand2b_1 _1113_ (.Y(_0255_),
    .B(_0254_),
    .A_N(_0253_));
 sg13g2_and3_1 _1114_ (.X(_0256_),
    .A(net175),
    .B(\system_inst.neuron.v_mem[3] ),
    .C(net6));
 sg13g2_nand3_1 _1115_ (.B(\system_inst.neuron.v_mem[3] ),
    .C(net6),
    .A(net175),
    .Y(_0257_));
 sg13g2_nand2_1 _1116_ (.Y(_0258_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net7));
 sg13g2_a21oi_1 _1117_ (.A1(net175),
    .A2(net6),
    .Y(_0259_),
    .B1(\system_inst.neuron.v_mem[3] ));
 sg13g2_nor2_1 _1118_ (.A(_0256_),
    .B(_0259_),
    .Y(_0260_));
 sg13g2_o21ai_1 _1119_ (.B1(_0257_),
    .Y(_0261_),
    .A1(_0258_),
    .A2(_0259_));
 sg13g2_xnor2_1 _1120_ (.Y(_0262_),
    .A(_0232_),
    .B(_0234_));
 sg13g2_nand2_1 _1121_ (.Y(_0263_),
    .A(_0261_),
    .B(_0262_));
 sg13g2_nand2_1 _1122_ (.Y(_0264_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net9));
 sg13g2_xnor2_1 _1123_ (.Y(_0265_),
    .A(_0261_),
    .B(_0262_));
 sg13g2_o21ai_1 _1124_ (.B1(_0263_),
    .Y(_0266_),
    .A1(_0264_),
    .A2(_0265_));
 sg13g2_inv_1 _1125_ (.Y(_0267_),
    .A(_0266_));
 sg13g2_xor2_1 _1126_ (.B(_0243_),
    .A(_0242_),
    .X(_0268_));
 sg13g2_inv_1 _1127_ (.Y(_0269_),
    .A(_0268_));
 sg13g2_nor2_1 _1128_ (.A(_0266_),
    .B(_0268_),
    .Y(_0270_));
 sg13g2_and3_1 _1129_ (.X(_0271_),
    .A(net175),
    .B(\system_inst.neuron.v_mem[2] ),
    .C(net5));
 sg13g2_nand2_1 _1130_ (.Y(_0272_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(net6));
 sg13g2_a21oi_1 _1131_ (.A1(net175),
    .A2(net5),
    .Y(_0273_),
    .B1(\system_inst.neuron.v_mem[2] ));
 sg13g2_or3_1 _1132_ (.A(_0271_),
    .B(_0272_),
    .C(_0273_),
    .X(_0274_));
 sg13g2_nand2b_1 _1133_ (.Y(_0275_),
    .B(_0274_),
    .A_N(_0271_));
 sg13g2_xnor2_1 _1134_ (.Y(_0276_),
    .A(_0258_),
    .B(_0260_));
 sg13g2_nand2_1 _1135_ (.Y(_0277_),
    .A(_0275_),
    .B(_0276_));
 sg13g2_nand2_1 _1136_ (.Y(_0278_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net8));
 sg13g2_xnor2_1 _1137_ (.Y(_0279_),
    .A(_0275_),
    .B(_0276_));
 sg13g2_o21ai_1 _1138_ (.B1(_0277_),
    .Y(_0280_),
    .A1(_0278_),
    .A2(_0279_));
 sg13g2_xor2_1 _1139_ (.B(_0265_),
    .A(_0264_),
    .X(_0281_));
 sg13g2_nand2_1 _1140_ (.Y(_0282_),
    .A(_0280_),
    .B(_0281_));
 sg13g2_xor2_1 _1141_ (.B(_0281_),
    .A(_0280_),
    .X(_0283_));
 sg13g2_nand2_1 _1142_ (.Y(_0284_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net5));
 sg13g2_or2_1 _1143_ (.X(_0285_),
    .B(_0284_),
    .A(_0008_));
 sg13g2_and3_1 _1144_ (.X(_0286_),
    .A(\system_inst.loader.weight_a[1] ),
    .B(\system_inst.neuron.v_mem[1] ),
    .C(net5));
 sg13g2_a21oi_1 _1145_ (.A1(\system_inst.loader.weight_a[1] ),
    .A2(net5),
    .Y(_0287_),
    .B1(\system_inst.neuron.v_mem[1] ));
 sg13g2_nand2_1 _1146_ (.Y(_0288_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net6));
 sg13g2_nor3_2 _1147_ (.A(_0286_),
    .B(_0287_),
    .C(_0288_),
    .Y(_0289_));
 sg13g2_o21ai_1 _1148_ (.B1(_0288_),
    .Y(_0290_),
    .A1(_0286_),
    .A2(_0287_));
 sg13g2_nor2b_2 _1149_ (.A(_0289_),
    .B_N(_0290_),
    .Y(_0291_));
 sg13g2_nor2b_1 _1150_ (.A(_0285_),
    .B_N(_0291_),
    .Y(_0292_));
 sg13g2_nand2_1 _1151_ (.Y(_0293_),
    .A(\system_inst.loader.weight_a[0] ),
    .B(net7));
 sg13g2_o21ai_1 _1152_ (.B1(_0272_),
    .Y(_0294_),
    .A1(_0271_),
    .A2(_0273_));
 sg13g2_and3_1 _1153_ (.X(_0295_),
    .A(_0274_),
    .B(_0286_),
    .C(_0294_));
 sg13g2_a21oi_1 _1154_ (.A1(_0274_),
    .A2(_0294_),
    .Y(_0296_),
    .B1(_0286_));
 sg13g2_or3_1 _1155_ (.A(_0293_),
    .B(_0295_),
    .C(_0296_),
    .X(_0297_));
 sg13g2_o21ai_1 _1156_ (.B1(_0293_),
    .Y(_0298_),
    .A1(_0295_),
    .A2(_0296_));
 sg13g2_and3_1 _1157_ (.X(_0299_),
    .A(_0289_),
    .B(_0297_),
    .C(_0298_));
 sg13g2_a21o_1 _1158_ (.A2(_0298_),
    .A1(_0297_),
    .B1(_0289_),
    .X(_0300_));
 sg13g2_nand2b_1 _1159_ (.Y(_0301_),
    .B(_0300_),
    .A_N(_0299_));
 sg13g2_nand2b_1 _1160_ (.Y(_0302_),
    .B(_0297_),
    .A_N(_0295_));
 sg13g2_xor2_1 _1161_ (.B(_0279_),
    .A(_0278_),
    .X(_0303_));
 sg13g2_a221oi_1 _1162_ (.B2(_0303_),
    .C1(_0299_),
    .B1(_0302_),
    .A1(_0292_),
    .Y(_0304_),
    .A2(_0300_));
 sg13g2_or2_1 _1163_ (.X(_0305_),
    .B(_0303_),
    .A(_0302_));
 sg13g2_nand2b_1 _1164_ (.Y(_0306_),
    .B(_0305_),
    .A_N(_0304_));
 sg13g2_nand3b_1 _1165_ (.B(_0305_),
    .C(_0283_),
    .Y(_0307_),
    .A_N(_0304_));
 sg13g2_nand2_1 _1166_ (.Y(_0308_),
    .A(_0266_),
    .B(_0268_));
 sg13g2_and2_1 _1167_ (.A(_0282_),
    .B(_0308_),
    .X(_0309_));
 sg13g2_a21oi_1 _1168_ (.A1(_0307_),
    .A2(_0309_),
    .Y(_0310_),
    .B1(_0270_));
 sg13g2_a221oi_1 _1169_ (.B2(_0309_),
    .C1(_0255_),
    .B1(_0307_),
    .A1(_0267_),
    .Y(_0311_),
    .A2(_0269_));
 sg13g2_o21ai_1 _1170_ (.B1(_0247_),
    .Y(_0312_),
    .A1(_0246_),
    .A2(_0249_));
 sg13g2_nand2_1 _1171_ (.Y(_0313_),
    .A(net174),
    .B(net10));
 sg13g2_nor2_1 _1172_ (.A(_0007_),
    .B(_0313_),
    .Y(_0314_));
 sg13g2_nand2_1 _1173_ (.Y(_0315_),
    .A(_0007_),
    .B(_0313_));
 sg13g2_nor2b_1 _1174_ (.A(_0314_),
    .B_N(_0315_),
    .Y(_0316_));
 sg13g2_xnor2_1 _1175_ (.Y(_0317_),
    .A(_0312_),
    .B(_0316_));
 sg13g2_xor2_1 _1176_ (.B(_0317_),
    .A(_0251_),
    .X(_0318_));
 sg13g2_o21ai_1 _1177_ (.B1(_0318_),
    .Y(_0319_),
    .A1(_0253_),
    .A2(_0311_));
 sg13g2_or3_1 _1178_ (.A(_0253_),
    .B(_0311_),
    .C(_0318_),
    .X(_0320_));
 sg13g2_and2_2 _1179_ (.A(_0319_),
    .B(_0320_),
    .X(_0321_));
 sg13g2_and2_1 _1180_ (.A(net161),
    .B(_0321_),
    .X(_0322_));
 sg13g2_xnor2_1 _1181_ (.Y(_0323_),
    .A(_0255_),
    .B(_0310_));
 sg13g2_xnor2_1 _1182_ (.Y(_0324_),
    .A(_0009_),
    .B(_0323_));
 sg13g2_nand2b_1 _1183_ (.Y(_0325_),
    .B(_0308_),
    .A_N(_0270_));
 sg13g2_nand3_1 _1184_ (.B(_0307_),
    .C(_0325_),
    .A(_0282_),
    .Y(_0326_));
 sg13g2_a21o_2 _1185_ (.A2(_0307_),
    .A1(_0282_),
    .B1(_0325_),
    .X(_0327_));
 sg13g2_nand2_2 _1186_ (.Y(_0328_),
    .A(_0326_),
    .B(_0327_));
 sg13g2_and2_1 _1187_ (.A(_0326_),
    .B(_0327_),
    .X(_0329_));
 sg13g2_a21oi_1 _1188_ (.A1(_0326_),
    .A2(_0327_),
    .Y(_0330_),
    .B1(_0010_));
 sg13g2_xor2_1 _1189_ (.B(_0306_),
    .A(_0283_),
    .X(_0331_));
 sg13g2_a21oi_1 _1190_ (.A1(_0163_),
    .A2(_0331_),
    .Y(_0332_),
    .B1(_0330_));
 sg13g2_nor2_1 _1191_ (.A(_0161_),
    .B(_0328_),
    .Y(_0333_));
 sg13g2_nand3_1 _1192_ (.B(_0326_),
    .C(_0327_),
    .A(_0010_),
    .Y(_0334_));
 sg13g2_xnor2_1 _1193_ (.Y(_0335_),
    .A(_0011_),
    .B(_0331_));
 sg13g2_nand3b_1 _1194_ (.B(_0334_),
    .C(_0335_),
    .Y(_0336_),
    .A_N(_0330_));
 sg13g2_nor3_1 _1195_ (.A(_0321_),
    .B(_0324_),
    .C(_0336_),
    .Y(_0337_));
 sg13g2_a21oi_1 _1196_ (.A1(_0292_),
    .A2(_0300_),
    .Y(_0338_),
    .B1(_0299_));
 sg13g2_xnor2_1 _1197_ (.Y(_0339_),
    .A(_0302_),
    .B(_0303_));
 sg13g2_xnor2_1 _1198_ (.Y(_0340_),
    .A(_0338_),
    .B(_0339_));
 sg13g2_inv_1 _1199_ (.Y(_0341_),
    .A(_0340_));
 sg13g2_or2_1 _1200_ (.X(_0342_),
    .B(_0340_),
    .A(\system_inst.neuron.threshold[4] ));
 sg13g2_xor2_1 _1201_ (.B(_0301_),
    .A(_0292_),
    .X(_0343_));
 sg13g2_inv_1 _1202_ (.Y(_0344_),
    .A(_0343_));
 sg13g2_xnor2_1 _1203_ (.Y(_0345_),
    .A(_0012_),
    .B(_0343_));
 sg13g2_nand2_1 _1204_ (.Y(_0346_),
    .A(\system_inst.neuron.threshold[4] ),
    .B(_0340_));
 sg13g2_and3_1 _1205_ (.X(_0347_),
    .A(_0342_),
    .B(_0345_),
    .C(_0346_));
 sg13g2_xnor2_1 _1206_ (.Y(_0348_),
    .A(_0285_),
    .B(_0291_));
 sg13g2_xor2_1 _1207_ (.B(_0291_),
    .A(_0285_),
    .X(_0349_));
 sg13g2_xor2_1 _1208_ (.B(_0284_),
    .A(_0008_),
    .X(_0350_));
 sg13g2_xnor2_1 _1209_ (.Y(_0351_),
    .A(_0013_),
    .B(_0348_));
 sg13g2_a21oi_1 _1210_ (.A1(_0169_),
    .A2(_0350_),
    .Y(_0352_),
    .B1(_0351_));
 sg13g2_a21o_1 _1211_ (.A2(_0349_),
    .A1(\system_inst.neuron.threshold[2] ),
    .B1(_0352_),
    .X(_0353_));
 sg13g2_o21ai_1 _1212_ (.B1(_0346_),
    .Y(_0354_),
    .A1(_0165_),
    .A2(_0344_));
 sg13g2_a22oi_1 _1213_ (.Y(_0355_),
    .B1(_0354_),
    .B2(_0342_),
    .A2(_0353_),
    .A1(_0347_));
 sg13g2_nor4_2 _1214_ (.A(_0321_),
    .B(_0324_),
    .C(_0336_),
    .Y(_0356_),
    .D(_0355_));
 sg13g2_nor4_2 _1215_ (.A(_0321_),
    .B(_0324_),
    .C(_0332_),
    .Y(_0357_),
    .D(_0333_));
 sg13g2_nor3_1 _1216_ (.A(_0159_),
    .B(_0321_),
    .C(_0323_),
    .Y(_0358_));
 sg13g2_nor3_2 _1217_ (.A(_0356_),
    .B(_0357_),
    .C(_0358_),
    .Y(_0359_));
 sg13g2_or3_2 _1218_ (.A(_0356_),
    .B(_0357_),
    .C(_0358_),
    .X(_0360_));
 sg13g2_xnor2_1 _1219_ (.Y(_0361_),
    .A(_0014_),
    .B(_0350_));
 sg13g2_nor2_1 _1220_ (.A(_0351_),
    .B(_0361_),
    .Y(_0362_));
 sg13g2_and2_1 _1221_ (.A(_0347_),
    .B(_0362_),
    .X(_0363_));
 sg13g2_o21ai_1 _1222_ (.B1(_0319_),
    .Y(_0364_),
    .A1(_0251_),
    .A2(_0317_));
 sg13g2_a21oi_1 _1223_ (.A1(_0312_),
    .A2(_0315_),
    .Y(_0365_),
    .B1(_0314_));
 sg13g2_xor2_1 _1224_ (.B(_0365_),
    .A(\system_inst.neuron.v_mem[8] ),
    .X(_0366_));
 sg13g2_xnor2_1 _1225_ (.Y(_0367_),
    .A(_0364_),
    .B(_0366_));
 sg13g2_a21oi_2 _1226_ (.B1(_0367_),
    .Y(_0368_),
    .A2(_0363_),
    .A1(_0337_));
 sg13g2_a21o_1 _1227_ (.A2(_0363_),
    .A1(_0337_),
    .B1(_0367_),
    .X(_0369_));
 sg13g2_nor2_2 _1228_ (.A(_0359_),
    .B(_0369_),
    .Y(_0370_));
 sg13g2_nor2_1 _1229_ (.A(\system_inst.leak_rate_1[1] ),
    .B(\system_inst.leak_rate_1[0] ),
    .Y(_0371_));
 sg13g2_nor3_1 _1230_ (.A(\system_inst.leak_rate_1[2] ),
    .B(\system_inst.leak_rate_1[1] ),
    .C(\system_inst.leak_rate_1[0] ),
    .Y(_0372_));
 sg13g2_nor2b_1 _1231_ (.A(\system_inst.leak_rate_1[3] ),
    .B_N(_0372_),
    .Y(_0373_));
 sg13g2_nor2b_1 _1232_ (.A(\system_inst.leak_rate_1[4] ),
    .B_N(_0373_),
    .Y(_0374_));
 sg13g2_nor2b_1 _1233_ (.A(\system_inst.leak_rate_1[5] ),
    .B_N(_0374_),
    .Y(_0375_));
 sg13g2_nand2b_1 _1234_ (.Y(_0376_),
    .B(_0375_),
    .A_N(\system_inst.leak_rate_1[6] ));
 sg13g2_nor2_1 _1235_ (.A(\system_inst.leak_rate_1[7] ),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_nor3_1 _1236_ (.A(_0359_),
    .B(_0369_),
    .C(_0377_),
    .Y(_0378_));
 sg13g2_nand2_1 _1237_ (.Y(_0379_),
    .A(\system_inst.leak_rate_1[7] ),
    .B(_0376_));
 sg13g2_nor2_1 _1238_ (.A(_0015_),
    .B(_0370_),
    .Y(_0380_));
 sg13g2_a21oi_1 _1239_ (.A1(_0378_),
    .A2(_0379_),
    .Y(_0381_),
    .B1(_0380_));
 sg13g2_nand2_1 _1240_ (.Y(_0382_),
    .A(_0321_),
    .B(_0381_));
 sg13g2_xnor2_1 _1241_ (.Y(_0383_),
    .A(_0321_),
    .B(_0381_));
 sg13g2_inv_1 _1242_ (.Y(_0384_),
    .A(_0383_));
 sg13g2_xnor2_1 _1243_ (.Y(_0385_),
    .A(\system_inst.leak_rate_1[6] ),
    .B(_0375_));
 sg13g2_nor2_1 _1244_ (.A(_0016_),
    .B(_0370_),
    .Y(_0386_));
 sg13g2_a21oi_1 _1245_ (.A1(_0370_),
    .A2(_0385_),
    .Y(_0387_),
    .B1(_0386_));
 sg13g2_nand2_1 _1246_ (.Y(_0388_),
    .A(_0323_),
    .B(_0387_));
 sg13g2_xnor2_1 _1247_ (.Y(_0389_),
    .A(_0323_),
    .B(_0387_));
 sg13g2_xnor2_1 _1248_ (.Y(_0390_),
    .A(\system_inst.leak_rate_1[3] ),
    .B(_0372_));
 sg13g2_a21o_1 _1249_ (.A2(_0368_),
    .A1(_0360_),
    .B1(_0019_),
    .X(_0391_));
 sg13g2_nand3_1 _1250_ (.B(_0368_),
    .C(_0390_),
    .A(_0360_),
    .Y(_0392_));
 sg13g2_a21oi_1 _1251_ (.A1(_0391_),
    .A2(_0392_),
    .Y(_0393_),
    .B1(_0341_));
 sg13g2_a21o_1 _1252_ (.A2(_0392_),
    .A1(_0391_),
    .B1(_0341_),
    .X(_0394_));
 sg13g2_xnor2_1 _1253_ (.Y(_0395_),
    .A(\system_inst.leak_rate_1[2] ),
    .B(_0371_));
 sg13g2_a21o_1 _1254_ (.A2(_0368_),
    .A1(_0360_),
    .B1(_0020_),
    .X(_0396_));
 sg13g2_nand3_1 _1255_ (.B(_0368_),
    .C(_0395_),
    .A(_0360_),
    .Y(_0397_));
 sg13g2_nand3_1 _1256_ (.B(_0396_),
    .C(_0397_),
    .A(_0344_),
    .Y(_0398_));
 sg13g2_nand3_1 _1257_ (.B(_0391_),
    .C(_0392_),
    .A(_0341_),
    .Y(_0399_));
 sg13g2_and2_1 _1258_ (.A(\system_inst.leak_rate_1[1] ),
    .B(\system_inst.leak_rate_1[0] ),
    .X(_0400_));
 sg13g2_a21oi_1 _1259_ (.A1(_0360_),
    .A2(_0368_),
    .Y(_0401_),
    .B1(_0021_));
 sg13g2_nor4_2 _1260_ (.A(_0359_),
    .B(_0369_),
    .C(_0371_),
    .Y(_0402_),
    .D(_0400_));
 sg13g2_nor3_1 _1261_ (.A(_0349_),
    .B(_0401_),
    .C(_0402_),
    .Y(_0403_));
 sg13g2_or3_1 _1262_ (.A(_0349_),
    .B(_0401_),
    .C(_0402_),
    .X(_0404_));
 sg13g2_nand2b_1 _1263_ (.Y(_0405_),
    .B(\system_inst.leak_rate_1[0] ),
    .A_N(_0350_));
 sg13g2_o21ai_1 _1264_ (.B1(_0349_),
    .Y(_0406_),
    .A1(_0401_),
    .A2(_0402_));
 sg13g2_nand3_1 _1265_ (.B(_0405_),
    .C(_0406_),
    .A(_0404_),
    .Y(_0407_));
 sg13g2_a21oi_2 _1266_ (.B1(_0403_),
    .Y(_0408_),
    .A2(_0406_),
    .A1(_0405_));
 sg13g2_a21o_1 _1267_ (.A2(_0397_),
    .A1(_0396_),
    .B1(_0344_),
    .X(_0409_));
 sg13g2_nand2_1 _1268_ (.Y(_0410_),
    .A(_0398_),
    .B(_0409_));
 sg13g2_nand2_1 _1269_ (.Y(_0411_),
    .A(_0394_),
    .B(_0399_));
 sg13g2_nand4_1 _1270_ (.B(_0398_),
    .C(_0399_),
    .A(_0394_),
    .Y(_0412_),
    .D(_0409_));
 sg13g2_a21o_1 _1271_ (.A2(_0399_),
    .A1(_0398_),
    .B1(_0393_),
    .X(_0413_));
 sg13g2_o21ai_1 _1272_ (.B1(_0413_),
    .Y(_0414_),
    .A1(_0408_),
    .A2(_0412_));
 sg13g2_xor2_1 _1273_ (.B(_0373_),
    .A(\system_inst.leak_rate_1[4] ),
    .X(_0415_));
 sg13g2_mux2_1 _1274_ (.A0(_0018_),
    .A1(_0415_),
    .S(_0370_),
    .X(_0416_));
 sg13g2_nor2b_1 _1275_ (.A(_0331_),
    .B_N(_0416_),
    .Y(_0417_));
 sg13g2_xnor2_1 _1276_ (.Y(_0418_),
    .A(_0331_),
    .B(_0416_));
 sg13g2_xnor2_1 _1277_ (.Y(_0419_),
    .A(\system_inst.leak_rate_1[5] ),
    .B(_0374_));
 sg13g2_nand3_1 _1278_ (.B(_0368_),
    .C(_0419_),
    .A(_0360_),
    .Y(_0420_));
 sg13g2_o21ai_1 _1279_ (.B1(_0420_),
    .Y(_0421_),
    .A1(_0017_),
    .A2(_0370_));
 sg13g2_nand2_1 _1280_ (.Y(_0422_),
    .A(_0328_),
    .B(_0421_));
 sg13g2_nor2_1 _1281_ (.A(_0328_),
    .B(_0421_),
    .Y(_0423_));
 sg13g2_xnor2_1 _1282_ (.Y(_0424_),
    .A(_0329_),
    .B(_0421_));
 sg13g2_and2_1 _1283_ (.A(_0418_),
    .B(_0424_),
    .X(_0425_));
 sg13g2_a221oi_1 _1284_ (.B2(_0414_),
    .C1(_0423_),
    .B1(_0425_),
    .A1(_0417_),
    .Y(_0426_),
    .A2(_0422_));
 sg13g2_o21ai_1 _1285_ (.B1(_0388_),
    .Y(_0427_),
    .A1(_0389_),
    .A2(_0426_));
 sg13g2_nand2b_1 _1286_ (.Y(_0428_),
    .B(_0383_),
    .A_N(_0427_));
 sg13g2_a21oi_2 _1287_ (.B1(net161),
    .Y(_0429_),
    .A2(_0427_),
    .A1(_0384_));
 sg13g2_a21oi_2 _1288_ (.B1(_0322_),
    .Y(_0430_),
    .A2(_0429_),
    .A1(_0428_));
 sg13g2_a21o_2 _1289_ (.A2(_0429_),
    .A1(_0428_),
    .B1(_0322_),
    .X(_0431_));
 sg13g2_or3_2 _1290_ (.A(\system_inst.leak_rate_2[2] ),
    .B(\system_inst.leak_rate_2[1] ),
    .C(\system_inst.leak_rate_2[0] ),
    .X(_0432_));
 sg13g2_nor2_1 _1291_ (.A(\system_inst.leak_rate_2[3] ),
    .B(_0432_),
    .Y(_0433_));
 sg13g2_nor3_1 _1292_ (.A(\system_inst.leak_rate_2[4] ),
    .B(\system_inst.leak_rate_2[3] ),
    .C(_0432_),
    .Y(_0434_));
 sg13g2_nor2b_1 _1293_ (.A(\system_inst.leak_rate_2[5] ),
    .B_N(_0434_),
    .Y(_0435_));
 sg13g2_nor2b_1 _1294_ (.A(\system_inst.leak_rate_2[6] ),
    .B_N(_0435_),
    .Y(_0436_));
 sg13g2_nand2b_1 _1295_ (.Y(_0437_),
    .B(\system_inst.leak_rate_2[7] ),
    .A_N(_0436_));
 sg13g2_and2_1 _1296_ (.A(net161),
    .B(_0323_),
    .X(_0438_));
 sg13g2_xor2_1 _1297_ (.B(_0426_),
    .A(_0389_),
    .X(_0439_));
 sg13g2_a21oi_2 _1298_ (.B1(_0438_),
    .Y(_0440_),
    .A2(_0439_),
    .A1(_0229_));
 sg13g2_nand2_1 _1299_ (.Y(_0441_),
    .A(\system_inst.neuron.threshold[7] ),
    .B(_0440_));
 sg13g2_nand2_1 _1300_ (.Y(_0442_),
    .A(net161),
    .B(_0328_));
 sg13g2_a21oi_1 _1301_ (.A1(_0414_),
    .A2(_0418_),
    .Y(_0443_),
    .B1(_0417_));
 sg13g2_xnor2_1 _1302_ (.Y(_0444_),
    .A(_0424_),
    .B(_0443_));
 sg13g2_mux2_2 _1303_ (.A0(_0329_),
    .A1(_0444_),
    .S(_0229_),
    .X(_0445_));
 sg13g2_o21ai_1 _1304_ (.B1(_0442_),
    .Y(_0446_),
    .A1(net161),
    .A2(_0444_));
 sg13g2_nand2_1 _1305_ (.Y(_0447_),
    .A(net161),
    .B(_0331_));
 sg13g2_xor2_1 _1306_ (.B(_0418_),
    .A(_0414_),
    .X(_0448_));
 sg13g2_o21ai_1 _1307_ (.B1(_0447_),
    .Y(_0449_),
    .A1(net161),
    .A2(_0448_));
 sg13g2_nand2_1 _1308_ (.Y(_0450_),
    .A(_0163_),
    .B(_0449_));
 sg13g2_a22oi_1 _1309_ (.Y(_0451_),
    .B1(_0449_),
    .B2(_0163_),
    .A2(_0446_),
    .A1(_0161_));
 sg13g2_o21ai_1 _1310_ (.B1(_0450_),
    .Y(_0452_),
    .A1(_0010_),
    .A2(_0445_));
 sg13g2_nor2_1 _1311_ (.A(_0229_),
    .B(_0340_),
    .Y(_0453_));
 sg13g2_o21ai_1 _1312_ (.B1(_0398_),
    .Y(_0454_),
    .A1(_0408_),
    .A2(_0410_));
 sg13g2_xnor2_1 _1313_ (.Y(_0455_),
    .A(_0411_),
    .B(_0454_));
 sg13g2_a21oi_2 _1314_ (.B1(_0453_),
    .Y(_0456_),
    .A2(_0455_),
    .A1(_0229_));
 sg13g2_a21o_2 _1315_ (.A2(_0455_),
    .A1(_0229_),
    .B1(_0453_),
    .X(_0457_));
 sg13g2_nand2_1 _1316_ (.Y(_0458_),
    .A(net162),
    .B(_0344_));
 sg13g2_xnor2_1 _1317_ (.Y(_0459_),
    .A(_0408_),
    .B(_0410_));
 sg13g2_o21ai_1 _1318_ (.B1(_0458_),
    .Y(_0460_),
    .A1(net162),
    .A2(_0459_));
 sg13g2_xnor2_1 _1319_ (.Y(_0461_),
    .A(_0012_),
    .B(_0460_));
 sg13g2_a21o_1 _1320_ (.A2(_0457_),
    .A1(_0164_),
    .B1(_0461_),
    .X(_0462_));
 sg13g2_and2_1 _1321_ (.A(\system_inst.leak_rate_1[0] ),
    .B(_0229_),
    .X(_0463_));
 sg13g2_xnor2_1 _1322_ (.Y(_0464_),
    .A(_0350_),
    .B(_0463_));
 sg13g2_or2_1 _1323_ (.X(_0465_),
    .B(_0464_),
    .A(\system_inst.neuron.threshold[1] ));
 sg13g2_a21o_1 _1324_ (.A2(_0406_),
    .A1(_0404_),
    .B1(_0405_),
    .X(_0466_));
 sg13g2_nor2_2 _1325_ (.A(_0229_),
    .B(_0348_),
    .Y(_0467_));
 sg13g2_a21oi_2 _1326_ (.B1(net161),
    .Y(_0468_),
    .A2(_0466_),
    .A1(_0407_));
 sg13g2_or2_2 _1327_ (.X(_0469_),
    .B(_0468_),
    .A(_0467_));
 sg13g2_nor2_1 _1328_ (.A(_0467_),
    .B(_0468_),
    .Y(_0470_));
 sg13g2_o21ai_1 _1329_ (.B1(_0168_),
    .Y(_0471_),
    .A1(_0467_),
    .A2(_0468_));
 sg13g2_or3_1 _1330_ (.A(_0168_),
    .B(_0467_),
    .C(_0468_),
    .X(_0472_));
 sg13g2_nand3_1 _1331_ (.B(_0471_),
    .C(_0472_),
    .A(_0465_),
    .Y(_0473_));
 sg13g2_nand2_1 _1332_ (.Y(_0474_),
    .A(\system_inst.neuron.threshold[2] ),
    .B(_0469_));
 sg13g2_a221oi_1 _1333_ (.B2(_0474_),
    .C1(_0461_),
    .B1(_0473_),
    .A1(_0164_),
    .Y(_0475_),
    .A2(_0457_));
 sg13g2_nor2_1 _1334_ (.A(_0164_),
    .B(_0457_),
    .Y(_0476_));
 sg13g2_nand2_1 _1335_ (.Y(_0477_),
    .A(\system_inst.neuron.threshold[4] ),
    .B(_0456_));
 sg13g2_nor2_1 _1336_ (.A(_0165_),
    .B(_0460_),
    .Y(_0478_));
 sg13g2_o21ai_1 _1337_ (.B1(_0478_),
    .Y(_0479_),
    .A1(\system_inst.neuron.threshold[4] ),
    .A2(_0456_));
 sg13g2_nand3b_1 _1338_ (.B(_0477_),
    .C(_0479_),
    .Y(_0480_),
    .A_N(_0475_));
 sg13g2_nor2_1 _1339_ (.A(_0163_),
    .B(_0449_),
    .Y(_0481_));
 sg13g2_inv_1 _1340_ (.Y(_0482_),
    .A(_0481_));
 sg13g2_a21oi_1 _1341_ (.A1(_0480_),
    .A2(_0482_),
    .Y(_0483_),
    .B1(_0452_));
 sg13g2_xor2_1 _1342_ (.B(_0440_),
    .A(_0009_),
    .X(_0484_));
 sg13g2_nor2_1 _1343_ (.A(_0161_),
    .B(_0446_),
    .Y(_0485_));
 sg13g2_or2_1 _1344_ (.X(_0486_),
    .B(_0485_),
    .A(_0484_));
 sg13g2_o21ai_1 _1345_ (.B1(_0441_),
    .Y(_0487_),
    .A1(_0483_),
    .A2(_0486_));
 sg13g2_xnor2_1 _1346_ (.Y(_0488_),
    .A(_0361_),
    .B(_0463_));
 sg13g2_nand3_1 _1347_ (.B(_0472_),
    .C(_0488_),
    .A(_0471_),
    .Y(_0489_));
 sg13g2_or4_1 _1348_ (.A(_0462_),
    .B(_0476_),
    .C(_0481_),
    .D(_0489_),
    .X(_0490_));
 sg13g2_nor4_1 _1349_ (.A(_0452_),
    .B(_0484_),
    .C(_0485_),
    .D(_0490_),
    .Y(_0491_));
 sg13g2_a21oi_1 _1350_ (.A1(_0229_),
    .A2(_0378_),
    .Y(_0492_),
    .B1(_0367_));
 sg13g2_and2_1 _1351_ (.A(_0382_),
    .B(_0429_),
    .X(_0493_));
 sg13g2_xnor2_1 _1352_ (.Y(_0494_),
    .A(_0492_),
    .B(_0493_));
 sg13g2_nor3_2 _1353_ (.A(_0431_),
    .B(_0491_),
    .C(_0494_),
    .Y(_0495_));
 sg13g2_nor2_1 _1354_ (.A(_0431_),
    .B(_0484_),
    .Y(_0496_));
 sg13g2_a21o_1 _1355_ (.A2(_0445_),
    .A1(_0010_),
    .B1(_0481_),
    .X(_0497_));
 sg13g2_nor4_1 _1356_ (.A(_0431_),
    .B(_0452_),
    .C(_0484_),
    .D(_0497_),
    .Y(_0498_));
 sg13g2_nor2_1 _1357_ (.A(_0451_),
    .B(_0485_),
    .Y(_0499_));
 sg13g2_nor2_1 _1358_ (.A(_0431_),
    .B(_0441_),
    .Y(_0500_));
 sg13g2_a221oi_1 _1359_ (.B2(_0496_),
    .C1(_0500_),
    .B1(_0499_),
    .A1(_0480_),
    .Y(_0501_),
    .A2(_0498_));
 sg13g2_nor3_1 _1360_ (.A(_0462_),
    .B(_0476_),
    .C(_0489_),
    .Y(_0502_));
 sg13g2_a21o_1 _1361_ (.A2(_0502_),
    .A1(_0498_),
    .B1(_0494_),
    .X(_0503_));
 sg13g2_nor2_2 _1362_ (.A(_0501_),
    .B(_0503_),
    .Y(_0504_));
 sg13g2_nand2b_1 _1363_ (.Y(_0505_),
    .B(_0436_),
    .A_N(\system_inst.leak_rate_2[7] ));
 sg13g2_and2_1 _1364_ (.A(_0504_),
    .B(_0505_),
    .X(_0506_));
 sg13g2_nor2_1 _1365_ (.A(_0022_),
    .B(_0504_),
    .Y(_0507_));
 sg13g2_a21oi_2 _1366_ (.B1(_0507_),
    .Y(_0508_),
    .A2(_0506_),
    .A1(_0437_));
 sg13g2_xnor2_1 _1367_ (.Y(_0509_),
    .A(_0430_),
    .B(_0508_));
 sg13g2_xnor2_1 _1368_ (.Y(_0510_),
    .A(\system_inst.leak_rate_2[1] ),
    .B(\system_inst.leak_rate_2[0] ));
 sg13g2_a21oi_1 _1369_ (.A1(_0487_),
    .A2(_0495_),
    .Y(_0511_),
    .B1(_0028_));
 sg13g2_a21o_1 _1370_ (.A2(_0495_),
    .A1(_0487_),
    .B1(_0028_),
    .X(_0512_));
 sg13g2_nor3_1 _1371_ (.A(_0501_),
    .B(_0503_),
    .C(_0510_),
    .Y(_0513_));
 sg13g2_or3_1 _1372_ (.A(_0501_),
    .B(_0503_),
    .C(_0510_),
    .X(_0514_));
 sg13g2_nor3_1 _1373_ (.A(_0469_),
    .B(_0511_),
    .C(_0513_),
    .Y(_0515_));
 sg13g2_nand3_1 _1374_ (.B(_0512_),
    .C(_0514_),
    .A(_0470_),
    .Y(_0516_));
 sg13g2_and2_1 _1375_ (.A(\system_inst.leak_rate_2[0] ),
    .B(_0464_),
    .X(_0517_));
 sg13g2_inv_1 _1376_ (.Y(_0518_),
    .A(_0517_));
 sg13g2_a21oi_1 _1377_ (.A1(_0512_),
    .A2(_0514_),
    .Y(_0519_),
    .B1(_0470_));
 sg13g2_o21ai_1 _1378_ (.B1(_0469_),
    .Y(_0520_),
    .A1(_0511_),
    .A2(_0513_));
 sg13g2_nand3_1 _1379_ (.B(_0518_),
    .C(_0520_),
    .A(_0516_),
    .Y(_0521_));
 sg13g2_a21oi_1 _1380_ (.A1(_0518_),
    .A2(_0520_),
    .Y(_0522_),
    .B1(_0515_));
 sg13g2_o21ai_1 _1381_ (.B1(_0516_),
    .Y(_0523_),
    .A1(_0517_),
    .A2(_0519_));
 sg13g2_a21oi_1 _1382_ (.A1(_0487_),
    .A2(_0495_),
    .Y(_0524_),
    .B1(_0026_));
 sg13g2_xnor2_1 _1383_ (.Y(_0525_),
    .A(\system_inst.leak_rate_2[3] ),
    .B(_0432_));
 sg13g2_nor3_1 _1384_ (.A(_0501_),
    .B(_0503_),
    .C(_0525_),
    .Y(_0526_));
 sg13g2_and3_1 _1385_ (.X(_0527_),
    .A(_0487_),
    .B(_0495_),
    .C(_0525_));
 sg13g2_a21oi_1 _1386_ (.A1(_0487_),
    .A2(_0495_),
    .Y(_0528_),
    .B1(_0170_));
 sg13g2_nor3_2 _1387_ (.A(_0457_),
    .B(_0527_),
    .C(_0528_),
    .Y(_0529_));
 sg13g2_nor3_1 _1388_ (.A(_0456_),
    .B(_0524_),
    .C(_0526_),
    .Y(_0530_));
 sg13g2_o21ai_1 _1389_ (.B1(_0457_),
    .Y(_0531_),
    .A1(_0527_),
    .A2(_0528_));
 sg13g2_nor2_1 _1390_ (.A(_0529_),
    .B(_0530_),
    .Y(_0532_));
 sg13g2_o21ai_1 _1391_ (.B1(\system_inst.leak_rate_2[2] ),
    .Y(_0533_),
    .A1(\system_inst.leak_rate_2[1] ),
    .A2(\system_inst.leak_rate_2[0] ));
 sg13g2_a21o_1 _1392_ (.A2(_0495_),
    .A1(_0487_),
    .B1(_0027_),
    .X(_0534_));
 sg13g2_nand4_1 _1393_ (.B(_0487_),
    .C(_0495_),
    .A(_0432_),
    .Y(_0535_),
    .D(_0533_));
 sg13g2_and3_1 _1394_ (.X(_0536_),
    .A(_0460_),
    .B(_0534_),
    .C(_0535_));
 sg13g2_nand3_1 _1395_ (.B(_0534_),
    .C(_0535_),
    .A(_0460_),
    .Y(_0537_));
 sg13g2_a21oi_1 _1396_ (.A1(_0534_),
    .A2(_0535_),
    .Y(_0538_),
    .B1(_0460_));
 sg13g2_nor2_1 _1397_ (.A(_0536_),
    .B(_0538_),
    .Y(_0539_));
 sg13g2_nor4_1 _1398_ (.A(_0529_),
    .B(_0530_),
    .C(_0536_),
    .D(_0538_),
    .Y(_0540_));
 sg13g2_a21oi_1 _1399_ (.A1(_0531_),
    .A2(_0537_),
    .Y(_0541_),
    .B1(_0529_));
 sg13g2_a21oi_1 _1400_ (.A1(_0523_),
    .A2(_0540_),
    .Y(_0542_),
    .B1(_0541_));
 sg13g2_a21o_1 _1401_ (.A2(_0540_),
    .A1(_0523_),
    .B1(_0541_),
    .X(_0543_));
 sg13g2_xor2_1 _1402_ (.B(_0433_),
    .A(\system_inst.leak_rate_2[4] ),
    .X(_0544_));
 sg13g2_mux2_1 _1403_ (.A0(_0025_),
    .A1(_0544_),
    .S(_0504_),
    .X(_0545_));
 sg13g2_nor2b_1 _1404_ (.A(_0449_),
    .B_N(_0545_),
    .Y(_0546_));
 sg13g2_xor2_1 _1405_ (.B(_0545_),
    .A(_0449_),
    .X(_0547_));
 sg13g2_inv_1 _1406_ (.Y(_0548_),
    .A(_0547_));
 sg13g2_xor2_1 _1407_ (.B(_0434_),
    .A(\system_inst.leak_rate_2[5] ),
    .X(_0549_));
 sg13g2_mux2_1 _1408_ (.A0(_0024_),
    .A1(_0549_),
    .S(_0504_),
    .X(_0550_));
 sg13g2_nand2b_1 _1409_ (.Y(_0551_),
    .B(_0446_),
    .A_N(_0550_));
 sg13g2_and2_1 _1410_ (.A(_0445_),
    .B(_0550_),
    .X(_0552_));
 sg13g2_xnor2_1 _1411_ (.Y(_0553_),
    .A(_0445_),
    .B(_0550_));
 sg13g2_or2_1 _1412_ (.X(_0554_),
    .B(_0553_),
    .A(_0547_));
 sg13g2_a21oi_1 _1413_ (.A1(_0546_),
    .A2(_0551_),
    .Y(_0555_),
    .B1(_0552_));
 sg13g2_o21ai_1 _1414_ (.B1(_0555_),
    .Y(_0556_),
    .A1(_0542_),
    .A2(_0554_));
 sg13g2_xor2_1 _1415_ (.B(_0435_),
    .A(\system_inst.leak_rate_2[6] ),
    .X(_0557_));
 sg13g2_mux2_1 _1416_ (.A0(_0023_),
    .A1(_0557_),
    .S(_0504_),
    .X(_0558_));
 sg13g2_nor2b_1 _1417_ (.A(_0440_),
    .B_N(_0558_),
    .Y(_0559_));
 sg13g2_xnor2_1 _1418_ (.Y(_0560_),
    .A(_0440_),
    .B(_0558_));
 sg13g2_and2_1 _1419_ (.A(_0509_),
    .B(_0560_),
    .X(_0561_));
 sg13g2_o21ai_1 _1420_ (.B1(_0559_),
    .Y(_0562_),
    .A1(_0431_),
    .A2(_0508_));
 sg13g2_a21oi_1 _1421_ (.A1(_0431_),
    .A2(_0508_),
    .Y(_0563_),
    .B1(net159));
 sg13g2_nand2_1 _1422_ (.Y(_0564_),
    .A(_0562_),
    .B(_0563_));
 sg13g2_a21oi_2 _1423_ (.B1(_0564_),
    .Y(_0565_),
    .A2(_0561_),
    .A1(_0556_));
 sg13g2_a21oi_2 _1424_ (.B1(_0494_),
    .Y(_0566_),
    .A2(_0506_),
    .A1(_0205_));
 sg13g2_xnor2_1 _1425_ (.Y(_0567_),
    .A(_0565_),
    .B(_0566_));
 sg13g2_xor2_1 _1426_ (.B(_0566_),
    .A(_0565_),
    .X(_0568_));
 sg13g2_xor2_1 _1427_ (.B(_0560_),
    .A(_0556_),
    .X(_0569_));
 sg13g2_nor2_1 _1428_ (.A(_0205_),
    .B(_0440_),
    .Y(_0570_));
 sg13g2_a21oi_1 _1429_ (.A1(_0205_),
    .A2(_0569_),
    .Y(_0571_),
    .B1(_0570_));
 sg13g2_nor2_2 _1430_ (.A(net152),
    .B(_0571_),
    .Y(_0572_));
 sg13g2_xnor2_1 _1431_ (.Y(_0573_),
    .A(_0160_),
    .B(_0572_));
 sg13g2_a21oi_1 _1432_ (.A1(_0556_),
    .A2(_0560_),
    .Y(_0574_),
    .B1(_0559_));
 sg13g2_or2_1 _1433_ (.X(_0575_),
    .B(_0574_),
    .A(_0509_));
 sg13g2_a21oi_1 _1434_ (.A1(_0509_),
    .A2(_0574_),
    .Y(_0576_),
    .B1(net159));
 sg13g2_a221oi_1 _1435_ (.B2(_0576_),
    .C1(net152),
    .B1(_0575_),
    .A1(net159),
    .Y(_0577_),
    .A2(_0430_));
 sg13g2_nand2_1 _1436_ (.Y(_0578_),
    .A(_0009_),
    .B(_0577_));
 sg13g2_xnor2_1 _1437_ (.Y(_0579_),
    .A(_0009_),
    .B(_0577_));
 sg13g2_nor2_1 _1438_ (.A(_0573_),
    .B(_0579_),
    .Y(_0580_));
 sg13g2_a21oi_1 _1439_ (.A1(_0543_),
    .A2(_0548_),
    .Y(_0581_),
    .B1(_0546_));
 sg13g2_xor2_1 _1440_ (.B(_0581_),
    .A(_0553_),
    .X(_0582_));
 sg13g2_nand2_1 _1441_ (.Y(_0583_),
    .A(net159),
    .B(_0446_));
 sg13g2_o21ai_1 _1442_ (.B1(_0583_),
    .Y(_0584_),
    .A1(net159),
    .A2(_0582_));
 sg13g2_nor2_2 _1443_ (.A(net152),
    .B(_0584_),
    .Y(_0585_));
 sg13g2_xnor2_1 _1444_ (.Y(_0586_),
    .A(_0011_),
    .B(_0585_));
 sg13g2_xnor2_1 _1445_ (.Y(_0587_),
    .A(_0542_),
    .B(_0548_));
 sg13g2_nand2_1 _1446_ (.Y(_0588_),
    .A(net159),
    .B(_0449_));
 sg13g2_o21ai_1 _1447_ (.B1(_0588_),
    .Y(_0589_),
    .A1(net159),
    .A2(_0587_));
 sg13g2_nor2_2 _1448_ (.A(net152),
    .B(_0589_),
    .Y(_0590_));
 sg13g2_o21ai_1 _1449_ (.B1(\system_inst.neuron.threshold[4] ),
    .Y(_0591_),
    .A1(net152),
    .A2(_0589_));
 sg13g2_xnor2_1 _1450_ (.Y(_0592_),
    .A(_0164_),
    .B(_0590_));
 sg13g2_or4_1 _1451_ (.A(_0573_),
    .B(_0579_),
    .C(_0586_),
    .D(_0592_),
    .X(_0593_));
 sg13g2_o21ai_1 _1452_ (.B1(_0537_),
    .Y(_0594_),
    .A1(_0522_),
    .A2(_0538_));
 sg13g2_nand2_1 _1453_ (.Y(_0595_),
    .A(_0532_),
    .B(_0594_));
 sg13g2_nor2_1 _1454_ (.A(_0532_),
    .B(_0594_),
    .Y(_0596_));
 sg13g2_nor2_1 _1455_ (.A(net160),
    .B(_0596_),
    .Y(_0597_));
 sg13g2_a22oi_1 _1456_ (.Y(_0598_),
    .B1(_0595_),
    .B2(_0597_),
    .A2(_0457_),
    .A1(net160));
 sg13g2_o21ai_1 _1457_ (.B1(_0166_),
    .Y(_0599_),
    .A1(net153),
    .A2(_0598_));
 sg13g2_nand3b_1 _1458_ (.B(_0012_),
    .C(_0568_),
    .Y(_0600_),
    .A_N(_0598_));
 sg13g2_xnor2_1 _1459_ (.Y(_0601_),
    .A(_0522_),
    .B(_0539_));
 sg13g2_mux2_1 _1460_ (.A0(_0460_),
    .A1(_0601_),
    .S(_0205_),
    .X(_0602_));
 sg13g2_inv_1 _1461_ (.Y(_0603_),
    .A(_0602_));
 sg13g2_nand3_1 _1462_ (.B(_0568_),
    .C(_0602_),
    .A(_0167_),
    .Y(_0604_));
 sg13g2_o21ai_1 _1463_ (.B1(\system_inst.neuron.threshold[2] ),
    .Y(_0605_),
    .A1(net153),
    .A2(_0603_));
 sg13g2_nand4_1 _1464_ (.B(_0600_),
    .C(_0604_),
    .A(_0599_),
    .Y(_0606_),
    .D(_0605_));
 sg13g2_nand2_1 _1465_ (.Y(_0607_),
    .A(\system_inst.leak_rate_2[0] ),
    .B(_0205_));
 sg13g2_xnor2_1 _1466_ (.Y(_0608_),
    .A(_0464_),
    .B(_0607_));
 sg13g2_nor2_1 _1467_ (.A(net153),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_nor3_1 _1468_ (.A(\system_inst.neuron.threshold[0] ),
    .B(net153),
    .C(_0608_),
    .Y(_0610_));
 sg13g2_o21ai_1 _1469_ (.B1(_0517_),
    .Y(_0611_),
    .A1(_0515_),
    .A2(_0519_));
 sg13g2_nand2_1 _1470_ (.Y(_0612_),
    .A(_0521_),
    .B(_0611_));
 sg13g2_mux2_1 _1471_ (.A0(_0469_),
    .A1(_0612_),
    .S(_0205_),
    .X(_0613_));
 sg13g2_nor2_1 _1472_ (.A(net153),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_o21ai_1 _1473_ (.B1(\system_inst.neuron.threshold[1] ),
    .Y(_0615_),
    .A1(net153),
    .A2(_0613_));
 sg13g2_nand3b_1 _1474_ (.B(_0568_),
    .C(_0169_),
    .Y(_0616_),
    .A_N(_0613_));
 sg13g2_nand2_1 _1475_ (.Y(_0617_),
    .A(_0615_),
    .B(_0616_));
 sg13g2_nand3b_1 _1476_ (.B(_0615_),
    .C(_0616_),
    .Y(_0618_),
    .A_N(_0610_));
 sg13g2_or2_1 _1477_ (.X(_0619_),
    .B(_0614_),
    .A(_0014_));
 sg13g2_a21o_1 _1478_ (.A2(_0619_),
    .A1(_0618_),
    .B1(_0606_),
    .X(_0620_));
 sg13g2_o21ai_1 _1479_ (.B1(_0168_),
    .Y(_0621_),
    .A1(net153),
    .A2(_0603_));
 sg13g2_nand2_1 _1480_ (.Y(_0622_),
    .A(_0599_),
    .B(_0621_));
 sg13g2_nand2_1 _1481_ (.Y(_0623_),
    .A(_0600_),
    .B(_0622_));
 sg13g2_a21o_1 _1482_ (.A2(_0623_),
    .A1(_0620_),
    .B1(_0593_),
    .X(_0624_));
 sg13g2_o21ai_1 _1483_ (.B1(\system_inst.neuron.threshold[5] ),
    .Y(_0625_),
    .A1(net152),
    .A2(_0584_));
 sg13g2_o21ai_1 _1484_ (.B1(_0625_),
    .Y(_0626_),
    .A1(_0586_),
    .A2(_0591_));
 sg13g2_o21ai_1 _1485_ (.B1(_0161_),
    .Y(_0627_),
    .A1(net152),
    .A2(_0571_));
 sg13g2_o21ai_1 _1486_ (.B1(_0627_),
    .Y(_0628_),
    .A1(_0009_),
    .A2(_0577_));
 sg13g2_a22oi_1 _1487_ (.Y(_0629_),
    .B1(_0628_),
    .B2(_0578_),
    .A2(_0626_),
    .A1(_0580_));
 sg13g2_xnor2_1 _1488_ (.Y(_0630_),
    .A(_0029_),
    .B(_0609_));
 sg13g2_nor4_1 _1489_ (.A(_0593_),
    .B(_0606_),
    .C(_0617_),
    .D(_0630_),
    .Y(_0631_));
 sg13g2_a21o_2 _1490_ (.A2(_0629_),
    .A1(_0624_),
    .B1(_0631_),
    .X(_0632_));
 sg13g2_nor2_2 _1491_ (.A(net181),
    .B(_0217_),
    .Y(_0633_));
 sg13g2_nand2_1 _1492_ (.Y(_0634_),
    .A(_0609_),
    .B(_0633_));
 sg13g2_o21ai_1 _1493_ (.B1(_0220_),
    .Y(_0043_),
    .A1(net151),
    .A2(_0634_));
 sg13g2_nand2_1 _1494_ (.Y(_0635_),
    .A(net126),
    .B(_0218_));
 sg13g2_nand2_1 _1495_ (.Y(_0636_),
    .A(_0614_),
    .B(_0633_));
 sg13g2_o21ai_1 _1496_ (.B1(_0635_),
    .Y(_0044_),
    .A1(net151),
    .A2(_0636_));
 sg13g2_nand2_1 _1497_ (.Y(_0637_),
    .A(net131),
    .B(net163));
 sg13g2_nand3_1 _1498_ (.B(_0602_),
    .C(_0633_),
    .A(_0568_),
    .Y(_0638_));
 sg13g2_o21ai_1 _1499_ (.B1(_0637_),
    .Y(_0045_),
    .A1(net151),
    .A2(_0638_));
 sg13g2_nand2_1 _1500_ (.Y(_0639_),
    .A(net198),
    .B(net163));
 sg13g2_or4_1 _1501_ (.A(net181),
    .B(_0217_),
    .C(net152),
    .D(_0598_),
    .X(_0640_));
 sg13g2_o21ai_1 _1502_ (.B1(_0639_),
    .Y(_0046_),
    .A1(net151),
    .A2(_0640_));
 sg13g2_nand2_1 _1503_ (.Y(_0641_),
    .A(net201),
    .B(net163));
 sg13g2_nand2_1 _1504_ (.Y(_0642_),
    .A(_0590_),
    .B(_0633_));
 sg13g2_o21ai_1 _1505_ (.B1(_0641_),
    .Y(_0047_),
    .A1(net151),
    .A2(_0642_));
 sg13g2_nand2_1 _1506_ (.Y(_0643_),
    .A(net200),
    .B(net163));
 sg13g2_nand2_1 _1507_ (.Y(_0644_),
    .A(_0585_),
    .B(_0633_));
 sg13g2_o21ai_1 _1508_ (.B1(_0643_),
    .Y(_0048_),
    .A1(net149),
    .A2(_0644_));
 sg13g2_nand2_1 _1509_ (.Y(_0645_),
    .A(net146),
    .B(net163));
 sg13g2_nand2_1 _1510_ (.Y(_0646_),
    .A(_0572_),
    .B(_0633_));
 sg13g2_o21ai_1 _1511_ (.B1(_0645_),
    .Y(_0049_),
    .A1(net149),
    .A2(_0646_));
 sg13g2_nand2_1 _1512_ (.Y(_0647_),
    .A(net109),
    .B(net163));
 sg13g2_nand2_1 _1513_ (.Y(_0648_),
    .A(_0577_),
    .B(_0633_));
 sg13g2_o21ai_1 _1514_ (.B1(_0647_),
    .Y(_0050_),
    .A1(net151),
    .A2(_0648_));
 sg13g2_and2_1 _1515_ (.A(net177),
    .B(net163),
    .X(_0051_));
 sg13g2_and2_1 _1516_ (.A(_0632_),
    .B(_0633_),
    .X(_0052_));
 sg13g2_nor2_2 _1517_ (.A(_0197_),
    .B(_0215_),
    .Y(_0649_));
 sg13g2_a21oi_2 _1518_ (.B1(_0649_),
    .Y(_0650_),
    .A2(_0632_),
    .A1(_0216_));
 sg13g2_nor2b_1 _1519_ (.A(_0650_),
    .B_N(net241),
    .Y(_0651_));
 sg13g2_o21ai_1 _1520_ (.B1(net191),
    .Y(_0652_),
    .A1(net241),
    .A2(_0649_));
 sg13g2_nor2_1 _1521_ (.A(_0651_),
    .B(_0652_),
    .Y(_0053_));
 sg13g2_xnor2_1 _1522_ (.Y(_0653_),
    .A(net196),
    .B(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_a22oi_1 _1523_ (.Y(_0654_),
    .B1(_0653_),
    .B2(_0649_),
    .A2(_0650_),
    .A1(net196));
 sg13g2_nor2_1 _1524_ (.A(net183),
    .B(net197),
    .Y(_0054_));
 sg13g2_nor3_1 _1525_ (.A(_0156_),
    .B(_0197_),
    .C(_0213_),
    .Y(_0655_));
 sg13g2_o21ai_1 _1526_ (.B1(_0156_),
    .Y(_0656_),
    .A1(_0213_),
    .A2(_0650_));
 sg13g2_nor2_1 _1527_ (.A(net183),
    .B(_0655_),
    .Y(_0657_));
 sg13g2_and2_1 _1528_ (.A(net262),
    .B(_0657_),
    .X(_0055_));
 sg13g2_nand2_1 _1529_ (.Y(_0658_),
    .A(net110),
    .B(net192));
 sg13g2_a21oi_1 _1530_ (.A1(_0196_),
    .A2(_0214_),
    .Y(_0056_),
    .B1(_0658_));
 sg13g2_nand2_1 _1531_ (.Y(_0659_),
    .A(\system_inst.neuron.threshold[3] ),
    .B(net176));
 sg13g2_nand4_1 _1532_ (.B(\system_inst.neuron.threshold[4] ),
    .C(\system_inst.neuron.threshold[3] ),
    .A(\system_inst.neuron.threshold[5] ),
    .Y(_0660_),
    .D(net176));
 sg13g2_nor2_1 _1533_ (.A(_0010_),
    .B(_0660_),
    .Y(_0661_));
 sg13g2_xnor2_1 _1534_ (.Y(_0662_),
    .A(_0009_),
    .B(_0661_));
 sg13g2_nor2_1 _1535_ (.A(_0034_),
    .B(_0659_),
    .Y(_0663_));
 sg13g2_xnor2_1 _1536_ (.Y(_0664_),
    .A(_0163_),
    .B(_0663_));
 sg13g2_nor2_1 _1537_ (.A(_0175_),
    .B(_0664_),
    .Y(_0665_));
 sg13g2_xnor2_1 _1538_ (.Y(_0666_),
    .A(_0161_),
    .B(_0660_));
 sg13g2_xnor2_1 _1539_ (.Y(_0667_),
    .A(_0032_),
    .B(_0666_));
 sg13g2_a21oi_1 _1540_ (.A1(_0175_),
    .A2(_0664_),
    .Y(_0668_),
    .B1(_0667_));
 sg13g2_xor2_1 _1541_ (.B(net176),
    .A(\system_inst.neuron.threshold[3] ),
    .X(_0669_));
 sg13g2_xnor2_1 _1542_ (.Y(_0670_),
    .A(_0034_),
    .B(_0659_));
 sg13g2_inv_1 _1543_ (.Y(_0671_),
    .A(_0670_));
 sg13g2_xnor2_1 _1544_ (.Y(_0672_),
    .A(_0035_),
    .B(_0670_));
 sg13g2_o21ai_1 _1545_ (.B1(_0672_),
    .Y(_0673_),
    .A1(_0036_),
    .A2(_0669_));
 sg13g2_nand2_1 _1546_ (.Y(_0674_),
    .A(_0036_),
    .B(_0669_));
 sg13g2_a22oi_1 _1547_ (.Y(_0675_),
    .B1(_0169_),
    .B2(\system_inst.loader.threshold_min[0] ),
    .A2(net176),
    .A1(net173));
 sg13g2_inv_1 _1548_ (.Y(_0676_),
    .A(_0675_));
 sg13g2_or2_1 _1549_ (.X(_0677_),
    .B(net176),
    .A(net173));
 sg13g2_nand2b_1 _1550_ (.Y(_0678_),
    .B(\system_inst.neuron.threshold[1] ),
    .A_N(\system_inst.loader.threshold_min[0] ));
 sg13g2_nand4_1 _1551_ (.B(_0675_),
    .C(_0677_),
    .A(_0674_),
    .Y(_0679_),
    .D(_0678_));
 sg13g2_nor2_1 _1552_ (.A(_0673_),
    .B(_0679_),
    .Y(_0680_));
 sg13g2_nand3_1 _1553_ (.B(_0668_),
    .C(_0680_),
    .A(_0029_),
    .Y(_0681_));
 sg13g2_and3_1 _1554_ (.X(_0682_),
    .A(_0674_),
    .B(_0676_),
    .C(_0677_));
 sg13g2_and2_1 _1555_ (.A(_0151_),
    .B(_0666_),
    .X(_0683_));
 sg13g2_a21oi_1 _1556_ (.A1(_0153_),
    .A2(_0671_),
    .Y(_0684_),
    .B1(_0683_));
 sg13g2_o21ai_1 _1557_ (.B1(_0684_),
    .Y(_0685_),
    .A1(_0673_),
    .A2(_0682_));
 sg13g2_a21oi_1 _1558_ (.A1(_0681_),
    .A2(_0685_),
    .Y(_0686_),
    .B1(_0665_));
 sg13g2_nor2_1 _1559_ (.A(_0668_),
    .B(_0683_),
    .Y(_0687_));
 sg13g2_nor2_1 _1560_ (.A(_0031_),
    .B(_0662_),
    .Y(_0688_));
 sg13g2_nor3_1 _1561_ (.A(_0686_),
    .B(_0687_),
    .C(_0688_),
    .Y(_0689_));
 sg13g2_nor2_1 _1562_ (.A(_0662_),
    .B(_0689_),
    .Y(_0690_));
 sg13g2_a21o_1 _1563_ (.A2(_0662_),
    .A1(_0031_),
    .B1(_0689_),
    .X(_0691_));
 sg13g2_nand2_1 _1564_ (.Y(_0692_),
    .A(net173),
    .B(net157));
 sg13g2_o21ai_1 _1565_ (.B1(_0692_),
    .Y(_0693_),
    .A1(_0168_),
    .A2(net157));
 sg13g2_nand2_1 _1566_ (.Y(_0694_),
    .A(net173),
    .B(\system_inst.loader.threshold_min[0] ));
 sg13g2_nand4_1 _1567_ (.B(\system_inst.loader.threshold_min[2] ),
    .C(net173),
    .A(\system_inst.loader.threshold_min[3] ),
    .Y(_0695_),
    .D(\system_inst.loader.threshold_min[0] ));
 sg13g2_nor3_1 _1568_ (.A(_0151_),
    .B(_0152_),
    .C(_0695_),
    .Y(_0696_));
 sg13g2_nand2_1 _1569_ (.Y(_0697_),
    .A(\system_inst.loader.threshold_min[6] ),
    .B(_0696_));
 sg13g2_xor2_1 _1570_ (.B(_0697_),
    .A(\system_inst.loader.threshold_min[7] ),
    .X(_0698_));
 sg13g2_nand2b_1 _1571_ (.Y(_0699_),
    .B(_0009_),
    .A_N(_0698_));
 sg13g2_xnor2_1 _1572_ (.Y(_0700_),
    .A(_0031_),
    .B(_0696_));
 sg13g2_nor2_1 _1573_ (.A(_0033_),
    .B(_0695_),
    .Y(_0701_));
 sg13g2_xnor2_1 _1574_ (.Y(_0702_),
    .A(_0032_),
    .B(_0701_));
 sg13g2_nand2_1 _1575_ (.Y(_0703_),
    .A(_0162_),
    .B(_0702_));
 sg13g2_xnor2_1 _1576_ (.Y(_0704_),
    .A(_0175_),
    .B(_0695_));
 sg13g2_nand2_2 _1577_ (.Y(_0705_),
    .A(_0169_),
    .B(_0171_));
 sg13g2_nand2_1 _1578_ (.Y(_0706_),
    .A(\system_inst.neuron.threshold[1] ),
    .B(\system_inst.neuron.threshold[0] ));
 sg13g2_and2_1 _1579_ (.A(_0678_),
    .B(_0706_),
    .X(_0707_));
 sg13g2_o21ai_1 _1580_ (.B1(_0694_),
    .Y(_0708_),
    .A1(net173),
    .A2(_0707_));
 sg13g2_nor2_1 _1581_ (.A(_0036_),
    .B(_0694_),
    .Y(_0709_));
 sg13g2_xor2_1 _1582_ (.B(_0694_),
    .A(_0036_),
    .X(_0710_));
 sg13g2_xnor2_1 _1583_ (.Y(_0711_),
    .A(_0013_),
    .B(_0710_));
 sg13g2_a21o_1 _1584_ (.A2(_0708_),
    .A1(_0705_),
    .B1(_0711_),
    .X(_0712_));
 sg13g2_xor2_1 _1585_ (.B(_0709_),
    .A(_0035_),
    .X(_0713_));
 sg13g2_nor2_1 _1586_ (.A(\system_inst.neuron.threshold[3] ),
    .B(_0713_),
    .Y(_0714_));
 sg13g2_a21oi_1 _1587_ (.A1(_0167_),
    .A2(_0710_),
    .Y(_0715_),
    .B1(_0714_));
 sg13g2_nor2_1 _1588_ (.A(_0034_),
    .B(_0704_),
    .Y(_0716_));
 sg13g2_a221oi_1 _1589_ (.B2(_0712_),
    .C1(_0716_),
    .B1(_0715_),
    .A1(\system_inst.neuron.threshold[3] ),
    .Y(_0717_),
    .A2(_0713_));
 sg13g2_a21oi_1 _1590_ (.A1(_0034_),
    .A2(_0704_),
    .Y(_0718_),
    .B1(_0717_));
 sg13g2_xnor2_1 _1591_ (.Y(_0719_),
    .A(_0011_),
    .B(_0702_));
 sg13g2_o21ai_1 _1592_ (.B1(_0703_),
    .Y(_0720_),
    .A1(_0718_),
    .A2(_0719_));
 sg13g2_xnor2_1 _1593_ (.Y(_0721_),
    .A(_0161_),
    .B(_0700_));
 sg13g2_a22oi_1 _1594_ (.Y(_0722_),
    .B1(_0720_),
    .B2(_0721_),
    .A2(_0700_),
    .A1(_0160_));
 sg13g2_xnor2_1 _1595_ (.Y(_0723_),
    .A(\system_inst.neuron.threshold[7] ),
    .B(_0698_));
 sg13g2_o21ai_1 _1596_ (.B1(_0699_),
    .Y(_0724_),
    .A1(_0722_),
    .A2(_0723_));
 sg13g2_nand2_1 _1597_ (.Y(_0725_),
    .A(\system_inst.loader.threshold_min[2] ),
    .B(net155));
 sg13g2_nor2_1 _1598_ (.A(net176),
    .B(_0705_),
    .Y(_0726_));
 sg13g2_xnor2_1 _1599_ (.Y(_0727_),
    .A(_0167_),
    .B(_0705_));
 sg13g2_o21ai_1 _1600_ (.B1(_0725_),
    .Y(_0728_),
    .A1(net155),
    .A2(_0727_));
 sg13g2_mux2_1 _1601_ (.A0(_0728_),
    .A1(_0693_),
    .S(net149),
    .X(_0729_));
 sg13g2_nand2_1 _1602_ (.Y(_0730_),
    .A(net186),
    .B(_0729_));
 sg13g2_nand2_1 _1603_ (.Y(_0731_),
    .A(net186),
    .B(net162));
 sg13g2_o21ai_1 _1604_ (.B1(_0219_),
    .Y(_0732_),
    .A1(net151),
    .A2(_0731_));
 sg13g2_a21oi_1 _1605_ (.A1(net265),
    .A2(net180),
    .Y(_0733_),
    .B1(net148));
 sg13g2_a22oi_1 _1606_ (.Y(_0057_),
    .B1(_0733_),
    .B2(_0730_),
    .A2(net148),
    .A1(_0167_));
 sg13g2_mux2_1 _1607_ (.A0(_0669_),
    .A1(\system_inst.loader.threshold_min[2] ),
    .S(net157),
    .X(_0734_));
 sg13g2_nand2_1 _1608_ (.Y(_0735_),
    .A(\system_inst.loader.threshold_min[3] ),
    .B(net155));
 sg13g2_nor3_1 _1609_ (.A(\system_inst.neuron.threshold[3] ),
    .B(net176),
    .C(_0705_),
    .Y(_0736_));
 sg13g2_xnor2_1 _1610_ (.Y(_0737_),
    .A(\system_inst.neuron.threshold[3] ),
    .B(_0726_));
 sg13g2_o21ai_1 _1611_ (.B1(_0735_),
    .Y(_0738_),
    .A1(net155),
    .A2(_0737_));
 sg13g2_mux2_1 _1612_ (.A0(_0738_),
    .A1(_0734_),
    .S(net149),
    .X(_0739_));
 sg13g2_nand2_1 _1613_ (.Y(_0740_),
    .A(net186),
    .B(_0739_));
 sg13g2_a21oi_1 _1614_ (.A1(net246),
    .A2(net180),
    .Y(_0741_),
    .B1(net148));
 sg13g2_a22oi_1 _1615_ (.Y(_0058_),
    .B1(_0740_),
    .B2(_0741_),
    .A2(net148),
    .A1(_0165_));
 sg13g2_nor2_1 _1616_ (.A(_0670_),
    .B(net156),
    .Y(_0742_));
 sg13g2_a21oi_1 _1617_ (.A1(net246),
    .A2(net156),
    .Y(_0743_),
    .B1(_0742_));
 sg13g2_nand2_1 _1618_ (.Y(_0744_),
    .A(\system_inst.loader.threshold_min[4] ),
    .B(net154));
 sg13g2_and2_1 _1619_ (.A(_0164_),
    .B(_0736_),
    .X(_0745_));
 sg13g2_xnor2_1 _1620_ (.Y(_0746_),
    .A(\system_inst.neuron.threshold[4] ),
    .B(_0736_));
 sg13g2_o21ai_1 _1621_ (.B1(_0744_),
    .Y(_0747_),
    .A1(net154),
    .A2(_0746_));
 sg13g2_o21ai_1 _1622_ (.B1(net186),
    .Y(_0748_),
    .A1(net150),
    .A2(_0747_));
 sg13g2_a21o_1 _1623_ (.A2(_0743_),
    .A1(net150),
    .B1(_0748_),
    .X(_0749_));
 sg13g2_a21oi_1 _1624_ (.A1(net230),
    .A2(net179),
    .Y(_0750_),
    .B1(net147));
 sg13g2_a22oi_1 _1625_ (.Y(_0059_),
    .B1(_0749_),
    .B2(_0750_),
    .A2(net147),
    .A1(_0164_));
 sg13g2_nor2_1 _1626_ (.A(_0664_),
    .B(net156),
    .Y(_0751_));
 sg13g2_a21oi_1 _1627_ (.A1(net230),
    .A2(net156),
    .Y(_0752_),
    .B1(_0751_));
 sg13g2_nand2_1 _1628_ (.Y(_0753_),
    .A(\system_inst.loader.threshold_min[5] ),
    .B(net154));
 sg13g2_and2_1 _1629_ (.A(_0162_),
    .B(_0745_),
    .X(_0754_));
 sg13g2_xnor2_1 _1630_ (.Y(_0755_),
    .A(\system_inst.neuron.threshold[5] ),
    .B(_0745_));
 sg13g2_o21ai_1 _1631_ (.B1(_0753_),
    .Y(_0756_),
    .A1(net154),
    .A2(_0755_));
 sg13g2_o21ai_1 _1632_ (.B1(net185),
    .Y(_0757_),
    .A1(net150),
    .A2(_0756_));
 sg13g2_a21o_1 _1633_ (.A2(_0752_),
    .A1(net150),
    .B1(_0757_),
    .X(_0758_));
 sg13g2_a21oi_1 _1634_ (.A1(net231),
    .A2(net179),
    .Y(_0759_),
    .B1(net147));
 sg13g2_a22oi_1 _1635_ (.Y(_0060_),
    .B1(_0758_),
    .B2(_0759_),
    .A2(net147),
    .A1(_0162_));
 sg13g2_nor2_1 _1636_ (.A(_0666_),
    .B(net156),
    .Y(_0760_));
 sg13g2_a21oi_1 _1637_ (.A1(_0151_),
    .A2(net156),
    .Y(_0761_),
    .B1(_0760_));
 sg13g2_nand2_1 _1638_ (.Y(_0762_),
    .A(\system_inst.loader.threshold_min[6] ),
    .B(net154));
 sg13g2_nand2_1 _1639_ (.Y(_0763_),
    .A(_0160_),
    .B(_0754_));
 sg13g2_xnor2_1 _1640_ (.Y(_0764_),
    .A(\system_inst.neuron.threshold[6] ),
    .B(_0754_));
 sg13g2_o21ai_1 _1641_ (.B1(_0762_),
    .Y(_0765_),
    .A1(net154),
    .A2(_0764_));
 sg13g2_mux2_1 _1642_ (.A0(_0765_),
    .A1(_0761_),
    .S(net150),
    .X(_0766_));
 sg13g2_nand2_1 _1643_ (.Y(_0767_),
    .A(net184),
    .B(_0766_));
 sg13g2_a21oi_1 _1644_ (.A1(net225),
    .A2(net179),
    .Y(_0768_),
    .B1(net147));
 sg13g2_a22oi_1 _1645_ (.Y(_0061_),
    .B1(_0767_),
    .B2(_0768_),
    .A2(net147),
    .A1(_0160_));
 sg13g2_xnor2_1 _1646_ (.Y(_0769_),
    .A(\system_inst.neuron.threshold[7] ),
    .B(_0763_));
 sg13g2_mux2_1 _1647_ (.A0(_0769_),
    .A1(\system_inst.loader.threshold_min[7] ),
    .S(net154),
    .X(_0770_));
 sg13g2_nor2b_1 _1648_ (.A(net225),
    .B_N(net156),
    .Y(_0771_));
 sg13g2_o21ai_1 _1649_ (.B1(net150),
    .Y(_0772_),
    .A1(_0690_),
    .A2(_0771_));
 sg13g2_o21ai_1 _1650_ (.B1(net184),
    .Y(_0773_),
    .A1(net150),
    .A2(_0770_));
 sg13g2_nand2b_1 _1651_ (.Y(_0774_),
    .B(_0772_),
    .A_N(_0773_));
 sg13g2_a21oi_1 _1652_ (.A1(net257),
    .A2(net179),
    .Y(_0775_),
    .B1(net147));
 sg13g2_a22oi_1 _1653_ (.Y(_0062_),
    .B1(_0774_),
    .B2(_0775_),
    .A2(net147),
    .A1(_0159_));
 sg13g2_nand3b_1 _1654_ (.B(net186),
    .C(net149),
    .Y(_0776_),
    .A_N(net157));
 sg13g2_nand2b_1 _1655_ (.Y(_0777_),
    .B(_0776_),
    .A_N(net148));
 sg13g2_nand2_1 _1656_ (.Y(_0778_),
    .A(_0038_),
    .B(net155));
 sg13g2_o21ai_1 _1657_ (.B1(_0778_),
    .Y(_0779_),
    .A1(_0171_),
    .A2(net154));
 sg13g2_nor3_1 _1658_ (.A(net180),
    .B(net149),
    .C(_0779_),
    .Y(_0780_));
 sg13g2_a21o_1 _1659_ (.A2(net179),
    .A1(\system_inst.loader.threshold_min[0] ),
    .B1(_0780_),
    .X(_0781_));
 sg13g2_mux2_1 _1660_ (.A0(_0781_),
    .A1(net234),
    .S(_0777_),
    .X(_0063_));
 sg13g2_nand2b_1 _1661_ (.Y(_0782_),
    .B(net156),
    .A_N(_0038_));
 sg13g2_and2_1 _1662_ (.A(net149),
    .B(_0782_),
    .X(_0783_));
 sg13g2_a21oi_1 _1663_ (.A1(_0705_),
    .A2(_0706_),
    .Y(_0784_),
    .B1(net155));
 sg13g2_a21o_1 _1664_ (.A2(net155),
    .A1(\system_inst.loader.threshold_min[1] ),
    .B1(_0784_),
    .X(_0785_));
 sg13g2_o21ai_1 _1665_ (.B1(net186),
    .Y(_0786_),
    .A1(net149),
    .A2(_0785_));
 sg13g2_nand2_1 _1666_ (.Y(_0787_),
    .A(net173),
    .B(net180));
 sg13g2_o21ai_1 _1667_ (.B1(_0787_),
    .Y(_0788_),
    .A1(_0783_),
    .A2(_0786_));
 sg13g2_mux2_1 _1668_ (.A0(_0788_),
    .A1(net267),
    .S(_0777_),
    .X(_0064_));
 sg13g2_or2_1 _1669_ (.X(_0789_),
    .B(\system_inst.loader.current_state[4] ),
    .A(\system_inst.loader.current_state[2] ));
 sg13g2_nor4_2 _1670_ (.A(\system_inst.loader.current_state[5] ),
    .B(\system_inst.loader.current_state[1] ),
    .C(\system_inst.loader.current_state[6] ),
    .Y(_0790_),
    .D(_0789_));
 sg13g2_nand2_1 _1671_ (.Y(_0791_),
    .A(_0037_),
    .B(_0790_));
 sg13g2_nor2_1 _1672_ (.A(net132),
    .B(_0791_),
    .Y(_0792_));
 sg13g2_o21ai_1 _1673_ (.B1(net1),
    .Y(_0793_),
    .A1(_0173_),
    .A2(net3));
 sg13g2_nor2_1 _1674_ (.A(_0792_),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_o21ai_1 _1675_ (.B1(_0790_),
    .Y(_0795_),
    .A1(_0174_),
    .A2(_0181_));
 sg13g2_nand2_1 _1676_ (.Y(_0796_),
    .A(net3),
    .B(_0795_));
 sg13g2_nand2_1 _1677_ (.Y(_0797_),
    .A(_0794_),
    .B(_0796_));
 sg13g2_and2_1 _1678_ (.A(_0174_),
    .B(_0790_),
    .X(_0798_));
 sg13g2_a21oi_1 _1679_ (.A1(net227),
    .A2(_0797_),
    .Y(_0799_),
    .B1(net182));
 sg13g2_o21ai_1 _1680_ (.B1(_0799_),
    .Y(_0065_),
    .A1(_0797_),
    .A2(_0798_));
 sg13g2_o21ai_1 _1681_ (.B1(net192),
    .Y(_0800_),
    .A1(net268),
    .A2(_0184_));
 sg13g2_a21oi_1 _1682_ (.A1(_0149_),
    .A2(_0184_),
    .Y(_0066_),
    .B1(_0800_));
 sg13g2_a21oi_1 _1683_ (.A1(\system_inst.loader.weight_a[1] ),
    .A2(_0183_),
    .Y(_0801_),
    .B1(net182));
 sg13g2_o21ai_1 _1684_ (.B1(_0801_),
    .Y(_0067_),
    .A1(_0146_),
    .A2(_0183_));
 sg13g2_o21ai_1 _1685_ (.B1(net192),
    .Y(_0802_),
    .A1(net175),
    .A2(_0184_));
 sg13g2_a21oi_1 _1686_ (.A1(_0145_),
    .A2(_0184_),
    .Y(_0068_),
    .B1(_0802_));
 sg13g2_o21ai_1 _1687_ (.B1(net193),
    .Y(_0803_),
    .A1(net259),
    .A2(net168));
 sg13g2_a21oi_1 _1688_ (.A1(_0149_),
    .A2(net168),
    .Y(_0069_),
    .B1(_0803_));
 sg13g2_a21oi_1 _1689_ (.A1(\system_inst.loader.shift_reg[0] ),
    .A2(net168),
    .Y(_0804_),
    .B1(net182));
 sg13g2_o21ai_1 _1690_ (.B1(_0804_),
    .Y(_0070_),
    .A1(_0155_),
    .A2(net168));
 sg13g2_o21ai_1 _1691_ (.B1(net190),
    .Y(_0805_),
    .A1(net228),
    .A2(_0192_));
 sg13g2_a21oi_1 _1692_ (.A1(_0145_),
    .A2(_0192_),
    .Y(_0071_),
    .B1(_0805_));
 sg13g2_o21ai_1 _1693_ (.B1(net190),
    .Y(_0806_),
    .A1(net232),
    .A2(net168));
 sg13g2_a21oi_1 _1694_ (.A1(_0144_),
    .A2(net168),
    .Y(_0072_),
    .B1(_0806_));
 sg13g2_o21ai_1 _1695_ (.B1(net187),
    .Y(_0807_),
    .A1(net238),
    .A2(net167));
 sg13g2_a21oi_1 _1696_ (.A1(_0143_),
    .A2(net167),
    .Y(_0073_),
    .B1(_0807_));
 sg13g2_o21ai_1 _1697_ (.B1(net187),
    .Y(_0808_),
    .A1(net222),
    .A2(net167));
 sg13g2_a21oi_1 _1698_ (.A1(_0142_),
    .A2(net167),
    .Y(_0074_),
    .B1(_0808_));
 sg13g2_o21ai_1 _1699_ (.B1(net187),
    .Y(_0809_),
    .A1(net207),
    .A2(net167));
 sg13g2_a21oi_1 _1700_ (.A1(_0141_),
    .A2(net167),
    .Y(_0075_),
    .B1(_0809_));
 sg13g2_o21ai_1 _1701_ (.B1(net187),
    .Y(_0810_),
    .A1(net209),
    .A2(net167));
 sg13g2_a21oi_1 _1702_ (.A1(_0140_),
    .A2(net167),
    .Y(_0076_),
    .B1(_0810_));
 sg13g2_a21oi_1 _1703_ (.A1(net4),
    .A2(net166),
    .Y(_0811_),
    .B1(net182));
 sg13g2_o21ai_1 _1704_ (.B1(_0811_),
    .Y(_0077_),
    .A1(_0154_),
    .A2(net166));
 sg13g2_o21ai_1 _1705_ (.B1(net185),
    .Y(_0812_),
    .A1(net242),
    .A2(net164));
 sg13g2_a21oi_1 _1706_ (.A1(_0146_),
    .A2(net164),
    .Y(_0078_),
    .B1(_0812_));
 sg13g2_o21ai_1 _1707_ (.B1(net185),
    .Y(_0813_),
    .A1(net205),
    .A2(net165));
 sg13g2_a21oi_1 _1708_ (.A1(_0145_),
    .A2(net165),
    .Y(_0079_),
    .B1(_0813_));
 sg13g2_o21ai_1 _1709_ (.B1(net185),
    .Y(_0814_),
    .A1(net248),
    .A2(net165));
 sg13g2_a21oi_1 _1710_ (.A1(_0144_),
    .A2(net165),
    .Y(_0080_),
    .B1(_0814_));
 sg13g2_o21ai_1 _1711_ (.B1(net185),
    .Y(_0815_),
    .A1(net237),
    .A2(net165));
 sg13g2_a21oi_1 _1712_ (.A1(_0143_),
    .A2(net165),
    .Y(_0081_),
    .B1(_0815_));
 sg13g2_o21ai_1 _1713_ (.B1(net184),
    .Y(_0816_),
    .A1(net236),
    .A2(net164));
 sg13g2_a21oi_1 _1714_ (.A1(_0142_),
    .A2(net164),
    .Y(_0082_),
    .B1(_0816_));
 sg13g2_o21ai_1 _1715_ (.B1(net184),
    .Y(_0817_),
    .A1(net219),
    .A2(net164));
 sg13g2_a21oi_1 _1716_ (.A1(_0141_),
    .A2(net164),
    .Y(_0083_),
    .B1(_0817_));
 sg13g2_o21ai_1 _1717_ (.B1(net184),
    .Y(_0818_),
    .A1(net217),
    .A2(net164));
 sg13g2_a21oi_1 _1718_ (.A1(_0140_),
    .A2(net164),
    .Y(_0084_),
    .B1(_0818_));
 sg13g2_o21ai_1 _1719_ (.B1(net186),
    .Y(_0819_),
    .A1(net256),
    .A2(net170));
 sg13g2_a21oi_1 _1720_ (.A1(_0149_),
    .A2(net170),
    .Y(_0085_),
    .B1(_0819_));
 sg13g2_a21oi_1 _1721_ (.A1(net173),
    .A2(_0190_),
    .Y(_0820_),
    .B1(net179));
 sg13g2_o21ai_1 _1722_ (.B1(_0820_),
    .Y(_0086_),
    .A1(_0146_),
    .A2(_0190_));
 sg13g2_a21oi_1 _1723_ (.A1(net265),
    .A2(_0190_),
    .Y(_0821_),
    .B1(net179));
 sg13g2_o21ai_1 _1724_ (.B1(_0821_),
    .Y(_0087_),
    .A1(_0145_),
    .A2(_0190_));
 sg13g2_a21oi_2 _1725_ (.B1(net182),
    .Y(_0822_),
    .A2(_0189_),
    .A1(\system_inst.loader.shift_reg[2] ));
 sg13g2_o21ai_1 _1726_ (.B1(_0822_),
    .Y(_0088_),
    .A1(_0153_),
    .A2(net170));
 sg13g2_a21oi_1 _1727_ (.A1(net226),
    .A2(net169),
    .Y(_0823_),
    .B1(net179));
 sg13g2_o21ai_1 _1728_ (.B1(_0823_),
    .Y(_0089_),
    .A1(_0152_),
    .A2(net169));
 sg13g2_o21ai_1 _1729_ (.B1(net184),
    .Y(_0824_),
    .A1(net231),
    .A2(net169));
 sg13g2_a21oi_1 _1730_ (.A1(_0142_),
    .A2(net169),
    .Y(_0090_),
    .B1(_0824_));
 sg13g2_o21ai_1 _1731_ (.B1(net184),
    .Y(_0825_),
    .A1(net225),
    .A2(net169));
 sg13g2_a21oi_1 _1732_ (.A1(_0141_),
    .A2(net169),
    .Y(_0091_),
    .B1(_0825_));
 sg13g2_o21ai_1 _1733_ (.B1(net184),
    .Y(_0826_),
    .A1(\system_inst.loader.threshold_min[7] ),
    .A2(net169));
 sg13g2_a21oi_1 _1734_ (.A1(_0140_),
    .A2(net169),
    .Y(_0092_),
    .B1(_0826_));
 sg13g2_o21ai_1 _1735_ (.B1(net189),
    .Y(_0827_),
    .A1(net143),
    .A2(net171));
 sg13g2_a21oi_1 _1736_ (.A1(_0149_),
    .A2(net171),
    .Y(_0093_),
    .B1(_0827_));
 sg13g2_a21oi_1 _1737_ (.A1(\system_inst.loader.shift_reg[0] ),
    .A2(net171),
    .Y(_0828_),
    .B1(net182));
 sg13g2_o21ai_1 _1738_ (.B1(_0828_),
    .Y(_0094_),
    .A1(_0150_),
    .A2(net171));
 sg13g2_o21ai_1 _1739_ (.B1(net189),
    .Y(_0829_),
    .A1(net220),
    .A2(net171));
 sg13g2_a21oi_1 _1740_ (.A1(_0145_),
    .A2(net171),
    .Y(_0095_),
    .B1(_0829_));
 sg13g2_o21ai_1 _1741_ (.B1(net188),
    .Y(_0830_),
    .A1(net223),
    .A2(net171));
 sg13g2_a21oi_1 _1742_ (.A1(_0144_),
    .A2(net171),
    .Y(_0096_),
    .B1(_0830_));
 sg13g2_and3_2 _1743_ (.X(_0831_),
    .A(net133),
    .B(net178),
    .C(net172));
 sg13g2_o21ai_1 _1744_ (.B1(net188),
    .Y(_0832_),
    .A1(net199),
    .A2(_0831_));
 sg13g2_a21oi_1 _1745_ (.A1(_0149_),
    .A2(_0831_),
    .Y(_0097_),
    .B1(_0832_));
 sg13g2_o21ai_1 _1746_ (.B1(net188),
    .Y(_0833_),
    .A1(net211),
    .A2(_0831_));
 sg13g2_a21oi_1 _1747_ (.A1(_0146_),
    .A2(_0831_),
    .Y(_0098_),
    .B1(_0833_));
 sg13g2_a21oi_1 _1748_ (.A1(\system_inst.loader.shift_reg[1] ),
    .A2(_0831_),
    .Y(_0834_),
    .B1(net182));
 sg13g2_o21ai_1 _1749_ (.B1(_0834_),
    .Y(_0099_),
    .A1(_0148_),
    .A2(_0831_));
 sg13g2_o21ai_1 _1750_ (.B1(net188),
    .Y(_0835_),
    .A1(net141),
    .A2(_0831_));
 sg13g2_a21oi_1 _1751_ (.A1(_0144_),
    .A2(_0831_),
    .Y(_0100_),
    .B1(_0835_));
 sg13g2_nor2_1 _1752_ (.A(net3),
    .B(_0798_),
    .Y(_0836_));
 sg13g2_nor2b_2 _1753_ (.A(_0836_),
    .B_N(_0794_),
    .Y(_0837_));
 sg13g2_nand2b_1 _1754_ (.Y(_0838_),
    .B(_0794_),
    .A_N(_0836_));
 sg13g2_o21ai_1 _1755_ (.B1(_0174_),
    .Y(_0839_),
    .A1(net172),
    .A2(_0790_));
 sg13g2_a21oi_1 _1756_ (.A1(net4),
    .A2(_0839_),
    .Y(_0840_),
    .B1(_0838_));
 sg13g2_o21ai_1 _1757_ (.B1(net189),
    .Y(_0841_),
    .A1(net250),
    .A2(_0837_));
 sg13g2_nor2_1 _1758_ (.A(_0840_),
    .B(_0841_),
    .Y(_0101_));
 sg13g2_a21oi_1 _1759_ (.A1(net250),
    .A2(_0839_),
    .Y(_0842_),
    .B1(net158));
 sg13g2_o21ai_1 _1760_ (.B1(net188),
    .Y(_0843_),
    .A1(net239),
    .A2(_0837_));
 sg13g2_nor2_1 _1761_ (.A(_0842_),
    .B(_0843_),
    .Y(_0102_));
 sg13g2_a21oi_1 _1762_ (.A1(net239),
    .A2(_0839_),
    .Y(_0844_),
    .B1(net158));
 sg13g2_o21ai_1 _1763_ (.B1(net188),
    .Y(_0115_),
    .A1(\system_inst.loader.shift_reg[2] ),
    .A2(_0837_));
 sg13g2_nor2_1 _1764_ (.A(_0844_),
    .B(_0115_),
    .Y(_0103_));
 sg13g2_a21oi_1 _1765_ (.A1(net263),
    .A2(_0839_),
    .Y(_0116_),
    .B1(net158));
 sg13g2_o21ai_1 _1766_ (.B1(net187),
    .Y(_0117_),
    .A1(net226),
    .A2(_0837_));
 sg13g2_nor2_1 _1767_ (.A(_0116_),
    .B(_0117_),
    .Y(_0104_));
 sg13g2_a21oi_1 _1768_ (.A1(net226),
    .A2(_0839_),
    .Y(_0118_),
    .B1(net158));
 sg13g2_o21ai_1 _1769_ (.B1(net187),
    .Y(_0119_),
    .A1(net204),
    .A2(_0837_));
 sg13g2_nor2_1 _1770_ (.A(_0118_),
    .B(_0119_),
    .Y(_0105_));
 sg13g2_a21oi_1 _1771_ (.A1(net204),
    .A2(_0839_),
    .Y(_0120_),
    .B1(net158));
 sg13g2_o21ai_1 _1772_ (.B1(net187),
    .Y(_0121_),
    .A1(net139),
    .A2(_0837_));
 sg13g2_nor2_1 _1773_ (.A(_0120_),
    .B(_0121_),
    .Y(_0106_));
 sg13g2_a21oi_1 _1774_ (.A1(net139),
    .A2(_0839_),
    .Y(_0122_),
    .B1(net158));
 sg13g2_o21ai_1 _1775_ (.B1(net187),
    .Y(_0123_),
    .A1(\system_inst.loader.shift_reg[6] ),
    .A2(_0837_));
 sg13g2_nor2_1 _1776_ (.A(_0122_),
    .B(_0123_),
    .Y(_0107_));
 sg13g2_nor2_1 _1777_ (.A(_0798_),
    .B(_0838_),
    .Y(_0124_));
 sg13g2_o21ai_1 _1778_ (.B1(net189),
    .Y(_0125_),
    .A1(net120),
    .A2(_0124_));
 sg13g2_a21oi_1 _1779_ (.A1(net120),
    .A2(_0837_),
    .Y(_0108_),
    .B1(_0125_));
 sg13g2_nand2_1 _1780_ (.Y(_0126_),
    .A(net124),
    .B(net158));
 sg13g2_nand3_1 _1781_ (.B(_0791_),
    .C(_0124_),
    .A(_0180_),
    .Y(_0127_));
 sg13g2_o21ai_1 _1782_ (.B1(net189),
    .Y(_0128_),
    .A1(net124),
    .A2(net120));
 sg13g2_a21oi_1 _1783_ (.A1(_0126_),
    .A2(_0127_),
    .Y(_0109_),
    .B1(_0128_));
 sg13g2_nand2_1 _1784_ (.Y(_0129_),
    .A(net112),
    .B(net158));
 sg13g2_a22oi_1 _1785_ (.Y(_0130_),
    .B1(_0790_),
    .B2(_0037_),
    .A2(_0180_),
    .A1(_0030_));
 sg13g2_nand3b_1 _1786_ (.B(_0124_),
    .C(_0130_),
    .Y(_0131_),
    .A_N(_0181_));
 sg13g2_a21oi_1 _1787_ (.A1(_0129_),
    .A2(_0131_),
    .Y(_0110_),
    .B1(net182));
 sg13g2_o21ai_1 _1788_ (.B1(net188),
    .Y(_0132_),
    .A1(_0197_),
    .A2(_0228_));
 sg13g2_xnor2_1 _1789_ (.Y(_0133_),
    .A(net215),
    .B(_0196_));
 sg13g2_nor2_1 _1790_ (.A(_0132_),
    .B(_0133_),
    .Y(_0111_));
 sg13g2_and3_1 _1791_ (.X(_0134_),
    .A(net121),
    .B(\system_inst.neuron.leak_counter_1[0] ),
    .C(_0196_));
 sg13g2_a21oi_1 _1792_ (.A1(\system_inst.neuron.leak_counter_1[0] ),
    .A2(_0196_),
    .Y(_0135_),
    .B1(net121));
 sg13g2_nor3_1 _1793_ (.A(_0132_),
    .B(_0134_),
    .C(net122),
    .Y(_0112_));
 sg13g2_nand2_1 _1794_ (.Y(_0136_),
    .A(net144),
    .B(_0134_));
 sg13g2_xnor2_1 _1795_ (.Y(_0137_),
    .A(net144),
    .B(_0134_));
 sg13g2_nor2_1 _1796_ (.A(_0132_),
    .B(net145),
    .Y(_0113_));
 sg13g2_xor2_1 _1797_ (.B(_0136_),
    .A(net208),
    .X(_0138_));
 sg13g2_nor2_1 _1798_ (.A(_0132_),
    .B(_0138_),
    .Y(_0114_));
 sg13g2_dfrbp_1 _1799_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net27),
    .D(_0000_),
    .Q_N(_0891_),
    .Q(\system_inst.loader.current_state[0] ));
 sg13g2_dfrbp_1 _1800_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net28),
    .D(_0001_),
    .Q_N(_0892_),
    .Q(\system_inst.loader.current_state[1] ));
 sg13g2_dfrbp_1 _1801_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net29),
    .D(_0002_),
    .Q_N(_0893_),
    .Q(\system_inst.loader.current_state[2] ));
 sg13g2_dfrbp_1 _1802_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net30),
    .D(_0003_),
    .Q_N(_0037_),
    .Q(\system_inst.loader.current_state[3] ));
 sg13g2_dfrbp_1 _1803_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net31),
    .D(net119),
    .Q_N(_0894_),
    .Q(\system_inst.loader.current_state[4] ));
 sg13g2_dfrbp_1 _1804_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net71),
    .D(_0005_),
    .Q_N(_0895_),
    .Q(\system_inst.loader.current_state[5] ));
 sg13g2_dfrbp_1 _1805_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net26),
    .D(_0006_),
    .Q_N(_0890_),
    .Q(\system_inst.loader.current_state[6] ));
 sg13g2_dfrbp_1 _1806_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net78),
    .D(_0039_),
    .Q_N(_0889_),
    .Q(\system_inst.neuron.leak_counter_2[0] ));
 sg13g2_dfrbp_1 _1807_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net76),
    .D(net117),
    .Q_N(_0888_),
    .Q(\system_inst.neuron.leak_counter_2[1] ));
 sg13g2_dfrbp_1 _1808_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net74),
    .D(_0041_),
    .Q_N(_0887_),
    .Q(\system_inst.neuron.leak_counter_2[2] ));
 sg13g2_dfrbp_1 _1809_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net72),
    .D(_0042_),
    .Q_N(_0886_),
    .Q(\system_inst.neuron.leak_counter_2[3] ));
 sg13g2_dfrbp_1 _1810_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net70),
    .D(_0043_),
    .Q_N(_0008_),
    .Q(\system_inst.neuron.v_mem[0] ));
 sg13g2_dfrbp_1 _1811_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net68),
    .D(_0044_),
    .Q_N(_0885_),
    .Q(\system_inst.neuron.v_mem[1] ));
 sg13g2_dfrbp_1 _1812_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net66),
    .D(_0045_),
    .Q_N(_0884_),
    .Q(\system_inst.neuron.v_mem[2] ));
 sg13g2_dfrbp_1 _1813_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net64),
    .D(_0046_),
    .Q_N(_0883_),
    .Q(\system_inst.neuron.v_mem[3] ));
 sg13g2_dfrbp_1 _1814_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net62),
    .D(_0047_),
    .Q_N(_0882_),
    .Q(\system_inst.neuron.v_mem[4] ));
 sg13g2_dfrbp_1 _1815_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net60),
    .D(_0048_),
    .Q_N(_0881_),
    .Q(\system_inst.neuron.v_mem[5] ));
 sg13g2_dfrbp_1 _1816_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net58),
    .D(_0049_),
    .Q_N(_0880_),
    .Q(\system_inst.neuron.v_mem[6] ));
 sg13g2_dfrbp_1 _1817_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net56),
    .D(_0050_),
    .Q_N(_0007_),
    .Q(\system_inst.neuron.v_mem[7] ));
 sg13g2_dfrbp_1 _1818_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net54),
    .D(_0051_),
    .Q_N(_0879_),
    .Q(\system_inst.neuron.v_mem[8] ));
 sg13g2_dfrbp_1 _1819_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net52),
    .D(_0052_),
    .Q_N(_0878_),
    .Q(spike_out));
 sg13g2_dfrbp_1 _1820_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net51),
    .D(_0053_),
    .Q_N(_0877_),
    .Q(\system_inst.neuron.refr_cnt[0] ));
 sg13g2_dfrbp_1 _1821_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net49),
    .D(_0054_),
    .Q_N(_0876_),
    .Q(\system_inst.neuron.refr_cnt[1] ));
 sg13g2_dfrbp_1 _1822_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net47),
    .D(_0055_),
    .Q_N(_0875_),
    .Q(\system_inst.neuron.refr_cnt[2] ));
 sg13g2_dfrbp_1 _1823_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net45),
    .D(net111),
    .Q_N(_0874_),
    .Q(\system_inst.neuron.refr_cnt[3] ));
 sg13g2_dfrbp_1 _1824_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net43),
    .D(_0057_),
    .Q_N(_0013_),
    .Q(\system_inst.neuron.threshold[2] ));
 sg13g2_dfrbp_1 _1825_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net42),
    .D(_0058_),
    .Q_N(_0012_),
    .Q(\system_inst.neuron.threshold[3] ));
 sg13g2_dfrbp_1 _1826_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net41),
    .D(_0059_),
    .Q_N(_0034_),
    .Q(\system_inst.neuron.threshold[4] ));
 sg13g2_dfrbp_1 _1827_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net40),
    .D(_0060_),
    .Q_N(_0011_),
    .Q(\system_inst.neuron.threshold[5] ));
 sg13g2_dfrbp_1 _1828_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net39),
    .D(net245),
    .Q_N(_0010_),
    .Q(\system_inst.neuron.threshold[6] ));
 sg13g2_dfrbp_1 _1829_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net38),
    .D(net258),
    .Q_N(_0009_),
    .Q(\system_inst.neuron.threshold[7] ));
 sg13g2_dfrbp_1 _1830_ (.CLK(clknet_4_5_0_clk),
    .RESET_B(net37),
    .D(net235),
    .Q_N(_0029_),
    .Q(\system_inst.neuron.threshold[0] ));
 sg13g2_dfrbp_1 _1831_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net36),
    .D(_0064_),
    .Q_N(_0014_),
    .Q(\system_inst.neuron.threshold[1] ));
 sg13g2_dfrbp_1 _1832_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net35),
    .D(_0065_),
    .Q_N(_0873_),
    .Q(params_ready));
 sg13g2_dfrbp_1 _1833_ (.CLK(clknet_4_15_0_clk),
    .RESET_B(net33),
    .D(_0066_),
    .Q_N(_0872_),
    .Q(\system_inst.loader.weight_a[0] ));
 sg13g2_dfrbp_1 _1834_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net25),
    .D(net251),
    .Q_N(_0871_),
    .Q(\system_inst.loader.weight_a[1] ));
 sg13g2_dfrbp_1 _1835_ (.CLK(clknet_4_14_0_clk),
    .RESET_B(net106),
    .D(_0068_),
    .Q_N(_0870_),
    .Q(\system_inst.loader.weight_a[2] ));
 sg13g2_dfrbp_1 _1836_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net104),
    .D(_0069_),
    .Q_N(_0869_),
    .Q(\system_inst.leak_rate_1[0] ));
 sg13g2_dfrbp_1 _1837_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net102),
    .D(net195),
    .Q_N(_0021_),
    .Q(\system_inst.leak_rate_1[1] ));
 sg13g2_dfrbp_1 _1838_ (.CLK(clknet_4_6_0_clk),
    .RESET_B(net100),
    .D(net229),
    .Q_N(_0020_),
    .Q(\system_inst.leak_rate_1[2] ));
 sg13g2_dfrbp_1 _1839_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net98),
    .D(net233),
    .Q_N(_0019_),
    .Q(\system_inst.leak_rate_1[3] ));
 sg13g2_dfrbp_1 _1840_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net96),
    .D(_0073_),
    .Q_N(_0018_),
    .Q(\system_inst.leak_rate_1[4] ));
 sg13g2_dfrbp_1 _1841_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net94),
    .D(_0074_),
    .Q_N(_0017_),
    .Q(\system_inst.leak_rate_1[5] ));
 sg13g2_dfrbp_1 _1842_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net92),
    .D(_0075_),
    .Q_N(_0016_),
    .Q(\system_inst.leak_rate_1[6] ));
 sg13g2_dfrbp_1 _1843_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net90),
    .D(net210),
    .Q_N(_0015_),
    .Q(\system_inst.leak_rate_1[7] ));
 sg13g2_dfrbp_1 _1844_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net88),
    .D(_0077_),
    .Q_N(_0868_),
    .Q(\system_inst.leak_rate_2[0] ));
 sg13g2_dfrbp_1 _1845_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net86),
    .D(net243),
    .Q_N(_0028_),
    .Q(\system_inst.leak_rate_2[1] ));
 sg13g2_dfrbp_1 _1846_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net84),
    .D(net206),
    .Q_N(_0027_),
    .Q(\system_inst.leak_rate_2[2] ));
 sg13g2_dfrbp_1 _1847_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net82),
    .D(net249),
    .Q_N(_0026_),
    .Q(\system_inst.leak_rate_2[3] ));
 sg13g2_dfrbp_1 _1848_ (.CLK(clknet_4_2_0_clk),
    .RESET_B(net80),
    .D(_0081_),
    .Q_N(_0025_),
    .Q(\system_inst.leak_rate_2[4] ));
 sg13g2_dfrbp_1 _1849_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net77),
    .D(_0082_),
    .Q_N(_0024_),
    .Q(\system_inst.leak_rate_2[5] ));
 sg13g2_dfrbp_1 _1850_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net73),
    .D(_0083_),
    .Q_N(_0023_),
    .Q(\system_inst.leak_rate_2[6] ));
 sg13g2_dfrbp_1 _1851_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net69),
    .D(net218),
    .Q_N(_0022_),
    .Q(\system_inst.leak_rate_2[7] ));
 sg13g2_dfrbp_1 _1852_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net65),
    .D(_0085_),
    .Q_N(_0038_),
    .Q(\system_inst.loader.threshold_min[0] ));
 sg13g2_dfrbp_1 _1853_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net61),
    .D(_0086_),
    .Q_N(_0867_),
    .Q(\system_inst.loader.threshold_min[1] ));
 sg13g2_dfrbp_1 _1854_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net57),
    .D(_0087_),
    .Q_N(_0036_),
    .Q(\system_inst.loader.threshold_min[2] ));
 sg13g2_dfrbp_1 _1855_ (.CLK(clknet_4_4_0_clk),
    .RESET_B(net53),
    .D(net247),
    .Q_N(_0035_),
    .Q(\system_inst.loader.threshold_min[3] ));
 sg13g2_dfrbp_1 _1856_ (.CLK(clknet_4_1_0_clk),
    .RESET_B(net48),
    .D(_0089_),
    .Q_N(_0033_),
    .Q(\system_inst.loader.threshold_min[4] ));
 sg13g2_dfrbp_1 _1857_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net44),
    .D(_0090_),
    .Q_N(_0032_),
    .Q(\system_inst.loader.threshold_min[5] ));
 sg13g2_dfrbp_1 _1858_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net32),
    .D(_0091_),
    .Q_N(_0031_),
    .Q(\system_inst.loader.threshold_min[6] ));
 sg13g2_dfrbp_1 _1859_ (.CLK(clknet_4_0_0_clk),
    .RESET_B(net105),
    .D(net255),
    .Q_N(_0866_),
    .Q(\system_inst.loader.threshold_min[7] ));
 sg13g2_dfrbp_1 _1860_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net101),
    .D(_0093_),
    .Q_N(_0865_),
    .Q(\system_inst.leak_cycles_1[0] ));
 sg13g2_dfrbp_1 _1861_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net97),
    .D(net129),
    .Q_N(_0864_),
    .Q(\system_inst.leak_cycles_1[1] ));
 sg13g2_dfrbp_1 _1862_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net93),
    .D(net221),
    .Q_N(_0863_),
    .Q(\system_inst.leak_cycles_1[2] ));
 sg13g2_dfrbp_1 _1863_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net89),
    .D(net224),
    .Q_N(_0862_),
    .Q(\system_inst.leak_cycles_1[3] ));
 sg13g2_dfrbp_1 _1864_ (.CLK(clknet_4_10_0_clk),
    .RESET_B(net85),
    .D(_0097_),
    .Q_N(_0861_),
    .Q(\system_inst.leak_cycles_2[0] ));
 sg13g2_dfrbp_1 _1865_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net81),
    .D(net212),
    .Q_N(_0860_),
    .Q(\system_inst.leak_cycles_2[1] ));
 sg13g2_dfrbp_1 _1866_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net75),
    .D(net136),
    .Q_N(_0859_),
    .Q(\system_inst.leak_cycles_2[2] ));
 sg13g2_dfrbp_1 _1867_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net67),
    .D(net142),
    .Q_N(_0858_),
    .Q(\system_inst.leak_cycles_2[3] ));
 sg13g2_dfrbp_1 _1868_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net59),
    .D(_0101_),
    .Q_N(_0857_),
    .Q(\system_inst.loader.shift_reg[0] ));
 sg13g2_dfrbp_1 _1869_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net50),
    .D(_0102_),
    .Q_N(_0856_),
    .Q(\system_inst.loader.shift_reg[1] ));
 sg13g2_dfrbp_1 _1870_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net34),
    .D(net240),
    .Q_N(_0855_),
    .Q(\system_inst.loader.shift_reg[2] ));
 sg13g2_dfrbp_1 _1871_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net103),
    .D(_0104_),
    .Q_N(_0854_),
    .Q(\system_inst.loader.shift_reg[3] ));
 sg13g2_dfrbp_1 _1872_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net95),
    .D(_0105_),
    .Q_N(_0853_),
    .Q(\system_inst.loader.shift_reg[4] ));
 sg13g2_dfrbp_1 _1873_ (.CLK(clknet_4_9_0_clk),
    .RESET_B(net87),
    .D(_0106_),
    .Q_N(_0852_),
    .Q(\system_inst.loader.shift_reg[5] ));
 sg13g2_dfrbp_1 _1874_ (.CLK(clknet_4_3_0_clk),
    .RESET_B(net79),
    .D(net140),
    .Q_N(_0851_),
    .Q(\system_inst.loader.shift_reg[6] ));
 sg13g2_dfrbp_1 _1875_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net63),
    .D(_0108_),
    .Q_N(_0850_),
    .Q(\system_inst.loader.bit_count[0] ));
 sg13g2_dfrbp_1 _1876_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net46),
    .D(net125),
    .Q_N(_0849_),
    .Q(\system_inst.loader.bit_count[1] ));
 sg13g2_dfrbp_1 _1877_ (.CLK(clknet_4_13_0_clk),
    .RESET_B(net99),
    .D(net113),
    .Q_N(_0030_),
    .Q(\system_inst.loader.bit_count[2] ));
 sg13g2_dfrbp_1 _1878_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net83),
    .D(_0111_),
    .Q_N(_0848_),
    .Q(\system_inst.neuron.leak_counter_1[0] ));
 sg13g2_dfrbp_1 _1879_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net55),
    .D(net123),
    .Q_N(_0847_),
    .Q(\system_inst.neuron.leak_counter_1[1] ));
 sg13g2_dfrbp_1 _1880_ (.CLK(clknet_4_11_0_clk),
    .RESET_B(net91),
    .D(_0113_),
    .Q_N(_0846_),
    .Q(\system_inst.neuron.leak_counter_1[2] ));
 sg13g2_dfrbp_1 _1881_ (.CLK(clknet_4_8_0_clk),
    .RESET_B(net107),
    .D(_0114_),
    .Q_N(_0845_),
    .Q(\system_inst.neuron.leak_counter_1[3] ));
 sg13g2_tiehi _1805__26 (.L_HI(net26));
 sg13g2_tiehi _1799__27 (.L_HI(net27));
 sg13g2_tiehi _1800__28 (.L_HI(net28));
 sg13g2_tiehi _1801__29 (.L_HI(net29));
 sg13g2_tiehi _1802__30 (.L_HI(net30));
 sg13g2_tiehi _1803__31 (.L_HI(net31));
 sg13g2_tiehi _1858__32 (.L_HI(net32));
 sg13g2_tiehi _1833__33 (.L_HI(net33));
 sg13g2_tiehi _1870__34 (.L_HI(net34));
 sg13g2_tiehi _1832__35 (.L_HI(net35));
 sg13g2_tiehi _1831__36 (.L_HI(net36));
 sg13g2_tiehi _1830__37 (.L_HI(net37));
 sg13g2_tiehi _1829__38 (.L_HI(net38));
 sg13g2_tiehi _1828__39 (.L_HI(net39));
 sg13g2_tiehi _1827__40 (.L_HI(net40));
 sg13g2_tiehi _1826__41 (.L_HI(net41));
 sg13g2_tiehi _1825__42 (.L_HI(net42));
 sg13g2_tiehi _1824__43 (.L_HI(net43));
 sg13g2_tiehi _1857__44 (.L_HI(net44));
 sg13g2_tiehi _1823__45 (.L_HI(net45));
 sg13g2_tiehi _1876__46 (.L_HI(net46));
 sg13g2_tiehi _1822__47 (.L_HI(net47));
 sg13g2_tiehi _1856__48 (.L_HI(net48));
 sg13g2_tiehi _1821__49 (.L_HI(net49));
 sg13g2_tiehi _1869__50 (.L_HI(net50));
 sg13g2_tiehi _1820__51 (.L_HI(net51));
 sg13g2_tiehi _1819__52 (.L_HI(net52));
 sg13g2_tiehi _1855__53 (.L_HI(net53));
 sg13g2_tiehi _1818__54 (.L_HI(net54));
 sg13g2_tiehi _1879__55 (.L_HI(net55));
 sg13g2_tiehi _1817__56 (.L_HI(net56));
 sg13g2_tiehi _1854__57 (.L_HI(net57));
 sg13g2_tiehi _1816__58 (.L_HI(net58));
 sg13g2_tiehi _1868__59 (.L_HI(net59));
 sg13g2_tiehi _1815__60 (.L_HI(net60));
 sg13g2_tiehi _1853__61 (.L_HI(net61));
 sg13g2_tiehi _1814__62 (.L_HI(net62));
 sg13g2_tiehi _1875__63 (.L_HI(net63));
 sg13g2_tiehi _1813__64 (.L_HI(net64));
 sg13g2_tiehi _1852__65 (.L_HI(net65));
 sg13g2_tiehi _1812__66 (.L_HI(net66));
 sg13g2_tiehi _1867__67 (.L_HI(net67));
 sg13g2_tiehi _1811__68 (.L_HI(net68));
 sg13g2_tiehi _1851__69 (.L_HI(net69));
 sg13g2_tiehi _1810__70 (.L_HI(net70));
 sg13g2_tiehi _1804__71 (.L_HI(net71));
 sg13g2_tiehi _1809__72 (.L_HI(net72));
 sg13g2_tiehi _1850__73 (.L_HI(net73));
 sg13g2_tiehi _1808__74 (.L_HI(net74));
 sg13g2_tiehi _1866__75 (.L_HI(net75));
 sg13g2_tiehi _1807__76 (.L_HI(net76));
 sg13g2_tiehi _1849__77 (.L_HI(net77));
 sg13g2_tiehi _1806__78 (.L_HI(net78));
 sg13g2_tiehi _1874__79 (.L_HI(net79));
 sg13g2_tiehi _1848__80 (.L_HI(net80));
 sg13g2_tiehi _1865__81 (.L_HI(net81));
 sg13g2_tiehi _1847__82 (.L_HI(net82));
 sg13g2_tiehi _1878__83 (.L_HI(net83));
 sg13g2_tiehi _1846__84 (.L_HI(net84));
 sg13g2_tiehi _1864__85 (.L_HI(net85));
 sg13g2_tiehi _1845__86 (.L_HI(net86));
 sg13g2_tiehi _1873__87 (.L_HI(net87));
 sg13g2_tiehi _1844__88 (.L_HI(net88));
 sg13g2_tiehi _1863__89 (.L_HI(net89));
 sg13g2_tiehi _1843__90 (.L_HI(net90));
 sg13g2_tiehi _1880__91 (.L_HI(net91));
 sg13g2_tiehi _1842__92 (.L_HI(net92));
 sg13g2_tiehi _1862__93 (.L_HI(net93));
 sg13g2_tiehi _1841__94 (.L_HI(net94));
 sg13g2_tiehi _1872__95 (.L_HI(net95));
 sg13g2_tiehi _1840__96 (.L_HI(net96));
 sg13g2_tiehi _1861__97 (.L_HI(net97));
 sg13g2_tiehi _1839__98 (.L_HI(net98));
 sg13g2_tiehi _1877__99 (.L_HI(net99));
 sg13g2_tiehi _1838__100 (.L_HI(net100));
 sg13g2_tiehi _1860__101 (.L_HI(net101));
 sg13g2_tiehi _1837__102 (.L_HI(net102));
 sg13g2_tiehi _1871__103 (.L_HI(net103));
 sg13g2_tiehi _1836__104 (.L_HI(net104));
 sg13g2_tiehi _1859__105 (.L_HI(net105));
 sg13g2_tiehi _1835__106 (.L_HI(net106));
 sg13g2_tiehi _1881__107 (.L_HI(net107));
 sg13g2_tiehi tt_um_alif_single_dualleak_108 (.L_HI(net108));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_alif_single_dualleak_12 (.L_LO(net12));
 sg13g2_tielo tt_um_alif_single_dualleak_13 (.L_LO(net13));
 sg13g2_tielo tt_um_alif_single_dualleak_14 (.L_LO(net14));
 sg13g2_tielo tt_um_alif_single_dualleak_15 (.L_LO(net15));
 sg13g2_tielo tt_um_alif_single_dualleak_16 (.L_LO(net16));
 sg13g2_tielo tt_um_alif_single_dualleak_17 (.L_LO(net17));
 sg13g2_tielo tt_um_alif_single_dualleak_18 (.L_LO(net18));
 sg13g2_tielo tt_um_alif_single_dualleak_19 (.L_LO(net19));
 sg13g2_tielo tt_um_alif_single_dualleak_20 (.L_LO(net20));
 sg13g2_tielo tt_um_alif_single_dualleak_21 (.L_LO(net21));
 sg13g2_tielo tt_um_alif_single_dualleak_22 (.L_LO(net22));
 sg13g2_tielo tt_um_alif_single_dualleak_23 (.L_LO(net23));
 sg13g2_tielo tt_um_alif_single_dualleak_24 (.L_LO(net24));
 sg13g2_tiehi _1834__25 (.L_HI(net25));
 sg13g2_buf_2 _1980_ (.A(params_ready),
    .X(uio_out[0]));
 sg13g2_buf_1 _1981_ (.A(spike_out),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout147 (.A(_0732_),
    .X(net147));
 sg13g2_buf_1 fanout148 (.A(_0732_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(net151));
 sg13g2_buf_2 fanout151 (.A(_0632_),
    .X(net151));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(_0567_));
 sg13g2_buf_2 fanout153 (.A(_0567_),
    .X(net153));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(_0724_));
 sg13g2_buf_2 fanout155 (.A(_0724_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_0691_),
    .X(net156));
 sg13g2_buf_1 fanout157 (.A(_0691_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_0838_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_0204_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_0228_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_0228_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_0218_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(net166),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_0194_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_0192_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_0189_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_0186_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_0181_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(net269),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(\system_inst.loader.weight_a[2] ),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(net260),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(\system_inst.neuron.threshold[2] ),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(net266),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_0176_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(net181),
    .X(net179));
 sg13g2_buf_1 fanout180 (.A(net181),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(net183),
    .X(net181));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(net183));
 sg13g2_buf_2 fanout183 (.A(_0172_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(net185),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_4 fanout186 (.X(net186),
    .A(rst_n));
 sg13g2_buf_2 fanout187 (.A(net190),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(net190),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(net190),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(net193),
    .X(net190));
 sg13g2_buf_4 fanout191 (.X(net191),
    .A(net193));
 sg13g2_buf_2 fanout192 (.A(net193),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(rst_n),
    .X(net193));
 sg13g2_buf_2 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_tielo tt_um_alif_single_dualleak_11 (.L_LO(net11));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\system_inst.neuron.v_mem[7] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold2 (.A(\system_inst.neuron.refr_cnt[3] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0056_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold4 (.A(\system_inst.loader.bit_count[2] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0110_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold6 (.A(\system_inst.neuron.v_mem[0] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold7 (.A(\system_inst.neuron.leak_counter_2[1] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0209_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0040_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold10 (.A(\system_inst.loader.current_state[4] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0004_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold12 (.A(\system_inst.loader.bit_count[0] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold13 (.A(\system_inst.neuron.leak_counter_1[1] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0135_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0112_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold16 (.A(\system_inst.loader.bit_count[1] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0109_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold18 (.A(\system_inst.neuron.v_mem[1] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold19 (.A(\system_inst.loader.current_state[2] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold20 (.A(\system_inst.leak_cycles_1[1] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0094_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold22 (.A(\system_inst.loader.current_state[6] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold23 (.A(\system_inst.neuron.v_mem[2] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold24 (.A(\system_inst.loader.current_state[0] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold25 (.A(\system_inst.loader.current_state[3] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0187_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold27 (.A(\system_inst.leak_cycles_2[2] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0099_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold29 (.A(\system_inst.loader.current_state[5] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0191_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold31 (.A(\system_inst.loader.shift_reg[5] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0107_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold33 (.A(\system_inst.leak_cycles_2[3] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0100_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold35 (.A(\system_inst.leak_cycles_1[0] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold36 (.A(\system_inst.neuron.leak_counter_1[2] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0137_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold38 (.A(\system_inst.neuron.v_mem[6] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold39 (.A(\system_inst.leak_rate_1[1] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0070_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold41 (.A(\system_inst.neuron.refr_cnt[1] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0654_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold43 (.A(\system_inst.neuron.v_mem[3] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold44 (.A(\system_inst.leak_cycles_2[0] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold45 (.A(\system_inst.neuron.v_mem[5] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold46 (.A(\system_inst.neuron.v_mem[4] ),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold47 (.A(\system_inst.loader.current_state[1] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold48 (.A(\system_inst.neuron.leak_counter_2[0] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold49 (.A(\system_inst.loader.shift_reg[4] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold50 (.A(\system_inst.leak_rate_2[2] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0079_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold52 (.A(\system_inst.leak_rate_1[6] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold53 (.A(\system_inst.neuron.leak_counter_1[3] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold54 (.A(\system_inst.leak_rate_1[7] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0076_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold56 (.A(\system_inst.leak_cycles_2[1] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0098_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold58 (.A(\system_inst.neuron.leak_counter_2[3] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0212_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold60 (.A(\system_inst.neuron.leak_counter_1[0] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold61 (.A(\system_inst.neuron.leak_counter_2[2] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold62 (.A(\system_inst.leak_rate_2[7] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0084_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold64 (.A(\system_inst.leak_rate_2[6] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold65 (.A(\system_inst.leak_cycles_1[2] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0095_),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold67 (.A(\system_inst.leak_rate_1[5] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold68 (.A(\system_inst.leak_cycles_1[3] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0096_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold70 (.A(\system_inst.loader.threshold_min[6] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold71 (.A(\system_inst.loader.shift_reg[3] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold72 (.A(params_ready),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold73 (.A(\system_inst.leak_rate_1[2] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0071_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold75 (.A(\system_inst.loader.threshold_min[4] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold76 (.A(\system_inst.loader.threshold_min[5] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold77 (.A(\system_inst.leak_rate_1[3] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0072_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold79 (.A(\system_inst.neuron.threshold[0] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0063_),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold81 (.A(\system_inst.leak_rate_2[5] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold82 (.A(\system_inst.leak_rate_2[4] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold83 (.A(\system_inst.leak_rate_1[4] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold84 (.A(\system_inst.loader.shift_reg[1] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0103_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold86 (.A(\system_inst.neuron.refr_cnt[0] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold87 (.A(\system_inst.leak_rate_2[1] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0078_),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold89 (.A(\system_inst.neuron.threshold[6] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0061_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold91 (.A(\system_inst.loader.threshold_min[3] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0088_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold93 (.A(\system_inst.leak_rate_2[3] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0080_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold95 (.A(\system_inst.loader.shift_reg[0] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0067_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold97 (.A(\system_inst.neuron.threshold[4] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold98 (.A(\system_inst.neuron.threshold[5] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold99 (.A(\system_inst.loader.shift_reg[6] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0092_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold101 (.A(\system_inst.loader.threshold_min[0] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold102 (.A(\system_inst.loader.threshold_min[7] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0062_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold104 (.A(\system_inst.leak_rate_1[0] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold105 (.A(\system_inst.loader.weight_a[2] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold106 (.A(\system_inst.neuron.refr_cnt[2] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0656_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold108 (.A(\system_inst.loader.shift_reg[2] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold109 (.A(\system_inst.leak_rate_2[0] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold110 (.A(\system_inst.loader.threshold_min[2] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold111 (.A(\system_inst.neuron.v_mem[8] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold112 (.A(\system_inst.neuron.threshold[1] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold113 (.A(\system_inst.loader.weight_a[0] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold114 (.A(\system_inst.loader.threshold_min[1] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold115 (.A(params_ready),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold116 (.A(params_ready),
    .X(net271));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_fill_2 FILLER_8_336 ();
 sg13g2_fill_1 FILLER_8_368 ();
 sg13g2_fill_1 FILLER_8_373 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_fill_1 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_4 FILLER_9_168 ();
 sg13g2_fill_1 FILLER_9_172 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_4 FILLER_9_231 ();
 sg13g2_fill_1 FILLER_9_235 ();
 sg13g2_decap_8 FILLER_9_262 ();
 sg13g2_decap_8 FILLER_9_269 ();
 sg13g2_decap_8 FILLER_9_276 ();
 sg13g2_decap_4 FILLER_9_283 ();
 sg13g2_fill_1 FILLER_9_287 ();
 sg13g2_fill_1 FILLER_9_314 ();
 sg13g2_fill_2 FILLER_9_360 ();
 sg13g2_fill_2 FILLER_9_370 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_fill_1 FILLER_10_84 ();
 sg13g2_decap_4 FILLER_10_90 ();
 sg13g2_fill_2 FILLER_10_94 ();
 sg13g2_decap_8 FILLER_10_100 ();
 sg13g2_decap_8 FILLER_10_107 ();
 sg13g2_decap_8 FILLER_10_114 ();
 sg13g2_decap_8 FILLER_10_121 ();
 sg13g2_decap_8 FILLER_10_128 ();
 sg13g2_decap_8 FILLER_10_135 ();
 sg13g2_decap_4 FILLER_10_142 ();
 sg13g2_fill_1 FILLER_10_146 ();
 sg13g2_fill_2 FILLER_10_152 ();
 sg13g2_fill_2 FILLER_10_180 ();
 sg13g2_decap_8 FILLER_10_208 ();
 sg13g2_decap_8 FILLER_10_215 ();
 sg13g2_fill_2 FILLER_10_222 ();
 sg13g2_fill_1 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_229 ();
 sg13g2_decap_8 FILLER_10_236 ();
 sg13g2_decap_4 FILLER_10_243 ();
 sg13g2_decap_4 FILLER_10_255 ();
 sg13g2_fill_2 FILLER_10_259 ();
 sg13g2_decap_4 FILLER_10_287 ();
 sg13g2_fill_1 FILLER_10_291 ();
 sg13g2_fill_2 FILLER_10_310 ();
 sg13g2_fill_2 FILLER_10_339 ();
 sg13g2_fill_1 FILLER_10_364 ();
 sg13g2_fill_2 FILLER_10_374 ();
 sg13g2_decap_4 FILLER_10_403 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_fill_2 FILLER_11_77 ();
 sg13g2_fill_1 FILLER_11_79 ();
 sg13g2_decap_4 FILLER_11_111 ();
 sg13g2_fill_1 FILLER_11_115 ();
 sg13g2_decap_4 FILLER_11_142 ();
 sg13g2_fill_2 FILLER_11_170 ();
 sg13g2_fill_1 FILLER_11_181 ();
 sg13g2_fill_2 FILLER_11_240 ();
 sg13g2_fill_1 FILLER_11_242 ();
 sg13g2_fill_1 FILLER_11_247 ();
 sg13g2_fill_2 FILLER_11_261 ();
 sg13g2_decap_8 FILLER_11_293 ();
 sg13g2_fill_1 FILLER_11_300 ();
 sg13g2_decap_8 FILLER_11_337 ();
 sg13g2_fill_2 FILLER_11_344 ();
 sg13g2_fill_1 FILLER_11_346 ();
 sg13g2_fill_1 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_fill_1 FILLER_12_70 ();
 sg13g2_decap_4 FILLER_12_109 ();
 sg13g2_fill_1 FILLER_12_133 ();
 sg13g2_fill_2 FILLER_12_224 ();
 sg13g2_fill_2 FILLER_12_304 ();
 sg13g2_fill_1 FILLER_12_306 ();
 sg13g2_fill_2 FILLER_12_321 ();
 sg13g2_decap_4 FILLER_12_360 ();
 sg13g2_fill_2 FILLER_12_364 ();
 sg13g2_fill_1 FILLER_12_369 ();
 sg13g2_fill_1 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_4 FILLER_13_96 ();
 sg13g2_decap_8 FILLER_13_120 ();
 sg13g2_fill_2 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_4 FILLER_13_168 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_decap_4 FILLER_13_180 ();
 sg13g2_fill_2 FILLER_13_184 ();
 sg13g2_fill_2 FILLER_13_201 ();
 sg13g2_fill_1 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_222 ();
 sg13g2_fill_2 FILLER_13_229 ();
 sg13g2_decap_8 FILLER_13_240 ();
 sg13g2_fill_2 FILLER_13_271 ();
 sg13g2_decap_4 FILLER_13_278 ();
 sg13g2_fill_1 FILLER_13_282 ();
 sg13g2_fill_1 FILLER_13_288 ();
 sg13g2_fill_2 FILLER_13_298 ();
 sg13g2_fill_2 FILLER_13_318 ();
 sg13g2_fill_2 FILLER_13_351 ();
 sg13g2_fill_1 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_decap_4 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_4 FILLER_14_21 ();
 sg13g2_fill_2 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_31 ();
 sg13g2_decap_4 FILLER_14_43 ();
 sg13g2_fill_1 FILLER_14_47 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_fill_2 FILLER_14_81 ();
 sg13g2_decap_4 FILLER_14_92 ();
 sg13g2_fill_2 FILLER_14_96 ();
 sg13g2_fill_2 FILLER_14_108 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_fill_1 FILLER_14_130 ();
 sg13g2_fill_2 FILLER_14_136 ();
 sg13g2_fill_1 FILLER_14_144 ();
 sg13g2_decap_4 FILLER_14_175 ();
 sg13g2_fill_2 FILLER_14_205 ();
 sg13g2_decap_8 FILLER_14_212 ();
 sg13g2_fill_2 FILLER_14_219 ();
 sg13g2_fill_2 FILLER_14_252 ();
 sg13g2_decap_4 FILLER_14_280 ();
 sg13g2_fill_1 FILLER_14_284 ();
 sg13g2_fill_2 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_fill_2 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_decap_4 FILLER_14_346 ();
 sg13g2_fill_2 FILLER_14_350 ();
 sg13g2_decap_4 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_402 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_16 ();
 sg13g2_fill_2 FILLER_15_48 ();
 sg13g2_decap_4 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_125 ();
 sg13g2_decap_4 FILLER_15_134 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_decap_8 FILLER_15_143 ();
 sg13g2_fill_1 FILLER_15_150 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_186 ();
 sg13g2_fill_1 FILLER_15_188 ();
 sg13g2_decap_8 FILLER_15_194 ();
 sg13g2_fill_1 FILLER_15_201 ();
 sg13g2_fill_2 FILLER_15_228 ();
 sg13g2_fill_2 FILLER_15_235 ();
 sg13g2_fill_1 FILLER_15_237 ();
 sg13g2_decap_4 FILLER_15_252 ();
 sg13g2_fill_1 FILLER_15_256 ();
 sg13g2_fill_2 FILLER_15_262 ();
 sg13g2_fill_1 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_289 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_fill_2 FILLER_15_319 ();
 sg13g2_fill_1 FILLER_15_321 ();
 sg13g2_fill_1 FILLER_15_328 ();
 sg13g2_fill_2 FILLER_15_381 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_4 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_15 ();
 sg13g2_decap_8 FILLER_16_22 ();
 sg13g2_decap_8 FILLER_16_29 ();
 sg13g2_fill_2 FILLER_16_36 ();
 sg13g2_fill_2 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_44 ();
 sg13g2_fill_2 FILLER_16_54 ();
 sg13g2_decap_4 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_72 ();
 sg13g2_fill_2 FILLER_16_79 ();
 sg13g2_decap_4 FILLER_16_99 ();
 sg13g2_fill_1 FILLER_16_103 ();
 sg13g2_decap_4 FILLER_16_108 ();
 sg13g2_fill_1 FILLER_16_112 ();
 sg13g2_decap_4 FILLER_16_118 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_decap_4 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_184 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_decap_8 FILLER_16_198 ();
 sg13g2_decap_8 FILLER_16_205 ();
 sg13g2_fill_1 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_230 ();
 sg13g2_fill_2 FILLER_16_240 ();
 sg13g2_fill_1 FILLER_16_242 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_fill_2 FILLER_16_286 ();
 sg13g2_fill_1 FILLER_16_293 ();
 sg13g2_decap_4 FILLER_16_335 ();
 sg13g2_fill_2 FILLER_16_343 ();
 sg13g2_fill_1 FILLER_16_345 ();
 sg13g2_fill_2 FILLER_16_366 ();
 sg13g2_fill_1 FILLER_17_26 ();
 sg13g2_fill_2 FILLER_17_42 ();
 sg13g2_fill_1 FILLER_17_44 ();
 sg13g2_fill_2 FILLER_17_75 ();
 sg13g2_fill_1 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_97 ();
 sg13g2_decap_4 FILLER_17_115 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_decap_4 FILLER_17_194 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_decap_4 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_decap_8 FILLER_17_244 ();
 sg13g2_fill_2 FILLER_17_251 ();
 sg13g2_fill_2 FILLER_17_258 ();
 sg13g2_fill_2 FILLER_17_265 ();
 sg13g2_fill_1 FILLER_17_267 ();
 sg13g2_fill_1 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_309 ();
 sg13g2_decap_4 FILLER_17_316 ();
 sg13g2_fill_2 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_18 ();
 sg13g2_fill_1 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_39 ();
 sg13g2_fill_2 FILLER_18_65 ();
 sg13g2_decap_8 FILLER_18_101 ();
 sg13g2_fill_2 FILLER_18_108 ();
 sg13g2_fill_1 FILLER_18_110 ();
 sg13g2_decap_8 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_132 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_decap_8 FILLER_18_162 ();
 sg13g2_decap_4 FILLER_18_169 ();
 sg13g2_fill_1 FILLER_18_178 ();
 sg13g2_fill_2 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_194 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_fill_1 FILLER_18_205 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_243 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_fill_2 FILLER_18_301 ();
 sg13g2_fill_1 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_317 ();
 sg13g2_fill_1 FILLER_18_359 ();
 sg13g2_fill_2 FILLER_18_395 ();
 sg13g2_fill_2 FILLER_19_43 ();
 sg13g2_fill_2 FILLER_19_54 ();
 sg13g2_fill_1 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_65 ();
 sg13g2_fill_1 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_4 FILLER_19_109 ();
 sg13g2_fill_1 FILLER_19_113 ();
 sg13g2_decap_4 FILLER_19_137 ();
 sg13g2_fill_2 FILLER_19_141 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_4 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_158 ();
 sg13g2_decap_4 FILLER_19_164 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_fill_2 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_183 ();
 sg13g2_decap_4 FILLER_19_193 ();
 sg13g2_fill_1 FILLER_19_197 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_fill_2 FILLER_19_218 ();
 sg13g2_decap_8 FILLER_19_246 ();
 sg13g2_fill_1 FILLER_19_253 ();
 sg13g2_decap_4 FILLER_19_266 ();
 sg13g2_fill_2 FILLER_19_270 ();
 sg13g2_decap_4 FILLER_19_298 ();
 sg13g2_fill_1 FILLER_19_328 ();
 sg13g2_fill_2 FILLER_19_352 ();
 sg13g2_fill_1 FILLER_19_373 ();
 sg13g2_decap_4 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_9 ();
 sg13g2_decap_4 FILLER_20_40 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_4 FILLER_20_76 ();
 sg13g2_fill_2 FILLER_20_80 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_4 FILLER_20_132 ();
 sg13g2_decap_4 FILLER_20_148 ();
 sg13g2_fill_1 FILLER_20_152 ();
 sg13g2_decap_8 FILLER_20_185 ();
 sg13g2_decap_8 FILLER_20_192 ();
 sg13g2_decap_4 FILLER_20_199 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_212 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_decap_8 FILLER_20_229 ();
 sg13g2_decap_8 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_4 FILLER_20_277 ();
 sg13g2_fill_2 FILLER_20_281 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_decap_4 FILLER_20_306 ();
 sg13g2_fill_2 FILLER_20_310 ();
 sg13g2_decap_8 FILLER_20_316 ();
 sg13g2_fill_2 FILLER_20_323 ();
 sg13g2_fill_1 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_26 ();
 sg13g2_fill_2 FILLER_21_61 ();
 sg13g2_fill_1 FILLER_21_63 ();
 sg13g2_fill_1 FILLER_21_69 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_4 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_4 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_109 ();
 sg13g2_fill_1 FILLER_21_120 ();
 sg13g2_fill_1 FILLER_21_126 ();
 sg13g2_fill_2 FILLER_21_135 ();
 sg13g2_fill_1 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_142 ();
 sg13g2_decap_8 FILLER_21_149 ();
 sg13g2_decap_4 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_decap_8 FILLER_21_185 ();
 sg13g2_decap_4 FILLER_21_192 ();
 sg13g2_fill_1 FILLER_21_216 ();
 sg13g2_decap_8 FILLER_21_232 ();
 sg13g2_decap_4 FILLER_21_239 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_decap_4 FILLER_21_265 ();
 sg13g2_fill_1 FILLER_21_274 ();
 sg13g2_fill_1 FILLER_21_280 ();
 sg13g2_fill_2 FILLER_21_289 ();
 sg13g2_fill_1 FILLER_21_291 ();
 sg13g2_fill_2 FILLER_21_318 ();
 sg13g2_fill_1 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_326 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_349 ();
 sg13g2_decap_4 FILLER_21_356 ();
 sg13g2_fill_2 FILLER_21_360 ();
 sg13g2_fill_2 FILLER_21_372 ();
 sg13g2_fill_1 FILLER_21_374 ();
 sg13g2_fill_1 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_28 ();
 sg13g2_fill_2 FILLER_22_36 ();
 sg13g2_decap_8 FILLER_22_43 ();
 sg13g2_decap_8 FILLER_22_58 ();
 sg13g2_decap_4 FILLER_22_65 ();
 sg13g2_fill_2 FILLER_22_69 ();
 sg13g2_decap_4 FILLER_22_89 ();
 sg13g2_fill_1 FILLER_22_93 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_4 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_117 ();
 sg13g2_fill_2 FILLER_22_124 ();
 sg13g2_fill_1 FILLER_22_134 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_fill_2 FILLER_22_147 ();
 sg13g2_fill_1 FILLER_22_149 ();
 sg13g2_decap_8 FILLER_22_160 ();
 sg13g2_decap_8 FILLER_22_185 ();
 sg13g2_decap_4 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_196 ();
 sg13g2_fill_2 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_216 ();
 sg13g2_decap_4 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_227 ();
 sg13g2_decap_8 FILLER_22_241 ();
 sg13g2_fill_2 FILLER_22_256 ();
 sg13g2_decap_4 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_266 ();
 sg13g2_fill_1 FILLER_22_272 ();
 sg13g2_decap_4 FILLER_22_285 ();
 sg13g2_fill_1 FILLER_22_289 ();
 sg13g2_decap_4 FILLER_22_311 ();
 sg13g2_fill_2 FILLER_22_331 ();
 sg13g2_decap_8 FILLER_22_359 ();
 sg13g2_decap_4 FILLER_22_366 ();
 sg13g2_fill_1 FILLER_22_370 ();
 sg13g2_fill_2 FILLER_22_380 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_11 ();
 sg13g2_fill_2 FILLER_23_30 ();
 sg13g2_fill_1 FILLER_23_32 ();
 sg13g2_decap_8 FILLER_23_37 ();
 sg13g2_fill_2 FILLER_23_44 ();
 sg13g2_decap_8 FILLER_23_54 ();
 sg13g2_decap_8 FILLER_23_61 ();
 sg13g2_fill_1 FILLER_23_68 ();
 sg13g2_fill_2 FILLER_23_77 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_decap_4 FILLER_23_106 ();
 sg13g2_decap_4 FILLER_23_121 ();
 sg13g2_decap_4 FILLER_23_141 ();
 sg13g2_fill_2 FILLER_23_145 ();
 sg13g2_fill_2 FILLER_23_166 ();
 sg13g2_fill_1 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_177 ();
 sg13g2_decap_4 FILLER_23_184 ();
 sg13g2_fill_1 FILLER_23_188 ();
 sg13g2_fill_2 FILLER_23_209 ();
 sg13g2_fill_1 FILLER_23_211 ();
 sg13g2_decap_4 FILLER_23_241 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_fill_1 FILLER_23_264 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_289 ();
 sg13g2_fill_2 FILLER_23_296 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_fill_1 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_fill_1 FILLER_23_359 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_17 ();
 sg13g2_fill_2 FILLER_24_24 ();
 sg13g2_fill_1 FILLER_24_26 ();
 sg13g2_fill_1 FILLER_24_37 ();
 sg13g2_fill_1 FILLER_24_43 ();
 sg13g2_fill_1 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_4 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_88 ();
 sg13g2_fill_2 FILLER_24_103 ();
 sg13g2_decap_8 FILLER_24_124 ();
 sg13g2_decap_4 FILLER_24_131 ();
 sg13g2_decap_8 FILLER_24_148 ();
 sg13g2_decap_8 FILLER_24_155 ();
 sg13g2_decap_8 FILLER_24_162 ();
 sg13g2_decap_8 FILLER_24_178 ();
 sg13g2_fill_2 FILLER_24_185 ();
 sg13g2_fill_2 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_204 ();
 sg13g2_decap_4 FILLER_24_230 ();
 sg13g2_fill_1 FILLER_24_234 ();
 sg13g2_decap_4 FILLER_24_247 ();
 sg13g2_fill_1 FILLER_24_251 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_fill_2 FILLER_24_354 ();
 sg13g2_fill_1 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_25_26 ();
 sg13g2_decap_4 FILLER_25_33 ();
 sg13g2_fill_2 FILLER_25_37 ();
 sg13g2_decap_8 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_61 ();
 sg13g2_fill_2 FILLER_25_81 ();
 sg13g2_fill_1 FILLER_25_92 ();
 sg13g2_decap_8 FILLER_25_101 ();
 sg13g2_fill_2 FILLER_25_108 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_decap_4 FILLER_25_127 ();
 sg13g2_fill_2 FILLER_25_131 ();
 sg13g2_fill_1 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_153 ();
 sg13g2_fill_1 FILLER_25_160 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_fill_2 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_183 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_decap_4 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_226 ();
 sg13g2_fill_2 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_fill_2 FILLER_25_249 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_283 ();
 sg13g2_decap_4 FILLER_25_290 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_fill_2 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_310 ();
 sg13g2_fill_1 FILLER_25_320 ();
 sg13g2_decap_4 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_335 ();
 sg13g2_decap_4 FILLER_25_346 ();
 sg13g2_fill_2 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_355 ();
 sg13g2_fill_1 FILLER_25_362 ();
 sg13g2_fill_1 FILLER_25_397 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_16 ();
 sg13g2_fill_1 FILLER_26_18 ();
 sg13g2_decap_4 FILLER_26_31 ();
 sg13g2_fill_1 FILLER_26_35 ();
 sg13g2_fill_1 FILLER_26_53 ();
 sg13g2_fill_2 FILLER_26_68 ();
 sg13g2_decap_8 FILLER_26_78 ();
 sg13g2_fill_1 FILLER_26_85 ();
 sg13g2_fill_2 FILLER_26_91 ();
 sg13g2_decap_4 FILLER_26_100 ();
 sg13g2_fill_2 FILLER_26_104 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_fill_2 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_143 ();
 sg13g2_fill_2 FILLER_26_150 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_184 ();
 sg13g2_fill_2 FILLER_26_191 ();
 sg13g2_fill_1 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_fill_1 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_fill_1 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_256 ();
 sg13g2_fill_2 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_265 ();
 sg13g2_decap_8 FILLER_26_274 ();
 sg13g2_decap_4 FILLER_26_281 ();
 sg13g2_fill_2 FILLER_26_311 ();
 sg13g2_fill_1 FILLER_26_313 ();
 sg13g2_fill_2 FILLER_26_328 ();
 sg13g2_fill_1 FILLER_26_345 ();
 sg13g2_fill_2 FILLER_26_380 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_15 ();
 sg13g2_fill_2 FILLER_27_19 ();
 sg13g2_decap_8 FILLER_27_25 ();
 sg13g2_decap_4 FILLER_27_32 ();
 sg13g2_fill_2 FILLER_27_40 ();
 sg13g2_decap_8 FILLER_27_47 ();
 sg13g2_decap_8 FILLER_27_54 ();
 sg13g2_fill_2 FILLER_27_61 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_decap_4 FILLER_27_69 ();
 sg13g2_fill_2 FILLER_27_73 ();
 sg13g2_fill_2 FILLER_27_80 ();
 sg13g2_decap_8 FILLER_27_108 ();
 sg13g2_fill_1 FILLER_27_115 ();
 sg13g2_decap_8 FILLER_27_124 ();
 sg13g2_decap_4 FILLER_27_131 ();
 sg13g2_decap_8 FILLER_27_150 ();
 sg13g2_decap_8 FILLER_27_157 ();
 sg13g2_decap_8 FILLER_27_170 ();
 sg13g2_fill_2 FILLER_27_177 ();
 sg13g2_fill_1 FILLER_27_179 ();
 sg13g2_decap_8 FILLER_27_184 ();
 sg13g2_fill_2 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_193 ();
 sg13g2_decap_8 FILLER_27_215 ();
 sg13g2_fill_2 FILLER_27_222 ();
 sg13g2_fill_1 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_260 ();
 sg13g2_decap_8 FILLER_27_292 ();
 sg13g2_fill_2 FILLER_27_299 ();
 sg13g2_fill_1 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_decap_8 FILLER_27_312 ();
 sg13g2_fill_1 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_329 ();
 sg13g2_fill_1 FILLER_27_340 ();
 sg13g2_fill_2 FILLER_27_362 ();
 sg13g2_fill_1 FILLER_27_364 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_2 FILLER_28_26 ();
 sg13g2_fill_2 FILLER_28_53 ();
 sg13g2_fill_2 FILLER_28_76 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_94 ();
 sg13g2_decap_4 FILLER_28_101 ();
 sg13g2_fill_1 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_decap_8 FILLER_28_116 ();
 sg13g2_decap_4 FILLER_28_123 ();
 sg13g2_decap_4 FILLER_28_151 ();
 sg13g2_decap_8 FILLER_28_185 ();
 sg13g2_decap_4 FILLER_28_192 ();
 sg13g2_fill_2 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_228 ();
 sg13g2_fill_2 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_decap_8 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_249 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_265 ();
 sg13g2_decap_4 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_289 ();
 sg13g2_fill_2 FILLER_28_362 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_fill_1 FILLER_28_382 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_decap_4 FILLER_29_30 ();
 sg13g2_fill_2 FILLER_29_48 ();
 sg13g2_fill_1 FILLER_29_50 ();
 sg13g2_decap_8 FILLER_29_55 ();
 sg13g2_fill_2 FILLER_29_62 ();
 sg13g2_decap_8 FILLER_29_74 ();
 sg13g2_fill_2 FILLER_29_81 ();
 sg13g2_fill_2 FILLER_29_92 ();
 sg13g2_fill_1 FILLER_29_94 ();
 sg13g2_decap_8 FILLER_29_121 ();
 sg13g2_decap_8 FILLER_29_143 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_165 ();
 sg13g2_decap_4 FILLER_29_171 ();
 sg13g2_fill_1 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_184 ();
 sg13g2_decap_8 FILLER_29_212 ();
 sg13g2_fill_2 FILLER_29_225 ();
 sg13g2_fill_1 FILLER_29_243 ();
 sg13g2_decap_4 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_256 ();
 sg13g2_decap_8 FILLER_29_275 ();
 sg13g2_fill_2 FILLER_29_282 ();
 sg13g2_fill_1 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_295 ();
 sg13g2_decap_8 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_fill_1 FILLER_29_322 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_355 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_24 ();
 sg13g2_fill_1 FILLER_30_26 ();
 sg13g2_decap_8 FILLER_30_37 ();
 sg13g2_fill_2 FILLER_30_44 ();
 sg13g2_fill_1 FILLER_30_46 ();
 sg13g2_decap_8 FILLER_30_65 ();
 sg13g2_decap_8 FILLER_30_72 ();
 sg13g2_fill_2 FILLER_30_79 ();
 sg13g2_fill_1 FILLER_30_81 ();
 sg13g2_decap_4 FILLER_30_98 ();
 sg13g2_fill_1 FILLER_30_102 ();
 sg13g2_decap_4 FILLER_30_108 ();
 sg13g2_decap_8 FILLER_30_115 ();
 sg13g2_decap_4 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_135 ();
 sg13g2_fill_1 FILLER_30_137 ();
 sg13g2_fill_1 FILLER_30_145 ();
 sg13g2_decap_4 FILLER_30_169 ();
 sg13g2_fill_2 FILLER_30_173 ();
 sg13g2_decap_8 FILLER_30_188 ();
 sg13g2_decap_4 FILLER_30_195 ();
 sg13g2_fill_1 FILLER_30_199 ();
 sg13g2_decap_8 FILLER_30_222 ();
 sg13g2_decap_4 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_233 ();
 sg13g2_decap_8 FILLER_30_240 ();
 sg13g2_decap_8 FILLER_30_247 ();
 sg13g2_decap_4 FILLER_30_254 ();
 sg13g2_decap_8 FILLER_30_271 ();
 sg13g2_fill_2 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_310 ();
 sg13g2_decap_4 FILLER_30_317 ();
 sg13g2_fill_2 FILLER_30_324 ();
 sg13g2_fill_1 FILLER_30_326 ();
 sg13g2_fill_2 FILLER_30_345 ();
 sg13g2_decap_4 FILLER_30_371 ();
 sg13g2_decap_4 FILLER_30_384 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_16 ();
 sg13g2_decap_4 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_25 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_4 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_60 ();
 sg13g2_fill_1 FILLER_31_78 ();
 sg13g2_decap_4 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_decap_8 FILLER_31_121 ();
 sg13g2_fill_2 FILLER_31_128 ();
 sg13g2_decap_4 FILLER_31_136 ();
 sg13g2_fill_1 FILLER_31_149 ();
 sg13g2_decap_8 FILLER_31_159 ();
 sg13g2_decap_8 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_201 ();
 sg13g2_decap_8 FILLER_31_208 ();
 sg13g2_decap_4 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_247 ();
 sg13g2_decap_8 FILLER_31_269 ();
 sg13g2_decap_4 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_decap_4 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_fill_2 FILLER_31_318 ();
 sg13g2_fill_1 FILLER_31_320 ();
 sg13g2_decap_4 FILLER_31_347 ();
 sg13g2_fill_1 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_381 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_30 ();
 sg13g2_decap_8 FILLER_32_47 ();
 sg13g2_decap_8 FILLER_32_71 ();
 sg13g2_fill_2 FILLER_32_78 ();
 sg13g2_fill_1 FILLER_32_80 ();
 sg13g2_fill_2 FILLER_32_86 ();
 sg13g2_decap_4 FILLER_32_100 ();
 sg13g2_decap_4 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_113 ();
 sg13g2_decap_4 FILLER_32_117 ();
 sg13g2_decap_4 FILLER_32_125 ();
 sg13g2_decap_4 FILLER_32_137 ();
 sg13g2_decap_4 FILLER_32_145 ();
 sg13g2_fill_2 FILLER_32_149 ();
 sg13g2_decap_4 FILLER_32_168 ();
 sg13g2_fill_1 FILLER_32_172 ();
 sg13g2_fill_2 FILLER_32_178 ();
 sg13g2_decap_4 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_209 ();
 sg13g2_decap_8 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_fill_1 FILLER_32_229 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_4 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_268 ();
 sg13g2_fill_1 FILLER_32_275 ();
 sg13g2_decap_8 FILLER_32_300 ();
 sg13g2_decap_8 FILLER_32_307 ();
 sg13g2_fill_2 FILLER_32_314 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_decap_8 FILLER_32_370 ();
 sg13g2_decap_8 FILLER_32_377 ();
 sg13g2_fill_2 FILLER_32_388 ();
 sg13g2_fill_1 FILLER_32_390 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_9 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_4 FILLER_33_21 ();
 sg13g2_fill_1 FILLER_33_25 ();
 sg13g2_fill_2 FILLER_33_30 ();
 sg13g2_fill_1 FILLER_33_32 ();
 sg13g2_decap_4 FILLER_33_43 ();
 sg13g2_fill_2 FILLER_33_52 ();
 sg13g2_fill_1 FILLER_33_54 ();
 sg13g2_fill_1 FILLER_33_72 ();
 sg13g2_decap_8 FILLER_33_78 ();
 sg13g2_fill_2 FILLER_33_94 ();
 sg13g2_fill_1 FILLER_33_109 ();
 sg13g2_decap_8 FILLER_33_136 ();
 sg13g2_fill_2 FILLER_33_143 ();
 sg13g2_fill_1 FILLER_33_145 ();
 sg13g2_decap_4 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_233 ();
 sg13g2_fill_1 FILLER_33_235 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_253 ();
 sg13g2_decap_4 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_decap_8 FILLER_33_310 ();
 sg13g2_fill_1 FILLER_33_317 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_343 ();
 sg13g2_fill_1 FILLER_33_345 ();
 sg13g2_decap_4 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_33_369 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_fill_2 FILLER_34_35 ();
 sg13g2_decap_4 FILLER_34_41 ();
 sg13g2_fill_2 FILLER_34_45 ();
 sg13g2_fill_1 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_69 ();
 sg13g2_decap_8 FILLER_34_76 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_decap_8 FILLER_34_135 ();
 sg13g2_fill_1 FILLER_34_142 ();
 sg13g2_decap_4 FILLER_34_151 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_decap_8 FILLER_34_197 ();
 sg13g2_decap_8 FILLER_34_220 ();
 sg13g2_decap_4 FILLER_34_227 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_255 ();
 sg13g2_decap_8 FILLER_34_262 ();
 sg13g2_decap_4 FILLER_34_269 ();
 sg13g2_fill_1 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_288 ();
 sg13g2_fill_2 FILLER_34_293 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_decap_8 FILLER_34_305 ();
 sg13g2_decap_4 FILLER_34_312 ();
 sg13g2_fill_1 FILLER_34_316 ();
 sg13g2_fill_1 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_337 ();
 sg13g2_decap_4 FILLER_34_352 ();
 sg13g2_fill_2 FILLER_34_364 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_11 ();
 sg13g2_decap_4 FILLER_35_17 ();
 sg13g2_fill_1 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_94 ();
 sg13g2_fill_1 FILLER_35_117 ();
 sg13g2_fill_2 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_147 ();
 sg13g2_decap_4 FILLER_35_185 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_fill_1 FILLER_35_201 ();
 sg13g2_fill_2 FILLER_35_228 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_fill_1 FILLER_35_246 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_1 FILLER_35_316 ();
 sg13g2_decap_4 FILLER_35_348 ();
 sg13g2_fill_1 FILLER_35_352 ();
 sg13g2_fill_2 FILLER_35_367 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_44 ();
 sg13g2_decap_4 FILLER_36_54 ();
 sg13g2_decap_8 FILLER_36_71 ();
 sg13g2_fill_2 FILLER_36_78 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_99 ();
 sg13g2_fill_1 FILLER_36_128 ();
 sg13g2_fill_1 FILLER_36_138 ();
 sg13g2_decap_8 FILLER_36_153 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_200 ();
 sg13g2_fill_2 FILLER_36_209 ();
 sg13g2_fill_1 FILLER_36_211 ();
 sg13g2_decap_8 FILLER_36_218 ();
 sg13g2_fill_2 FILLER_36_225 ();
 sg13g2_fill_1 FILLER_36_227 ();
 sg13g2_decap_8 FILLER_36_240 ();
 sg13g2_fill_2 FILLER_36_247 ();
 sg13g2_decap_4 FILLER_36_253 ();
 sg13g2_fill_2 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_decap_8 FILLER_36_277 ();
 sg13g2_fill_2 FILLER_36_284 ();
 sg13g2_fill_1 FILLER_36_286 ();
 sg13g2_decap_4 FILLER_36_296 ();
 sg13g2_fill_2 FILLER_36_300 ();
 sg13g2_fill_2 FILLER_36_307 ();
 sg13g2_fill_1 FILLER_36_309 ();
 sg13g2_fill_2 FILLER_36_324 ();
 sg13g2_fill_1 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_36_340 ();
 sg13g2_decap_8 FILLER_36_347 ();
 sg13g2_fill_1 FILLER_36_354 ();
 sg13g2_fill_2 FILLER_36_376 ();
 sg13g2_fill_1 FILLER_36_378 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_fill_1 FILLER_37_71 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_fill_1 FILLER_37_173 ();
 sg13g2_decap_4 FILLER_37_226 ();
 sg13g2_fill_2 FILLER_37_254 ();
 sg13g2_fill_2 FILLER_37_276 ();
 sg13g2_fill_1 FILLER_37_278 ();
 sg13g2_fill_2 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_49 ();
 sg13g2_fill_1 FILLER_38_51 ();
 sg13g2_fill_2 FILLER_38_82 ();
 sg13g2_fill_1 FILLER_38_84 ();
 sg13g2_fill_1 FILLER_38_123 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_179 ();
 sg13g2_fill_2 FILLER_38_183 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_219 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_decap_4 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_4 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_270 ();
 sg13g2_decap_8 FILLER_38_277 ();
 sg13g2_decap_4 FILLER_38_284 ();
 sg13g2_fill_2 FILLER_38_288 ();
 sg13g2_decap_8 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_302 ();
 sg13g2_fill_1 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_332 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_2 FILLER_38_349 ();
 sg13g2_fill_2 FILLER_38_377 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net108;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net12;
 assign uio_oe[3] = net13;
 assign uio_oe[4] = net14;
 assign uio_oe[5] = net15;
 assign uio_oe[6] = net16;
 assign uio_oe[7] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule
