VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_oscillating_bones
  CLASS BLOCK ;
  FOREIGN tt_um_oscillating_bones ;
  ORIGIN 0.000 0.000 ;
  SIZE 202.080 BY 313.740 ;
  PIN ena
    PORT
      LAYER Metal5 ;
        RECT 190.890 312.740 191.190 313.740 ;
    END
  END ena
  PIN clk
    PORT
      LAYER Metal5 ;
        RECT 187.050 312.740 187.350 313.740 ;
    END
  END clk
  PIN rst_n
    PORT
      LAYER Metal5 ;
        RECT 183.210 312.740 183.510 313.740 ;
    END
  END rst_n
  PIN ui_in[0]
    PORT
      LAYER Metal5 ;
        RECT 179.370 312.740 179.670 313.740 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER Metal5 ;
        RECT 175.530 312.740 175.830 313.740 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER Metal5 ;
        RECT 171.690 312.740 171.990 313.740 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER Metal5 ;
        RECT 167.850 312.740 168.150 313.740 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER Metal5 ;
        RECT 164.010 312.740 164.310 313.740 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER Metal5 ;
        RECT 160.170 312.740 160.470 313.740 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER Metal5 ;
        RECT 156.330 312.740 156.630 313.740 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER Metal5 ;
        RECT 152.490 312.740 152.790 313.740 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER Metal5 ;
        RECT 148.650 312.740 148.950 313.740 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER Metal5 ;
        RECT 144.810 312.740 145.110 313.740 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER Metal5 ;
        RECT 140.970 312.740 141.270 313.740 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER Metal5 ;
        RECT 137.130 312.740 137.430 313.740 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER Metal5 ;
        RECT 133.290 312.740 133.590 313.740 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER Metal5 ;
        RECT 129.450 312.740 129.750 313.740 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER Metal5 ;
        RECT 125.610 312.740 125.910 313.740 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER Metal5 ;
        RECT 121.770 312.740 122.070 313.740 ;
    END
  END uio_in[7]
  PIN uo_out[0]
    ANTENNAGATEAREA 3.481800 ;
    ANTENNADIFFAREA 12.700800 ;
    PORT
      LAYER Metal5 ;
        RECT 117.930 312.740 118.230 313.740 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 0.241800 ;
    ANTENNADIFFAREA 0.712400 ;
    PORT
      LAYER Metal5 ;
        RECT 114.090 312.740 114.390 313.740 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNAGATEAREA 0.241800 ;
    ANTENNADIFFAREA 0.712400 ;
    PORT
      LAYER Metal5 ;
        RECT 110.250 312.740 110.550 313.740 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 0.712400 ;
    PORT
      LAYER Metal5 ;
        RECT 106.410 312.740 106.710 313.740 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 102.570 312.740 102.870 313.740 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 98.730 312.740 99.030 313.740 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 94.890 312.740 95.190 313.740 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 91.050 312.740 91.350 313.740 ;
    END
  END uo_out[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 87.210 312.740 87.510 313.740 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 83.370 312.740 83.670 313.740 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 79.530 312.740 79.830 313.740 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 75.690 312.740 75.990 313.740 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 71.850 312.740 72.150 313.740 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 68.010 312.740 68.310 313.740 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 64.170 312.740 64.470 313.740 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 60.330 312.740 60.630 313.740 ;
    END
  END uio_out[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 56.490 312.740 56.790 313.740 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 52.650 312.740 52.950 313.740 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 48.810 312.740 49.110 313.740 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 44.970 312.740 45.270 313.740 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 41.130 312.740 41.430 313.740 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 37.290 312.740 37.590 313.740 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 33.450 312.740 33.750 313.740 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 119.649071 ;
    PORT
      LAYER Metal5 ;
        RECT 29.610 312.740 29.910 313.740 ;
    END
  END uio_oe[7]
  PIN VGND
    ANTENNADIFFAREA 119.649071 ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 5.900 0.000 8.100 310.000 ;
    END
  END VGND
  PIN VDPWR
    ANTENNADIFFAREA 126.628197 ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 9.900 0.000 12.100 310.000 ;
    END
  END VDPWR
  OBS
      LAYER GatPoly ;
        RECT 28.200 59.385 185.850 309.725 ;
      LAYER Metal1 ;
        RECT 28.200 59.385 185.850 309.795 ;
      LAYER Metal2 ;
        RECT 25.480 57.840 187.730 312.715 ;
      LAYER Metal3 ;
        RECT 6.065 51.470 196.625 312.715 ;
      LAYER Metal4 ;
        RECT 6.080 51.470 196.625 312.715 ;
      LAYER Metal5 ;
        RECT 6.550 312.530 29.400 312.875 ;
        RECT 30.120 312.530 33.240 312.875 ;
        RECT 33.960 312.530 37.080 312.875 ;
        RECT 37.800 312.530 40.920 312.875 ;
        RECT 41.640 312.530 44.760 312.875 ;
        RECT 45.480 312.530 48.600 312.875 ;
        RECT 49.320 312.530 52.440 312.875 ;
        RECT 53.160 312.530 56.280 312.875 ;
        RECT 57.000 312.530 60.120 312.875 ;
        RECT 60.840 312.530 63.960 312.875 ;
        RECT 64.680 312.530 67.800 312.875 ;
        RECT 68.520 312.530 71.640 312.875 ;
        RECT 72.360 312.530 75.480 312.875 ;
        RECT 76.200 312.530 79.320 312.875 ;
        RECT 80.040 312.530 83.160 312.875 ;
        RECT 83.880 312.530 87.000 312.875 ;
        RECT 87.720 312.530 90.840 312.875 ;
        RECT 91.560 312.530 94.680 312.875 ;
        RECT 95.400 312.530 98.520 312.875 ;
        RECT 99.240 312.530 102.360 312.875 ;
        RECT 103.080 312.530 106.200 312.875 ;
        RECT 106.920 312.530 110.040 312.875 ;
        RECT 110.760 312.530 113.880 312.875 ;
        RECT 114.600 312.530 117.720 312.875 ;
        RECT 118.440 312.530 121.560 312.875 ;
        RECT 122.280 312.530 125.400 312.875 ;
        RECT 126.120 312.530 129.240 312.875 ;
        RECT 129.960 312.530 133.080 312.875 ;
        RECT 133.800 312.530 136.920 312.875 ;
        RECT 137.640 312.530 140.760 312.875 ;
        RECT 141.480 312.530 144.600 312.875 ;
        RECT 145.320 312.530 148.440 312.875 ;
        RECT 149.160 312.530 152.280 312.875 ;
        RECT 153.000 312.530 156.120 312.875 ;
        RECT 156.840 312.530 159.960 312.875 ;
        RECT 160.680 312.530 163.800 312.875 ;
        RECT 164.520 312.530 167.640 312.875 ;
        RECT 168.360 312.530 171.480 312.875 ;
        RECT 172.200 312.530 175.320 312.875 ;
        RECT 176.040 312.530 179.160 312.875 ;
        RECT 179.880 312.530 183.000 312.875 ;
        RECT 183.720 312.530 186.840 312.875 ;
        RECT 187.560 312.530 190.680 312.875 ;
        RECT 191.400 312.530 196.625 312.875 ;
        RECT 6.550 310.210 196.625 312.530 ;
        RECT 8.310 51.470 9.690 310.210 ;
        RECT 12.310 51.470 196.625 310.210 ;
      LAYER TopMetal1 ;
        RECT 16.625 51.470 196.625 231.470 ;
      LAYER TopMetal2 ;
        RECT 28.300 59.235 185.650 223.905 ;
  END
END tt_um_oscillating_bones
END LIBRARY

